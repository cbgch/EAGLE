//Key = 1011101001110100110100000001000101001110001101010110100111110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376;

XNOR2_X1 U762 ( .A(G107), .B(n1055), .ZN(G9) );
NOR2_X1 U763 ( .A1(n1056), .A2(n1057), .ZN(G75) );
NOR4_X1 U764 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1057) );
XOR2_X1 U765 ( .A(n1062), .B(KEYINPUT28), .Z(n1061) );
NAND2_X1 U766 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U767 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NAND3_X1 U768 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1063) );
NAND2_X1 U769 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NAND2_X1 U770 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND3_X1 U772 ( .A1(n1077), .A2(n1066), .A3(n1078), .ZN(n1076) );
NAND2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1075) );
NAND4_X1 U774 ( .A1(n1081), .A2(n1079), .A3(n1082), .A4(n1066), .ZN(n1071) );
AND2_X1 U775 ( .A1(n1083), .A2(n1067), .ZN(n1060) );
AND3_X1 U776 ( .A1(n1079), .A2(n1073), .A3(n1070), .ZN(n1067) );
NAND3_X1 U777 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1058) );
NAND4_X1 U778 ( .A1(n1070), .A2(n1066), .A3(n1068), .A4(n1087), .ZN(n1086) );
NAND2_X1 U779 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U780 ( .A1(n1073), .A2(n1090), .ZN(n1089) );
NAND2_X1 U781 ( .A1(n1079), .A2(n1091), .ZN(n1088) );
INV_X1 U782 ( .A(n1092), .ZN(n1070) );
NOR3_X1 U783 ( .A1(n1093), .A2(G953), .A3(G952), .ZN(n1056) );
INV_X1 U784 ( .A(n1084), .ZN(n1093) );
NAND4_X1 U785 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1084) );
NOR4_X1 U786 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
XOR2_X1 U787 ( .A(KEYINPUT40), .B(n1102), .Z(n1101) );
XNOR2_X1 U788 ( .A(G478), .B(n1103), .ZN(n1098) );
NOR2_X1 U789 ( .A1(KEYINPUT22), .A2(n1104), .ZN(n1103) );
XNOR2_X1 U790 ( .A(n1105), .B(KEYINPUT56), .ZN(n1104) );
NOR3_X1 U791 ( .A1(n1106), .A2(n1078), .A3(n1107), .ZN(n1096) );
XOR2_X1 U792 ( .A(n1108), .B(n1109), .Z(G72) );
XOR2_X1 U793 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND3_X1 U794 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
NAND2_X1 U795 ( .A1(G953), .A2(n1115), .ZN(n1114) );
NAND2_X1 U796 ( .A1(n1116), .A2(n1117), .ZN(n1113) );
NAND2_X1 U797 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XOR2_X1 U798 ( .A(n1120), .B(n1121), .Z(n1116) );
NAND2_X1 U799 ( .A1(KEYINPUT3), .A2(n1122), .ZN(n1121) );
NAND3_X1 U800 ( .A1(n1118), .A2(n1119), .A3(n1123), .ZN(n1112) );
XOR2_X1 U801 ( .A(n1120), .B(n1124), .Z(n1123) );
NAND2_X1 U802 ( .A1(KEYINPUT3), .A2(n1125), .ZN(n1124) );
INV_X1 U803 ( .A(n1122), .ZN(n1125) );
XOR2_X1 U804 ( .A(n1126), .B(KEYINPUT14), .Z(n1122) );
NAND2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1120) );
NAND2_X1 U806 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XOR2_X1 U807 ( .A(n1131), .B(KEYINPUT12), .Z(n1127) );
OR2_X1 U808 ( .A1(n1130), .A2(n1129), .ZN(n1131) );
XNOR2_X1 U809 ( .A(n1132), .B(n1133), .ZN(n1130) );
XNOR2_X1 U810 ( .A(G131), .B(KEYINPUT7), .ZN(n1132) );
INV_X1 U811 ( .A(KEYINPUT41), .ZN(n1119) );
NAND2_X1 U812 ( .A1(n1085), .A2(n1134), .ZN(n1110) );
NAND2_X1 U813 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U814 ( .A(n1137), .B(KEYINPUT48), .Z(n1135) );
NOR2_X1 U815 ( .A1(n1138), .A2(n1085), .ZN(n1108) );
AND2_X1 U816 ( .A1(G227), .A2(G900), .ZN(n1138) );
XOR2_X1 U817 ( .A(n1139), .B(n1140), .Z(G69) );
NAND2_X1 U818 ( .A1(G953), .A2(n1141), .ZN(n1140) );
NAND2_X1 U819 ( .A1(G898), .A2(G224), .ZN(n1141) );
NAND2_X1 U820 ( .A1(KEYINPUT16), .A2(n1142), .ZN(n1139) );
XOR2_X1 U821 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U822 ( .A1(n1145), .A2(n1085), .ZN(n1144) );
XOR2_X1 U823 ( .A(KEYINPUT19), .B(n1146), .Z(n1145) );
NOR2_X1 U824 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U825 ( .A1(n1149), .A2(n1150), .ZN(n1143) );
NAND2_X1 U826 ( .A1(G953), .A2(n1151), .ZN(n1150) );
XOR2_X1 U827 ( .A(n1152), .B(n1153), .Z(n1149) );
NOR2_X1 U828 ( .A1(n1154), .A2(n1155), .ZN(G66) );
XOR2_X1 U829 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND3_X1 U830 ( .A1(n1158), .A2(G217), .A3(KEYINPUT62), .ZN(n1156) );
NOR2_X1 U831 ( .A1(n1154), .A2(n1159), .ZN(G63) );
NOR3_X1 U832 ( .A1(n1105), .A2(n1160), .A3(n1161), .ZN(n1159) );
AND3_X1 U833 ( .A1(n1162), .A2(G478), .A3(n1158), .ZN(n1161) );
NOR2_X1 U834 ( .A1(n1163), .A2(n1162), .ZN(n1160) );
AND2_X1 U835 ( .A1(n1059), .A2(G478), .ZN(n1163) );
NOR2_X1 U836 ( .A1(n1154), .A2(n1164), .ZN(G60) );
XOR2_X1 U837 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U838 ( .A(KEYINPUT33), .B(n1167), .Z(n1166) );
NOR2_X1 U839 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XNOR2_X1 U840 ( .A(G104), .B(n1170), .ZN(G6) );
NAND3_X1 U841 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1170) );
XOR2_X1 U842 ( .A(KEYINPUT23), .B(n1066), .Z(n1172) );
NOR2_X1 U843 ( .A1(n1154), .A2(n1174), .ZN(G57) );
NOR2_X1 U844 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XOR2_X1 U845 ( .A(n1177), .B(KEYINPUT42), .Z(n1176) );
NAND2_X1 U846 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NOR2_X1 U847 ( .A1(n1178), .A2(n1179), .ZN(n1175) );
XNOR2_X1 U848 ( .A(n1180), .B(n1181), .ZN(n1179) );
XOR2_X1 U849 ( .A(n1129), .B(n1182), .Z(n1181) );
XOR2_X1 U850 ( .A(n1183), .B(n1184), .Z(n1180) );
AND2_X1 U851 ( .A1(G472), .A2(n1158), .ZN(n1184) );
NAND2_X1 U852 ( .A1(KEYINPUT47), .A2(n1185), .ZN(n1183) );
XOR2_X1 U853 ( .A(n1186), .B(n1187), .Z(n1178) );
NAND2_X1 U854 ( .A1(KEYINPUT10), .A2(n1188), .ZN(n1186) );
NAND2_X1 U855 ( .A1(n1189), .A2(G210), .ZN(n1188) );
NOR2_X1 U856 ( .A1(n1154), .A2(n1190), .ZN(G54) );
XOR2_X1 U857 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U858 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U859 ( .A(n1195), .B(n1185), .Z(n1194) );
NOR2_X1 U860 ( .A1(KEYINPUT51), .A2(n1196), .ZN(n1195) );
AND2_X1 U861 ( .A1(G469), .A2(n1158), .ZN(n1193) );
INV_X1 U862 ( .A(n1169), .ZN(n1158) );
XOR2_X1 U863 ( .A(n1197), .B(n1198), .Z(n1191) );
NOR3_X1 U864 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1198) );
NOR2_X1 U865 ( .A1(KEYINPUT25), .A2(n1202), .ZN(n1201) );
NOR2_X1 U866 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
AND3_X1 U867 ( .A1(KEYINPUT37), .A2(n1205), .A3(G140), .ZN(n1204) );
NOR2_X1 U868 ( .A1(KEYINPUT37), .A2(G140), .ZN(n1203) );
NOR2_X1 U869 ( .A1(n1206), .A2(n1207), .ZN(n1200) );
INV_X1 U870 ( .A(KEYINPUT25), .ZN(n1207) );
NOR2_X1 U871 ( .A1(G110), .A2(n1208), .ZN(n1206) );
XOR2_X1 U872 ( .A(KEYINPUT37), .B(G140), .Z(n1208) );
INV_X1 U873 ( .A(n1209), .ZN(n1199) );
NAND3_X1 U874 ( .A1(G227), .A2(n1085), .A3(KEYINPUT6), .ZN(n1197) );
NOR2_X1 U875 ( .A1(n1154), .A2(n1210), .ZN(G51) );
XOR2_X1 U876 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U877 ( .A(KEYINPUT31), .B(n1213), .Z(n1212) );
NOR2_X1 U878 ( .A1(n1214), .A2(n1169), .ZN(n1213) );
NAND2_X1 U879 ( .A1(G902), .A2(n1059), .ZN(n1169) );
NAND4_X1 U880 ( .A1(n1215), .A2(n1136), .A3(n1216), .A4(n1137), .ZN(n1059) );
OR2_X1 U881 ( .A1(n1217), .A2(n1100), .ZN(n1137) );
INV_X1 U882 ( .A(n1148), .ZN(n1216) );
NAND3_X1 U883 ( .A1(n1218), .A2(n1055), .A3(n1219), .ZN(n1148) );
NAND2_X1 U884 ( .A1(n1171), .A2(n1083), .ZN(n1219) );
NAND2_X1 U885 ( .A1(n1220), .A2(n1221), .ZN(n1083) );
NAND2_X1 U886 ( .A1(n1173), .A2(n1066), .ZN(n1221) );
NAND2_X1 U887 ( .A1(n1222), .A2(n1068), .ZN(n1220) );
NAND3_X1 U888 ( .A1(n1065), .A2(n1066), .A3(n1171), .ZN(n1055) );
AND4_X1 U889 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1136) );
AND4_X1 U890 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1226) );
NAND3_X1 U891 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1225) );
INV_X1 U892 ( .A(n1234), .ZN(n1233) );
XOR2_X1 U893 ( .A(KEYINPUT29), .B(n1090), .Z(n1231) );
XOR2_X1 U894 ( .A(n1147), .B(KEYINPUT4), .Z(n1215) );
NAND4_X1 U895 ( .A1(n1235), .A2(n1236), .A3(n1237), .A4(n1238), .ZN(n1147) );
XOR2_X1 U896 ( .A(n1239), .B(n1240), .Z(n1211) );
NOR2_X1 U897 ( .A1(n1085), .A2(G952), .ZN(n1154) );
XNOR2_X1 U898 ( .A(G146), .B(n1223), .ZN(G48) );
NAND4_X1 U899 ( .A1(n1241), .A2(n1242), .A3(n1173), .A4(n1091), .ZN(n1223) );
XOR2_X1 U900 ( .A(n1224), .B(n1243), .Z(G45) );
XOR2_X1 U901 ( .A(KEYINPUT2), .B(G143), .Z(n1243) );
NAND3_X1 U902 ( .A1(n1244), .A2(n1091), .A3(n1245), .ZN(n1224) );
XOR2_X1 U903 ( .A(n1126), .B(n1246), .Z(G42) );
NAND3_X1 U904 ( .A1(KEYINPUT9), .A2(n1073), .A3(n1247), .ZN(n1246) );
XOR2_X1 U905 ( .A(n1217), .B(KEYINPUT52), .Z(n1247) );
NAND3_X1 U906 ( .A1(n1173), .A2(n1080), .A3(n1242), .ZN(n1217) );
XNOR2_X1 U907 ( .A(G137), .B(n1230), .ZN(G39) );
NAND4_X1 U908 ( .A1(n1241), .A2(n1242), .A3(n1073), .A4(n1068), .ZN(n1230) );
XOR2_X1 U909 ( .A(n1248), .B(n1229), .Z(G36) );
NAND3_X1 U910 ( .A1(n1073), .A2(n1065), .A3(n1244), .ZN(n1229) );
XNOR2_X1 U911 ( .A(G131), .B(n1228), .ZN(G33) );
NAND3_X1 U912 ( .A1(n1173), .A2(n1073), .A3(n1244), .ZN(n1228) );
AND2_X1 U913 ( .A1(n1222), .A2(n1242), .ZN(n1244) );
INV_X1 U914 ( .A(n1249), .ZN(n1242) );
INV_X1 U915 ( .A(n1100), .ZN(n1073) );
NAND2_X1 U916 ( .A1(n1082), .A2(n1250), .ZN(n1100) );
XOR2_X1 U917 ( .A(G128), .B(n1251), .Z(G30) );
NOR2_X1 U918 ( .A1(n1249), .A2(n1234), .ZN(n1251) );
NAND3_X1 U919 ( .A1(n1065), .A2(n1091), .A3(n1241), .ZN(n1234) );
NAND2_X1 U920 ( .A1(n1090), .A2(n1232), .ZN(n1249) );
XOR2_X1 U921 ( .A(n1187), .B(n1252), .Z(G3) );
NOR2_X1 U922 ( .A1(n1253), .A2(KEYINPUT60), .ZN(n1252) );
AND3_X1 U923 ( .A1(n1222), .A2(n1068), .A3(n1171), .ZN(n1253) );
XOR2_X1 U924 ( .A(n1118), .B(n1227), .Z(G27) );
NAND4_X1 U925 ( .A1(n1173), .A2(n1079), .A3(n1254), .A4(n1080), .ZN(n1227) );
AND2_X1 U926 ( .A1(n1232), .A2(n1091), .ZN(n1254) );
NAND2_X1 U927 ( .A1(n1092), .A2(n1255), .ZN(n1232) );
NAND4_X1 U928 ( .A1(G953), .A2(G902), .A3(n1256), .A4(n1115), .ZN(n1255) );
INV_X1 U929 ( .A(G900), .ZN(n1115) );
INV_X1 U930 ( .A(G125), .ZN(n1118) );
XOR2_X1 U931 ( .A(n1257), .B(n1235), .Z(G24) );
NAND3_X1 U932 ( .A1(n1245), .A2(n1066), .A3(n1258), .ZN(n1235) );
NOR2_X1 U933 ( .A1(n1259), .A2(n1099), .ZN(n1066) );
AND2_X1 U934 ( .A1(n1260), .A2(n1261), .ZN(n1245) );
XOR2_X1 U935 ( .A(n1262), .B(KEYINPUT54), .Z(n1260) );
XNOR2_X1 U936 ( .A(G119), .B(n1236), .ZN(G21) );
NAND3_X1 U937 ( .A1(n1241), .A2(n1068), .A3(n1258), .ZN(n1236) );
AND2_X1 U938 ( .A1(n1263), .A2(n1099), .ZN(n1241) );
INV_X1 U939 ( .A(n1264), .ZN(n1099) );
XOR2_X1 U940 ( .A(KEYINPUT61), .B(n1265), .Z(n1263) );
XOR2_X1 U941 ( .A(n1237), .B(n1266), .Z(G18) );
XOR2_X1 U942 ( .A(n1267), .B(KEYINPUT39), .Z(n1266) );
NAND3_X1 U943 ( .A1(n1222), .A2(n1065), .A3(n1258), .ZN(n1237) );
XNOR2_X1 U944 ( .A(G113), .B(n1238), .ZN(G15) );
NAND3_X1 U945 ( .A1(n1222), .A2(n1173), .A3(n1258), .ZN(n1238) );
AND3_X1 U946 ( .A1(n1091), .A2(n1268), .A3(n1079), .ZN(n1258) );
NOR2_X1 U947 ( .A1(n1102), .A2(n1078), .ZN(n1079) );
INV_X1 U948 ( .A(n1077), .ZN(n1102) );
AND2_X1 U949 ( .A1(n1269), .A2(n1262), .ZN(n1173) );
NOR2_X1 U950 ( .A1(n1259), .A2(n1264), .ZN(n1222) );
XOR2_X1 U951 ( .A(n1205), .B(n1218), .Z(G12) );
NAND3_X1 U952 ( .A1(n1171), .A2(n1068), .A3(n1080), .ZN(n1218) );
AND2_X1 U953 ( .A1(n1264), .A2(n1265), .ZN(n1080) );
XNOR2_X1 U954 ( .A(n1259), .B(KEYINPUT38), .ZN(n1265) );
NAND2_X1 U955 ( .A1(n1270), .A2(n1094), .ZN(n1259) );
NAND2_X1 U956 ( .A1(G217), .A2(n1271), .ZN(n1094) );
NAND2_X1 U957 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
OR2_X1 U958 ( .A1(n1274), .A2(G234), .ZN(n1273) );
XNOR2_X1 U959 ( .A(n1107), .B(KEYINPUT30), .ZN(n1270) );
AND3_X1 U960 ( .A1(n1275), .A2(n1272), .A3(n1274), .ZN(n1107) );
XOR2_X1 U961 ( .A(n1157), .B(KEYINPUT24), .Z(n1274) );
XNOR2_X1 U962 ( .A(n1276), .B(n1277), .ZN(n1157) );
XOR2_X1 U963 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U964 ( .A(G119), .B(G110), .Z(n1279) );
XOR2_X1 U965 ( .A(KEYINPUT15), .B(G140), .Z(n1278) );
XOR2_X1 U966 ( .A(n1280), .B(n1281), .Z(n1276) );
XOR2_X1 U967 ( .A(n1282), .B(n1283), .Z(n1280) );
NOR2_X1 U968 ( .A1(G125), .A2(KEYINPUT44), .ZN(n1283) );
NAND2_X1 U969 ( .A1(n1284), .A2(n1285), .ZN(n1282) );
NAND4_X1 U970 ( .A1(G137), .A2(G221), .A3(G234), .A4(n1085), .ZN(n1285) );
NAND2_X1 U971 ( .A1(n1286), .A2(n1287), .ZN(n1284) );
NAND3_X1 U972 ( .A1(G234), .A2(n1085), .A3(G221), .ZN(n1287) );
XOR2_X1 U973 ( .A(KEYINPUT0), .B(G137), .Z(n1286) );
NAND2_X1 U974 ( .A1(G217), .A2(n1288), .ZN(n1275) );
INV_X1 U975 ( .A(G234), .ZN(n1288) );
XOR2_X1 U976 ( .A(n1289), .B(G472), .Z(n1264) );
NAND2_X1 U977 ( .A1(n1290), .A2(n1272), .ZN(n1289) );
NAND2_X1 U978 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
OR2_X1 U979 ( .A1(n1293), .A2(KEYINPUT57), .ZN(n1292) );
XOR2_X1 U980 ( .A(n1294), .B(n1295), .Z(n1291) );
XOR2_X1 U981 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U982 ( .A(n1298), .B(KEYINPUT8), .Z(n1297) );
NAND2_X1 U983 ( .A1(KEYINPUT57), .A2(n1293), .ZN(n1296) );
XNOR2_X1 U984 ( .A(n1187), .B(n1299), .ZN(n1293) );
AND3_X1 U985 ( .A1(n1189), .A2(n1300), .A3(G210), .ZN(n1299) );
INV_X1 U986 ( .A(KEYINPUT1), .ZN(n1300) );
XOR2_X1 U987 ( .A(n1182), .B(n1240), .Z(n1294) );
XOR2_X1 U988 ( .A(n1301), .B(KEYINPUT55), .Z(n1182) );
NAND2_X1 U989 ( .A1(n1302), .A2(n1303), .ZN(n1068) );
OR3_X1 U990 ( .A1(n1262), .A2(n1261), .A3(KEYINPUT20), .ZN(n1303) );
NAND2_X1 U991 ( .A1(KEYINPUT20), .A2(n1065), .ZN(n1302) );
NOR2_X1 U992 ( .A1(n1262), .A2(n1269), .ZN(n1065) );
INV_X1 U993 ( .A(n1261), .ZN(n1269) );
XOR2_X1 U994 ( .A(n1105), .B(G478), .Z(n1261) );
NOR2_X1 U995 ( .A1(n1162), .A2(G902), .ZN(n1105) );
XNOR2_X1 U996 ( .A(n1304), .B(n1305), .ZN(n1162) );
XOR2_X1 U997 ( .A(G128), .B(n1306), .Z(n1305) );
XOR2_X1 U998 ( .A(KEYINPUT63), .B(G143), .Z(n1306) );
XOR2_X1 U999 ( .A(n1307), .B(n1308), .Z(n1304) );
AND3_X1 U1000 ( .A1(G217), .A2(n1085), .A3(G234), .ZN(n1308) );
XNOR2_X1 U1001 ( .A(n1309), .B(n1310), .ZN(n1307) );
NAND2_X1 U1002 ( .A1(KEYINPUT49), .A2(n1248), .ZN(n1310) );
INV_X1 U1003 ( .A(G134), .ZN(n1248) );
NAND2_X1 U1004 ( .A1(n1311), .A2(KEYINPUT59), .ZN(n1309) );
XOR2_X1 U1005 ( .A(n1312), .B(G107), .Z(n1311) );
NAND3_X1 U1006 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1312) );
NAND2_X1 U1007 ( .A1(KEYINPUT53), .A2(G122), .ZN(n1315) );
NAND3_X1 U1008 ( .A1(n1257), .A2(n1316), .A3(G116), .ZN(n1314) );
NAND2_X1 U1009 ( .A1(n1317), .A2(n1267), .ZN(n1313) );
INV_X1 U1010 ( .A(G116), .ZN(n1267) );
NAND2_X1 U1011 ( .A1(n1318), .A2(n1316), .ZN(n1317) );
INV_X1 U1012 ( .A(KEYINPUT53), .ZN(n1316) );
XOR2_X1 U1013 ( .A(KEYINPUT13), .B(G122), .Z(n1318) );
NAND2_X1 U1014 ( .A1(n1319), .A2(n1095), .ZN(n1262) );
NAND3_X1 U1015 ( .A1(n1168), .A2(n1272), .A3(n1165), .ZN(n1095) );
INV_X1 U1016 ( .A(G475), .ZN(n1168) );
XNOR2_X1 U1017 ( .A(n1106), .B(KEYINPUT21), .ZN(n1319) );
AND2_X1 U1018 ( .A1(G475), .A2(n1320), .ZN(n1106) );
NAND2_X1 U1019 ( .A1(n1165), .A2(n1272), .ZN(n1320) );
XNOR2_X1 U1020 ( .A(n1321), .B(n1322), .ZN(n1165) );
XOR2_X1 U1021 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1022 ( .A(G113), .B(G104), .Z(n1324) );
XOR2_X1 U1023 ( .A(G125), .B(G122), .Z(n1323) );
XNOR2_X1 U1024 ( .A(n1325), .B(n1326), .ZN(n1321) );
XNOR2_X1 U1025 ( .A(n1327), .B(n1328), .ZN(n1326) );
NOR2_X1 U1026 ( .A1(G140), .A2(KEYINPUT18), .ZN(n1328) );
NAND2_X1 U1027 ( .A1(KEYINPUT58), .A2(n1329), .ZN(n1327) );
XOR2_X1 U1028 ( .A(n1330), .B(n1331), .Z(n1329) );
XOR2_X1 U1029 ( .A(G131), .B(n1332), .Z(n1331) );
NAND2_X1 U1030 ( .A1(n1189), .A2(G214), .ZN(n1330) );
NOR2_X1 U1031 ( .A1(G953), .A2(G237), .ZN(n1189) );
AND3_X1 U1032 ( .A1(n1091), .A2(n1268), .A3(n1090), .ZN(n1171) );
NOR2_X1 U1033 ( .A1(n1077), .A2(n1078), .ZN(n1090) );
AND2_X1 U1034 ( .A1(G221), .A2(n1333), .ZN(n1078) );
NAND2_X1 U1035 ( .A1(G234), .A2(n1272), .ZN(n1333) );
XNOR2_X1 U1036 ( .A(G469), .B(n1334), .ZN(n1077) );
NOR2_X1 U1037 ( .A1(G902), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1038 ( .A(n1336), .B(n1337), .Z(n1335) );
NAND2_X1 U1039 ( .A1(n1338), .A2(KEYINPUT36), .ZN(n1337) );
XOR2_X1 U1040 ( .A(n1339), .B(n1340), .Z(n1338) );
NOR2_X1 U1041 ( .A1(G227), .A2(KEYINPUT34), .ZN(n1340) );
NAND3_X1 U1042 ( .A1(n1341), .A2(n1342), .A3(n1209), .ZN(n1339) );
NAND2_X1 U1043 ( .A1(G110), .A2(n1126), .ZN(n1209) );
INV_X1 U1044 ( .A(G140), .ZN(n1126) );
OR2_X1 U1045 ( .A1(G140), .A2(KEYINPUT50), .ZN(n1342) );
NAND3_X1 U1046 ( .A1(G140), .A2(n1205), .A3(KEYINPUT50), .ZN(n1341) );
NAND2_X1 U1047 ( .A1(n1343), .A2(n1344), .ZN(n1336) );
NAND2_X1 U1048 ( .A1(n1185), .A2(n1196), .ZN(n1344) );
XOR2_X1 U1049 ( .A(n1345), .B(KEYINPUT5), .Z(n1343) );
OR2_X1 U1050 ( .A1(n1196), .A2(n1185), .ZN(n1345) );
INV_X1 U1051 ( .A(n1298), .ZN(n1185) );
NAND2_X1 U1052 ( .A1(n1346), .A2(n1347), .ZN(n1298) );
NAND2_X1 U1053 ( .A1(G131), .A2(n1133), .ZN(n1347) );
XOR2_X1 U1054 ( .A(n1348), .B(KEYINPUT26), .Z(n1346) );
OR2_X1 U1055 ( .A1(n1133), .A2(G131), .ZN(n1348) );
XOR2_X1 U1056 ( .A(G134), .B(G137), .Z(n1133) );
XNOR2_X1 U1057 ( .A(n1349), .B(n1240), .ZN(n1196) );
NAND2_X1 U1058 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
NAND2_X1 U1059 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
NAND2_X1 U1060 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NAND2_X1 U1061 ( .A1(G101), .A2(n1356), .ZN(n1355) );
INV_X1 U1062 ( .A(KEYINPUT32), .ZN(n1354) );
NAND2_X1 U1063 ( .A1(n1357), .A2(n1187), .ZN(n1350) );
INV_X1 U1064 ( .A(G101), .ZN(n1187) );
NAND2_X1 U1065 ( .A1(n1356), .A2(n1358), .ZN(n1357) );
OR2_X1 U1066 ( .A1(n1352), .A2(KEYINPUT32), .ZN(n1358) );
XOR2_X1 U1067 ( .A(n1359), .B(G107), .Z(n1352) );
NAND2_X1 U1068 ( .A1(KEYINPUT11), .A2(G104), .ZN(n1359) );
INV_X1 U1069 ( .A(KEYINPUT46), .ZN(n1356) );
NAND2_X1 U1070 ( .A1(n1092), .A2(n1360), .ZN(n1268) );
NAND4_X1 U1071 ( .A1(G953), .A2(G902), .A3(n1256), .A4(n1151), .ZN(n1360) );
INV_X1 U1072 ( .A(G898), .ZN(n1151) );
NAND3_X1 U1073 ( .A1(n1256), .A2(n1085), .A3(G952), .ZN(n1092) );
NAND2_X1 U1074 ( .A1(G237), .A2(G234), .ZN(n1256) );
NOR2_X1 U1075 ( .A1(n1082), .A2(n1081), .ZN(n1091) );
INV_X1 U1076 ( .A(n1250), .ZN(n1081) );
NAND2_X1 U1077 ( .A1(G214), .A2(n1361), .ZN(n1250) );
XNOR2_X1 U1078 ( .A(n1362), .B(n1214), .ZN(n1082) );
NAND2_X1 U1079 ( .A1(G210), .A2(n1361), .ZN(n1214) );
NAND2_X1 U1080 ( .A1(n1363), .A2(n1272), .ZN(n1361) );
INV_X1 U1081 ( .A(G237), .ZN(n1363) );
NAND3_X1 U1082 ( .A1(n1364), .A2(n1365), .A3(n1272), .ZN(n1362) );
INV_X1 U1083 ( .A(G902), .ZN(n1272) );
NAND2_X1 U1084 ( .A1(n1366), .A2(n1129), .ZN(n1365) );
NAND2_X1 U1085 ( .A1(n1367), .A2(n1240), .ZN(n1364) );
INV_X1 U1086 ( .A(n1129), .ZN(n1240) );
XOR2_X1 U1087 ( .A(n1332), .B(n1281), .Z(n1129) );
XOR2_X1 U1088 ( .A(G128), .B(n1325), .Z(n1281) );
XOR2_X1 U1089 ( .A(G146), .B(KEYINPUT17), .Z(n1325) );
INV_X1 U1090 ( .A(G143), .ZN(n1332) );
XOR2_X1 U1091 ( .A(KEYINPUT45), .B(n1366), .Z(n1367) );
INV_X1 U1092 ( .A(n1239), .ZN(n1366) );
XOR2_X1 U1093 ( .A(n1368), .B(n1369), .Z(n1239) );
XNOR2_X1 U1094 ( .A(n1370), .B(n1153), .ZN(n1369) );
XOR2_X1 U1095 ( .A(n1205), .B(n1257), .Z(n1153) );
INV_X1 U1096 ( .A(G122), .ZN(n1257) );
NAND2_X1 U1097 ( .A1(KEYINPUT27), .A2(n1152), .ZN(n1370) );
XOR2_X1 U1098 ( .A(n1371), .B(n1372), .Z(n1152) );
XOR2_X1 U1099 ( .A(G104), .B(n1373), .Z(n1372) );
XOR2_X1 U1100 ( .A(KEYINPUT35), .B(G107), .Z(n1373) );
XOR2_X1 U1101 ( .A(n1301), .B(G101), .Z(n1371) );
XNOR2_X1 U1102 ( .A(G113), .B(n1374), .ZN(n1301) );
XOR2_X1 U1103 ( .A(G119), .B(G116), .Z(n1374) );
XOR2_X1 U1104 ( .A(n1375), .B(n1376), .Z(n1368) );
XOR2_X1 U1105 ( .A(KEYINPUT43), .B(G125), .Z(n1376) );
NAND2_X1 U1106 ( .A1(G224), .A2(n1085), .ZN(n1375) );
INV_X1 U1107 ( .A(G953), .ZN(n1085) );
INV_X1 U1108 ( .A(G110), .ZN(n1205) );
endmodule


