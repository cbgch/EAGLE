//Key = 0101100001000100000010010000111100001000101010110000111000000011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426;

XOR2_X1 U778 ( .A(G107), .B(n1077), .Z(G9) );
AND2_X1 U779 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U780 ( .A1(n1080), .A2(n1081), .ZN(G75) );
NOR3_X1 U781 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NOR2_X1 U782 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NOR3_X1 U783 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1085) );
NAND3_X1 U784 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1087) );
NAND3_X1 U785 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1082) );
NAND2_X1 U786 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U787 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND3_X1 U788 ( .A1(n1091), .A2(n1100), .A3(n1101), .ZN(n1099) );
NAND2_X1 U789 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NAND2_X1 U790 ( .A1(n1092), .A2(n1104), .ZN(n1103) );
NAND2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U792 ( .A1(n1090), .A2(n1086), .ZN(n1106) );
INV_X1 U793 ( .A(KEYINPUT48), .ZN(n1086) );
INV_X1 U794 ( .A(n1107), .ZN(n1105) );
NAND2_X1 U795 ( .A1(n1108), .A2(n1109), .ZN(n1102) );
NAND2_X1 U796 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND3_X1 U798 ( .A1(n1108), .A2(n1114), .A3(n1092), .ZN(n1098) );
NAND2_X1 U799 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U800 ( .A1(n1101), .A2(n1117), .ZN(n1116) );
NAND2_X1 U801 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
OR2_X1 U802 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U803 ( .A1(n1091), .A2(n1122), .ZN(n1115) );
OR2_X1 U804 ( .A1(n1123), .A2(n1079), .ZN(n1122) );
INV_X1 U805 ( .A(n1089), .ZN(n1096) );
NOR3_X1 U806 ( .A1(n1124), .A2(G953), .A3(G952), .ZN(n1080) );
INV_X1 U807 ( .A(n1093), .ZN(n1124) );
NAND4_X1 U808 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1093) );
NOR4_X1 U809 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1128) );
XOR2_X1 U810 ( .A(G475), .B(n1133), .Z(n1132) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(n1131) );
NOR2_X1 U812 ( .A1(KEYINPUT59), .A2(n1136), .ZN(n1135) );
NOR2_X1 U813 ( .A1(n1137), .A2(n1112), .ZN(n1127) );
XNOR2_X1 U814 ( .A(n1138), .B(n1139), .ZN(n1126) );
NOR2_X1 U815 ( .A1(G469), .A2(KEYINPUT24), .ZN(n1139) );
XOR2_X1 U816 ( .A(n1140), .B(n1141), .Z(n1125) );
XNOR2_X1 U817 ( .A(G472), .B(n1142), .ZN(n1141) );
XOR2_X1 U818 ( .A(KEYINPUT45), .B(KEYINPUT31), .Z(n1140) );
XOR2_X1 U819 ( .A(n1143), .B(n1144), .Z(G72) );
NOR2_X1 U820 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XNOR2_X1 U821 ( .A(G953), .B(KEYINPUT18), .ZN(n1146) );
AND2_X1 U822 ( .A1(G227), .A2(G900), .ZN(n1145) );
NAND2_X1 U823 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
NAND2_X1 U824 ( .A1(n1149), .A2(n1094), .ZN(n1148) );
XNOR2_X1 U825 ( .A(n1150), .B(n1151), .ZN(n1149) );
NOR2_X1 U826 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U827 ( .A(n1154), .B(KEYINPUT39), .Z(n1152) );
NAND3_X1 U828 ( .A1(G900), .A2(n1150), .A3(G953), .ZN(n1147) );
XNOR2_X1 U829 ( .A(n1155), .B(n1156), .ZN(n1150) );
XNOR2_X1 U830 ( .A(n1157), .B(n1158), .ZN(n1156) );
XOR2_X1 U831 ( .A(n1159), .B(n1160), .Z(n1155) );
XNOR2_X1 U832 ( .A(G137), .B(KEYINPUT26), .ZN(n1159) );
XOR2_X1 U833 ( .A(n1161), .B(n1162), .Z(G69) );
XOR2_X1 U834 ( .A(n1163), .B(n1164), .Z(n1162) );
NAND2_X1 U835 ( .A1(G953), .A2(n1165), .ZN(n1164) );
NAND2_X1 U836 ( .A1(G898), .A2(G224), .ZN(n1165) );
NAND2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(n1163) );
NAND2_X1 U838 ( .A1(G953), .A2(n1168), .ZN(n1167) );
XOR2_X1 U839 ( .A(n1169), .B(n1170), .Z(n1166) );
XOR2_X1 U840 ( .A(n1171), .B(n1172), .Z(n1170) );
XNOR2_X1 U841 ( .A(KEYINPUT12), .B(n1173), .ZN(n1169) );
AND2_X1 U842 ( .A1(n1174), .A2(n1094), .ZN(n1161) );
NOR2_X1 U843 ( .A1(n1175), .A2(n1176), .ZN(G66) );
NOR3_X1 U844 ( .A1(n1134), .A2(n1177), .A3(n1178), .ZN(n1176) );
AND3_X1 U845 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1178) );
INV_X1 U846 ( .A(n1136), .ZN(n1180) );
NOR2_X1 U847 ( .A1(n1182), .A2(n1179), .ZN(n1177) );
NOR2_X1 U848 ( .A1(n1183), .A2(n1136), .ZN(n1182) );
NOR2_X1 U849 ( .A1(n1175), .A2(n1184), .ZN(G63) );
XNOR2_X1 U850 ( .A(n1185), .B(n1186), .ZN(n1184) );
XOR2_X1 U851 ( .A(KEYINPUT34), .B(n1187), .Z(n1186) );
AND2_X1 U852 ( .A1(G478), .A2(n1181), .ZN(n1187) );
NOR2_X1 U853 ( .A1(n1175), .A2(n1188), .ZN(G60) );
NOR3_X1 U854 ( .A1(n1133), .A2(n1189), .A3(n1190), .ZN(n1188) );
AND3_X1 U855 ( .A1(n1191), .A2(G475), .A3(n1181), .ZN(n1190) );
NOR2_X1 U856 ( .A1(n1192), .A2(n1191), .ZN(n1189) );
AND2_X1 U857 ( .A1(n1084), .A2(G475), .ZN(n1192) );
INV_X1 U858 ( .A(n1183), .ZN(n1084) );
XNOR2_X1 U859 ( .A(n1193), .B(n1194), .ZN(G6) );
NAND2_X1 U860 ( .A1(KEYINPUT28), .A2(n1195), .ZN(n1193) );
XNOR2_X1 U861 ( .A(KEYINPUT9), .B(n1196), .ZN(n1195) );
NOR2_X1 U862 ( .A1(n1175), .A2(n1197), .ZN(G57) );
XOR2_X1 U863 ( .A(n1198), .B(n1199), .Z(n1197) );
XNOR2_X1 U864 ( .A(n1200), .B(n1201), .ZN(n1199) );
AND2_X1 U865 ( .A1(G472), .A2(n1181), .ZN(n1201) );
NOR2_X1 U866 ( .A1(n1175), .A2(n1202), .ZN(G54) );
NOR2_X1 U867 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
XOR2_X1 U868 ( .A(n1205), .B(n1206), .Z(n1204) );
NOR2_X1 U869 ( .A1(KEYINPUT5), .A2(n1207), .ZN(n1206) );
AND2_X1 U870 ( .A1(G469), .A2(n1181), .ZN(n1205) );
AND2_X1 U871 ( .A1(n1207), .A2(KEYINPUT5), .ZN(n1203) );
NOR2_X1 U872 ( .A1(n1175), .A2(n1208), .ZN(G51) );
XOR2_X1 U873 ( .A(n1209), .B(n1210), .Z(n1208) );
XNOR2_X1 U874 ( .A(n1211), .B(n1212), .ZN(n1210) );
NAND3_X1 U875 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1209) );
NAND2_X1 U876 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND3_X1 U877 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1214) );
INV_X1 U878 ( .A(n1217), .ZN(n1218) );
NAND2_X1 U879 ( .A1(n1221), .A2(G125), .ZN(n1213) );
XNOR2_X1 U880 ( .A(n1217), .B(n1219), .ZN(n1221) );
NAND2_X1 U881 ( .A1(n1181), .A2(n1222), .ZN(n1217) );
NOR2_X1 U882 ( .A1(n1223), .A2(n1183), .ZN(n1181) );
NOR3_X1 U883 ( .A1(n1154), .A2(n1174), .A3(n1153), .ZN(n1183) );
NAND4_X1 U884 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1153) );
NAND3_X1 U885 ( .A1(n1228), .A2(n1123), .A3(n1229), .ZN(n1224) );
NAND4_X1 U886 ( .A1(n1194), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1174) );
AND4_X1 U887 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1232) );
NOR3_X1 U888 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1231) );
NOR3_X1 U889 ( .A1(n1240), .A2(n1241), .A3(n1110), .ZN(n1239) );
NOR4_X1 U890 ( .A1(n1242), .A2(n1118), .A3(n1243), .A4(n1244), .ZN(n1241) );
INV_X1 U891 ( .A(KEYINPUT60), .ZN(n1240) );
NOR4_X1 U892 ( .A1(KEYINPUT60), .A2(n1243), .A3(n1245), .A4(n1244), .ZN(n1238) );
XNOR2_X1 U893 ( .A(n1088), .B(KEYINPUT3), .ZN(n1244) );
NOR4_X1 U894 ( .A1(n1246), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1237) );
INV_X1 U895 ( .A(n1079), .ZN(n1249) );
NOR2_X1 U896 ( .A1(n1250), .A2(n1251), .ZN(n1247) );
INV_X1 U897 ( .A(KEYINPUT7), .ZN(n1251) );
NOR3_X1 U898 ( .A1(n1118), .A2(n1242), .A3(n1252), .ZN(n1250) );
NOR2_X1 U899 ( .A1(KEYINPUT7), .A2(n1253), .ZN(n1246) );
NAND2_X1 U900 ( .A1(n1123), .A2(n1078), .ZN(n1194) );
NOR2_X1 U901 ( .A1(n1245), .A2(n1248), .ZN(n1078) );
INV_X1 U902 ( .A(n1108), .ZN(n1248) );
NAND3_X1 U903 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1154) );
NAND2_X1 U904 ( .A1(n1092), .A2(n1257), .ZN(n1256) );
NAND2_X1 U905 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XOR2_X1 U906 ( .A(KEYINPUT47), .B(n1260), .Z(n1258) );
NOR2_X1 U907 ( .A1(n1094), .A2(G952), .ZN(n1175) );
XNOR2_X1 U908 ( .A(G146), .B(n1261), .ZN(G48) );
NAND3_X1 U909 ( .A1(n1123), .A2(n1262), .A3(n1229), .ZN(n1261) );
XOR2_X1 U910 ( .A(KEYINPUT0), .B(n1228), .Z(n1262) );
XNOR2_X1 U911 ( .A(G143), .B(n1225), .ZN(G45) );
NAND4_X1 U912 ( .A1(n1107), .A2(n1229), .A3(n1263), .A4(n1130), .ZN(n1225) );
XNOR2_X1 U913 ( .A(n1264), .B(n1265), .ZN(G42) );
NAND2_X1 U914 ( .A1(KEYINPUT63), .A2(n1227), .ZN(n1264) );
NAND4_X1 U915 ( .A1(n1123), .A2(n1266), .A3(n1092), .A4(n1090), .ZN(n1227) );
XNOR2_X1 U916 ( .A(G137), .B(n1226), .ZN(G39) );
NAND4_X1 U917 ( .A1(n1101), .A2(n1228), .A3(n1266), .A4(n1092), .ZN(n1226) );
XNOR2_X1 U918 ( .A(n1267), .B(n1268), .ZN(G36) );
NOR2_X1 U919 ( .A1(n1269), .A2(n1259), .ZN(n1268) );
NAND3_X1 U920 ( .A1(n1266), .A2(n1079), .A3(n1107), .ZN(n1259) );
XNOR2_X1 U921 ( .A(n1092), .B(KEYINPUT22), .ZN(n1269) );
NAND2_X1 U922 ( .A1(n1270), .A2(n1271), .ZN(G33) );
NAND3_X1 U923 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n1271) );
INV_X1 U924 ( .A(G131), .ZN(n1274) );
NAND2_X1 U925 ( .A1(G131), .A2(n1275), .ZN(n1270) );
NAND2_X1 U926 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND2_X1 U927 ( .A1(KEYINPUT10), .A2(n1272), .ZN(n1277) );
NAND2_X1 U928 ( .A1(n1278), .A2(n1279), .ZN(n1276) );
INV_X1 U929 ( .A(KEYINPUT10), .ZN(n1279) );
NAND2_X1 U930 ( .A1(n1272), .A2(n1273), .ZN(n1278) );
INV_X1 U931 ( .A(KEYINPUT35), .ZN(n1273) );
AND2_X1 U932 ( .A1(n1092), .A2(n1280), .ZN(n1272) );
XOR2_X1 U933 ( .A(KEYINPUT6), .B(n1260), .Z(n1280) );
AND3_X1 U934 ( .A1(n1123), .A2(n1266), .A3(n1107), .ZN(n1260) );
AND2_X1 U935 ( .A1(n1113), .A2(n1281), .ZN(n1092) );
XNOR2_X1 U936 ( .A(G128), .B(n1254), .ZN(G30) );
NAND3_X1 U937 ( .A1(n1228), .A2(n1079), .A3(n1229), .ZN(n1254) );
AND2_X1 U938 ( .A1(n1266), .A2(n1252), .ZN(n1229) );
NOR2_X1 U939 ( .A1(n1118), .A2(n1282), .ZN(n1266) );
XNOR2_X1 U940 ( .A(G101), .B(n1230), .ZN(G3) );
NAND2_X1 U941 ( .A1(n1283), .A2(n1107), .ZN(n1230) );
XNOR2_X1 U942 ( .A(G125), .B(n1255), .ZN(G27) );
NAND3_X1 U943 ( .A1(n1123), .A2(n1090), .A3(n1284), .ZN(n1255) );
NOR3_X1 U944 ( .A1(n1110), .A2(n1282), .A3(n1285), .ZN(n1284) );
AND2_X1 U945 ( .A1(n1089), .A2(n1286), .ZN(n1282) );
NAND4_X1 U946 ( .A1(G953), .A2(G902), .A3(n1287), .A4(n1288), .ZN(n1286) );
INV_X1 U947 ( .A(G900), .ZN(n1288) );
XNOR2_X1 U948 ( .A(G122), .B(n1236), .ZN(G24) );
NAND4_X1 U949 ( .A1(n1263), .A2(n1289), .A3(n1108), .A4(n1130), .ZN(n1236) );
NOR2_X1 U950 ( .A1(n1290), .A2(n1291), .ZN(n1108) );
NAND2_X1 U951 ( .A1(n1292), .A2(n1293), .ZN(G21) );
NAND2_X1 U952 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
XNOR2_X1 U953 ( .A(KEYINPUT58), .B(n1235), .ZN(n1294) );
NAND2_X1 U954 ( .A1(n1296), .A2(G119), .ZN(n1292) );
XOR2_X1 U955 ( .A(n1235), .B(KEYINPUT25), .Z(n1296) );
NAND3_X1 U956 ( .A1(n1101), .A2(n1228), .A3(n1289), .ZN(n1235) );
AND2_X1 U957 ( .A1(n1291), .A2(n1290), .ZN(n1228) );
INV_X1 U958 ( .A(n1297), .ZN(n1291) );
XNOR2_X1 U959 ( .A(G116), .B(n1234), .ZN(G18) );
NAND3_X1 U960 ( .A1(n1107), .A2(n1079), .A3(n1289), .ZN(n1234) );
NOR2_X1 U961 ( .A1(n1263), .A2(n1298), .ZN(n1079) );
INV_X1 U962 ( .A(n1130), .ZN(n1298) );
XOR2_X1 U963 ( .A(n1233), .B(n1299), .Z(G15) );
NOR2_X1 U964 ( .A1(G113), .A2(KEYINPUT55), .ZN(n1299) );
NAND3_X1 U965 ( .A1(n1107), .A2(n1123), .A3(n1289), .ZN(n1233) );
NOR3_X1 U966 ( .A1(n1285), .A2(n1242), .A3(n1110), .ZN(n1289) );
NOR2_X1 U967 ( .A1(n1300), .A2(n1130), .ZN(n1123) );
NOR2_X1 U968 ( .A1(n1297), .A2(n1290), .ZN(n1107) );
XOR2_X1 U969 ( .A(n1301), .B(n1302), .Z(G12) );
AND2_X1 U970 ( .A1(n1090), .A2(n1283), .ZN(n1302) );
NOR2_X1 U971 ( .A1(n1088), .A2(n1245), .ZN(n1283) );
INV_X1 U972 ( .A(n1253), .ZN(n1245) );
NOR3_X1 U973 ( .A1(n1118), .A2(n1242), .A3(n1110), .ZN(n1253) );
INV_X1 U974 ( .A(n1252), .ZN(n1110) );
NOR2_X1 U975 ( .A1(n1113), .A2(n1112), .ZN(n1252) );
INV_X1 U976 ( .A(n1281), .ZN(n1112) );
NAND2_X1 U977 ( .A1(G214), .A2(n1303), .ZN(n1281) );
XOR2_X1 U978 ( .A(n1129), .B(n1304), .Z(n1113) );
XOR2_X1 U979 ( .A(KEYINPUT44), .B(KEYINPUT41), .Z(n1304) );
XNOR2_X1 U980 ( .A(n1305), .B(n1222), .ZN(n1129) );
AND2_X1 U981 ( .A1(G210), .A2(n1303), .ZN(n1222) );
NAND2_X1 U982 ( .A1(n1306), .A2(n1223), .ZN(n1303) );
NAND2_X1 U983 ( .A1(n1307), .A2(n1223), .ZN(n1305) );
XOR2_X1 U984 ( .A(n1211), .B(n1308), .Z(n1307) );
NOR2_X1 U985 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XOR2_X1 U986 ( .A(KEYINPUT32), .B(n1311), .Z(n1310) );
NOR3_X1 U987 ( .A1(n1212), .A2(n1216), .A3(n1312), .ZN(n1311) );
NOR2_X1 U988 ( .A1(n1313), .A2(n1314), .ZN(n1309) );
INV_X1 U989 ( .A(n1212), .ZN(n1314) );
NAND2_X1 U990 ( .A1(G224), .A2(n1094), .ZN(n1212) );
NOR2_X1 U991 ( .A1(n1216), .A2(n1312), .ZN(n1313) );
NAND2_X1 U992 ( .A1(n1315), .A2(n1316), .ZN(n1312) );
OR2_X1 U993 ( .A1(G125), .A2(KEYINPUT62), .ZN(n1316) );
NAND3_X1 U994 ( .A1(G125), .A2(n1219), .A3(KEYINPUT62), .ZN(n1315) );
NOR2_X1 U995 ( .A1(n1219), .A2(G125), .ZN(n1216) );
XOR2_X1 U996 ( .A(n1317), .B(n1318), .Z(n1219) );
NAND3_X1 U997 ( .A1(n1319), .A2(n1320), .A3(n1321), .ZN(n1211) );
NAND2_X1 U998 ( .A1(KEYINPUT21), .A2(n1322), .ZN(n1321) );
NAND3_X1 U999 ( .A1(n1323), .A2(n1324), .A3(n1325), .ZN(n1320) );
INV_X1 U1000 ( .A(KEYINPUT21), .ZN(n1324) );
OR2_X1 U1001 ( .A1(n1325), .A2(n1323), .ZN(n1319) );
NOR2_X1 U1002 ( .A1(KEYINPUT43), .A2(n1322), .ZN(n1323) );
XNOR2_X1 U1003 ( .A(n1173), .B(G122), .ZN(n1322) );
XNOR2_X1 U1004 ( .A(n1326), .B(n1171), .ZN(n1325) );
XNOR2_X1 U1005 ( .A(n1327), .B(n1328), .ZN(n1171) );
XNOR2_X1 U1006 ( .A(G101), .B(n1329), .ZN(n1328) );
NAND2_X1 U1007 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
XOR2_X1 U1008 ( .A(n1332), .B(KEYINPUT11), .Z(n1330) );
NAND2_X1 U1009 ( .A1(n1333), .A2(G119), .ZN(n1332) );
XNOR2_X1 U1010 ( .A(G116), .B(KEYINPUT2), .ZN(n1333) );
NAND2_X1 U1011 ( .A1(n1334), .A2(n1335), .ZN(n1327) );
XNOR2_X1 U1012 ( .A(KEYINPUT4), .B(KEYINPUT36), .ZN(n1334) );
XNOR2_X1 U1013 ( .A(G113), .B(KEYINPUT14), .ZN(n1326) );
AND2_X1 U1014 ( .A1(n1336), .A2(n1089), .ZN(n1242) );
NAND3_X1 U1015 ( .A1(n1287), .A2(n1094), .A3(G952), .ZN(n1089) );
NAND4_X1 U1016 ( .A1(G953), .A2(G902), .A3(n1287), .A4(n1168), .ZN(n1336) );
INV_X1 U1017 ( .A(G898), .ZN(n1168) );
NAND2_X1 U1018 ( .A1(G237), .A2(G234), .ZN(n1287) );
AND2_X1 U1019 ( .A1(n1337), .A2(n1338), .ZN(n1118) );
OR2_X1 U1020 ( .A1(n1285), .A2(KEYINPUT40), .ZN(n1338) );
INV_X1 U1021 ( .A(n1091), .ZN(n1285) );
NOR2_X1 U1022 ( .A1(n1121), .A2(n1137), .ZN(n1091) );
INV_X1 U1023 ( .A(n1120), .ZN(n1137) );
NAND3_X1 U1024 ( .A1(n1121), .A2(n1120), .A3(KEYINPUT40), .ZN(n1337) );
NAND2_X1 U1025 ( .A1(G221), .A2(n1339), .ZN(n1120) );
XNOR2_X1 U1026 ( .A(n1138), .B(G469), .ZN(n1121) );
NAND3_X1 U1027 ( .A1(n1340), .A2(n1341), .A3(n1223), .ZN(n1138) );
NAND2_X1 U1028 ( .A1(n1207), .A2(n1342), .ZN(n1341) );
INV_X1 U1029 ( .A(KEYINPUT15), .ZN(n1342) );
XOR2_X1 U1030 ( .A(n1343), .B(n1344), .Z(n1207) );
NAND3_X1 U1031 ( .A1(n1344), .A2(n1343), .A3(KEYINPUT15), .ZN(n1340) );
XOR2_X1 U1032 ( .A(n1345), .B(n1346), .Z(n1343) );
XNOR2_X1 U1033 ( .A(n1265), .B(G110), .ZN(n1346) );
NAND2_X1 U1034 ( .A1(G227), .A2(n1094), .ZN(n1345) );
XNOR2_X1 U1035 ( .A(n1347), .B(n1348), .ZN(n1344) );
XOR2_X1 U1036 ( .A(n1349), .B(n1350), .Z(n1348) );
XNOR2_X1 U1037 ( .A(KEYINPUT51), .B(n1200), .ZN(n1350) );
XOR2_X1 U1038 ( .A(n1157), .B(n1335), .Z(n1347) );
XNOR2_X1 U1039 ( .A(n1196), .B(G107), .ZN(n1335) );
INV_X1 U1040 ( .A(G104), .ZN(n1196) );
XNOR2_X1 U1041 ( .A(KEYINPUT1), .B(n1351), .ZN(n1157) );
NOR2_X1 U1042 ( .A1(KEYINPUT8), .A2(n1318), .ZN(n1351) );
INV_X1 U1043 ( .A(n1101), .ZN(n1088) );
NOR2_X1 U1044 ( .A1(n1130), .A2(n1263), .ZN(n1101) );
INV_X1 U1045 ( .A(n1300), .ZN(n1263) );
XOR2_X1 U1046 ( .A(n1133), .B(n1352), .Z(n1300) );
NOR2_X1 U1047 ( .A1(G475), .A2(KEYINPUT38), .ZN(n1352) );
NOR2_X1 U1048 ( .A1(n1191), .A2(G902), .ZN(n1133) );
XOR2_X1 U1049 ( .A(n1353), .B(n1354), .Z(n1191) );
XOR2_X1 U1050 ( .A(n1355), .B(n1356), .Z(n1354) );
XNOR2_X1 U1051 ( .A(n1357), .B(G131), .ZN(n1356) );
XOR2_X1 U1052 ( .A(KEYINPUT56), .B(G146), .Z(n1355) );
XOR2_X1 U1053 ( .A(n1358), .B(n1158), .Z(n1353) );
XOR2_X1 U1054 ( .A(G140), .B(G125), .Z(n1158) );
XOR2_X1 U1055 ( .A(n1359), .B(n1360), .Z(n1358) );
NOR2_X1 U1056 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
INV_X1 U1057 ( .A(G214), .ZN(n1362) );
NAND3_X1 U1058 ( .A1(n1363), .A2(n1364), .A3(n1365), .ZN(n1359) );
NAND2_X1 U1059 ( .A1(KEYINPUT50), .A2(G104), .ZN(n1365) );
OR3_X1 U1060 ( .A1(G104), .A2(KEYINPUT50), .A3(n1172), .ZN(n1364) );
NAND2_X1 U1061 ( .A1(n1172), .A2(n1366), .ZN(n1363) );
NAND2_X1 U1062 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
INV_X1 U1063 ( .A(KEYINPUT50), .ZN(n1368) );
XNOR2_X1 U1064 ( .A(G104), .B(KEYINPUT17), .ZN(n1367) );
XOR2_X1 U1065 ( .A(G113), .B(G122), .Z(n1172) );
XNOR2_X1 U1066 ( .A(n1369), .B(G478), .ZN(n1130) );
NAND2_X1 U1067 ( .A1(n1185), .A2(n1223), .ZN(n1369) );
XNOR2_X1 U1068 ( .A(n1370), .B(n1371), .ZN(n1185) );
NOR2_X1 U1069 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
INV_X1 U1070 ( .A(G217), .ZN(n1373) );
XOR2_X1 U1071 ( .A(n1374), .B(n1375), .Z(n1370) );
NOR2_X1 U1072 ( .A1(KEYINPUT37), .A2(n1376), .ZN(n1375) );
XOR2_X1 U1073 ( .A(n1377), .B(n1378), .Z(n1376) );
XNOR2_X1 U1074 ( .A(n1379), .B(n1380), .ZN(n1378) );
INV_X1 U1075 ( .A(G128), .ZN(n1380) );
NAND2_X1 U1076 ( .A1(KEYINPUT53), .A2(n1357), .ZN(n1379) );
NAND2_X1 U1077 ( .A1(KEYINPUT30), .A2(n1267), .ZN(n1377) );
INV_X1 U1078 ( .A(G134), .ZN(n1267) );
NAND3_X1 U1079 ( .A1(n1381), .A2(n1382), .A3(n1383), .ZN(n1374) );
NAND2_X1 U1080 ( .A1(KEYINPUT27), .A2(n1384), .ZN(n1383) );
NAND3_X1 U1081 ( .A1(G107), .A2(n1385), .A3(n1386), .ZN(n1382) );
INV_X1 U1082 ( .A(KEYINPUT27), .ZN(n1385) );
OR2_X1 U1083 ( .A1(n1386), .A2(G107), .ZN(n1381) );
NOR2_X1 U1084 ( .A1(n1387), .A2(n1384), .ZN(n1386) );
XNOR2_X1 U1085 ( .A(G122), .B(n1388), .ZN(n1384) );
INV_X1 U1086 ( .A(KEYINPUT42), .ZN(n1387) );
INV_X1 U1087 ( .A(n1243), .ZN(n1090) );
NAND2_X1 U1088 ( .A1(n1297), .A2(n1290), .ZN(n1243) );
XNOR2_X1 U1089 ( .A(n1134), .B(n1136), .ZN(n1290) );
NAND2_X1 U1090 ( .A1(G217), .A2(n1339), .ZN(n1136) );
NAND2_X1 U1091 ( .A1(G234), .A2(n1223), .ZN(n1339) );
NOR2_X1 U1092 ( .A1(n1179), .A2(G902), .ZN(n1134) );
XNOR2_X1 U1093 ( .A(n1389), .B(n1390), .ZN(n1179) );
XOR2_X1 U1094 ( .A(n1391), .B(n1392), .Z(n1390) );
XNOR2_X1 U1095 ( .A(G110), .B(G119), .ZN(n1392) );
NAND3_X1 U1096 ( .A1(n1393), .A2(n1394), .A3(n1395), .ZN(n1391) );
NAND2_X1 U1097 ( .A1(G125), .A2(n1265), .ZN(n1395) );
INV_X1 U1098 ( .A(G140), .ZN(n1265) );
NAND2_X1 U1099 ( .A1(n1396), .A2(n1397), .ZN(n1394) );
INV_X1 U1100 ( .A(KEYINPUT23), .ZN(n1397) );
NAND2_X1 U1101 ( .A1(n1398), .A2(n1220), .ZN(n1396) );
XNOR2_X1 U1102 ( .A(KEYINPUT13), .B(G140), .ZN(n1398) );
NAND2_X1 U1103 ( .A1(KEYINPUT23), .A2(n1399), .ZN(n1393) );
NAND2_X1 U1104 ( .A1(n1400), .A2(n1401), .ZN(n1399) );
OR2_X1 U1105 ( .A1(G140), .A2(KEYINPUT13), .ZN(n1401) );
NAND3_X1 U1106 ( .A1(G140), .A2(n1220), .A3(KEYINPUT13), .ZN(n1400) );
INV_X1 U1107 ( .A(G125), .ZN(n1220) );
XNOR2_X1 U1108 ( .A(n1402), .B(n1403), .ZN(n1389) );
NAND2_X1 U1109 ( .A1(KEYINPUT20), .A2(n1404), .ZN(n1402) );
XNOR2_X1 U1110 ( .A(n1405), .B(n1406), .ZN(n1404) );
NOR2_X1 U1111 ( .A1(n1372), .A2(n1407), .ZN(n1406) );
INV_X1 U1112 ( .A(G221), .ZN(n1407) );
NAND2_X1 U1113 ( .A1(n1408), .A2(n1094), .ZN(n1372) );
XOR2_X1 U1114 ( .A(KEYINPUT33), .B(G234), .Z(n1408) );
INV_X1 U1115 ( .A(G137), .ZN(n1405) );
XNOR2_X1 U1116 ( .A(n1142), .B(n1409), .ZN(n1297) );
NOR2_X1 U1117 ( .A1(G472), .A2(n1410), .ZN(n1409) );
XNOR2_X1 U1118 ( .A(KEYINPUT57), .B(KEYINPUT29), .ZN(n1410) );
NAND2_X1 U1119 ( .A1(n1411), .A2(n1223), .ZN(n1142) );
INV_X1 U1120 ( .A(G902), .ZN(n1223) );
XOR2_X1 U1121 ( .A(n1412), .B(n1198), .Z(n1411) );
XNOR2_X1 U1122 ( .A(n1413), .B(n1318), .ZN(n1198) );
XNOR2_X1 U1123 ( .A(n1357), .B(KEYINPUT52), .ZN(n1318) );
INV_X1 U1124 ( .A(G143), .ZN(n1357) );
XOR2_X1 U1125 ( .A(n1414), .B(n1415), .Z(n1413) );
NOR2_X1 U1126 ( .A1(n1361), .A2(n1416), .ZN(n1415) );
INV_X1 U1127 ( .A(G210), .ZN(n1416) );
NAND2_X1 U1128 ( .A1(n1094), .A2(n1306), .ZN(n1361) );
INV_X1 U1129 ( .A(G237), .ZN(n1306) );
INV_X1 U1130 ( .A(G953), .ZN(n1094) );
NAND3_X1 U1131 ( .A1(n1417), .A2(n1418), .A3(n1419), .ZN(n1414) );
OR2_X1 U1132 ( .A1(n1331), .A2(n1420), .ZN(n1419) );
NAND2_X1 U1133 ( .A1(G116), .A2(n1295), .ZN(n1331) );
NAND3_X1 U1134 ( .A1(n1420), .A2(n1388), .A3(n1295), .ZN(n1418) );
INV_X1 U1135 ( .A(G119), .ZN(n1295) );
INV_X1 U1136 ( .A(G116), .ZN(n1388) );
NAND2_X1 U1137 ( .A1(n1421), .A2(G119), .ZN(n1417) );
XNOR2_X1 U1138 ( .A(n1420), .B(G116), .ZN(n1421) );
XOR2_X1 U1139 ( .A(G113), .B(n1349), .Z(n1420) );
XOR2_X1 U1140 ( .A(n1160), .B(n1422), .Z(n1349) );
XNOR2_X1 U1141 ( .A(n1423), .B(KEYINPUT49), .ZN(n1422) );
NAND2_X1 U1142 ( .A1(n1424), .A2(KEYINPUT54), .ZN(n1423) );
XNOR2_X1 U1143 ( .A(G137), .B(KEYINPUT61), .ZN(n1424) );
XOR2_X1 U1144 ( .A(n1425), .B(n1403), .Z(n1160) );
INV_X1 U1145 ( .A(n1317), .ZN(n1403) );
XOR2_X1 U1146 ( .A(G128), .B(G146), .Z(n1317) );
XNOR2_X1 U1147 ( .A(G134), .B(G131), .ZN(n1425) );
NAND2_X1 U1148 ( .A1(KEYINPUT46), .A2(n1426), .ZN(n1412) );
XNOR2_X1 U1149 ( .A(KEYINPUT19), .B(n1200), .ZN(n1426) );
INV_X1 U1150 ( .A(G101), .ZN(n1200) );
NOR2_X1 U1151 ( .A1(KEYINPUT16), .A2(n1173), .ZN(n1301) );
INV_X1 U1152 ( .A(G110), .ZN(n1173) );
endmodule


