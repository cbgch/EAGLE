//Key = 0000010101110101001111110100101111001110100010001111110011101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349;

XNOR2_X1 U754 ( .A(G107), .B(n1034), .ZN(G9) );
NOR2_X1 U755 ( .A1(n1035), .A2(n1036), .ZN(G75) );
NOR4_X1 U756 ( .A1(n1037), .A2(n1038), .A3(G953), .A4(n1039), .ZN(n1036) );
NOR3_X1 U757 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1038) );
NOR2_X1 U758 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR3_X1 U759 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NOR3_X1 U760 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1043) );
NOR2_X1 U761 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U762 ( .A1(n1053), .A2(n1045), .ZN(n1052) );
NOR2_X1 U763 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U764 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U765 ( .A1(n1058), .A2(n1047), .ZN(n1051) );
NOR2_X1 U766 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND3_X1 U767 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1037) );
NAND4_X1 U768 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1062) );
NOR3_X1 U769 ( .A1(n1045), .A2(n1048), .A3(n1047), .ZN(n1067) );
INV_X1 U770 ( .A(n1068), .ZN(n1048) );
INV_X1 U771 ( .A(n1069), .ZN(n1045) );
INV_X1 U772 ( .A(n1040), .ZN(n1066) );
NAND2_X1 U773 ( .A1(n1049), .A2(n1042), .ZN(n1065) );
INV_X1 U774 ( .A(n1070), .ZN(n1042) );
NAND3_X1 U775 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1064) );
NOR3_X1 U776 ( .A1(n1039), .A2(G953), .A3(G952), .ZN(n1035) );
AND4_X1 U777 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1039) );
NOR4_X1 U778 ( .A1(n1078), .A2(n1079), .A3(n1047), .A4(n1080), .ZN(n1077) );
XNOR2_X1 U779 ( .A(KEYINPUT41), .B(n1081), .ZN(n1080) );
XOR2_X1 U780 ( .A(n1082), .B(n1083), .Z(n1078) );
NOR2_X1 U781 ( .A1(KEYINPUT8), .A2(n1084), .ZN(n1083) );
XOR2_X1 U782 ( .A(KEYINPUT26), .B(G472), .Z(n1084) );
NOR3_X1 U783 ( .A1(n1085), .A2(n1086), .A3(n1049), .ZN(n1076) );
AND2_X1 U784 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NAND2_X1 U785 ( .A1(G478), .A2(n1089), .ZN(n1075) );
XOR2_X1 U786 ( .A(KEYINPUT52), .B(n1090), .Z(n1074) );
NOR2_X1 U787 ( .A1(n1088), .A2(n1091), .ZN(n1090) );
XOR2_X1 U788 ( .A(n1087), .B(KEYINPUT34), .Z(n1091) );
XOR2_X1 U789 ( .A(n1092), .B(n1093), .Z(G72) );
NAND2_X1 U790 ( .A1(G953), .A2(n1094), .ZN(n1093) );
NAND2_X1 U791 ( .A1(G900), .A2(G227), .ZN(n1094) );
NAND2_X1 U792 ( .A1(KEYINPUT48), .A2(n1095), .ZN(n1092) );
XOR2_X1 U793 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U794 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U795 ( .A1(n1100), .A2(n1101), .ZN(n1096) );
NAND2_X1 U796 ( .A1(G953), .A2(n1102), .ZN(n1101) );
XOR2_X1 U797 ( .A(n1103), .B(n1104), .Z(n1100) );
XOR2_X1 U798 ( .A(KEYINPUT47), .B(KEYINPUT45), .Z(n1104) );
XNOR2_X1 U799 ( .A(n1105), .B(n1106), .ZN(n1103) );
XOR2_X1 U800 ( .A(n1107), .B(n1108), .Z(G69) );
NOR2_X1 U801 ( .A1(n1109), .A2(n1098), .ZN(n1108) );
AND2_X1 U802 ( .A1(G224), .A2(G898), .ZN(n1109) );
NAND2_X1 U803 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
NAND2_X1 U804 ( .A1(n1112), .A2(n1098), .ZN(n1111) );
XNOR2_X1 U805 ( .A(n1113), .B(n1063), .ZN(n1112) );
NAND3_X1 U806 ( .A1(G898), .A2(n1113), .A3(G953), .ZN(n1110) );
XNOR2_X1 U807 ( .A(n1114), .B(n1115), .ZN(n1113) );
XOR2_X1 U808 ( .A(n1116), .B(KEYINPUT57), .Z(n1114) );
NAND2_X1 U809 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NOR2_X1 U810 ( .A1(n1119), .A2(n1120), .ZN(G66) );
XOR2_X1 U811 ( .A(n1121), .B(n1122), .Z(n1120) );
NAND2_X1 U812 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
NOR2_X1 U813 ( .A1(n1119), .A2(n1125), .ZN(G63) );
XNOR2_X1 U814 ( .A(n1126), .B(n1127), .ZN(n1125) );
NAND2_X1 U815 ( .A1(n1123), .A2(G478), .ZN(n1126) );
NOR2_X1 U816 ( .A1(n1119), .A2(n1128), .ZN(G60) );
XOR2_X1 U817 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U818 ( .A(KEYINPUT49), .B(n1131), .Z(n1130) );
NOR2_X1 U819 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XOR2_X1 U820 ( .A(KEYINPUT9), .B(G475), .Z(n1133) );
XNOR2_X1 U821 ( .A(G104), .B(n1134), .ZN(G6) );
NOR2_X1 U822 ( .A1(n1119), .A2(n1135), .ZN(G57) );
XOR2_X1 U823 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U824 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U825 ( .A(n1140), .B(n1141), .Z(n1139) );
AND2_X1 U826 ( .A1(G472), .A2(n1123), .ZN(n1141) );
INV_X1 U827 ( .A(n1132), .ZN(n1123) );
NAND2_X1 U828 ( .A1(KEYINPUT21), .A2(n1142), .ZN(n1140) );
XNOR2_X1 U829 ( .A(KEYINPUT31), .B(n1143), .ZN(n1142) );
XOR2_X1 U830 ( .A(n1144), .B(KEYINPUT60), .Z(n1138) );
XNOR2_X1 U831 ( .A(n1145), .B(n1146), .ZN(n1136) );
XNOR2_X1 U832 ( .A(n1147), .B(n1148), .ZN(n1145) );
NOR2_X1 U833 ( .A1(n1119), .A2(n1149), .ZN(G54) );
XOR2_X1 U834 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U835 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U836 ( .A(n1154), .B(n1155), .Z(n1150) );
XNOR2_X1 U837 ( .A(KEYINPUT29), .B(n1156), .ZN(n1155) );
NOR3_X1 U838 ( .A1(n1132), .A2(KEYINPUT61), .A3(n1157), .ZN(n1156) );
NOR2_X1 U839 ( .A1(n1119), .A2(n1158), .ZN(G51) );
XOR2_X1 U840 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U841 ( .A(KEYINPUT56), .B(n1161), .Z(n1160) );
NOR2_X1 U842 ( .A1(n1087), .A2(n1132), .ZN(n1161) );
NAND2_X1 U843 ( .A1(G902), .A2(n1162), .ZN(n1132) );
NAND2_X1 U844 ( .A1(n1063), .A2(n1061), .ZN(n1162) );
INV_X1 U845 ( .A(n1099), .ZN(n1061) );
NAND4_X1 U846 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1099) );
NOR4_X1 U847 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
NOR3_X1 U848 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1165) );
NOR2_X1 U849 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
INV_X1 U850 ( .A(KEYINPUT44), .ZN(n1174) );
NOR4_X1 U851 ( .A1(KEYINPUT44), .A2(n1176), .A3(n1081), .A4(n1177), .ZN(n1172) );
NAND2_X1 U852 ( .A1(n1072), .A2(n1178), .ZN(n1176) );
INV_X1 U853 ( .A(n1179), .ZN(n1072) );
NOR3_X1 U854 ( .A1(n1180), .A2(n1071), .A3(n1181), .ZN(n1171) );
XOR2_X1 U855 ( .A(KEYINPUT18), .B(n1060), .Z(n1181) );
NAND3_X1 U856 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1180) );
AND4_X1 U857 ( .A1(n1185), .A2(n1034), .A3(n1186), .A4(n1187), .ZN(n1063) );
NOR4_X1 U858 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187) );
NOR2_X1 U859 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XNOR2_X1 U860 ( .A(n1194), .B(KEYINPUT43), .ZN(n1192) );
NOR2_X1 U861 ( .A1(n1046), .A2(n1195), .ZN(n1190) );
INV_X1 U862 ( .A(n1182), .ZN(n1046) );
INV_X1 U863 ( .A(n1134), .ZN(n1189) );
NAND3_X1 U864 ( .A1(n1070), .A2(n1196), .A3(n1060), .ZN(n1134) );
INV_X1 U865 ( .A(n1197), .ZN(n1188) );
NOR2_X1 U866 ( .A1(n1198), .A2(n1199), .ZN(n1186) );
NAND3_X1 U867 ( .A1(n1070), .A2(n1196), .A3(n1059), .ZN(n1034) );
NOR2_X1 U868 ( .A1(n1098), .A2(G952), .ZN(n1119) );
XNOR2_X1 U869 ( .A(G146), .B(n1163), .ZN(G48) );
NAND3_X1 U870 ( .A1(n1194), .A2(n1060), .A3(n1200), .ZN(n1163) );
XOR2_X1 U871 ( .A(n1175), .B(n1201), .Z(G45) );
XOR2_X1 U872 ( .A(KEYINPUT19), .B(G143), .Z(n1201) );
NAND4_X1 U873 ( .A1(n1200), .A2(n1179), .A3(n1202), .A4(n1178), .ZN(n1175) );
XNOR2_X1 U874 ( .A(n1164), .B(n1203), .ZN(G42) );
NOR2_X1 U875 ( .A1(KEYINPUT1), .A2(n1204), .ZN(n1203) );
NAND3_X1 U876 ( .A1(n1205), .A2(n1060), .A3(n1206), .ZN(n1164) );
XNOR2_X1 U877 ( .A(n1207), .B(n1170), .ZN(G39) );
AND3_X1 U878 ( .A1(n1194), .A2(n1069), .A3(n1206), .ZN(n1170) );
XOR2_X1 U879 ( .A(G134), .B(n1169), .Z(G36) );
AND3_X1 U880 ( .A1(n1179), .A2(n1059), .A3(n1206), .ZN(n1169) );
XOR2_X1 U881 ( .A(G131), .B(n1168), .Z(G33) );
AND3_X1 U882 ( .A1(n1060), .A2(n1179), .A3(n1206), .ZN(n1168) );
AND4_X1 U883 ( .A1(n1055), .A2(n1068), .A3(n1183), .A4(n1073), .ZN(n1206) );
XOR2_X1 U884 ( .A(G128), .B(n1167), .Z(G30) );
AND3_X1 U885 ( .A1(n1194), .A2(n1059), .A3(n1200), .ZN(n1167) );
INV_X1 U886 ( .A(n1177), .ZN(n1200) );
NAND3_X1 U887 ( .A1(n1182), .A2(n1183), .A3(n1055), .ZN(n1177) );
XNOR2_X1 U888 ( .A(n1143), .B(n1208), .ZN(G3) );
NOR2_X1 U889 ( .A1(KEYINPUT14), .A2(n1197), .ZN(n1208) );
NAND3_X1 U890 ( .A1(n1179), .A2(n1196), .A3(n1069), .ZN(n1197) );
AND3_X1 U891 ( .A1(n1182), .A2(n1209), .A3(n1055), .ZN(n1196) );
NAND2_X1 U892 ( .A1(n1210), .A2(n1211), .ZN(G27) );
NAND2_X1 U893 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NAND2_X1 U894 ( .A1(G125), .A2(n1214), .ZN(n1210) );
NAND2_X1 U895 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND2_X1 U896 ( .A1(KEYINPUT24), .A2(n1217), .ZN(n1216) );
INV_X1 U897 ( .A(n1218), .ZN(n1217) );
OR2_X1 U898 ( .A1(n1212), .A2(KEYINPUT24), .ZN(n1215) );
NOR2_X1 U899 ( .A1(KEYINPUT3), .A2(n1218), .ZN(n1212) );
NAND4_X1 U900 ( .A1(n1182), .A2(n1183), .A3(n1060), .A4(n1219), .ZN(n1218) );
NOR2_X1 U901 ( .A1(n1071), .A2(n1220), .ZN(n1219) );
XNOR2_X1 U902 ( .A(KEYINPUT40), .B(n1047), .ZN(n1220) );
INV_X1 U903 ( .A(n1184), .ZN(n1047) );
INV_X1 U904 ( .A(n1205), .ZN(n1071) );
NAND2_X1 U905 ( .A1(n1040), .A2(n1221), .ZN(n1183) );
NAND4_X1 U906 ( .A1(G953), .A2(G902), .A3(n1222), .A4(n1102), .ZN(n1221) );
INV_X1 U907 ( .A(G900), .ZN(n1102) );
XNOR2_X1 U908 ( .A(G122), .B(n1185), .ZN(G24) );
NAND4_X1 U909 ( .A1(n1223), .A2(n1070), .A3(n1202), .A4(n1178), .ZN(n1185) );
NOR2_X1 U910 ( .A1(n1224), .A2(n1079), .ZN(n1070) );
XOR2_X1 U911 ( .A(n1225), .B(n1226), .Z(G21) );
NOR2_X1 U912 ( .A1(n1227), .A2(n1193), .ZN(n1226) );
NAND2_X1 U913 ( .A1(n1069), .A2(n1223), .ZN(n1193) );
INV_X1 U914 ( .A(n1194), .ZN(n1227) );
NOR2_X1 U915 ( .A1(n1228), .A2(n1229), .ZN(n1194) );
NOR2_X1 U916 ( .A1(KEYINPUT55), .A2(n1230), .ZN(n1225) );
XOR2_X1 U917 ( .A(n1199), .B(n1231), .Z(G18) );
NOR2_X1 U918 ( .A1(KEYINPUT42), .A2(n1232), .ZN(n1231) );
AND3_X1 U919 ( .A1(n1223), .A2(n1059), .A3(n1179), .ZN(n1199) );
NOR2_X1 U920 ( .A1(n1202), .A2(n1233), .ZN(n1059) );
XNOR2_X1 U921 ( .A(n1234), .B(n1198), .ZN(G15) );
AND3_X1 U922 ( .A1(n1179), .A2(n1223), .A3(n1060), .ZN(n1198) );
NOR2_X1 U923 ( .A1(n1178), .A2(n1081), .ZN(n1060) );
INV_X1 U924 ( .A(n1202), .ZN(n1081) );
AND3_X1 U925 ( .A1(n1182), .A2(n1209), .A3(n1184), .ZN(n1223) );
NOR2_X1 U926 ( .A1(n1056), .A2(n1235), .ZN(n1184) );
INV_X1 U927 ( .A(n1057), .ZN(n1235) );
NOR2_X1 U928 ( .A1(n1079), .A2(n1229), .ZN(n1179) );
INV_X1 U929 ( .A(n1224), .ZN(n1229) );
XOR2_X1 U930 ( .A(n1236), .B(n1237), .Z(G12) );
NAND2_X1 U931 ( .A1(KEYINPUT10), .A2(G110), .ZN(n1237) );
NAND2_X1 U932 ( .A1(n1238), .A2(n1182), .ZN(n1236) );
NOR2_X1 U933 ( .A1(n1068), .A2(n1049), .ZN(n1182) );
INV_X1 U934 ( .A(n1073), .ZN(n1049) );
NAND2_X1 U935 ( .A1(G214), .A2(n1239), .ZN(n1073) );
XNOR2_X1 U936 ( .A(n1240), .B(n1088), .ZN(n1068) );
AND2_X1 U937 ( .A1(n1159), .A2(n1241), .ZN(n1088) );
XOR2_X1 U938 ( .A(n1242), .B(n1243), .Z(n1159) );
XNOR2_X1 U939 ( .A(n1244), .B(n1245), .ZN(n1243) );
NAND2_X1 U940 ( .A1(G224), .A2(n1098), .ZN(n1244) );
XOR2_X1 U941 ( .A(n1246), .B(n1247), .Z(n1242) );
NOR2_X1 U942 ( .A1(KEYINPUT27), .A2(n1115), .ZN(n1247) );
XNOR2_X1 U943 ( .A(G110), .B(n1248), .ZN(n1115) );
XNOR2_X1 U944 ( .A(n1249), .B(n1213), .ZN(n1246) );
INV_X1 U945 ( .A(G125), .ZN(n1213) );
NAND2_X1 U946 ( .A1(n1250), .A2(n1118), .ZN(n1249) );
NAND3_X1 U947 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1118) );
XNOR2_X1 U948 ( .A(G113), .B(n1254), .ZN(n1253) );
NAND2_X1 U949 ( .A1(n1255), .A2(n1143), .ZN(n1252) );
NAND2_X1 U950 ( .A1(G101), .A2(n1256), .ZN(n1251) );
XOR2_X1 U951 ( .A(n1117), .B(KEYINPUT39), .Z(n1250) );
NAND3_X1 U952 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1117) );
XNOR2_X1 U953 ( .A(n1254), .B(n1234), .ZN(n1259) );
NAND2_X1 U954 ( .A1(KEYINPUT23), .A2(n1260), .ZN(n1254) );
XNOR2_X1 U955 ( .A(n1230), .B(G116), .ZN(n1260) );
OR2_X1 U956 ( .A1(n1256), .A2(n1143), .ZN(n1258) );
OR2_X1 U957 ( .A1(n1255), .A2(G101), .ZN(n1257) );
XNOR2_X1 U958 ( .A(n1261), .B(n1256), .ZN(n1255) );
XOR2_X1 U959 ( .A(G104), .B(G107), .Z(n1256) );
XNOR2_X1 U960 ( .A(KEYINPUT6), .B(KEYINPUT22), .ZN(n1261) );
NAND2_X1 U961 ( .A1(KEYINPUT7), .A2(n1087), .ZN(n1240) );
NAND2_X1 U962 ( .A1(G210), .A2(n1239), .ZN(n1087) );
NAND2_X1 U963 ( .A1(n1262), .A2(n1241), .ZN(n1239) );
XOR2_X1 U964 ( .A(n1195), .B(KEYINPUT36), .Z(n1238) );
NAND4_X1 U965 ( .A1(n1205), .A2(n1069), .A3(n1055), .A4(n1209), .ZN(n1195) );
NAND2_X1 U966 ( .A1(n1263), .A2(n1040), .ZN(n1209) );
NAND3_X1 U967 ( .A1(n1222), .A2(n1098), .A3(G952), .ZN(n1040) );
XOR2_X1 U968 ( .A(KEYINPUT38), .B(n1264), .Z(n1263) );
NOR4_X1 U969 ( .A1(G898), .A2(n1265), .A3(n1241), .A4(n1098), .ZN(n1264) );
INV_X1 U970 ( .A(n1222), .ZN(n1265) );
NAND2_X1 U971 ( .A1(G237), .A2(G234), .ZN(n1222) );
AND2_X1 U972 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U973 ( .A1(G221), .A2(n1266), .ZN(n1057) );
XOR2_X1 U974 ( .A(n1267), .B(n1157), .Z(n1056) );
INV_X1 U975 ( .A(G469), .ZN(n1157) );
NAND2_X1 U976 ( .A1(n1268), .A2(n1241), .ZN(n1267) );
XOR2_X1 U977 ( .A(n1152), .B(n1269), .Z(n1268) );
XNOR2_X1 U978 ( .A(n1154), .B(n1270), .ZN(n1269) );
NOR2_X1 U979 ( .A1(KEYINPUT16), .A2(n1153), .ZN(n1270) );
XNOR2_X1 U980 ( .A(G110), .B(G140), .ZN(n1153) );
NAND2_X1 U981 ( .A1(G227), .A2(n1098), .ZN(n1154) );
XNOR2_X1 U982 ( .A(n1271), .B(n1272), .ZN(n1152) );
INV_X1 U983 ( .A(n1105), .ZN(n1272) );
XOR2_X1 U984 ( .A(n1273), .B(n1274), .Z(n1105) );
XNOR2_X1 U985 ( .A(G146), .B(n1275), .ZN(n1273) );
XOR2_X1 U986 ( .A(n1276), .B(KEYINPUT5), .Z(n1271) );
NAND2_X1 U987 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND2_X1 U988 ( .A1(G101), .A2(n1279), .ZN(n1278) );
XOR2_X1 U989 ( .A(KEYINPUT33), .B(n1280), .Z(n1277) );
NOR2_X1 U990 ( .A1(G101), .A2(n1279), .ZN(n1280) );
XNOR2_X1 U991 ( .A(n1281), .B(n1282), .ZN(n1279) );
NOR2_X1 U992 ( .A1(KEYINPUT35), .A2(n1283), .ZN(n1282) );
INV_X1 U993 ( .A(G104), .ZN(n1283) );
NOR2_X1 U994 ( .A1(n1178), .A2(n1202), .ZN(n1069) );
XNOR2_X1 U995 ( .A(n1284), .B(G475), .ZN(n1202) );
NAND2_X1 U996 ( .A1(n1129), .A2(n1241), .ZN(n1284) );
XNOR2_X1 U997 ( .A(n1285), .B(n1286), .ZN(n1129) );
XOR2_X1 U998 ( .A(n1287), .B(n1288), .Z(n1286) );
XNOR2_X1 U999 ( .A(G131), .B(n1248), .ZN(n1288) );
XNOR2_X1 U1000 ( .A(n1289), .B(G143), .ZN(n1287) );
XOR2_X1 U1001 ( .A(n1290), .B(n1291), .Z(n1285) );
XNOR2_X1 U1002 ( .A(n1234), .B(n1292), .ZN(n1291) );
NOR2_X1 U1003 ( .A1(KEYINPUT12), .A2(n1293), .ZN(n1292) );
XOR2_X1 U1004 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U1005 ( .A(G125), .B(KEYINPUT17), .ZN(n1295) );
NAND2_X1 U1006 ( .A1(KEYINPUT53), .A2(n1204), .ZN(n1294) );
XOR2_X1 U1007 ( .A(n1296), .B(n1297), .Z(n1290) );
NOR4_X1 U1008 ( .A1(KEYINPUT2), .A2(G953), .A3(G237), .A4(n1298), .ZN(n1297) );
INV_X1 U1009 ( .A(G214), .ZN(n1298) );
NAND2_X1 U1010 ( .A1(KEYINPUT63), .A2(G104), .ZN(n1296) );
INV_X1 U1011 ( .A(n1233), .ZN(n1178) );
NOR2_X1 U1012 ( .A1(n1299), .A2(n1086), .ZN(n1233) );
NOR2_X1 U1013 ( .A1(n1089), .A2(G478), .ZN(n1086) );
AND2_X1 U1014 ( .A1(n1300), .A2(n1089), .ZN(n1299) );
NAND2_X1 U1015 ( .A1(n1301), .A2(n1241), .ZN(n1089) );
XNOR2_X1 U1016 ( .A(KEYINPUT28), .B(n1302), .ZN(n1301) );
INV_X1 U1017 ( .A(n1127), .ZN(n1302) );
XNOR2_X1 U1018 ( .A(n1303), .B(n1304), .ZN(n1127) );
XOR2_X1 U1019 ( .A(n1305), .B(n1306), .Z(n1304) );
NAND3_X1 U1020 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1306) );
NAND2_X1 U1021 ( .A1(G134), .A2(n1310), .ZN(n1309) );
OR3_X1 U1022 ( .A1(n1310), .A2(G134), .A3(n1311), .ZN(n1308) );
INV_X1 U1023 ( .A(KEYINPUT50), .ZN(n1310) );
NAND2_X1 U1024 ( .A1(n1311), .A2(n1312), .ZN(n1307) );
NAND2_X1 U1025 ( .A1(n1313), .A2(KEYINPUT50), .ZN(n1312) );
XNOR2_X1 U1026 ( .A(G134), .B(KEYINPUT4), .ZN(n1313) );
XOR2_X1 U1027 ( .A(n1275), .B(KEYINPUT59), .Z(n1311) );
NAND3_X1 U1028 ( .A1(G217), .A2(n1098), .A3(G234), .ZN(n1305) );
NAND2_X1 U1029 ( .A1(n1314), .A2(n1315), .ZN(n1303) );
NAND2_X1 U1030 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XNOR2_X1 U1031 ( .A(KEYINPUT25), .B(n1281), .ZN(n1316) );
OR2_X1 U1032 ( .A1(n1281), .A2(n1317), .ZN(n1314) );
XNOR2_X1 U1033 ( .A(n1318), .B(n1232), .ZN(n1317) );
NAND2_X1 U1034 ( .A1(KEYINPUT11), .A2(n1248), .ZN(n1318) );
INV_X1 U1035 ( .A(G122), .ZN(n1248) );
INV_X1 U1036 ( .A(G107), .ZN(n1281) );
XNOR2_X1 U1037 ( .A(G478), .B(KEYINPUT62), .ZN(n1300) );
NOR2_X1 U1038 ( .A1(n1224), .A2(n1228), .ZN(n1205) );
INV_X1 U1039 ( .A(n1079), .ZN(n1228) );
XNOR2_X1 U1040 ( .A(n1319), .B(n1124), .ZN(n1079) );
AND2_X1 U1041 ( .A1(G217), .A2(n1266), .ZN(n1124) );
NAND2_X1 U1042 ( .A1(G234), .A2(n1241), .ZN(n1266) );
NAND2_X1 U1043 ( .A1(n1122), .A2(n1241), .ZN(n1319) );
XOR2_X1 U1044 ( .A(n1320), .B(n1321), .Z(n1122) );
XOR2_X1 U1045 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U1046 ( .A(n1324), .B(G110), .Z(n1323) );
NAND2_X1 U1047 ( .A1(n1325), .A2(KEYINPUT58), .ZN(n1324) );
XNOR2_X1 U1048 ( .A(n1326), .B(n1230), .ZN(n1325) );
INV_X1 U1049 ( .A(G119), .ZN(n1230) );
NAND2_X1 U1050 ( .A1(n1327), .A2(KEYINPUT20), .ZN(n1326) );
XNOR2_X1 U1051 ( .A(G128), .B(KEYINPUT0), .ZN(n1327) );
NAND2_X1 U1052 ( .A1(n1328), .A2(n1329), .ZN(n1322) );
NAND2_X1 U1053 ( .A1(G146), .A2(n1106), .ZN(n1329) );
XOR2_X1 U1054 ( .A(n1330), .B(KEYINPUT54), .Z(n1328) );
OR2_X1 U1055 ( .A1(n1106), .A2(G146), .ZN(n1330) );
XNOR2_X1 U1056 ( .A(G125), .B(n1204), .ZN(n1106) );
INV_X1 U1057 ( .A(G140), .ZN(n1204) );
XOR2_X1 U1058 ( .A(n1331), .B(n1332), .Z(n1320) );
AND3_X1 U1059 ( .A1(G221), .A2(n1098), .A3(G234), .ZN(n1332) );
NAND2_X1 U1060 ( .A1(KEYINPUT51), .A2(n1207), .ZN(n1331) );
XNOR2_X1 U1061 ( .A(n1082), .B(G472), .ZN(n1224) );
NAND2_X1 U1062 ( .A1(n1333), .A2(n1241), .ZN(n1082) );
INV_X1 U1063 ( .A(G902), .ZN(n1241) );
XOR2_X1 U1064 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1065 ( .A(n1336), .B(n1148), .Z(n1335) );
XNOR2_X1 U1066 ( .A(n1337), .B(n1338), .ZN(n1148) );
XNOR2_X1 U1067 ( .A(G119), .B(n1339), .ZN(n1338) );
NAND2_X1 U1068 ( .A1(KEYINPUT15), .A2(n1232), .ZN(n1339) );
INV_X1 U1069 ( .A(G116), .ZN(n1232) );
NAND2_X1 U1070 ( .A1(KEYINPUT37), .A2(n1234), .ZN(n1337) );
INV_X1 U1071 ( .A(G113), .ZN(n1234) );
XNOR2_X1 U1072 ( .A(n1340), .B(n1144), .ZN(n1336) );
NAND3_X1 U1073 ( .A1(n1262), .A2(n1098), .A3(G210), .ZN(n1144) );
INV_X1 U1074 ( .A(G953), .ZN(n1098) );
INV_X1 U1075 ( .A(G237), .ZN(n1262) );
NAND2_X1 U1076 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
NAND2_X1 U1077 ( .A1(n1245), .A2(n1147), .ZN(n1342) );
INV_X1 U1078 ( .A(n1146), .ZN(n1245) );
XOR2_X1 U1079 ( .A(n1343), .B(KEYINPUT46), .Z(n1341) );
NAND2_X1 U1080 ( .A1(n1274), .A2(n1146), .ZN(n1343) );
NAND2_X1 U1081 ( .A1(n1344), .A2(n1345), .ZN(n1146) );
NAND2_X1 U1082 ( .A1(n1346), .A2(n1289), .ZN(n1345) );
INV_X1 U1083 ( .A(G146), .ZN(n1289) );
XNOR2_X1 U1084 ( .A(KEYINPUT13), .B(n1347), .ZN(n1346) );
INV_X1 U1085 ( .A(n1275), .ZN(n1347) );
NAND2_X1 U1086 ( .A1(n1275), .A2(G146), .ZN(n1344) );
XOR2_X1 U1087 ( .A(G128), .B(G143), .Z(n1275) );
INV_X1 U1088 ( .A(n1147), .ZN(n1274) );
XOR2_X1 U1089 ( .A(G131), .B(n1348), .Z(n1147) );
XNOR2_X1 U1090 ( .A(n1207), .B(G134), .ZN(n1348) );
INV_X1 U1091 ( .A(G137), .ZN(n1207) );
XNOR2_X1 U1092 ( .A(n1349), .B(n1143), .ZN(n1334) );
INV_X1 U1093 ( .A(G101), .ZN(n1143) );
XNOR2_X1 U1094 ( .A(KEYINPUT32), .B(KEYINPUT30), .ZN(n1349) );
endmodule


