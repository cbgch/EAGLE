//Key = 0000011011111001110111101111101000011111011101010000110011111110


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
n2164, n2165, n2166, n2167;

OR2_X1 U1219 ( .A1(n1776), .A2(STATO_REG_0__SCAN_IN), .ZN(n1634) );
INV_X2 U1220 ( .A(n1634), .ZN(n1635) );
INV_X2 U1221 ( .A(U280), .ZN(n1779) );
INV_X1 U1222 ( .A(n1636), .ZN(U375) );
NAND2_X1 U1223 ( .A1(n1637), .A2(n1638), .ZN(U344) );
NAND2_X1 U1224 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1639), .ZN(n1638) );
NAND2_X1 U1225 ( .A1(n1640), .A2(DATA_IN_7_), .ZN(n1637) );
NAND2_X1 U1226 ( .A1(n1641), .A2(n1642), .ZN(U343) );
NAND2_X1 U1227 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1639), .ZN(n1642) );
NAND2_X1 U1228 ( .A1(n1640), .A2(DATA_IN_6_), .ZN(n1641) );
NAND2_X1 U1229 ( .A1(n1643), .A2(n1644), .ZN(U342) );
NAND2_X1 U1230 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1639), .ZN(n1644) );
NAND2_X1 U1231 ( .A1(n1640), .A2(DATA_IN_5_), .ZN(n1643) );
NAND2_X1 U1232 ( .A1(n1645), .A2(n1646), .ZN(U341) );
NAND2_X1 U1233 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1639), .ZN(n1646) );
NAND2_X1 U1234 ( .A1(n1640), .A2(DATA_IN_4_), .ZN(n1645) );
NAND2_X1 U1235 ( .A1(n1647), .A2(n1648), .ZN(U340) );
NAND2_X1 U1236 ( .A1(n1649), .A2(n1639), .ZN(n1648) );
XOR2_X1 U1237 ( .A(n1650), .B(KEYINPUT12), .Z(n1649) );
NAND2_X1 U1238 ( .A1(n1640), .A2(DATA_IN_3_), .ZN(n1647) );
NAND2_X1 U1239 ( .A1(n1651), .A2(n1652), .ZN(U339) );
NAND2_X1 U1240 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1639), .ZN(n1652) );
NAND2_X1 U1241 ( .A1(n1640), .A2(DATA_IN_2_), .ZN(n1651) );
NAND2_X1 U1242 ( .A1(n1653), .A2(n1654), .ZN(U338) );
NAND2_X1 U1243 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1639), .ZN(n1654) );
NAND2_X1 U1244 ( .A1(n1640), .A2(DATA_IN_1_), .ZN(n1653) );
NAND2_X1 U1245 ( .A1(n1655), .A2(n1656), .ZN(U337) );
NAND2_X1 U1246 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1639), .ZN(n1656) );
NAND2_X1 U1247 ( .A1(n1657), .A2(n1658), .ZN(n1639) );
XOR2_X1 U1248 ( .A(n1636), .B(KEYINPUT63), .Z(n1657) );
NAND2_X1 U1249 ( .A1(n1640), .A2(DATA_IN_0_), .ZN(n1655) );
AND2_X1 U1250 ( .A1(n1658), .A2(n1636), .ZN(n1640) );
NAND2_X1 U1251 ( .A1(n1659), .A2(n1660), .ZN(n1658) );
NAND2_X1 U1252 ( .A1(n1661), .A2(n1662), .ZN(U336) );
NAND2_X1 U1253 ( .A1(n1663), .A2(n1664), .ZN(n1662) );
XOR2_X1 U1254 ( .A(RMIN_REG_7__SCAN_IN), .B(KEYINPUT33), .Z(n1663) );
NAND2_X1 U1255 ( .A1(n1665), .A2(DATA_IN_7_), .ZN(n1661) );
NAND2_X1 U1256 ( .A1(n1666), .A2(n1667), .ZN(U335) );
NAND2_X1 U1257 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1664), .ZN(n1667) );
NAND2_X1 U1258 ( .A1(n1665), .A2(DATA_IN_6_), .ZN(n1666) );
NAND2_X1 U1259 ( .A1(n1668), .A2(n1669), .ZN(U334) );
NAND2_X1 U1260 ( .A1(n1670), .A2(DATA_IN_5_), .ZN(n1669) );
XOR2_X1 U1261 ( .A(n1664), .B(KEYINPUT36), .Z(n1670) );
NAND2_X1 U1262 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1664), .ZN(n1668) );
NAND2_X1 U1263 ( .A1(n1671), .A2(n1672), .ZN(U333) );
NAND2_X1 U1264 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1664), .ZN(n1672) );
NAND2_X1 U1265 ( .A1(n1665), .A2(DATA_IN_4_), .ZN(n1671) );
NAND2_X1 U1266 ( .A1(n1673), .A2(n1674), .ZN(U332) );
NAND2_X1 U1267 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1664), .ZN(n1674) );
NAND2_X1 U1268 ( .A1(n1675), .A2(n1665), .ZN(n1673) );
XOR2_X1 U1269 ( .A(n1676), .B(KEYINPUT25), .Z(n1675) );
NAND2_X1 U1270 ( .A1(n1677), .A2(n1678), .ZN(U331) );
NAND2_X1 U1271 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1664), .ZN(n1678) );
XOR2_X1 U1272 ( .A(KEYINPUT39), .B(n1679), .Z(n1677) );
NOR2_X1 U1273 ( .A1(n1680), .A2(n1664), .ZN(n1679) );
NAND2_X1 U1274 ( .A1(n1681), .A2(n1682), .ZN(U330) );
NAND2_X1 U1275 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1664), .ZN(n1682) );
NAND2_X1 U1276 ( .A1(n1665), .A2(DATA_IN_1_), .ZN(n1681) );
NAND2_X1 U1277 ( .A1(n1683), .A2(n1684), .ZN(U329) );
NAND2_X1 U1278 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1664), .ZN(n1684) );
NAND2_X1 U1279 ( .A1(n1665), .A2(DATA_IN_0_), .ZN(n1683) );
INV_X1 U1280 ( .A(n1664), .ZN(n1665) );
NAND2_X1 U1281 ( .A1(n1636), .A2(n1685), .ZN(n1664) );
NAND2_X1 U1282 ( .A1(n1686), .A2(n1660), .ZN(n1685) );
NAND2_X1 U1283 ( .A1(n1659), .A2(n1687), .ZN(n1686) );
NAND2_X1 U1284 ( .A1(n1688), .A2(n1689), .ZN(n1687) );
NAND3_X1 U1285 ( .A1(n1690), .A2(n1691), .A3(n1692), .ZN(n1689) );
NAND2_X1 U1286 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1693), .ZN(n1692) );
NAND3_X1 U1287 ( .A1(n1694), .A2(n1695), .A3(n1696), .ZN(n1691) );
NAND2_X1 U1288 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1697), .ZN(n1696) );
NAND3_X1 U1289 ( .A1(n1698), .A2(n1699), .A3(n1700), .ZN(n1695) );
NAND2_X1 U1290 ( .A1(DATA_IN_5_), .A2(n1701), .ZN(n1700) );
NAND3_X1 U1291 ( .A1(n1702), .A2(n1703), .A3(n1704), .ZN(n1699) );
NAND2_X1 U1292 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1705), .ZN(n1704) );
NAND3_X1 U1293 ( .A1(n1706), .A2(n1707), .A3(n1708), .ZN(n1703) );
NAND2_X1 U1294 ( .A1(DATA_IN_3_), .A2(n1709), .ZN(n1708) );
NAND3_X1 U1295 ( .A1(n1710), .A2(n1711), .A3(n1712), .ZN(n1707) );
NAND2_X1 U1296 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1713), .ZN(n1712) );
NAND2_X1 U1297 ( .A1(n1714), .A2(n1715), .ZN(n1711) );
XOR2_X1 U1298 ( .A(KEYINPUT58), .B(DATA_IN_2_), .Z(n1715) );
XOR2_X1 U1299 ( .A(n1716), .B(KEYINPUT26), .Z(n1714) );
NAND3_X1 U1300 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1717), .A3(n1718), .ZN(n1710) );
XNOR2_X1 U1301 ( .A(DATA_IN_0_), .B(KEYINPUT14), .ZN(n1718) );
NAND2_X1 U1302 ( .A1(DATA_IN_1_), .A2(n1719), .ZN(n1717) );
NAND2_X1 U1303 ( .A1(DATA_IN_2_), .A2(n1716), .ZN(n1706) );
NAND2_X1 U1304 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1676), .ZN(n1702) );
NAND2_X1 U1305 ( .A1(DATA_IN_4_), .A2(n1720), .ZN(n1698) );
NAND2_X1 U1306 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1721), .ZN(n1694) );
OR2_X1 U1307 ( .A1(n1697), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1690) );
NAND2_X1 U1308 ( .A1(DATA_IN_7_), .A2(n1722), .ZN(n1688) );
AND2_X1 U1309 ( .A1(n1723), .A2(n1724), .ZN(n1659) );
NAND2_X1 U1310 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1693), .ZN(n1724) );
INV_X1 U1311 ( .A(DATA_IN_7_), .ZN(n1693) );
NAND3_X1 U1312 ( .A1(n1725), .A2(n1726), .A3(n1727), .ZN(n1723) );
NAND2_X1 U1313 ( .A1(DATA_IN_7_), .A2(n1728), .ZN(n1727) );
NAND3_X1 U1314 ( .A1(n1729), .A2(n1730), .A3(n1731), .ZN(n1726) );
NAND2_X1 U1315 ( .A1(DATA_IN_6_), .A2(n1732), .ZN(n1731) );
NAND3_X1 U1316 ( .A1(n1733), .A2(n1734), .A3(n1735), .ZN(n1730) );
NAND2_X1 U1317 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1721), .ZN(n1735) );
NAND3_X1 U1318 ( .A1(n1736), .A2(n1737), .A3(n1738), .ZN(n1734) );
NAND2_X1 U1319 ( .A1(DATA_IN_4_), .A2(n1739), .ZN(n1738) );
NAND3_X1 U1320 ( .A1(n1740), .A2(n1741), .A3(n1742), .ZN(n1737) );
NAND2_X1 U1321 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1676), .ZN(n1742) );
NAND3_X1 U1322 ( .A1(n1743), .A2(n1744), .A3(n1745), .ZN(n1741) );
NAND2_X1 U1323 ( .A1(DATA_IN_2_), .A2(n1746), .ZN(n1745) );
NAND3_X1 U1324 ( .A1(n1747), .A2(n1748), .A3(DATA_IN_0_), .ZN(n1744) );
NAND2_X1 U1325 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1749), .ZN(n1747) );
XOR2_X1 U1326 ( .A(KEYINPUT28), .B(DATA_IN_1_), .Z(n1749) );
NAND2_X1 U1327 ( .A1(n1750), .A2(DATA_IN_1_), .ZN(n1743) );
XOR2_X1 U1328 ( .A(n1751), .B(KEYINPUT55), .Z(n1750) );
NAND2_X1 U1329 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1680), .ZN(n1740) );
NAND2_X1 U1330 ( .A1(DATA_IN_3_), .A2(n1650), .ZN(n1736) );
NAND2_X1 U1331 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1705), .ZN(n1733) );
NAND2_X1 U1332 ( .A1(DATA_IN_5_), .A2(n1752), .ZN(n1729) );
NAND2_X1 U1333 ( .A1(n1753), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1725) );
XOR2_X1 U1334 ( .A(n1697), .B(KEYINPUT40), .Z(n1753) );
INV_X1 U1335 ( .A(DATA_IN_6_), .ZN(n1697) );
NAND2_X1 U1336 ( .A1(n1754), .A2(n1755), .ZN(U328) );
NAND2_X1 U1337 ( .A1(n1756), .A2(DATA_IN_7_), .ZN(n1755) );
NAND2_X1 U1338 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1757), .ZN(n1754) );
NAND2_X1 U1339 ( .A1(n1758), .A2(n1759), .ZN(U327) );
NAND2_X1 U1340 ( .A1(n1756), .A2(DATA_IN_6_), .ZN(n1759) );
NAND2_X1 U1341 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1757), .ZN(n1758) );
NAND2_X1 U1342 ( .A1(n1760), .A2(n1761), .ZN(U326) );
NAND2_X1 U1343 ( .A1(n1756), .A2(DATA_IN_5_), .ZN(n1761) );
NAND2_X1 U1344 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1757), .ZN(n1760) );
NAND2_X1 U1345 ( .A1(n1762), .A2(n1763), .ZN(U325) );
NAND2_X1 U1346 ( .A1(n1756), .A2(DATA_IN_4_), .ZN(n1763) );
XOR2_X1 U1347 ( .A(n1764), .B(KEYINPUT50), .Z(n1762) );
NAND2_X1 U1348 ( .A1(n1765), .A2(n1757), .ZN(n1764) );
XOR2_X1 U1349 ( .A(RLAST_REG_4__SCAN_IN), .B(KEYINPUT2), .Z(n1765) );
NAND2_X1 U1350 ( .A1(n1766), .A2(n1767), .ZN(U324) );
NAND2_X1 U1351 ( .A1(n1756), .A2(DATA_IN_3_), .ZN(n1767) );
NAND2_X1 U1352 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1757), .ZN(n1766) );
NAND2_X1 U1353 ( .A1(n1768), .A2(n1769), .ZN(U323) );
NAND2_X1 U1354 ( .A1(n1756), .A2(DATA_IN_2_), .ZN(n1769) );
NAND2_X1 U1355 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1757), .ZN(n1768) );
NAND2_X1 U1356 ( .A1(n1770), .A2(n1771), .ZN(U322) );
NAND2_X1 U1357 ( .A1(n1756), .A2(DATA_IN_1_), .ZN(n1771) );
NAND2_X1 U1358 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1757), .ZN(n1770) );
NAND2_X1 U1359 ( .A1(n1772), .A2(n1773), .ZN(U321) );
NAND2_X1 U1360 ( .A1(n1756), .A2(DATA_IN_0_), .ZN(n1773) );
AND2_X1 U1361 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1774), .ZN(n1756) );
NAND2_X1 U1362 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1757), .ZN(n1772) );
NAND2_X1 U1363 ( .A1(n1636), .A2(n1774), .ZN(n1757) );
NAND2_X1 U1364 ( .A1(n1660), .A2(n1775), .ZN(n1774) );
NAND2_X1 U1365 ( .A1(n1660), .A2(n1776), .ZN(n1636) );
NAND2_X1 U1366 ( .A1(n1777), .A2(n1778), .ZN(U320) );
NAND2_X1 U1367 ( .A1(n1635), .A2(DATA_IN_7_), .ZN(n1778) );
NAND2_X1 U1368 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1779), .ZN(n1777) );
NAND2_X1 U1369 ( .A1(n1780), .A2(n1781), .ZN(U319) );
NAND2_X1 U1370 ( .A1(n1635), .A2(DATA_IN_6_), .ZN(n1781) );
NAND2_X1 U1371 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1779), .ZN(n1780) );
NAND2_X1 U1372 ( .A1(n1782), .A2(n1783), .ZN(U318) );
NAND2_X1 U1373 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1779), .ZN(n1783) );
XOR2_X1 U1374 ( .A(KEYINPUT17), .B(n1784), .Z(n1782) );
NOR2_X1 U1375 ( .A1(n1721), .A2(n1634), .ZN(n1784) );
NAND2_X1 U1376 ( .A1(n1785), .A2(n1786), .ZN(U317) );
NAND2_X1 U1377 ( .A1(n1635), .A2(DATA_IN_4_), .ZN(n1786) );
NAND2_X1 U1378 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1779), .ZN(n1785) );
NAND2_X1 U1379 ( .A1(n1787), .A2(n1788), .ZN(U316) );
NAND2_X1 U1380 ( .A1(n1635), .A2(DATA_IN_3_), .ZN(n1788) );
NAND2_X1 U1381 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1779), .ZN(n1787) );
NAND2_X1 U1382 ( .A1(n1789), .A2(n1790), .ZN(U315) );
NAND2_X1 U1383 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1791), .ZN(n1790) );
XOR2_X1 U1384 ( .A(KEYINPUT48), .B(n1779), .Z(n1791) );
NAND2_X1 U1385 ( .A1(n1635), .A2(DATA_IN_2_), .ZN(n1789) );
NAND2_X1 U1386 ( .A1(n1792), .A2(n1793), .ZN(U314) );
NAND2_X1 U1387 ( .A1(n1635), .A2(DATA_IN_1_), .ZN(n1793) );
NAND2_X1 U1388 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1779), .ZN(n1792) );
NAND2_X1 U1389 ( .A1(n1794), .A2(n1795), .ZN(U313) );
NAND2_X1 U1390 ( .A1(n1635), .A2(DATA_IN_0_), .ZN(n1795) );
NAND2_X1 U1391 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1779), .ZN(n1794) );
NAND2_X1 U1392 ( .A1(n1796), .A2(n1797), .ZN(U312) );
NAND2_X1 U1393 ( .A1(n1798), .A2(n1635), .ZN(n1797) );
XNOR2_X1 U1394 ( .A(REG1_REG_7__SCAN_IN), .B(KEYINPUT41), .ZN(n1798) );
NAND2_X1 U1395 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1779), .ZN(n1796) );
NAND2_X1 U1396 ( .A1(n1799), .A2(n1800), .ZN(U311) );
NAND2_X1 U1397 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1779), .ZN(n1800) );
XOR2_X1 U1398 ( .A(KEYINPUT5), .B(n1801), .Z(n1799) );
AND2_X1 U1399 ( .A1(n1635), .A2(REG1_REG_6__SCAN_IN), .ZN(n1801) );
NAND2_X1 U1400 ( .A1(n1802), .A2(n1803), .ZN(U310) );
NAND2_X1 U1401 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1635), .ZN(n1803) );
NAND2_X1 U1402 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1779), .ZN(n1802) );
NAND2_X1 U1403 ( .A1(n1804), .A2(n1805), .ZN(U309) );
NAND2_X1 U1404 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1635), .ZN(n1805) );
NAND2_X1 U1405 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1779), .ZN(n1804) );
NAND2_X1 U1406 ( .A1(n1806), .A2(n1807), .ZN(U308) );
NAND2_X1 U1407 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1635), .ZN(n1807) );
NAND2_X1 U1408 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1779), .ZN(n1806) );
NAND2_X1 U1409 ( .A1(n1808), .A2(n1809), .ZN(U307) );
NAND2_X1 U1410 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1635), .ZN(n1809) );
NAND2_X1 U1411 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1779), .ZN(n1808) );
NAND2_X1 U1412 ( .A1(n1810), .A2(n1811), .ZN(U306) );
NAND2_X1 U1413 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1635), .ZN(n1811) );
NAND2_X1 U1414 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1779), .ZN(n1810) );
NAND2_X1 U1415 ( .A1(n1812), .A2(n1813), .ZN(U305) );
NAND2_X1 U1416 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1635), .ZN(n1813) );
NAND2_X1 U1417 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1779), .ZN(n1812) );
NAND2_X1 U1418 ( .A1(n1814), .A2(n1815), .ZN(U304) );
NAND2_X1 U1419 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1635), .ZN(n1815) );
NAND2_X1 U1420 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1779), .ZN(n1814) );
NAND2_X1 U1421 ( .A1(n1816), .A2(n1817), .ZN(U303) );
NAND2_X1 U1422 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1635), .ZN(n1817) );
NAND2_X1 U1423 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1779), .ZN(n1816) );
NAND2_X1 U1424 ( .A1(n1818), .A2(n1819), .ZN(U302) );
NAND2_X1 U1425 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1635), .ZN(n1819) );
NAND2_X1 U1426 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1779), .ZN(n1818) );
NAND2_X1 U1427 ( .A1(n1820), .A2(n1821), .ZN(U301) );
NAND2_X1 U1428 ( .A1(n1822), .A2(n1635), .ZN(n1821) );
XNOR2_X1 U1429 ( .A(REG2_REG_4__SCAN_IN), .B(KEYINPUT60), .ZN(n1822) );
NAND2_X1 U1430 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1779), .ZN(n1820) );
NAND2_X1 U1431 ( .A1(n1823), .A2(n1824), .ZN(U300) );
NAND2_X1 U1432 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1825), .ZN(n1824) );
XOR2_X1 U1433 ( .A(KEYINPUT54), .B(n1779), .Z(n1825) );
NAND2_X1 U1434 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1635), .ZN(n1823) );
NAND2_X1 U1435 ( .A1(n1826), .A2(n1827), .ZN(U299) );
NAND2_X1 U1436 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1635), .ZN(n1827) );
XOR2_X1 U1437 ( .A(n1828), .B(KEYINPUT29), .Z(n1826) );
NAND2_X1 U1438 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1779), .ZN(n1828) );
NAND2_X1 U1439 ( .A1(n1829), .A2(n1830), .ZN(U298) );
NAND2_X1 U1440 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1635), .ZN(n1830) );
NAND2_X1 U1441 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1779), .ZN(n1829) );
NAND2_X1 U1442 ( .A1(n1831), .A2(n1832), .ZN(U297) );
NAND2_X1 U1443 ( .A1(n1833), .A2(REG2_REG_0__SCAN_IN), .ZN(n1832) );
XOR2_X1 U1444 ( .A(n1634), .B(KEYINPUT47), .Z(n1833) );
NAND2_X1 U1445 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1779), .ZN(n1831) );
NAND2_X1 U1446 ( .A1(n1834), .A2(n1835), .ZN(U296) );
NAND2_X1 U1447 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1635), .ZN(n1835) );
NAND2_X1 U1448 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1779), .ZN(n1834) );
NAND2_X1 U1449 ( .A1(n1836), .A2(n1837), .ZN(U295) );
NAND2_X1 U1450 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1635), .ZN(n1837) );
NAND2_X1 U1451 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1779), .ZN(n1836) );
NAND2_X1 U1452 ( .A1(n1838), .A2(n1839), .ZN(U294) );
NAND2_X1 U1453 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1779), .ZN(n1839) );
XOR2_X1 U1454 ( .A(KEYINPUT20), .B(n1840), .Z(n1838) );
AND2_X1 U1455 ( .A1(n1635), .A2(REG3_REG_5__SCAN_IN), .ZN(n1840) );
NAND2_X1 U1456 ( .A1(n1841), .A2(n1842), .ZN(U293) );
NAND2_X1 U1457 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1635), .ZN(n1842) );
NAND2_X1 U1458 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1779), .ZN(n1841) );
NAND2_X1 U1459 ( .A1(n1843), .A2(n1844), .ZN(U292) );
NAND2_X1 U1460 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1635), .ZN(n1844) );
NAND2_X1 U1461 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1779), .ZN(n1843) );
NAND2_X1 U1462 ( .A1(n1845), .A2(n1846), .ZN(U291) );
NAND2_X1 U1463 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1847), .ZN(n1846) );
XOR2_X1 U1464 ( .A(KEYINPUT31), .B(n1779), .Z(n1847) );
NAND2_X1 U1465 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1635), .ZN(n1845) );
NAND2_X1 U1466 ( .A1(n1848), .A2(n1849), .ZN(U290) );
NAND2_X1 U1467 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1635), .ZN(n1849) );
NAND2_X1 U1468 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1779), .ZN(n1848) );
NAND2_X1 U1469 ( .A1(n1850), .A2(n1851), .ZN(U289) );
NAND2_X1 U1470 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1635), .ZN(n1851) );
NAND2_X1 U1471 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1779), .ZN(n1850) );
NAND3_X1 U1472 ( .A1(n1852), .A2(n1853), .A3(n1854), .ZN(U288) );
NAND2_X1 U1473 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1779), .ZN(n1854) );
NAND2_X1 U1474 ( .A1(n1855), .A2(REG4_REG_7__SCAN_IN), .ZN(n1853) );
NAND2_X1 U1475 ( .A1(n1856), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1852) );
NAND3_X1 U1476 ( .A1(n1857), .A2(n1858), .A3(n1859), .ZN(U287) );
NOR3_X1 U1477 ( .A1(n1860), .A2(n1861), .A3(n1862), .ZN(n1859) );
NOR4_X1 U1478 ( .A1(n1863), .A2(n1864), .A3(n1865), .A4(n1866), .ZN(n1862));
NOR4_X1 U1479 ( .A1(n1867), .A2(n1868), .A3(n1869), .A4(n1870), .ZN(n1861));
XOR2_X1 U1480 ( .A(KEYINPUT27), .B(n1871), .Z(n1870) );
NOR2_X1 U1481 ( .A1(n1872), .A2(n1873), .ZN(n1860) );
XOR2_X1 U1482 ( .A(RLAST_REG_6__SCAN_IN), .B(KEYINPUT16), .Z(n1873) );
NAND2_X1 U1483 ( .A1(n1855), .A2(REG4_REG_6__SCAN_IN), .ZN(n1858) );
NAND2_X1 U1484 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1779), .ZN(n1857) );
NAND4_X1 U1485 ( .A1(n1874), .A2(n1875), .A3(n1876), .A4(n1877), .ZN(U286));
NOR3_X1 U1486 ( .A1(n1878), .A2(n1879), .A3(n1880), .ZN(n1877) );
NOR2_X1 U1487 ( .A1(n1866), .A2(n1881), .ZN(n1880) );
XNOR2_X1 U1488 ( .A(n1864), .B(n1865), .ZN(n1881) );
NOR2_X1 U1489 ( .A1(n1882), .A2(n1863), .ZN(n1864) );
NOR3_X1 U1490 ( .A1(n1883), .A2(n1884), .A3(n1885), .ZN(n1863) );
AND2_X1 U1491 ( .A1(n1884), .A2(n1886), .ZN(n1882) );
NAND2_X1 U1492 ( .A1(n1887), .A2(n1888), .ZN(n1886) );
NOR2_X1 U1493 ( .A1(n1889), .A2(n1890), .ZN(n1879) );
XNOR2_X1 U1494 ( .A(n1867), .B(n1869), .ZN(n1890) );
NOR2_X1 U1495 ( .A1(n1891), .A2(n1868), .ZN(n1867) );
NOR3_X1 U1496 ( .A1(n1892), .A2(n1884), .A3(n1883), .ZN(n1868) );
AND2_X1 U1497 ( .A1(n1884), .A2(n1893), .ZN(n1891) );
OR2_X1 U1498 ( .A1(n1883), .A2(n1892), .ZN(n1893) );
INV_X1 U1499 ( .A(n1894), .ZN(n1884) );
NOR2_X1 U1500 ( .A1(n1894), .A2(n1895), .ZN(n1878) );
NAND2_X1 U1501 ( .A1(n1896), .A2(n1897), .ZN(n1894) );
NAND3_X1 U1502 ( .A1(n1898), .A2(n1899), .A3(n1900), .ZN(n1897) );
XOR2_X1 U1503 ( .A(n1901), .B(n1902), .Z(n1900) );
NAND2_X1 U1504 ( .A1(n1903), .A2(n1904), .ZN(n1899) );
NAND3_X1 U1505 ( .A1(n1904), .A2(n1905), .A3(n1906), .ZN(n1896) );
XOR2_X1 U1506 ( .A(n1907), .B(n1901), .Z(n1906) );
NAND2_X1 U1507 ( .A1(n1908), .A2(n1909), .ZN(n1901) );
NAND2_X1 U1508 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1910), .ZN(n1909) );
NAND2_X1 U1509 ( .A1(RESTART), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1908) );
NAND2_X1 U1510 ( .A1(KEYINPUT21), .A2(n1902), .ZN(n1907) );
NAND2_X1 U1511 ( .A1(n1911), .A2(n1912), .ZN(n1902) );
NAND2_X1 U1512 ( .A1(RESTART), .A2(n1732), .ZN(n1912) );
NAND2_X1 U1513 ( .A1(n1913), .A2(n1910), .ZN(n1911) );
XOR2_X1 U1514 ( .A(KEYINPUT59), .B(DATA_IN_6_), .Z(n1913) );
NAND2_X1 U1515 ( .A1(n1898), .A2(n1914), .ZN(n1905) );
NAND2_X1 U1516 ( .A1(n1915), .A2(n1916), .ZN(n1898) );
NAND2_X1 U1517 ( .A1(n1917), .A2(n1918), .ZN(n1904) );
NAND2_X1 U1518 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1779), .ZN(n1876) );
NAND2_X1 U1519 ( .A1(n1855), .A2(REG4_REG_5__SCAN_IN), .ZN(n1875) );
NAND2_X1 U1520 ( .A1(n1856), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1874) );
NAND4_X1 U1521 ( .A1(n1919), .A2(n1920), .A3(n1921), .A4(n1922), .ZN(U285));
NOR3_X1 U1522 ( .A1(n1923), .A2(n1924), .A3(n1925), .ZN(n1922) );
NOR2_X1 U1523 ( .A1(n1926), .A2(n1927), .ZN(n1925) );
NOR2_X1 U1524 ( .A1(n1888), .A2(n1895), .ZN(n1924) );
XNOR2_X1 U1525 ( .A(n1928), .B(KEYINPUT49), .ZN(n1923) );
NAND2_X1 U1526 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1779), .ZN(n1928) );
NAND2_X1 U1527 ( .A1(n1929), .A2(RLAST_REG_4__SCAN_IN), .ZN(n1921) );
XOR2_X1 U1528 ( .A(n1872), .B(KEYINPUT53), .Z(n1929) );
NAND3_X1 U1529 ( .A1(n1930), .A2(n1865), .A3(n1931), .ZN(n1920) );
NAND3_X1 U1530 ( .A1(n1932), .A2(n1933), .A3(n1934), .ZN(n1865) );
XOR2_X1 U1531 ( .A(n1888), .B(n1935), .Z(n1932) );
NAND2_X1 U1532 ( .A1(n1936), .A2(n1937), .ZN(n1930) );
NAND2_X1 U1533 ( .A1(n1934), .A2(n1933), .ZN(n1937) );
XOR2_X1 U1534 ( .A(n1883), .B(n1935), .Z(n1936) );
NOR2_X1 U1535 ( .A1(KEYINPUT32), .A2(n1887), .ZN(n1935) );
INV_X1 U1536 ( .A(n1885), .ZN(n1887) );
NAND2_X1 U1537 ( .A1(n1938), .A2(n1871), .ZN(n1919) );
XOR2_X1 U1538 ( .A(n1939), .B(KEYINPUT6), .Z(n1938) );
NAND3_X1 U1539 ( .A1(n1940), .A2(n1941), .A3(n1942), .ZN(n1939) );
XNOR2_X1 U1540 ( .A(KEYINPUT9), .B(n1869), .ZN(n1942) );
OR3_X1 U1541 ( .A1(n1943), .A2(n1944), .A3(n1945), .ZN(n1869) );
NAND2_X1 U1542 ( .A1(n1944), .A2(n1888), .ZN(n1941) );
INV_X1 U1543 ( .A(n1883), .ZN(n1888) );
INV_X1 U1544 ( .A(n1946), .ZN(n1944) );
NAND2_X1 U1545 ( .A1(n1943), .A2(n1945), .ZN(n1940) );
XOR2_X1 U1546 ( .A(n1892), .B(n1883), .Z(n1943) );
NAND2_X1 U1547 ( .A1(n1947), .A2(n1948), .ZN(n1883) );
NAND2_X1 U1548 ( .A1(n1903), .A2(n1949), .ZN(n1948) );
XOR2_X1 U1549 ( .A(n1917), .B(n1950), .Z(n1949) );
NOR2_X1 U1550 ( .A1(n1918), .A2(n1951), .ZN(n1950) );
XOR2_X1 U1551 ( .A(KEYINPUT35), .B(n1952), .Z(n1947) );
NOR2_X1 U1552 ( .A1(n1903), .A2(n1953), .ZN(n1952) );
XOR2_X1 U1553 ( .A(n1954), .B(n1955), .Z(n1953) );
XOR2_X1 U1554 ( .A(KEYINPUT18), .B(n1915), .Z(n1955) );
INV_X1 U1555 ( .A(n1917), .ZN(n1915) );
NAND2_X1 U1556 ( .A1(n1956), .A2(n1957), .ZN(n1917) );
NAND2_X1 U1557 ( .A1(RESTART), .A2(n1701), .ZN(n1957) );
NAND2_X1 U1558 ( .A1(n1958), .A2(n1910), .ZN(n1956) );
NAND2_X1 U1559 ( .A1(n1959), .A2(n1960), .ZN(n1954) );
NAND2_X1 U1560 ( .A1(KEYINPUT30), .A2(n1918), .ZN(n1960) );
NAND2_X1 U1561 ( .A1(n1916), .A2(n1951), .ZN(n1959) );
INV_X1 U1562 ( .A(KEYINPUT10), .ZN(n1951) );
INV_X1 U1563 ( .A(n1918), .ZN(n1916) );
NAND2_X1 U1564 ( .A1(n1961), .A2(n1962), .ZN(n1918) );
NAND2_X1 U1565 ( .A1(RESTART), .A2(n1752), .ZN(n1962) );
INV_X1 U1566 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1752) );
NAND2_X1 U1567 ( .A1(n1721), .A2(n1910), .ZN(n1961) );
INV_X1 U1568 ( .A(n1914), .ZN(n1903) );
NAND2_X1 U1569 ( .A1(n1963), .A2(n1964), .ZN(n1914) );
NAND2_X1 U1570 ( .A1(n1965), .A2(n1966), .ZN(n1964) );
NAND2_X1 U1571 ( .A1(n1967), .A2(n1968), .ZN(n1965) );
OR2_X1 U1572 ( .A1(n1968), .A2(n1967), .ZN(n1963) );
NAND4_X1 U1573 ( .A1(n1969), .A2(n1970), .A3(n1971), .A4(n1972), .ZN(U284));
NAND2_X1 U1574 ( .A1(n1871), .A2(n1973), .ZN(n1972) );
XOR2_X1 U1575 ( .A(n1945), .B(n1974), .Z(n1973) );
NAND2_X1 U1576 ( .A1(KEYINPUT42), .A2(n1946), .ZN(n1974) );
NAND2_X1 U1577 ( .A1(n1975), .A2(n1892), .ZN(n1946) );
NAND2_X1 U1578 ( .A1(n1976), .A2(n1977), .ZN(n1892) );
XNOR2_X1 U1579 ( .A(n1978), .B(KEYINPUT57), .ZN(n1976) );
INV_X1 U1580 ( .A(n1934), .ZN(n1945) );
INV_X1 U1581 ( .A(n1889), .ZN(n1871) );
NAND2_X1 U1582 ( .A1(n1979), .A2(n1931), .ZN(n1971) );
XOR2_X1 U1583 ( .A(n1934), .B(n1933), .Z(n1979) );
NAND2_X1 U1584 ( .A1(n1975), .A2(n1885), .ZN(n1933) );
NAND2_X1 U1585 ( .A1(n1977), .A2(n1978), .ZN(n1885) );
OR2_X1 U1586 ( .A1(n1978), .A2(n1977), .ZN(n1975) );
NAND2_X1 U1587 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1779), .ZN(n1970) );
XOR2_X1 U1588 ( .A(KEYINPUT23), .B(n1980), .Z(n1969) );
NOR3_X1 U1589 ( .A1(n1981), .A2(n1982), .A3(n1983), .ZN(n1980) );
NOR2_X1 U1590 ( .A1(n1984), .A2(n1927), .ZN(n1983) );
AND2_X1 U1591 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1856), .ZN(n1982) );
NOR2_X1 U1592 ( .A1(n1978), .A2(n1895), .ZN(n1981) );
XNOR2_X1 U1593 ( .A(n1985), .B(n1986), .ZN(n1978) );
XOR2_X1 U1594 ( .A(n1968), .B(n1966), .Z(n1986) );
NAND2_X1 U1595 ( .A1(n1987), .A2(n1988), .ZN(n1966) );
NAND2_X1 U1596 ( .A1(n1989), .A2(n1990), .ZN(n1988) );
OR2_X1 U1597 ( .A1(n1991), .A2(n1992), .ZN(n1989) );
NAND2_X1 U1598 ( .A1(n1992), .A2(n1991), .ZN(n1987) );
NAND3_X1 U1599 ( .A1(n1993), .A2(n1994), .A3(n1995), .ZN(n1968) );
NAND2_X1 U1600 ( .A1(KEYINPUT34), .A2(n1720), .ZN(n1995) );
NAND3_X1 U1601 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1996), .A3(RESTART), .ZN(n1994) );
NAND2_X1 U1602 ( .A1(n1997), .A2(n1910), .ZN(n1993) );
NAND2_X1 U1603 ( .A1(n1996), .A2(n1926), .ZN(n1997) );
INV_X1 U1604 ( .A(KEYINPUT34), .ZN(n1996) );
NAND2_X1 U1605 ( .A1(KEYINPUT62), .A2(n1967), .ZN(n1985) );
AND2_X1 U1606 ( .A1(n1998), .A2(n1999), .ZN(n1967) );
NAND2_X1 U1607 ( .A1(RESTART), .A2(n1739), .ZN(n1999) );
NAND2_X1 U1608 ( .A1(n1705), .A2(n1910), .ZN(n1998) );
NAND4_X1 U1609 ( .A1(n2000), .A2(n2001), .A3(n2002), .A4(n2003), .ZN(U283));
NAND2_X1 U1610 ( .A1(n2004), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2003) );
XOR2_X1 U1611 ( .A(n1872), .B(KEYINPUT38), .Z(n2004) );
NOR2_X1 U1612 ( .A1(n2005), .A2(n2006), .ZN(n2002) );
NOR2_X1 U1613 ( .A1(n2007), .A2(n1895), .ZN(n2006) );
XNOR2_X1 U1614 ( .A(KEYINPUT4), .B(n2008), .ZN(n2007) );
NOR2_X1 U1615 ( .A1(n1934), .A2(n2009), .ZN(n2005) );
NOR2_X1 U1616 ( .A1(n2010), .A2(n2011), .ZN(n2009) );
NOR2_X1 U1617 ( .A1(n2012), .A2(n1866), .ZN(n2011) );
NOR2_X1 U1618 ( .A1(n1889), .A2(n2013), .ZN(n2010) );
XOR2_X1 U1619 ( .A(KEYINPUT0), .B(n2012), .Z(n2013) );
AND2_X1 U1620 ( .A1(n2014), .A2(n2015), .ZN(n2012) );
OR2_X1 U1621 ( .A1(n2016), .A2(n2017), .ZN(n2015) );
NOR3_X1 U1622 ( .A1(n2014), .A2(n2017), .A3(n2016), .ZN(n1934) );
NOR2_X1 U1623 ( .A1(n1977), .A2(n2018), .ZN(n2014) );
AND2_X1 U1624 ( .A1(n2008), .A2(n2019), .ZN(n2018) );
NAND2_X1 U1625 ( .A1(n2020), .A2(n2021), .ZN(n2019) );
NOR3_X1 U1626 ( .A1(n2022), .A2(n2008), .A3(n2023), .ZN(n1977) );
XOR2_X1 U1627 ( .A(n2024), .B(n1992), .Z(n2008) );
AND3_X1 U1628 ( .A1(n2025), .A2(n2026), .A3(n2027), .ZN(n1992) );
NAND2_X1 U1629 ( .A1(RESTART), .A2(n2028), .ZN(n2027) );
NAND2_X1 U1630 ( .A1(KEYINPUT56), .A2(n2029), .ZN(n2028) );
XOR2_X1 U1631 ( .A(RMIN_REG_3__SCAN_IN), .B(KEYINPUT61), .Z(n2029) );
NAND3_X1 U1632 ( .A1(KEYINPUT56), .A2(n1910), .A3(REG4_REG_3__SCAN_IN), .ZN(n2026) );
OR2_X1 U1633 ( .A1(KEYINPUT56), .A2(REG4_REG_3__SCAN_IN), .ZN(n2025) );
NAND2_X1 U1634 ( .A1(n2030), .A2(n2031), .ZN(n2024) );
NAND2_X1 U1635 ( .A1(n2032), .A2(n2033), .ZN(n2031) );
NAND2_X1 U1636 ( .A1(KEYINPUT37), .A2(n1991), .ZN(n2033) );
INV_X1 U1637 ( .A(n1990), .ZN(n2032) );
NAND2_X1 U1638 ( .A1(n1991), .A2(n1990), .ZN(n2030) );
NAND2_X1 U1639 ( .A1(n2034), .A2(n2035), .ZN(n1990) );
NAND2_X1 U1640 ( .A1(n2036), .A2(n2037), .ZN(n2035) );
OR2_X1 U1641 ( .A1(n2038), .A2(n2039), .ZN(n2036) );
NAND2_X1 U1642 ( .A1(n2039), .A2(n2038), .ZN(n2034) );
NAND2_X1 U1643 ( .A1(n2040), .A2(n2041), .ZN(n1991) );
NAND2_X1 U1644 ( .A1(RESTART), .A2(n1650), .ZN(n2041) );
NAND2_X1 U1645 ( .A1(n1676), .A2(n1910), .ZN(n2040) );
NAND2_X1 U1646 ( .A1(n1855), .A2(REG4_REG_2__SCAN_IN), .ZN(n2001) );
NAND2_X1 U1647 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1779), .ZN(n2000) );
NAND4_X1 U1648 ( .A1(n2042), .A2(n2043), .A3(n2044), .A4(n2045), .ZN(U282));
NOR3_X1 U1649 ( .A1(n2046), .A2(n2047), .A3(n2048), .ZN(n2045) );
NOR2_X1 U1650 ( .A1(n1889), .A2(n2049), .ZN(n2048) );
NOR2_X1 U1651 ( .A1(n1866), .A2(n2050), .ZN(n2047) );
XOR2_X1 U1652 ( .A(n2049), .B(KEYINPUT3), .Z(n2050) );
XNOR2_X1 U1653 ( .A(n2016), .B(n2017), .ZN(n2049) );
XOR2_X1 U1654 ( .A(n2022), .B(n2023), .Z(n2016) );
NOR2_X1 U1655 ( .A1(n2021), .A2(n1895), .ZN(n2046) );
INV_X1 U1656 ( .A(n2022), .ZN(n2021) );
NAND2_X1 U1657 ( .A1(n2051), .A2(n2052), .ZN(n2022) );
NAND3_X1 U1658 ( .A1(n2053), .A2(n2054), .A3(n2055), .ZN(n2052) );
INV_X1 U1659 ( .A(n2056), .ZN(n2055) );
XOR2_X1 U1660 ( .A(KEYINPUT44), .B(n2039), .Z(n2053) );
NAND2_X1 U1661 ( .A1(n2056), .A2(n2057), .ZN(n2051) );
NAND2_X1 U1662 ( .A1(n2039), .A2(n2058), .ZN(n2057) );
OR2_X1 U1663 ( .A1(n2054), .A2(KEYINPUT44), .ZN(n2058) );
INV_X1 U1664 ( .A(KEYINPUT46), .ZN(n2054) );
AND2_X1 U1665 ( .A1(n2059), .A2(n2060), .ZN(n2039) );
XOR2_X1 U1666 ( .A(n2061), .B(KEYINPUT51), .Z(n2059) );
NAND2_X1 U1667 ( .A1(n2062), .A2(n2063), .ZN(n2061) );
XNOR2_X1 U1668 ( .A(n2037), .B(n2038), .ZN(n2056) );
NAND2_X1 U1669 ( .A1(n2064), .A2(n2065), .ZN(n2038) );
NAND2_X1 U1670 ( .A1(RESTART), .A2(n1716), .ZN(n2065) );
INV_X1 U1671 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1716) );
NAND2_X1 U1672 ( .A1(n2066), .A2(n1910), .ZN(n2064) );
NAND2_X1 U1673 ( .A1(n2067), .A2(n2068), .ZN(n2037) );
NAND2_X1 U1674 ( .A1(n2069), .A2(n1910), .ZN(n2068) );
NAND2_X1 U1675 ( .A1(DATA_IN_2_), .A2(n2070), .ZN(n2069) );
NAND2_X1 U1676 ( .A1(n2071), .A2(n1746), .ZN(n2067) );
NAND2_X1 U1677 ( .A1(DATA_IN_2_), .A2(n2072), .ZN(n2071) );
NAND2_X1 U1678 ( .A1(RESTART), .A2(n2070), .ZN(n2072) );
INV_X1 U1679 ( .A(KEYINPUT13), .ZN(n2070) );
NAND2_X1 U1680 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1779), .ZN(n2044) );
NAND2_X1 U1681 ( .A1(n1855), .A2(REG4_REG_1__SCAN_IN), .ZN(n2043) );
NAND2_X1 U1682 ( .A1(n1856), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2042) );
NAND4_X1 U1683 ( .A1(n2073), .A2(n2074), .A3(n2075), .A4(n2076), .ZN(U281));
NOR2_X1 U1684 ( .A1(n2077), .A2(n2078), .ZN(n2076) );
AND2_X1 U1685 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1856), .ZN(n2078) );
INV_X1 U1686 ( .A(n1872), .ZN(n1856) );
NAND2_X1 U1687 ( .A1(n2079), .A2(n1775), .ZN(n1872) );
INV_X1 U1688 ( .A(ENABLE), .ZN(n1775) );
NOR2_X1 U1689 ( .A1(n2080), .A2(n1895), .ZN(n2077) );
NAND4_X1 U1690 ( .A1(STATO_REG_1__SCAN_IN), .A2(n2081), .A3(n2082), .A4(U280), .ZN(n1895) );
NAND2_X1 U1691 ( .A1(n2083), .A2(n1910), .ZN(n2081) );
NAND3_X1 U1692 ( .A1(n2084), .A2(n2085), .A3(n2086), .ZN(n2083) );
INV_X1 U1693 ( .A(n2087), .ZN(n2080) );
NAND2_X1 U1694 ( .A1(n1855), .A2(REG4_REG_0__SCAN_IN), .ZN(n2075) );
INV_X1 U1695 ( .A(n1927), .ZN(n1855) );
NAND3_X1 U1696 ( .A1(AVERAGE), .A2(n2079), .A3(ENABLE), .ZN(n1927) );
NAND2_X1 U1697 ( .A1(n2088), .A2(DATA_OUT_REG_0__SCAN_IN), .ZN(n2074) );
XOR2_X1 U1698 ( .A(U280), .B(KEYINPUT15), .Z(n2088) );
NAND2_X1 U1699 ( .A1(n2017), .A2(n2089), .ZN(n2073) );
NAND2_X1 U1700 ( .A1(n2090), .A2(n1866), .ZN(n2089) );
INV_X1 U1701 ( .A(n1931), .ZN(n1866) );
NOR3_X1 U1702 ( .A1(n1776), .A2(n1779), .A3(n2082), .ZN(n1931) );
NAND3_X1 U1703 ( .A1(n2091), .A2(n2092), .A3(RESTART), .ZN(n2082) );
NAND2_X1 U1704 ( .A1(n2093), .A2(n1722), .ZN(n2092) );
INV_X1 U1705 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1722) );
OR2_X1 U1706 ( .A1(n2094), .A2(n1728), .ZN(n2093) );
NAND2_X1 U1707 ( .A1(n2094), .A2(n1728), .ZN(n2091) );
INV_X1 U1708 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1728) );
NAND2_X1 U1709 ( .A1(n2095), .A2(n2096), .ZN(n2094) );
NAND2_X1 U1710 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n2097), .ZN(n2096) );
NAND2_X1 U1711 ( .A1(n2098), .A2(n1732), .ZN(n2097) );
INV_X1 U1712 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1732) );
XOR2_X1 U1713 ( .A(KEYINPUT8), .B(n2099), .Z(n2098) );
NAND2_X1 U1714 ( .A1(n2099), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2095) );
AND2_X1 U1715 ( .A1(n2100), .A2(n2101), .ZN(n2099) );
NAND2_X1 U1716 ( .A1(n1701), .A2(n2102), .ZN(n2101) );
NAND2_X1 U1717 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n2103), .ZN(n2102) );
INV_X1 U1718 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1701) );
OR2_X1 U1719 ( .A1(n2103), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2100) );
NAND2_X1 U1720 ( .A1(n2104), .A2(n2105), .ZN(n2103) );
NAND2_X1 U1721 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2105) );
NAND3_X1 U1722 ( .A1(n2106), .A2(n2107), .A3(n2108), .ZN(n2104) );
NAND2_X1 U1723 ( .A1(n1739), .A2(n1720), .ZN(n2108) );
INV_X1 U1724 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1720) );
INV_X1 U1725 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1739) );
NAND3_X1 U1726 ( .A1(n2109), .A2(n2110), .A3(n2111), .ZN(n2107) );
NAND2_X1 U1727 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2111) );
NAND3_X1 U1728 ( .A1(n2112), .A2(n2113), .A3(n2114), .ZN(n2110) );
XOR2_X1 U1729 ( .A(KEYINPUT45), .B(n2115), .Z(n2114) );
NOR2_X1 U1730 ( .A1(n2116), .A2(n2117), .ZN(n2115) );
NOR2_X1 U1731 ( .A1(n1751), .A2(n1719), .ZN(n2117) );
NAND2_X1 U1732 ( .A1(n2118), .A2(n1746), .ZN(n2113) );
INV_X1 U1733 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1746) );
XOR2_X1 U1734 ( .A(RMIN_REG_2__SCAN_IN), .B(KEYINPUT24), .Z(n2118) );
NAND2_X1 U1735 ( .A1(n1751), .A2(n1719), .ZN(n2112) );
INV_X1 U1736 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1719) );
NAND2_X1 U1737 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2109) );
NAND2_X1 U1738 ( .A1(n1650), .A2(n1709), .ZN(n2106) );
INV_X1 U1739 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1709) );
INV_X1 U1740 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1650) );
XOR2_X1 U1741 ( .A(n1889), .B(KEYINPUT7), .Z(n2090) );
NAND3_X1 U1742 ( .A1(n2079), .A2(n2119), .A3(n2086), .ZN(n1889) );
AND2_X1 U1743 ( .A1(ENABLE), .A2(n2120), .ZN(n2086) );
XOR2_X1 U1744 ( .A(KEYINPUT52), .B(AVERAGE), .Z(n2120) );
NAND2_X1 U1745 ( .A1(n2084), .A2(n2085), .ZN(n2119) );
NAND3_X1 U1746 ( .A1(n2121), .A2(n2122), .A3(n2123), .ZN(n2085) );
OR2_X1 U1747 ( .A1(DATA_IN_7_), .A2(REG4_REG_7__SCAN_IN), .ZN(n2123) );
NAND3_X1 U1748 ( .A1(n2124), .A2(n2125), .A3(n2126), .ZN(n2122) );
OR2_X1 U1749 ( .A1(DATA_IN_6_), .A2(REG4_REG_6__SCAN_IN), .ZN(n2126) );
NAND3_X1 U1750 ( .A1(n2127), .A2(n2128), .A3(n2129), .ZN(n2125) );
NAND2_X1 U1751 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2129) );
NAND3_X1 U1752 ( .A1(n2130), .A2(n2131), .A3(n2132), .ZN(n2128) );
NAND2_X1 U1753 ( .A1(n1705), .A2(n1926), .ZN(n2132) );
INV_X1 U1754 ( .A(REG4_REG_4__SCAN_IN), .ZN(n1926) );
INV_X1 U1755 ( .A(DATA_IN_4_), .ZN(n1705) );
NAND3_X1 U1756 ( .A1(n2133), .A2(n2134), .A3(n2135), .ZN(n2131) );
NAND2_X1 U1757 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2135) );
NAND3_X1 U1758 ( .A1(n2136), .A2(n2137), .A3(n2138), .ZN(n2134) );
NAND2_X1 U1759 ( .A1(n1680), .A2(n2066), .ZN(n2138) );
INV_X1 U1760 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2066) );
INV_X1 U1761 ( .A(DATA_IN_2_), .ZN(n1680) );
NAND2_X1 U1762 ( .A1(n2139), .A2(n2140), .ZN(n2137) );
XOR2_X1 U1763 ( .A(KEYINPUT43), .B(n2141), .Z(n2139) );
NOR2_X1 U1764 ( .A1(n1713), .A2(n2142), .ZN(n2141) );
NAND2_X1 U1765 ( .A1(n1713), .A2(n2142), .ZN(n2136) );
INV_X1 U1766 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2142) );
INV_X1 U1767 ( .A(DATA_IN_1_), .ZN(n1713) );
NAND2_X1 U1768 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2133) );
NAND2_X1 U1769 ( .A1(n1676), .A2(n1984), .ZN(n2130) );
INV_X1 U1770 ( .A(REG4_REG_3__SCAN_IN), .ZN(n1984) );
INV_X1 U1771 ( .A(DATA_IN_3_), .ZN(n1676) );
NAND2_X1 U1772 ( .A1(REG4_REG_5__SCAN_IN), .A2(n2143), .ZN(n2127) );
XOR2_X1 U1773 ( .A(KEYINPUT1), .B(DATA_IN_5_), .Z(n2143) );
NAND2_X1 U1774 ( .A1(n1721), .A2(n1958), .ZN(n2124) );
INV_X1 U1775 ( .A(REG4_REG_5__SCAN_IN), .ZN(n1958) );
INV_X1 U1776 ( .A(DATA_IN_5_), .ZN(n1721) );
NAND2_X1 U1777 ( .A1(REG4_REG_6__SCAN_IN), .A2(DATA_IN_6_), .ZN(n2121) );
NAND2_X1 U1778 ( .A1(REG4_REG_7__SCAN_IN), .A2(DATA_IN_7_), .ZN(n2084) );
NOR3_X1 U1779 ( .A1(n1779), .A2(RESTART), .A3(n1776), .ZN(n2079) );
AND2_X1 U1780 ( .A1(n2023), .A2(n2144), .ZN(n2017) );
NAND2_X1 U1781 ( .A1(n2145), .A2(n2087), .ZN(n2144) );
INV_X1 U1782 ( .A(n2020), .ZN(n2023) );
NOR2_X1 U1783 ( .A1(n2087), .A2(n2145), .ZN(n2020) );
AND3_X1 U1784 ( .A1(n2146), .A2(n2147), .A3(n2148), .ZN(n2145) );
OR3_X1 U1785 ( .A1(DATA_IN_0_), .A2(REG4_REG_0__SCAN_IN), .A3(RESTART), .ZN(n2147) );
NAND3_X1 U1786 ( .A1(n1748), .A2(n2149), .A3(RESTART), .ZN(n2146) );
NAND2_X1 U1787 ( .A1(n2150), .A2(n2151), .ZN(n2087) );
NAND2_X1 U1788 ( .A1(n2062), .A2(n2152), .ZN(n2151) );
NAND2_X1 U1789 ( .A1(n2063), .A2(n2060), .ZN(n2152) );
NAND2_X1 U1790 ( .A1(n2153), .A2(n2154), .ZN(n2060) );
INV_X1 U1791 ( .A(n2155), .ZN(n2154) );
INV_X1 U1792 ( .A(n2148), .ZN(n2153) );
NAND2_X1 U1793 ( .A1(n2155), .A2(n2148), .ZN(n2063) );
NAND2_X1 U1794 ( .A1(n2156), .A2(n2157), .ZN(n2150) );
INV_X1 U1795 ( .A(n2062), .ZN(n2157) );
NAND2_X1 U1796 ( .A1(n2158), .A2(n2159), .ZN(n2062) );
NAND2_X1 U1797 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1910), .ZN(n2159) );
NAND2_X1 U1798 ( .A1(RESTART), .A2(RMIN_REG_1__SCAN_IN), .ZN(n2158) );
XOR2_X1 U1799 ( .A(n2148), .B(n2155), .Z(n2156) );
NAND2_X1 U1800 ( .A1(n2160), .A2(n2161), .ZN(n2155) );
NAND2_X1 U1801 ( .A1(RESTART), .A2(n1751), .ZN(n2161) );
INV_X1 U1802 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1751) );
NAND2_X1 U1803 ( .A1(n2162), .A2(n1910), .ZN(n2160) );
XOR2_X1 U1804 ( .A(KEYINPUT22), .B(DATA_IN_1_), .Z(n2162) );
NAND2_X1 U1805 ( .A1(n2163), .A2(n2164), .ZN(n2148) );
OR2_X1 U1806 ( .A1(n1910), .A2(n2116), .ZN(n2164) );
NOR2_X1 U1807 ( .A1(n2149), .A2(n1748), .ZN(n2116) );
INV_X1 U1808 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1748) );
INV_X1 U1809 ( .A(RMIN_REG_0__SCAN_IN), .ZN(n2149) );
NAND2_X1 U1810 ( .A1(n2140), .A2(n1910), .ZN(n2163) );
INV_X1 U1811 ( .A(RESTART), .ZN(n1910) );
NAND2_X1 U1812 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2140) );
NAND2_X1 U1813 ( .A1(n2165), .A2(n1634), .ZN(U280) );
XOR2_X1 U1814 ( .A(KEYINPUT11), .B(n2166), .Z(n2165) );
NOR2_X1 U1815 ( .A1(n2167), .A2(n1660), .ZN(n2166) );
INV_X1 U1816 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1660) );
XOR2_X1 U1817 ( .A(n1776), .B(KEYINPUT19), .Z(n2167) );
INV_X1 U1818 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1776) );
endmodule


