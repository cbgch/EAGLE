//Key = 0110001011001100101001010011100101010000001011011001010100110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322;

XNOR2_X1 U735 ( .A(G107), .B(n1005), .ZN(G9) );
NAND4_X1 U736 ( .A1(KEYINPUT6), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1005) );
NOR2_X1 U737 ( .A1(n1009), .A2(n1010), .ZN(G75) );
XOR2_X1 U738 ( .A(n1011), .B(KEYINPUT47), .Z(n1010) );
NAND3_X1 U739 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1011) );
NAND2_X1 U740 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NAND2_X1 U741 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND3_X1 U742 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NAND2_X1 U743 ( .A1(n1022), .A2(n1023), .ZN(n1019) );
NAND3_X1 U744 ( .A1(n1007), .A2(n1024), .A3(n1025), .ZN(n1023) );
NAND2_X1 U745 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NAND2_X1 U746 ( .A1(n1028), .A2(n1029), .ZN(n1022) );
NAND2_X1 U747 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U748 ( .A1(n1025), .A2(n1032), .ZN(n1031) );
OR2_X1 U749 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U750 ( .A1(n1007), .A2(n1035), .ZN(n1030) );
NAND2_X1 U751 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U752 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NAND4_X1 U753 ( .A1(n1041), .A2(n1042), .A3(n1028), .A4(n1043), .ZN(n1017) );
NOR2_X1 U754 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U755 ( .A1(n1025), .A2(n1046), .ZN(n1044) );
NAND2_X1 U756 ( .A1(n1047), .A2(n1020), .ZN(n1042) );
NAND2_X1 U757 ( .A1(n1025), .A2(n1048), .ZN(n1047) );
NAND2_X1 U758 ( .A1(n1021), .A2(n1039), .ZN(n1048) );
INV_X1 U759 ( .A(KEYINPUT29), .ZN(n1039) );
NAND2_X1 U760 ( .A1(n1049), .A2(n1050), .ZN(n1041) );
NAND2_X1 U761 ( .A1(n1021), .A2(n1051), .ZN(n1050) );
NAND2_X1 U762 ( .A1(n1025), .A2(n1046), .ZN(n1051) );
INV_X1 U763 ( .A(KEYINPUT45), .ZN(n1046) );
INV_X1 U764 ( .A(n1052), .ZN(n1025) );
INV_X1 U765 ( .A(n1053), .ZN(n1015) );
INV_X1 U766 ( .A(n1054), .ZN(n1012) );
NOR2_X1 U767 ( .A1(G952), .A2(n1054), .ZN(n1009) );
NAND2_X1 U768 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND4_X1 U769 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
NOR4_X1 U770 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1060) );
NOR2_X1 U771 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U772 ( .A1(KEYINPUT25), .A2(n1067), .ZN(n1065) );
XOR2_X1 U773 ( .A(n1068), .B(KEYINPUT52), .Z(n1067) );
NOR3_X1 U774 ( .A1(G469), .A2(KEYINPUT25), .A3(n1068), .ZN(n1063) );
XOR2_X1 U775 ( .A(KEYINPUT39), .B(n1069), .Z(n1062) );
NAND3_X1 U776 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1061) );
XOR2_X1 U777 ( .A(n1038), .B(KEYINPUT20), .Z(n1072) );
NAND2_X1 U778 ( .A1(KEYINPUT25), .A2(n1068), .ZN(n1071) );
NOR3_X1 U779 ( .A1(n1073), .A2(n1040), .A3(n1049), .ZN(n1059) );
NOR2_X1 U780 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XOR2_X1 U781 ( .A(n1076), .B(KEYINPUT32), .Z(n1075) );
XOR2_X1 U782 ( .A(n1077), .B(n1078), .Z(n1057) );
NAND2_X1 U783 ( .A1(KEYINPUT2), .A2(n1079), .ZN(n1078) );
XOR2_X1 U784 ( .A(n1080), .B(n1081), .Z(G72) );
NOR2_X1 U785 ( .A1(n1082), .A2(n1055), .ZN(n1081) );
NOR2_X1 U786 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U787 ( .A1(n1085), .A2(n1086), .ZN(n1080) );
NAND2_X1 U788 ( .A1(n1087), .A2(n1055), .ZN(n1086) );
XOR2_X1 U789 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U790 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
XOR2_X1 U791 ( .A(KEYINPUT17), .B(n1092), .Z(n1091) );
NOR2_X1 U792 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U793 ( .A(KEYINPUT56), .B(n1095), .Z(n1094) );
INV_X1 U794 ( .A(n1096), .ZN(n1090) );
NAND3_X1 U795 ( .A1(G900), .A2(n1089), .A3(G953), .ZN(n1085) );
XOR2_X1 U796 ( .A(n1097), .B(n1098), .Z(n1089) );
XNOR2_X1 U797 ( .A(n1099), .B(n1100), .ZN(n1098) );
NAND2_X1 U798 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
OR2_X1 U799 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XOR2_X1 U800 ( .A(n1105), .B(KEYINPUT0), .Z(n1101) );
NAND2_X1 U801 ( .A1(n1104), .A2(n1103), .ZN(n1105) );
XOR2_X1 U802 ( .A(G134), .B(G137), .Z(n1103) );
XOR2_X1 U803 ( .A(n1106), .B(n1107), .Z(n1097) );
NOR2_X1 U804 ( .A1(KEYINPUT22), .A2(n1108), .ZN(n1107) );
XOR2_X1 U805 ( .A(n1109), .B(n1110), .Z(n1108) );
XOR2_X1 U806 ( .A(KEYINPUT31), .B(G140), .Z(n1110) );
XOR2_X1 U807 ( .A(n1111), .B(n1112), .Z(G69) );
XOR2_X1 U808 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U809 ( .A1(n1115), .A2(n1055), .ZN(n1114) );
AND2_X1 U810 ( .A1(G224), .A2(G898), .ZN(n1115) );
NAND2_X1 U811 ( .A1(n1116), .A2(n1117), .ZN(n1113) );
NAND2_X1 U812 ( .A1(G953), .A2(n1118), .ZN(n1117) );
XNOR2_X1 U813 ( .A(n1119), .B(n1120), .ZN(n1116) );
NAND2_X1 U814 ( .A1(n1055), .A2(n1121), .ZN(n1111) );
NOR2_X1 U815 ( .A1(n1122), .A2(n1123), .ZN(G66) );
XNOR2_X1 U816 ( .A(n1124), .B(KEYINPUT58), .ZN(n1123) );
NOR3_X1 U817 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1122) );
NOR3_X1 U818 ( .A1(n1128), .A2(n1077), .A3(n1129), .ZN(n1127) );
NOR2_X1 U819 ( .A1(n1130), .A2(n1131), .ZN(n1126) );
NOR2_X1 U820 ( .A1(n1014), .A2(n1077), .ZN(n1130) );
INV_X1 U821 ( .A(n1079), .ZN(n1125) );
NOR2_X1 U822 ( .A1(n1124), .A2(n1132), .ZN(G63) );
XOR2_X1 U823 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U824 ( .A1(n1076), .A2(n1129), .ZN(n1134) );
NOR3_X1 U825 ( .A1(n1124), .A2(n1135), .A3(n1136), .ZN(G60) );
NOR4_X1 U826 ( .A1(n1137), .A2(n1129), .A3(KEYINPUT50), .A4(n1138), .ZN(n1136) );
NOR2_X1 U827 ( .A1(n1139), .A2(n1140), .ZN(n1135) );
NOR3_X1 U828 ( .A1(n1129), .A2(n1141), .A3(n1138), .ZN(n1140) );
INV_X1 U829 ( .A(G475), .ZN(n1138) );
NOR2_X1 U830 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
INV_X1 U831 ( .A(KEYINPUT50), .ZN(n1143) );
INV_X1 U832 ( .A(n1137), .ZN(n1139) );
NAND2_X1 U833 ( .A1(KEYINPUT26), .A2(n1142), .ZN(n1137) );
XOR2_X1 U834 ( .A(G104), .B(n1144), .Z(G6) );
NOR2_X1 U835 ( .A1(n1124), .A2(n1145), .ZN(G57) );
XOR2_X1 U836 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U837 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U838 ( .A(n1150), .B(n1151), .Z(n1146) );
XOR2_X1 U839 ( .A(KEYINPUT34), .B(n1152), .Z(n1151) );
NOR2_X1 U840 ( .A1(n1153), .A2(n1129), .ZN(n1150) );
INV_X1 U841 ( .A(G472), .ZN(n1153) );
NOR2_X1 U842 ( .A1(n1124), .A2(n1154), .ZN(G54) );
XOR2_X1 U843 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U844 ( .A(KEYINPUT24), .B(n1157), .Z(n1156) );
NOR2_X1 U845 ( .A1(n1066), .A2(n1129), .ZN(n1157) );
NOR2_X1 U846 ( .A1(n1055), .A2(G952), .ZN(n1124) );
NOR2_X1 U847 ( .A1(n1158), .A2(n1159), .ZN(G51) );
XOR2_X1 U848 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U849 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U850 ( .A1(n1164), .A2(n1129), .ZN(n1163) );
OR2_X1 U851 ( .A1(n1165), .A2(n1014), .ZN(n1129) );
NOR4_X1 U852 ( .A1(n1121), .A2(n1096), .A3(n1093), .A4(n1095), .ZN(n1014) );
NAND3_X1 U853 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1093) );
NAND2_X1 U854 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
XOR2_X1 U855 ( .A(n1171), .B(KEYINPUT42), .Z(n1169) );
NAND3_X1 U856 ( .A1(n1172), .A2(n1173), .A3(n1028), .ZN(n1166) );
XOR2_X1 U857 ( .A(KEYINPUT40), .B(n1174), .Z(n1173) );
NAND4_X1 U858 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1096) );
NAND4_X1 U859 ( .A1(n1179), .A2(n1174), .A3(n1180), .A4(n1008), .ZN(n1176) );
XOR2_X1 U860 ( .A(n1036), .B(KEYINPUT21), .Z(n1179) );
NAND3_X1 U861 ( .A1(n1181), .A2(n1172), .A3(n1033), .ZN(n1175) );
OR4_X1 U862 ( .A1(n1144), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1121) );
OR4_X1 U863 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1184) );
AND2_X1 U864 ( .A1(n1008), .A2(n1189), .ZN(n1183) );
NAND2_X1 U865 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND3_X1 U866 ( .A1(n1192), .A2(n1193), .A3(n1007), .ZN(n1191) );
OR2_X1 U867 ( .A1(n1006), .A2(KEYINPUT3), .ZN(n1193) );
NAND2_X1 U868 ( .A1(KEYINPUT3), .A2(n1194), .ZN(n1192) );
NAND3_X1 U869 ( .A1(n1036), .A2(n1195), .A3(n1196), .ZN(n1194) );
NAND3_X1 U870 ( .A1(n1197), .A2(n1198), .A3(n1033), .ZN(n1190) );
NAND2_X1 U871 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
INV_X1 U872 ( .A(KEYINPUT49), .ZN(n1200) );
NAND2_X1 U873 ( .A1(KEYINPUT49), .A2(n1201), .ZN(n1197) );
NAND2_X1 U874 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
INV_X1 U875 ( .A(n1195), .ZN(n1202) );
NOR3_X1 U876 ( .A1(n1204), .A2(n1045), .A3(n1026), .ZN(n1144) );
NAND2_X1 U877 ( .A1(n1205), .A2(n1206), .ZN(n1162) );
NAND2_X1 U878 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
INV_X1 U879 ( .A(n1209), .ZN(n1205) );
NOR2_X1 U880 ( .A1(n1210), .A2(n1055), .ZN(n1158) );
XNOR2_X1 U881 ( .A(G952), .B(KEYINPUT1), .ZN(n1210) );
XOR2_X1 U882 ( .A(n1106), .B(n1167), .Z(G48) );
NAND4_X1 U883 ( .A1(n1174), .A2(n1181), .A3(n1180), .A4(n1170), .ZN(n1167) );
XOR2_X1 U884 ( .A(G143), .B(n1211), .Z(G45) );
NOR2_X1 U885 ( .A1(n1036), .A2(n1171), .ZN(n1211) );
NAND4_X1 U886 ( .A1(n1033), .A2(n1180), .A3(n1212), .A4(n1213), .ZN(n1171) );
INV_X1 U887 ( .A(n1214), .ZN(n1180) );
XOR2_X1 U888 ( .A(G140), .B(n1095), .Z(G42) );
AND3_X1 U889 ( .A1(n1172), .A2(n1034), .A3(n1181), .ZN(n1095) );
XNOR2_X1 U890 ( .A(G137), .B(n1215), .ZN(G39) );
NAND3_X1 U891 ( .A1(n1174), .A2(n1172), .A3(n1216), .ZN(n1215) );
XOR2_X1 U892 ( .A(n1217), .B(KEYINPUT9), .Z(n1216) );
INV_X1 U893 ( .A(n1218), .ZN(n1174) );
XOR2_X1 U894 ( .A(n1219), .B(n1177), .Z(G36) );
NAND3_X1 U895 ( .A1(n1172), .A2(n1008), .A3(n1033), .ZN(n1177) );
INV_X1 U896 ( .A(n1220), .ZN(n1033) );
INV_X1 U897 ( .A(n1027), .ZN(n1008) );
NOR2_X1 U898 ( .A1(n1214), .A2(n1052), .ZN(n1172) );
XOR2_X1 U899 ( .A(G131), .B(n1221), .Z(G33) );
NOR4_X1 U900 ( .A1(n1222), .A2(n1214), .A3(n1026), .A4(n1220), .ZN(n1221) );
XOR2_X1 U901 ( .A(n1052), .B(KEYINPUT14), .Z(n1222) );
NAND2_X1 U902 ( .A1(n1038), .A2(n1223), .ZN(n1052) );
XOR2_X1 U903 ( .A(G128), .B(n1224), .Z(G30) );
NOR4_X1 U904 ( .A1(n1036), .A2(n1027), .A3(n1214), .A4(n1218), .ZN(n1224) );
NAND2_X1 U905 ( .A1(n1196), .A2(n1225), .ZN(n1214) );
INV_X1 U906 ( .A(n1170), .ZN(n1036) );
XOR2_X1 U907 ( .A(G101), .B(n1182), .Z(G3) );
NOR3_X1 U908 ( .A1(n1217), .A2(n1204), .A3(n1220), .ZN(n1182) );
XOR2_X1 U909 ( .A(n1109), .B(n1178), .Z(G27) );
NAND4_X1 U910 ( .A1(n1203), .A2(n1181), .A3(n1034), .A4(n1225), .ZN(n1178) );
NAND2_X1 U911 ( .A1(n1053), .A2(n1226), .ZN(n1225) );
NAND4_X1 U912 ( .A1(G953), .A2(G902), .A3(n1227), .A4(n1084), .ZN(n1226) );
INV_X1 U913 ( .A(G900), .ZN(n1084) );
INV_X1 U914 ( .A(n1026), .ZN(n1181) );
XNOR2_X1 U915 ( .A(n1188), .B(n1228), .ZN(G24) );
NAND2_X1 U916 ( .A1(KEYINPUT53), .A2(G122), .ZN(n1228) );
NOR4_X1 U917 ( .A1(n1199), .A2(n1045), .A3(n1229), .A4(n1230), .ZN(n1188) );
INV_X1 U918 ( .A(n1007), .ZN(n1045) );
NOR2_X1 U919 ( .A1(n1231), .A2(n1232), .ZN(n1007) );
XOR2_X1 U920 ( .A(G119), .B(n1187), .Z(G21) );
NOR3_X1 U921 ( .A1(n1199), .A2(n1217), .A3(n1218), .ZN(n1187) );
NAND2_X1 U922 ( .A1(n1232), .A2(n1231), .ZN(n1218) );
XOR2_X1 U923 ( .A(G116), .B(n1233), .Z(G18) );
NOR4_X1 U924 ( .A1(KEYINPUT4), .A2(n1027), .A3(n1199), .A4(n1220), .ZN(n1233) );
NAND2_X1 U925 ( .A1(n1234), .A2(n1213), .ZN(n1027) );
INV_X1 U926 ( .A(n1230), .ZN(n1213) );
XOR2_X1 U927 ( .A(KEYINPUT27), .B(n1212), .Z(n1234) );
XOR2_X1 U928 ( .A(G113), .B(n1186), .Z(G15) );
NOR3_X1 U929 ( .A1(n1199), .A2(n1026), .A3(n1220), .ZN(n1186) );
NAND2_X1 U930 ( .A1(n1231), .A2(n1235), .ZN(n1220) );
NAND2_X1 U931 ( .A1(n1230), .A2(n1212), .ZN(n1026) );
INV_X1 U932 ( .A(n1229), .ZN(n1212) );
NAND2_X1 U933 ( .A1(n1203), .A2(n1195), .ZN(n1199) );
AND3_X1 U934 ( .A1(n1021), .A2(n1020), .A3(n1170), .ZN(n1203) );
XOR2_X1 U935 ( .A(G110), .B(n1185), .Z(G12) );
AND3_X1 U936 ( .A1(n1034), .A2(n1006), .A3(n1028), .ZN(n1185) );
INV_X1 U937 ( .A(n1217), .ZN(n1028) );
NAND2_X1 U938 ( .A1(n1230), .A2(n1229), .ZN(n1217) );
XOR2_X1 U939 ( .A(n1070), .B(KEYINPUT62), .Z(n1229) );
XOR2_X1 U940 ( .A(n1236), .B(G475), .Z(n1070) );
NAND2_X1 U941 ( .A1(n1142), .A2(n1165), .ZN(n1236) );
XNOR2_X1 U942 ( .A(n1237), .B(n1238), .ZN(n1142) );
XOR2_X1 U943 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U944 ( .A(n1241), .B(n1242), .Z(n1240) );
NOR2_X1 U945 ( .A1(G143), .A2(KEYINPUT10), .ZN(n1242) );
AND3_X1 U946 ( .A1(G214), .A2(n1055), .A3(n1243), .ZN(n1241) );
XOR2_X1 U947 ( .A(n1244), .B(n1245), .Z(n1237) );
XOR2_X1 U948 ( .A(G131), .B(G125), .Z(n1245) );
XOR2_X1 U949 ( .A(n1246), .B(G104), .Z(n1244) );
NAND2_X1 U950 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND2_X1 U951 ( .A1(n1249), .A2(G113), .ZN(n1248) );
XOR2_X1 U952 ( .A(KEYINPUT12), .B(n1250), .Z(n1247) );
NOR2_X1 U953 ( .A1(G113), .A2(n1249), .ZN(n1250) );
NOR2_X1 U954 ( .A1(n1069), .A2(n1251), .ZN(n1230) );
NOR2_X1 U955 ( .A1(n1076), .A2(n1074), .ZN(n1251) );
AND2_X1 U956 ( .A1(n1074), .A2(n1076), .ZN(n1069) );
INV_X1 U957 ( .A(G478), .ZN(n1076) );
NOR2_X1 U958 ( .A1(n1133), .A2(G902), .ZN(n1074) );
XOR2_X1 U959 ( .A(n1252), .B(n1253), .Z(n1133) );
XOR2_X1 U960 ( .A(G128), .B(n1254), .Z(n1253) );
XOR2_X1 U961 ( .A(G143), .B(G134), .Z(n1254) );
XOR2_X1 U962 ( .A(n1255), .B(n1256), .Z(n1252) );
AND3_X1 U963 ( .A1(G217), .A2(n1055), .A3(G234), .ZN(n1256) );
XNOR2_X1 U964 ( .A(G107), .B(n1257), .ZN(n1255) );
NOR2_X1 U965 ( .A1(KEYINPUT15), .A2(n1258), .ZN(n1257) );
XOR2_X1 U966 ( .A(n1259), .B(n1249), .Z(n1258) );
NAND2_X1 U967 ( .A1(KEYINPUT33), .A2(n1260), .ZN(n1259) );
INV_X1 U968 ( .A(G116), .ZN(n1260) );
INV_X1 U969 ( .A(n1204), .ZN(n1006) );
NAND3_X1 U970 ( .A1(n1196), .A2(n1195), .A3(n1170), .ZN(n1204) );
NOR2_X1 U971 ( .A1(n1038), .A2(n1040), .ZN(n1170) );
INV_X1 U972 ( .A(n1223), .ZN(n1040) );
NAND2_X1 U973 ( .A1(G214), .A2(n1261), .ZN(n1223) );
XNOR2_X1 U974 ( .A(n1262), .B(n1164), .ZN(n1038) );
NAND2_X1 U975 ( .A1(G210), .A2(n1261), .ZN(n1164) );
NAND2_X1 U976 ( .A1(n1243), .A2(n1165), .ZN(n1261) );
INV_X1 U977 ( .A(G237), .ZN(n1243) );
NAND2_X1 U978 ( .A1(n1263), .A2(n1165), .ZN(n1262) );
XOR2_X1 U979 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U980 ( .A(KEYINPUT18), .B(n1266), .Z(n1265) );
NOR2_X1 U981 ( .A1(n1267), .A2(n1209), .ZN(n1266) );
NOR2_X1 U982 ( .A1(n1208), .A2(n1207), .ZN(n1209) );
NAND2_X1 U983 ( .A1(G224), .A2(n1055), .ZN(n1208) );
NOR2_X1 U984 ( .A1(G224), .A2(n1268), .ZN(n1267) );
XNOR2_X1 U985 ( .A(KEYINPUT7), .B(n1207), .ZN(n1268) );
XNOR2_X1 U986 ( .A(n1269), .B(n1109), .ZN(n1207) );
INV_X1 U987 ( .A(G125), .ZN(n1109) );
INV_X1 U988 ( .A(n1160), .ZN(n1264) );
XOR2_X1 U989 ( .A(n1270), .B(n1120), .Z(n1160) );
XNOR2_X1 U990 ( .A(G110), .B(n1249), .ZN(n1120) );
XNOR2_X1 U991 ( .A(G122), .B(KEYINPUT30), .ZN(n1249) );
NAND2_X1 U992 ( .A1(KEYINPUT63), .A2(n1119), .ZN(n1270) );
XNOR2_X1 U993 ( .A(n1271), .B(n1272), .ZN(n1119) );
XOR2_X1 U994 ( .A(n1273), .B(n1274), .Z(n1272) );
NOR2_X1 U995 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
XOR2_X1 U996 ( .A(KEYINPUT57), .B(n1277), .Z(n1276) );
NOR2_X1 U997 ( .A1(G113), .A2(n1278), .ZN(n1277) );
AND2_X1 U998 ( .A1(n1278), .A2(G113), .ZN(n1275) );
NAND2_X1 U999 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND2_X1 U1000 ( .A1(G116), .A2(n1281), .ZN(n1280) );
XOR2_X1 U1001 ( .A(KEYINPUT48), .B(n1282), .Z(n1279) );
NOR2_X1 U1002 ( .A1(G116), .A2(n1281), .ZN(n1282) );
INV_X1 U1003 ( .A(G119), .ZN(n1281) );
XOR2_X1 U1004 ( .A(n1283), .B(n1284), .Z(n1271) );
NOR2_X1 U1005 ( .A1(G101), .A2(KEYINPUT46), .ZN(n1284) );
XNOR2_X1 U1006 ( .A(KEYINPUT55), .B(KEYINPUT37), .ZN(n1283) );
NAND2_X1 U1007 ( .A1(n1285), .A2(n1053), .ZN(n1195) );
NAND3_X1 U1008 ( .A1(n1227), .A2(n1055), .A3(G952), .ZN(n1053) );
NAND4_X1 U1009 ( .A1(G953), .A2(G902), .A3(n1227), .A4(n1118), .ZN(n1285) );
INV_X1 U1010 ( .A(G898), .ZN(n1118) );
NAND2_X1 U1011 ( .A1(G237), .A2(G234), .ZN(n1227) );
NOR2_X1 U1012 ( .A1(n1021), .A2(n1049), .ZN(n1196) );
INV_X1 U1013 ( .A(n1020), .ZN(n1049) );
NAND2_X1 U1014 ( .A1(G221), .A2(n1286), .ZN(n1020) );
XOR2_X1 U1015 ( .A(n1287), .B(n1068), .Z(n1021) );
NAND2_X1 U1016 ( .A1(n1288), .A2(n1165), .ZN(n1068) );
XNOR2_X1 U1017 ( .A(n1155), .B(KEYINPUT60), .ZN(n1288) );
XNOR2_X1 U1018 ( .A(n1289), .B(n1290), .ZN(n1155) );
XNOR2_X1 U1019 ( .A(n1274), .B(n1291), .ZN(n1290) );
XNOR2_X1 U1020 ( .A(n1292), .B(n1293), .ZN(n1291) );
NOR2_X1 U1021 ( .A1(G953), .A2(n1083), .ZN(n1293) );
INV_X1 U1022 ( .A(G227), .ZN(n1083) );
XOR2_X1 U1023 ( .A(G104), .B(G107), .Z(n1274) );
XNOR2_X1 U1024 ( .A(n1149), .B(n1100), .ZN(n1289) );
XOR2_X1 U1025 ( .A(n1294), .B(n1295), .Z(n1100) );
NOR2_X1 U1026 ( .A1(G143), .A2(KEYINPUT54), .ZN(n1295) );
XOR2_X1 U1027 ( .A(G101), .B(n1296), .Z(n1149) );
NAND2_X1 U1028 ( .A1(KEYINPUT13), .A2(n1066), .ZN(n1287) );
INV_X1 U1029 ( .A(G469), .ZN(n1066) );
NOR2_X1 U1030 ( .A1(n1235), .A2(n1231), .ZN(n1034) );
XOR2_X1 U1031 ( .A(n1058), .B(KEYINPUT44), .Z(n1231) );
XNOR2_X1 U1032 ( .A(n1297), .B(n1298), .ZN(n1058) );
XOR2_X1 U1033 ( .A(KEYINPUT51), .B(G472), .Z(n1298) );
NAND2_X1 U1034 ( .A1(n1299), .A2(n1165), .ZN(n1297) );
XOR2_X1 U1035 ( .A(n1148), .B(n1300), .Z(n1299) );
XNOR2_X1 U1036 ( .A(n1301), .B(n1302), .ZN(n1300) );
NOR2_X1 U1037 ( .A1(KEYINPUT19), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1038 ( .A(KEYINPUT35), .B(n1296), .Z(n1303) );
XNOR2_X1 U1039 ( .A(n1304), .B(n1305), .ZN(n1296) );
NOR2_X1 U1040 ( .A1(G137), .A2(KEYINPUT38), .ZN(n1305) );
XOR2_X1 U1041 ( .A(n1219), .B(n1306), .Z(n1304) );
NOR2_X1 U1042 ( .A1(KEYINPUT43), .A2(n1104), .ZN(n1306) );
XNOR2_X1 U1043 ( .A(G131), .B(KEYINPUT28), .ZN(n1104) );
INV_X1 U1044 ( .A(G134), .ZN(n1219) );
NAND2_X1 U1045 ( .A1(KEYINPUT8), .A2(n1307), .ZN(n1301) );
XOR2_X1 U1046 ( .A(G101), .B(n1308), .Z(n1307) );
NOR2_X1 U1047 ( .A1(n1152), .A2(KEYINPUT11), .ZN(n1308) );
AND3_X1 U1048 ( .A1(n1309), .A2(n1055), .A3(G210), .ZN(n1152) );
XOR2_X1 U1049 ( .A(KEYINPUT16), .B(G237), .Z(n1309) );
XNOR2_X1 U1050 ( .A(n1310), .B(n1311), .ZN(n1148) );
XOR2_X1 U1051 ( .A(G116), .B(n1312), .Z(n1311) );
XOR2_X1 U1052 ( .A(KEYINPUT5), .B(G119), .Z(n1312) );
XOR2_X1 U1053 ( .A(n1269), .B(G113), .Z(n1310) );
XOR2_X1 U1054 ( .A(n1313), .B(n1294), .Z(n1269) );
XOR2_X1 U1055 ( .A(G128), .B(KEYINPUT36), .Z(n1294) );
XOR2_X1 U1056 ( .A(n1314), .B(G143), .Z(n1313) );
NAND2_X1 U1057 ( .A1(KEYINPUT59), .A2(n1106), .ZN(n1314) );
INV_X1 U1058 ( .A(G146), .ZN(n1106) );
INV_X1 U1059 ( .A(n1232), .ZN(n1235) );
XOR2_X1 U1060 ( .A(n1079), .B(n1315), .Z(n1232) );
NOR2_X1 U1061 ( .A1(n1316), .A2(KEYINPUT41), .ZN(n1315) );
INV_X1 U1062 ( .A(n1077), .ZN(n1316) );
NAND2_X1 U1063 ( .A1(G217), .A2(n1286), .ZN(n1077) );
NAND2_X1 U1064 ( .A1(G234), .A2(n1165), .ZN(n1286) );
NAND2_X1 U1065 ( .A1(n1128), .A2(n1165), .ZN(n1079) );
INV_X1 U1066 ( .A(G902), .ZN(n1165) );
INV_X1 U1067 ( .A(n1131), .ZN(n1128) );
XOR2_X1 U1068 ( .A(n1317), .B(n1318), .Z(n1131) );
XOR2_X1 U1069 ( .A(n1319), .B(n1320), .Z(n1318) );
XOR2_X1 U1070 ( .A(G128), .B(G125), .Z(n1320) );
XOR2_X1 U1071 ( .A(KEYINPUT61), .B(G137), .Z(n1319) );
XOR2_X1 U1072 ( .A(n1321), .B(n1292), .Z(n1317) );
XOR2_X1 U1073 ( .A(G110), .B(n1239), .Z(n1292) );
XOR2_X1 U1074 ( .A(G140), .B(G146), .Z(n1239) );
XOR2_X1 U1075 ( .A(n1322), .B(G119), .Z(n1321) );
NAND4_X1 U1076 ( .A1(KEYINPUT23), .A2(G221), .A3(G234), .A4(n1055), .ZN(n1322) );
INV_X1 U1077 ( .A(G953), .ZN(n1055) );
endmodule


