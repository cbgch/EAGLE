//Key = 0110101100111001101010100110000110110001000001000110111010001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291;

XNOR2_X1 U722 ( .A(G107), .B(n982), .ZN(G9) );
NAND4_X1 U723 ( .A1(n983), .A2(n984), .A3(n985), .A4(n986), .ZN(n982) );
XNOR2_X1 U724 ( .A(KEYINPUT36), .B(n987), .ZN(n986) );
NOR2_X1 U725 ( .A1(n988), .A2(n989), .ZN(G75) );
NOR4_X1 U726 ( .A1(n990), .A2(n991), .A3(G953), .A4(n992), .ZN(n989) );
NOR2_X1 U727 ( .A1(n993), .A2(n987), .ZN(n991) );
XOR2_X1 U728 ( .A(n994), .B(KEYINPUT47), .Z(n993) );
NAND2_X1 U729 ( .A1(n995), .A2(n996), .ZN(n990) );
NAND3_X1 U730 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n996) );
NAND2_X1 U731 ( .A1(n1000), .A2(n994), .ZN(n998) );
NAND4_X1 U732 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n985), .ZN(n994) );
NAND2_X1 U733 ( .A1(n1004), .A2(n1005), .ZN(n997) );
NAND2_X1 U734 ( .A1(n1001), .A2(n1006), .ZN(n1004) );
NAND2_X1 U735 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND3_X1 U736 ( .A1(n985), .A2(n1009), .A3(n1003), .ZN(n1008) );
NAND2_X1 U737 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND2_X1 U738 ( .A1(n1002), .A2(n1012), .ZN(n1007) );
NAND2_X1 U739 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U740 ( .A1(n985), .A2(n1015), .ZN(n1014) );
NAND2_X1 U741 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U742 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND2_X1 U743 ( .A1(n1003), .A2(n1020), .ZN(n1013) );
NAND2_X1 U744 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
INV_X1 U745 ( .A(n1023), .ZN(n1001) );
NOR3_X1 U746 ( .A1(n992), .A2(G953), .A3(G952), .ZN(n988) );
AND4_X1 U747 ( .A1(n1024), .A2(n1005), .A3(n1025), .A4(n1026), .ZN(n992) );
NOR4_X1 U748 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
XNOR2_X1 U749 ( .A(KEYINPUT44), .B(n1031), .ZN(n1030) );
XNOR2_X1 U750 ( .A(n1032), .B(KEYINPUT49), .ZN(n1027) );
NOR3_X1 U751 ( .A1(n1033), .A2(n1034), .A3(n1018), .ZN(n1025) );
XOR2_X1 U752 ( .A(n1035), .B(n1036), .Z(n1024) );
NOR2_X1 U753 ( .A1(n1037), .A2(KEYINPUT9), .ZN(n1036) );
INV_X1 U754 ( .A(n1038), .ZN(n1037) );
XOR2_X1 U755 ( .A(n1039), .B(n1040), .Z(G72) );
NOR2_X1 U756 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR2_X1 U757 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
XOR2_X1 U758 ( .A(n1045), .B(KEYINPUT26), .Z(n1044) );
NOR2_X1 U759 ( .A1(n1046), .A2(n1045), .ZN(n1041) );
NAND2_X1 U760 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
INV_X1 U761 ( .A(n1043), .ZN(n1046) );
NAND2_X1 U762 ( .A1(n1049), .A2(n1050), .ZN(n1043) );
NAND2_X1 U763 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XNOR2_X1 U764 ( .A(KEYINPUT5), .B(n1047), .ZN(n1051) );
XOR2_X1 U765 ( .A(n1053), .B(n1054), .Z(n1049) );
XNOR2_X1 U766 ( .A(n1055), .B(n1056), .ZN(n1054) );
XNOR2_X1 U767 ( .A(G125), .B(n1057), .ZN(n1053) );
XNOR2_X1 U768 ( .A(KEYINPUT33), .B(n1058), .ZN(n1057) );
INV_X1 U769 ( .A(G134), .ZN(n1058) );
NAND2_X1 U770 ( .A1(G953), .A2(n1059), .ZN(n1039) );
NAND2_X1 U771 ( .A1(G900), .A2(G227), .ZN(n1059) );
XOR2_X1 U772 ( .A(n1060), .B(n1061), .Z(G69) );
NOR3_X1 U773 ( .A1(n1047), .A2(KEYINPUT38), .A3(n1062), .ZN(n1061) );
AND2_X1 U774 ( .A1(G224), .A2(G898), .ZN(n1062) );
NAND2_X1 U775 ( .A1(n1063), .A2(n1064), .ZN(n1060) );
NAND2_X1 U776 ( .A1(n1065), .A2(n1047), .ZN(n1064) );
XOR2_X1 U777 ( .A(n1066), .B(n1067), .Z(n1065) );
NAND3_X1 U778 ( .A1(G898), .A2(n1067), .A3(G953), .ZN(n1063) );
NOR2_X1 U779 ( .A1(n1068), .A2(n1069), .ZN(G66) );
XNOR2_X1 U780 ( .A(n1070), .B(n1071), .ZN(n1069) );
NOR3_X1 U781 ( .A1(n1072), .A2(n995), .A3(n1038), .ZN(n1071) );
XNOR2_X1 U782 ( .A(KEYINPUT32), .B(n1073), .ZN(n1072) );
NOR2_X1 U783 ( .A1(n1068), .A2(n1074), .ZN(G63) );
XOR2_X1 U784 ( .A(n1075), .B(n1076), .Z(n1074) );
NOR2_X1 U785 ( .A1(n1077), .A2(KEYINPUT0), .ZN(n1075) );
AND2_X1 U786 ( .A1(G478), .A2(n1078), .ZN(n1077) );
NOR2_X1 U787 ( .A1(n1068), .A2(n1079), .ZN(G60) );
XOR2_X1 U788 ( .A(n1080), .B(n1081), .Z(n1079) );
NAND2_X1 U789 ( .A1(n1078), .A2(G475), .ZN(n1080) );
XNOR2_X1 U790 ( .A(G104), .B(n1082), .ZN(G6) );
NOR2_X1 U791 ( .A1(n1068), .A2(n1083), .ZN(G57) );
XOR2_X1 U792 ( .A(n1084), .B(n1085), .Z(n1083) );
XNOR2_X1 U793 ( .A(n1086), .B(n1087), .ZN(n1085) );
NAND2_X1 U794 ( .A1(n1078), .A2(G472), .ZN(n1086) );
XOR2_X1 U795 ( .A(n1088), .B(n1089), .Z(n1084) );
NAND2_X1 U796 ( .A1(KEYINPUT11), .A2(n1090), .ZN(n1089) );
XNOR2_X1 U797 ( .A(n1091), .B(n1092), .ZN(n1090) );
XNOR2_X1 U798 ( .A(n1093), .B(KEYINPUT13), .ZN(n1092) );
NAND2_X1 U799 ( .A1(KEYINPUT45), .A2(n1094), .ZN(n1093) );
XOR2_X1 U800 ( .A(KEYINPUT25), .B(n1095), .Z(n1094) );
NAND2_X1 U801 ( .A1(n1096), .A2(n1097), .ZN(n1088) );
NAND2_X1 U802 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U803 ( .A(n1100), .B(KEYINPUT41), .Z(n1096) );
OR2_X1 U804 ( .A1(n1098), .A2(n1099), .ZN(n1100) );
NOR2_X1 U805 ( .A1(n1068), .A2(n1101), .ZN(G54) );
XOR2_X1 U806 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U807 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U808 ( .A(n1106), .B(n1107), .Z(n1102) );
NAND2_X1 U809 ( .A1(n1078), .A2(G469), .ZN(n1106) );
NOR2_X1 U810 ( .A1(n1068), .A2(n1108), .ZN(G51) );
XOR2_X1 U811 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U812 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U813 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
INV_X1 U814 ( .A(n1115), .ZN(n1114) );
XNOR2_X1 U815 ( .A(KEYINPUT24), .B(n1116), .ZN(n1113) );
NOR2_X1 U816 ( .A1(n1115), .A2(n1116), .ZN(n1111) );
XOR2_X1 U817 ( .A(n1117), .B(n1067), .Z(n1109) );
NAND2_X1 U818 ( .A1(n1078), .A2(n1118), .ZN(n1117) );
NOR2_X1 U819 ( .A1(n1073), .A2(n995), .ZN(n1078) );
NOR2_X1 U820 ( .A1(n1048), .A2(n1066), .ZN(n995) );
NAND4_X1 U821 ( .A1(n1082), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1066) );
NOR4_X1 U822 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1121) );
NAND2_X1 U823 ( .A1(n1126), .A2(n1127), .ZN(n1120) );
NAND2_X1 U824 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND3_X1 U825 ( .A1(n984), .A2(n985), .A3(n983), .ZN(n1129) );
XOR2_X1 U826 ( .A(n1130), .B(KEYINPUT57), .Z(n1128) );
NAND4_X1 U827 ( .A1(n1131), .A2(n983), .A3(n1126), .A4(n985), .ZN(n1082) );
NAND4_X1 U828 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1048) );
NOR4_X1 U829 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1135) );
NOR2_X1 U830 ( .A1(n1140), .A2(n1141), .ZN(n1134) );
NOR3_X1 U831 ( .A1(n1142), .A2(n1022), .A3(n1010), .ZN(n1141) );
NOR4_X1 U832 ( .A1(n1143), .A2(n1144), .A3(n1011), .A4(n1145), .ZN(n1140) );
INV_X1 U833 ( .A(n1146), .ZN(n1144) );
XNOR2_X1 U834 ( .A(n1147), .B(KEYINPUT46), .ZN(n1143) );
NOR2_X1 U835 ( .A1(n1047), .A2(G952), .ZN(n1068) );
NAND2_X1 U836 ( .A1(n1148), .A2(n1149), .ZN(G48) );
NAND2_X1 U837 ( .A1(n1150), .A2(n1133), .ZN(n1149) );
NAND2_X1 U838 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
OR2_X1 U839 ( .A1(KEYINPUT58), .A2(KEYINPUT60), .ZN(n1152) );
NAND3_X1 U840 ( .A1(n1153), .A2(n1154), .A3(KEYINPUT60), .ZN(n1148) );
OR2_X1 U841 ( .A1(n1151), .A2(KEYINPUT58), .ZN(n1154) );
NAND2_X1 U842 ( .A1(n1155), .A2(n1151), .ZN(n1153) );
OR2_X1 U843 ( .A1(n1133), .A2(KEYINPUT58), .ZN(n1155) );
NAND4_X1 U844 ( .A1(n1156), .A2(n1131), .A3(n1157), .A4(n1147), .ZN(n1133) );
XNOR2_X1 U845 ( .A(G143), .B(n1132), .ZN(G45) );
NAND3_X1 U846 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1132) );
NOR3_X1 U847 ( .A1(n1022), .A2(n1031), .A3(n1159), .ZN(n1158) );
XOR2_X1 U848 ( .A(G140), .B(n1139), .Z(G42) );
NOR3_X1 U849 ( .A1(n1010), .A2(n1021), .A3(n1142), .ZN(n1139) );
INV_X1 U850 ( .A(n1160), .ZN(n1021) );
XOR2_X1 U851 ( .A(G137), .B(n1138), .Z(G39) );
NOR3_X1 U852 ( .A1(n1142), .A2(n1161), .A3(n1162), .ZN(n1138) );
INV_X1 U853 ( .A(n1147), .ZN(n1161) );
XOR2_X1 U854 ( .A(n1163), .B(n1137), .Z(G36) );
NOR3_X1 U855 ( .A1(n1011), .A2(n1022), .A3(n1142), .ZN(n1137) );
XNOR2_X1 U856 ( .A(G134), .B(KEYINPUT39), .ZN(n1163) );
XOR2_X1 U857 ( .A(G131), .B(n1164), .Z(G33) );
NOR4_X1 U858 ( .A1(KEYINPUT43), .A2(n1022), .A3(n1010), .A4(n1142), .ZN(n1164) );
NAND4_X1 U859 ( .A1(n1156), .A2(n999), .A3(n1165), .A4(n1005), .ZN(n1142) );
INV_X1 U860 ( .A(n1016), .ZN(n1156) );
XOR2_X1 U861 ( .A(n1146), .B(KEYINPUT4), .Z(n1016) );
INV_X1 U862 ( .A(n1131), .ZN(n1010) );
INV_X1 U863 ( .A(n1166), .ZN(n1022) );
XNOR2_X1 U864 ( .A(G128), .B(n1167), .ZN(G30) );
NAND4_X1 U865 ( .A1(n1157), .A2(n1147), .A3(n984), .A4(n1146), .ZN(n1167) );
XNOR2_X1 U866 ( .A(G101), .B(n1119), .ZN(G3) );
NAND4_X1 U867 ( .A1(n1002), .A2(n983), .A3(n1166), .A4(n1126), .ZN(n1119) );
XOR2_X1 U868 ( .A(G125), .B(n1136), .Z(G27) );
AND4_X1 U869 ( .A1(n1131), .A2(n1003), .A3(n1157), .A4(n1160), .ZN(n1136) );
INV_X1 U870 ( .A(n1145), .ZN(n1157) );
NAND2_X1 U871 ( .A1(n1126), .A2(n1165), .ZN(n1145) );
NAND2_X1 U872 ( .A1(n1023), .A2(n1168), .ZN(n1165) );
NAND4_X1 U873 ( .A1(G953), .A2(G902), .A3(n1169), .A4(n1052), .ZN(n1168) );
INV_X1 U874 ( .A(G900), .ZN(n1052) );
XOR2_X1 U875 ( .A(G122), .B(n1125), .Z(G24) );
AND4_X1 U876 ( .A1(n1170), .A2(n985), .A3(n1028), .A4(n1171), .ZN(n1125) );
NAND2_X1 U877 ( .A1(n1172), .A2(n1173), .ZN(n985) );
NAND2_X1 U878 ( .A1(n1166), .A2(n1174), .ZN(n1173) );
NAND3_X1 U879 ( .A1(n1175), .A2(n1176), .A3(KEYINPUT53), .ZN(n1172) );
XNOR2_X1 U880 ( .A(n1177), .B(n1124), .ZN(G21) );
AND3_X1 U881 ( .A1(n1002), .A2(n1147), .A3(n1170), .ZN(n1124) );
XOR2_X1 U882 ( .A(G116), .B(n1123), .Z(G18) );
AND3_X1 U883 ( .A1(n984), .A2(n1166), .A3(n1170), .ZN(n1123) );
INV_X1 U884 ( .A(n1011), .ZN(n984) );
NAND2_X1 U885 ( .A1(n1031), .A2(n1178), .ZN(n1011) );
XNOR2_X1 U886 ( .A(KEYINPUT28), .B(n1159), .ZN(n1178) );
XNOR2_X1 U887 ( .A(n1122), .B(n1179), .ZN(G15) );
NAND2_X1 U888 ( .A1(KEYINPUT12), .A2(G113), .ZN(n1179) );
AND3_X1 U889 ( .A1(n1131), .A2(n1166), .A3(n1170), .ZN(n1122) );
AND3_X1 U890 ( .A1(n1126), .A2(n1180), .A3(n1003), .ZN(n1170) );
AND2_X1 U891 ( .A1(n1019), .A2(n1181), .ZN(n1003) );
NOR2_X1 U892 ( .A1(n1182), .A2(n1176), .ZN(n1166) );
NOR2_X1 U893 ( .A1(n1028), .A2(n1031), .ZN(n1131) );
XNOR2_X1 U894 ( .A(G110), .B(n1183), .ZN(G12) );
NOR2_X1 U895 ( .A1(n1184), .A2(KEYINPUT61), .ZN(n1183) );
NOR2_X1 U896 ( .A1(n987), .A2(n1130), .ZN(n1184) );
NAND3_X1 U897 ( .A1(n983), .A2(n1160), .A3(n1002), .ZN(n1130) );
INV_X1 U898 ( .A(n1162), .ZN(n1002) );
NAND2_X1 U899 ( .A1(n1031), .A2(n1159), .ZN(n1162) );
INV_X1 U900 ( .A(n1028), .ZN(n1159) );
XOR2_X1 U901 ( .A(G478), .B(n1185), .Z(n1028) );
AND2_X1 U902 ( .A1(n1073), .A2(n1076), .ZN(n1185) );
XNOR2_X1 U903 ( .A(n1186), .B(n1187), .ZN(n1076) );
XOR2_X1 U904 ( .A(n1188), .B(n1189), .Z(n1187) );
NAND2_X1 U905 ( .A1(G217), .A2(n1190), .ZN(n1189) );
NAND3_X1 U906 ( .A1(n1191), .A2(n1192), .A3(KEYINPUT63), .ZN(n1188) );
NAND2_X1 U907 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
INV_X1 U908 ( .A(KEYINPUT62), .ZN(n1194) );
XNOR2_X1 U909 ( .A(n1195), .B(n1196), .ZN(n1193) );
NAND2_X1 U910 ( .A1(KEYINPUT2), .A2(G128), .ZN(n1195) );
NAND3_X1 U911 ( .A1(G143), .A2(n1197), .A3(KEYINPUT62), .ZN(n1191) );
XOR2_X1 U912 ( .A(n1198), .B(n1199), .Z(n1186) );
NOR2_X1 U913 ( .A1(KEYINPUT21), .A2(n1200), .ZN(n1199) );
XNOR2_X1 U914 ( .A(n1201), .B(n1202), .ZN(n1200) );
XOR2_X1 U915 ( .A(G122), .B(G116), .Z(n1202) );
XNOR2_X1 U916 ( .A(G134), .B(KEYINPUT10), .ZN(n1198) );
INV_X1 U917 ( .A(n1171), .ZN(n1031) );
XNOR2_X1 U918 ( .A(n1203), .B(G475), .ZN(n1171) );
NAND2_X1 U919 ( .A1(n1081), .A2(n1073), .ZN(n1203) );
XNOR2_X1 U920 ( .A(n1204), .B(n1205), .ZN(n1081) );
XOR2_X1 U921 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U922 ( .A(n1208), .B(n1209), .Z(n1204) );
XNOR2_X1 U923 ( .A(n1210), .B(n1211), .ZN(n1208) );
NAND2_X1 U924 ( .A1(n1212), .A2(n1213), .ZN(n1210) );
NAND4_X1 U925 ( .A1(G214), .A2(G143), .A3(n1214), .A4(n1047), .ZN(n1213) );
XOR2_X1 U926 ( .A(n1215), .B(KEYINPUT30), .Z(n1212) );
NAND2_X1 U927 ( .A1(n1196), .A2(n1216), .ZN(n1215) );
NAND3_X1 U928 ( .A1(n1214), .A2(n1047), .A3(G214), .ZN(n1216) );
XNOR2_X1 U929 ( .A(n1217), .B(KEYINPUT1), .ZN(n1214) );
NAND2_X1 U930 ( .A1(n1218), .A2(n1219), .ZN(n1160) );
NAND2_X1 U931 ( .A1(n1147), .A2(n1174), .ZN(n1219) );
INV_X1 U932 ( .A(KEYINPUT53), .ZN(n1174) );
NOR2_X1 U933 ( .A1(n1175), .A2(n1176), .ZN(n1147) );
NAND3_X1 U934 ( .A1(n1176), .A2(n1182), .A3(KEYINPUT53), .ZN(n1218) );
INV_X1 U935 ( .A(n1175), .ZN(n1182) );
XOR2_X1 U936 ( .A(n1220), .B(n1038), .Z(n1175) );
NAND2_X1 U937 ( .A1(G217), .A2(n1221), .ZN(n1038) );
XNOR2_X1 U938 ( .A(n1035), .B(KEYINPUT16), .ZN(n1220) );
AND2_X1 U939 ( .A1(n1073), .A2(n1070), .ZN(n1035) );
NAND3_X1 U940 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1070) );
NAND2_X1 U941 ( .A1(KEYINPUT55), .A2(n1225), .ZN(n1224) );
OR3_X1 U942 ( .A1(n1225), .A2(KEYINPUT55), .A3(n1226), .ZN(n1223) );
NAND2_X1 U943 ( .A1(n1226), .A2(n1227), .ZN(n1222) );
NAND2_X1 U944 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
INV_X1 U945 ( .A(KEYINPUT55), .ZN(n1229) );
XOR2_X1 U946 ( .A(KEYINPUT20), .B(n1225), .Z(n1228) );
XNOR2_X1 U947 ( .A(n1230), .B(n1231), .ZN(n1225) );
XOR2_X1 U948 ( .A(n1206), .B(n1232), .Z(n1231) );
XOR2_X1 U949 ( .A(n1233), .B(n1234), .Z(n1232) );
NOR2_X1 U950 ( .A1(G140), .A2(KEYINPUT40), .ZN(n1233) );
XOR2_X1 U951 ( .A(n1235), .B(KEYINPUT3), .Z(n1206) );
XNOR2_X1 U952 ( .A(G119), .B(n1236), .ZN(n1230) );
XNOR2_X1 U953 ( .A(KEYINPUT19), .B(n1197), .ZN(n1236) );
INV_X1 U954 ( .A(G128), .ZN(n1197) );
XOR2_X1 U955 ( .A(n1237), .B(n1238), .Z(n1226) );
XOR2_X1 U956 ( .A(KEYINPUT29), .B(G137), .Z(n1238) );
NAND2_X1 U957 ( .A1(n1190), .A2(G221), .ZN(n1237) );
AND2_X1 U958 ( .A1(G234), .A2(n1047), .ZN(n1190) );
INV_X1 U959 ( .A(n1032), .ZN(n1176) );
XNOR2_X1 U960 ( .A(n1239), .B(G472), .ZN(n1032) );
NAND2_X1 U961 ( .A1(n1240), .A2(n1073), .ZN(n1239) );
XNOR2_X1 U962 ( .A(n1241), .B(n1242), .ZN(n1240) );
INV_X1 U963 ( .A(n1087), .ZN(n1242) );
XOR2_X1 U964 ( .A(n1243), .B(n1211), .Z(n1087) );
NAND2_X1 U965 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XNOR2_X1 U966 ( .A(n1246), .B(n1247), .ZN(n1241) );
NAND2_X1 U967 ( .A1(KEYINPUT34), .A2(n1248), .ZN(n1247) );
XOR2_X1 U968 ( .A(n1098), .B(n1249), .Z(n1248) );
XNOR2_X1 U969 ( .A(G101), .B(KEYINPUT51), .ZN(n1249) );
NAND3_X1 U970 ( .A1(n1217), .A2(n1047), .A3(G210), .ZN(n1098) );
NAND2_X1 U971 ( .A1(n1250), .A2(KEYINPUT50), .ZN(n1246) );
XNOR2_X1 U972 ( .A(n1095), .B(n1251), .ZN(n1250) );
NOR2_X1 U973 ( .A1(KEYINPUT42), .A2(n1091), .ZN(n1251) );
XOR2_X1 U974 ( .A(n1252), .B(G146), .Z(n1091) );
XNOR2_X1 U975 ( .A(n1253), .B(G131), .ZN(n1095) );
AND2_X1 U976 ( .A1(n1146), .A2(n1180), .ZN(n983) );
NAND2_X1 U977 ( .A1(n1023), .A2(n1254), .ZN(n1180) );
NAND4_X1 U978 ( .A1(G953), .A2(G902), .A3(n1169), .A4(n1255), .ZN(n1254) );
INV_X1 U979 ( .A(G898), .ZN(n1255) );
NAND3_X1 U980 ( .A1(n1169), .A2(n1047), .A3(G952), .ZN(n1023) );
NAND2_X1 U981 ( .A1(G237), .A2(G234), .ZN(n1169) );
NOR2_X1 U982 ( .A1(n1018), .A2(n1019), .ZN(n1146) );
NOR2_X1 U983 ( .A1(n1256), .A2(n1033), .ZN(n1019) );
NOR2_X1 U984 ( .A1(n1257), .A2(n1258), .ZN(n1033) );
AND2_X1 U985 ( .A1(n1259), .A2(n1073), .ZN(n1258) );
XOR2_X1 U986 ( .A(n1034), .B(KEYINPUT23), .Z(n1256) );
AND3_X1 U987 ( .A1(n1257), .A2(n1073), .A3(n1259), .ZN(n1034) );
XOR2_X1 U988 ( .A(n1260), .B(n1261), .Z(n1259) );
XNOR2_X1 U989 ( .A(n1262), .B(KEYINPUT37), .ZN(n1261) );
NAND2_X1 U990 ( .A1(n1263), .A2(KEYINPUT35), .ZN(n1262) );
XOR2_X1 U991 ( .A(n1264), .B(n1107), .Z(n1263) );
NOR2_X1 U992 ( .A1(KEYINPUT17), .A2(n1265), .ZN(n1107) );
XNOR2_X1 U993 ( .A(n1201), .B(n1266), .ZN(n1265) );
XNOR2_X1 U994 ( .A(G101), .B(KEYINPUT15), .ZN(n1264) );
XOR2_X1 U995 ( .A(n1104), .B(n1234), .Z(n1260) );
XNOR2_X1 U996 ( .A(n1267), .B(n1268), .ZN(n1104) );
INV_X1 U997 ( .A(n1055), .ZN(n1268) );
XOR2_X1 U998 ( .A(n1207), .B(n1269), .Z(n1055) );
XNOR2_X1 U999 ( .A(G128), .B(n1270), .ZN(n1269) );
NAND2_X1 U1000 ( .A1(n1271), .A2(KEYINPUT6), .ZN(n1270) );
XNOR2_X1 U1001 ( .A(n1272), .B(n1196), .ZN(n1271) );
NAND2_X1 U1002 ( .A1(KEYINPUT22), .A2(n1151), .ZN(n1272) );
XOR2_X1 U1003 ( .A(G131), .B(G140), .Z(n1207) );
XOR2_X1 U1004 ( .A(n1253), .B(n1273), .Z(n1267) );
AND2_X1 U1005 ( .A1(n1047), .A2(G227), .ZN(n1273) );
XOR2_X1 U1006 ( .A(n1274), .B(n1056), .Z(n1253) );
XOR2_X1 U1007 ( .A(G137), .B(KEYINPUT56), .Z(n1056) );
NAND2_X1 U1008 ( .A1(KEYINPUT31), .A2(G134), .ZN(n1274) );
XOR2_X1 U1009 ( .A(G469), .B(KEYINPUT52), .Z(n1257) );
INV_X1 U1010 ( .A(n1181), .ZN(n1018) );
NAND2_X1 U1011 ( .A1(G221), .A2(n1221), .ZN(n1181) );
NAND2_X1 U1012 ( .A1(G234), .A2(n1073), .ZN(n1221) );
INV_X1 U1013 ( .A(n1126), .ZN(n987) );
NOR2_X1 U1014 ( .A1(n999), .A2(n1000), .ZN(n1126) );
INV_X1 U1015 ( .A(n1005), .ZN(n1000) );
NAND2_X1 U1016 ( .A1(G214), .A2(n1275), .ZN(n1005) );
INV_X1 U1017 ( .A(n1029), .ZN(n999) );
XNOR2_X1 U1018 ( .A(n1276), .B(n1118), .ZN(n1029) );
AND2_X1 U1019 ( .A1(G210), .A2(n1275), .ZN(n1118) );
NAND2_X1 U1020 ( .A1(n1217), .A2(n1073), .ZN(n1275) );
INV_X1 U1021 ( .A(G237), .ZN(n1217) );
NAND2_X1 U1022 ( .A1(n1277), .A2(n1073), .ZN(n1276) );
INV_X1 U1023 ( .A(G902), .ZN(n1073) );
XOR2_X1 U1024 ( .A(n1278), .B(n1279), .Z(n1277) );
XNOR2_X1 U1025 ( .A(KEYINPUT48), .B(n1116), .ZN(n1279) );
NAND2_X1 U1026 ( .A1(G224), .A2(n1047), .ZN(n1116) );
INV_X1 U1027 ( .A(G953), .ZN(n1047) );
XNOR2_X1 U1028 ( .A(n1067), .B(n1115), .ZN(n1278) );
XNOR2_X1 U1029 ( .A(n1252), .B(n1235), .ZN(n1115) );
XNOR2_X1 U1030 ( .A(G125), .B(n1151), .ZN(n1235) );
INV_X1 U1031 ( .A(G146), .ZN(n1151) );
XNOR2_X1 U1032 ( .A(G128), .B(n1280), .ZN(n1252) );
XNOR2_X1 U1033 ( .A(KEYINPUT59), .B(n1196), .ZN(n1280) );
INV_X1 U1034 ( .A(G143), .ZN(n1196) );
XNOR2_X1 U1035 ( .A(n1281), .B(n1282), .ZN(n1067) );
XOR2_X1 U1036 ( .A(n1209), .B(n1105), .Z(n1282) );
XNOR2_X1 U1037 ( .A(n1099), .B(n1234), .ZN(n1105) );
XOR2_X1 U1038 ( .A(G110), .B(KEYINPUT54), .Z(n1234) );
INV_X1 U1039 ( .A(G101), .ZN(n1099) );
XOR2_X1 U1040 ( .A(G122), .B(n1266), .Z(n1209) );
XOR2_X1 U1041 ( .A(G104), .B(KEYINPUT8), .Z(n1266) );
XOR2_X1 U1042 ( .A(n1283), .B(n1284), .Z(n1281) );
NOR2_X1 U1043 ( .A1(KEYINPUT27), .A2(n1201), .ZN(n1284) );
INV_X1 U1044 ( .A(G107), .ZN(n1201) );
NAND2_X1 U1045 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
NAND3_X1 U1046 ( .A1(n1245), .A2(n1211), .A3(n1287), .ZN(n1286) );
INV_X1 U1047 ( .A(G113), .ZN(n1211) );
NAND2_X1 U1048 ( .A1(n1288), .A2(n1289), .ZN(n1285) );
NAND2_X1 U1049 ( .A1(n1287), .A2(n1245), .ZN(n1289) );
NAND2_X1 U1050 ( .A1(n1290), .A2(n1177), .ZN(n1245) );
INV_X1 U1051 ( .A(G119), .ZN(n1177) );
XNOR2_X1 U1052 ( .A(KEYINPUT18), .B(G116), .ZN(n1290) );
XOR2_X1 U1053 ( .A(n1244), .B(KEYINPUT14), .Z(n1287) );
NAND2_X1 U1054 ( .A1(G119), .A2(n1291), .ZN(n1244) );
XOR2_X1 U1055 ( .A(KEYINPUT18), .B(G116), .Z(n1291) );
XNOR2_X1 U1056 ( .A(G113), .B(KEYINPUT7), .ZN(n1288) );
endmodule


