//Key = 0001000101111010001100011001001001011110100101110011000011001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285;

XNOR2_X1 U708 ( .A(G107), .B(n982), .ZN(G9) );
NOR2_X1 U709 ( .A1(n983), .A2(n984), .ZN(G75) );
NOR3_X1 U710 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n984) );
NOR2_X1 U711 ( .A1(n988), .A2(n989), .ZN(n986) );
NOR3_X1 U712 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n988) );
NOR3_X1 U713 ( .A1(n993), .A2(n994), .A3(n995), .ZN(n992) );
NOR2_X1 U714 ( .A1(n996), .A2(n997), .ZN(n994) );
AND2_X1 U715 ( .A1(n998), .A2(n999), .ZN(n997) );
NOR2_X1 U716 ( .A1(n1000), .A2(n1001), .ZN(n996) );
INV_X1 U717 ( .A(n1002), .ZN(n1001) );
NOR2_X1 U718 ( .A1(n1003), .A2(n1004), .ZN(n1000) );
XNOR2_X1 U719 ( .A(n1005), .B(KEYINPUT14), .ZN(n1004) );
NOR3_X1 U720 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n991) );
NOR2_X1 U721 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
XOR2_X1 U722 ( .A(KEYINPUT26), .B(n1011), .Z(n990) );
NOR3_X1 U723 ( .A1(n1012), .A2(n995), .A3(n1006), .ZN(n1011) );
INV_X1 U724 ( .A(n1013), .ZN(n1006) );
INV_X1 U725 ( .A(n1014), .ZN(n995) );
NAND3_X1 U726 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n985) );
NAND4_X1 U727 ( .A1(n1013), .A2(n1014), .A3(n1018), .A4(n1012), .ZN(n1017) );
NAND2_X1 U728 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND2_X1 U729 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
XOR2_X1 U730 ( .A(KEYINPUT47), .B(n1023), .Z(n1019) );
NOR3_X1 U731 ( .A1(n1024), .A2(n1025), .A3(n993), .ZN(n1013) );
INV_X1 U732 ( .A(n999), .ZN(n1025) );
NOR3_X1 U733 ( .A1(n1026), .A2(G953), .A3(G952), .ZN(n983) );
INV_X1 U734 ( .A(n1015), .ZN(n1026) );
NAND4_X1 U735 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1015) );
NOR4_X1 U736 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
XNOR2_X1 U737 ( .A(KEYINPUT29), .B(n1035), .ZN(n1034) );
NOR3_X1 U738 ( .A1(n1007), .A2(n1021), .A3(n1036), .ZN(n1029) );
NAND2_X1 U739 ( .A1(n1037), .A2(n1038), .ZN(n1028) );
XOR2_X1 U740 ( .A(n1039), .B(n1040), .Z(n1027) );
NOR2_X1 U741 ( .A1(G478), .A2(KEYINPUT32), .ZN(n1040) );
XOR2_X1 U742 ( .A(n1041), .B(n1042), .Z(G72) );
XOR2_X1 U743 ( .A(n1043), .B(n1044), .Z(n1042) );
NOR2_X1 U744 ( .A1(n1016), .A2(n1045), .ZN(n1044) );
XOR2_X1 U745 ( .A(KEYINPUT52), .B(n1046), .Z(n1045) );
NOR2_X1 U746 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U747 ( .A1(n1049), .A2(n1050), .ZN(n1043) );
NAND2_X1 U748 ( .A1(G953), .A2(n1051), .ZN(n1050) );
XNOR2_X1 U749 ( .A(KEYINPUT7), .B(n1048), .ZN(n1051) );
XOR2_X1 U750 ( .A(n1052), .B(n1053), .Z(n1049) );
XOR2_X1 U751 ( .A(n1054), .B(n1055), .Z(n1053) );
XOR2_X1 U752 ( .A(n1056), .B(G125), .Z(n1055) );
NAND2_X1 U753 ( .A1(KEYINPUT3), .A2(n1057), .ZN(n1056) );
NAND2_X1 U754 ( .A1(KEYINPUT56), .A2(n1058), .ZN(n1054) );
NAND2_X1 U755 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U756 ( .A1(G134), .A2(n1061), .ZN(n1060) );
XOR2_X1 U757 ( .A(n1062), .B(KEYINPUT31), .Z(n1059) );
OR2_X1 U758 ( .A1(n1061), .A2(G134), .ZN(n1062) );
XOR2_X1 U759 ( .A(G137), .B(KEYINPUT35), .Z(n1061) );
XNOR2_X1 U760 ( .A(n1063), .B(n1064), .ZN(n1052) );
NOR2_X1 U761 ( .A1(KEYINPUT63), .A2(n1065), .ZN(n1064) );
NAND2_X1 U762 ( .A1(n1016), .A2(n1066), .ZN(n1041) );
NAND2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XOR2_X1 U764 ( .A(n1069), .B(KEYINPUT1), .Z(n1067) );
XOR2_X1 U765 ( .A(n1070), .B(n1071), .Z(G69) );
NOR2_X1 U766 ( .A1(n1072), .A2(n1016), .ZN(n1071) );
NOR2_X1 U767 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U768 ( .A1(KEYINPUT4), .A2(n1075), .ZN(n1070) );
NOR2_X1 U769 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U770 ( .A(KEYINPUT42), .B(n1078), .Z(n1077) );
AND2_X1 U771 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U772 ( .A1(n1080), .A2(n1079), .ZN(n1076) );
NAND2_X1 U773 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NAND2_X1 U774 ( .A1(G953), .A2(n1074), .ZN(n1082) );
XNOR2_X1 U775 ( .A(n1083), .B(n1084), .ZN(n1081) );
XOR2_X1 U776 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U777 ( .A1(G953), .A2(n1087), .ZN(n1080) );
NOR2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(G66) );
XOR2_X1 U779 ( .A(n1090), .B(n1091), .Z(n1089) );
XOR2_X1 U780 ( .A(KEYINPUT27), .B(n1092), .Z(n1091) );
NOR2_X1 U781 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(G63) );
XOR2_X1 U783 ( .A(n1097), .B(n1098), .Z(n1096) );
XOR2_X1 U784 ( .A(KEYINPUT53), .B(n1099), .Z(n1098) );
NOR2_X1 U785 ( .A1(n1094), .A2(n1100), .ZN(n1099) );
INV_X1 U786 ( .A(G478), .ZN(n1100) );
NOR2_X1 U787 ( .A1(G952), .A2(n1101), .ZN(n1095) );
XNOR2_X1 U788 ( .A(G953), .B(KEYINPUT2), .ZN(n1101) );
NOR2_X1 U789 ( .A1(n1088), .A2(n1102), .ZN(G60) );
XOR2_X1 U790 ( .A(n1103), .B(n1104), .Z(n1102) );
XOR2_X1 U791 ( .A(KEYINPUT0), .B(n1105), .Z(n1104) );
NOR2_X1 U792 ( .A1(n1106), .A2(n1094), .ZN(n1105) );
XOR2_X1 U793 ( .A(n1107), .B(n1108), .Z(G6) );
XNOR2_X1 U794 ( .A(G104), .B(KEYINPUT58), .ZN(n1108) );
NOR2_X1 U795 ( .A1(n1088), .A2(n1109), .ZN(G57) );
XOR2_X1 U796 ( .A(n1110), .B(n1111), .Z(n1109) );
XNOR2_X1 U797 ( .A(n1112), .B(n1113), .ZN(n1111) );
XOR2_X1 U798 ( .A(n1086), .B(n1114), .Z(n1110) );
NOR2_X1 U799 ( .A1(n1115), .A2(n1094), .ZN(n1114) );
NOR2_X1 U800 ( .A1(n1116), .A2(n1117), .ZN(G54) );
XOR2_X1 U801 ( .A(KEYINPUT16), .B(n1088), .Z(n1117) );
XOR2_X1 U802 ( .A(n1118), .B(n1119), .Z(n1116) );
XNOR2_X1 U803 ( .A(n1120), .B(n1121), .ZN(n1119) );
XOR2_X1 U804 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U805 ( .A1(n1124), .A2(n1094), .ZN(n1123) );
NAND2_X1 U806 ( .A1(KEYINPUT51), .A2(n1057), .ZN(n1122) );
XOR2_X1 U807 ( .A(n1125), .B(n1126), .Z(n1118) );
NOR3_X1 U808 ( .A1(n1088), .A2(n1127), .A3(n1128), .ZN(G51) );
NOR2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XOR2_X1 U810 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U811 ( .A1(KEYINPUT55), .A2(n1133), .ZN(n1132) );
INV_X1 U812 ( .A(KEYINPUT25), .ZN(n1129) );
NOR2_X1 U813 ( .A1(KEYINPUT25), .A2(n1134), .ZN(n1127) );
XOR2_X1 U814 ( .A(n1131), .B(n1135), .Z(n1134) );
NOR2_X1 U815 ( .A1(KEYINPUT55), .A2(n1136), .ZN(n1135) );
XOR2_X1 U816 ( .A(n1137), .B(n1138), .Z(n1131) );
NOR2_X1 U817 ( .A1(n1139), .A2(n1094), .ZN(n1138) );
NAND2_X1 U818 ( .A1(G902), .A2(n987), .ZN(n1094) );
NAND3_X1 U819 ( .A1(n1068), .A2(n1069), .A3(n1087), .ZN(n987) );
AND2_X1 U820 ( .A1(n1140), .A2(n1141), .ZN(n1087) );
AND4_X1 U821 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1141) );
AND4_X1 U822 ( .A1(n1107), .A2(n982), .A3(n1146), .A4(n1147), .ZN(n1140) );
NAND3_X1 U823 ( .A1(n1014), .A2(n1148), .A3(n1005), .ZN(n982) );
NAND3_X1 U824 ( .A1(n1014), .A2(n1148), .A3(n1003), .ZN(n1107) );
AND4_X1 U825 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1068) );
NOR4_X1 U826 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1152) );
NAND3_X1 U827 ( .A1(n1157), .A2(n1005), .A3(n1158), .ZN(n1151) );
NOR2_X1 U828 ( .A1(n1016), .A2(G952), .ZN(n1088) );
XNOR2_X1 U829 ( .A(G146), .B(n1149), .ZN(G48) );
NAND3_X1 U830 ( .A1(n1003), .A2(n1023), .A3(n1159), .ZN(n1149) );
XNOR2_X1 U831 ( .A(G143), .B(n1150), .ZN(G45) );
NAND4_X1 U832 ( .A1(n1158), .A2(n1023), .A3(n1160), .A4(n1032), .ZN(n1150) );
XOR2_X1 U833 ( .A(n1161), .B(n1156), .Z(G42) );
AND3_X1 U834 ( .A1(n1157), .A2(n998), .A3(n1162), .ZN(n1156) );
NAND2_X1 U835 ( .A1(KEYINPUT33), .A2(n1163), .ZN(n1161) );
XOR2_X1 U836 ( .A(G137), .B(n1164), .Z(G39) );
NOR2_X1 U837 ( .A1(KEYINPUT48), .A2(n1069), .ZN(n1164) );
NAND3_X1 U838 ( .A1(n1157), .A2(n999), .A3(n1159), .ZN(n1069) );
XOR2_X1 U839 ( .A(G134), .B(n1165), .Z(G36) );
NOR3_X1 U840 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1165) );
INV_X1 U841 ( .A(n1005), .ZN(n1168) );
XNOR2_X1 U842 ( .A(n1157), .B(KEYINPUT17), .ZN(n1167) );
XOR2_X1 U843 ( .A(G131), .B(n1155), .Z(G33) );
AND3_X1 U844 ( .A1(n1157), .A2(n1003), .A3(n1158), .ZN(n1155) );
INV_X1 U845 ( .A(n1166), .ZN(n1158) );
NAND3_X1 U846 ( .A1(n998), .A2(n1169), .A3(n1010), .ZN(n1166) );
INV_X1 U847 ( .A(n989), .ZN(n1157) );
NAND2_X1 U848 ( .A1(n1022), .A2(n1170), .ZN(n989) );
NAND2_X1 U849 ( .A1(n1171), .A2(n1172), .ZN(G30) );
NAND2_X1 U850 ( .A1(n1154), .A2(n1173), .ZN(n1172) );
XOR2_X1 U851 ( .A(KEYINPUT60), .B(n1174), .Z(n1171) );
NOR2_X1 U852 ( .A1(n1154), .A2(n1173), .ZN(n1174) );
AND3_X1 U853 ( .A1(n1005), .A2(n1023), .A3(n1159), .ZN(n1154) );
AND4_X1 U854 ( .A1(n998), .A2(n1175), .A3(n1033), .A4(n1169), .ZN(n1159) );
XNOR2_X1 U855 ( .A(G101), .B(n1145), .ZN(G3) );
NAND3_X1 U856 ( .A1(n999), .A2(n1148), .A3(n1010), .ZN(n1145) );
XOR2_X1 U857 ( .A(G125), .B(n1153), .Z(G27) );
AND3_X1 U858 ( .A1(n1002), .A2(n1023), .A3(n1162), .ZN(n1153) );
AND3_X1 U859 ( .A1(n1009), .A2(n1169), .A3(n1003), .ZN(n1162) );
NAND2_X1 U860 ( .A1(n993), .A2(n1176), .ZN(n1169) );
NAND4_X1 U861 ( .A1(G953), .A2(G902), .A3(n1177), .A4(n1048), .ZN(n1176) );
INV_X1 U862 ( .A(G900), .ZN(n1048) );
XNOR2_X1 U863 ( .A(G122), .B(n1144), .ZN(G24) );
NAND4_X1 U864 ( .A1(n1178), .A2(n1014), .A3(n1160), .A4(n1032), .ZN(n1144) );
NOR2_X1 U865 ( .A1(n1033), .A2(n1179), .ZN(n1014) );
XNOR2_X1 U866 ( .A(G119), .B(n1147), .ZN(G21) );
NAND4_X1 U867 ( .A1(n1178), .A2(n999), .A3(n1175), .A4(n1033), .ZN(n1147) );
XNOR2_X1 U868 ( .A(G116), .B(n1143), .ZN(G18) );
NAND3_X1 U869 ( .A1(n1178), .A2(n1005), .A3(n1010), .ZN(n1143) );
NOR2_X1 U870 ( .A1(n1032), .A2(n1180), .ZN(n1005) );
NAND3_X1 U871 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(G15) );
NAND2_X1 U872 ( .A1(G113), .A2(n1184), .ZN(n1183) );
OR3_X1 U873 ( .A1(n1184), .A2(G113), .A3(n1146), .ZN(n1182) );
INV_X1 U874 ( .A(KEYINPUT12), .ZN(n1184) );
NAND2_X1 U875 ( .A1(n1185), .A2(n1146), .ZN(n1181) );
NAND3_X1 U876 ( .A1(n1010), .A2(n1178), .A3(n1003), .ZN(n1146) );
AND2_X1 U877 ( .A1(n1180), .A2(n1032), .ZN(n1003) );
AND2_X1 U878 ( .A1(n1002), .A2(n1186), .ZN(n1178) );
NOR2_X1 U879 ( .A1(n1024), .A2(n1007), .ZN(n1002) );
AND2_X1 U880 ( .A1(n1187), .A2(n1175), .ZN(n1010) );
XNOR2_X1 U881 ( .A(n1179), .B(KEYINPUT50), .ZN(n1175) );
NAND2_X1 U882 ( .A1(n1188), .A2(KEYINPUT12), .ZN(n1185) );
XNOR2_X1 U883 ( .A(G113), .B(KEYINPUT20), .ZN(n1188) );
XOR2_X1 U884 ( .A(n1142), .B(n1189), .Z(G12) );
XNOR2_X1 U885 ( .A(G110), .B(KEYINPUT15), .ZN(n1189) );
NAND3_X1 U886 ( .A1(n1009), .A2(n1148), .A3(n999), .ZN(n1142) );
NOR2_X1 U887 ( .A1(n1032), .A2(n1160), .ZN(n999) );
INV_X1 U888 ( .A(n1180), .ZN(n1160) );
XOR2_X1 U889 ( .A(n1039), .B(n1190), .Z(n1180) );
NOR2_X1 U890 ( .A1(G478), .A2(KEYINPUT49), .ZN(n1190) );
NOR2_X1 U891 ( .A1(n1097), .A2(G902), .ZN(n1039) );
XOR2_X1 U892 ( .A(n1191), .B(n1192), .Z(n1097) );
XNOR2_X1 U893 ( .A(n1173), .B(n1193), .ZN(n1192) );
XNOR2_X1 U894 ( .A(n1194), .B(G134), .ZN(n1193) );
XOR2_X1 U895 ( .A(n1195), .B(n1196), .Z(n1191) );
AND2_X1 U896 ( .A1(n1197), .A2(G217), .ZN(n1196) );
NAND2_X1 U897 ( .A1(n1198), .A2(n1199), .ZN(n1195) );
NAND2_X1 U898 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U899 ( .A(KEYINPUT57), .B(n1202), .Z(n1198) );
NOR2_X1 U900 ( .A1(n1200), .A2(n1201), .ZN(n1202) );
INV_X1 U901 ( .A(G107), .ZN(n1201) );
XNOR2_X1 U902 ( .A(n1203), .B(n1204), .ZN(n1200) );
XNOR2_X1 U903 ( .A(G116), .B(KEYINPUT23), .ZN(n1203) );
XOR2_X1 U904 ( .A(n1205), .B(n1106), .Z(n1032) );
INV_X1 U905 ( .A(G475), .ZN(n1106) );
OR2_X1 U906 ( .A1(n1103), .A2(G902), .ZN(n1205) );
XNOR2_X1 U907 ( .A(n1206), .B(n1207), .ZN(n1103) );
XOR2_X1 U908 ( .A(n1208), .B(n1209), .Z(n1206) );
NOR2_X1 U909 ( .A1(KEYINPUT44), .A2(n1210), .ZN(n1209) );
XNOR2_X1 U910 ( .A(G113), .B(n1204), .ZN(n1210) );
NAND2_X1 U911 ( .A1(n1211), .A2(n1212), .ZN(n1208) );
NAND2_X1 U912 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XOR2_X1 U913 ( .A(KEYINPUT43), .B(n1215), .Z(n1211) );
NOR2_X1 U914 ( .A1(n1213), .A2(n1214), .ZN(n1215) );
XOR2_X1 U915 ( .A(n1216), .B(n1217), .Z(n1214) );
XNOR2_X1 U916 ( .A(n1194), .B(G131), .ZN(n1217) );
NAND2_X1 U917 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
XOR2_X1 U918 ( .A(KEYINPUT59), .B(G214), .Z(n1219) );
XNOR2_X1 U919 ( .A(n1220), .B(n1221), .ZN(n1213) );
XNOR2_X1 U920 ( .A(KEYINPUT62), .B(n1222), .ZN(n1221) );
AND2_X1 U921 ( .A1(n1186), .A2(n998), .ZN(n1148) );
NOR2_X1 U922 ( .A1(n1035), .A2(n1007), .ZN(n998) );
INV_X1 U923 ( .A(n1012), .ZN(n1007) );
NAND2_X1 U924 ( .A1(G221), .A2(n1223), .ZN(n1012) );
INV_X1 U925 ( .A(n1024), .ZN(n1035) );
XOR2_X1 U926 ( .A(n1224), .B(n1124), .Z(n1024) );
INV_X1 U927 ( .A(G469), .ZN(n1124) );
NAND2_X1 U928 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XNOR2_X1 U929 ( .A(n1227), .B(n1228), .ZN(n1225) );
XNOR2_X1 U930 ( .A(n1229), .B(n1230), .ZN(n1227) );
NOR2_X1 U931 ( .A1(KEYINPUT22), .A2(n1126), .ZN(n1230) );
XOR2_X1 U932 ( .A(n1065), .B(n1231), .Z(n1126) );
XNOR2_X1 U933 ( .A(n1232), .B(n1233), .ZN(n1231) );
NOR2_X1 U934 ( .A1(G953), .A2(n1047), .ZN(n1233) );
INV_X1 U935 ( .A(G227), .ZN(n1047) );
NOR2_X1 U936 ( .A1(KEYINPUT41), .A2(n1234), .ZN(n1229) );
XOR2_X1 U937 ( .A(n1125), .B(n1057), .Z(n1234) );
XNOR2_X1 U938 ( .A(n1235), .B(n1236), .ZN(n1057) );
XNOR2_X1 U939 ( .A(G146), .B(n1237), .ZN(n1236) );
NAND2_X1 U940 ( .A1(KEYINPUT37), .A2(n1194), .ZN(n1237) );
INV_X1 U941 ( .A(G143), .ZN(n1194) );
NAND2_X1 U942 ( .A1(KEYINPUT46), .A2(n1173), .ZN(n1235) );
XNOR2_X1 U943 ( .A(G107), .B(n1238), .ZN(n1125) );
AND2_X1 U944 ( .A1(n1023), .A2(n1239), .ZN(n1186) );
NAND2_X1 U945 ( .A1(n993), .A2(n1240), .ZN(n1239) );
NAND4_X1 U946 ( .A1(G953), .A2(G902), .A3(n1177), .A4(n1074), .ZN(n1240) );
INV_X1 U947 ( .A(G898), .ZN(n1074) );
NAND3_X1 U948 ( .A1(n1177), .A2(n1016), .A3(G952), .ZN(n993) );
NAND2_X1 U949 ( .A1(G237), .A2(G234), .ZN(n1177) );
NOR2_X1 U950 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
INV_X1 U951 ( .A(n1170), .ZN(n1021) );
NAND2_X1 U952 ( .A1(G214), .A2(n1241), .ZN(n1170) );
NOR2_X1 U953 ( .A1(n1036), .A2(n1242), .ZN(n1022) );
AND2_X1 U954 ( .A1(n1243), .A2(n1038), .ZN(n1242) );
XNOR2_X1 U955 ( .A(KEYINPUT8), .B(n1139), .ZN(n1243) );
NOR2_X1 U956 ( .A1(n1038), .A2(n1037), .ZN(n1036) );
INV_X1 U957 ( .A(n1139), .ZN(n1037) );
NAND2_X1 U958 ( .A1(G210), .A2(n1241), .ZN(n1139) );
NAND2_X1 U959 ( .A1(n1244), .A2(n1226), .ZN(n1241) );
INV_X1 U960 ( .A(G237), .ZN(n1244) );
NAND2_X1 U961 ( .A1(n1245), .A2(n1246), .ZN(n1038) );
XNOR2_X1 U962 ( .A(n1133), .B(n1247), .ZN(n1246) );
XOR2_X1 U963 ( .A(n1137), .B(KEYINPUT19), .Z(n1247) );
XOR2_X1 U964 ( .A(n1248), .B(n1249), .Z(n1137) );
XNOR2_X1 U965 ( .A(G125), .B(n1250), .ZN(n1248) );
NOR2_X1 U966 ( .A1(G953), .A2(n1073), .ZN(n1250) );
INV_X1 U967 ( .A(G224), .ZN(n1073) );
INV_X1 U968 ( .A(n1136), .ZN(n1133) );
NAND2_X1 U969 ( .A1(n1251), .A2(n1252), .ZN(n1136) );
NAND2_X1 U970 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
INV_X1 U971 ( .A(n1083), .ZN(n1254) );
XOR2_X1 U972 ( .A(KEYINPUT38), .B(n1255), .Z(n1253) );
NAND2_X1 U973 ( .A1(n1255), .A2(n1083), .ZN(n1251) );
XNOR2_X1 U974 ( .A(n1256), .B(n1238), .ZN(n1083) );
XNOR2_X1 U975 ( .A(n1257), .B(n1207), .ZN(n1238) );
XOR2_X1 U976 ( .A(G104), .B(KEYINPUT36), .Z(n1207) );
NAND2_X1 U977 ( .A1(KEYINPUT30), .A2(G107), .ZN(n1256) );
XOR2_X1 U978 ( .A(n1258), .B(n1086), .Z(n1255) );
NAND2_X1 U979 ( .A1(KEYINPUT45), .A2(n1085), .ZN(n1258) );
XOR2_X1 U980 ( .A(G110), .B(n1204), .Z(n1085) );
XOR2_X1 U981 ( .A(G122), .B(KEYINPUT39), .Z(n1204) );
XNOR2_X1 U982 ( .A(G902), .B(KEYINPUT61), .ZN(n1245) );
NOR2_X1 U983 ( .A1(n1179), .A2(n1187), .ZN(n1009) );
INV_X1 U984 ( .A(n1033), .ZN(n1187) );
XOR2_X1 U985 ( .A(n1259), .B(n1093), .Z(n1033) );
NAND2_X1 U986 ( .A1(G217), .A2(n1223), .ZN(n1093) );
NAND2_X1 U987 ( .A1(G234), .A2(n1226), .ZN(n1223) );
NAND2_X1 U988 ( .A1(n1090), .A2(n1226), .ZN(n1259) );
XOR2_X1 U989 ( .A(n1260), .B(n1261), .Z(n1090) );
XOR2_X1 U990 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U991 ( .A(n1264), .B(n1265), .Z(n1263) );
NOR2_X1 U992 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XOR2_X1 U993 ( .A(n1268), .B(KEYINPUT9), .Z(n1267) );
NAND2_X1 U994 ( .A1(n1269), .A2(n1232), .ZN(n1268) );
NOR2_X1 U995 ( .A1(n1269), .A2(n1232), .ZN(n1266) );
INV_X1 U996 ( .A(G110), .ZN(n1232) );
XNOR2_X1 U997 ( .A(G119), .B(n1270), .ZN(n1269) );
XNOR2_X1 U998 ( .A(KEYINPUT5), .B(n1173), .ZN(n1270) );
INV_X1 U999 ( .A(G128), .ZN(n1173) );
NAND2_X1 U1000 ( .A1(KEYINPUT11), .A2(n1220), .ZN(n1264) );
XOR2_X1 U1001 ( .A(G125), .B(n1065), .Z(n1220) );
XNOR2_X1 U1002 ( .A(n1163), .B(KEYINPUT6), .ZN(n1065) );
INV_X1 U1003 ( .A(G140), .ZN(n1163) );
NAND2_X1 U1004 ( .A1(G221), .A2(n1197), .ZN(n1262) );
AND2_X1 U1005 ( .A1(G234), .A2(n1016), .ZN(n1197) );
INV_X1 U1006 ( .A(G953), .ZN(n1016) );
XNOR2_X1 U1007 ( .A(G137), .B(n1271), .ZN(n1260) );
XNOR2_X1 U1008 ( .A(KEYINPUT40), .B(n1222), .ZN(n1271) );
INV_X1 U1009 ( .A(G146), .ZN(n1222) );
XNOR2_X1 U1010 ( .A(n1031), .B(KEYINPUT24), .ZN(n1179) );
XOR2_X1 U1011 ( .A(n1272), .B(n1115), .Z(n1031) );
INV_X1 U1012 ( .A(G472), .ZN(n1115) );
NAND2_X1 U1013 ( .A1(n1273), .A2(n1226), .ZN(n1272) );
INV_X1 U1014 ( .A(G902), .ZN(n1226) );
XOR2_X1 U1015 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U1016 ( .A(n1112), .B(n1276), .Z(n1275) );
NOR2_X1 U1017 ( .A1(KEYINPUT28), .A2(n1086), .ZN(n1276) );
XNOR2_X1 U1018 ( .A(G113), .B(n1277), .ZN(n1086) );
XNOR2_X1 U1019 ( .A(n1278), .B(G116), .ZN(n1277) );
INV_X1 U1020 ( .A(G119), .ZN(n1278) );
XNOR2_X1 U1021 ( .A(n1249), .B(n1279), .ZN(n1112) );
XNOR2_X1 U1022 ( .A(KEYINPUT34), .B(n1228), .ZN(n1279) );
INV_X1 U1023 ( .A(n1120), .ZN(n1228) );
XOR2_X1 U1024 ( .A(n1280), .B(n1281), .Z(n1120) );
INV_X1 U1025 ( .A(n1063), .ZN(n1281) );
XOR2_X1 U1026 ( .A(G131), .B(KEYINPUT10), .Z(n1063) );
XNOR2_X1 U1027 ( .A(G134), .B(G137), .ZN(n1280) );
XOR2_X1 U1028 ( .A(G128), .B(n1282), .Z(n1249) );
NOR2_X1 U1029 ( .A1(KEYINPUT21), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U1030 ( .A(G143), .B(G146), .ZN(n1283) );
XNOR2_X1 U1031 ( .A(KEYINPUT18), .B(n1284), .ZN(n1274) );
NOR2_X1 U1032 ( .A1(KEYINPUT54), .A2(n1113), .ZN(n1284) );
XNOR2_X1 U1033 ( .A(n1285), .B(n1257), .ZN(n1113) );
XNOR2_X1 U1034 ( .A(G101), .B(KEYINPUT13), .ZN(n1257) );
NAND2_X1 U1035 ( .A1(G210), .A2(n1218), .ZN(n1285) );
NOR2_X1 U1036 ( .A1(G953), .A2(G237), .ZN(n1218) );
endmodule


