//Key = 1110010100011011111001110110000000010110111101101100101111111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345;

XNOR2_X1 U742 ( .A(G107), .B(n1033), .ZN(G9) );
NOR2_X1 U743 ( .A1(n1034), .A2(n1035), .ZN(G75) );
NOR3_X1 U744 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
XOR2_X1 U745 ( .A(KEYINPUT54), .B(n1039), .Z(n1038) );
NOR2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR4_X1 U747 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1041) );
NOR3_X1 U748 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1042) );
NOR2_X1 U749 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
XNOR2_X1 U750 ( .A(KEYINPUT52), .B(n1051), .ZN(n1050) );
NOR3_X1 U751 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1047) );
NOR2_X1 U752 ( .A1(n1055), .A2(n1056), .ZN(n1046) );
INV_X1 U753 ( .A(n1057), .ZN(n1056) );
XNOR2_X1 U754 ( .A(n1058), .B(KEYINPUT36), .ZN(n1055) );
NOR3_X1 U755 ( .A1(n1045), .A2(n1059), .A3(n1053), .ZN(n1040) );
NOR2_X1 U756 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U757 ( .A1(n1062), .A2(n1051), .ZN(n1061) );
NOR2_X1 U758 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U759 ( .A1(n1065), .A2(n1044), .ZN(n1064) );
NOR2_X1 U760 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U762 ( .A1(n1070), .A2(n1043), .ZN(n1063) );
NOR2_X1 U763 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR3_X1 U764 ( .A1(n1044), .A2(n1073), .A3(n1043), .ZN(n1060) );
INV_X1 U765 ( .A(n1074), .ZN(n1043) );
NAND3_X1 U766 ( .A1(n1075), .A2(n1076), .A3(G952), .ZN(n1036) );
NOR3_X1 U767 ( .A1(n1077), .A2(G953), .A3(n1078), .ZN(n1034) );
INV_X1 U768 ( .A(n1075), .ZN(n1078) );
NAND4_X1 U769 ( .A1(n1079), .A2(n1080), .A3(n1058), .A4(n1081), .ZN(n1075) );
NOR4_X1 U770 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1081) );
XNOR2_X1 U771 ( .A(G469), .B(n1086), .ZN(n1085) );
NOR2_X1 U772 ( .A1(n1087), .A2(KEYINPUT32), .ZN(n1086) );
XNOR2_X1 U773 ( .A(n1088), .B(KEYINPUT41), .ZN(n1084) );
XOR2_X1 U774 ( .A(n1089), .B(n1090), .Z(n1083) );
NAND2_X1 U775 ( .A1(KEYINPUT15), .A2(n1091), .ZN(n1089) );
XNOR2_X1 U776 ( .A(G478), .B(n1092), .ZN(n1080) );
NAND2_X1 U777 ( .A1(KEYINPUT57), .A2(n1093), .ZN(n1092) );
XNOR2_X1 U778 ( .A(G952), .B(KEYINPUT61), .ZN(n1077) );
XOR2_X1 U779 ( .A(n1094), .B(n1095), .Z(G72) );
XOR2_X1 U780 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U782 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U783 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U784 ( .A1(KEYINPUT50), .A2(n1104), .ZN(n1103) );
XOR2_X1 U785 ( .A(n1105), .B(KEYINPUT9), .Z(n1100) );
NAND2_X1 U786 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND4_X1 U787 ( .A1(n1108), .A2(n1109), .A3(n1110), .A4(n1111), .ZN(n1107) );
XOR2_X1 U788 ( .A(n1112), .B(KEYINPUT33), .Z(n1106) );
NAND2_X1 U789 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND3_X1 U790 ( .A1(n1110), .A2(n1111), .A3(n1109), .ZN(n1114) );
NAND2_X1 U791 ( .A1(n1115), .A2(n1116), .ZN(n1109) );
XNOR2_X1 U792 ( .A(n1117), .B(n1118), .ZN(n1115) );
AND2_X1 U793 ( .A1(n1119), .A2(KEYINPUT58), .ZN(n1118) );
NAND3_X1 U794 ( .A1(G131), .A2(n1119), .A3(n1120), .ZN(n1110) );
XNOR2_X1 U795 ( .A(KEYINPUT58), .B(G134), .ZN(n1120) );
XNOR2_X1 U796 ( .A(n1121), .B(KEYINPUT18), .ZN(n1098) );
NAND2_X1 U797 ( .A1(n1122), .A2(n1076), .ZN(n1096) );
NAND2_X1 U798 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XNOR2_X1 U799 ( .A(KEYINPUT35), .B(n1125), .ZN(n1124) );
NAND2_X1 U800 ( .A1(G953), .A2(n1126), .ZN(n1094) );
NAND2_X1 U801 ( .A1(G900), .A2(G227), .ZN(n1126) );
NAND2_X1 U802 ( .A1(n1127), .A2(n1128), .ZN(G69) );
OR3_X1 U803 ( .A1(n1129), .A2(KEYINPUT19), .A3(n1130), .ZN(n1128) );
NAND2_X1 U804 ( .A1(n1130), .A2(n1131), .ZN(n1127) );
NAND2_X1 U805 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
OR2_X1 U806 ( .A1(n1134), .A2(KEYINPUT13), .ZN(n1133) );
NAND2_X1 U807 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
OR2_X1 U808 ( .A1(KEYINPUT13), .A2(KEYINPUT19), .ZN(n1135) );
INV_X1 U809 ( .A(n1129), .ZN(n1134) );
NAND2_X1 U810 ( .A1(G953), .A2(n1136), .ZN(n1129) );
XOR2_X1 U811 ( .A(KEYINPUT7), .B(n1137), .Z(n1136) );
AND2_X1 U812 ( .A1(G224), .A2(G898), .ZN(n1137) );
XNOR2_X1 U813 ( .A(n1138), .B(n1139), .ZN(n1130) );
NOR2_X1 U814 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XNOR2_X1 U815 ( .A(n1142), .B(n1143), .ZN(n1141) );
NAND2_X1 U816 ( .A1(n1076), .A2(n1144), .ZN(n1138) );
NOR2_X1 U817 ( .A1(n1145), .A2(n1146), .ZN(G66) );
NOR3_X1 U818 ( .A1(n1090), .A2(n1147), .A3(n1148), .ZN(n1146) );
NOR3_X1 U819 ( .A1(n1149), .A2(n1091), .A3(n1150), .ZN(n1148) );
INV_X1 U820 ( .A(n1151), .ZN(n1149) );
NOR2_X1 U821 ( .A1(n1152), .A2(n1151), .ZN(n1147) );
NOR2_X1 U822 ( .A1(n1153), .A2(n1091), .ZN(n1152) );
NOR2_X1 U823 ( .A1(n1145), .A2(n1154), .ZN(G63) );
XOR2_X1 U824 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U825 ( .A1(n1157), .A2(KEYINPUT39), .ZN(n1156) );
NAND2_X1 U826 ( .A1(n1158), .A2(G478), .ZN(n1155) );
NOR2_X1 U827 ( .A1(n1145), .A2(n1159), .ZN(G60) );
XNOR2_X1 U828 ( .A(n1160), .B(n1161), .ZN(n1159) );
AND2_X1 U829 ( .A1(G475), .A2(n1158), .ZN(n1161) );
XNOR2_X1 U830 ( .A(G104), .B(n1162), .ZN(G6) );
NOR2_X1 U831 ( .A1(n1145), .A2(n1163), .ZN(G57) );
XOR2_X1 U832 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U833 ( .A(n1166), .B(n1167), .Z(n1165) );
AND2_X1 U834 ( .A1(G472), .A2(n1158), .ZN(n1166) );
XOR2_X1 U835 ( .A(n1168), .B(n1169), .Z(n1164) );
XNOR2_X1 U836 ( .A(KEYINPUT37), .B(n1170), .ZN(n1169) );
NOR2_X1 U837 ( .A1(KEYINPUT20), .A2(n1171), .ZN(n1170) );
NOR2_X1 U838 ( .A1(n1145), .A2(n1172), .ZN(G54) );
XOR2_X1 U839 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U840 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U841 ( .A1(n1177), .A2(n1150), .ZN(n1175) );
XOR2_X1 U842 ( .A(KEYINPUT30), .B(KEYINPUT12), .Z(n1173) );
NOR2_X1 U843 ( .A1(n1145), .A2(n1178), .ZN(G51) );
XOR2_X1 U844 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U845 ( .A(KEYINPUT22), .B(n1181), .Z(n1180) );
NOR2_X1 U846 ( .A1(n1182), .A2(n1150), .ZN(n1181) );
INV_X1 U847 ( .A(n1158), .ZN(n1150) );
NOR2_X1 U848 ( .A1(n1183), .A2(n1153), .ZN(n1158) );
INV_X1 U849 ( .A(n1037), .ZN(n1153) );
NAND3_X1 U850 ( .A1(n1184), .A2(n1125), .A3(n1123), .ZN(n1037) );
AND4_X1 U851 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1123) );
NOR4_X1 U852 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1188) );
NOR2_X1 U853 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NOR2_X1 U854 ( .A1(n1195), .A2(n1196), .ZN(n1193) );
XNOR2_X1 U855 ( .A(n1057), .B(KEYINPUT40), .ZN(n1196) );
AND4_X1 U856 ( .A1(KEYINPUT4), .A2(n1197), .A3(n1049), .A4(n1198), .ZN(n1190) );
NOR2_X1 U857 ( .A1(KEYINPUT4), .A2(n1199), .ZN(n1189) );
INV_X1 U858 ( .A(n1144), .ZN(n1184) );
NAND2_X1 U859 ( .A1(n1200), .A2(n1201), .ZN(n1144) );
AND4_X1 U860 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1162), .ZN(n1201) );
NAND3_X1 U861 ( .A1(n1205), .A2(n1206), .A3(n1072), .ZN(n1162) );
AND4_X1 U862 ( .A1(n1033), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1200) );
NAND3_X1 U863 ( .A1(n1071), .A2(n1206), .A3(n1205), .ZN(n1033) );
XOR2_X1 U864 ( .A(n1210), .B(n1211), .Z(n1179) );
NOR2_X1 U865 ( .A1(n1076), .A2(G952), .ZN(n1145) );
XNOR2_X1 U866 ( .A(n1191), .B(n1212), .ZN(G48) );
NAND2_X1 U867 ( .A1(KEYINPUT38), .A2(G146), .ZN(n1212) );
AND3_X1 U868 ( .A1(n1072), .A2(n1213), .A3(n1214), .ZN(n1191) );
XNOR2_X1 U869 ( .A(G143), .B(n1199), .ZN(G45) );
NAND3_X1 U870 ( .A1(n1195), .A2(n1198), .A3(n1197), .ZN(n1199) );
NOR3_X1 U871 ( .A1(n1215), .A2(n1079), .A3(n1073), .ZN(n1197) );
XNOR2_X1 U872 ( .A(G140), .B(n1216), .ZN(G42) );
NAND3_X1 U873 ( .A1(n1217), .A2(n1057), .A3(KEYINPUT5), .ZN(n1216) );
INV_X1 U874 ( .A(n1194), .ZN(n1217) );
NAND3_X1 U875 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(G39) );
NAND2_X1 U876 ( .A1(KEYINPUT29), .A2(n1119), .ZN(n1220) );
NAND3_X1 U877 ( .A1(G137), .A2(n1221), .A3(n1187), .ZN(n1219) );
NAND2_X1 U878 ( .A1(n1222), .A2(n1223), .ZN(n1218) );
NAND2_X1 U879 ( .A1(n1224), .A2(n1221), .ZN(n1223) );
INV_X1 U880 ( .A(KEYINPUT29), .ZN(n1221) );
XNOR2_X1 U881 ( .A(G137), .B(KEYINPUT55), .ZN(n1224) );
INV_X1 U882 ( .A(n1187), .ZN(n1222) );
NAND3_X1 U883 ( .A1(n1214), .A2(n1058), .A3(n1225), .ZN(n1187) );
XNOR2_X1 U884 ( .A(G134), .B(n1125), .ZN(G36) );
NAND4_X1 U885 ( .A1(n1195), .A2(n1198), .A3(n1058), .A4(n1071), .ZN(n1125) );
XNOR2_X1 U886 ( .A(n1116), .B(n1226), .ZN(G33) );
NOR2_X1 U887 ( .A1(n1049), .A2(n1194), .ZN(n1226) );
NAND3_X1 U888 ( .A1(n1198), .A2(n1058), .A3(n1072), .ZN(n1194) );
INV_X1 U889 ( .A(n1051), .ZN(n1058) );
NAND2_X1 U890 ( .A1(n1227), .A2(n1052), .ZN(n1051) );
INV_X1 U891 ( .A(n1054), .ZN(n1227) );
INV_X1 U892 ( .A(n1228), .ZN(n1198) );
XNOR2_X1 U893 ( .A(G128), .B(n1185), .ZN(G30) );
NAND3_X1 U894 ( .A1(n1071), .A2(n1213), .A3(n1214), .ZN(n1185) );
NOR3_X1 U895 ( .A1(n1229), .A2(n1230), .A3(n1228), .ZN(n1214) );
NAND2_X1 U896 ( .A1(n1067), .A2(n1231), .ZN(n1228) );
XNOR2_X1 U897 ( .A(G101), .B(n1209), .ZN(G3) );
NAND3_X1 U898 ( .A1(n1195), .A2(n1205), .A3(n1225), .ZN(n1209) );
XNOR2_X1 U899 ( .A(G125), .B(n1186), .ZN(G27) );
NAND4_X1 U900 ( .A1(n1074), .A2(n1057), .A3(n1232), .A4(n1072), .ZN(n1186) );
AND2_X1 U901 ( .A1(n1231), .A2(n1213), .ZN(n1232) );
NAND2_X1 U902 ( .A1(n1045), .A2(n1233), .ZN(n1231) );
NAND2_X1 U903 ( .A1(n1121), .A2(n1234), .ZN(n1233) );
NOR2_X1 U904 ( .A1(n1076), .A2(G900), .ZN(n1121) );
XNOR2_X1 U905 ( .A(G122), .B(n1208), .ZN(G24) );
NAND4_X1 U906 ( .A1(n1074), .A2(n1206), .A3(n1235), .A4(n1236), .ZN(n1208) );
NOR2_X1 U907 ( .A1(n1079), .A2(n1215), .ZN(n1235) );
INV_X1 U908 ( .A(n1053), .ZN(n1206) );
NAND2_X1 U909 ( .A1(n1230), .A2(n1229), .ZN(n1053) );
XNOR2_X1 U910 ( .A(G119), .B(n1204), .ZN(G21) );
NAND4_X1 U911 ( .A1(n1225), .A2(n1074), .A3(n1237), .A4(n1236), .ZN(n1204) );
NOR2_X1 U912 ( .A1(n1230), .A2(n1229), .ZN(n1237) );
INV_X1 U913 ( .A(n1088), .ZN(n1229) );
XNOR2_X1 U914 ( .A(n1238), .B(n1239), .ZN(G18) );
NAND2_X1 U915 ( .A1(KEYINPUT2), .A2(n1207), .ZN(n1238) );
NAND2_X1 U916 ( .A1(n1240), .A2(n1071), .ZN(n1207) );
NOR2_X1 U917 ( .A1(n1241), .A2(n1215), .ZN(n1071) );
XNOR2_X1 U918 ( .A(n1203), .B(n1242), .ZN(G15) );
XOR2_X1 U919 ( .A(KEYINPUT6), .B(G113), .Z(n1242) );
NAND2_X1 U920 ( .A1(n1240), .A2(n1072), .ZN(n1203) );
AND2_X1 U921 ( .A1(n1243), .A2(n1241), .ZN(n1072) );
XNOR2_X1 U922 ( .A(KEYINPUT42), .B(n1215), .ZN(n1243) );
AND3_X1 U923 ( .A1(n1195), .A2(n1236), .A3(n1074), .ZN(n1240) );
NOR2_X1 U924 ( .A1(n1068), .A2(n1082), .ZN(n1074) );
INV_X1 U925 ( .A(n1069), .ZN(n1082) );
INV_X1 U926 ( .A(n1049), .ZN(n1195) );
NAND2_X1 U927 ( .A1(n1230), .A2(n1088), .ZN(n1049) );
XNOR2_X1 U928 ( .A(G110), .B(n1202), .ZN(G12) );
NAND3_X1 U929 ( .A1(n1057), .A2(n1205), .A3(n1225), .ZN(n1202) );
INV_X1 U930 ( .A(n1044), .ZN(n1225) );
NAND2_X1 U931 ( .A1(n1215), .A2(n1079), .ZN(n1044) );
INV_X1 U932 ( .A(n1241), .ZN(n1079) );
XNOR2_X1 U933 ( .A(n1244), .B(G475), .ZN(n1241) );
NAND2_X1 U934 ( .A1(n1160), .A2(n1183), .ZN(n1244) );
XNOR2_X1 U935 ( .A(n1245), .B(n1246), .ZN(n1160) );
XOR2_X1 U936 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U937 ( .A(n1249), .B(n1250), .Z(n1248) );
NAND2_X1 U938 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U939 ( .A1(G113), .A2(n1253), .ZN(n1252) );
XOR2_X1 U940 ( .A(KEYINPUT45), .B(n1254), .Z(n1251) );
NOR2_X1 U941 ( .A1(G113), .A2(n1253), .ZN(n1254) );
NAND2_X1 U942 ( .A1(n1255), .A2(n1256), .ZN(n1249) );
NAND4_X1 U943 ( .A1(G143), .A2(G214), .A3(n1257), .A4(n1076), .ZN(n1256) );
XOR2_X1 U944 ( .A(n1258), .B(KEYINPUT53), .Z(n1255) );
NAND2_X1 U945 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NAND3_X1 U946 ( .A1(n1257), .A2(n1076), .A3(G214), .ZN(n1260) );
XOR2_X1 U947 ( .A(n1261), .B(n1262), .Z(n1245) );
XNOR2_X1 U948 ( .A(G146), .B(n1116), .ZN(n1262) );
XNOR2_X1 U949 ( .A(G125), .B(n1263), .ZN(n1261) );
NOR2_X1 U950 ( .A1(KEYINPUT8), .A2(n1264), .ZN(n1263) );
XOR2_X1 U951 ( .A(n1102), .B(KEYINPUT17), .Z(n1264) );
XNOR2_X1 U952 ( .A(n1265), .B(n1093), .ZN(n1215) );
OR2_X1 U953 ( .A1(G902), .A2(n1157), .ZN(n1093) );
AND2_X1 U954 ( .A1(n1266), .A2(n1267), .ZN(n1157) );
NAND4_X1 U955 ( .A1(n1268), .A2(G217), .A3(G234), .A4(n1269), .ZN(n1267) );
XNOR2_X1 U956 ( .A(n1270), .B(n1271), .ZN(n1269) );
NAND2_X1 U957 ( .A1(n1272), .A2(n1273), .ZN(n1266) );
NAND3_X1 U958 ( .A1(n1268), .A2(G234), .A3(G217), .ZN(n1273) );
XNOR2_X1 U959 ( .A(G953), .B(KEYINPUT34), .ZN(n1268) );
XNOR2_X1 U960 ( .A(n1270), .B(n1274), .ZN(n1272) );
INV_X1 U961 ( .A(n1271), .ZN(n1274) );
XOR2_X1 U962 ( .A(G107), .B(n1275), .Z(n1271) );
XNOR2_X1 U963 ( .A(n1117), .B(G122), .ZN(n1275) );
XNOR2_X1 U964 ( .A(n1276), .B(n1277), .ZN(n1270) );
NAND2_X1 U965 ( .A1(KEYINPUT21), .A2(n1239), .ZN(n1277) );
NAND2_X1 U966 ( .A1(KEYINPUT60), .A2(n1278), .ZN(n1276) );
XNOR2_X1 U967 ( .A(n1259), .B(G128), .ZN(n1278) );
INV_X1 U968 ( .A(G143), .ZN(n1259) );
NAND2_X1 U969 ( .A1(KEYINPUT56), .A2(G478), .ZN(n1265) );
AND2_X1 U970 ( .A1(n1236), .A2(n1067), .ZN(n1205) );
AND2_X1 U971 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U972 ( .A1(G221), .A2(n1279), .ZN(n1069) );
XNOR2_X1 U973 ( .A(n1087), .B(n1177), .ZN(n1068) );
INV_X1 U974 ( .A(G469), .ZN(n1177) );
AND3_X1 U975 ( .A1(n1280), .A2(n1281), .A3(n1183), .ZN(n1087) );
OR2_X1 U976 ( .A1(n1176), .A2(KEYINPUT44), .ZN(n1281) );
XNOR2_X1 U977 ( .A(n1282), .B(n1283), .ZN(n1176) );
NAND3_X1 U978 ( .A1(n1282), .A2(n1283), .A3(KEYINPUT44), .ZN(n1280) );
XOR2_X1 U979 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U980 ( .A(n1286), .B(n1113), .ZN(n1285) );
INV_X1 U981 ( .A(n1108), .ZN(n1113) );
XNOR2_X1 U982 ( .A(n1287), .B(n1288), .ZN(n1108) );
NAND2_X1 U983 ( .A1(KEYINPUT49), .A2(n1289), .ZN(n1287) );
XNOR2_X1 U984 ( .A(G146), .B(n1290), .ZN(n1289) );
NAND2_X1 U985 ( .A1(KEYINPUT25), .A2(G143), .ZN(n1290) );
XOR2_X1 U986 ( .A(n1291), .B(KEYINPUT24), .Z(n1284) );
XNOR2_X1 U987 ( .A(n1102), .B(n1292), .ZN(n1282) );
XOR2_X1 U988 ( .A(G110), .B(n1293), .Z(n1292) );
AND2_X1 U989 ( .A1(n1076), .A2(G227), .ZN(n1293) );
AND2_X1 U990 ( .A1(n1213), .A2(n1294), .ZN(n1236) );
NAND2_X1 U991 ( .A1(n1045), .A2(n1295), .ZN(n1294) );
NAND2_X1 U992 ( .A1(n1140), .A2(n1234), .ZN(n1295) );
AND2_X1 U993 ( .A1(n1296), .A2(n1297), .ZN(n1234) );
XNOR2_X1 U994 ( .A(G902), .B(KEYINPUT59), .ZN(n1296) );
NOR2_X1 U995 ( .A1(n1076), .A2(G898), .ZN(n1140) );
NAND3_X1 U996 ( .A1(n1297), .A2(n1076), .A3(G952), .ZN(n1045) );
NAND2_X1 U997 ( .A1(G237), .A2(G234), .ZN(n1297) );
INV_X1 U998 ( .A(n1073), .ZN(n1213) );
NAND2_X1 U999 ( .A1(n1054), .A2(n1052), .ZN(n1073) );
NAND2_X1 U1000 ( .A1(G214), .A2(n1298), .ZN(n1052) );
XOR2_X1 U1001 ( .A(n1299), .B(n1182), .Z(n1054) );
NAND2_X1 U1002 ( .A1(G210), .A2(n1298), .ZN(n1182) );
NAND2_X1 U1003 ( .A1(n1257), .A2(n1183), .ZN(n1298) );
NAND2_X1 U1004 ( .A1(n1300), .A2(n1183), .ZN(n1299) );
XOR2_X1 U1005 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1006 ( .A(n1210), .B(n1303), .Z(n1302) );
NOR2_X1 U1007 ( .A1(KEYINPUT51), .A2(n1211), .ZN(n1303) );
XOR2_X1 U1008 ( .A(n1304), .B(n1305), .Z(n1210) );
XOR2_X1 U1009 ( .A(n1306), .B(n1307), .Z(n1305) );
XNOR2_X1 U1010 ( .A(KEYINPUT46), .B(n1104), .ZN(n1307) );
INV_X1 U1011 ( .A(G125), .ZN(n1104) );
AND2_X1 U1012 ( .A1(n1076), .A2(G224), .ZN(n1306) );
XOR2_X1 U1013 ( .A(n1142), .B(n1308), .Z(n1304) );
NOR2_X1 U1014 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
NOR2_X1 U1015 ( .A1(KEYINPUT48), .A2(n1311), .ZN(n1310) );
NOR2_X1 U1016 ( .A1(KEYINPUT27), .A2(n1143), .ZN(n1309) );
INV_X1 U1017 ( .A(n1311), .ZN(n1143) );
XNOR2_X1 U1018 ( .A(n1312), .B(n1313), .ZN(n1311) );
XNOR2_X1 U1019 ( .A(n1253), .B(G110), .ZN(n1313) );
INV_X1 U1020 ( .A(G122), .ZN(n1253) );
XNOR2_X1 U1021 ( .A(KEYINPUT62), .B(KEYINPUT43), .ZN(n1312) );
XOR2_X1 U1022 ( .A(n1314), .B(n1286), .Z(n1142) );
XNOR2_X1 U1023 ( .A(n1315), .B(n1247), .ZN(n1286) );
XOR2_X1 U1024 ( .A(G104), .B(KEYINPUT31), .Z(n1247) );
XNOR2_X1 U1025 ( .A(G107), .B(G101), .ZN(n1315) );
XNOR2_X1 U1026 ( .A(KEYINPUT23), .B(KEYINPUT1), .ZN(n1301) );
NOR2_X1 U1027 ( .A1(n1088), .A2(n1230), .ZN(n1057) );
XOR2_X1 U1028 ( .A(n1090), .B(n1091), .Z(n1230) );
NAND2_X1 U1029 ( .A1(G217), .A2(n1279), .ZN(n1091) );
NAND2_X1 U1030 ( .A1(G234), .A2(n1183), .ZN(n1279) );
NOR2_X1 U1031 ( .A1(n1151), .A2(G902), .ZN(n1090) );
XNOR2_X1 U1032 ( .A(n1316), .B(n1317), .ZN(n1151) );
NOR2_X1 U1033 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
XOR2_X1 U1034 ( .A(n1320), .B(KEYINPUT63), .Z(n1319) );
NAND2_X1 U1035 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NOR2_X1 U1036 ( .A1(n1322), .A2(n1321), .ZN(n1318) );
XNOR2_X1 U1037 ( .A(G146), .B(n1323), .ZN(n1321) );
NAND2_X1 U1038 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
NAND2_X1 U1039 ( .A1(n1102), .A2(G125), .ZN(n1325) );
XOR2_X1 U1040 ( .A(KEYINPUT26), .B(n1326), .Z(n1324) );
NOR2_X1 U1041 ( .A1(G125), .A2(n1102), .ZN(n1326) );
XNOR2_X1 U1042 ( .A(G140), .B(KEYINPUT3), .ZN(n1102) );
XNOR2_X1 U1043 ( .A(n1327), .B(n1328), .ZN(n1322) );
XOR2_X1 U1044 ( .A(G119), .B(G110), .Z(n1328) );
NAND2_X1 U1045 ( .A1(KEYINPUT0), .A2(G128), .ZN(n1327) );
NAND2_X1 U1046 ( .A1(KEYINPUT14), .A2(n1329), .ZN(n1316) );
XNOR2_X1 U1047 ( .A(n1119), .B(n1330), .ZN(n1329) );
AND3_X1 U1048 ( .A1(G221), .A2(n1076), .A3(G234), .ZN(n1330) );
XNOR2_X1 U1049 ( .A(n1331), .B(G472), .ZN(n1088) );
NAND2_X1 U1050 ( .A1(n1332), .A2(n1183), .ZN(n1331) );
INV_X1 U1051 ( .A(G902), .ZN(n1183) );
XOR2_X1 U1052 ( .A(n1333), .B(n1334), .Z(n1332) );
NAND2_X1 U1053 ( .A1(KEYINPUT16), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1054 ( .A(KEYINPUT47), .B(n1167), .Z(n1335) );
XOR2_X1 U1055 ( .A(n1211), .B(n1336), .Z(n1167) );
XOR2_X1 U1056 ( .A(n1314), .B(n1291), .Z(n1336) );
XOR2_X1 U1057 ( .A(n1337), .B(KEYINPUT10), .Z(n1291) );
NAND3_X1 U1058 ( .A1(n1338), .A2(n1339), .A3(n1111), .ZN(n1337) );
NAND3_X1 U1059 ( .A1(G131), .A2(n1117), .A3(G137), .ZN(n1111) );
INV_X1 U1060 ( .A(G134), .ZN(n1117) );
NAND2_X1 U1061 ( .A1(n1340), .A2(n1119), .ZN(n1339) );
INV_X1 U1062 ( .A(G137), .ZN(n1119) );
XNOR2_X1 U1063 ( .A(G131), .B(G134), .ZN(n1340) );
NAND3_X1 U1064 ( .A1(G134), .A2(n1116), .A3(G137), .ZN(n1338) );
INV_X1 U1065 ( .A(G131), .ZN(n1116) );
XNOR2_X1 U1066 ( .A(G113), .B(n1341), .ZN(n1314) );
XNOR2_X1 U1067 ( .A(G119), .B(n1239), .ZN(n1341) );
INV_X1 U1068 ( .A(G116), .ZN(n1239) );
XNOR2_X1 U1069 ( .A(n1342), .B(n1288), .ZN(n1211) );
XOR2_X1 U1070 ( .A(G128), .B(KEYINPUT28), .Z(n1288) );
XNOR2_X1 U1071 ( .A(G143), .B(G146), .ZN(n1342) );
NAND2_X1 U1072 ( .A1(n1343), .A2(n1344), .ZN(n1333) );
NAND2_X1 U1073 ( .A1(n1168), .A2(n1171), .ZN(n1344) );
XOR2_X1 U1074 ( .A(KEYINPUT11), .B(n1345), .Z(n1343) );
NOR2_X1 U1075 ( .A1(n1171), .A2(n1168), .ZN(n1345) );
NAND3_X1 U1076 ( .A1(n1257), .A2(n1076), .A3(G210), .ZN(n1168) );
INV_X1 U1077 ( .A(G953), .ZN(n1076) );
INV_X1 U1078 ( .A(G237), .ZN(n1257) );
INV_X1 U1079 ( .A(G101), .ZN(n1171) );
endmodule


