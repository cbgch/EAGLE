//Key = 1010011111111100100011011011100110101011111011001110000101000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319;

XNOR2_X1 U726 ( .A(G107), .B(n1002), .ZN(G9) );
NAND4_X1 U727 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(G75) );
NOR3_X1 U728 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1006) );
NAND2_X1 U729 ( .A1(n1010), .A2(n1011), .ZN(n1005) );
NAND2_X1 U730 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND3_X1 U731 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NAND2_X1 U732 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NAND2_X1 U733 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
OR2_X1 U734 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U735 ( .A1(n1023), .A2(n1024), .ZN(n1017) );
NAND2_X1 U736 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U737 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
XNOR2_X1 U738 ( .A(n1029), .B(KEYINPUT24), .ZN(n1027) );
NAND3_X1 U739 ( .A1(n1023), .A2(n1030), .A3(n1019), .ZN(n1012) );
NAND2_X1 U740 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND3_X1 U741 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1032) );
OR2_X1 U742 ( .A1(n1036), .A2(n1014), .ZN(n1034) );
OR3_X1 U743 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1033) );
NAND2_X1 U744 ( .A1(n1040), .A2(n1014), .ZN(n1031) );
INV_X1 U745 ( .A(n1041), .ZN(n1010) );
NAND4_X1 U746 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1003) );
NOR3_X1 U747 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
XNOR2_X1 U748 ( .A(n1049), .B(n1050), .ZN(n1048) );
NOR2_X1 U749 ( .A1(KEYINPUT46), .A2(n1051), .ZN(n1050) );
NAND3_X1 U750 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1046) );
XNOR2_X1 U751 ( .A(n1055), .B(n1056), .ZN(n1054) );
OR3_X1 U752 ( .A1(G472), .A2(KEYINPUT52), .A3(n1057), .ZN(n1053) );
NAND2_X1 U753 ( .A1(n1058), .A2(n1057), .ZN(n1052) );
NAND2_X1 U754 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
INV_X1 U755 ( .A(KEYINPUT52), .ZN(n1060) );
XNOR2_X1 U756 ( .A(KEYINPUT5), .B(n1061), .ZN(n1059) );
NOR3_X1 U757 ( .A1(n1062), .A2(n1029), .A3(n1039), .ZN(n1044) );
INV_X1 U758 ( .A(n1063), .ZN(n1029) );
XNOR2_X1 U759 ( .A(n1064), .B(KEYINPUT2), .ZN(n1062) );
NAND2_X1 U760 ( .A1(KEYINPUT52), .A2(G472), .ZN(n1043) );
NAND3_X1 U761 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(G72) );
XOR2_X1 U762 ( .A(n1068), .B(KEYINPUT51), .Z(n1067) );
NAND2_X1 U763 ( .A1(G953), .A2(n1069), .ZN(n1068) );
NAND2_X1 U764 ( .A1(G900), .A2(n1070), .ZN(n1069) );
OR2_X1 U765 ( .A1(n1071), .A2(G227), .ZN(n1070) );
NAND2_X1 U766 ( .A1(n1072), .A2(n1004), .ZN(n1066) );
XOR2_X1 U767 ( .A(n1071), .B(n1007), .Z(n1072) );
NAND4_X1 U768 ( .A1(G227), .A2(n1071), .A3(G900), .A4(G953), .ZN(n1065) );
XNOR2_X1 U769 ( .A(n1073), .B(n1074), .ZN(n1071) );
XOR2_X1 U770 ( .A(n1075), .B(n1076), .Z(n1074) );
XNOR2_X1 U771 ( .A(n1077), .B(n1078), .ZN(n1073) );
NAND2_X1 U772 ( .A1(n1079), .A2(KEYINPUT31), .ZN(n1078) );
XNOR2_X1 U773 ( .A(G125), .B(KEYINPUT4), .ZN(n1079) );
NAND2_X1 U774 ( .A1(n1080), .A2(KEYINPUT27), .ZN(n1077) );
XNOR2_X1 U775 ( .A(G134), .B(n1081), .ZN(n1080) );
XNOR2_X1 U776 ( .A(KEYINPUT48), .B(n1082), .ZN(n1081) );
XOR2_X1 U777 ( .A(n1083), .B(n1084), .Z(G69) );
NOR2_X1 U778 ( .A1(n1085), .A2(n1004), .ZN(n1084) );
NOR2_X1 U779 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR4_X1 U780 ( .A1(n1088), .A2(n1089), .A3(KEYINPUT17), .A4(n1090), .ZN(n1083) );
AND2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR2_X1 U782 ( .A1(n1093), .A2(n1094), .ZN(n1089) );
NOR2_X1 U783 ( .A1(KEYINPUT1), .A2(n1092), .ZN(n1094) );
INV_X1 U784 ( .A(n1095), .ZN(n1093) );
NOR4_X1 U785 ( .A1(n1095), .A2(n1091), .A3(KEYINPUT1), .A4(n1092), .ZN(n1088) );
NAND3_X1 U786 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1092) );
XOR2_X1 U787 ( .A(KEYINPUT44), .B(n1099), .Z(n1098) );
NOR2_X1 U788 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U789 ( .A1(n1101), .A2(n1100), .ZN(n1097) );
NAND2_X1 U790 ( .A1(G953), .A2(n1087), .ZN(n1096) );
INV_X1 U791 ( .A(KEYINPUT50), .ZN(n1091) );
NAND2_X1 U792 ( .A1(n1102), .A2(n1103), .ZN(n1095) );
NAND2_X1 U793 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XNOR2_X1 U794 ( .A(KEYINPUT14), .B(n1009), .ZN(n1105) );
INV_X1 U795 ( .A(n1008), .ZN(n1104) );
XNOR2_X1 U796 ( .A(KEYINPUT6), .B(n1004), .ZN(n1102) );
NOR2_X1 U797 ( .A1(n1106), .A2(n1107), .ZN(G66) );
XOR2_X1 U798 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U799 ( .A1(KEYINPUT54), .A2(n1110), .ZN(n1109) );
NOR2_X1 U800 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
NOR2_X1 U801 ( .A1(n1106), .A2(n1113), .ZN(G63) );
XOR2_X1 U802 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U803 ( .A(KEYINPUT32), .B(n1116), .Z(n1115) );
NOR2_X1 U804 ( .A1(n1056), .A2(n1112), .ZN(n1116) );
NOR2_X1 U805 ( .A1(n1106), .A2(n1117), .ZN(G60) );
XOR2_X1 U806 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U807 ( .A1(n1120), .A2(n1112), .ZN(n1118) );
XNOR2_X1 U808 ( .A(G104), .B(n1121), .ZN(G6) );
NOR2_X1 U809 ( .A1(n1106), .A2(n1122), .ZN(G57) );
XNOR2_X1 U810 ( .A(n1123), .B(n1124), .ZN(n1122) );
XOR2_X1 U811 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U812 ( .A1(n1061), .A2(n1112), .ZN(n1126) );
NOR2_X1 U813 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
XOR2_X1 U814 ( .A(n1129), .B(KEYINPUT39), .Z(n1128) );
NAND2_X1 U815 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U816 ( .A1(n1131), .A2(n1130), .ZN(n1127) );
XNOR2_X1 U817 ( .A(KEYINPUT8), .B(n1132), .ZN(n1130) );
NOR2_X1 U818 ( .A1(n1106), .A2(n1133), .ZN(G54) );
XOR2_X1 U819 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U820 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U821 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U822 ( .A1(KEYINPUT49), .A2(n1140), .ZN(n1138) );
XNOR2_X1 U823 ( .A(n1141), .B(n1142), .ZN(n1140) );
XOR2_X1 U824 ( .A(n1143), .B(n1144), .Z(n1134) );
XNOR2_X1 U825 ( .A(n1145), .B(G131), .ZN(n1144) );
XNOR2_X1 U826 ( .A(G110), .B(n1146), .ZN(n1143) );
NOR2_X1 U827 ( .A1(n1051), .A2(n1112), .ZN(n1146) );
NOR2_X1 U828 ( .A1(n1106), .A2(n1147), .ZN(G51) );
XOR2_X1 U829 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U830 ( .A(KEYINPUT18), .B(n1150), .Z(n1149) );
NOR2_X1 U831 ( .A1(n1151), .A2(n1112), .ZN(n1150) );
NAND2_X1 U832 ( .A1(G902), .A2(n1152), .ZN(n1112) );
OR3_X1 U833 ( .A1(n1009), .A2(n1008), .A3(n1007), .ZN(n1152) );
NAND4_X1 U834 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1007) );
AND4_X1 U835 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1156) );
AND2_X1 U836 ( .A1(n1161), .A2(n1162), .ZN(n1155) );
NAND2_X1 U837 ( .A1(n1163), .A2(n1019), .ZN(n1153) );
NAND4_X1 U838 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1008) );
NAND4_X1 U839 ( .A1(n1016), .A2(n1021), .A3(n1168), .A4(n1037), .ZN(n1165) );
NOR2_X1 U840 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
XNOR2_X1 U841 ( .A(n1171), .B(KEYINPUT15), .ZN(n1170) );
INV_X1 U842 ( .A(n1172), .ZN(n1169) );
NOR2_X1 U843 ( .A1(n1173), .A2(n1174), .ZN(n1164) );
AND4_X1 U844 ( .A1(KEYINPUT60), .A2(n1175), .A3(n1176), .A4(n1023), .ZN(n1174) );
NAND2_X1 U845 ( .A1(n1064), .A2(n1177), .ZN(n1176) );
NOR3_X1 U846 ( .A1(KEYINPUT60), .A2(n1025), .A3(n1178), .ZN(n1173) );
NAND4_X1 U847 ( .A1(n1179), .A2(n1180), .A3(n1121), .A4(n1002), .ZN(n1009) );
NAND2_X1 U848 ( .A1(n1037), .A2(n1181), .ZN(n1002) );
NAND2_X1 U849 ( .A1(n1038), .A2(n1181), .ZN(n1121) );
AND4_X1 U850 ( .A1(n1182), .A2(n1023), .A3(n1171), .A4(n1172), .ZN(n1181) );
NAND3_X1 U851 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1180) );
NAND2_X1 U852 ( .A1(n1171), .A2(n1186), .ZN(n1184) );
NAND2_X1 U853 ( .A1(n1187), .A2(n1025), .ZN(n1183) );
NAND2_X1 U854 ( .A1(KEYINPUT62), .A2(n1022), .ZN(n1187) );
NAND2_X1 U855 ( .A1(n1188), .A2(n1189), .ZN(n1179) );
INV_X1 U856 ( .A(KEYINPUT62), .ZN(n1189) );
AND2_X1 U857 ( .A1(G953), .A2(n1190), .ZN(n1106) );
XOR2_X1 U858 ( .A(KEYINPUT57), .B(G952), .Z(n1190) );
XNOR2_X1 U859 ( .A(G146), .B(n1159), .ZN(G48) );
NAND4_X1 U860 ( .A1(n1191), .A2(n1038), .A3(n1171), .A4(n1040), .ZN(n1159) );
XOR2_X1 U861 ( .A(n1154), .B(n1192), .Z(G45) );
NAND2_X1 U862 ( .A1(KEYINPUT9), .A2(G143), .ZN(n1192) );
NAND4_X1 U863 ( .A1(n1193), .A2(n1171), .A3(n1177), .A4(n1064), .ZN(n1154) );
XNOR2_X1 U864 ( .A(G140), .B(n1194), .ZN(G42) );
NAND2_X1 U865 ( .A1(n1195), .A2(n1019), .ZN(n1194) );
XNOR2_X1 U866 ( .A(n1163), .B(KEYINPUT23), .ZN(n1195) );
AND2_X1 U867 ( .A1(n1196), .A2(n1040), .ZN(n1163) );
XNOR2_X1 U868 ( .A(n1158), .B(n1197), .ZN(G39) );
NOR2_X1 U869 ( .A1(KEYINPUT53), .A2(n1082), .ZN(n1197) );
NAND4_X1 U870 ( .A1(n1191), .A2(n1019), .A3(n1040), .A4(n1014), .ZN(n1158) );
XOR2_X1 U871 ( .A(n1157), .B(n1198), .Z(G36) );
XNOR2_X1 U872 ( .A(G134), .B(KEYINPUT37), .ZN(n1198) );
NAND3_X1 U873 ( .A1(n1193), .A2(n1037), .A3(n1019), .ZN(n1157) );
XNOR2_X1 U874 ( .A(G131), .B(n1162), .ZN(G33) );
NAND3_X1 U875 ( .A1(n1019), .A2(n1193), .A3(n1038), .ZN(n1162) );
AND3_X1 U876 ( .A1(n1040), .A2(n1199), .A3(n1021), .ZN(n1193) );
XOR2_X1 U877 ( .A(n1182), .B(KEYINPUT47), .Z(n1040) );
AND2_X1 U878 ( .A1(n1028), .A2(n1200), .ZN(n1019) );
INV_X1 U879 ( .A(n1047), .ZN(n1028) );
XNOR2_X1 U880 ( .A(G128), .B(n1161), .ZN(G30) );
NAND4_X1 U881 ( .A1(n1191), .A2(n1037), .A3(n1182), .A4(n1171), .ZN(n1161) );
INV_X1 U882 ( .A(n1201), .ZN(n1037) );
AND3_X1 U883 ( .A1(n1202), .A2(n1199), .A3(n1203), .ZN(n1191) );
XNOR2_X1 U884 ( .A(G101), .B(n1204), .ZN(G3) );
NOR2_X1 U885 ( .A1(KEYINPUT58), .A2(n1205), .ZN(n1204) );
NOR3_X1 U886 ( .A1(n1206), .A2(n1186), .A3(n1207), .ZN(n1205) );
XNOR2_X1 U887 ( .A(KEYINPUT21), .B(n1025), .ZN(n1206) );
XNOR2_X1 U888 ( .A(G125), .B(n1160), .ZN(G27) );
NAND3_X1 U889 ( .A1(n1196), .A2(n1171), .A3(n1016), .ZN(n1160) );
AND3_X1 U890 ( .A1(n1038), .A2(n1199), .A3(n1022), .ZN(n1196) );
NAND2_X1 U891 ( .A1(n1041), .A2(n1208), .ZN(n1199) );
NAND4_X1 U892 ( .A1(G953), .A2(G902), .A3(n1209), .A4(n1210), .ZN(n1208) );
INV_X1 U893 ( .A(G900), .ZN(n1210) );
XOR2_X1 U894 ( .A(G122), .B(n1211), .Z(G24) );
NOR2_X1 U895 ( .A1(n1212), .A2(n1025), .ZN(n1211) );
XOR2_X1 U896 ( .A(n1178), .B(KEYINPUT59), .Z(n1212) );
NAND3_X1 U897 ( .A1(n1016), .A2(n1023), .A3(n1213), .ZN(n1178) );
AND3_X1 U898 ( .A1(n1177), .A2(n1172), .A3(n1064), .ZN(n1213) );
NOR2_X1 U899 ( .A1(n1202), .A2(n1203), .ZN(n1023) );
XNOR2_X1 U900 ( .A(G119), .B(n1214), .ZN(G21) );
NAND2_X1 U901 ( .A1(KEYINPUT34), .A2(n1215), .ZN(n1214) );
INV_X1 U902 ( .A(n1166), .ZN(n1215) );
NAND4_X1 U903 ( .A1(n1175), .A2(n1014), .A3(n1203), .A4(n1202), .ZN(n1166) );
XNOR2_X1 U904 ( .A(n1216), .B(n1217), .ZN(G18) );
NOR4_X1 U905 ( .A1(KEYINPUT3), .A2(n1201), .A3(n1186), .A4(n1218), .ZN(n1217) );
NAND2_X1 U906 ( .A1(n1219), .A2(n1177), .ZN(n1201) );
XNOR2_X1 U907 ( .A(n1064), .B(KEYINPUT25), .ZN(n1219) );
XNOR2_X1 U908 ( .A(G113), .B(n1167), .ZN(G15) );
NAND3_X1 U909 ( .A1(n1038), .A2(n1021), .A3(n1175), .ZN(n1167) );
INV_X1 U910 ( .A(n1218), .ZN(n1175) );
NAND3_X1 U911 ( .A1(n1171), .A2(n1172), .A3(n1016), .ZN(n1218) );
AND2_X1 U912 ( .A1(n1035), .A2(n1036), .ZN(n1016) );
INV_X1 U913 ( .A(n1186), .ZN(n1021) );
NAND2_X1 U914 ( .A1(n1042), .A2(n1202), .ZN(n1186) );
XOR2_X1 U915 ( .A(G110), .B(n1188), .Z(G12) );
AND3_X1 U916 ( .A1(n1022), .A2(n1171), .A3(n1185), .ZN(n1188) );
INV_X1 U917 ( .A(n1207), .ZN(n1185) );
NAND3_X1 U918 ( .A1(n1014), .A2(n1172), .A3(n1182), .ZN(n1207) );
NOR2_X1 U919 ( .A1(n1035), .A2(n1039), .ZN(n1182) );
INV_X1 U920 ( .A(n1036), .ZN(n1039) );
NAND2_X1 U921 ( .A1(G221), .A2(n1220), .ZN(n1036) );
XNOR2_X1 U922 ( .A(n1049), .B(n1051), .ZN(n1035) );
INV_X1 U923 ( .A(G469), .ZN(n1051) );
NAND2_X1 U924 ( .A1(n1221), .A2(n1222), .ZN(n1049) );
XOR2_X1 U925 ( .A(n1223), .B(n1224), .Z(n1221) );
XNOR2_X1 U926 ( .A(n1136), .B(n1142), .ZN(n1224) );
XOR2_X1 U927 ( .A(n1225), .B(n1226), .Z(n1142) );
XNOR2_X1 U928 ( .A(n1227), .B(G101), .ZN(n1226) );
NAND3_X1 U929 ( .A1(n1228), .A2(n1229), .A3(KEYINPUT45), .ZN(n1225) );
NAND2_X1 U930 ( .A1(G104), .A2(n1230), .ZN(n1229) );
NAND2_X1 U931 ( .A1(G107), .A2(n1231), .ZN(n1230) );
OR2_X1 U932 ( .A1(n1232), .A2(KEYINPUT36), .ZN(n1231) );
NAND3_X1 U933 ( .A1(n1233), .A2(n1234), .A3(KEYINPUT36), .ZN(n1228) );
NAND2_X1 U934 ( .A1(G107), .A2(n1232), .ZN(n1234) );
INV_X1 U935 ( .A(KEYINPUT26), .ZN(n1232) );
NAND2_X1 U936 ( .A1(KEYINPUT26), .A2(n1235), .ZN(n1233) );
NAND2_X1 U937 ( .A1(G107), .A2(n1236), .ZN(n1235) );
XNOR2_X1 U938 ( .A(n1237), .B(KEYINPUT61), .ZN(n1136) );
NAND2_X1 U939 ( .A1(G227), .A2(n1004), .ZN(n1237) );
XNOR2_X1 U940 ( .A(n1238), .B(n1239), .ZN(n1223) );
INV_X1 U941 ( .A(n1240), .ZN(n1239) );
NAND3_X1 U942 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1238) );
NAND2_X1 U943 ( .A1(KEYINPUT33), .A2(n1244), .ZN(n1243) );
NAND3_X1 U944 ( .A1(n1245), .A2(n1246), .A3(G140), .ZN(n1242) );
NAND2_X1 U945 ( .A1(n1247), .A2(n1145), .ZN(n1241) );
NAND2_X1 U946 ( .A1(n1248), .A2(n1246), .ZN(n1247) );
INV_X1 U947 ( .A(KEYINPUT33), .ZN(n1246) );
XNOR2_X1 U948 ( .A(KEYINPUT30), .B(n1244), .ZN(n1248) );
INV_X1 U949 ( .A(n1245), .ZN(n1244) );
XOR2_X1 U950 ( .A(G110), .B(KEYINPUT41), .Z(n1245) );
NAND2_X1 U951 ( .A1(n1041), .A2(n1249), .ZN(n1172) );
NAND4_X1 U952 ( .A1(G953), .A2(G902), .A3(n1209), .A4(n1087), .ZN(n1249) );
INV_X1 U953 ( .A(G898), .ZN(n1087) );
NAND3_X1 U954 ( .A1(n1209), .A2(n1004), .A3(G952), .ZN(n1041) );
NAND2_X1 U955 ( .A1(G237), .A2(G234), .ZN(n1209) );
NAND2_X1 U956 ( .A1(n1250), .A2(n1251), .ZN(n1014) );
OR3_X1 U957 ( .A1(n1177), .A2(n1064), .A3(KEYINPUT25), .ZN(n1251) );
NAND2_X1 U958 ( .A1(KEYINPUT25), .A2(n1038), .ZN(n1250) );
NOR2_X1 U959 ( .A1(n1252), .A2(n1177), .ZN(n1038) );
XNOR2_X1 U960 ( .A(n1253), .B(n1055), .ZN(n1177) );
NAND2_X1 U961 ( .A1(n1114), .A2(n1222), .ZN(n1055) );
XNOR2_X1 U962 ( .A(n1254), .B(n1255), .ZN(n1114) );
XOR2_X1 U963 ( .A(G107), .B(n1256), .Z(n1255) );
XNOR2_X1 U964 ( .A(G122), .B(n1216), .ZN(n1256) );
XOR2_X1 U965 ( .A(n1257), .B(n1258), .Z(n1254) );
AND2_X1 U966 ( .A1(n1259), .A2(G217), .ZN(n1258) );
NAND2_X1 U967 ( .A1(n1260), .A2(n1261), .ZN(n1257) );
NAND2_X1 U968 ( .A1(G134), .A2(n1262), .ZN(n1261) );
XOR2_X1 U969 ( .A(KEYINPUT10), .B(n1263), .Z(n1260) );
NOR2_X1 U970 ( .A1(G134), .A2(n1262), .ZN(n1263) );
NAND2_X1 U971 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
NAND2_X1 U972 ( .A1(G143), .A2(n1227), .ZN(n1265) );
XOR2_X1 U973 ( .A(KEYINPUT16), .B(n1266), .Z(n1264) );
NOR2_X1 U974 ( .A1(G143), .A2(n1227), .ZN(n1266) );
NAND2_X1 U975 ( .A1(KEYINPUT28), .A2(n1056), .ZN(n1253) );
INV_X1 U976 ( .A(G478), .ZN(n1056) );
INV_X1 U977 ( .A(n1064), .ZN(n1252) );
XOR2_X1 U978 ( .A(n1267), .B(n1120), .Z(n1064) );
INV_X1 U979 ( .A(G475), .ZN(n1120) );
OR2_X1 U980 ( .A1(n1119), .A2(G902), .ZN(n1267) );
XOR2_X1 U981 ( .A(n1268), .B(n1269), .Z(n1119) );
XOR2_X1 U982 ( .A(G122), .B(n1270), .Z(n1269) );
NOR2_X1 U983 ( .A1(KEYINPUT63), .A2(n1271), .ZN(n1270) );
XOR2_X1 U984 ( .A(n1076), .B(n1272), .Z(n1271) );
XOR2_X1 U985 ( .A(n1273), .B(n1274), .Z(n1272) );
NAND2_X1 U986 ( .A1(G214), .A2(n1275), .ZN(n1274) );
NAND2_X1 U987 ( .A1(KEYINPUT55), .A2(n1276), .ZN(n1273) );
XNOR2_X1 U988 ( .A(n1145), .B(G125), .ZN(n1276) );
INV_X1 U989 ( .A(G140), .ZN(n1145) );
INV_X1 U990 ( .A(n1025), .ZN(n1171) );
NAND2_X1 U991 ( .A1(n1047), .A2(n1200), .ZN(n1025) );
XNOR2_X1 U992 ( .A(n1063), .B(KEYINPUT0), .ZN(n1200) );
NAND2_X1 U993 ( .A1(G214), .A2(n1277), .ZN(n1063) );
XNOR2_X1 U994 ( .A(n1151), .B(n1278), .ZN(n1047) );
NOR2_X1 U995 ( .A1(G902), .A2(n1148), .ZN(n1278) );
XNOR2_X1 U996 ( .A(n1279), .B(n1280), .ZN(n1148) );
XNOR2_X1 U997 ( .A(n1141), .B(n1281), .ZN(n1280) );
XNOR2_X1 U998 ( .A(n1101), .B(n1282), .ZN(n1281) );
NOR2_X1 U999 ( .A1(G953), .A2(n1086), .ZN(n1282) );
INV_X1 U1000 ( .A(G224), .ZN(n1086) );
XOR2_X1 U1001 ( .A(G110), .B(n1283), .Z(n1101) );
XOR2_X1 U1002 ( .A(KEYINPUT20), .B(G122), .Z(n1283) );
XOR2_X1 U1003 ( .A(n1284), .B(n1285), .Z(n1279) );
NOR2_X1 U1004 ( .A1(KEYINPUT43), .A2(n1100), .ZN(n1285) );
XNOR2_X1 U1005 ( .A(n1286), .B(n1287), .ZN(n1100) );
XOR2_X1 U1006 ( .A(n1288), .B(n1268), .Z(n1287) );
XNOR2_X1 U1007 ( .A(G113), .B(n1236), .ZN(n1268) );
INV_X1 U1008 ( .A(G104), .ZN(n1236) );
NOR2_X1 U1009 ( .A1(KEYINPUT35), .A2(n1216), .ZN(n1288) );
XNOR2_X1 U1010 ( .A(G101), .B(n1289), .ZN(n1286) );
XNOR2_X1 U1011 ( .A(n1290), .B(G107), .ZN(n1289) );
XNOR2_X1 U1012 ( .A(G125), .B(n1291), .ZN(n1284) );
NAND2_X1 U1013 ( .A1(G210), .A2(n1277), .ZN(n1151) );
NAND2_X1 U1014 ( .A1(n1292), .A2(n1222), .ZN(n1277) );
INV_X1 U1015 ( .A(G237), .ZN(n1292) );
NOR2_X1 U1016 ( .A1(n1202), .A2(n1042), .ZN(n1022) );
INV_X1 U1017 ( .A(n1203), .ZN(n1042) );
XOR2_X1 U1018 ( .A(n1293), .B(n1111), .Z(n1203) );
NAND2_X1 U1019 ( .A1(G217), .A2(n1220), .ZN(n1111) );
NAND2_X1 U1020 ( .A1(G234), .A2(n1222), .ZN(n1220) );
NAND2_X1 U1021 ( .A1(n1110), .A2(n1222), .ZN(n1293) );
XNOR2_X1 U1022 ( .A(n1294), .B(n1295), .ZN(n1110) );
XOR2_X1 U1023 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U1024 ( .A(n1298), .B(n1075), .Z(n1297) );
XNOR2_X1 U1025 ( .A(n1227), .B(G140), .ZN(n1075) );
INV_X1 U1026 ( .A(G128), .ZN(n1227) );
NAND2_X1 U1027 ( .A1(KEYINPUT42), .A2(G146), .ZN(n1298) );
XOR2_X1 U1028 ( .A(n1299), .B(n1300), .Z(n1296) );
NOR2_X1 U1029 ( .A1(G137), .A2(KEYINPUT19), .ZN(n1300) );
NAND2_X1 U1030 ( .A1(G221), .A2(n1259), .ZN(n1299) );
AND2_X1 U1031 ( .A1(G234), .A2(n1004), .ZN(n1259) );
INV_X1 U1032 ( .A(G953), .ZN(n1004) );
XOR2_X1 U1033 ( .A(n1301), .B(n1302), .Z(n1294) );
XOR2_X1 U1034 ( .A(KEYINPUT38), .B(G125), .Z(n1302) );
XNOR2_X1 U1035 ( .A(G110), .B(G119), .ZN(n1301) );
XOR2_X1 U1036 ( .A(n1057), .B(n1061), .Z(n1202) );
INV_X1 U1037 ( .A(G472), .ZN(n1061) );
NAND3_X1 U1038 ( .A1(n1303), .A2(n1304), .A3(n1222), .ZN(n1057) );
INV_X1 U1039 ( .A(G902), .ZN(n1222) );
NAND2_X1 U1040 ( .A1(KEYINPUT11), .A2(n1305), .ZN(n1304) );
XOR2_X1 U1041 ( .A(n1123), .B(n1306), .Z(n1305) );
OR3_X1 U1042 ( .A1(n1123), .A2(n1306), .A3(KEYINPUT11), .ZN(n1303) );
XOR2_X1 U1043 ( .A(n1307), .B(n1131), .Z(n1306) );
INV_X1 U1044 ( .A(G101), .ZN(n1131) );
NAND2_X1 U1045 ( .A1(KEYINPUT12), .A2(n1132), .ZN(n1307) );
NAND2_X1 U1046 ( .A1(G210), .A2(n1275), .ZN(n1132) );
NOR2_X1 U1047 ( .A1(G953), .A2(G237), .ZN(n1275) );
XOR2_X1 U1048 ( .A(n1308), .B(n1309), .Z(n1123) );
XNOR2_X1 U1049 ( .A(G113), .B(n1310), .ZN(n1309) );
NAND2_X1 U1050 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NAND4_X1 U1051 ( .A1(KEYINPUT13), .A2(n1216), .A3(n1290), .A4(n1313), .ZN(n1312) );
NAND2_X1 U1052 ( .A1(n1314), .A2(n1315), .ZN(n1311) );
NAND2_X1 U1053 ( .A1(n1316), .A2(n1290), .ZN(n1315) );
INV_X1 U1054 ( .A(G119), .ZN(n1290) );
OR2_X1 U1055 ( .A1(n1216), .A2(KEYINPUT13), .ZN(n1316) );
NAND2_X1 U1056 ( .A1(n1216), .A2(n1313), .ZN(n1314) );
INV_X1 U1057 ( .A(KEYINPUT22), .ZN(n1313) );
INV_X1 U1058 ( .A(G116), .ZN(n1216) );
XNOR2_X1 U1059 ( .A(n1240), .B(n1291), .ZN(n1308) );
NOR2_X1 U1060 ( .A1(KEYINPUT29), .A2(G128), .ZN(n1291) );
XNOR2_X1 U1061 ( .A(n1139), .B(n1076), .ZN(n1240) );
XOR2_X1 U1062 ( .A(G131), .B(n1141), .Z(n1076) );
XOR2_X1 U1063 ( .A(G146), .B(G143), .Z(n1141) );
XOR2_X1 U1064 ( .A(n1317), .B(n1318), .Z(n1139) );
XNOR2_X1 U1065 ( .A(KEYINPUT56), .B(n1082), .ZN(n1318) );
INV_X1 U1066 ( .A(G137), .ZN(n1082) );
NAND2_X1 U1067 ( .A1(n1319), .A2(KEYINPUT7), .ZN(n1317) );
XNOR2_X1 U1068 ( .A(G134), .B(KEYINPUT40), .ZN(n1319) );
endmodule


