//Key = 0101000000000101111001010011101011100110010110111010011110000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349;

XNOR2_X1 U749 ( .A(G107), .B(n1034), .ZN(G9) );
NOR2_X1 U750 ( .A1(n1035), .A2(n1036), .ZN(G75) );
NOR4_X1 U751 ( .A1(G953), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1036) );
NOR2_X1 U752 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U753 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR3_X1 U754 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NAND3_X1 U755 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1044) );
NAND2_X1 U756 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
OR3_X1 U757 ( .A1(n1052), .A2(n1053), .A3(n1050), .ZN(n1047) );
NOR4_X1 U758 ( .A1(n1054), .A2(n1055), .A3(n1050), .A4(n1051), .ZN(n1042) );
NOR4_X1 U759 ( .A1(n1046), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1055) );
NOR2_X1 U760 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR2_X1 U761 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR3_X1 U762 ( .A1(n1063), .A2(n1064), .A3(n1045), .ZN(n1057) );
NOR2_X1 U763 ( .A1(n1065), .A2(n1066), .ZN(n1056) );
XOR2_X1 U764 ( .A(KEYINPUT33), .B(n1067), .Z(n1066) );
NOR2_X1 U765 ( .A1(n1068), .A2(n1069), .ZN(n1054) );
NOR2_X1 U766 ( .A1(n1045), .A2(n1060), .ZN(n1069) );
NOR3_X1 U767 ( .A1(n1037), .A2(G953), .A3(G952), .ZN(n1035) );
AND4_X1 U768 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1037) );
NOR4_X1 U769 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1050), .ZN(n1073) );
INV_X1 U770 ( .A(n1077), .ZN(n1050) );
NOR2_X1 U771 ( .A1(n1078), .A2(n1079), .ZN(n1072) );
XOR2_X1 U772 ( .A(n1080), .B(n1081), .Z(n1078) );
NAND2_X1 U773 ( .A1(KEYINPUT48), .A2(n1082), .ZN(n1080) );
XOR2_X1 U774 ( .A(n1083), .B(G469), .Z(n1070) );
XOR2_X1 U775 ( .A(n1084), .B(n1085), .Z(G72) );
NAND2_X1 U776 ( .A1(G953), .A2(n1086), .ZN(n1085) );
NAND2_X1 U777 ( .A1(G900), .A2(G227), .ZN(n1086) );
NAND2_X1 U778 ( .A1(KEYINPUT23), .A2(n1087), .ZN(n1084) );
XOR2_X1 U779 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U780 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U781 ( .A(n1092), .B(n1093), .Z(n1091) );
XOR2_X1 U782 ( .A(G131), .B(n1094), .Z(n1093) );
XOR2_X1 U783 ( .A(KEYINPUT55), .B(G140), .Z(n1094) );
XOR2_X1 U784 ( .A(n1095), .B(n1096), .Z(n1092) );
XOR2_X1 U785 ( .A(G125), .B(n1097), .Z(n1096) );
NOR2_X1 U786 ( .A1(KEYINPUT9), .A2(n1098), .ZN(n1097) );
XNOR2_X1 U787 ( .A(G134), .B(n1099), .ZN(n1098) );
NOR2_X1 U788 ( .A1(KEYINPUT5), .A2(n1100), .ZN(n1099) );
NAND2_X1 U789 ( .A1(n1101), .A2(KEYINPUT53), .ZN(n1095) );
XOR2_X1 U790 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR3_X1 U791 ( .A1(n1104), .A2(KEYINPUT49), .A3(G953), .ZN(n1088) );
XOR2_X1 U792 ( .A(KEYINPUT40), .B(n1105), .Z(n1104) );
NOR2_X1 U793 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U794 ( .A(n1108), .B(n1109), .Z(G69) );
NOR2_X1 U795 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U796 ( .A(n1112), .B(KEYINPUT51), .Z(n1111) );
AND2_X1 U797 ( .A1(G224), .A2(G898), .ZN(n1110) );
NAND2_X1 U798 ( .A1(n1113), .A2(n1114), .ZN(n1108) );
NAND3_X1 U799 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
INV_X1 U800 ( .A(n1118), .ZN(n1116) );
OR2_X1 U801 ( .A1(n1115), .A2(n1117), .ZN(n1113) );
NAND2_X1 U802 ( .A1(n1112), .A2(n1119), .ZN(n1117) );
NAND4_X1 U803 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1119) );
NOR2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XNOR2_X1 U805 ( .A(n1126), .B(KEYINPUT6), .ZN(n1125) );
XOR2_X1 U806 ( .A(n1127), .B(KEYINPUT50), .Z(n1124) );
XOR2_X1 U807 ( .A(n1128), .B(n1129), .Z(n1115) );
XNOR2_X1 U808 ( .A(n1130), .B(KEYINPUT42), .ZN(n1129) );
NAND2_X1 U809 ( .A1(KEYINPUT54), .A2(n1131), .ZN(n1130) );
XNOR2_X1 U810 ( .A(n1132), .B(n1133), .ZN(n1128) );
NOR2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(G66) );
XOR2_X1 U812 ( .A(n1136), .B(n1137), .Z(n1135) );
NOR2_X1 U813 ( .A1(KEYINPUT0), .A2(n1138), .ZN(n1137) );
NAND2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1134), .A2(n1141), .ZN(G63) );
XOR2_X1 U816 ( .A(n1142), .B(n1143), .Z(n1141) );
AND2_X1 U817 ( .A1(G478), .A2(n1139), .ZN(n1142) );
NOR2_X1 U818 ( .A1(n1134), .A2(n1144), .ZN(G60) );
NOR2_X1 U819 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U820 ( .A(KEYINPUT14), .B(n1147), .Z(n1146) );
NOR2_X1 U821 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
AND2_X1 U822 ( .A1(n1149), .A2(n1148), .ZN(n1145) );
NAND2_X1 U823 ( .A1(n1139), .A2(G475), .ZN(n1149) );
XNOR2_X1 U824 ( .A(G104), .B(n1150), .ZN(G6) );
NOR2_X1 U825 ( .A1(n1134), .A2(n1151), .ZN(G57) );
XOR2_X1 U826 ( .A(n1152), .B(KEYINPUT38), .Z(n1151) );
NAND2_X1 U827 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND2_X1 U828 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U829 ( .A(KEYINPUT8), .B(n1157), .Z(n1155) );
NAND2_X1 U830 ( .A1(n1158), .A2(n1159), .ZN(n1153) );
XOR2_X1 U831 ( .A(KEYINPUT56), .B(n1157), .Z(n1158) );
AND2_X1 U832 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NAND2_X1 U833 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U834 ( .A1(n1139), .A2(G472), .ZN(n1163) );
INV_X1 U835 ( .A(n1164), .ZN(n1162) );
NAND3_X1 U836 ( .A1(n1139), .A2(G472), .A3(n1164), .ZN(n1160) );
XOR2_X1 U837 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U838 ( .A(KEYINPUT21), .B(n1167), .Z(n1166) );
NOR2_X1 U839 ( .A1(n1134), .A2(n1168), .ZN(G54) );
NOR3_X1 U840 ( .A1(n1169), .A2(n1170), .A3(n1171), .ZN(n1168) );
NOR2_X1 U841 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XOR2_X1 U842 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR3_X1 U843 ( .A1(n1176), .A2(n1177), .A3(n1175), .ZN(n1170) );
INV_X1 U844 ( .A(n1172), .ZN(n1176) );
AND2_X1 U845 ( .A1(n1175), .A2(n1178), .ZN(n1169) );
XNOR2_X1 U846 ( .A(n1179), .B(n1180), .ZN(n1175) );
NOR3_X1 U847 ( .A1(n1181), .A2(KEYINPUT57), .A3(G953), .ZN(n1180) );
INV_X1 U848 ( .A(G227), .ZN(n1181) );
NAND2_X1 U849 ( .A1(n1139), .A2(G469), .ZN(n1179) );
INV_X1 U850 ( .A(n1182), .ZN(n1139) );
NOR2_X1 U851 ( .A1(n1183), .A2(n1184), .ZN(G51) );
XOR2_X1 U852 ( .A(KEYINPUT61), .B(n1134), .Z(n1184) );
NOR2_X1 U853 ( .A1(n1112), .A2(G952), .ZN(n1134) );
XOR2_X1 U854 ( .A(n1185), .B(n1186), .Z(n1183) );
OR2_X1 U855 ( .A1(n1182), .A2(n1082), .ZN(n1186) );
NAND2_X1 U856 ( .A1(G902), .A2(n1039), .ZN(n1182) );
NAND4_X1 U857 ( .A1(n1187), .A2(n1188), .A3(n1126), .A4(n1189), .ZN(n1039) );
AND4_X1 U858 ( .A1(n1127), .A2(n1121), .A3(n1120), .A4(n1122), .ZN(n1189) );
AND4_X1 U859 ( .A1(n1150), .A2(n1190), .A3(n1191), .A4(n1034), .ZN(n1126) );
NAND3_X1 U860 ( .A1(n1053), .A2(n1067), .A3(n1192), .ZN(n1034) );
NAND3_X1 U861 ( .A1(n1192), .A2(n1067), .A3(n1052), .ZN(n1150) );
XNOR2_X1 U862 ( .A(KEYINPUT29), .B(n1106), .ZN(n1188) );
NAND3_X1 U863 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1106) );
NAND2_X1 U864 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
XOR2_X1 U865 ( .A(KEYINPUT62), .B(n1198), .Z(n1197) );
NAND3_X1 U866 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1193) );
NAND2_X1 U867 ( .A1(n1202), .A2(n1203), .ZN(n1200) );
NAND2_X1 U868 ( .A1(n1204), .A2(n1071), .ZN(n1203) );
XOR2_X1 U869 ( .A(n1060), .B(KEYINPUT41), .Z(n1204) );
INV_X1 U870 ( .A(n1049), .ZN(n1060) );
INV_X1 U871 ( .A(n1107), .ZN(n1187) );
NAND4_X1 U872 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1107) );
NAND2_X1 U873 ( .A1(n1209), .A2(n1210), .ZN(n1206) );
INV_X1 U874 ( .A(n1202), .ZN(n1209) );
NAND3_X1 U875 ( .A1(n1062), .A2(n1053), .A3(n1211), .ZN(n1205) );
NAND2_X1 U876 ( .A1(KEYINPUT30), .A2(n1212), .ZN(n1185) );
XOR2_X1 U877 ( .A(n1213), .B(n1214), .Z(n1212) );
NOR2_X1 U878 ( .A1(KEYINPUT39), .A2(n1215), .ZN(n1213) );
XOR2_X1 U879 ( .A(n1102), .B(G125), .Z(n1215) );
XOR2_X1 U880 ( .A(n1216), .B(n1217), .Z(G48) );
NOR2_X1 U881 ( .A1(KEYINPUT20), .A2(n1218), .ZN(n1217) );
NOR4_X1 U882 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1202), .ZN(n1216) );
NAND2_X1 U883 ( .A1(n1052), .A2(n1196), .ZN(n1202) );
NOR2_X1 U884 ( .A1(KEYINPUT34), .A2(n1222), .ZN(n1220) );
NOR2_X1 U885 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
NOR2_X1 U886 ( .A1(n1201), .A2(n1225), .ZN(n1219) );
INV_X1 U887 ( .A(KEYINPUT34), .ZN(n1225) );
XNOR2_X1 U888 ( .A(G143), .B(n1226), .ZN(G45) );
NAND2_X1 U889 ( .A1(n1198), .A2(n1196), .ZN(n1226) );
AND4_X1 U890 ( .A1(n1201), .A2(n1062), .A3(n1227), .A4(n1228), .ZN(n1198) );
XOR2_X1 U891 ( .A(n1229), .B(n1194), .Z(G42) );
NAND3_X1 U892 ( .A1(n1052), .A2(n1061), .A3(n1211), .ZN(n1194) );
XOR2_X1 U893 ( .A(n1100), .B(n1230), .Z(G39) );
NAND2_X1 U894 ( .A1(n1211), .A2(n1231), .ZN(n1230) );
INV_X1 U895 ( .A(G137), .ZN(n1100) );
XNOR2_X1 U896 ( .A(G134), .B(n1232), .ZN(G36) );
NAND4_X1 U897 ( .A1(KEYINPUT15), .A2(n1211), .A3(n1062), .A4(n1053), .ZN(n1232) );
XNOR2_X1 U898 ( .A(G131), .B(n1207), .ZN(G33) );
NAND3_X1 U899 ( .A1(n1052), .A2(n1062), .A3(n1211), .ZN(n1207) );
AND2_X1 U900 ( .A1(n1049), .A2(n1201), .ZN(n1211) );
NOR2_X1 U901 ( .A1(n1064), .A2(n1076), .ZN(n1049) );
INV_X1 U902 ( .A(n1063), .ZN(n1076) );
NAND3_X1 U903 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(G30) );
NAND2_X1 U904 ( .A1(KEYINPUT52), .A2(G128), .ZN(n1235) );
OR3_X1 U905 ( .A1(G128), .A2(KEYINPUT52), .A3(n1208), .ZN(n1234) );
NAND2_X1 U906 ( .A1(n1236), .A2(n1208), .ZN(n1233) );
NAND4_X1 U907 ( .A1(n1201), .A2(n1199), .A3(n1053), .A4(n1196), .ZN(n1208) );
AND2_X1 U908 ( .A1(n1237), .A2(n1224), .ZN(n1201) );
NAND2_X1 U909 ( .A1(n1238), .A2(n1239), .ZN(n1236) );
INV_X1 U910 ( .A(KEYINPUT52), .ZN(n1239) );
XOR2_X1 U911 ( .A(KEYINPUT27), .B(G128), .Z(n1238) );
XOR2_X1 U912 ( .A(n1190), .B(n1240), .Z(G3) );
NOR2_X1 U913 ( .A1(G101), .A2(KEYINPUT45), .ZN(n1240) );
NAND3_X1 U914 ( .A1(n1071), .A2(n1192), .A3(n1062), .ZN(n1190) );
XNOR2_X1 U915 ( .A(G125), .B(n1241), .ZN(G27) );
NAND4_X1 U916 ( .A1(n1242), .A2(KEYINPUT3), .A3(n1210), .A4(n1052), .ZN(n1241) );
AND4_X1 U917 ( .A1(n1068), .A2(n1061), .A3(n1224), .A4(n1077), .ZN(n1210) );
NAND2_X1 U918 ( .A1(n1041), .A2(n1243), .ZN(n1224) );
NAND3_X1 U919 ( .A1(G902), .A2(n1244), .A3(n1090), .ZN(n1243) );
NOR2_X1 U920 ( .A1(n1112), .A2(G900), .ZN(n1090) );
XOR2_X1 U921 ( .A(n1065), .B(KEYINPUT13), .Z(n1242) );
XNOR2_X1 U922 ( .A(n1122), .B(n1245), .ZN(G24) );
NOR2_X1 U923 ( .A1(KEYINPUT11), .A2(n1246), .ZN(n1245) );
NAND4_X1 U924 ( .A1(n1247), .A2(n1067), .A3(n1227), .A4(n1228), .ZN(n1122) );
INV_X1 U925 ( .A(n1045), .ZN(n1067) );
NAND2_X1 U926 ( .A1(n1248), .A2(n1249), .ZN(n1045) );
XOR2_X1 U927 ( .A(n1250), .B(n1120), .Z(G21) );
NAND2_X1 U928 ( .A1(n1231), .A2(n1247), .ZN(n1120) );
NOR2_X1 U929 ( .A1(n1221), .A2(n1051), .ZN(n1231) );
INV_X1 U930 ( .A(n1071), .ZN(n1051) );
INV_X1 U931 ( .A(n1199), .ZN(n1221) );
NOR2_X1 U932 ( .A1(n1249), .A2(n1248), .ZN(n1199) );
XNOR2_X1 U933 ( .A(G116), .B(n1121), .ZN(G18) );
NAND3_X1 U934 ( .A1(n1062), .A2(n1053), .A3(n1247), .ZN(n1121) );
NOR2_X1 U935 ( .A1(n1227), .A2(n1251), .ZN(n1053) );
XOR2_X1 U936 ( .A(n1252), .B(n1127), .Z(G15) );
NAND3_X1 U937 ( .A1(n1052), .A2(n1062), .A3(n1247), .ZN(n1127) );
AND3_X1 U938 ( .A1(n1253), .A2(n1077), .A3(n1068), .ZN(n1247) );
INV_X1 U939 ( .A(n1046), .ZN(n1068) );
NOR2_X1 U940 ( .A1(n1079), .A2(n1248), .ZN(n1062) );
AND2_X1 U941 ( .A1(n1251), .A2(n1227), .ZN(n1052) );
XOR2_X1 U942 ( .A(G110), .B(n1254), .Z(G12) );
NOR2_X1 U943 ( .A1(KEYINPUT36), .A2(n1191), .ZN(n1254) );
NAND3_X1 U944 ( .A1(n1071), .A2(n1192), .A3(n1061), .ZN(n1191) );
AND2_X1 U945 ( .A1(n1248), .A2(n1079), .ZN(n1061) );
INV_X1 U946 ( .A(n1249), .ZN(n1079) );
XOR2_X1 U947 ( .A(n1255), .B(n1140), .Z(n1249) );
AND2_X1 U948 ( .A1(G217), .A2(n1256), .ZN(n1140) );
OR2_X1 U949 ( .A1(n1138), .A2(G902), .ZN(n1255) );
XOR2_X1 U950 ( .A(n1257), .B(n1258), .Z(n1138) );
XOR2_X1 U951 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U952 ( .A(G125), .B(G110), .Z(n1260) );
XOR2_X1 U953 ( .A(G146), .B(G137), .Z(n1259) );
XOR2_X1 U954 ( .A(n1261), .B(n1262), .Z(n1257) );
XOR2_X1 U955 ( .A(n1263), .B(n1264), .Z(n1262) );
NAND2_X1 U956 ( .A1(KEYINPUT37), .A2(n1229), .ZN(n1264) );
INV_X1 U957 ( .A(G140), .ZN(n1229) );
NAND2_X1 U958 ( .A1(KEYINPUT18), .A2(n1250), .ZN(n1263) );
INV_X1 U959 ( .A(G119), .ZN(n1250) );
XOR2_X1 U960 ( .A(n1265), .B(n1266), .Z(n1261) );
NAND2_X1 U961 ( .A1(n1267), .A2(G221), .ZN(n1265) );
NOR2_X1 U962 ( .A1(n1268), .A2(n1075), .ZN(n1248) );
NOR3_X1 U963 ( .A1(G472), .A2(G902), .A3(n1269), .ZN(n1075) );
INV_X1 U964 ( .A(n1270), .ZN(n1269) );
XOR2_X1 U965 ( .A(n1074), .B(KEYINPUT2), .Z(n1268) );
AND2_X1 U966 ( .A1(G472), .A2(n1271), .ZN(n1074) );
NAND2_X1 U967 ( .A1(n1272), .A2(n1270), .ZN(n1271) );
NAND2_X1 U968 ( .A1(n1273), .A2(n1274), .ZN(n1270) );
NAND2_X1 U969 ( .A1(n1275), .A2(n1159), .ZN(n1274) );
XOR2_X1 U970 ( .A(n1276), .B(KEYINPUT25), .Z(n1273) );
OR2_X1 U971 ( .A1(n1159), .A2(n1275), .ZN(n1276) );
XNOR2_X1 U972 ( .A(n1277), .B(n1167), .ZN(n1275) );
XNOR2_X1 U973 ( .A(n1278), .B(n1279), .ZN(n1167) );
XOR2_X1 U974 ( .A(G119), .B(n1280), .Z(n1279) );
NOR2_X1 U975 ( .A1(G116), .A2(KEYINPUT35), .ZN(n1280) );
NAND2_X1 U976 ( .A1(KEYINPUT46), .A2(n1252), .ZN(n1278) );
INV_X1 U977 ( .A(G113), .ZN(n1252) );
NAND2_X1 U978 ( .A1(KEYINPUT17), .A2(n1165), .ZN(n1277) );
INV_X1 U979 ( .A(n1156), .ZN(n1159) );
XOR2_X1 U980 ( .A(n1281), .B(G101), .Z(n1156) );
NAND2_X1 U981 ( .A1(n1282), .A2(G210), .ZN(n1281) );
AND2_X1 U982 ( .A1(n1253), .A2(n1237), .ZN(n1192) );
INV_X1 U983 ( .A(n1223), .ZN(n1237) );
NAND2_X1 U984 ( .A1(n1077), .A2(n1046), .ZN(n1223) );
NAND3_X1 U985 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1046) );
OR2_X1 U986 ( .A1(n1083), .A2(KEYINPUT43), .ZN(n1285) );
NAND3_X1 U987 ( .A1(KEYINPUT43), .A2(n1083), .A3(G469), .ZN(n1284) );
NAND2_X1 U988 ( .A1(n1286), .A2(n1287), .ZN(n1283) );
INV_X1 U989 ( .A(G469), .ZN(n1287) );
NAND2_X1 U990 ( .A1(KEYINPUT43), .A2(n1288), .ZN(n1286) );
XNOR2_X1 U991 ( .A(KEYINPUT32), .B(n1083), .ZN(n1288) );
NAND4_X1 U992 ( .A1(n1289), .A2(n1272), .A3(n1290), .A4(n1291), .ZN(n1083) );
NAND2_X1 U993 ( .A1(n1178), .A2(n1292), .ZN(n1291) );
INV_X1 U994 ( .A(n1293), .ZN(n1178) );
NAND4_X1 U995 ( .A1(n1294), .A2(n1112), .A3(G227), .A4(n1293), .ZN(n1290) );
NAND2_X1 U996 ( .A1(n1172), .A2(n1177), .ZN(n1293) );
NOR2_X1 U997 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
AND3_X1 U998 ( .A1(n1177), .A2(KEYINPUT44), .A3(KEYINPUT63), .ZN(n1296) );
NOR2_X1 U999 ( .A1(n1297), .A2(n1177), .ZN(n1295) );
NOR2_X1 U1000 ( .A1(n1298), .A2(n1292), .ZN(n1297) );
NOR2_X1 U1001 ( .A1(KEYINPUT63), .A2(n1172), .ZN(n1298) );
NAND2_X1 U1002 ( .A1(n1299), .A2(n1300), .ZN(n1289) );
NAND2_X1 U1003 ( .A1(G227), .A2(n1112), .ZN(n1300) );
XOR2_X1 U1004 ( .A(n1301), .B(n1177), .Z(n1299) );
INV_X1 U1005 ( .A(n1174), .ZN(n1177) );
XOR2_X1 U1006 ( .A(n1302), .B(n1303), .Z(n1174) );
XOR2_X1 U1007 ( .A(n1304), .B(n1305), .Z(n1303) );
INV_X1 U1008 ( .A(n1165), .ZN(n1305) );
XOR2_X1 U1009 ( .A(n1306), .B(n1307), .Z(n1165) );
XOR2_X1 U1010 ( .A(G137), .B(G134), .Z(n1307) );
XOR2_X1 U1011 ( .A(n1102), .B(G131), .Z(n1306) );
NOR2_X1 U1012 ( .A1(G101), .A2(KEYINPUT19), .ZN(n1304) );
XNOR2_X1 U1013 ( .A(n1103), .B(n1308), .ZN(n1302) );
XOR2_X1 U1014 ( .A(KEYINPUT26), .B(KEYINPUT10), .Z(n1103) );
NOR3_X1 U1015 ( .A1(n1292), .A2(KEYINPUT63), .A3(n1172), .ZN(n1301) );
XOR2_X1 U1016 ( .A(G110), .B(G140), .Z(n1172) );
INV_X1 U1017 ( .A(KEYINPUT44), .ZN(n1292) );
NAND2_X1 U1018 ( .A1(G221), .A2(n1256), .ZN(n1077) );
NAND2_X1 U1019 ( .A1(G234), .A2(n1309), .ZN(n1256) );
AND2_X1 U1020 ( .A1(n1196), .A2(n1310), .ZN(n1253) );
NAND2_X1 U1021 ( .A1(n1041), .A2(n1311), .ZN(n1310) );
NAND3_X1 U1022 ( .A1(G902), .A2(n1244), .A3(n1118), .ZN(n1311) );
NOR2_X1 U1023 ( .A1(n1112), .A2(G898), .ZN(n1118) );
NAND3_X1 U1024 ( .A1(n1244), .A2(n1112), .A3(G952), .ZN(n1041) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1244) );
INV_X1 U1026 ( .A(n1065), .ZN(n1196) );
NAND2_X1 U1027 ( .A1(n1064), .A2(n1063), .ZN(n1065) );
NAND2_X1 U1028 ( .A1(G214), .A2(n1312), .ZN(n1063) );
XNOR2_X1 U1029 ( .A(n1313), .B(n1082), .ZN(n1064) );
NAND2_X1 U1030 ( .A1(G210), .A2(n1312), .ZN(n1082) );
NAND2_X1 U1031 ( .A1(n1309), .A2(n1314), .ZN(n1312) );
INV_X1 U1032 ( .A(G237), .ZN(n1314) );
XOR2_X1 U1033 ( .A(n1272), .B(KEYINPUT58), .Z(n1309) );
NAND2_X1 U1034 ( .A1(KEYINPUT16), .A2(n1315), .ZN(n1313) );
XOR2_X1 U1035 ( .A(KEYINPUT28), .B(n1081), .Z(n1315) );
AND2_X1 U1036 ( .A1(n1316), .A2(n1272), .ZN(n1081) );
XOR2_X1 U1037 ( .A(n1317), .B(n1214), .Z(n1316) );
XNOR2_X1 U1038 ( .A(n1318), .B(n1319), .ZN(n1214) );
AND2_X1 U1039 ( .A1(n1112), .A2(G224), .ZN(n1319) );
NAND2_X1 U1040 ( .A1(n1320), .A2(n1321), .ZN(n1318) );
NAND2_X1 U1041 ( .A1(n1133), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1042 ( .A(n1323), .B(KEYINPUT7), .Z(n1320) );
OR2_X1 U1043 ( .A1(n1322), .A2(n1133), .ZN(n1323) );
XNOR2_X1 U1044 ( .A(G110), .B(G122), .ZN(n1133) );
XNOR2_X1 U1045 ( .A(n1131), .B(n1132), .ZN(n1322) );
XNOR2_X1 U1046 ( .A(G113), .B(n1324), .ZN(n1132) );
XOR2_X1 U1047 ( .A(G119), .B(G116), .Z(n1324) );
XOR2_X1 U1048 ( .A(G101), .B(n1308), .Z(n1131) );
XOR2_X1 U1049 ( .A(G104), .B(G107), .Z(n1308) );
XOR2_X1 U1050 ( .A(n1325), .B(n1326), .Z(n1317) );
INV_X1 U1051 ( .A(n1102), .ZN(n1326) );
XOR2_X1 U1052 ( .A(n1327), .B(n1328), .Z(n1102) );
XOR2_X1 U1053 ( .A(n1218), .B(KEYINPUT60), .Z(n1327) );
INV_X1 U1054 ( .A(G146), .ZN(n1218) );
NAND2_X1 U1055 ( .A1(KEYINPUT47), .A2(G125), .ZN(n1325) );
NOR2_X1 U1056 ( .A1(n1228), .A2(n1227), .ZN(n1071) );
XNOR2_X1 U1057 ( .A(n1329), .B(G475), .ZN(n1227) );
NAND2_X1 U1058 ( .A1(n1148), .A2(n1272), .ZN(n1329) );
INV_X1 U1059 ( .A(G902), .ZN(n1272) );
XNOR2_X1 U1060 ( .A(G143), .B(n1330), .ZN(n1148) );
XOR2_X1 U1061 ( .A(n1331), .B(n1332), .Z(n1330) );
XOR2_X1 U1062 ( .A(n1333), .B(n1334), .Z(n1332) );
XOR2_X1 U1063 ( .A(n1335), .B(n1336), .Z(n1334) );
NOR2_X1 U1064 ( .A1(G146), .A2(KEYINPUT22), .ZN(n1336) );
NAND2_X1 U1065 ( .A1(n1282), .A2(G214), .ZN(n1335) );
NOR2_X1 U1066 ( .A1(G953), .A2(G237), .ZN(n1282) );
XNOR2_X1 U1067 ( .A(n1337), .B(n1338), .ZN(n1333) );
NOR2_X1 U1068 ( .A1(KEYINPUT59), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1069 ( .A(n1246), .B(KEYINPUT1), .Z(n1339) );
INV_X1 U1070 ( .A(G122), .ZN(n1246) );
NOR2_X1 U1071 ( .A1(KEYINPUT4), .A2(G140), .ZN(n1337) );
XOR2_X1 U1072 ( .A(n1340), .B(n1341), .Z(n1331) );
XOR2_X1 U1073 ( .A(G113), .B(G104), .Z(n1341) );
XOR2_X1 U1074 ( .A(G131), .B(G125), .Z(n1340) );
INV_X1 U1075 ( .A(n1251), .ZN(n1228) );
XOR2_X1 U1076 ( .A(n1342), .B(G478), .Z(n1251) );
OR2_X1 U1077 ( .A1(n1143), .A2(G902), .ZN(n1342) );
XNOR2_X1 U1078 ( .A(n1343), .B(n1344), .ZN(n1143) );
XOR2_X1 U1079 ( .A(n1345), .B(n1328), .Z(n1344) );
XOR2_X1 U1080 ( .A(G143), .B(n1266), .Z(n1328) );
XOR2_X1 U1081 ( .A(G128), .B(KEYINPUT31), .Z(n1266) );
AND2_X1 U1082 ( .A1(n1267), .A2(G217), .ZN(n1345) );
AND2_X1 U1083 ( .A1(G234), .A2(n1112), .ZN(n1267) );
INV_X1 U1084 ( .A(G953), .ZN(n1112) );
XOR2_X1 U1085 ( .A(n1346), .B(n1347), .Z(n1343) );
NOR2_X1 U1086 ( .A1(KEYINPUT24), .A2(n1348), .ZN(n1347) );
XOR2_X1 U1087 ( .A(G107), .B(n1349), .Z(n1348) );
XOR2_X1 U1088 ( .A(G122), .B(G116), .Z(n1349) );
XNOR2_X1 U1089 ( .A(G134), .B(KEYINPUT12), .ZN(n1346) );
endmodule


