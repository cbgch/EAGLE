//Key = 1001111101111010000010111101110000100111101001110100110100111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296;

XOR2_X1 U727 ( .A(n993), .B(n994), .Z(G9) );
NAND2_X1 U728 ( .A1(KEYINPUT34), .A2(G107), .ZN(n994) );
NAND3_X1 U729 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n993) );
XNOR2_X1 U730 ( .A(n998), .B(KEYINPUT45), .ZN(n997) );
NOR2_X1 U731 ( .A1(n999), .A2(n1000), .ZN(G75) );
NOR4_X1 U732 ( .A1(n1001), .A2(n1002), .A3(G953), .A4(n1003), .ZN(n1000) );
NOR4_X1 U733 ( .A1(n1004), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n1002) );
NOR2_X1 U734 ( .A1(n1008), .A2(n1009), .ZN(n1004) );
NOR2_X1 U735 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NAND3_X1 U736 ( .A1(n1012), .A2(n1013), .A3(KEYINPUT49), .ZN(n1001) );
NAND2_X1 U737 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND3_X1 U738 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1015) );
XOR2_X1 U739 ( .A(KEYINPUT28), .B(n1019), .Z(n1018) );
NOR3_X1 U740 ( .A1(n1006), .A2(n1020), .A3(n1005), .ZN(n1019) );
INV_X1 U741 ( .A(n998), .ZN(n1005) );
NAND3_X1 U742 ( .A1(n1020), .A2(n998), .A3(n1021), .ZN(n1017) );
NOR3_X1 U743 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1021) );
NOR3_X1 U744 ( .A1(n1025), .A2(n1026), .A3(n995), .ZN(n1024) );
INV_X1 U745 ( .A(n1027), .ZN(n1025) );
NOR2_X1 U746 ( .A1(n1028), .A2(n1027), .ZN(n1023) );
NAND3_X1 U747 ( .A1(n1020), .A2(n1029), .A3(n1030), .ZN(n1016) );
INV_X1 U748 ( .A(n1006), .ZN(n1030) );
NAND3_X1 U749 ( .A1(n1028), .A2(n1027), .A3(n1031), .ZN(n1006) );
INV_X1 U750 ( .A(n1022), .ZN(n1031) );
NAND2_X1 U751 ( .A1(n1032), .A2(n1033), .ZN(n1029) );
NAND2_X1 U752 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR3_X1 U753 ( .A1(n1003), .A2(G953), .A3(G952), .ZN(n999) );
AND4_X1 U754 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1003) );
AND4_X1 U755 ( .A1(n1027), .A2(n1040), .A3(n1014), .A4(n1034), .ZN(n1039) );
XOR2_X1 U756 ( .A(n1041), .B(KEYINPUT56), .Z(n1038) );
XNOR2_X1 U757 ( .A(n1042), .B(G478), .ZN(n1037) );
XNOR2_X1 U758 ( .A(n1007), .B(KEYINPUT50), .ZN(n1036) );
NAND2_X1 U759 ( .A1(n1043), .A2(n1044), .ZN(G72) );
NAND2_X1 U760 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U761 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND2_X1 U762 ( .A1(KEYINPUT54), .A2(KEYINPUT11), .ZN(n1048) );
OR3_X1 U763 ( .A1(n1049), .A2(KEYINPUT54), .A3(n1046), .ZN(n1043) );
NAND2_X1 U764 ( .A1(G953), .A2(n1050), .ZN(n1046) );
NAND2_X1 U765 ( .A1(G900), .A2(G227), .ZN(n1050) );
XOR2_X1 U766 ( .A(n1047), .B(KEYINPUT11), .Z(n1049) );
AND2_X1 U767 ( .A1(n1051), .A2(n1052), .ZN(n1047) );
NAND3_X1 U768 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
XNOR2_X1 U769 ( .A(n1056), .B(n1057), .ZN(n1055) );
NAND2_X1 U770 ( .A1(G953), .A2(n1058), .ZN(n1054) );
NAND2_X1 U771 ( .A1(n1059), .A2(n1060), .ZN(n1053) );
NAND3_X1 U772 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1051) );
XNOR2_X1 U773 ( .A(n1057), .B(n1062), .ZN(n1061) );
INV_X1 U774 ( .A(n1056), .ZN(n1062) );
XOR2_X1 U775 ( .A(n1063), .B(n1064), .Z(G69) );
XOR2_X1 U776 ( .A(n1065), .B(n1066), .Z(n1064) );
NAND2_X1 U777 ( .A1(G953), .A2(n1067), .ZN(n1066) );
NAND2_X1 U778 ( .A1(G898), .A2(G224), .ZN(n1067) );
NAND2_X1 U779 ( .A1(n1068), .A2(n1069), .ZN(n1065) );
NAND2_X1 U780 ( .A1(G953), .A2(n1070), .ZN(n1069) );
XNOR2_X1 U781 ( .A(n1071), .B(n1072), .ZN(n1068) );
XNOR2_X1 U782 ( .A(n1073), .B(n1074), .ZN(n1071) );
NAND2_X1 U783 ( .A1(KEYINPUT23), .A2(n1075), .ZN(n1074) );
NAND2_X1 U784 ( .A1(KEYINPUT63), .A2(n1076), .ZN(n1073) );
AND2_X1 U785 ( .A1(n1077), .A2(n1060), .ZN(n1063) );
NOR2_X1 U786 ( .A1(n1078), .A2(n1079), .ZN(G66) );
NOR2_X1 U787 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U788 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U789 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
AND2_X1 U790 ( .A1(n1086), .A2(KEYINPUT12), .ZN(n1082) );
NOR2_X1 U791 ( .A1(KEYINPUT12), .A2(n1086), .ZN(n1080) );
NOR2_X1 U792 ( .A1(n1078), .A2(n1087), .ZN(G63) );
NOR3_X1 U793 ( .A1(n1042), .A2(n1088), .A3(n1089), .ZN(n1087) );
AND3_X1 U794 ( .A1(n1090), .A2(n1091), .A3(G902), .ZN(n1089) );
NOR2_X1 U795 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR3_X1 U796 ( .A1(KEYINPUT2), .A2(n1092), .A3(n1093), .ZN(n1090) );
INV_X1 U797 ( .A(G478), .ZN(n1093) );
XNOR2_X1 U798 ( .A(n1012), .B(KEYINPUT3), .ZN(n1092) );
NOR2_X1 U799 ( .A1(n1078), .A2(n1094), .ZN(G60) );
XOR2_X1 U800 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U801 ( .A1(n1097), .A2(n1085), .ZN(n1096) );
NAND2_X1 U802 ( .A1(KEYINPUT9), .A2(n1098), .ZN(n1095) );
XNOR2_X1 U803 ( .A(n1099), .B(n1100), .ZN(G6) );
NOR2_X1 U804 ( .A1(n1078), .A2(n1101), .ZN(G57) );
XOR2_X1 U805 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U806 ( .A(n1104), .B(G101), .Z(n1103) );
NAND2_X1 U807 ( .A1(KEYINPUT40), .A2(n1105), .ZN(n1102) );
XOR2_X1 U808 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U809 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U810 ( .A1(n1110), .A2(n1085), .ZN(n1109) );
NAND2_X1 U811 ( .A1(n1111), .A2(KEYINPUT25), .ZN(n1108) );
XNOR2_X1 U812 ( .A(n1112), .B(n1113), .ZN(n1111) );
NOR2_X1 U813 ( .A1(KEYINPUT18), .A2(n1114), .ZN(n1113) );
NOR2_X1 U814 ( .A1(n1078), .A2(n1115), .ZN(G54) );
XOR2_X1 U815 ( .A(n1116), .B(n1117), .Z(n1115) );
XNOR2_X1 U816 ( .A(n1118), .B(n1056), .ZN(n1117) );
XOR2_X1 U817 ( .A(n1119), .B(n1120), .Z(n1056) );
XOR2_X1 U818 ( .A(n1121), .B(n1122), .Z(n1116) );
NOR2_X1 U819 ( .A1(n1123), .A2(n1085), .ZN(n1121) );
NOR2_X1 U820 ( .A1(n1078), .A2(n1124), .ZN(G51) );
XOR2_X1 U821 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U822 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U823 ( .A1(n1129), .A2(n1085), .ZN(n1128) );
OR2_X1 U824 ( .A1(n1130), .A2(n1012), .ZN(n1085) );
NOR2_X1 U825 ( .A1(n1077), .A2(n1059), .ZN(n1012) );
NAND4_X1 U826 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1059) );
NOR4_X1 U827 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1134) );
AND2_X1 U828 ( .A1(n1139), .A2(n1140), .ZN(n1133) );
NAND2_X1 U829 ( .A1(n1141), .A2(n1009), .ZN(n1131) );
XOR2_X1 U830 ( .A(n1142), .B(KEYINPUT27), .Z(n1141) );
NAND4_X1 U831 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1077) );
NOR4_X1 U832 ( .A1(n1147), .A2(n1148), .A3(n1100), .A4(n1149), .ZN(n1146) );
INV_X1 U833 ( .A(n1150), .ZN(n1149) );
AND3_X1 U834 ( .A1(n996), .A2(n998), .A3(n1026), .ZN(n1100) );
NAND2_X1 U835 ( .A1(n996), .A2(n1151), .ZN(n1145) );
NAND2_X1 U836 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U837 ( .A1(n1154), .A2(n995), .ZN(n1153) );
XNOR2_X1 U838 ( .A(n998), .B(KEYINPUT59), .ZN(n1154) );
NAND2_X1 U839 ( .A1(n1028), .A2(n1155), .ZN(n1152) );
NAND2_X1 U840 ( .A1(n1156), .A2(n1155), .ZN(n1143) );
NAND3_X1 U841 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1127) );
OR2_X1 U842 ( .A1(n1160), .A2(KEYINPUT22), .ZN(n1159) );
NAND3_X1 U843 ( .A1(KEYINPUT22), .A2(n1160), .A3(n1161), .ZN(n1158) );
NAND2_X1 U844 ( .A1(n1162), .A2(n1163), .ZN(n1157) );
NAND2_X1 U845 ( .A1(n1164), .A2(KEYINPUT22), .ZN(n1163) );
XNOR2_X1 U846 ( .A(n1160), .B(KEYINPUT0), .ZN(n1164) );
AND2_X1 U847 ( .A1(n1165), .A2(n1166), .ZN(n1160) );
NAND2_X1 U848 ( .A1(n1112), .A2(n1167), .ZN(n1166) );
NAND2_X1 U849 ( .A1(KEYINPUT60), .A2(n1168), .ZN(n1167) );
NAND2_X1 U850 ( .A1(KEYINPUT53), .A2(n1169), .ZN(n1168) );
NAND2_X1 U851 ( .A1(G125), .A2(n1170), .ZN(n1165) );
NAND2_X1 U852 ( .A1(KEYINPUT53), .A2(n1171), .ZN(n1170) );
NAND2_X1 U853 ( .A1(KEYINPUT60), .A2(n1172), .ZN(n1171) );
NOR2_X1 U854 ( .A1(n1060), .A2(G952), .ZN(n1078) );
XOR2_X1 U855 ( .A(G146), .B(n1135), .Z(G48) );
AND4_X1 U856 ( .A1(n1173), .A2(n1026), .A3(n1009), .A4(n1174), .ZN(n1135) );
XNOR2_X1 U857 ( .A(n1175), .B(n1132), .ZN(G45) );
NAND4_X1 U858 ( .A1(n1176), .A2(n1009), .A3(n1177), .A4(n1178), .ZN(n1132) );
NAND2_X1 U859 ( .A1(KEYINPUT52), .A2(n1179), .ZN(n1175) );
XOR2_X1 U860 ( .A(n1140), .B(n1180), .Z(G42) );
XOR2_X1 U861 ( .A(KEYINPUT14), .B(G140), .Z(n1180) );
NAND4_X1 U862 ( .A1(n1173), .A2(n1026), .A3(n1034), .A4(n1014), .ZN(n1140) );
XNOR2_X1 U863 ( .A(G137), .B(n1139), .ZN(G39) );
NAND4_X1 U864 ( .A1(n1173), .A2(n1028), .A3(n1014), .A4(n1174), .ZN(n1139) );
XOR2_X1 U865 ( .A(G134), .B(n1138), .Z(G36) );
AND3_X1 U866 ( .A1(n1014), .A2(n995), .A3(n1176), .ZN(n1138) );
XNOR2_X1 U867 ( .A(n1181), .B(n1137), .ZN(G33) );
AND3_X1 U868 ( .A1(n1026), .A2(n1014), .A3(n1176), .ZN(n1137) );
AND4_X1 U869 ( .A1(n1155), .A2(n1007), .A3(n1182), .A4(n1027), .ZN(n1176) );
NOR2_X1 U870 ( .A1(n1010), .A2(n1183), .ZN(n1014) );
INV_X1 U871 ( .A(n1011), .ZN(n1183) );
XNOR2_X1 U872 ( .A(n1136), .B(n1184), .ZN(G30) );
NAND2_X1 U873 ( .A1(KEYINPUT47), .A2(G128), .ZN(n1184) );
AND4_X1 U874 ( .A1(n1173), .A2(n995), .A3(n1009), .A4(n1174), .ZN(n1136) );
AND4_X1 U875 ( .A1(n1007), .A2(n1035), .A3(n1182), .A4(n1027), .ZN(n1173) );
XOR2_X1 U876 ( .A(G101), .B(n1185), .Z(G3) );
NOR3_X1 U877 ( .A1(n1032), .A2(n1186), .A3(n1187), .ZN(n1185) );
XNOR2_X1 U878 ( .A(n1028), .B(KEYINPUT51), .ZN(n1186) );
XNOR2_X1 U879 ( .A(n1169), .B(n1188), .ZN(G27) );
NOR2_X1 U880 ( .A1(n1189), .A2(n1142), .ZN(n1188) );
NAND4_X1 U881 ( .A1(n1020), .A2(n1034), .A3(n1026), .A4(n1190), .ZN(n1142) );
AND3_X1 U882 ( .A1(n1035), .A2(n1027), .A3(n1182), .ZN(n1190) );
NAND2_X1 U883 ( .A1(n1022), .A2(n1191), .ZN(n1182) );
NAND4_X1 U884 ( .A1(G953), .A2(G902), .A3(n1192), .A4(n1058), .ZN(n1191) );
INV_X1 U885 ( .A(G900), .ZN(n1058) );
XNOR2_X1 U886 ( .A(n1148), .B(n1193), .ZN(G24) );
XNOR2_X1 U887 ( .A(G122), .B(KEYINPUT21), .ZN(n1193) );
AND4_X1 U888 ( .A1(n1194), .A2(n998), .A3(n1177), .A4(n1178), .ZN(n1148) );
NOR2_X1 U889 ( .A1(n1174), .A2(n1035), .ZN(n998) );
XNOR2_X1 U890 ( .A(G119), .B(n1195), .ZN(G21) );
NOR2_X1 U891 ( .A1(KEYINPUT26), .A2(n1196), .ZN(n1195) );
INV_X1 U892 ( .A(n1144), .ZN(n1196) );
NAND4_X1 U893 ( .A1(n1028), .A2(n1194), .A3(n1035), .A4(n1174), .ZN(n1144) );
XOR2_X1 U894 ( .A(G116), .B(n1147), .Z(G18) );
AND3_X1 U895 ( .A1(n1155), .A2(n995), .A3(n1194), .ZN(n1147) );
AND2_X1 U896 ( .A1(n1040), .A2(n1177), .ZN(n995) );
NAND2_X1 U897 ( .A1(n1197), .A2(n1198), .ZN(G15) );
NAND3_X1 U898 ( .A1(n1199), .A2(n1200), .A3(n1156), .ZN(n1198) );
XOR2_X1 U899 ( .A(n1201), .B(KEYINPUT61), .Z(n1197) );
NAND2_X1 U900 ( .A1(G113), .A2(n1202), .ZN(n1201) );
NAND2_X1 U901 ( .A1(n1156), .A2(n1199), .ZN(n1202) );
XNOR2_X1 U902 ( .A(n1032), .B(KEYINPUT35), .ZN(n1199) );
INV_X1 U903 ( .A(n1155), .ZN(n1032) );
NOR2_X1 U904 ( .A1(n1035), .A2(n1034), .ZN(n1155) );
AND2_X1 U905 ( .A1(n1026), .A2(n1194), .ZN(n1156) );
AND4_X1 U906 ( .A1(n1020), .A2(n1009), .A3(n1027), .A4(n1203), .ZN(n1194) );
INV_X1 U907 ( .A(n1007), .ZN(n1020) );
NOR2_X1 U908 ( .A1(n1177), .A2(n1040), .ZN(n1026) );
INV_X1 U909 ( .A(n1178), .ZN(n1040) );
XOR2_X1 U910 ( .A(G110), .B(n1204), .Z(G12) );
NOR2_X1 U911 ( .A1(KEYINPUT33), .A2(n1150), .ZN(n1204) );
NAND4_X1 U912 ( .A1(n1028), .A2(n996), .A3(n1034), .A4(n1035), .ZN(n1150) );
XNOR2_X1 U913 ( .A(n1041), .B(KEYINPUT43), .ZN(n1035) );
XNOR2_X1 U914 ( .A(n1205), .B(n1084), .ZN(n1041) );
NAND2_X1 U915 ( .A1(G217), .A2(n1206), .ZN(n1084) );
NAND2_X1 U916 ( .A1(n1086), .A2(n1130), .ZN(n1205) );
XOR2_X1 U917 ( .A(n1207), .B(n1208), .Z(n1086) );
XOR2_X1 U918 ( .A(n1209), .B(n1210), .Z(n1208) );
XNOR2_X1 U919 ( .A(n1211), .B(n1212), .ZN(n1210) );
NOR2_X1 U920 ( .A1(G110), .A2(KEYINPUT17), .ZN(n1212) );
NOR2_X1 U921 ( .A1(KEYINPUT57), .A2(n1213), .ZN(n1211) );
XNOR2_X1 U922 ( .A(KEYINPUT4), .B(n1214), .ZN(n1213) );
NAND2_X1 U923 ( .A1(G221), .A2(n1215), .ZN(n1209) );
XNOR2_X1 U924 ( .A(G119), .B(n1216), .ZN(n1207) );
XOR2_X1 U925 ( .A(G137), .B(G128), .Z(n1216) );
INV_X1 U926 ( .A(n1174), .ZN(n1034) );
XOR2_X1 U927 ( .A(n1217), .B(n1110), .Z(n1174) );
INV_X1 U928 ( .A(G472), .ZN(n1110) );
NAND2_X1 U929 ( .A1(n1218), .A2(n1130), .ZN(n1217) );
XOR2_X1 U930 ( .A(n1219), .B(n1220), .Z(n1218) );
XNOR2_X1 U931 ( .A(n1114), .B(n1221), .ZN(n1220) );
XNOR2_X1 U932 ( .A(n1104), .B(n1222), .ZN(n1221) );
NOR2_X1 U933 ( .A1(G101), .A2(KEYINPUT48), .ZN(n1222) );
NAND3_X1 U934 ( .A1(n1223), .A2(n1060), .A3(G210), .ZN(n1104) );
INV_X1 U935 ( .A(n1119), .ZN(n1114) );
XNOR2_X1 U936 ( .A(n1106), .B(n1172), .ZN(n1219) );
INV_X1 U937 ( .A(n1112), .ZN(n1172) );
XNOR2_X1 U938 ( .A(n1224), .B(n1225), .ZN(n1106) );
XOR2_X1 U939 ( .A(n1226), .B(G119), .Z(n1224) );
NAND2_X1 U940 ( .A1(KEYINPUT20), .A2(G116), .ZN(n1226) );
INV_X1 U941 ( .A(n1187), .ZN(n996) );
NAND4_X1 U942 ( .A1(n1009), .A2(n1007), .A3(n1027), .A4(n1203), .ZN(n1187) );
NAND2_X1 U943 ( .A1(n1022), .A2(n1227), .ZN(n1203) );
NAND4_X1 U944 ( .A1(G953), .A2(G902), .A3(n1192), .A4(n1070), .ZN(n1227) );
INV_X1 U945 ( .A(G898), .ZN(n1070) );
NAND3_X1 U946 ( .A1(n1192), .A2(n1060), .A3(G952), .ZN(n1022) );
NAND2_X1 U947 ( .A1(G237), .A2(G234), .ZN(n1192) );
NAND2_X1 U948 ( .A1(G221), .A2(n1206), .ZN(n1027) );
NAND2_X1 U949 ( .A1(G234), .A2(n1130), .ZN(n1206) );
XOR2_X1 U950 ( .A(n1228), .B(n1123), .Z(n1007) );
INV_X1 U951 ( .A(G469), .ZN(n1123) );
NAND2_X1 U952 ( .A1(n1229), .A2(n1130), .ZN(n1228) );
XNOR2_X1 U953 ( .A(n1122), .B(n1230), .ZN(n1229) );
XOR2_X1 U954 ( .A(n1231), .B(KEYINPUT13), .Z(n1230) );
NAND2_X1 U955 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
OR2_X1 U956 ( .A1(n1119), .A2(n1234), .ZN(n1233) );
XOR2_X1 U957 ( .A(n1235), .B(KEYINPUT31), .Z(n1232) );
NAND2_X1 U958 ( .A1(n1234), .A2(n1119), .ZN(n1235) );
XOR2_X1 U959 ( .A(G131), .B(n1236), .Z(n1119) );
XOR2_X1 U960 ( .A(G137), .B(G134), .Z(n1236) );
XNOR2_X1 U961 ( .A(n1237), .B(n1120), .ZN(n1234) );
XOR2_X1 U962 ( .A(G128), .B(n1238), .Z(n1120) );
NOR2_X1 U963 ( .A1(KEYINPUT19), .A2(n1239), .ZN(n1238) );
NAND2_X1 U964 ( .A1(KEYINPUT37), .A2(n1118), .ZN(n1237) );
XOR2_X1 U965 ( .A(n1240), .B(G104), .Z(n1118) );
XNOR2_X1 U966 ( .A(n1241), .B(n1242), .ZN(n1122) );
XOR2_X1 U967 ( .A(G140), .B(G110), .Z(n1242) );
NAND2_X1 U968 ( .A1(G227), .A2(n1060), .ZN(n1241) );
INV_X1 U969 ( .A(n1189), .ZN(n1009) );
NAND2_X1 U970 ( .A1(n1010), .A2(n1011), .ZN(n1189) );
NAND2_X1 U971 ( .A1(n1243), .A2(n1244), .ZN(n1011) );
XNOR2_X1 U972 ( .A(G214), .B(KEYINPUT42), .ZN(n1243) );
XNOR2_X1 U973 ( .A(n1129), .B(n1245), .ZN(n1010) );
NOR2_X1 U974 ( .A1(G902), .A2(n1246), .ZN(n1245) );
XOR2_X1 U975 ( .A(n1125), .B(n1247), .Z(n1246) );
NOR3_X1 U976 ( .A1(KEYINPUT1), .A2(n1248), .A3(n1249), .ZN(n1247) );
NOR2_X1 U977 ( .A1(n1169), .A2(n1250), .ZN(n1249) );
XNOR2_X1 U978 ( .A(n1251), .B(KEYINPUT7), .ZN(n1250) );
INV_X1 U979 ( .A(G125), .ZN(n1169) );
NOR2_X1 U980 ( .A1(G125), .A2(n1252), .ZN(n1248) );
XOR2_X1 U981 ( .A(n1251), .B(n1253), .Z(n1252) );
XOR2_X1 U982 ( .A(KEYINPUT36), .B(KEYINPUT29), .Z(n1253) );
XOR2_X1 U983 ( .A(n1162), .B(n1112), .Z(n1251) );
XOR2_X1 U984 ( .A(n1254), .B(n1239), .Z(n1112) );
XNOR2_X1 U985 ( .A(G146), .B(G143), .ZN(n1239) );
XNOR2_X1 U986 ( .A(G128), .B(KEYINPUT58), .ZN(n1254) );
INV_X1 U987 ( .A(n1161), .ZN(n1162) );
NAND2_X1 U988 ( .A1(G224), .A2(n1060), .ZN(n1161) );
XOR2_X1 U989 ( .A(n1072), .B(n1255), .Z(n1125) );
XOR2_X1 U990 ( .A(n1076), .B(n1075), .Z(n1255) );
XNOR2_X1 U991 ( .A(G110), .B(n1256), .ZN(n1075) );
XNOR2_X1 U992 ( .A(KEYINPUT39), .B(n1257), .ZN(n1256) );
NAND2_X1 U993 ( .A1(n1258), .A2(n1259), .ZN(n1076) );
NAND2_X1 U994 ( .A1(n1225), .A2(n1260), .ZN(n1259) );
XOR2_X1 U995 ( .A(n1261), .B(KEYINPUT44), .Z(n1258) );
OR2_X1 U996 ( .A1(n1260), .A2(n1225), .ZN(n1261) );
XOR2_X1 U997 ( .A(G116), .B(G119), .Z(n1260) );
NAND2_X1 U998 ( .A1(n1262), .A2(n1263), .ZN(n1072) );
NAND2_X1 U999 ( .A1(n1264), .A2(n1099), .ZN(n1263) );
INV_X1 U1000 ( .A(G104), .ZN(n1099) );
XOR2_X1 U1001 ( .A(n1240), .B(KEYINPUT32), .Z(n1264) );
NAND2_X1 U1002 ( .A1(G104), .A2(n1265), .ZN(n1262) );
XOR2_X1 U1003 ( .A(n1240), .B(KEYINPUT46), .Z(n1265) );
XOR2_X1 U1004 ( .A(G101), .B(n1266), .Z(n1240) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1244), .ZN(n1129) );
NAND2_X1 U1006 ( .A1(n1223), .A2(n1130), .ZN(n1244) );
NOR2_X1 U1007 ( .A1(n1178), .A2(n1177), .ZN(n1028) );
XNOR2_X1 U1008 ( .A(n1042), .B(n1267), .ZN(n1177) );
NOR2_X1 U1009 ( .A1(G478), .A2(KEYINPUT15), .ZN(n1267) );
NOR2_X1 U1010 ( .A1(n1091), .A2(G902), .ZN(n1042) );
XNOR2_X1 U1011 ( .A(n1268), .B(n1269), .ZN(n1091) );
XOR2_X1 U1012 ( .A(n1270), .B(n1271), .Z(n1269) );
NAND2_X1 U1013 ( .A1(G217), .A2(n1215), .ZN(n1271) );
AND2_X1 U1014 ( .A1(G234), .A2(n1060), .ZN(n1215) );
NAND2_X1 U1015 ( .A1(n1272), .A2(KEYINPUT5), .ZN(n1270) );
XOR2_X1 U1016 ( .A(n1273), .B(n1274), .Z(n1272) );
NOR2_X1 U1017 ( .A1(KEYINPUT16), .A2(n1266), .ZN(n1274) );
XNOR2_X1 U1018 ( .A(G107), .B(KEYINPUT55), .ZN(n1266) );
NAND2_X1 U1019 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
NAND2_X1 U1020 ( .A1(G116), .A2(n1257), .ZN(n1276) );
XOR2_X1 U1021 ( .A(KEYINPUT24), .B(n1277), .Z(n1275) );
NOR2_X1 U1022 ( .A1(G116), .A2(n1257), .ZN(n1277) );
XNOR2_X1 U1023 ( .A(G128), .B(n1278), .ZN(n1268) );
XNOR2_X1 U1024 ( .A(n1179), .B(G134), .ZN(n1278) );
XNOR2_X1 U1025 ( .A(n1279), .B(n1280), .ZN(n1178) );
XNOR2_X1 U1026 ( .A(KEYINPUT30), .B(n1097), .ZN(n1280) );
INV_X1 U1027 ( .A(G475), .ZN(n1097) );
NAND2_X1 U1028 ( .A1(n1098), .A2(n1130), .ZN(n1279) );
INV_X1 U1029 ( .A(G902), .ZN(n1130) );
XOR2_X1 U1030 ( .A(n1281), .B(n1282), .Z(n1098) );
XOR2_X1 U1031 ( .A(n1283), .B(n1284), .Z(n1282) );
XNOR2_X1 U1032 ( .A(n1257), .B(G104), .ZN(n1284) );
INV_X1 U1033 ( .A(G122), .ZN(n1257) );
XNOR2_X1 U1034 ( .A(KEYINPUT8), .B(n1181), .ZN(n1283) );
INV_X1 U1035 ( .A(G131), .ZN(n1181) );
XNOR2_X1 U1036 ( .A(n1285), .B(n1225), .ZN(n1281) );
XOR2_X1 U1037 ( .A(n1200), .B(KEYINPUT38), .Z(n1225) );
INV_X1 U1038 ( .A(G113), .ZN(n1200) );
XNOR2_X1 U1039 ( .A(n1286), .B(n1287), .ZN(n1285) );
NAND2_X1 U1040 ( .A1(KEYINPUT10), .A2(n1214), .ZN(n1287) );
XNOR2_X1 U1041 ( .A(G146), .B(n1057), .ZN(n1214) );
XOR2_X1 U1042 ( .A(G140), .B(G125), .Z(n1057) );
NAND3_X1 U1043 ( .A1(n1288), .A2(n1289), .A3(KEYINPUT6), .ZN(n1286) );
NAND2_X1 U1044 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
INV_X1 U1045 ( .A(KEYINPUT41), .ZN(n1291) );
NAND2_X1 U1046 ( .A1(n1292), .A2(n1293), .ZN(n1290) );
NAND2_X1 U1047 ( .A1(n1294), .A2(n1179), .ZN(n1293) );
INV_X1 U1048 ( .A(G143), .ZN(n1179) );
NAND2_X1 U1049 ( .A1(n1295), .A2(n1296), .ZN(n1292) );
XNOR2_X1 U1050 ( .A(G143), .B(KEYINPUT62), .ZN(n1295) );
NAND3_X1 U1051 ( .A1(G143), .A2(n1294), .A3(KEYINPUT41), .ZN(n1288) );
INV_X1 U1052 ( .A(n1296), .ZN(n1294) );
NAND3_X1 U1053 ( .A1(n1223), .A2(n1060), .A3(G214), .ZN(n1296) );
INV_X1 U1054 ( .A(G953), .ZN(n1060) );
INV_X1 U1055 ( .A(G237), .ZN(n1223) );
endmodule


