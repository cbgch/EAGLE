//Key = 0101010110101010101010111110000011111011000000101101101001100011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276;

XNOR2_X1 U699 ( .A(G107), .B(n972), .ZN(G9) );
NAND3_X1 U700 ( .A1(n973), .A2(n974), .A3(n975), .ZN(n972) );
XNOR2_X1 U701 ( .A(n976), .B(KEYINPUT38), .ZN(n975) );
NOR2_X1 U702 ( .A1(n977), .A2(n978), .ZN(G75) );
NOR4_X1 U703 ( .A1(n979), .A2(n980), .A3(n981), .A4(n982), .ZN(n978) );
XOR2_X1 U704 ( .A(n983), .B(KEYINPUT45), .Z(n982) );
NAND2_X1 U705 ( .A1(n984), .A2(n985), .ZN(n983) );
NAND3_X1 U706 ( .A1(n986), .A2(n987), .A3(n988), .ZN(n985) );
NAND3_X1 U707 ( .A1(n989), .A2(n990), .A3(n991), .ZN(n987) );
NAND3_X1 U708 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
NAND4_X1 U709 ( .A1(n995), .A2(n996), .A3(n974), .A4(n997), .ZN(n990) );
XOR2_X1 U710 ( .A(KEYINPUT40), .B(n994), .Z(n997) );
OR3_X1 U711 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n989) );
NAND2_X1 U712 ( .A1(n1001), .A2(n976), .ZN(n984) );
AND2_X1 U713 ( .A1(n1002), .A2(n1001), .ZN(n981) );
NOR3_X1 U714 ( .A1(n1003), .A2(n998), .A3(n1004), .ZN(n1001) );
NAND3_X1 U715 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n979) );
NAND3_X1 U716 ( .A1(n986), .A2(n1008), .A3(n988), .ZN(n1007) );
INV_X1 U717 ( .A(n1004), .ZN(n988) );
NAND2_X1 U718 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND2_X1 U719 ( .A1(n994), .A2(n1011), .ZN(n1010) );
NAND2_X1 U720 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND2_X1 U721 ( .A1(n974), .A2(n1014), .ZN(n1013) );
NAND2_X1 U722 ( .A1(n1015), .A2(n1016), .ZN(n1012) );
XOR2_X1 U723 ( .A(KEYINPUT4), .B(n993), .Z(n1015) );
NAND2_X1 U724 ( .A1(n1017), .A2(n1018), .ZN(n1009) );
INV_X1 U725 ( .A(n998), .ZN(n1017) );
NOR3_X1 U726 ( .A1(n1019), .A2(G953), .A3(G952), .ZN(n977) );
INV_X1 U727 ( .A(n1005), .ZN(n1019) );
NAND4_X1 U728 ( .A1(n1020), .A2(n999), .A3(n1021), .A4(n1022), .ZN(n1005) );
NOR2_X1 U729 ( .A1(n998), .A2(n1023), .ZN(n1022) );
XOR2_X1 U730 ( .A(G478), .B(n1024), .Z(n1023) );
NAND2_X1 U731 ( .A1(n993), .A2(n974), .ZN(n998) );
XOR2_X1 U732 ( .A(KEYINPUT57), .B(n1025), .Z(n1020) );
XOR2_X1 U733 ( .A(n1026), .B(n1027), .Z(G72) );
NOR3_X1 U734 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
NOR2_X1 U735 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
XOR2_X1 U736 ( .A(n1033), .B(KEYINPUT23), .Z(n1028) );
NAND2_X1 U737 ( .A1(n1031), .A2(n1032), .ZN(n1033) );
XOR2_X1 U738 ( .A(n1034), .B(n1035), .Z(n1032) );
NOR2_X1 U739 ( .A1(G131), .A2(KEYINPUT43), .ZN(n1035) );
XNOR2_X1 U740 ( .A(n1036), .B(n1037), .ZN(n1031) );
XNOR2_X1 U741 ( .A(G140), .B(KEYINPUT30), .ZN(n1036) );
NAND2_X1 U742 ( .A1(n1038), .A2(n1039), .ZN(n1026) );
NAND2_X1 U743 ( .A1(n1040), .A2(n1006), .ZN(n1039) );
NAND2_X1 U744 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
XNOR2_X1 U745 ( .A(n1043), .B(KEYINPUT3), .ZN(n1041) );
NAND2_X1 U746 ( .A1(n1044), .A2(G953), .ZN(n1038) );
XOR2_X1 U747 ( .A(KEYINPUT62), .B(n1045), .Z(n1044) );
NOR2_X1 U748 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
XOR2_X1 U749 ( .A(n1048), .B(n1049), .Z(G69) );
XOR2_X1 U750 ( .A(n1050), .B(n1051), .Z(n1049) );
NOR2_X1 U751 ( .A1(G953), .A2(n1052), .ZN(n1051) );
NAND3_X1 U752 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1050) );
XOR2_X1 U753 ( .A(n1056), .B(KEYINPUT6), .Z(n1055) );
NAND2_X1 U754 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
OR2_X1 U755 ( .A1(n1058), .A2(n1057), .ZN(n1054) );
XOR2_X1 U756 ( .A(n1059), .B(n1060), .Z(n1057) );
NAND2_X1 U757 ( .A1(n1061), .A2(n1062), .ZN(n1053) );
NAND2_X1 U758 ( .A1(G953), .A2(n1063), .ZN(n1048) );
NAND2_X1 U759 ( .A1(G898), .A2(G224), .ZN(n1063) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(G66) );
XOR2_X1 U761 ( .A(n1066), .B(n1067), .Z(n1065) );
NOR2_X1 U762 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U763 ( .A1(n1064), .A2(n1070), .ZN(G63) );
NOR3_X1 U764 ( .A1(n1024), .A2(n1071), .A3(n1072), .ZN(n1070) );
AND3_X1 U765 ( .A1(n1073), .A2(G478), .A3(n1074), .ZN(n1072) );
NOR2_X1 U766 ( .A1(n1075), .A2(n1073), .ZN(n1071) );
AND2_X1 U767 ( .A1(n980), .A2(G478), .ZN(n1075) );
NOR2_X1 U768 ( .A1(n1064), .A2(n1076), .ZN(G60) );
XOR2_X1 U769 ( .A(n1077), .B(n1078), .Z(n1076) );
NAND3_X1 U770 ( .A1(n1074), .A2(G475), .A3(KEYINPUT36), .ZN(n1077) );
NAND2_X1 U771 ( .A1(n1079), .A2(n1080), .ZN(G6) );
NAND2_X1 U772 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U773 ( .A1(G104), .A2(n1083), .ZN(n1079) );
NAND2_X1 U774 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U775 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
OR2_X1 U776 ( .A1(n1087), .A2(n1081), .ZN(n1084) );
NOR2_X1 U777 ( .A1(KEYINPUT50), .A2(n1088), .ZN(n1081) );
INV_X1 U778 ( .A(KEYINPUT18), .ZN(n1087) );
NOR2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(G57) );
XNOR2_X1 U780 ( .A(n1091), .B(n1092), .ZN(n1090) );
XOR2_X1 U781 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U782 ( .A1(n1095), .A2(KEYINPUT15), .ZN(n1094) );
AND2_X1 U783 ( .A1(G472), .A2(n1074), .ZN(n1095) );
NOR2_X1 U784 ( .A1(G952), .A2(n1096), .ZN(n1089) );
XOR2_X1 U785 ( .A(n1006), .B(KEYINPUT13), .Z(n1096) );
NOR2_X1 U786 ( .A1(n1064), .A2(n1097), .ZN(G54) );
NOR2_X1 U787 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U788 ( .A(n1100), .B(KEYINPUT26), .Z(n1099) );
NAND2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U790 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
XNOR2_X1 U791 ( .A(n1103), .B(n1104), .ZN(n1102) );
NAND2_X1 U792 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NAND2_X1 U793 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U794 ( .A1(G227), .A2(n1006), .ZN(n1108) );
XOR2_X1 U795 ( .A(KEYINPUT63), .B(n1109), .Z(n1105) );
AND2_X1 U796 ( .A1(n1074), .A2(G469), .ZN(n1101) );
NOR2_X1 U797 ( .A1(n1064), .A2(n1110), .ZN(G51) );
XOR2_X1 U798 ( .A(n1111), .B(n1112), .Z(n1110) );
NAND2_X1 U799 ( .A1(n1074), .A2(n1113), .ZN(n1112) );
INV_X1 U800 ( .A(n1069), .ZN(n1074) );
NAND2_X1 U801 ( .A1(G902), .A2(n980), .ZN(n1069) );
NAND3_X1 U802 ( .A1(n1052), .A2(n1042), .A3(n1043), .ZN(n980) );
AND4_X1 U803 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1043) );
NAND2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
INV_X1 U805 ( .A(n1120), .ZN(n1119) );
XOR2_X1 U806 ( .A(n1121), .B(KEYINPUT46), .Z(n1118) );
NAND3_X1 U807 ( .A1(n1014), .A2(n1122), .A3(n1123), .ZN(n1114) );
XOR2_X1 U808 ( .A(KEYINPUT19), .B(n994), .Z(n1122) );
AND4_X1 U809 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1042) );
AND2_X1 U810 ( .A1(n1128), .A2(n1129), .ZN(n1052) );
AND4_X1 U811 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1129) );
NOR4_X1 U812 ( .A1(n1134), .A2(n1086), .A3(n1135), .A4(n1136), .ZN(n1128) );
NOR2_X1 U813 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U814 ( .A(KEYINPUT5), .B(n1018), .Z(n1138) );
AND3_X1 U815 ( .A1(n973), .A2(n976), .A3(n974), .ZN(n1135) );
INV_X1 U816 ( .A(n1088), .ZN(n1086) );
NAND3_X1 U817 ( .A1(n973), .A2(n974), .A3(n1002), .ZN(n1088) );
INV_X1 U818 ( .A(n1139), .ZN(n1134) );
NAND2_X1 U819 ( .A1(n1140), .A2(n1141), .ZN(n1111) );
NAND2_X1 U820 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XOR2_X1 U821 ( .A(KEYINPUT11), .B(n1144), .Z(n1143) );
XOR2_X1 U822 ( .A(KEYINPUT52), .B(n1145), .Z(n1140) );
NOR2_X1 U823 ( .A1(n1142), .A2(n1144), .ZN(n1145) );
XOR2_X1 U824 ( .A(n1146), .B(KEYINPUT47), .Z(n1144) );
NOR2_X1 U825 ( .A1(n1006), .A2(G952), .ZN(n1064) );
XOR2_X1 U826 ( .A(n1147), .B(n1116), .Z(G48) );
NAND3_X1 U827 ( .A1(n1148), .A2(n1018), .A3(n1002), .ZN(n1116) );
XNOR2_X1 U828 ( .A(n1149), .B(n1117), .ZN(G45) );
NAND4_X1 U829 ( .A1(n1150), .A2(n1151), .A3(n1018), .A4(n1152), .ZN(n1117) );
NOR2_X1 U830 ( .A1(KEYINPUT0), .A2(n1153), .ZN(n1149) );
XOR2_X1 U831 ( .A(n1154), .B(KEYINPUT42), .Z(n1153) );
XNOR2_X1 U832 ( .A(G140), .B(n1155), .ZN(G42) );
NAND3_X1 U833 ( .A1(n1123), .A2(n1014), .A3(n1156), .ZN(n1155) );
XOR2_X1 U834 ( .A(n1003), .B(KEYINPUT51), .Z(n1156) );
INV_X1 U835 ( .A(n994), .ZN(n1003) );
XOR2_X1 U836 ( .A(G137), .B(n1157), .Z(G39) );
NOR2_X1 U837 ( .A1(n1121), .A2(n1120), .ZN(n1157) );
NAND2_X1 U838 ( .A1(n994), .A2(n1148), .ZN(n1120) );
NAND2_X1 U839 ( .A1(n1158), .A2(n1159), .ZN(G36) );
NAND2_X1 U840 ( .A1(n1160), .A2(n1124), .ZN(n1159) );
XOR2_X1 U841 ( .A(n1161), .B(KEYINPUT37), .Z(n1158) );
OR2_X1 U842 ( .A1(n1124), .A2(n1160), .ZN(n1161) );
XNOR2_X1 U843 ( .A(G134), .B(KEYINPUT20), .ZN(n1160) );
NAND3_X1 U844 ( .A1(n1151), .A2(n976), .A3(n994), .ZN(n1124) );
XOR2_X1 U845 ( .A(n1162), .B(n1125), .Z(G33) );
NAND3_X1 U846 ( .A1(n1002), .A2(n1151), .A3(n994), .ZN(n1125) );
NOR2_X1 U847 ( .A1(n1000), .A2(n1163), .ZN(n994) );
AND3_X1 U848 ( .A1(n1016), .A2(n1164), .A3(n1014), .ZN(n1151) );
XOR2_X1 U849 ( .A(G128), .B(n1165), .Z(G30) );
NOR2_X1 U850 ( .A1(KEYINPUT27), .A2(n1126), .ZN(n1165) );
NAND3_X1 U851 ( .A1(n976), .A2(n1018), .A3(n1148), .ZN(n1126) );
AND3_X1 U852 ( .A1(n1166), .A2(n1164), .A3(n1014), .ZN(n1148) );
XOR2_X1 U853 ( .A(n1167), .B(n1139), .Z(G3) );
NAND3_X1 U854 ( .A1(n973), .A2(n1016), .A3(n986), .ZN(n1139) );
XNOR2_X1 U855 ( .A(G125), .B(n1127), .ZN(G27) );
NAND3_X1 U856 ( .A1(n993), .A2(n1018), .A3(n1123), .ZN(n1127) );
AND3_X1 U857 ( .A1(n992), .A2(n1164), .A3(n1002), .ZN(n1123) );
NAND2_X1 U858 ( .A1(n1004), .A2(n1168), .ZN(n1164) );
NAND3_X1 U859 ( .A1(G902), .A2(n1169), .A3(n1029), .ZN(n1168) );
AND2_X1 U860 ( .A1(n1061), .A2(n1047), .ZN(n1029) );
INV_X1 U861 ( .A(G900), .ZN(n1047) );
XOR2_X1 U862 ( .A(n1170), .B(n1133), .Z(G24) );
NAND4_X1 U863 ( .A1(n1171), .A2(n974), .A3(n1150), .A4(n1152), .ZN(n1133) );
XOR2_X1 U864 ( .A(G119), .B(n1172), .Z(G21) );
NOR2_X1 U865 ( .A1(KEYINPUT28), .A2(n1132), .ZN(n1172) );
NAND3_X1 U866 ( .A1(n986), .A2(n1166), .A3(n1171), .ZN(n1132) );
NAND2_X1 U867 ( .A1(n1173), .A2(n1174), .ZN(n1166) );
NAND3_X1 U868 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1174) );
INV_X1 U869 ( .A(KEYINPUT61), .ZN(n1177) );
NAND2_X1 U870 ( .A1(KEYINPUT61), .A2(n992), .ZN(n1173) );
NAND2_X1 U871 ( .A1(n1178), .A2(n1179), .ZN(G18) );
NAND2_X1 U872 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U873 ( .A(KEYINPUT49), .B(n1182), .Z(n1178) );
NOR2_X1 U874 ( .A1(n1180), .A2(n1181), .ZN(n1182) );
AND2_X1 U875 ( .A1(n1183), .A2(n1018), .ZN(n1180) );
XOR2_X1 U876 ( .A(n1137), .B(KEYINPUT33), .Z(n1183) );
NAND4_X1 U877 ( .A1(n993), .A2(n976), .A3(n1016), .A4(n1184), .ZN(n1137) );
AND2_X1 U878 ( .A1(n1150), .A2(n1185), .ZN(n976) );
XOR2_X1 U879 ( .A(n1186), .B(G113), .Z(G15) );
NAND2_X1 U880 ( .A1(KEYINPUT48), .A2(n1131), .ZN(n1186) );
NAND3_X1 U881 ( .A1(n1002), .A2(n1016), .A3(n1171), .ZN(n1131) );
AND3_X1 U882 ( .A1(n1018), .A2(n1184), .A3(n993), .ZN(n1171) );
NOR2_X1 U883 ( .A1(n1187), .A2(n996), .ZN(n993) );
INV_X1 U884 ( .A(n995), .ZN(n1187) );
NAND2_X1 U885 ( .A1(n1188), .A2(n1189), .ZN(n1016) );
OR3_X1 U886 ( .A1(n1190), .A2(n1175), .A3(KEYINPUT61), .ZN(n1189) );
NAND2_X1 U887 ( .A1(KEYINPUT61), .A2(n974), .ZN(n1188) );
NOR2_X1 U888 ( .A1(n1176), .A2(n1175), .ZN(n974) );
INV_X1 U889 ( .A(n1190), .ZN(n1176) );
AND2_X1 U890 ( .A1(n1152), .A2(n1191), .ZN(n1002) );
XNOR2_X1 U891 ( .A(n1185), .B(KEYINPUT55), .ZN(n1152) );
XNOR2_X1 U892 ( .A(G110), .B(n1130), .ZN(G12) );
NAND3_X1 U893 ( .A1(n992), .A2(n973), .A3(n986), .ZN(n1130) );
INV_X1 U894 ( .A(n1121), .ZN(n986) );
NAND2_X1 U895 ( .A1(n1185), .A2(n1191), .ZN(n1121) );
INV_X1 U896 ( .A(n1150), .ZN(n1191) );
XNOR2_X1 U897 ( .A(n1024), .B(n1192), .ZN(n1150) );
NOR2_X1 U898 ( .A1(G478), .A2(KEYINPUT17), .ZN(n1192) );
NOR2_X1 U899 ( .A1(n1073), .A2(G902), .ZN(n1024) );
AND2_X1 U900 ( .A1(n1193), .A2(n1194), .ZN(n1073) );
NAND2_X1 U901 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NAND2_X1 U902 ( .A1(n1197), .A2(G217), .ZN(n1196) );
NAND3_X1 U903 ( .A1(n1197), .A2(G217), .A3(n1198), .ZN(n1193) );
INV_X1 U904 ( .A(n1195), .ZN(n1198) );
XOR2_X1 U905 ( .A(n1199), .B(n1200), .Z(n1195) );
XOR2_X1 U906 ( .A(G134), .B(n1201), .Z(n1200) );
XOR2_X1 U907 ( .A(KEYINPUT9), .B(G143), .Z(n1201) );
XOR2_X1 U908 ( .A(n1202), .B(n1203), .Z(n1199) );
NOR2_X1 U909 ( .A1(G128), .A2(KEYINPUT31), .ZN(n1203) );
NAND2_X1 U910 ( .A1(n1204), .A2(n1205), .ZN(n1202) );
OR2_X1 U911 ( .A1(n1206), .A2(G107), .ZN(n1205) );
XOR2_X1 U912 ( .A(n1207), .B(KEYINPUT60), .Z(n1204) );
NAND2_X1 U913 ( .A1(G107), .A2(n1206), .ZN(n1207) );
NAND3_X1 U914 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1206) );
NAND2_X1 U915 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
OR3_X1 U916 ( .A1(n1212), .A2(n1211), .A3(n1181), .ZN(n1209) );
INV_X1 U917 ( .A(KEYINPUT32), .ZN(n1212) );
NAND2_X1 U918 ( .A1(n1213), .A2(n1181), .ZN(n1208) );
NAND2_X1 U919 ( .A1(n1214), .A2(KEYINPUT32), .ZN(n1213) );
XNOR2_X1 U920 ( .A(n1211), .B(KEYINPUT41), .ZN(n1214) );
XNOR2_X1 U921 ( .A(n1170), .B(KEYINPUT29), .ZN(n1211) );
INV_X1 U922 ( .A(G122), .ZN(n1170) );
XNOR2_X1 U923 ( .A(n1025), .B(KEYINPUT44), .ZN(n1185) );
XNOR2_X1 U924 ( .A(n1215), .B(G475), .ZN(n1025) );
NAND2_X1 U925 ( .A1(n1078), .A2(n1216), .ZN(n1215) );
XOR2_X1 U926 ( .A(n1217), .B(n1218), .Z(n1078) );
NOR2_X1 U927 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
XOR2_X1 U928 ( .A(n1221), .B(KEYINPUT24), .Z(n1220) );
NAND2_X1 U929 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
XOR2_X1 U930 ( .A(n1082), .B(KEYINPUT12), .Z(n1222) );
INV_X1 U931 ( .A(G104), .ZN(n1082) );
NOR2_X1 U932 ( .A1(G104), .A2(n1223), .ZN(n1219) );
XOR2_X1 U933 ( .A(n1224), .B(G122), .Z(n1223) );
NAND2_X1 U934 ( .A1(KEYINPUT35), .A2(n1225), .ZN(n1224) );
XOR2_X1 U935 ( .A(KEYINPUT1), .B(n1226), .Z(n1225) );
NAND2_X1 U936 ( .A1(KEYINPUT22), .A2(n1227), .ZN(n1217) );
XOR2_X1 U937 ( .A(n1228), .B(n1229), .Z(n1227) );
XOR2_X1 U938 ( .A(n1230), .B(n1231), .Z(n1229) );
NOR2_X1 U939 ( .A1(G143), .A2(KEYINPUT2), .ZN(n1231) );
AND3_X1 U940 ( .A1(G214), .A2(n1006), .A3(n1232), .ZN(n1230) );
XOR2_X1 U941 ( .A(G131), .B(n1233), .Z(n1228) );
NOR2_X1 U942 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U943 ( .A(n1236), .B(KEYINPUT39), .Z(n1235) );
NAND2_X1 U944 ( .A1(n1237), .A2(n1147), .ZN(n1236) );
NOR2_X1 U945 ( .A1(n1238), .A2(n1237), .ZN(n1234) );
XNOR2_X1 U946 ( .A(n1239), .B(n1240), .ZN(n1237) );
XOR2_X1 U947 ( .A(KEYINPUT16), .B(G140), .Z(n1240) );
NAND2_X1 U948 ( .A1(KEYINPUT14), .A2(n1037), .ZN(n1239) );
XOR2_X1 U949 ( .A(n1147), .B(KEYINPUT56), .Z(n1238) );
AND3_X1 U950 ( .A1(n1018), .A2(n1184), .A3(n1014), .ZN(n973) );
NOR2_X1 U951 ( .A1(n995), .A2(n996), .ZN(n1014) );
AND2_X1 U952 ( .A1(G221), .A2(n1241), .ZN(n996) );
XOR2_X1 U953 ( .A(n1242), .B(G469), .Z(n995) );
NAND2_X1 U954 ( .A1(n1243), .A2(n1216), .ZN(n1242) );
XNOR2_X1 U955 ( .A(n1104), .B(n1244), .ZN(n1243) );
NOR2_X1 U956 ( .A1(n1109), .A2(n1245), .ZN(n1244) );
AND2_X1 U957 ( .A1(n1046), .A2(n1107), .ZN(n1245) );
NOR3_X1 U958 ( .A1(n1107), .A2(G953), .A3(n1046), .ZN(n1109) );
INV_X1 U959 ( .A(G227), .ZN(n1046) );
XNOR2_X1 U960 ( .A(n1246), .B(n1060), .ZN(n1104) );
NAND2_X1 U961 ( .A1(n1004), .A2(n1247), .ZN(n1184) );
NAND4_X1 U962 ( .A1(n1061), .A2(G902), .A3(n1169), .A4(n1062), .ZN(n1247) );
INV_X1 U963 ( .A(G898), .ZN(n1062) );
XOR2_X1 U964 ( .A(n1006), .B(KEYINPUT10), .Z(n1061) );
NAND3_X1 U965 ( .A1(n1169), .A2(n1006), .A3(G952), .ZN(n1004) );
NAND2_X1 U966 ( .A1(G237), .A2(G234), .ZN(n1169) );
AND2_X1 U967 ( .A1(n1248), .A2(n1000), .ZN(n1018) );
XNOR2_X1 U968 ( .A(n1021), .B(KEYINPUT53), .ZN(n1000) );
XOR2_X1 U969 ( .A(n1249), .B(n1113), .Z(n1021) );
AND2_X1 U970 ( .A1(G210), .A2(n1250), .ZN(n1113) );
NAND2_X1 U971 ( .A1(n1251), .A2(n1216), .ZN(n1249) );
XNOR2_X1 U972 ( .A(n1142), .B(n1146), .ZN(n1251) );
XNOR2_X1 U973 ( .A(n1252), .B(n1253), .ZN(n1146) );
INV_X1 U974 ( .A(n1254), .ZN(n1253) );
XNOR2_X1 U975 ( .A(n1255), .B(n1037), .ZN(n1252) );
NAND2_X1 U976 ( .A1(G224), .A2(n1006), .ZN(n1255) );
XNOR2_X1 U977 ( .A(n1060), .B(n1256), .ZN(n1142) );
XNOR2_X1 U978 ( .A(n1257), .B(n1058), .ZN(n1256) );
XOR2_X1 U979 ( .A(G110), .B(G122), .Z(n1058) );
NAND2_X1 U980 ( .A1(KEYINPUT58), .A2(n1059), .ZN(n1257) );
XNOR2_X1 U981 ( .A(n1167), .B(n1258), .ZN(n1060) );
XOR2_X1 U982 ( .A(G107), .B(G104), .Z(n1258) );
XOR2_X1 U983 ( .A(KEYINPUT25), .B(n1163), .Z(n1248) );
INV_X1 U984 ( .A(n999), .ZN(n1163) );
NAND2_X1 U985 ( .A1(G214), .A2(n1250), .ZN(n999) );
NAND2_X1 U986 ( .A1(n1232), .A2(n1216), .ZN(n1250) );
AND2_X1 U987 ( .A1(n1190), .A2(n1175), .ZN(n992) );
XOR2_X1 U988 ( .A(n1259), .B(n1068), .Z(n1175) );
NAND2_X1 U989 ( .A1(G217), .A2(n1241), .ZN(n1068) );
NAND2_X1 U990 ( .A1(G234), .A2(n1216), .ZN(n1241) );
OR2_X1 U991 ( .A1(n1067), .A2(G902), .ZN(n1259) );
XNOR2_X1 U992 ( .A(n1260), .B(n1261), .ZN(n1067) );
XOR2_X1 U993 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U994 ( .A(G137), .B(G119), .Z(n1263) );
XOR2_X1 U995 ( .A(KEYINPUT8), .B(KEYINPUT54), .Z(n1262) );
XOR2_X1 U996 ( .A(n1264), .B(n1265), .Z(n1260) );
XOR2_X1 U997 ( .A(n1266), .B(n1107), .Z(n1265) );
XOR2_X1 U998 ( .A(G110), .B(G140), .Z(n1107) );
XNOR2_X1 U999 ( .A(n1267), .B(n1037), .ZN(n1264) );
XNOR2_X1 U1000 ( .A(G125), .B(KEYINPUT34), .ZN(n1037) );
NAND2_X1 U1001 ( .A1(n1197), .A2(G221), .ZN(n1267) );
AND2_X1 U1002 ( .A1(G234), .A2(n1006), .ZN(n1197) );
XOR2_X1 U1003 ( .A(n1268), .B(G472), .Z(n1190) );
NAND2_X1 U1004 ( .A1(n1269), .A2(n1216), .ZN(n1268) );
INV_X1 U1005 ( .A(G902), .ZN(n1216) );
XOR2_X1 U1006 ( .A(n1270), .B(n1093), .Z(n1269) );
XNOR2_X1 U1007 ( .A(n1246), .B(n1059), .ZN(n1093) );
XOR2_X1 U1008 ( .A(n1271), .B(n1272), .Z(n1059) );
XOR2_X1 U1009 ( .A(KEYINPUT59), .B(G119), .Z(n1272) );
XOR2_X1 U1010 ( .A(n1181), .B(n1226), .Z(n1271) );
XOR2_X1 U1011 ( .A(G113), .B(KEYINPUT21), .Z(n1226) );
INV_X1 U1012 ( .A(G116), .ZN(n1181) );
XOR2_X1 U1013 ( .A(n1162), .B(n1034), .Z(n1246) );
XNOR2_X1 U1014 ( .A(n1254), .B(n1273), .ZN(n1034) );
XOR2_X1 U1015 ( .A(G137), .B(G134), .Z(n1273) );
XOR2_X1 U1016 ( .A(n1154), .B(n1266), .Z(n1254) );
XNOR2_X1 U1017 ( .A(G128), .B(n1147), .ZN(n1266) );
INV_X1 U1018 ( .A(G146), .ZN(n1147) );
INV_X1 U1019 ( .A(G143), .ZN(n1154) );
INV_X1 U1020 ( .A(G131), .ZN(n1162) );
NAND2_X1 U1021 ( .A1(KEYINPUT7), .A2(n1091), .ZN(n1270) );
AND2_X1 U1022 ( .A1(n1274), .A2(n1275), .ZN(n1091) );
NAND2_X1 U1023 ( .A1(n1276), .A2(n1167), .ZN(n1275) );
INV_X1 U1024 ( .A(G101), .ZN(n1167) );
NAND3_X1 U1025 ( .A1(n1232), .A2(n1006), .A3(G210), .ZN(n1276) );
NAND4_X1 U1026 ( .A1(n1232), .A2(n1006), .A3(G210), .A4(G101), .ZN(n1274) );
INV_X1 U1027 ( .A(G953), .ZN(n1006) );
INV_X1 U1028 ( .A(G237), .ZN(n1232) );
endmodule


