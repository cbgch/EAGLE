//Key = 0011110000101001110111001000001111101110010010110001000111100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284;

NOR4_X2 U704 ( .A1(n988), .A2(n1012), .A3(n1200), .A4(n1201), .ZN(n1086) );
XNOR2_X1 U705 ( .A(G107), .B(n973), .ZN(G9) );
NOR2_X1 U706 ( .A1(n974), .A2(n975), .ZN(G75) );
NOR4_X1 U707 ( .A1(n976), .A2(n977), .A3(G953), .A4(n978), .ZN(n975) );
NOR2_X1 U708 ( .A1(n979), .A2(n980), .ZN(n977) );
NOR2_X1 U709 ( .A1(n981), .A2(n982), .ZN(n979) );
NOR3_X1 U710 ( .A1(n983), .A2(n984), .A3(n985), .ZN(n982) );
NOR2_X1 U711 ( .A1(n986), .A2(n987), .ZN(n984) );
NOR2_X1 U712 ( .A1(n988), .A2(n989), .ZN(n987) );
NOR3_X1 U713 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n986) );
NOR3_X1 U714 ( .A1(n993), .A2(n994), .A3(n995), .ZN(n992) );
NOR2_X1 U715 ( .A1(n996), .A2(n997), .ZN(n991) );
NOR4_X1 U716 ( .A1(n993), .A2(n998), .A3(n989), .A4(n990), .ZN(n981) );
NOR2_X1 U717 ( .A1(n999), .A2(n1000), .ZN(n998) );
NOR2_X1 U718 ( .A1(n1001), .A2(n983), .ZN(n1000) );
NOR3_X1 U719 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(n1001) );
AND2_X1 U720 ( .A1(n1005), .A2(KEYINPUT53), .ZN(n1004) );
XNOR2_X1 U721 ( .A(KEYINPUT22), .B(n1006), .ZN(n1002) );
NOR3_X1 U722 ( .A1(n985), .A2(n1007), .A3(n1008), .ZN(n999) );
NOR2_X1 U723 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NOR2_X1 U724 ( .A1(KEYINPUT53), .A2(n1011), .ZN(n1009) );
NOR2_X1 U725 ( .A1(n1012), .A2(n1011), .ZN(n1007) );
INV_X1 U726 ( .A(n1005), .ZN(n985) );
NAND3_X1 U727 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n976) );
XNOR2_X1 U728 ( .A(n1016), .B(KEYINPUT41), .ZN(n1015) );
NOR3_X1 U729 ( .A1(n978), .A2(G953), .A3(G952), .ZN(n974) );
AND4_X1 U730 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n978) );
NOR4_X1 U731 ( .A1(n993), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1020) );
XOR2_X1 U732 ( .A(n1024), .B(G472), .Z(n1019) );
XOR2_X1 U733 ( .A(n1025), .B(KEYINPUT7), .Z(n1017) );
XOR2_X1 U734 ( .A(n1026), .B(n1027), .Z(G72) );
NOR2_X1 U735 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR2_X1 U736 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
XNOR2_X1 U737 ( .A(G227), .B(KEYINPUT1), .ZN(n1030) );
NAND2_X1 U738 ( .A1(n1032), .A2(n1033), .ZN(n1026) );
OR2_X1 U739 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
XOR2_X1 U740 ( .A(n1036), .B(KEYINPUT23), .Z(n1032) );
NAND2_X1 U741 ( .A1(n1037), .A2(n1035), .ZN(n1036) );
NOR2_X1 U742 ( .A1(G953), .A2(n1016), .ZN(n1035) );
XOR2_X1 U743 ( .A(n1034), .B(KEYINPUT27), .Z(n1037) );
NAND2_X1 U744 ( .A1(n1038), .A2(n1039), .ZN(n1034) );
NAND2_X1 U745 ( .A1(G953), .A2(n1031), .ZN(n1039) );
XOR2_X1 U746 ( .A(n1040), .B(n1041), .Z(n1038) );
XOR2_X1 U747 ( .A(n1042), .B(n1043), .Z(n1041) );
NAND2_X1 U748 ( .A1(KEYINPUT4), .A2(n1044), .ZN(n1042) );
XOR2_X1 U749 ( .A(n1045), .B(n1046), .Z(n1040) );
NOR2_X1 U750 ( .A1(G131), .A2(KEYINPUT6), .ZN(n1046) );
NOR2_X1 U751 ( .A1(KEYINPUT54), .A2(n1047), .ZN(n1045) );
XOR2_X1 U752 ( .A(G140), .B(n1048), .Z(n1047) );
NAND2_X1 U753 ( .A1(n1049), .A2(n1050), .ZN(G69) );
NAND2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U755 ( .A(n1053), .B(n1054), .Z(n1049) );
NOR2_X1 U756 ( .A1(n1052), .A2(n1055), .ZN(n1054) );
XOR2_X1 U757 ( .A(KEYINPUT26), .B(n1056), .Z(n1055) );
AND2_X1 U758 ( .A1(n1051), .A2(n1029), .ZN(n1056) );
NAND3_X1 U759 ( .A1(n1057), .A2(n1058), .A3(n1013), .ZN(n1051) );
NAND3_X1 U760 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1052) );
XOR2_X1 U761 ( .A(n1062), .B(KEYINPUT45), .Z(n1061) );
NAND2_X1 U762 ( .A1(G953), .A2(n1063), .ZN(n1062) );
NAND2_X1 U763 ( .A1(n1064), .A2(n1065), .ZN(n1060) );
NAND2_X1 U764 ( .A1(n1066), .A2(n1067), .ZN(n1059) );
XOR2_X1 U765 ( .A(KEYINPUT19), .B(n1064), .Z(n1066) );
NAND2_X1 U766 ( .A1(G953), .A2(n1068), .ZN(n1053) );
NAND2_X1 U767 ( .A1(G898), .A2(G224), .ZN(n1068) );
NOR2_X1 U768 ( .A1(n1069), .A2(n1070), .ZN(G66) );
XNOR2_X1 U769 ( .A(n1071), .B(n1072), .ZN(n1070) );
NOR2_X1 U770 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U771 ( .A1(n1069), .A2(n1075), .ZN(G63) );
XOR2_X1 U772 ( .A(n1076), .B(n1077), .Z(n1075) );
NOR3_X1 U773 ( .A1(n1074), .A2(KEYINPUT13), .A3(n1078), .ZN(n1076) );
INV_X1 U774 ( .A(G478), .ZN(n1078) );
NOR2_X1 U775 ( .A1(n1069), .A2(n1079), .ZN(G60) );
XOR2_X1 U776 ( .A(n1080), .B(n1081), .Z(n1079) );
XOR2_X1 U777 ( .A(KEYINPUT36), .B(n1082), .Z(n1081) );
AND2_X1 U778 ( .A1(G475), .A2(n1083), .ZN(n1082) );
XNOR2_X1 U779 ( .A(G104), .B(n1084), .ZN(G6) );
NAND4_X1 U780 ( .A1(n1085), .A2(KEYINPUT58), .A3(n1086), .A4(n1005), .ZN(n1084) );
XOR2_X1 U781 ( .A(n1087), .B(KEYINPUT21), .Z(n1085) );
NOR2_X1 U782 ( .A1(n1069), .A2(n1088), .ZN(G57) );
XOR2_X1 U783 ( .A(n1089), .B(n1090), .Z(n1088) );
XOR2_X1 U784 ( .A(KEYINPUT25), .B(n1091), .Z(n1090) );
NOR2_X1 U785 ( .A1(KEYINPUT50), .A2(n1092), .ZN(n1091) );
NOR2_X1 U786 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U787 ( .A(KEYINPUT14), .B(n1095), .Z(n1094) );
AND2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U789 ( .A1(n1097), .A2(n1096), .ZN(n1093) );
XOR2_X1 U790 ( .A(n1098), .B(n1099), .Z(n1089) );
NAND3_X1 U791 ( .A1(n1083), .A2(G472), .A3(KEYINPUT17), .ZN(n1098) );
NOR2_X1 U792 ( .A1(n1100), .A2(n1101), .ZN(G54) );
XOR2_X1 U793 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U794 ( .A(KEYINPUT55), .B(n1104), .Z(n1103) );
NOR2_X1 U795 ( .A1(KEYINPUT28), .A2(n1105), .ZN(n1104) );
XOR2_X1 U796 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U797 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND3_X1 U798 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND2_X1 U800 ( .A1(n1115), .A2(n1116), .ZN(n1111) );
INV_X1 U801 ( .A(KEYINPUT15), .ZN(n1116) );
NAND2_X1 U802 ( .A1(n1117), .A2(n1118), .ZN(n1115) );
XOR2_X1 U803 ( .A(KEYINPUT34), .B(n1113), .Z(n1117) );
NAND2_X1 U804 ( .A1(KEYINPUT15), .A2(n1119), .ZN(n1110) );
NAND2_X1 U805 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
OR2_X1 U806 ( .A1(n1122), .A2(KEYINPUT34), .ZN(n1121) );
NAND3_X1 U807 ( .A1(n1118), .A2(n1122), .A3(KEYINPUT34), .ZN(n1120) );
INV_X1 U808 ( .A(n1114), .ZN(n1118) );
NOR2_X1 U809 ( .A1(n1074), .A2(n1123), .ZN(n1102) );
XOR2_X1 U810 ( .A(KEYINPUT37), .B(G469), .Z(n1123) );
NOR2_X1 U811 ( .A1(G952), .A2(n1124), .ZN(n1100) );
XOR2_X1 U812 ( .A(n1029), .B(KEYINPUT60), .Z(n1124) );
NOR3_X1 U813 ( .A1(n1069), .A2(n1125), .A3(n1126), .ZN(G51) );
NOR3_X1 U814 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1126) );
INV_X1 U815 ( .A(n1130), .ZN(n1127) );
NOR2_X1 U816 ( .A1(n1131), .A2(n1130), .ZN(n1125) );
NAND2_X1 U817 ( .A1(n1083), .A2(n1132), .ZN(n1130) );
INV_X1 U818 ( .A(n1074), .ZN(n1083) );
NAND2_X1 U819 ( .A1(G902), .A2(n1133), .ZN(n1074) );
NAND3_X1 U820 ( .A1(n1014), .A2(n1016), .A3(n1013), .ZN(n1133) );
AND2_X1 U821 ( .A1(n973), .A2(n1134), .ZN(n1013) );
NAND3_X1 U822 ( .A1(n1086), .A2(n1135), .A3(n996), .ZN(n1134) );
NAND2_X1 U823 ( .A1(n1006), .A2(n1136), .ZN(n1135) );
NAND3_X1 U824 ( .A1(n994), .A2(n1005), .A3(n1086), .ZN(n973) );
AND4_X1 U825 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1016) );
NOR4_X1 U826 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1140) );
AND2_X1 U827 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NOR3_X1 U828 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1143) );
XNOR2_X1 U829 ( .A(KEYINPUT5), .B(n1136), .ZN(n1147) );
INV_X1 U830 ( .A(n1150), .ZN(n1142) );
INV_X1 U831 ( .A(n1151), .ZN(n1141) );
AND2_X1 U832 ( .A1(n1152), .A2(n1153), .ZN(n1139) );
NAND3_X1 U833 ( .A1(n1154), .A2(n994), .A3(n1155), .ZN(n1138) );
XNOR2_X1 U834 ( .A(n1156), .B(KEYINPUT12), .ZN(n1155) );
AND2_X1 U835 ( .A1(n1157), .A2(n1058), .ZN(n1014) );
NAND3_X1 U836 ( .A1(n1086), .A2(n1005), .A3(n995), .ZN(n1058) );
XOR2_X1 U837 ( .A(KEYINPUT29), .B(n1057), .Z(n1157) );
AND4_X1 U838 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1057) );
NOR2_X1 U839 ( .A1(n1128), .A2(n1129), .ZN(n1131) );
XNOR2_X1 U840 ( .A(n1162), .B(KEYINPUT62), .ZN(n1129) );
NAND2_X1 U841 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U842 ( .A1(n1164), .A2(n1163), .ZN(n1128) );
NAND2_X1 U843 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NOR2_X1 U844 ( .A1(n1029), .A2(G952), .ZN(n1069) );
XOR2_X1 U845 ( .A(n1167), .B(n1150), .Z(G48) );
NAND3_X1 U846 ( .A1(n1156), .A2(n995), .A3(n1154), .ZN(n1150) );
XOR2_X1 U847 ( .A(n1168), .B(n1151), .Z(G45) );
NAND4_X1 U848 ( .A1(n1154), .A2(n1003), .A3(n1021), .A4(n1023), .ZN(n1151) );
AND2_X1 U849 ( .A1(n1169), .A2(n1170), .ZN(n1154) );
XNOR2_X1 U850 ( .A(G140), .B(n1171), .ZN(G42) );
NAND4_X1 U851 ( .A1(n1145), .A2(n1018), .A3(n1172), .A4(n1173), .ZN(n1171) );
XOR2_X1 U852 ( .A(KEYINPUT42), .B(n1170), .Z(n1172) );
XOR2_X1 U853 ( .A(n1153), .B(n1174), .Z(G39) );
NAND2_X1 U854 ( .A1(KEYINPUT33), .A2(G137), .ZN(n1174) );
NAND3_X1 U855 ( .A1(n1156), .A2(n996), .A3(n1146), .ZN(n1153) );
XOR2_X1 U856 ( .A(n1175), .B(n1176), .Z(G36) );
AND2_X1 U857 ( .A1(n1177), .A2(n1146), .ZN(n1176) );
NOR2_X1 U858 ( .A1(KEYINPUT49), .A2(n1178), .ZN(n1175) );
NAND2_X1 U859 ( .A1(n1179), .A2(n1180), .ZN(G33) );
NAND2_X1 U860 ( .A1(G131), .A2(n1152), .ZN(n1180) );
XOR2_X1 U861 ( .A(KEYINPUT38), .B(n1181), .Z(n1179) );
NOR2_X1 U862 ( .A1(G131), .A2(n1152), .ZN(n1181) );
NAND3_X1 U863 ( .A1(n995), .A2(n1003), .A3(n1146), .ZN(n1152) );
INV_X1 U864 ( .A(n1149), .ZN(n1146) );
NAND3_X1 U865 ( .A1(n1170), .A2(n1173), .A3(n1018), .ZN(n1149) );
INV_X1 U866 ( .A(n983), .ZN(n1018) );
NAND2_X1 U867 ( .A1(n1012), .A2(n1011), .ZN(n983) );
XOR2_X1 U868 ( .A(n1182), .B(n1183), .Z(G30) );
NAND4_X1 U869 ( .A1(n1169), .A2(n1156), .A3(n994), .A4(n1184), .ZN(n1183) );
XOR2_X1 U870 ( .A(KEYINPUT35), .B(n1170), .Z(n1184) );
INV_X1 U871 ( .A(n988), .ZN(n1170) );
INV_X1 U872 ( .A(n1148), .ZN(n994) );
NAND2_X1 U873 ( .A1(n1185), .A2(n1186), .ZN(G3) );
NAND2_X1 U874 ( .A1(G101), .A2(n1187), .ZN(n1186) );
XOR2_X1 U875 ( .A(KEYINPUT32), .B(n1188), .Z(n1185) );
NOR2_X1 U876 ( .A1(G101), .A2(n1187), .ZN(n1188) );
NAND3_X1 U877 ( .A1(n1086), .A2(n1003), .A3(n996), .ZN(n1187) );
XOR2_X1 U878 ( .A(n1048), .B(n1137), .Z(G27) );
NAND4_X1 U879 ( .A1(n1145), .A2(n1169), .A3(n1025), .A4(n997), .ZN(n1137) );
AND3_X1 U880 ( .A1(n1173), .A2(n1011), .A3(n1010), .ZN(n1169) );
NAND2_X1 U881 ( .A1(n980), .A2(n1189), .ZN(n1173) );
NAND4_X1 U882 ( .A1(G902), .A2(G953), .A3(n1190), .A4(n1031), .ZN(n1189) );
INV_X1 U883 ( .A(G900), .ZN(n1031) );
NOR2_X1 U884 ( .A1(n1006), .A2(n1087), .ZN(n1145) );
XOR2_X1 U885 ( .A(n1191), .B(n1158), .Z(G24) );
NAND4_X1 U886 ( .A1(n1192), .A2(n1005), .A3(n1021), .A4(n1023), .ZN(n1158) );
NAND2_X1 U887 ( .A1(n1193), .A2(n1194), .ZN(n1005) );
OR2_X1 U888 ( .A1(n1136), .A2(KEYINPUT47), .ZN(n1194) );
NAND3_X1 U889 ( .A1(n1195), .A2(n1196), .A3(KEYINPUT47), .ZN(n1193) );
XOR2_X1 U890 ( .A(n1159), .B(n1197), .Z(G21) );
XNOR2_X1 U891 ( .A(G119), .B(KEYINPUT61), .ZN(n1197) );
NAND3_X1 U892 ( .A1(n1192), .A2(n996), .A3(n1156), .ZN(n1159) );
NOR2_X1 U893 ( .A1(n1195), .A2(n1196), .ZN(n1156) );
INV_X1 U894 ( .A(n989), .ZN(n996) );
XNOR2_X1 U895 ( .A(G116), .B(n1160), .ZN(G18) );
NAND2_X1 U896 ( .A1(n1177), .A2(n1192), .ZN(n1160) );
NOR2_X1 U897 ( .A1(n1148), .A2(n1136), .ZN(n1177) );
INV_X1 U898 ( .A(n1003), .ZN(n1136) );
NAND2_X1 U899 ( .A1(n1198), .A2(n1023), .ZN(n1148) );
XNOR2_X1 U900 ( .A(G113), .B(n1161), .ZN(G15) );
NAND3_X1 U901 ( .A1(n995), .A2(n1003), .A3(n1192), .ZN(n1161) );
AND3_X1 U902 ( .A1(n1025), .A2(n1010), .A3(n1199), .ZN(n1192) );
NOR3_X1 U903 ( .A1(n1200), .A2(n993), .A3(n1201), .ZN(n1199) );
INV_X1 U904 ( .A(n997), .ZN(n993) );
INV_X1 U905 ( .A(n1012), .ZN(n1010) );
NOR2_X1 U906 ( .A1(n1195), .A2(n1022), .ZN(n1003) );
INV_X1 U907 ( .A(n1087), .ZN(n995) );
NAND2_X1 U908 ( .A1(n1202), .A2(n1021), .ZN(n1087) );
XOR2_X1 U909 ( .A(G110), .B(n1203), .Z(G12) );
NOR4_X1 U910 ( .A1(KEYINPUT11), .A2(n1204), .A3(n989), .A4(n1006), .ZN(n1203) );
NAND2_X1 U911 ( .A1(n1205), .A2(n1022), .ZN(n1006) );
INV_X1 U912 ( .A(n1196), .ZN(n1022) );
XNOR2_X1 U913 ( .A(n1206), .B(n1073), .ZN(n1196) );
NAND2_X1 U914 ( .A1(G217), .A2(n1207), .ZN(n1073) );
NAND2_X1 U915 ( .A1(n1071), .A2(n1208), .ZN(n1206) );
XNOR2_X1 U916 ( .A(n1209), .B(n1210), .ZN(n1071) );
XOR2_X1 U917 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U918 ( .A(G128), .B(G125), .Z(n1212) );
XOR2_X1 U919 ( .A(G146), .B(G137), .Z(n1211) );
XNOR2_X1 U920 ( .A(n1213), .B(n1106), .ZN(n1209) );
XOR2_X1 U921 ( .A(n1214), .B(G119), .Z(n1213) );
NAND2_X1 U922 ( .A1(n1215), .A2(G221), .ZN(n1214) );
XNOR2_X1 U923 ( .A(KEYINPUT47), .B(n1195), .ZN(n1205) );
XNOR2_X1 U924 ( .A(n1216), .B(n1217), .ZN(n1195) );
XNOR2_X1 U925 ( .A(KEYINPUT44), .B(n1024), .ZN(n1217) );
NAND2_X1 U926 ( .A1(n1218), .A2(n1208), .ZN(n1024) );
XOR2_X1 U927 ( .A(n1219), .B(n1220), .Z(n1218) );
XNOR2_X1 U928 ( .A(n1099), .B(n1221), .ZN(n1220) );
NOR2_X1 U929 ( .A1(KEYINPUT18), .A2(n1096), .ZN(n1221) );
NAND2_X1 U930 ( .A1(n1222), .A2(G210), .ZN(n1096) );
XOR2_X1 U931 ( .A(n1223), .B(n1224), .Z(n1099) );
XOR2_X1 U932 ( .A(n1225), .B(n1113), .Z(n1224) );
NAND2_X1 U933 ( .A1(KEYINPUT20), .A2(G472), .ZN(n1216) );
NAND2_X1 U934 ( .A1(n1198), .A2(n1202), .ZN(n989) );
XOR2_X1 U935 ( .A(n1023), .B(KEYINPUT31), .Z(n1202) );
XNOR2_X1 U936 ( .A(n1226), .B(G478), .ZN(n1023) );
OR2_X1 U937 ( .A1(n1077), .A2(G902), .ZN(n1226) );
XNOR2_X1 U938 ( .A(n1227), .B(n1228), .ZN(n1077) );
XOR2_X1 U939 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U940 ( .A(G128), .B(G122), .Z(n1230) );
XOR2_X1 U941 ( .A(G143), .B(G134), .Z(n1229) );
XOR2_X1 U942 ( .A(n1231), .B(n1232), .Z(n1227) );
XOR2_X1 U943 ( .A(G107), .B(n1233), .Z(n1232) );
NOR2_X1 U944 ( .A1(KEYINPUT9), .A2(n1234), .ZN(n1233) );
XNOR2_X1 U945 ( .A(G116), .B(KEYINPUT56), .ZN(n1234) );
NAND2_X1 U946 ( .A1(G217), .A2(n1215), .ZN(n1231) );
AND2_X1 U947 ( .A1(n1235), .A2(G234), .ZN(n1215) );
INV_X1 U948 ( .A(n1021), .ZN(n1198) );
XNOR2_X1 U949 ( .A(n1236), .B(G475), .ZN(n1021) );
NAND2_X1 U950 ( .A1(n1237), .A2(n1208), .ZN(n1236) );
XNOR2_X1 U951 ( .A(n1080), .B(KEYINPUT2), .ZN(n1237) );
XNOR2_X1 U952 ( .A(n1238), .B(n1239), .ZN(n1080) );
XOR2_X1 U953 ( .A(n1240), .B(n1241), .Z(n1239) );
XNOR2_X1 U954 ( .A(n1242), .B(n1243), .ZN(n1241) );
NAND2_X1 U955 ( .A1(n1222), .A2(G214), .ZN(n1242) );
NOR2_X1 U956 ( .A1(n1244), .A2(G237), .ZN(n1222) );
INV_X1 U957 ( .A(n1235), .ZN(n1244) );
XOR2_X1 U958 ( .A(n1245), .B(n1246), .Z(n1240) );
NAND2_X1 U959 ( .A1(KEYINPUT57), .A2(G113), .ZN(n1246) );
NAND3_X1 U960 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(n1245) );
NAND2_X1 U961 ( .A1(G140), .A2(n1250), .ZN(n1249) );
OR3_X1 U962 ( .A1(n1250), .A2(G140), .A3(KEYINPUT8), .ZN(n1248) );
OR2_X1 U963 ( .A1(KEYINPUT0), .A2(n1251), .ZN(n1250) );
NAND2_X1 U964 ( .A1(KEYINPUT8), .A2(n1251), .ZN(n1247) );
XOR2_X1 U965 ( .A(n1048), .B(KEYINPUT24), .Z(n1251) );
XOR2_X1 U966 ( .A(n1252), .B(n1253), .Z(n1238) );
XOR2_X1 U967 ( .A(KEYINPUT39), .B(G131), .Z(n1253) );
XOR2_X1 U968 ( .A(G104), .B(n1191), .Z(n1252) );
INV_X1 U969 ( .A(G122), .ZN(n1191) );
INV_X1 U970 ( .A(n1086), .ZN(n1204) );
AND2_X1 U971 ( .A1(n980), .A2(n1254), .ZN(n1201) );
NAND4_X1 U972 ( .A1(G902), .A2(G953), .A3(n1190), .A4(n1063), .ZN(n1254) );
INV_X1 U973 ( .A(G898), .ZN(n1063) );
NAND3_X1 U974 ( .A1(n1190), .A2(n1029), .A3(G952), .ZN(n980) );
NAND2_X1 U975 ( .A1(G237), .A2(G234), .ZN(n1190) );
INV_X1 U976 ( .A(n1011), .ZN(n1200) );
NAND2_X1 U977 ( .A1(G214), .A2(n1255), .ZN(n1011) );
XOR2_X1 U978 ( .A(n1256), .B(n1132), .Z(n1012) );
AND2_X1 U979 ( .A1(G210), .A2(n1255), .ZN(n1132) );
NAND2_X1 U980 ( .A1(n1257), .A2(n1208), .ZN(n1255) );
INV_X1 U981 ( .A(G237), .ZN(n1257) );
NAND3_X1 U982 ( .A1(n1258), .A2(n1208), .A3(n1259), .ZN(n1256) );
NAND3_X1 U983 ( .A1(n1260), .A2(n1166), .A3(n1163), .ZN(n1259) );
NAND2_X1 U984 ( .A1(n1261), .A2(n1262), .ZN(n1258) );
NAND2_X1 U985 ( .A1(n1260), .A2(n1166), .ZN(n1262) );
NAND3_X1 U986 ( .A1(G224), .A2(n1263), .A3(n1264), .ZN(n1166) );
XOR2_X1 U987 ( .A(G125), .B(n1223), .Z(n1263) );
XNOR2_X1 U988 ( .A(n1165), .B(KEYINPUT3), .ZN(n1260) );
NAND2_X1 U989 ( .A1(n1265), .A2(n1266), .ZN(n1165) );
NAND2_X1 U990 ( .A1(n1264), .A2(G224), .ZN(n1266) );
XOR2_X1 U991 ( .A(KEYINPUT40), .B(n1235), .Z(n1264) );
XOR2_X1 U992 ( .A(n1048), .B(n1223), .Z(n1265) );
XOR2_X1 U993 ( .A(n1243), .B(n1267), .Z(n1223) );
INV_X1 U994 ( .A(n1268), .ZN(n1267) );
INV_X1 U995 ( .A(G125), .ZN(n1048) );
XOR2_X1 U996 ( .A(KEYINPUT46), .B(n1163), .Z(n1261) );
XOR2_X1 U997 ( .A(n1065), .B(n1064), .Z(n1163) );
XNOR2_X1 U998 ( .A(n1225), .B(n1269), .ZN(n1064) );
XOR2_X1 U999 ( .A(G122), .B(G110), .Z(n1269) );
XNOR2_X1 U1000 ( .A(G113), .B(n1270), .ZN(n1225) );
XOR2_X1 U1001 ( .A(G119), .B(G116), .Z(n1270) );
INV_X1 U1002 ( .A(n1067), .ZN(n1065) );
NAND2_X1 U1003 ( .A1(n1271), .A2(n1272), .ZN(n1067) );
OR2_X1 U1004 ( .A1(n1273), .A2(KEYINPUT48), .ZN(n1272) );
NAND3_X1 U1005 ( .A1(n1274), .A2(n1219), .A3(KEYINPUT48), .ZN(n1271) );
NAND2_X1 U1006 ( .A1(n990), .A2(n997), .ZN(n988) );
NAND2_X1 U1007 ( .A1(G221), .A2(n1207), .ZN(n997) );
NAND2_X1 U1008 ( .A1(G234), .A2(n1208), .ZN(n1207) );
INV_X1 U1009 ( .A(n1025), .ZN(n990) );
XOR2_X1 U1010 ( .A(n1275), .B(G469), .Z(n1025) );
NAND2_X1 U1011 ( .A1(n1276), .A2(n1208), .ZN(n1275) );
INV_X1 U1012 ( .A(G902), .ZN(n1208) );
XOR2_X1 U1013 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U1014 ( .A(n1113), .B(n1114), .Z(n1278) );
XOR2_X1 U1015 ( .A(n1044), .B(n1279), .Z(n1114) );
XOR2_X1 U1016 ( .A(KEYINPUT43), .B(n1273), .Z(n1279) );
XOR2_X1 U1017 ( .A(n1274), .B(n1097), .Z(n1273) );
INV_X1 U1018 ( .A(n1219), .ZN(n1097) );
XNOR2_X1 U1019 ( .A(G101), .B(KEYINPUT51), .ZN(n1219) );
XOR2_X1 U1020 ( .A(G104), .B(G107), .Z(n1274) );
XOR2_X1 U1021 ( .A(n1268), .B(n1280), .Z(n1044) );
NOR2_X1 U1022 ( .A1(KEYINPUT52), .A2(n1281), .ZN(n1280) );
XOR2_X1 U1023 ( .A(n1282), .B(n1243), .Z(n1281) );
XOR2_X1 U1024 ( .A(n1168), .B(n1167), .Z(n1243) );
INV_X1 U1025 ( .A(G146), .ZN(n1167) );
INV_X1 U1026 ( .A(G143), .ZN(n1168) );
XNOR2_X1 U1027 ( .A(KEYINPUT16), .B(KEYINPUT10), .ZN(n1282) );
XOR2_X1 U1028 ( .A(n1182), .B(KEYINPUT30), .Z(n1268) );
INV_X1 U1029 ( .A(G128), .ZN(n1182) );
INV_X1 U1030 ( .A(n1122), .ZN(n1113) );
XOR2_X1 U1031 ( .A(G131), .B(n1283), .Z(n1122) );
INV_X1 U1032 ( .A(n1043), .ZN(n1283) );
XOR2_X1 U1033 ( .A(n1178), .B(G137), .Z(n1043) );
INV_X1 U1034 ( .A(G134), .ZN(n1178) );
XNOR2_X1 U1035 ( .A(n1108), .B(n1284), .ZN(n1277) );
NOR2_X1 U1036 ( .A1(KEYINPUT59), .A2(n1106), .ZN(n1284) );
XNOR2_X1 U1037 ( .A(G110), .B(G140), .ZN(n1106) );
NAND2_X1 U1038 ( .A1(G227), .A2(n1235), .ZN(n1108) );
XOR2_X1 U1039 ( .A(n1029), .B(KEYINPUT63), .Z(n1235) );
INV_X1 U1040 ( .A(G953), .ZN(n1029) );
endmodule


