//Key = 1100010000000101110101110010111000011001111101011100110001110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304;

XNOR2_X1 U720 ( .A(G107), .B(n989), .ZN(G9) );
NOR2_X1 U721 ( .A1(n990), .A2(n991), .ZN(G75) );
NOR4_X1 U722 ( .A1(n992), .A2(n993), .A3(G953), .A4(n994), .ZN(n991) );
NOR3_X1 U723 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n993) );
NOR2_X1 U724 ( .A1(n998), .A2(n999), .ZN(n997) );
NOR2_X1 U725 ( .A1(n1000), .A2(n1001), .ZN(n998) );
NOR2_X1 U726 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NOR2_X1 U727 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NOR2_X1 U728 ( .A1(n1006), .A2(n1007), .ZN(n1002) );
NOR2_X1 U729 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
NOR2_X1 U730 ( .A1(n1010), .A2(n1011), .ZN(n996) );
NOR4_X1 U731 ( .A1(KEYINPUT35), .A2(n1012), .A3(n1005), .A4(n1007), .ZN(n1011) );
NAND3_X1 U732 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n992) );
NAND2_X1 U733 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NAND2_X1 U734 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND2_X1 U735 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
XOR2_X1 U736 ( .A(n1022), .B(KEYINPUT6), .Z(n1018) );
NAND4_X1 U737 ( .A1(n1023), .A2(n1010), .A3(n1024), .A4(n1025), .ZN(n1022) );
NOR2_X1 U738 ( .A1(n995), .A2(n1005), .ZN(n1024) );
INV_X1 U739 ( .A(n1026), .ZN(n995) );
INV_X1 U740 ( .A(n999), .ZN(n1010) );
NAND2_X1 U741 ( .A1(n1020), .A2(n1027), .ZN(n1013) );
NAND2_X1 U742 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U743 ( .A1(n1026), .A2(n1030), .ZN(n1029) );
NAND2_X1 U744 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U745 ( .A1(KEYINPUT35), .A2(n1033), .ZN(n1032) );
NAND2_X1 U746 ( .A1(n1034), .A2(n1035), .ZN(n1031) );
NAND2_X1 U747 ( .A1(n1036), .A2(n1037), .ZN(n1028) );
XOR2_X1 U748 ( .A(n1001), .B(KEYINPUT5), .Z(n1036) );
NOR3_X1 U749 ( .A1(n1007), .A2(n1005), .A3(n999), .ZN(n1020) );
INV_X1 U750 ( .A(n1038), .ZN(n1007) );
NOR3_X1 U751 ( .A1(n994), .A2(G953), .A3(G952), .ZN(n990) );
AND4_X1 U752 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n994) );
NOR4_X1 U753 ( .A1(n1034), .A2(n1023), .A3(n1043), .A4(n1044), .ZN(n1042) );
NOR2_X1 U754 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
XOR2_X1 U755 ( .A(KEYINPUT41), .B(G478), .Z(n1046) );
INV_X1 U756 ( .A(n1047), .ZN(n1043) );
NOR3_X1 U757 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1041) );
NOR2_X1 U758 ( .A1(n1021), .A2(n1051), .ZN(n1050) );
INV_X1 U759 ( .A(KEYINPUT62), .ZN(n1051) );
NOR2_X1 U760 ( .A1(KEYINPUT62), .A2(n1026), .ZN(n1049) );
XOR2_X1 U761 ( .A(KEYINPUT31), .B(n1052), .Z(n1048) );
XOR2_X1 U762 ( .A(n1053), .B(n1054), .Z(n1039) );
XOR2_X1 U763 ( .A(KEYINPUT8), .B(G469), .Z(n1054) );
XOR2_X1 U764 ( .A(n1055), .B(n1056), .Z(G72) );
XOR2_X1 U765 ( .A(n1057), .B(n1058), .Z(n1056) );
NAND2_X1 U766 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
INV_X1 U767 ( .A(n1061), .ZN(n1060) );
XOR2_X1 U768 ( .A(n1062), .B(n1063), .Z(n1059) );
NOR2_X1 U769 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
XOR2_X1 U770 ( .A(n1066), .B(KEYINPUT57), .Z(n1065) );
NAND2_X1 U771 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U772 ( .A1(n1067), .A2(n1068), .ZN(n1064) );
XNOR2_X1 U773 ( .A(G125), .B(G140), .ZN(n1062) );
NAND2_X1 U774 ( .A1(n1069), .A2(n1070), .ZN(n1057) );
NAND2_X1 U775 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR2_X1 U776 ( .A1(n1073), .A2(n1070), .ZN(n1055) );
AND2_X1 U777 ( .A1(G227), .A2(G900), .ZN(n1073) );
XOR2_X1 U778 ( .A(n1074), .B(n1075), .Z(G69) );
NOR2_X1 U779 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U780 ( .A(n1078), .B(KEYINPUT59), .Z(n1077) );
NAND2_X1 U781 ( .A1(G953), .A2(n1079), .ZN(n1078) );
NAND2_X1 U782 ( .A1(G898), .A2(G224), .ZN(n1079) );
NOR2_X1 U783 ( .A1(n1080), .A2(G953), .ZN(n1076) );
NOR2_X1 U784 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U785 ( .A1(n1083), .A2(n1084), .ZN(n1074) );
INV_X1 U786 ( .A(n1085), .ZN(n1084) );
NOR2_X1 U787 ( .A1(n1086), .A2(n1087), .ZN(G66) );
XOR2_X1 U788 ( .A(n1088), .B(n1089), .Z(n1087) );
XOR2_X1 U789 ( .A(n1090), .B(KEYINPUT16), .Z(n1088) );
NAND2_X1 U790 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR2_X1 U791 ( .A1(n1093), .A2(n1070), .ZN(n1086) );
XNOR2_X1 U792 ( .A(G952), .B(KEYINPUT52), .ZN(n1093) );
NOR2_X1 U793 ( .A1(n1094), .A2(n1095), .ZN(G63) );
XOR2_X1 U794 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U795 ( .A1(KEYINPUT26), .A2(n1098), .ZN(n1097) );
NAND2_X1 U796 ( .A1(n1091), .A2(G478), .ZN(n1096) );
NOR3_X1 U797 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(G60) );
AND3_X1 U798 ( .A1(KEYINPUT33), .A2(G953), .A3(G952), .ZN(n1101) );
NOR2_X1 U799 ( .A1(KEYINPUT33), .A2(n1102), .ZN(n1100) );
INV_X1 U800 ( .A(n1094), .ZN(n1102) );
XOR2_X1 U801 ( .A(n1103), .B(n1104), .Z(n1099) );
NAND2_X1 U802 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
OR2_X1 U803 ( .A1(KEYINPUT50), .A2(n1107), .ZN(n1106) );
NAND2_X1 U804 ( .A1(KEYINPUT44), .A2(n1107), .ZN(n1105) );
XOR2_X1 U805 ( .A(n1108), .B(KEYINPUT36), .Z(n1107) );
NAND2_X1 U806 ( .A1(n1091), .A2(G475), .ZN(n1103) );
XOR2_X1 U807 ( .A(n1109), .B(n1110), .Z(G6) );
XOR2_X1 U808 ( .A(n1111), .B(KEYINPUT51), .Z(n1110) );
NOR2_X1 U809 ( .A1(n1094), .A2(n1112), .ZN(G57) );
XOR2_X1 U810 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U811 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U812 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U813 ( .A1(n1091), .A2(G472), .ZN(n1117) );
XOR2_X1 U814 ( .A(n1119), .B(n1120), .Z(n1113) );
XOR2_X1 U815 ( .A(KEYINPUT30), .B(KEYINPUT1), .Z(n1120) );
NAND2_X1 U816 ( .A1(KEYINPUT48), .A2(n1121), .ZN(n1119) );
NOR2_X1 U817 ( .A1(n1094), .A2(n1122), .ZN(G54) );
XOR2_X1 U818 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U819 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U820 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR3_X1 U821 ( .A1(n1129), .A2(KEYINPUT7), .A3(G953), .ZN(n1128) );
INV_X1 U822 ( .A(G227), .ZN(n1129) );
NAND2_X1 U823 ( .A1(n1091), .A2(G469), .ZN(n1125) );
XOR2_X1 U824 ( .A(n1130), .B(n1131), .Z(n1123) );
XOR2_X1 U825 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U826 ( .A1(n1094), .A2(n1134), .ZN(G51) );
XOR2_X1 U827 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U828 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U829 ( .A1(n1091), .A2(n1139), .ZN(n1137) );
NOR2_X1 U830 ( .A1(n1140), .A2(n1015), .ZN(n1091) );
AND4_X1 U831 ( .A1(n1141), .A2(n1071), .A3(n1142), .A4(n1143), .ZN(n1015) );
XNOR2_X1 U832 ( .A(KEYINPUT12), .B(n1081), .ZN(n1143) );
NAND4_X1 U833 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1081) );
NAND2_X1 U834 ( .A1(n1148), .A2(n1149), .ZN(n1144) );
XNOR2_X1 U835 ( .A(KEYINPUT56), .B(n1150), .ZN(n1148) );
XOR2_X1 U836 ( .A(KEYINPUT11), .B(n1072), .Z(n1142) );
AND4_X1 U837 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1072) );
AND2_X1 U838 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
OR2_X1 U839 ( .A1(n1157), .A2(KEYINPUT24), .ZN(n1152) );
NAND3_X1 U840 ( .A1(n1158), .A2(n1159), .A3(KEYINPUT24), .ZN(n1151) );
AND4_X1 U841 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1071) );
AND2_X1 U842 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U843 ( .A1(n1166), .A2(n1016), .ZN(n1162) );
NAND2_X1 U844 ( .A1(n1167), .A2(n1168), .ZN(n1161) );
INV_X1 U845 ( .A(KEYINPUT25), .ZN(n1168) );
NAND4_X1 U846 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(KEYINPUT25), .ZN(n1160) );
INV_X1 U847 ( .A(n1082), .ZN(n1141) );
NAND4_X1 U848 ( .A1(n1109), .A2(n1172), .A3(n1173), .A4(n989), .ZN(n1082) );
NAND3_X1 U849 ( .A1(n1026), .A2(n1008), .A3(n1174), .ZN(n989) );
NAND3_X1 U850 ( .A1(n1174), .A2(n1026), .A3(n1009), .ZN(n1109) );
NOR2_X1 U851 ( .A1(n1070), .A2(G952), .ZN(n1094) );
XOR2_X1 U852 ( .A(n1175), .B(n1165), .Z(G48) );
NAND3_X1 U853 ( .A1(n1009), .A2(n1033), .A3(n1176), .ZN(n1165) );
XOR2_X1 U854 ( .A(G143), .B(n1167), .Z(G45) );
AND2_X1 U855 ( .A1(n1169), .A2(n1177), .ZN(n1167) );
AND4_X1 U856 ( .A1(n1178), .A2(n1037), .A3(n1033), .A4(n1179), .ZN(n1169) );
XNOR2_X1 U857 ( .A(G140), .B(n1164), .ZN(G42) );
NAND2_X1 U858 ( .A1(n1180), .A2(n1021), .ZN(n1164) );
XOR2_X1 U859 ( .A(G137), .B(n1181), .Z(G39) );
NOR2_X1 U860 ( .A1(n1001), .A2(n1182), .ZN(n1181) );
XOR2_X1 U861 ( .A(KEYINPUT49), .B(n1166), .Z(n1182) );
AND2_X1 U862 ( .A1(n1176), .A2(n1183), .ZN(n1166) );
INV_X1 U863 ( .A(n1016), .ZN(n1001) );
XNOR2_X1 U864 ( .A(G134), .B(n1153), .ZN(G36) );
NAND4_X1 U865 ( .A1(n1177), .A2(n1016), .A3(n1037), .A4(n1008), .ZN(n1153) );
XNOR2_X1 U866 ( .A(G131), .B(n1156), .ZN(G33) );
NAND2_X1 U867 ( .A1(n1180), .A2(n1037), .ZN(n1156) );
AND3_X1 U868 ( .A1(n1016), .A2(n1009), .A3(n1177), .ZN(n1180) );
NOR2_X1 U869 ( .A1(n1052), .A2(n1034), .ZN(n1016) );
INV_X1 U870 ( .A(n1035), .ZN(n1052) );
XOR2_X1 U871 ( .A(n1155), .B(n1184), .Z(G30) );
NOR2_X1 U872 ( .A1(G128), .A2(KEYINPUT2), .ZN(n1184) );
NAND3_X1 U873 ( .A1(n1008), .A2(n1033), .A3(n1176), .ZN(n1155) );
AND3_X1 U874 ( .A1(n1185), .A2(n1186), .A3(n1177), .ZN(n1176) );
NOR2_X1 U875 ( .A1(n1004), .A2(n1171), .ZN(n1177) );
INV_X1 U876 ( .A(n1187), .ZN(n1171) );
INV_X1 U877 ( .A(n1170), .ZN(n1004) );
XOR2_X1 U878 ( .A(n1121), .B(n1172), .Z(G3) );
NAND3_X1 U879 ( .A1(n1183), .A2(n1174), .A3(n1037), .ZN(n1172) );
XOR2_X1 U880 ( .A(n1157), .B(n1188), .Z(G27) );
NAND2_X1 U881 ( .A1(KEYINPUT39), .A2(G125), .ZN(n1188) );
NAND2_X1 U882 ( .A1(n1158), .A2(n1009), .ZN(n1157) );
AND4_X1 U883 ( .A1(n1038), .A2(n1021), .A3(n1033), .A4(n1187), .ZN(n1158) );
NAND2_X1 U884 ( .A1(n999), .A2(n1189), .ZN(n1187) );
NAND3_X1 U885 ( .A1(G902), .A2(n1190), .A3(n1061), .ZN(n1189) );
NOR2_X1 U886 ( .A1(n1070), .A2(G900), .ZN(n1061) );
XOR2_X1 U887 ( .A(n1191), .B(n1145), .Z(G24) );
NAND4_X1 U888 ( .A1(n1192), .A2(n1026), .A3(n1178), .A4(n1179), .ZN(n1145) );
NOR2_X1 U889 ( .A1(n1186), .A2(n1185), .ZN(n1026) );
XOR2_X1 U890 ( .A(n1193), .B(n1146), .Z(G21) );
NAND4_X1 U891 ( .A1(n1192), .A2(n1183), .A3(n1185), .A4(n1186), .ZN(n1146) );
INV_X1 U892 ( .A(n1194), .ZN(n1185) );
NAND2_X1 U893 ( .A1(n1195), .A2(n1196), .ZN(G18) );
OR2_X1 U894 ( .A1(n1147), .A2(G116), .ZN(n1196) );
XOR2_X1 U895 ( .A(n1197), .B(KEYINPUT37), .Z(n1195) );
NAND2_X1 U896 ( .A1(G116), .A2(n1147), .ZN(n1197) );
NAND3_X1 U897 ( .A1(n1037), .A2(n1008), .A3(n1192), .ZN(n1147) );
AND3_X1 U898 ( .A1(n1033), .A2(n1198), .A3(n1038), .ZN(n1192) );
AND2_X1 U899 ( .A1(n1178), .A2(n1040), .ZN(n1008) );
XOR2_X1 U900 ( .A(n1199), .B(KEYINPUT63), .Z(n1178) );
XOR2_X1 U901 ( .A(G113), .B(n1200), .Z(G15) );
NOR3_X1 U902 ( .A1(n1150), .A2(KEYINPUT55), .A3(n1201), .ZN(n1200) );
NAND4_X1 U903 ( .A1(n1038), .A2(n1009), .A3(n1037), .A4(n1198), .ZN(n1150) );
AND2_X1 U904 ( .A1(n1194), .A2(n1186), .ZN(n1037) );
INV_X1 U905 ( .A(n1159), .ZN(n1009) );
NAND2_X1 U906 ( .A1(n1202), .A2(n1179), .ZN(n1159) );
INV_X1 U907 ( .A(n1040), .ZN(n1179) );
NOR2_X1 U908 ( .A1(n1203), .A2(n1023), .ZN(n1038) );
XNOR2_X1 U909 ( .A(n1173), .B(n1204), .ZN(G12) );
NOR2_X1 U910 ( .A1(KEYINPUT61), .A2(n1205), .ZN(n1204) );
NAND3_X1 U911 ( .A1(n1183), .A2(n1174), .A3(n1021), .ZN(n1173) );
NOR2_X1 U912 ( .A1(n1186), .A2(n1194), .ZN(n1021) );
XOR2_X1 U913 ( .A(n1206), .B(n1092), .Z(n1194) );
AND2_X1 U914 ( .A1(G217), .A2(n1207), .ZN(n1092) );
OR2_X1 U915 ( .A1(n1089), .A2(G902), .ZN(n1206) );
XNOR2_X1 U916 ( .A(n1208), .B(n1209), .ZN(n1089) );
XOR2_X1 U917 ( .A(G137), .B(n1210), .Z(n1209) );
AND3_X1 U918 ( .A1(n1211), .A2(G234), .A3(G221), .ZN(n1210) );
XOR2_X1 U919 ( .A(KEYINPUT54), .B(n1070), .Z(n1211) );
NAND2_X1 U920 ( .A1(n1212), .A2(n1213), .ZN(n1208) );
OR2_X1 U921 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U922 ( .A(n1216), .B(KEYINPUT32), .Z(n1212) );
NAND2_X1 U923 ( .A1(n1215), .A2(n1214), .ZN(n1216) );
XNOR2_X1 U924 ( .A(n1217), .B(n1218), .ZN(n1214) );
XOR2_X1 U925 ( .A(n1205), .B(G119), .Z(n1217) );
XOR2_X1 U926 ( .A(G140), .B(n1219), .Z(n1215) );
XNOR2_X1 U927 ( .A(n1220), .B(G472), .ZN(n1186) );
NAND2_X1 U928 ( .A1(n1221), .A2(n1140), .ZN(n1220) );
XOR2_X1 U929 ( .A(n1118), .B(n1222), .Z(n1221) );
XOR2_X1 U930 ( .A(G101), .B(n1223), .Z(n1222) );
NOR2_X1 U931 ( .A1(KEYINPUT60), .A2(n1067), .ZN(n1223) );
XOR2_X1 U932 ( .A(n1224), .B(n1225), .Z(n1118) );
XOR2_X1 U933 ( .A(G119), .B(n1226), .Z(n1225) );
XOR2_X1 U934 ( .A(KEYINPUT18), .B(G146), .Z(n1226) );
XOR2_X1 U935 ( .A(n1227), .B(n1228), .Z(n1224) );
XOR2_X1 U936 ( .A(n1229), .B(n1230), .Z(n1227) );
INV_X1 U937 ( .A(n1231), .ZN(n1230) );
NAND2_X1 U938 ( .A1(n1232), .A2(G210), .ZN(n1229) );
AND3_X1 U939 ( .A1(n1149), .A2(n1198), .A3(n1170), .ZN(n1174) );
NOR2_X1 U940 ( .A1(n1025), .A2(n1023), .ZN(n1170) );
AND2_X1 U941 ( .A1(G221), .A2(n1207), .ZN(n1023) );
NAND2_X1 U942 ( .A1(G234), .A2(n1140), .ZN(n1207) );
INV_X1 U943 ( .A(n1203), .ZN(n1025) );
NAND2_X1 U944 ( .A1(n1233), .A2(n1234), .ZN(n1203) );
OR2_X1 U945 ( .A1(n1053), .A2(G469), .ZN(n1234) );
XOR2_X1 U946 ( .A(n1235), .B(KEYINPUT3), .Z(n1233) );
NAND2_X1 U947 ( .A1(G469), .A2(n1053), .ZN(n1235) );
NAND2_X1 U948 ( .A1(n1236), .A2(n1140), .ZN(n1053) );
XOR2_X1 U949 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U950 ( .A(n1130), .B(n1239), .Z(n1238) );
XOR2_X1 U951 ( .A(n1240), .B(n1241), .Z(n1130) );
XOR2_X1 U952 ( .A(G101), .B(n1068), .Z(n1241) );
XNOR2_X1 U953 ( .A(n1242), .B(n1243), .ZN(n1068) );
NOR3_X1 U954 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1243) );
NOR2_X1 U955 ( .A1(n1247), .A2(n1175), .ZN(n1246) );
AND3_X1 U956 ( .A1(n1175), .A2(n1247), .A3(KEYINPUT22), .ZN(n1245) );
AND2_X1 U957 ( .A1(KEYINPUT13), .A2(n1248), .ZN(n1247) );
INV_X1 U958 ( .A(G146), .ZN(n1175) );
NOR2_X1 U959 ( .A1(KEYINPUT22), .A2(n1248), .ZN(n1244) );
NAND2_X1 U960 ( .A1(KEYINPUT43), .A2(n1218), .ZN(n1242) );
XOR2_X1 U961 ( .A(n1205), .B(KEYINPUT28), .Z(n1240) );
XOR2_X1 U962 ( .A(n1249), .B(n1250), .Z(n1237) );
XNOR2_X1 U963 ( .A(G107), .B(n1251), .ZN(n1250) );
NAND2_X1 U964 ( .A1(KEYINPUT19), .A2(n1115), .ZN(n1251) );
INV_X1 U965 ( .A(n1067), .ZN(n1115) );
XNOR2_X1 U966 ( .A(n1252), .B(n1253), .ZN(n1067) );
XOR2_X1 U967 ( .A(G134), .B(n1127), .Z(n1252) );
INV_X1 U968 ( .A(G137), .ZN(n1127) );
NAND2_X1 U969 ( .A1(KEYINPUT58), .A2(G227), .ZN(n1249) );
NAND2_X1 U970 ( .A1(n999), .A2(n1254), .ZN(n1198) );
NAND3_X1 U971 ( .A1(n1085), .A2(n1190), .A3(G902), .ZN(n1254) );
NOR2_X1 U972 ( .A1(n1070), .A2(G898), .ZN(n1085) );
NAND3_X1 U973 ( .A1(n1190), .A2(n1070), .A3(G952), .ZN(n999) );
NAND2_X1 U974 ( .A1(G237), .A2(G234), .ZN(n1190) );
INV_X1 U975 ( .A(n1201), .ZN(n1149) );
XOR2_X1 U976 ( .A(n1012), .B(KEYINPUT20), .Z(n1201) );
INV_X1 U977 ( .A(n1033), .ZN(n1012) );
NOR2_X1 U978 ( .A1(n1035), .A2(n1034), .ZN(n1033) );
AND2_X1 U979 ( .A1(G214), .A2(n1255), .ZN(n1034) );
XNOR2_X1 U980 ( .A(KEYINPUT0), .B(n1256), .ZN(n1255) );
XOR2_X1 U981 ( .A(n1257), .B(n1139), .Z(n1035) );
AND2_X1 U982 ( .A1(G210), .A2(n1256), .ZN(n1139) );
NAND2_X1 U983 ( .A1(n1258), .A2(n1140), .ZN(n1256) );
XOR2_X1 U984 ( .A(KEYINPUT40), .B(G237), .Z(n1258) );
NAND2_X1 U985 ( .A1(n1259), .A2(n1140), .ZN(n1257) );
XOR2_X1 U986 ( .A(n1260), .B(n1261), .Z(n1259) );
INV_X1 U987 ( .A(n1138), .ZN(n1261) );
XOR2_X1 U988 ( .A(n1231), .B(n1262), .Z(n1138) );
XNOR2_X1 U989 ( .A(n1263), .B(n1219), .ZN(n1262) );
NAND2_X1 U990 ( .A1(G224), .A2(n1264), .ZN(n1263) );
XOR2_X1 U991 ( .A(KEYINPUT15), .B(G953), .Z(n1264) );
XOR2_X1 U992 ( .A(n1265), .B(n1266), .Z(n1231) );
NOR2_X1 U993 ( .A1(KEYINPUT9), .A2(n1267), .ZN(n1266) );
XOR2_X1 U994 ( .A(n1248), .B(KEYINPUT27), .Z(n1265) );
INV_X1 U995 ( .A(G143), .ZN(n1248) );
NAND2_X1 U996 ( .A1(KEYINPUT47), .A2(n1135), .ZN(n1260) );
XOR2_X1 U997 ( .A(n1083), .B(KEYINPUT21), .Z(n1135) );
XNOR2_X1 U998 ( .A(n1268), .B(n1269), .ZN(n1083) );
XOR2_X1 U999 ( .A(n1270), .B(n1271), .Z(n1269) );
NAND2_X1 U1000 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NAND2_X1 U1001 ( .A1(n1228), .A2(G119), .ZN(n1273) );
NAND2_X1 U1002 ( .A1(n1274), .A2(n1193), .ZN(n1272) );
INV_X1 U1003 ( .A(G119), .ZN(n1193) );
XNOR2_X1 U1004 ( .A(n1228), .B(KEYINPUT34), .ZN(n1274) );
XOR2_X1 U1005 ( .A(G113), .B(G116), .Z(n1228) );
NAND2_X1 U1006 ( .A1(n1275), .A2(n1276), .ZN(n1270) );
NAND3_X1 U1007 ( .A1(KEYINPUT29), .A2(n1111), .A3(n1277), .ZN(n1276) );
XOR2_X1 U1008 ( .A(n1278), .B(G101), .Z(n1277) );
NAND2_X1 U1009 ( .A1(G107), .A2(n1279), .ZN(n1278) );
INV_X1 U1010 ( .A(KEYINPUT10), .ZN(n1279) );
NAND2_X1 U1011 ( .A1(n1280), .A2(n1281), .ZN(n1275) );
NAND2_X1 U1012 ( .A1(KEYINPUT29), .A2(n1111), .ZN(n1281) );
INV_X1 U1013 ( .A(G104), .ZN(n1111) );
XOR2_X1 U1014 ( .A(n1121), .B(n1282), .Z(n1280) );
NOR2_X1 U1015 ( .A1(G107), .A2(KEYINPUT10), .ZN(n1282) );
INV_X1 U1016 ( .A(G101), .ZN(n1121) );
XOR2_X1 U1017 ( .A(n1205), .B(n1283), .Z(n1268) );
XOR2_X1 U1018 ( .A(KEYINPUT42), .B(G122), .Z(n1283) );
INV_X1 U1019 ( .A(G110), .ZN(n1205) );
INV_X1 U1020 ( .A(n1005), .ZN(n1183) );
NAND2_X1 U1021 ( .A1(n1202), .A2(n1040), .ZN(n1005) );
XOR2_X1 U1022 ( .A(n1284), .B(G475), .Z(n1040) );
NAND2_X1 U1023 ( .A1(n1108), .A2(n1140), .ZN(n1284) );
INV_X1 U1024 ( .A(G902), .ZN(n1140) );
XOR2_X1 U1025 ( .A(n1285), .B(n1286), .Z(n1108) );
XOR2_X1 U1026 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U1027 ( .A(G113), .B(n1191), .Z(n1288) );
INV_X1 U1028 ( .A(G122), .ZN(n1191) );
NAND2_X1 U1029 ( .A1(n1289), .A2(KEYINPUT45), .ZN(n1287) );
XOR2_X1 U1030 ( .A(n1290), .B(G143), .Z(n1289) );
NAND2_X1 U1031 ( .A1(n1232), .A2(G214), .ZN(n1290) );
NOR2_X1 U1032 ( .A1(G953), .A2(G237), .ZN(n1232) );
XNOR2_X1 U1033 ( .A(n1219), .B(n1132), .ZN(n1285) );
XNOR2_X1 U1034 ( .A(n1253), .B(n1239), .ZN(n1132) );
XOR2_X1 U1035 ( .A(G104), .B(G140), .Z(n1239) );
XNOR2_X1 U1036 ( .A(G131), .B(KEYINPUT46), .ZN(n1253) );
XOR2_X1 U1037 ( .A(G125), .B(G146), .Z(n1219) );
XOR2_X1 U1038 ( .A(n1199), .B(KEYINPUT23), .Z(n1202) );
NAND3_X1 U1039 ( .A1(n1291), .A2(n1292), .A3(n1047), .ZN(n1199) );
NAND2_X1 U1040 ( .A1(n1045), .A2(n1293), .ZN(n1047) );
OR3_X1 U1041 ( .A1(n1293), .A2(n1045), .A3(KEYINPUT38), .ZN(n1292) );
INV_X1 U1042 ( .A(G478), .ZN(n1293) );
NAND2_X1 U1043 ( .A1(KEYINPUT38), .A2(n1045), .ZN(n1291) );
NOR2_X1 U1044 ( .A1(G902), .A2(n1098), .ZN(n1045) );
AND2_X1 U1045 ( .A1(n1294), .A2(n1295), .ZN(n1098) );
NAND2_X1 U1046 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
NAND3_X1 U1047 ( .A1(G234), .A2(n1070), .A3(G217), .ZN(n1297) );
XOR2_X1 U1048 ( .A(n1298), .B(KEYINPUT14), .Z(n1294) );
NAND4_X1 U1049 ( .A1(G217), .A2(G234), .A3(n1299), .A4(n1070), .ZN(n1298) );
INV_X1 U1050 ( .A(G953), .ZN(n1070) );
INV_X1 U1051 ( .A(n1296), .ZN(n1299) );
XOR2_X1 U1052 ( .A(n1300), .B(n1301), .Z(n1296) );
XNOR2_X1 U1053 ( .A(n1302), .B(n1133), .ZN(n1301) );
XOR2_X1 U1054 ( .A(G134), .B(G107), .Z(n1133) );
NAND2_X1 U1055 ( .A1(KEYINPUT17), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1056 ( .A(KEYINPUT4), .B(n1218), .Z(n1303) );
INV_X1 U1057 ( .A(n1267), .ZN(n1218) );
XNOR2_X1 U1058 ( .A(G128), .B(KEYINPUT53), .ZN(n1267) );
XNOR2_X1 U1059 ( .A(G116), .B(n1304), .ZN(n1300) );
XOR2_X1 U1060 ( .A(G143), .B(G122), .Z(n1304) );
endmodule


