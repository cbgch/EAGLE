//Key = 1110010010101111100001101010101000000101011000100010000011001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310;

XOR2_X1 U721 ( .A(n987), .B(n988), .Z(G9) );
NAND2_X1 U722 ( .A1(n989), .A2(KEYINPUT5), .ZN(n987) );
XNOR2_X1 U723 ( .A(G107), .B(KEYINPUT20), .ZN(n989) );
NOR2_X1 U724 ( .A1(n990), .A2(n991), .ZN(G75) );
NOR4_X1 U725 ( .A1(n992), .A2(n993), .A3(G953), .A4(n994), .ZN(n991) );
NOR2_X1 U726 ( .A1(n995), .A2(n996), .ZN(n993) );
NOR2_X1 U727 ( .A1(n997), .A2(n998), .ZN(n995) );
NOR3_X1 U728 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n998) );
NOR2_X1 U729 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NOR2_X1 U730 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NOR2_X1 U731 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NOR2_X1 U732 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NOR2_X1 U733 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NOR2_X1 U734 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NOR2_X1 U735 ( .A1(n1014), .A2(n1015), .ZN(n1006) );
NOR2_X1 U736 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR2_X1 U737 ( .A1(KEYINPUT48), .A2(n1018), .ZN(n1016) );
INV_X1 U738 ( .A(n1019), .ZN(n1018) );
NOR2_X1 U739 ( .A1(n1020), .A2(n1015), .ZN(n1002) );
NOR2_X1 U740 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U741 ( .A1(n1023), .A2(n1009), .ZN(n1022) );
NOR2_X1 U742 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
XNOR2_X1 U743 ( .A(n1026), .B(KEYINPUT46), .ZN(n1025) );
AND3_X1 U744 ( .A1(KEYINPUT48), .A2(n1005), .A3(n1019), .ZN(n1021) );
NOR4_X1 U745 ( .A1(n1027), .A2(n1009), .A3(n1015), .A4(n1005), .ZN(n997) );
INV_X1 U746 ( .A(n1028), .ZN(n1005) );
NOR2_X1 U747 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U748 ( .A1(n999), .A2(n1031), .ZN(n1029) );
INV_X1 U749 ( .A(n1032), .ZN(n999) );
NAND2_X1 U750 ( .A1(n1033), .A2(n1034), .ZN(n992) );
XOR2_X1 U751 ( .A(KEYINPUT52), .B(n1035), .Z(n1034) );
NOR3_X1 U752 ( .A1(n994), .A2(G953), .A3(G952), .ZN(n990) );
AND4_X1 U753 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n994) );
NOR4_X1 U754 ( .A1(n1040), .A2(n1041), .A3(n1015), .A4(n1042), .ZN(n1039) );
XNOR2_X1 U755 ( .A(G469), .B(n1043), .ZN(n1042) );
XNOR2_X1 U756 ( .A(n1044), .B(n1045), .ZN(n1040) );
NOR2_X1 U757 ( .A1(G478), .A2(KEYINPUT34), .ZN(n1045) );
NOR3_X1 U758 ( .A1(n1046), .A2(n1047), .A3(n1000), .ZN(n1038) );
NAND2_X1 U759 ( .A1(n1048), .A2(n1049), .ZN(n1036) );
XOR2_X1 U760 ( .A(n1050), .B(n1051), .Z(G72) );
NOR2_X1 U761 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U762 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NAND2_X1 U763 ( .A1(n1056), .A2(n1057), .ZN(n1050) );
NAND2_X1 U764 ( .A1(n1058), .A2(n1053), .ZN(n1057) );
XOR2_X1 U765 ( .A(n1059), .B(n1035), .Z(n1058) );
OR3_X1 U766 ( .A1(n1059), .A2(n1055), .A3(n1053), .ZN(n1056) );
NAND2_X1 U767 ( .A1(KEYINPUT26), .A2(n1060), .ZN(n1059) );
XOR2_X1 U768 ( .A(n1061), .B(n1062), .Z(n1060) );
XOR2_X1 U769 ( .A(n1063), .B(n1064), .Z(n1062) );
XOR2_X1 U770 ( .A(n1065), .B(n1066), .Z(n1061) );
NAND2_X1 U771 ( .A1(KEYINPUT61), .A2(n1067), .ZN(n1065) );
XOR2_X1 U772 ( .A(n1068), .B(n1069), .Z(G69) );
XOR2_X1 U773 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND2_X1 U774 ( .A1(G953), .A2(n1072), .ZN(n1071) );
NAND2_X1 U775 ( .A1(G898), .A2(G224), .ZN(n1072) );
NAND3_X1 U776 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1070) );
NAND2_X1 U777 ( .A1(G953), .A2(n1076), .ZN(n1075) );
NAND2_X1 U778 ( .A1(n1077), .A2(n1078), .ZN(n1074) );
XNOR2_X1 U779 ( .A(n1079), .B(n1080), .ZN(n1078) );
XOR2_X1 U780 ( .A(KEYINPUT2), .B(KEYINPUT10), .Z(n1080) );
XNOR2_X1 U781 ( .A(n1081), .B(n1082), .ZN(n1077) );
XOR2_X1 U782 ( .A(n1083), .B(n1084), .Z(n1082) );
NAND2_X1 U783 ( .A1(n1085), .A2(n1086), .ZN(n1073) );
XOR2_X1 U784 ( .A(n1087), .B(n1088), .Z(n1086) );
XNOR2_X1 U785 ( .A(n1089), .B(KEYINPUT63), .ZN(n1085) );
NOR2_X1 U786 ( .A1(n1033), .A2(G953), .ZN(n1068) );
NOR2_X1 U787 ( .A1(n1090), .A2(n1091), .ZN(G66) );
XOR2_X1 U788 ( .A(KEYINPUT9), .B(n1092), .Z(n1091) );
NOR3_X1 U789 ( .A1(n1048), .A2(n1093), .A3(n1094), .ZN(n1090) );
AND2_X1 U790 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR3_X1 U791 ( .A1(n1096), .A2(n1097), .A3(n1095), .ZN(n1093) );
NAND3_X1 U792 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1095) );
XNOR2_X1 U793 ( .A(G217), .B(KEYINPUT24), .ZN(n1100) );
NOR2_X1 U794 ( .A1(n1092), .A2(n1101), .ZN(G63) );
NOR3_X1 U795 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
AND2_X1 U796 ( .A1(KEYINPUT31), .A2(n1105), .ZN(n1104) );
NOR2_X1 U797 ( .A1(KEYINPUT31), .A2(n1106), .ZN(n1103) );
NOR2_X1 U798 ( .A1(n1107), .A2(n1044), .ZN(n1106) );
NOR2_X1 U799 ( .A1(n1108), .A2(n1105), .ZN(n1107) );
AND2_X1 U800 ( .A1(n1098), .A2(G478), .ZN(n1108) );
NOR3_X1 U801 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1102) );
INV_X1 U802 ( .A(G478), .ZN(n1111) );
NOR2_X1 U803 ( .A1(KEYINPUT31), .A2(n1105), .ZN(n1110) );
NOR2_X1 U804 ( .A1(n1092), .A2(n1112), .ZN(G60) );
XNOR2_X1 U805 ( .A(n1113), .B(n1114), .ZN(n1112) );
XOR2_X1 U806 ( .A(KEYINPUT25), .B(n1115), .Z(n1114) );
NOR2_X1 U807 ( .A1(n1116), .A2(n1109), .ZN(n1115) );
XOR2_X1 U808 ( .A(G104), .B(n1117), .Z(G6) );
NOR2_X1 U809 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XOR2_X1 U810 ( .A(n1120), .B(KEYINPUT28), .Z(n1119) );
NAND2_X1 U811 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U812 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
INV_X1 U813 ( .A(KEYINPUT47), .ZN(n1124) );
NAND3_X1 U814 ( .A1(n1125), .A2(n1009), .A3(KEYINPUT47), .ZN(n1121) );
NOR2_X1 U815 ( .A1(n1092), .A2(n1126), .ZN(G57) );
XOR2_X1 U816 ( .A(n1127), .B(n1128), .Z(n1126) );
XNOR2_X1 U817 ( .A(n1129), .B(n1130), .ZN(n1128) );
XOR2_X1 U818 ( .A(KEYINPUT59), .B(n1131), .Z(n1130) );
NOR2_X1 U819 ( .A1(n1132), .A2(n1109), .ZN(n1131) );
XOR2_X1 U820 ( .A(n1063), .B(n1133), .Z(n1127) );
NOR2_X1 U821 ( .A1(n1092), .A2(n1134), .ZN(G54) );
XOR2_X1 U822 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U823 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U824 ( .A1(KEYINPUT33), .A2(n1139), .ZN(n1138) );
NAND2_X1 U825 ( .A1(KEYINPUT21), .A2(n1140), .ZN(n1137) );
XOR2_X1 U826 ( .A(n1141), .B(n1142), .Z(n1135) );
NOR2_X1 U827 ( .A1(n1143), .A2(n1109), .ZN(n1142) );
INV_X1 U828 ( .A(G469), .ZN(n1143) );
XNOR2_X1 U829 ( .A(G140), .B(G110), .ZN(n1141) );
NOR2_X1 U830 ( .A1(n1092), .A2(n1144), .ZN(G51) );
XOR2_X1 U831 ( .A(n1145), .B(n1146), .Z(n1144) );
XNOR2_X1 U832 ( .A(n1147), .B(n1148), .ZN(n1146) );
NOR3_X1 U833 ( .A1(n1149), .A2(n1150), .A3(n1109), .ZN(n1148) );
NAND2_X1 U834 ( .A1(G902), .A2(n1098), .ZN(n1109) );
NAND2_X1 U835 ( .A1(n1033), .A2(n1151), .ZN(n1098) );
XOR2_X1 U836 ( .A(KEYINPUT51), .B(n1035), .Z(n1151) );
AND4_X1 U837 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1035) );
AND4_X1 U838 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
NOR2_X1 U839 ( .A1(n1160), .A2(n1161), .ZN(n1154) );
INV_X1 U840 ( .A(n1162), .ZN(n1161) );
NAND3_X1 U841 ( .A1(n1163), .A2(n1026), .A3(n1164), .ZN(n1152) );
AND4_X1 U842 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1033) );
NOR4_X1 U843 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1168) );
NOR2_X1 U844 ( .A1(n1173), .A2(n988), .ZN(n1167) );
AND4_X1 U845 ( .A1(n1174), .A2(n1024), .A3(n1175), .A4(n1176), .ZN(n988) );
NAND2_X1 U846 ( .A1(n1011), .A2(n1177), .ZN(n1165) );
XOR2_X1 U847 ( .A(KEYINPUT6), .B(n1123), .Z(n1177) );
AND2_X1 U848 ( .A1(n1125), .A2(n1175), .ZN(n1123) );
AND3_X1 U849 ( .A1(n1030), .A2(n1176), .A3(n1026), .ZN(n1125) );
INV_X1 U850 ( .A(G210), .ZN(n1150) );
XNOR2_X1 U851 ( .A(KEYINPUT49), .B(n1178), .ZN(n1149) );
XNOR2_X1 U852 ( .A(n1179), .B(n1180), .ZN(n1145) );
NOR2_X1 U853 ( .A1(n1053), .A2(G952), .ZN(n1092) );
XNOR2_X1 U854 ( .A(G146), .B(n1181), .ZN(G48) );
NAND3_X1 U855 ( .A1(n1164), .A2(n1026), .A3(n1182), .ZN(n1181) );
XNOR2_X1 U856 ( .A(n1163), .B(KEYINPUT42), .ZN(n1182) );
XNOR2_X1 U857 ( .A(G143), .B(n1153), .ZN(G45) );
NAND4_X1 U858 ( .A1(n1164), .A2(n1017), .A3(n1183), .A4(n1184), .ZN(n1153) );
XOR2_X1 U859 ( .A(n1157), .B(n1185), .Z(G42) );
NAND2_X1 U860 ( .A1(KEYINPUT39), .A2(G140), .ZN(n1185) );
NAND3_X1 U861 ( .A1(n1026), .A2(n1019), .A3(n1186), .ZN(n1157) );
XNOR2_X1 U862 ( .A(G137), .B(n1156), .ZN(G39) );
NAND3_X1 U863 ( .A1(n1163), .A2(n1028), .A3(n1186), .ZN(n1156) );
NAND2_X1 U864 ( .A1(n1187), .A2(n1188), .ZN(G36) );
NAND2_X1 U865 ( .A1(G134), .A2(n1162), .ZN(n1188) );
XOR2_X1 U866 ( .A(KEYINPUT57), .B(n1189), .Z(n1187) );
NOR2_X1 U867 ( .A1(G134), .A2(n1162), .ZN(n1189) );
NAND3_X1 U868 ( .A1(n1017), .A2(n1024), .A3(n1186), .ZN(n1162) );
XOR2_X1 U869 ( .A(n1160), .B(n1190), .Z(G33) );
XNOR2_X1 U870 ( .A(KEYINPUT27), .B(n1067), .ZN(n1190) );
INV_X1 U871 ( .A(G131), .ZN(n1067) );
AND3_X1 U872 ( .A1(n1017), .A2(n1026), .A3(n1186), .ZN(n1160) );
AND3_X1 U873 ( .A1(n1030), .A2(n1191), .A3(n1192), .ZN(n1186) );
INV_X1 U874 ( .A(n1015), .ZN(n1192) );
NAND2_X1 U875 ( .A1(n1193), .A2(n1013), .ZN(n1015) );
INV_X1 U876 ( .A(n1012), .ZN(n1193) );
XOR2_X1 U877 ( .A(n1159), .B(n1194), .Z(G30) );
NAND2_X1 U878 ( .A1(KEYINPUT37), .A2(G128), .ZN(n1194) );
NAND3_X1 U879 ( .A1(n1163), .A2(n1024), .A3(n1164), .ZN(n1159) );
AND2_X1 U880 ( .A1(n1174), .A2(n1191), .ZN(n1164) );
NAND2_X1 U881 ( .A1(n1195), .A2(n1196), .ZN(G3) );
NAND2_X1 U882 ( .A1(G101), .A2(n1166), .ZN(n1196) );
XOR2_X1 U883 ( .A(n1197), .B(KEYINPUT58), .Z(n1195) );
OR2_X1 U884 ( .A1(n1166), .A2(G101), .ZN(n1197) );
NAND4_X1 U885 ( .A1(n1017), .A2(n1028), .A3(n1174), .A4(n1176), .ZN(n1166) );
XNOR2_X1 U886 ( .A(n1198), .B(n1199), .ZN(G27) );
NOR2_X1 U887 ( .A1(KEYINPUT17), .A2(n1158), .ZN(n1199) );
NAND4_X1 U888 ( .A1(n1019), .A2(n1011), .A3(n1026), .A4(n1200), .ZN(n1158) );
AND3_X1 U889 ( .A1(n1032), .A2(n1031), .A3(n1191), .ZN(n1200) );
NAND2_X1 U890 ( .A1(n996), .A2(n1201), .ZN(n1191) );
NAND4_X1 U891 ( .A1(G953), .A2(G902), .A3(n1202), .A4(n1055), .ZN(n1201) );
INV_X1 U892 ( .A(G900), .ZN(n1055) );
XOR2_X1 U893 ( .A(G122), .B(n1173), .Z(G24) );
AND4_X1 U894 ( .A1(n1203), .A2(n1175), .A3(n1183), .A4(n1184), .ZN(n1173) );
INV_X1 U895 ( .A(n1009), .ZN(n1175) );
NAND2_X1 U896 ( .A1(n1204), .A2(n1205), .ZN(n1009) );
XOR2_X1 U897 ( .A(G119), .B(n1172), .Z(G21) );
AND3_X1 U898 ( .A1(n1203), .A2(n1028), .A3(n1163), .ZN(n1172) );
NOR2_X1 U899 ( .A1(n1205), .A2(n1204), .ZN(n1163) );
INV_X1 U900 ( .A(n1041), .ZN(n1205) );
XNOR2_X1 U901 ( .A(n1206), .B(n1171), .ZN(G18) );
AND3_X1 U902 ( .A1(n1203), .A2(n1024), .A3(n1017), .ZN(n1171) );
AND2_X1 U903 ( .A1(n1207), .A2(n1183), .ZN(n1024) );
XNOR2_X1 U904 ( .A(G113), .B(n1208), .ZN(G15) );
NOR2_X1 U905 ( .A1(n1170), .A2(KEYINPUT40), .ZN(n1208) );
AND3_X1 U906 ( .A1(n1026), .A2(n1203), .A3(n1017), .ZN(n1170) );
AND2_X1 U907 ( .A1(n1204), .A2(n1041), .ZN(n1017) );
AND4_X1 U908 ( .A1(n1011), .A2(n1032), .A3(n1176), .A4(n1031), .ZN(n1203) );
NOR2_X1 U909 ( .A1(n1183), .A2(n1207), .ZN(n1026) );
INV_X1 U910 ( .A(n1184), .ZN(n1207) );
XNOR2_X1 U911 ( .A(n1169), .B(n1209), .ZN(G12) );
NAND2_X1 U912 ( .A1(KEYINPUT30), .A2(G110), .ZN(n1209) );
AND4_X1 U913 ( .A1(n1028), .A2(n1019), .A3(n1174), .A4(n1176), .ZN(n1169) );
NAND2_X1 U914 ( .A1(n996), .A2(n1210), .ZN(n1176) );
NAND4_X1 U915 ( .A1(G953), .A2(G902), .A3(n1202), .A4(n1076), .ZN(n1210) );
INV_X1 U916 ( .A(G898), .ZN(n1076) );
NAND3_X1 U917 ( .A1(n1202), .A2(n1053), .A3(G952), .ZN(n996) );
NAND2_X1 U918 ( .A1(G237), .A2(G234), .ZN(n1202) );
AND2_X1 U919 ( .A1(n1030), .A2(n1011), .ZN(n1174) );
INV_X1 U920 ( .A(n1118), .ZN(n1011) );
NAND2_X1 U921 ( .A1(n1012), .A2(n1013), .ZN(n1118) );
NAND2_X1 U922 ( .A1(G214), .A2(n1178), .ZN(n1013) );
XNOR2_X1 U923 ( .A(n1211), .B(n1212), .ZN(n1012) );
AND2_X1 U924 ( .A1(n1178), .A2(G210), .ZN(n1212) );
NAND2_X1 U925 ( .A1(n1213), .A2(n1214), .ZN(n1178) );
XNOR2_X1 U926 ( .A(G237), .B(KEYINPUT44), .ZN(n1213) );
NAND4_X1 U927 ( .A1(n1215), .A2(n1097), .A3(n1216), .A4(n1217), .ZN(n1211) );
NAND4_X1 U928 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(KEYINPUT0), .ZN(n1217) );
NAND2_X1 U929 ( .A1(n1221), .A2(n1222), .ZN(n1216) );
NAND2_X1 U930 ( .A1(n1220), .A2(n1223), .ZN(n1221) );
NAND2_X1 U931 ( .A1(KEYINPUT29), .A2(n1218), .ZN(n1223) );
INV_X1 U932 ( .A(n1179), .ZN(n1218) );
NAND2_X1 U933 ( .A1(n1179), .A2(n1224), .ZN(n1215) );
NAND3_X1 U934 ( .A1(n1225), .A2(n1226), .A3(n1227), .ZN(n1224) );
NAND2_X1 U935 ( .A1(n1222), .A2(n1219), .ZN(n1227) );
INV_X1 U936 ( .A(KEYINPUT29), .ZN(n1219) );
INV_X1 U937 ( .A(KEYINPUT0), .ZN(n1222) );
NAND2_X1 U938 ( .A1(n1228), .A2(n1229), .ZN(n1226) );
INV_X1 U939 ( .A(KEYINPUT38), .ZN(n1229) );
NAND2_X1 U940 ( .A1(n1220), .A2(n1230), .ZN(n1228) );
NAND2_X1 U941 ( .A1(KEYINPUT0), .A2(KEYINPUT29), .ZN(n1230) );
NAND2_X1 U942 ( .A1(KEYINPUT38), .A2(n1220), .ZN(n1225) );
XNOR2_X1 U943 ( .A(n1231), .B(n1232), .ZN(n1220) );
NOR2_X1 U944 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NOR3_X1 U945 ( .A1(KEYINPUT12), .A2(n1235), .A3(n1198), .ZN(n1234) );
NOR2_X1 U946 ( .A1(n1180), .A2(n1236), .ZN(n1233) );
INV_X1 U947 ( .A(KEYINPUT12), .ZN(n1236) );
XOR2_X1 U948 ( .A(n1235), .B(G125), .Z(n1180) );
NAND2_X1 U949 ( .A1(KEYINPUT14), .A2(n1147), .ZN(n1231) );
NAND2_X1 U950 ( .A1(G224), .A2(n1053), .ZN(n1147) );
XOR2_X1 U951 ( .A(n1237), .B(n1079), .Z(n1179) );
INV_X1 U952 ( .A(n1089), .ZN(n1079) );
XNOR2_X1 U953 ( .A(G110), .B(n1238), .ZN(n1089) );
XOR2_X1 U954 ( .A(n1239), .B(n1087), .Z(n1237) );
XOR2_X1 U955 ( .A(G119), .B(n1081), .Z(n1087) );
XNOR2_X1 U956 ( .A(G113), .B(n1206), .ZN(n1081) );
NAND2_X1 U957 ( .A1(KEYINPUT56), .A2(n1088), .ZN(n1239) );
XNOR2_X1 U958 ( .A(n1083), .B(G101), .ZN(n1088) );
NAND2_X1 U959 ( .A1(KEYINPUT60), .A2(n1240), .ZN(n1083) );
XNOR2_X1 U960 ( .A(n1241), .B(G104), .ZN(n1240) );
NOR2_X1 U961 ( .A1(n1032), .A2(n1000), .ZN(n1030) );
INV_X1 U962 ( .A(n1031), .ZN(n1000) );
NAND2_X1 U963 ( .A1(G221), .A2(n1099), .ZN(n1031) );
XNOR2_X1 U964 ( .A(n1043), .B(n1242), .ZN(n1032) );
NOR2_X1 U965 ( .A1(G469), .A2(KEYINPUT53), .ZN(n1242) );
NAND2_X1 U966 ( .A1(n1243), .A2(n1097), .ZN(n1043) );
XOR2_X1 U967 ( .A(n1244), .B(n1245), .Z(n1243) );
XOR2_X1 U968 ( .A(n1140), .B(n1246), .Z(n1245) );
NAND2_X1 U969 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND2_X1 U970 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
INV_X1 U971 ( .A(G140), .ZN(n1250) );
XNOR2_X1 U972 ( .A(KEYINPUT8), .B(n1251), .ZN(n1249) );
NAND2_X1 U973 ( .A1(n1252), .A2(G140), .ZN(n1247) );
XNOR2_X1 U974 ( .A(G110), .B(KEYINPUT16), .ZN(n1252) );
XOR2_X1 U975 ( .A(n1253), .B(n1254), .Z(n1140) );
XNOR2_X1 U976 ( .A(n1241), .B(n1255), .ZN(n1254) );
NOR2_X1 U977 ( .A1(G101), .A2(KEYINPUT4), .ZN(n1255) );
INV_X1 U978 ( .A(G107), .ZN(n1241) );
XOR2_X1 U979 ( .A(n1063), .B(n1256), .Z(n1253) );
XNOR2_X1 U980 ( .A(n1257), .B(G137), .ZN(n1063) );
XOR2_X1 U981 ( .A(KEYINPUT22), .B(n1139), .Z(n1244) );
NOR2_X1 U982 ( .A1(n1054), .A2(G953), .ZN(n1139) );
INV_X1 U983 ( .A(G227), .ZN(n1054) );
NOR2_X1 U984 ( .A1(n1041), .A2(n1204), .ZN(n1019) );
NOR2_X1 U985 ( .A1(n1258), .A2(n1047), .ZN(n1204) );
NOR2_X1 U986 ( .A1(n1049), .A2(n1048), .ZN(n1047) );
AND2_X1 U987 ( .A1(n1259), .A2(n1049), .ZN(n1258) );
NAND2_X1 U988 ( .A1(G217), .A2(n1099), .ZN(n1049) );
NAND2_X1 U989 ( .A1(G234), .A2(n1214), .ZN(n1099) );
XNOR2_X1 U990 ( .A(G902), .B(KEYINPUT55), .ZN(n1214) );
XOR2_X1 U991 ( .A(KEYINPUT45), .B(n1048), .Z(n1259) );
AND2_X1 U992 ( .A1(n1096), .A2(n1097), .ZN(n1048) );
XNOR2_X1 U993 ( .A(n1260), .B(n1261), .ZN(n1096) );
XOR2_X1 U994 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U995 ( .A(G137), .B(G119), .Z(n1263) );
XNOR2_X1 U996 ( .A(KEYINPUT7), .B(n1264), .ZN(n1262) );
XOR2_X1 U997 ( .A(n1265), .B(n1266), .Z(n1260) );
XOR2_X1 U998 ( .A(n1267), .B(n1066), .Z(n1266) );
XNOR2_X1 U999 ( .A(n1268), .B(n1251), .ZN(n1265) );
INV_X1 U1000 ( .A(G110), .ZN(n1251) );
NAND2_X1 U1001 ( .A1(n1269), .A2(G221), .ZN(n1268) );
XOR2_X1 U1002 ( .A(n1270), .B(n1132), .Z(n1041) );
INV_X1 U1003 ( .A(G472), .ZN(n1132) );
NAND2_X1 U1004 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XNOR2_X1 U1005 ( .A(KEYINPUT41), .B(n1097), .ZN(n1272) );
INV_X1 U1006 ( .A(G902), .ZN(n1097) );
XOR2_X1 U1007 ( .A(n1273), .B(n1274), .Z(n1271) );
XOR2_X1 U1008 ( .A(G137), .B(G134), .Z(n1274) );
XNOR2_X1 U1009 ( .A(n1133), .B(n1275), .ZN(n1273) );
NOR2_X1 U1010 ( .A1(KEYINPUT54), .A2(n1235), .ZN(n1275) );
XNOR2_X1 U1011 ( .A(n1129), .B(n1267), .ZN(n1235) );
NAND3_X1 U1012 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1129) );
OR2_X1 U1013 ( .A1(n1279), .A2(KEYINPUT50), .ZN(n1278) );
NAND3_X1 U1014 ( .A1(KEYINPUT50), .A2(n1280), .A3(n1264), .ZN(n1277) );
OR2_X1 U1015 ( .A1(n1264), .A2(n1280), .ZN(n1276) );
NOR2_X1 U1016 ( .A1(G143), .A2(KEYINPUT32), .ZN(n1280) );
INV_X1 U1017 ( .A(G146), .ZN(n1264) );
XNOR2_X1 U1018 ( .A(n1281), .B(n1282), .ZN(n1133) );
XOR2_X1 U1019 ( .A(n1283), .B(n1084), .Z(n1282) );
XNOR2_X1 U1020 ( .A(G101), .B(G119), .ZN(n1084) );
NAND2_X1 U1021 ( .A1(KEYINPUT1), .A2(n1206), .ZN(n1283) );
INV_X1 U1022 ( .A(G116), .ZN(n1206) );
XOR2_X1 U1023 ( .A(n1284), .B(n1285), .Z(n1281) );
XNOR2_X1 U1024 ( .A(G131), .B(n1286), .ZN(n1285) );
NAND2_X1 U1025 ( .A1(n1287), .A2(G210), .ZN(n1286) );
NAND2_X1 U1026 ( .A1(KEYINPUT15), .A2(n1288), .ZN(n1284) );
NOR2_X1 U1027 ( .A1(n1184), .A2(n1183), .ZN(n1028) );
XNOR2_X1 U1028 ( .A(G478), .B(n1289), .ZN(n1183) );
NOR2_X1 U1029 ( .A1(n1044), .A2(KEYINPUT43), .ZN(n1289) );
NOR2_X1 U1030 ( .A1(n1105), .A2(G902), .ZN(n1044) );
XNOR2_X1 U1031 ( .A(n1290), .B(n1291), .ZN(n1105) );
XOR2_X1 U1032 ( .A(n1257), .B(n1292), .Z(n1291) );
XOR2_X1 U1033 ( .A(n1293), .B(n1294), .Z(n1292) );
AND2_X1 U1034 ( .A1(n1269), .A2(G217), .ZN(n1294) );
AND2_X1 U1035 ( .A1(G234), .A2(n1053), .ZN(n1269) );
INV_X1 U1036 ( .A(G953), .ZN(n1053) );
NOR2_X1 U1037 ( .A1(KEYINPUT18), .A2(n1295), .ZN(n1293) );
XNOR2_X1 U1038 ( .A(n1296), .B(KEYINPUT13), .ZN(n1295) );
XOR2_X1 U1039 ( .A(G134), .B(n1267), .Z(n1257) );
XOR2_X1 U1040 ( .A(G128), .B(KEYINPUT19), .Z(n1267) );
XOR2_X1 U1041 ( .A(n1297), .B(n1298), .Z(n1290) );
XNOR2_X1 U1042 ( .A(KEYINPUT35), .B(n1279), .ZN(n1298) );
XNOR2_X1 U1043 ( .A(G107), .B(G116), .ZN(n1297) );
NAND3_X1 U1044 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1184) );
INV_X1 U1045 ( .A(n1046), .ZN(n1301) );
NOR2_X1 U1046 ( .A1(n1302), .A2(G475), .ZN(n1046) );
OR2_X1 U1047 ( .A1(n1037), .A2(KEYINPUT11), .ZN(n1300) );
NAND2_X1 U1048 ( .A1(G475), .A2(n1302), .ZN(n1037) );
NAND2_X1 U1049 ( .A1(n1303), .A2(n1113), .ZN(n1302) );
XNOR2_X1 U1050 ( .A(n1304), .B(n1305), .ZN(n1113) );
XOR2_X1 U1051 ( .A(n1256), .B(n1306), .Z(n1305) );
XNOR2_X1 U1052 ( .A(n1066), .B(n1238), .ZN(n1306) );
INV_X1 U1053 ( .A(n1296), .ZN(n1238) );
XOR2_X1 U1054 ( .A(G122), .B(KEYINPUT62), .Z(n1296) );
XNOR2_X1 U1055 ( .A(n1198), .B(G140), .ZN(n1066) );
INV_X1 U1056 ( .A(G125), .ZN(n1198) );
XNOR2_X1 U1057 ( .A(n1307), .B(n1064), .ZN(n1256) );
XNOR2_X1 U1058 ( .A(n1279), .B(G146), .ZN(n1064) );
INV_X1 U1059 ( .A(G143), .ZN(n1279) );
XNOR2_X1 U1060 ( .A(G104), .B(G131), .ZN(n1307) );
XOR2_X1 U1061 ( .A(n1308), .B(n1309), .Z(n1304) );
NOR2_X1 U1062 ( .A1(KEYINPUT23), .A2(n1288), .ZN(n1309) );
INV_X1 U1063 ( .A(G113), .ZN(n1288) );
XOR2_X1 U1064 ( .A(n1310), .B(KEYINPUT3), .Z(n1308) );
NAND2_X1 U1065 ( .A1(n1287), .A2(G214), .ZN(n1310) );
NOR2_X1 U1066 ( .A1(G953), .A2(G237), .ZN(n1287) );
XNOR2_X1 U1067 ( .A(G902), .B(KEYINPUT36), .ZN(n1303) );
NAND2_X1 U1068 ( .A1(KEYINPUT11), .A2(n1116), .ZN(n1299) );
INV_X1 U1069 ( .A(G475), .ZN(n1116) );
endmodule


