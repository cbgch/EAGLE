//Key = 1011010101100010001011101011000010111000100010011000101101010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328;

XNOR2_X1 U743 ( .A(G107), .B(n1023), .ZN(G9) );
NAND3_X1 U744 ( .A1(n1024), .A2(n1025), .A3(KEYINPUT14), .ZN(n1023) );
INV_X1 U745 ( .A(n1026), .ZN(n1025) );
NOR2_X1 U746 ( .A1(n1027), .A2(n1028), .ZN(G75) );
NOR3_X1 U747 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NAND3_X1 U748 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1029) );
NAND3_X1 U749 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NAND2_X1 U750 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NAND4_X1 U751 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1035) );
XOR2_X1 U752 ( .A(n1044), .B(KEYINPUT42), .Z(n1042) );
NAND2_X1 U753 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND3_X1 U754 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1041) );
NAND2_X1 U755 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND2_X1 U756 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U757 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U758 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U759 ( .A1(n1058), .A2(n1059), .ZN(n1050) );
INV_X1 U760 ( .A(n1060), .ZN(n1059) );
NAND2_X1 U761 ( .A1(n1045), .A2(n1061), .ZN(n1040) );
NAND2_X1 U762 ( .A1(n1062), .A2(n1063), .ZN(n1032) );
XOR2_X1 U763 ( .A(n1039), .B(KEYINPUT5), .Z(n1062) );
NAND2_X1 U764 ( .A1(n1045), .A2(n1047), .ZN(n1039) );
AND3_X1 U765 ( .A1(n1058), .A2(n1052), .A3(n1049), .ZN(n1045) );
INV_X1 U766 ( .A(n1064), .ZN(n1049) );
NOR3_X1 U767 ( .A1(n1030), .A2(G952), .A3(n1065), .ZN(n1027) );
INV_X1 U768 ( .A(n1033), .ZN(n1065) );
NAND4_X1 U769 ( .A1(n1066), .A2(n1052), .A3(n1067), .A4(n1068), .ZN(n1033) );
NOR4_X1 U770 ( .A1(n1038), .A2(n1056), .A3(n1069), .A4(n1070), .ZN(n1068) );
XNOR2_X1 U771 ( .A(n1071), .B(n1072), .ZN(n1070) );
NAND2_X1 U772 ( .A1(KEYINPUT44), .A2(n1073), .ZN(n1071) );
INV_X1 U773 ( .A(n1074), .ZN(n1056) );
XOR2_X1 U774 ( .A(n1075), .B(n1076), .Z(n1067) );
XOR2_X1 U775 ( .A(KEYINPUT36), .B(KEYINPUT3), .Z(n1076) );
XNOR2_X1 U776 ( .A(n1077), .B(n1078), .ZN(n1075) );
XNOR2_X1 U777 ( .A(n1079), .B(KEYINPUT43), .ZN(n1066) );
INV_X1 U778 ( .A(n1080), .ZN(n1030) );
XOR2_X1 U779 ( .A(n1081), .B(n1082), .Z(G72) );
XOR2_X1 U780 ( .A(n1083), .B(n1084), .Z(n1082) );
NOR3_X1 U781 ( .A1(n1085), .A2(KEYINPUT29), .A3(G953), .ZN(n1084) );
NOR2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XNOR2_X1 U783 ( .A(KEYINPUT17), .B(n1088), .ZN(n1087) );
NOR2_X1 U784 ( .A1(n1089), .A2(n1090), .ZN(n1083) );
XOR2_X1 U785 ( .A(n1091), .B(n1092), .Z(n1090) );
XOR2_X1 U786 ( .A(n1093), .B(n1094), .Z(n1092) );
XNOR2_X1 U787 ( .A(G131), .B(KEYINPUT59), .ZN(n1094) );
NAND2_X1 U788 ( .A1(KEYINPUT26), .A2(n1095), .ZN(n1093) );
XNOR2_X1 U789 ( .A(n1096), .B(n1097), .ZN(n1091) );
NOR2_X1 U790 ( .A1(G900), .A2(n1098), .ZN(n1089) );
NOR2_X1 U791 ( .A1(n1099), .A2(n1098), .ZN(n1081) );
NOR2_X1 U792 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XOR2_X1 U793 ( .A(n1102), .B(n1103), .Z(G69) );
XOR2_X1 U794 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U795 ( .A1(n1106), .A2(G953), .ZN(n1105) );
NOR2_X1 U796 ( .A1(n1107), .A2(n1108), .ZN(n1104) );
XNOR2_X1 U797 ( .A(n1109), .B(n1110), .ZN(n1108) );
XOR2_X1 U798 ( .A(n1111), .B(KEYINPUT10), .Z(n1107) );
NAND2_X1 U799 ( .A1(G953), .A2(n1112), .ZN(n1111) );
NOR2_X1 U800 ( .A1(n1113), .A2(n1098), .ZN(n1102) );
NOR2_X1 U801 ( .A1(n1114), .A2(n1112), .ZN(n1113) );
NOR2_X1 U802 ( .A1(n1115), .A2(n1116), .ZN(G66) );
XOR2_X1 U803 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U804 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NOR2_X1 U805 ( .A1(n1115), .A2(n1121), .ZN(G63) );
XOR2_X1 U806 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U807 ( .A1(n1124), .A2(n1120), .ZN(n1123) );
INV_X1 U808 ( .A(G478), .ZN(n1124) );
NOR2_X1 U809 ( .A1(n1115), .A2(n1125), .ZN(G60) );
XNOR2_X1 U810 ( .A(n1126), .B(n1127), .ZN(n1125) );
XOR2_X1 U811 ( .A(KEYINPUT4), .B(n1128), .Z(n1127) );
NOR2_X1 U812 ( .A1(n1129), .A2(n1120), .ZN(n1128) );
XOR2_X1 U813 ( .A(n1130), .B(n1131), .Z(G6) );
NOR2_X1 U814 ( .A1(KEYINPUT45), .A2(n1132), .ZN(n1131) );
NOR2_X1 U815 ( .A1(n1133), .A2(n1026), .ZN(n1130) );
XNOR2_X1 U816 ( .A(n1134), .B(KEYINPUT19), .ZN(n1133) );
NOR2_X1 U817 ( .A1(n1115), .A2(n1135), .ZN(G57) );
XOR2_X1 U818 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U819 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U820 ( .A(n1140), .B(n1141), .Z(n1136) );
NOR2_X1 U821 ( .A1(n1078), .A2(n1120), .ZN(n1141) );
INV_X1 U822 ( .A(G472), .ZN(n1078) );
XNOR2_X1 U823 ( .A(n1142), .B(n1143), .ZN(n1140) );
NOR2_X1 U824 ( .A1(G101), .A2(KEYINPUT28), .ZN(n1143) );
NOR2_X1 U825 ( .A1(n1115), .A2(n1144), .ZN(G54) );
XOR2_X1 U826 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U827 ( .A(n1147), .B(n1148), .Z(n1145) );
NOR2_X1 U828 ( .A1(n1149), .A2(n1120), .ZN(n1148) );
XOR2_X1 U829 ( .A(n1150), .B(G140), .Z(n1147) );
NAND2_X1 U830 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XNOR2_X1 U831 ( .A(KEYINPUT2), .B(n1153), .ZN(n1151) );
NOR2_X1 U832 ( .A1(n1115), .A2(n1154), .ZN(G51) );
XOR2_X1 U833 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U834 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U835 ( .A1(n1072), .A2(n1120), .ZN(n1158) );
NAND2_X1 U836 ( .A1(G902), .A2(n1031), .ZN(n1120) );
NAND3_X1 U837 ( .A1(n1159), .A2(n1088), .A3(n1106), .ZN(n1031) );
AND4_X1 U838 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1106) );
NOR4_X1 U839 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1163) );
NOR2_X1 U840 ( .A1(n1060), .A2(n1026), .ZN(n1167) );
NAND2_X1 U841 ( .A1(n1168), .A2(n1047), .ZN(n1026) );
NOR2_X1 U842 ( .A1(n1134), .A2(n1024), .ZN(n1060) );
NOR2_X1 U843 ( .A1(n1169), .A2(n1170), .ZN(n1165) );
NAND4_X1 U844 ( .A1(n1171), .A2(n1058), .A3(n1172), .A4(n1063), .ZN(n1170) );
INV_X1 U845 ( .A(n1173), .ZN(n1171) );
INV_X1 U846 ( .A(KEYINPUT49), .ZN(n1169) );
NOR2_X1 U847 ( .A1(KEYINPUT49), .A2(n1174), .ZN(n1164) );
NOR2_X1 U848 ( .A1(n1175), .A2(n1176), .ZN(n1162) );
INV_X1 U849 ( .A(n1086), .ZN(n1159) );
NAND4_X1 U850 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1086) );
NOR4_X1 U851 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1180) );
NAND2_X1 U852 ( .A1(KEYINPUT55), .A2(n1185), .ZN(n1155) );
NOR2_X1 U853 ( .A1(n1098), .A2(G952), .ZN(n1115) );
XNOR2_X1 U854 ( .A(G146), .B(n1179), .ZN(G48) );
NAND2_X1 U855 ( .A1(n1186), .A2(n1134), .ZN(n1179) );
XNOR2_X1 U856 ( .A(G143), .B(n1177), .ZN(G45) );
NAND3_X1 U857 ( .A1(n1046), .A2(n1187), .A3(n1188), .ZN(n1177) );
NOR3_X1 U858 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1188) );
XNOR2_X1 U859 ( .A(G140), .B(n1178), .ZN(G42) );
NAND3_X1 U860 ( .A1(n1134), .A2(n1192), .A3(n1061), .ZN(n1178) );
XOR2_X1 U861 ( .A(n1088), .B(n1193), .Z(G39) );
NOR2_X1 U862 ( .A1(G137), .A2(KEYINPUT13), .ZN(n1193) );
NAND2_X1 U863 ( .A1(n1192), .A2(n1172), .ZN(n1088) );
NAND2_X1 U864 ( .A1(n1194), .A2(n1195), .ZN(G36) );
OR2_X1 U865 ( .A1(n1196), .A2(G134), .ZN(n1195) );
NAND2_X1 U866 ( .A1(G134), .A2(n1197), .ZN(n1194) );
NAND2_X1 U867 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NAND2_X1 U868 ( .A1(n1184), .A2(n1200), .ZN(n1199) );
INV_X1 U869 ( .A(KEYINPUT7), .ZN(n1200) );
NAND2_X1 U870 ( .A1(KEYINPUT7), .A2(n1196), .ZN(n1198) );
NAND2_X1 U871 ( .A1(KEYINPUT40), .A2(n1184), .ZN(n1196) );
AND3_X1 U872 ( .A1(n1192), .A2(n1024), .A3(n1046), .ZN(n1184) );
XNOR2_X1 U873 ( .A(n1201), .B(n1183), .ZN(G33) );
AND3_X1 U874 ( .A1(n1134), .A2(n1192), .A3(n1046), .ZN(n1183) );
NOR4_X1 U875 ( .A1(n1202), .A2(n1054), .A3(n1190), .A4(n1038), .ZN(n1192) );
XOR2_X1 U876 ( .A(n1182), .B(n1203), .Z(G30) );
NOR2_X1 U877 ( .A1(KEYINPUT58), .A2(n1204), .ZN(n1203) );
AND2_X1 U878 ( .A1(n1186), .A2(n1024), .ZN(n1182) );
AND4_X1 U879 ( .A1(n1187), .A2(n1079), .A3(n1205), .A4(n1206), .ZN(n1186) );
XNOR2_X1 U880 ( .A(n1166), .B(n1207), .ZN(G3) );
XNOR2_X1 U881 ( .A(KEYINPUT0), .B(n1208), .ZN(n1207) );
AND3_X1 U882 ( .A1(n1052), .A2(n1168), .A3(n1046), .ZN(n1166) );
XOR2_X1 U883 ( .A(G125), .B(n1181), .Z(G27) );
AND4_X1 U884 ( .A1(n1061), .A2(n1134), .A3(n1209), .A4(n1058), .ZN(n1181) );
NOR2_X1 U885 ( .A1(n1190), .A2(n1210), .ZN(n1209) );
INV_X1 U886 ( .A(n1205), .ZN(n1190) );
NAND2_X1 U887 ( .A1(n1064), .A2(n1211), .ZN(n1205) );
NAND4_X1 U888 ( .A1(G953), .A2(G902), .A3(n1212), .A4(n1101), .ZN(n1211) );
INV_X1 U889 ( .A(G900), .ZN(n1101) );
XNOR2_X1 U890 ( .A(G122), .B(n1161), .ZN(G24) );
NAND4_X1 U891 ( .A1(n1213), .A2(n1047), .A3(n1214), .A4(n1215), .ZN(n1161) );
NOR2_X1 U892 ( .A1(n1206), .A2(n1079), .ZN(n1047) );
XNOR2_X1 U893 ( .A(n1216), .B(n1174), .ZN(G21) );
NAND2_X1 U894 ( .A1(n1213), .A2(n1172), .ZN(n1174) );
AND3_X1 U895 ( .A1(n1079), .A2(n1206), .A3(n1052), .ZN(n1172) );
XNOR2_X1 U896 ( .A(G119), .B(KEYINPUT18), .ZN(n1216) );
XOR2_X1 U897 ( .A(G116), .B(n1176), .Z(G18) );
AND3_X1 U898 ( .A1(n1213), .A2(n1024), .A3(n1046), .ZN(n1176) );
NOR2_X1 U899 ( .A1(n1215), .A2(n1189), .ZN(n1024) );
INV_X1 U900 ( .A(n1214), .ZN(n1189) );
XOR2_X1 U901 ( .A(n1175), .B(n1217), .Z(G15) );
XOR2_X1 U902 ( .A(KEYINPUT6), .B(G113), .Z(n1217) );
AND3_X1 U903 ( .A1(n1134), .A2(n1213), .A3(n1046), .ZN(n1175) );
AND2_X1 U904 ( .A1(n1218), .A2(n1206), .ZN(n1046) );
AND3_X1 U905 ( .A1(n1063), .A2(n1173), .A3(n1058), .ZN(n1213) );
AND2_X1 U906 ( .A1(n1219), .A2(n1074), .ZN(n1058) );
XNOR2_X1 U907 ( .A(KEYINPUT50), .B(n1069), .ZN(n1219) );
INV_X1 U908 ( .A(n1057), .ZN(n1069) );
NOR2_X1 U909 ( .A1(n1214), .A2(n1191), .ZN(n1134) );
INV_X1 U910 ( .A(n1215), .ZN(n1191) );
XNOR2_X1 U911 ( .A(G110), .B(n1160), .ZN(G12) );
NAND3_X1 U912 ( .A1(n1052), .A2(n1168), .A3(n1061), .ZN(n1160) );
NOR2_X1 U913 ( .A1(n1206), .A2(n1218), .ZN(n1061) );
INV_X1 U914 ( .A(n1079), .ZN(n1218) );
XOR2_X1 U915 ( .A(n1220), .B(n1119), .Z(n1079) );
NAND2_X1 U916 ( .A1(G217), .A2(n1221), .ZN(n1119) );
NAND2_X1 U917 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
XNOR2_X1 U918 ( .A(n1118), .B(KEYINPUT11), .ZN(n1222) );
XNOR2_X1 U919 ( .A(n1224), .B(n1225), .ZN(n1118) );
XOR2_X1 U920 ( .A(n1226), .B(n1227), .Z(n1225) );
XNOR2_X1 U921 ( .A(n1228), .B(n1229), .ZN(n1227) );
NOR2_X1 U922 ( .A1(KEYINPUT33), .A2(n1230), .ZN(n1228) );
XOR2_X1 U923 ( .A(n1231), .B(n1232), .Z(n1224) );
XNOR2_X1 U924 ( .A(n1233), .B(G110), .ZN(n1232) );
XOR2_X1 U925 ( .A(n1234), .B(n1235), .Z(n1231) );
NOR2_X1 U926 ( .A1(KEYINPUT60), .A2(n1204), .ZN(n1235) );
NAND3_X1 U927 ( .A1(n1236), .A2(n1098), .A3(G221), .ZN(n1234) );
XOR2_X1 U928 ( .A(KEYINPUT37), .B(n1237), .Z(n1236) );
NAND2_X1 U929 ( .A1(n1238), .A2(n1239), .ZN(n1206) );
NAND2_X1 U930 ( .A1(G472), .A2(n1077), .ZN(n1239) );
XOR2_X1 U931 ( .A(KEYINPUT47), .B(n1240), .Z(n1238) );
NOR2_X1 U932 ( .A1(G472), .A2(n1077), .ZN(n1240) );
NAND2_X1 U933 ( .A1(n1241), .A2(n1223), .ZN(n1077) );
XOR2_X1 U934 ( .A(n1242), .B(n1243), .Z(n1241) );
NOR2_X1 U935 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XOR2_X1 U936 ( .A(KEYINPUT16), .B(n1246), .Z(n1245) );
NOR2_X1 U937 ( .A1(n1142), .A2(n1247), .ZN(n1246) );
AND2_X1 U938 ( .A1(n1247), .A2(n1142), .ZN(n1244) );
NOR3_X1 U939 ( .A1(G237), .A2(G953), .A3(n1248), .ZN(n1142) );
XOR2_X1 U940 ( .A(G101), .B(KEYINPUT12), .Z(n1247) );
NOR2_X1 U941 ( .A1(KEYINPUT38), .A2(n1249), .ZN(n1242) );
XNOR2_X1 U942 ( .A(n1250), .B(n1139), .ZN(n1249) );
XOR2_X1 U943 ( .A(G113), .B(n1251), .Z(n1139) );
XNOR2_X1 U944 ( .A(n1233), .B(G116), .ZN(n1251) );
NAND2_X1 U945 ( .A1(n1252), .A2(n1253), .ZN(n1250) );
OR2_X1 U946 ( .A1(n1138), .A2(KEYINPUT15), .ZN(n1253) );
XNOR2_X1 U947 ( .A(n1254), .B(n1255), .ZN(n1138) );
NAND3_X1 U948 ( .A1(n1255), .A2(n1254), .A3(KEYINPUT15), .ZN(n1252) );
XOR2_X1 U949 ( .A(n1256), .B(KEYINPUT8), .Z(n1255) );
AND2_X1 U950 ( .A1(n1187), .A2(n1173), .ZN(n1168) );
NAND2_X1 U951 ( .A1(n1064), .A2(n1257), .ZN(n1173) );
NAND4_X1 U952 ( .A1(G953), .A2(G902), .A3(n1212), .A4(n1112), .ZN(n1257) );
INV_X1 U953 ( .A(G898), .ZN(n1112) );
NAND3_X1 U954 ( .A1(n1080), .A2(n1212), .A3(G952), .ZN(n1064) );
NAND2_X1 U955 ( .A1(G237), .A2(G234), .ZN(n1212) );
XOR2_X1 U956 ( .A(G953), .B(KEYINPUT62), .Z(n1080) );
NOR2_X1 U957 ( .A1(n1210), .A2(n1054), .ZN(n1187) );
NAND2_X1 U958 ( .A1(n1258), .A2(n1074), .ZN(n1054) );
NAND2_X1 U959 ( .A1(G221), .A2(n1221), .ZN(n1074) );
NAND2_X1 U960 ( .A1(G234), .A2(n1223), .ZN(n1221) );
XNOR2_X1 U961 ( .A(n1057), .B(KEYINPUT23), .ZN(n1258) );
XNOR2_X1 U962 ( .A(n1259), .B(n1260), .ZN(n1057) );
XNOR2_X1 U963 ( .A(KEYINPUT57), .B(n1149), .ZN(n1260) );
INV_X1 U964 ( .A(G469), .ZN(n1149) );
NAND2_X1 U965 ( .A1(n1261), .A2(n1223), .ZN(n1259) );
XOR2_X1 U966 ( .A(n1262), .B(n1146), .Z(n1261) );
XOR2_X1 U967 ( .A(n1254), .B(n1263), .Z(n1146) );
XNOR2_X1 U968 ( .A(n1264), .B(n1265), .ZN(n1263) );
NOR2_X1 U969 ( .A1(G953), .A2(n1100), .ZN(n1265) );
INV_X1 U970 ( .A(G227), .ZN(n1100) );
INV_X1 U971 ( .A(G110), .ZN(n1264) );
XOR2_X1 U972 ( .A(n1266), .B(n1095), .Z(n1254) );
XOR2_X1 U973 ( .A(G134), .B(n1226), .Z(n1095) );
XOR2_X1 U974 ( .A(G137), .B(KEYINPUT25), .Z(n1226) );
XNOR2_X1 U975 ( .A(G131), .B(KEYINPUT20), .ZN(n1266) );
XOR2_X1 U976 ( .A(n1267), .B(n1268), .Z(n1262) );
NOR2_X1 U977 ( .A1(G140), .A2(KEYINPUT31), .ZN(n1268) );
NAND2_X1 U978 ( .A1(n1152), .A2(n1153), .ZN(n1267) );
OR2_X1 U979 ( .A1(n1269), .A2(n1097), .ZN(n1153) );
NAND2_X1 U980 ( .A1(n1269), .A2(n1097), .ZN(n1152) );
XNOR2_X1 U981 ( .A(n1270), .B(KEYINPUT35), .ZN(n1097) );
XNOR2_X1 U982 ( .A(n1271), .B(n1272), .ZN(n1269) );
XOR2_X1 U983 ( .A(G104), .B(n1273), .Z(n1272) );
NOR2_X1 U984 ( .A1(G107), .A2(KEYINPUT61), .ZN(n1273) );
NAND2_X1 U985 ( .A1(KEYINPUT22), .A2(n1208), .ZN(n1271) );
INV_X1 U986 ( .A(n1063), .ZN(n1210) );
NOR2_X1 U987 ( .A1(n1037), .A2(n1038), .ZN(n1063) );
INV_X1 U988 ( .A(n1043), .ZN(n1038) );
NAND2_X1 U989 ( .A1(G214), .A2(n1274), .ZN(n1043) );
XOR2_X1 U990 ( .A(KEYINPUT24), .B(n1275), .Z(n1274) );
INV_X1 U991 ( .A(n1202), .ZN(n1037) );
XOR2_X1 U992 ( .A(n1073), .B(n1072), .Z(n1202) );
OR2_X1 U993 ( .A1(n1248), .A2(n1275), .ZN(n1072) );
NOR2_X1 U994 ( .A1(G902), .A2(G237), .ZN(n1275) );
INV_X1 U995 ( .A(G210), .ZN(n1248) );
NAND2_X1 U996 ( .A1(n1276), .A2(n1223), .ZN(n1073) );
XOR2_X1 U997 ( .A(n1277), .B(n1185), .Z(n1276) );
XNOR2_X1 U998 ( .A(n1278), .B(n1256), .ZN(n1185) );
XNOR2_X1 U999 ( .A(n1270), .B(KEYINPUT21), .ZN(n1256) );
XNOR2_X1 U1000 ( .A(n1279), .B(n1230), .ZN(n1270) );
XNOR2_X1 U1001 ( .A(G128), .B(G143), .ZN(n1279) );
XNOR2_X1 U1002 ( .A(G125), .B(n1280), .ZN(n1278) );
NOR2_X1 U1003 ( .A1(G953), .A2(n1114), .ZN(n1280) );
INV_X1 U1004 ( .A(G224), .ZN(n1114) );
XOR2_X1 U1005 ( .A(n1157), .B(KEYINPUT41), .Z(n1277) );
NAND3_X1 U1006 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1157) );
NAND2_X1 U1007 ( .A1(KEYINPUT56), .A2(n1284), .ZN(n1283) );
NAND2_X1 U1008 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND3_X1 U1009 ( .A1(n1287), .A2(n1288), .A3(n1285), .ZN(n1282) );
INV_X1 U1010 ( .A(n1110), .ZN(n1285) );
INV_X1 U1011 ( .A(KEYINPUT56), .ZN(n1288) );
NAND2_X1 U1012 ( .A1(KEYINPUT9), .A2(n1109), .ZN(n1287) );
NAND3_X1 U1013 ( .A1(KEYINPUT9), .A2(n1109), .A3(n1110), .ZN(n1281) );
XOR2_X1 U1014 ( .A(G110), .B(n1289), .Z(n1110) );
XNOR2_X1 U1015 ( .A(KEYINPUT1), .B(n1290), .ZN(n1289) );
INV_X1 U1016 ( .A(n1286), .ZN(n1109) );
NAND2_X1 U1017 ( .A1(n1291), .A2(n1292), .ZN(n1286) );
NAND2_X1 U1018 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XNOR2_X1 U1019 ( .A(G104), .B(G107), .ZN(n1293) );
NAND2_X1 U1020 ( .A1(n1295), .A2(n1296), .ZN(n1291) );
XOR2_X1 U1021 ( .A(KEYINPUT32), .B(n1294), .Z(n1296) );
XNOR2_X1 U1022 ( .A(n1208), .B(n1297), .ZN(n1294) );
NOR2_X1 U1023 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
XOR2_X1 U1024 ( .A(n1300), .B(KEYINPUT52), .Z(n1299) );
NAND2_X1 U1025 ( .A1(n1301), .A2(G113), .ZN(n1300) );
NOR2_X1 U1026 ( .A1(G113), .A2(n1301), .ZN(n1298) );
XOR2_X1 U1027 ( .A(n1302), .B(G116), .Z(n1301) );
NAND2_X1 U1028 ( .A1(KEYINPUT54), .A2(n1233), .ZN(n1302) );
INV_X1 U1029 ( .A(G119), .ZN(n1233) );
INV_X1 U1030 ( .A(G101), .ZN(n1208) );
XNOR2_X1 U1031 ( .A(n1303), .B(G104), .ZN(n1295) );
INV_X1 U1032 ( .A(G107), .ZN(n1303) );
NOR2_X1 U1033 ( .A1(n1214), .A2(n1215), .ZN(n1052) );
XOR2_X1 U1034 ( .A(n1304), .B(n1129), .Z(n1215) );
INV_X1 U1035 ( .A(G475), .ZN(n1129) );
NAND2_X1 U1036 ( .A1(n1126), .A2(n1223), .ZN(n1304) );
INV_X1 U1037 ( .A(G902), .ZN(n1223) );
XNOR2_X1 U1038 ( .A(n1305), .B(n1306), .ZN(n1126) );
XNOR2_X1 U1039 ( .A(n1229), .B(n1307), .ZN(n1306) );
XNOR2_X1 U1040 ( .A(n1308), .B(n1309), .ZN(n1307) );
NOR2_X1 U1041 ( .A1(KEYINPUT39), .A2(n1230), .ZN(n1309) );
XNOR2_X1 U1042 ( .A(G146), .B(KEYINPUT27), .ZN(n1230) );
NAND2_X1 U1043 ( .A1(KEYINPUT34), .A2(n1290), .ZN(n1308) );
INV_X1 U1044 ( .A(n1096), .ZN(n1229) );
XOR2_X1 U1045 ( .A(G125), .B(G140), .Z(n1096) );
XOR2_X1 U1046 ( .A(n1310), .B(n1311), .Z(n1305) );
XNOR2_X1 U1047 ( .A(G113), .B(n1312), .ZN(n1311) );
NAND2_X1 U1048 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
NAND2_X1 U1049 ( .A1(n1315), .A2(n1201), .ZN(n1314) );
XOR2_X1 U1050 ( .A(n1316), .B(KEYINPUT63), .Z(n1313) );
OR2_X1 U1051 ( .A1(n1201), .A2(n1315), .ZN(n1316) );
XNOR2_X1 U1052 ( .A(n1317), .B(G143), .ZN(n1315) );
NAND3_X1 U1053 ( .A1(n1318), .A2(n1098), .A3(G214), .ZN(n1317) );
INV_X1 U1054 ( .A(G237), .ZN(n1318) );
INV_X1 U1055 ( .A(G131), .ZN(n1201) );
NAND2_X1 U1056 ( .A1(KEYINPUT48), .A2(n1132), .ZN(n1310) );
INV_X1 U1057 ( .A(G104), .ZN(n1132) );
XOR2_X1 U1058 ( .A(G478), .B(n1319), .Z(n1214) );
NOR2_X1 U1059 ( .A1(G902), .A2(n1122), .ZN(n1319) );
XOR2_X1 U1060 ( .A(n1320), .B(n1321), .Z(n1122) );
NOR2_X1 U1061 ( .A1(KEYINPUT46), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1062 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1063 ( .A(n1325), .B(n1326), .Z(n1324) );
NOR2_X1 U1064 ( .A1(G143), .A2(KEYINPUT53), .ZN(n1326) );
XNOR2_X1 U1065 ( .A(G107), .B(n1327), .ZN(n1325) );
NOR2_X1 U1066 ( .A1(KEYINPUT30), .A2(n1290), .ZN(n1327) );
INV_X1 U1067 ( .A(G122), .ZN(n1290) );
XNOR2_X1 U1068 ( .A(G116), .B(n1328), .ZN(n1323) );
XNOR2_X1 U1069 ( .A(G134), .B(n1204), .ZN(n1328) );
INV_X1 U1070 ( .A(G128), .ZN(n1204) );
NAND3_X1 U1071 ( .A1(n1237), .A2(n1098), .A3(G217), .ZN(n1320) );
INV_X1 U1072 ( .A(G953), .ZN(n1098) );
XOR2_X1 U1073 ( .A(G234), .B(KEYINPUT51), .Z(n1237) );
endmodule


