//Key = 0110111011111000101110111101010101001111100010111000100100100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412;

NAND2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(G9) );
NAND2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U769 ( .A(KEYINPUT27), .B(n1074), .Z(n1070) );
NOR2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1074) );
NOR2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(G75) );
NOR3_X1 U772 ( .A1(n1077), .A2(G953), .A3(n1078), .ZN(n1076) );
XOR2_X1 U773 ( .A(KEYINPUT29), .B(n1079), .Z(n1077) );
NOR3_X1 U774 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NOR2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NOR2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NOR2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U778 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR2_X1 U780 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NOR2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U782 ( .A1(n1097), .A2(n1098), .ZN(n1093) );
NOR2_X1 U783 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NOR3_X1 U784 ( .A1(n1096), .A2(n1098), .A3(n1101), .ZN(n1089) );
NOR2_X1 U785 ( .A1(n1102), .A2(n1096), .ZN(n1085) );
NOR2_X1 U786 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U787 ( .A1(n1105), .A2(n1092), .ZN(n1104) );
NOR2_X1 U788 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR2_X1 U789 ( .A1(n1108), .A2(n1098), .ZN(n1107) );
NOR2_X1 U790 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U791 ( .A1(n1111), .A2(n1112), .ZN(n1109) );
XNOR2_X1 U792 ( .A(KEYINPUT47), .B(n1113), .ZN(n1111) );
NOR3_X1 U793 ( .A1(n1114), .A2(n1088), .A3(n1115), .ZN(n1106) );
NOR3_X1 U794 ( .A1(n1098), .A2(n1088), .A3(n1116), .ZN(n1103) );
NOR3_X1 U795 ( .A1(n1078), .A2(G953), .A3(G952), .ZN(n1075) );
AND4_X1 U796 ( .A1(n1117), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1078) );
NOR4_X1 U797 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1120) );
XOR2_X1 U798 ( .A(n1125), .B(KEYINPUT13), .Z(n1123) );
NAND2_X1 U799 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U800 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U801 ( .A(KEYINPUT23), .B(n1130), .Z(n1126) );
NOR2_X1 U802 ( .A1(n1128), .A2(n1129), .ZN(n1130) );
XNOR2_X1 U803 ( .A(n1131), .B(KEYINPUT61), .ZN(n1129) );
XNOR2_X1 U804 ( .A(n1132), .B(KEYINPUT0), .ZN(n1128) );
XOR2_X1 U805 ( .A(n1133), .B(n1134), .Z(n1122) );
XOR2_X1 U806 ( .A(KEYINPUT52), .B(n1135), .Z(n1134) );
NOR2_X1 U807 ( .A1(KEYINPUT54), .A2(n1136), .ZN(n1135) );
XOR2_X1 U808 ( .A(n1137), .B(n1138), .Z(G72) );
XOR2_X1 U809 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U810 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NOR2_X1 U811 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
XOR2_X1 U812 ( .A(KEYINPUT20), .B(G227), .Z(n1144) );
NAND2_X1 U813 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
NAND2_X1 U814 ( .A1(G953), .A2(n1143), .ZN(n1146) );
XOR2_X1 U815 ( .A(n1147), .B(n1148), .Z(n1145) );
XNOR2_X1 U816 ( .A(G125), .B(n1149), .ZN(n1148) );
XNOR2_X1 U817 ( .A(KEYINPUT14), .B(KEYINPUT1), .ZN(n1149) );
XOR2_X1 U818 ( .A(n1150), .B(n1151), .Z(n1147) );
XNOR2_X1 U819 ( .A(n1152), .B(n1153), .ZN(n1150) );
NOR2_X1 U820 ( .A1(G140), .A2(KEYINPUT56), .ZN(n1153) );
NAND2_X1 U821 ( .A1(n1142), .A2(n1080), .ZN(n1137) );
NAND2_X1 U822 ( .A1(n1154), .A2(n1155), .ZN(G69) );
NAND2_X1 U823 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U824 ( .A1(n1158), .A2(n1159), .ZN(n1154) );
NAND2_X1 U825 ( .A1(n1160), .A2(n1157), .ZN(n1159) );
NAND2_X1 U826 ( .A1(G953), .A2(n1161), .ZN(n1157) );
INV_X1 U827 ( .A(n1156), .ZN(n1158) );
XNOR2_X1 U828 ( .A(n1162), .B(n1163), .ZN(n1156) );
AND2_X1 U829 ( .A1(n1082), .A2(n1142), .ZN(n1163) );
NAND2_X1 U830 ( .A1(n1164), .A2(n1160), .ZN(n1162) );
INV_X1 U831 ( .A(n1165), .ZN(n1160) );
XOR2_X1 U832 ( .A(n1166), .B(n1167), .Z(n1164) );
NAND2_X1 U833 ( .A1(n1168), .A2(KEYINPUT44), .ZN(n1166) );
XNOR2_X1 U834 ( .A(n1169), .B(n1170), .ZN(n1168) );
NOR2_X1 U835 ( .A1(n1171), .A2(n1172), .ZN(G66) );
XOR2_X1 U836 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U837 ( .A1(n1175), .A2(n1176), .ZN(n1173) );
NOR2_X1 U838 ( .A1(n1171), .A2(n1177), .ZN(G63) );
XOR2_X1 U839 ( .A(n1178), .B(n1179), .Z(n1177) );
NOR2_X1 U840 ( .A1(n1180), .A2(n1176), .ZN(n1178) );
NOR2_X1 U841 ( .A1(n1171), .A2(n1181), .ZN(G60) );
NOR3_X1 U842 ( .A1(n1132), .A2(n1182), .A3(n1183), .ZN(n1181) );
NOR3_X1 U843 ( .A1(n1184), .A2(n1131), .A3(n1176), .ZN(n1183) );
NOR2_X1 U844 ( .A1(n1185), .A2(n1186), .ZN(n1182) );
NOR2_X1 U845 ( .A1(n1187), .A2(n1131), .ZN(n1185) );
NOR2_X1 U846 ( .A1(n1082), .A2(n1080), .ZN(n1187) );
XNOR2_X1 U847 ( .A(G104), .B(n1188), .ZN(G6) );
NOR2_X1 U848 ( .A1(n1171), .A2(n1189), .ZN(G57) );
XNOR2_X1 U849 ( .A(n1190), .B(n1191), .ZN(n1189) );
XOR2_X1 U850 ( .A(n1192), .B(KEYINPUT48), .Z(n1191) );
OR2_X1 U851 ( .A1(n1176), .A2(n1136), .ZN(n1192) );
NOR2_X1 U852 ( .A1(n1171), .A2(n1193), .ZN(G54) );
XOR2_X1 U853 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U854 ( .A(n1196), .B(n1197), .Z(n1195) );
NOR2_X1 U855 ( .A1(n1198), .A2(n1176), .ZN(n1196) );
XOR2_X1 U856 ( .A(n1199), .B(G140), .Z(n1194) );
NAND2_X1 U857 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND2_X1 U858 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XNOR2_X1 U859 ( .A(n1152), .B(KEYINPUT45), .ZN(n1203) );
XOR2_X1 U860 ( .A(n1204), .B(KEYINPUT30), .Z(n1202) );
XOR2_X1 U861 ( .A(KEYINPUT25), .B(n1205), .Z(n1200) );
NOR2_X1 U862 ( .A1(n1206), .A2(n1204), .ZN(n1205) );
NOR2_X1 U863 ( .A1(n1171), .A2(n1207), .ZN(G51) );
XOR2_X1 U864 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U865 ( .A(n1210), .B(n1211), .Z(n1209) );
NOR2_X1 U866 ( .A1(KEYINPUT49), .A2(n1212), .ZN(n1211) );
XNOR2_X1 U867 ( .A(n1213), .B(n1214), .ZN(n1208) );
NOR2_X1 U868 ( .A1(n1215), .A2(n1176), .ZN(n1214) );
NAND2_X1 U869 ( .A1(G902), .A2(n1216), .ZN(n1176) );
OR2_X1 U870 ( .A1(n1080), .A2(n1082), .ZN(n1216) );
NAND4_X1 U871 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1082) );
AND4_X1 U872 ( .A1(n1221), .A2(n1188), .A3(n1222), .A4(n1223), .ZN(n1220) );
INV_X1 U873 ( .A(n1072), .ZN(n1222) );
NOR3_X1 U874 ( .A1(n1224), .A2(n1092), .A3(n1225), .ZN(n1072) );
INV_X1 U875 ( .A(n1226), .ZN(n1092) );
NAND3_X1 U876 ( .A1(n1227), .A2(n1226), .A3(n1100), .ZN(n1188) );
NOR3_X1 U877 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1219) );
NOR4_X1 U878 ( .A1(n1231), .A2(n1232), .A3(n1225), .A4(n1101), .ZN(n1230) );
NAND3_X1 U879 ( .A1(n1088), .A2(n1233), .A3(n1234), .ZN(n1232) );
INV_X1 U880 ( .A(KEYINPUT28), .ZN(n1231) );
NOR2_X1 U881 ( .A1(KEYINPUT28), .A2(n1235), .ZN(n1229) );
NOR3_X1 U882 ( .A1(n1096), .A2(n1116), .A3(n1224), .ZN(n1228) );
INV_X1 U883 ( .A(n1236), .ZN(n1116) );
INV_X1 U884 ( .A(n1237), .ZN(n1096) );
NAND4_X1 U885 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1080) );
AND4_X1 U886 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1241) );
NAND2_X1 U887 ( .A1(n1246), .A2(n1247), .ZN(n1240) );
XNOR2_X1 U888 ( .A(KEYINPUT51), .B(n1225), .ZN(n1247) );
NAND3_X1 U889 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1238) );
NAND2_X1 U890 ( .A1(n1251), .A2(n1252), .ZN(n1249) );
NAND3_X1 U891 ( .A1(n1253), .A2(n1254), .A3(n1234), .ZN(n1252) );
NAND2_X1 U892 ( .A1(n1100), .A2(n1119), .ZN(n1251) );
NOR2_X1 U893 ( .A1(n1142), .A2(G952), .ZN(n1171) );
NAND2_X1 U894 ( .A1(n1255), .A2(n1256), .ZN(G48) );
NAND2_X1 U895 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XOR2_X1 U896 ( .A(KEYINPUT11), .B(n1259), .Z(n1255) );
NOR2_X1 U897 ( .A1(n1257), .A2(n1258), .ZN(n1259) );
INV_X1 U898 ( .A(n1239), .ZN(n1257) );
NAND2_X1 U899 ( .A1(n1246), .A2(n1100), .ZN(n1239) );
INV_X1 U900 ( .A(n1260), .ZN(n1246) );
XNOR2_X1 U901 ( .A(G143), .B(n1261), .ZN(G45) );
NAND4_X1 U902 ( .A1(n1250), .A2(n1234), .A3(n1262), .A4(n1263), .ZN(n1261) );
NOR3_X1 U903 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1263) );
XNOR2_X1 U904 ( .A(n1110), .B(KEYINPUT24), .ZN(n1262) );
XNOR2_X1 U905 ( .A(G140), .B(n1245), .ZN(G42) );
NAND3_X1 U906 ( .A1(n1100), .A2(n1236), .A3(n1267), .ZN(n1245) );
XNOR2_X1 U907 ( .A(G137), .B(n1244), .ZN(G39) );
NAND2_X1 U908 ( .A1(n1268), .A2(n1267), .ZN(n1244) );
XOR2_X1 U909 ( .A(G134), .B(n1269), .Z(G36) );
NOR2_X1 U910 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
AND2_X1 U911 ( .A1(KEYINPUT12), .A2(n1243), .ZN(n1271) );
NOR2_X1 U912 ( .A1(KEYINPUT33), .A2(n1243), .ZN(n1270) );
NAND3_X1 U913 ( .A1(n1267), .A2(n1099), .A3(n1250), .ZN(n1243) );
NAND2_X1 U914 ( .A1(n1272), .A2(n1273), .ZN(G33) );
NAND2_X1 U915 ( .A1(KEYINPUT32), .A2(n1274), .ZN(n1273) );
XOR2_X1 U916 ( .A(n1275), .B(n1276), .Z(n1272) );
NOR2_X1 U917 ( .A1(KEYINPUT32), .A2(n1274), .ZN(n1276) );
XNOR2_X1 U918 ( .A(n1277), .B(KEYINPUT19), .ZN(n1274) );
NAND3_X1 U919 ( .A1(n1267), .A2(n1100), .A3(n1278), .ZN(n1275) );
XNOR2_X1 U920 ( .A(n1250), .B(KEYINPUT55), .ZN(n1278) );
AND2_X1 U921 ( .A1(n1248), .A2(n1119), .ZN(n1267) );
INV_X1 U922 ( .A(n1098), .ZN(n1119) );
NAND2_X1 U923 ( .A1(n1279), .A2(n1114), .ZN(n1098) );
INV_X1 U924 ( .A(n1115), .ZN(n1279) );
XNOR2_X1 U925 ( .A(n1280), .B(n1281), .ZN(G30) );
NOR2_X1 U926 ( .A1(n1225), .A2(n1260), .ZN(n1281) );
NAND4_X1 U927 ( .A1(n1248), .A2(n1234), .A3(n1282), .A4(n1283), .ZN(n1260) );
NOR2_X1 U928 ( .A1(n1284), .A2(n1265), .ZN(n1248) );
INV_X1 U929 ( .A(n1099), .ZN(n1225) );
XNOR2_X1 U930 ( .A(G101), .B(n1221), .ZN(G3) );
NAND3_X1 U931 ( .A1(n1250), .A2(n1227), .A3(n1237), .ZN(n1221) );
XNOR2_X1 U932 ( .A(G125), .B(n1242), .ZN(G27) );
NAND3_X1 U933 ( .A1(n1100), .A2(n1236), .A3(n1285), .ZN(n1242) );
NOR3_X1 U934 ( .A1(n1095), .A2(n1265), .A3(n1088), .ZN(n1285) );
INV_X1 U935 ( .A(n1286), .ZN(n1088) );
AND2_X1 U936 ( .A1(n1084), .A2(n1287), .ZN(n1265) );
NAND4_X1 U937 ( .A1(G902), .A2(G953), .A3(n1288), .A4(n1143), .ZN(n1287) );
INV_X1 U938 ( .A(G900), .ZN(n1143) );
NAND2_X1 U939 ( .A1(n1289), .A2(n1290), .ZN(G24) );
NAND2_X1 U940 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
INV_X1 U941 ( .A(G122), .ZN(n1292) );
XNOR2_X1 U942 ( .A(KEYINPUT15), .B(n1217), .ZN(n1291) );
NAND2_X1 U943 ( .A1(G122), .A2(n1293), .ZN(n1289) );
XOR2_X1 U944 ( .A(n1217), .B(KEYINPUT42), .Z(n1293) );
NAND4_X1 U945 ( .A1(n1253), .A2(n1294), .A3(n1226), .A4(n1254), .ZN(n1217) );
NAND2_X1 U946 ( .A1(n1295), .A2(n1296), .ZN(n1226) );
OR3_X1 U947 ( .A1(n1283), .A2(n1282), .A3(KEYINPUT7), .ZN(n1296) );
NAND2_X1 U948 ( .A1(KEYINPUT7), .A2(n1236), .ZN(n1295) );
XNOR2_X1 U949 ( .A(G119), .B(n1218), .ZN(G21) );
NAND2_X1 U950 ( .A1(n1294), .A2(n1268), .ZN(n1218) );
AND3_X1 U951 ( .A1(n1282), .A2(n1283), .A3(n1237), .ZN(n1268) );
XOR2_X1 U952 ( .A(n1235), .B(n1297), .Z(G18) );
NAND2_X1 U953 ( .A1(n1298), .A2(KEYINPUT39), .ZN(n1297) );
XNOR2_X1 U954 ( .A(G116), .B(KEYINPUT22), .ZN(n1298) );
NAND3_X1 U955 ( .A1(n1250), .A2(n1099), .A3(n1294), .ZN(n1235) );
AND3_X1 U956 ( .A1(n1286), .A2(n1233), .A3(n1234), .ZN(n1294) );
NOR2_X1 U957 ( .A1(n1254), .A2(n1264), .ZN(n1099) );
XNOR2_X1 U958 ( .A(G113), .B(n1223), .ZN(G15) );
NAND4_X1 U959 ( .A1(n1250), .A2(n1100), .A3(n1299), .A4(n1286), .ZN(n1223) );
NAND2_X1 U960 ( .A1(n1300), .A2(n1301), .ZN(n1286) );
OR2_X1 U961 ( .A1(n1284), .A2(KEYINPUT47), .ZN(n1301) );
INV_X1 U962 ( .A(n1110), .ZN(n1284) );
NAND3_X1 U963 ( .A1(n1117), .A2(n1112), .A3(KEYINPUT47), .ZN(n1300) );
NOR2_X1 U964 ( .A1(n1253), .A2(n1266), .ZN(n1100) );
INV_X1 U965 ( .A(n1101), .ZN(n1250) );
NAND2_X1 U966 ( .A1(n1302), .A2(n1283), .ZN(n1101) );
XNOR2_X1 U967 ( .A(KEYINPUT7), .B(n1282), .ZN(n1302) );
XNOR2_X1 U968 ( .A(G110), .B(n1303), .ZN(G12) );
NAND4_X1 U969 ( .A1(KEYINPUT40), .A2(n1237), .A3(n1227), .A4(n1236), .ZN(n1303) );
NOR2_X1 U970 ( .A1(n1283), .A2(n1118), .ZN(n1236) );
INV_X1 U971 ( .A(n1282), .ZN(n1118) );
XOR2_X1 U972 ( .A(n1304), .B(n1175), .Z(n1282) );
NAND2_X1 U973 ( .A1(G217), .A2(n1305), .ZN(n1175) );
OR2_X1 U974 ( .A1(n1174), .A2(G902), .ZN(n1304) );
XNOR2_X1 U975 ( .A(n1306), .B(n1307), .ZN(n1174) );
XNOR2_X1 U976 ( .A(n1308), .B(n1309), .ZN(n1307) );
XNOR2_X1 U977 ( .A(n1258), .B(G137), .ZN(n1309) );
INV_X1 U978 ( .A(G146), .ZN(n1258) );
INV_X1 U979 ( .A(G110), .ZN(n1308) );
XOR2_X1 U980 ( .A(n1310), .B(n1311), .Z(n1306) );
XOR2_X1 U981 ( .A(n1312), .B(n1313), .Z(n1310) );
AND2_X1 U982 ( .A1(n1314), .A2(G221), .ZN(n1313) );
NAND2_X1 U983 ( .A1(n1315), .A2(n1316), .ZN(n1312) );
NAND2_X1 U984 ( .A1(G119), .A2(n1280), .ZN(n1316) );
XOR2_X1 U985 ( .A(KEYINPUT4), .B(n1317), .Z(n1315) );
NOR2_X1 U986 ( .A1(G119), .A2(n1280), .ZN(n1317) );
NAND3_X1 U987 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1283) );
OR2_X1 U988 ( .A1(n1321), .A2(n1133), .ZN(n1320) );
NAND3_X1 U989 ( .A1(n1133), .A2(n1321), .A3(G472), .ZN(n1319) );
NAND2_X1 U990 ( .A1(n1322), .A2(n1136), .ZN(n1318) );
INV_X1 U991 ( .A(G472), .ZN(n1136) );
NAND2_X1 U992 ( .A1(n1323), .A2(n1321), .ZN(n1322) );
INV_X1 U993 ( .A(KEYINPUT59), .ZN(n1321) );
XNOR2_X1 U994 ( .A(KEYINPUT9), .B(n1133), .ZN(n1323) );
NAND2_X1 U995 ( .A1(n1324), .A2(n1190), .ZN(n1133) );
XNOR2_X1 U996 ( .A(n1325), .B(n1326), .ZN(n1190) );
XOR2_X1 U997 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U998 ( .A(n1152), .B(n1329), .ZN(n1328) );
AND2_X1 U999 ( .A1(n1330), .A2(G210), .ZN(n1329) );
XNOR2_X1 U1000 ( .A(n1331), .B(n1332), .ZN(n1325) );
XNOR2_X1 U1001 ( .A(G101), .B(G113), .ZN(n1331) );
XNOR2_X1 U1002 ( .A(KEYINPUT37), .B(n1333), .ZN(n1324) );
INV_X1 U1003 ( .A(n1224), .ZN(n1227) );
NAND2_X1 U1004 ( .A1(n1110), .A2(n1299), .ZN(n1224) );
AND2_X1 U1005 ( .A1(n1334), .A2(n1233), .ZN(n1299) );
NAND2_X1 U1006 ( .A1(n1084), .A2(n1335), .ZN(n1233) );
NAND3_X1 U1007 ( .A1(n1165), .A2(n1288), .A3(G902), .ZN(n1335) );
NOR2_X1 U1008 ( .A1(G898), .A2(n1142), .ZN(n1165) );
NAND3_X1 U1009 ( .A1(n1288), .A2(n1142), .A3(G952), .ZN(n1084) );
NAND2_X1 U1010 ( .A1(G237), .A2(G234), .ZN(n1288) );
XNOR2_X1 U1011 ( .A(n1234), .B(KEYINPUT8), .ZN(n1334) );
INV_X1 U1012 ( .A(n1095), .ZN(n1234) );
NAND2_X1 U1013 ( .A1(n1115), .A2(n1114), .ZN(n1095) );
NAND2_X1 U1014 ( .A1(G214), .A2(n1336), .ZN(n1114) );
XOR2_X1 U1015 ( .A(n1337), .B(n1215), .Z(n1115) );
NAND2_X1 U1016 ( .A1(G210), .A2(n1336), .ZN(n1215) );
NAND2_X1 U1017 ( .A1(n1338), .A2(n1333), .ZN(n1336) );
INV_X1 U1018 ( .A(G237), .ZN(n1338) );
NAND2_X1 U1019 ( .A1(n1339), .A2(n1333), .ZN(n1337) );
XOR2_X1 U1020 ( .A(n1340), .B(n1341), .Z(n1339) );
XNOR2_X1 U1021 ( .A(n1213), .B(n1210), .ZN(n1341) );
XOR2_X1 U1022 ( .A(n1342), .B(n1343), .Z(n1210) );
NOR2_X1 U1023 ( .A1(G953), .A2(n1161), .ZN(n1343) );
INV_X1 U1024 ( .A(G224), .ZN(n1161) );
NAND2_X1 U1025 ( .A1(n1344), .A2(n1345), .ZN(n1342) );
NAND3_X1 U1026 ( .A1(n1346), .A2(n1169), .A3(KEYINPUT38), .ZN(n1345) );
XOR2_X1 U1027 ( .A(n1347), .B(n1348), .Z(n1346) );
NAND2_X1 U1028 ( .A1(n1349), .A2(n1350), .ZN(n1347) );
OR2_X1 U1029 ( .A1(n1170), .A2(KEYINPUT5), .ZN(n1350) );
OR2_X1 U1030 ( .A1(n1351), .A2(KEYINPUT60), .ZN(n1349) );
NAND2_X1 U1031 ( .A1(n1352), .A2(n1353), .ZN(n1344) );
NAND2_X1 U1032 ( .A1(KEYINPUT38), .A2(n1169), .ZN(n1353) );
NAND2_X1 U1033 ( .A1(n1354), .A2(n1355), .ZN(n1169) );
NAND2_X1 U1034 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
XOR2_X1 U1035 ( .A(KEYINPUT10), .B(n1358), .Z(n1354) );
NOR2_X1 U1036 ( .A1(n1357), .A2(n1356), .ZN(n1358) );
NAND2_X1 U1037 ( .A1(n1359), .A2(n1360), .ZN(n1356) );
NAND2_X1 U1038 ( .A1(KEYINPUT62), .A2(n1327), .ZN(n1360) );
XOR2_X1 U1039 ( .A(G119), .B(n1361), .Z(n1327) );
OR3_X1 U1040 ( .A1(n1361), .A2(G119), .A3(KEYINPUT62), .ZN(n1359) );
XNOR2_X1 U1041 ( .A(G116), .B(KEYINPUT50), .ZN(n1361) );
XNOR2_X1 U1042 ( .A(n1362), .B(n1348), .ZN(n1352) );
XNOR2_X1 U1043 ( .A(n1167), .B(KEYINPUT31), .ZN(n1348) );
XNOR2_X1 U1044 ( .A(G110), .B(n1363), .ZN(n1167) );
NAND2_X1 U1045 ( .A1(n1364), .A2(n1365), .ZN(n1362) );
NAND2_X1 U1046 ( .A1(n1170), .A2(KEYINPUT5), .ZN(n1365) );
INV_X1 U1047 ( .A(n1351), .ZN(n1170) );
NAND2_X1 U1048 ( .A1(n1351), .A2(KEYINPUT60), .ZN(n1364) );
XNOR2_X1 U1049 ( .A(n1366), .B(G101), .ZN(n1351) );
NAND2_X1 U1050 ( .A1(KEYINPUT6), .A2(n1367), .ZN(n1366) );
INV_X1 U1051 ( .A(n1332), .ZN(n1213) );
NAND2_X1 U1052 ( .A1(n1368), .A2(n1369), .ZN(n1332) );
NAND2_X1 U1053 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
XOR2_X1 U1054 ( .A(n1372), .B(KEYINPUT35), .Z(n1370) );
XOR2_X1 U1055 ( .A(KEYINPUT58), .B(n1373), .Z(n1368) );
NOR2_X1 U1056 ( .A1(n1372), .A2(n1374), .ZN(n1373) );
XOR2_X1 U1057 ( .A(n1371), .B(KEYINPUT3), .Z(n1374) );
XNOR2_X1 U1058 ( .A(KEYINPUT18), .B(n1212), .ZN(n1340) );
NOR2_X1 U1059 ( .A1(n1117), .A2(n1121), .ZN(n1110) );
INV_X1 U1060 ( .A(n1112), .ZN(n1121) );
NAND2_X1 U1061 ( .A1(G221), .A2(n1305), .ZN(n1112) );
NAND2_X1 U1062 ( .A1(G234), .A2(n1333), .ZN(n1305) );
INV_X1 U1063 ( .A(n1113), .ZN(n1117) );
XNOR2_X1 U1064 ( .A(n1375), .B(n1376), .ZN(n1113) );
XNOR2_X1 U1065 ( .A(KEYINPUT21), .B(n1198), .ZN(n1376) );
INV_X1 U1066 ( .A(G469), .ZN(n1198) );
NAND2_X1 U1067 ( .A1(n1377), .A2(n1333), .ZN(n1375) );
INV_X1 U1068 ( .A(G902), .ZN(n1333) );
XOR2_X1 U1069 ( .A(n1378), .B(n1379), .Z(n1377) );
XNOR2_X1 U1070 ( .A(n1204), .B(n1197), .ZN(n1379) );
XOR2_X1 U1071 ( .A(G110), .B(n1380), .Z(n1197) );
AND2_X1 U1072 ( .A1(n1142), .A2(G227), .ZN(n1380) );
XOR2_X1 U1073 ( .A(n1381), .B(n1382), .Z(n1204) );
XOR2_X1 U1074 ( .A(KEYINPUT26), .B(G101), .Z(n1382) );
XNOR2_X1 U1075 ( .A(n1367), .B(n1151), .ZN(n1381) );
XOR2_X1 U1076 ( .A(n1371), .B(n1372), .Z(n1151) );
XOR2_X1 U1077 ( .A(n1383), .B(G146), .Z(n1372) );
XNOR2_X1 U1078 ( .A(G128), .B(KEYINPUT41), .ZN(n1371) );
XNOR2_X1 U1079 ( .A(G104), .B(n1073), .ZN(n1367) );
INV_X1 U1080 ( .A(G107), .ZN(n1073) );
XNOR2_X1 U1081 ( .A(n1206), .B(n1384), .ZN(n1378) );
XOR2_X1 U1082 ( .A(KEYINPUT2), .B(n1385), .Z(n1384) );
NOR2_X1 U1083 ( .A1(G140), .A2(KEYINPUT43), .ZN(n1385) );
INV_X1 U1084 ( .A(n1152), .ZN(n1206) );
XOR2_X1 U1085 ( .A(G131), .B(n1386), .Z(n1152) );
XOR2_X1 U1086 ( .A(G137), .B(G134), .Z(n1386) );
NOR2_X1 U1087 ( .A1(n1254), .A2(n1253), .ZN(n1237) );
INV_X1 U1088 ( .A(n1264), .ZN(n1253) );
XOR2_X1 U1089 ( .A(n1124), .B(KEYINPUT46), .Z(n1264) );
XOR2_X1 U1090 ( .A(n1387), .B(n1180), .Z(n1124) );
INV_X1 U1091 ( .A(G478), .ZN(n1180) );
OR2_X1 U1092 ( .A1(n1179), .A2(G902), .ZN(n1387) );
XNOR2_X1 U1093 ( .A(n1388), .B(n1389), .ZN(n1179) );
NOR3_X1 U1094 ( .A1(n1390), .A2(KEYINPUT53), .A3(n1391), .ZN(n1389) );
NOR2_X1 U1095 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
XOR2_X1 U1096 ( .A(n1394), .B(KEYINPUT36), .Z(n1390) );
NAND2_X1 U1097 ( .A1(n1392), .A2(n1393), .ZN(n1394) );
XNOR2_X1 U1098 ( .A(n1280), .B(n1395), .ZN(n1393) );
XNOR2_X1 U1099 ( .A(n1383), .B(G134), .ZN(n1395) );
INV_X1 U1100 ( .A(G143), .ZN(n1383) );
INV_X1 U1101 ( .A(G128), .ZN(n1280) );
XOR2_X1 U1102 ( .A(n1363), .B(n1396), .Z(n1392) );
XOR2_X1 U1103 ( .A(G116), .B(n1397), .Z(n1396) );
NOR2_X1 U1104 ( .A1(G107), .A2(KEYINPUT17), .ZN(n1397) );
NAND2_X1 U1105 ( .A1(G217), .A2(n1314), .ZN(n1388) );
AND2_X1 U1106 ( .A1(G234), .A2(n1142), .ZN(n1314) );
INV_X1 U1107 ( .A(G953), .ZN(n1142) );
INV_X1 U1108 ( .A(n1266), .ZN(n1254) );
XOR2_X1 U1109 ( .A(n1132), .B(n1131), .Z(n1266) );
INV_X1 U1110 ( .A(G475), .ZN(n1131) );
NOR2_X1 U1111 ( .A1(n1186), .A2(G902), .ZN(n1132) );
INV_X1 U1112 ( .A(n1184), .ZN(n1186) );
XNOR2_X1 U1113 ( .A(n1398), .B(n1399), .ZN(n1184) );
XNOR2_X1 U1114 ( .A(n1400), .B(n1363), .ZN(n1399) );
XOR2_X1 U1115 ( .A(G122), .B(KEYINPUT34), .Z(n1363) );
NAND2_X1 U1116 ( .A1(n1401), .A2(n1402), .ZN(n1400) );
NAND2_X1 U1117 ( .A1(G146), .A2(n1311), .ZN(n1402) );
XOR2_X1 U1118 ( .A(KEYINPUT16), .B(n1403), .Z(n1401) );
NOR2_X1 U1119 ( .A1(G146), .A2(n1311), .ZN(n1403) );
XNOR2_X1 U1120 ( .A(n1212), .B(G140), .ZN(n1311) );
INV_X1 U1121 ( .A(G125), .ZN(n1212) );
XOR2_X1 U1122 ( .A(n1404), .B(n1405), .Z(n1398) );
XNOR2_X1 U1123 ( .A(n1357), .B(G104), .ZN(n1405) );
INV_X1 U1124 ( .A(G113), .ZN(n1357) );
NAND3_X1 U1125 ( .A1(n1406), .A2(n1407), .A3(n1408), .ZN(n1404) );
NAND2_X1 U1126 ( .A1(KEYINPUT63), .A2(n1409), .ZN(n1408) );
NAND3_X1 U1127 ( .A1(n1410), .A2(n1411), .A3(n1277), .ZN(n1407) );
INV_X1 U1128 ( .A(KEYINPUT63), .ZN(n1411) );
OR2_X1 U1129 ( .A1(n1277), .A2(n1410), .ZN(n1406) );
NOR2_X1 U1130 ( .A1(KEYINPUT57), .A2(n1409), .ZN(n1410) );
XNOR2_X1 U1131 ( .A(n1412), .B(G143), .ZN(n1409) );
NAND2_X1 U1132 ( .A1(G214), .A2(n1330), .ZN(n1412) );
NOR2_X1 U1133 ( .A1(G953), .A2(G237), .ZN(n1330) );
INV_X1 U1134 ( .A(G131), .ZN(n1277) );
endmodule


