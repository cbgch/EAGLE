//Key = 0100000110110110110001001000011110011000010101101011010110110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
n1441, n1442, n1443;

XOR2_X1 U786 ( .A(n1091), .B(n1092), .Z(G9) );
NAND4_X1 U787 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(G75) );
NAND4_X1 U788 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1095) );
NAND2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND3_X1 U790 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1101) );
INV_X1 U791 ( .A(KEYINPUT10), .ZN(n1104) );
NAND3_X1 U792 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1099) );
NAND2_X1 U793 ( .A1(n1105), .A2(n1109), .ZN(n1107) );
NAND2_X1 U794 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U795 ( .A1(KEYINPUT10), .A2(n1103), .ZN(n1111) );
NAND2_X1 U796 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NAND2_X1 U797 ( .A1(n1114), .A2(n1115), .ZN(n1106) );
NAND2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U799 ( .A(KEYINPUT46), .B(n1118), .Z(n1116) );
NAND2_X1 U800 ( .A1(n1105), .A2(n1119), .ZN(n1094) );
NAND2_X1 U801 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND3_X1 U802 ( .A1(n1114), .A2(n1122), .A3(n1097), .ZN(n1121) );
INV_X1 U803 ( .A(n1123), .ZN(n1097) );
NAND2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
NAND2_X1 U805 ( .A1(n1098), .A2(n1126), .ZN(n1125) );
NAND2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U807 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U808 ( .A1(n1108), .A2(n1131), .ZN(n1124) );
NAND2_X1 U809 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XOR2_X1 U810 ( .A(KEYINPUT53), .B(n1134), .Z(n1132) );
NAND4_X1 U811 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1114), .ZN(n1120) );
NOR2_X1 U812 ( .A1(n1129), .A2(n1138), .ZN(n1137) );
XOR2_X1 U813 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U814 ( .A1(n1141), .A2(KEYINPUT60), .ZN(n1140) );
INV_X1 U815 ( .A(n1142), .ZN(n1141) );
XNOR2_X1 U816 ( .A(n1143), .B(n1144), .ZN(n1136) );
NOR2_X1 U817 ( .A1(KEYINPUT42), .A2(n1145), .ZN(n1144) );
XOR2_X1 U818 ( .A(n1146), .B(KEYINPUT25), .Z(n1135) );
XOR2_X1 U819 ( .A(n1147), .B(n1148), .Z(G72) );
NOR2_X1 U820 ( .A1(n1149), .A2(n1096), .ZN(n1148) );
NOR2_X1 U821 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND2_X1 U822 ( .A1(n1152), .A2(n1153), .ZN(n1147) );
NAND3_X1 U823 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1153) );
NAND2_X1 U824 ( .A1(G953), .A2(n1151), .ZN(n1155) );
XOR2_X1 U825 ( .A(n1157), .B(KEYINPUT56), .Z(n1154) );
NAND3_X1 U826 ( .A1(n1157), .A2(n1096), .A3(n1158), .ZN(n1152) );
INV_X1 U827 ( .A(n1156), .ZN(n1158) );
XOR2_X1 U828 ( .A(n1159), .B(n1160), .Z(n1156) );
XOR2_X1 U829 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U830 ( .A(KEYINPUT54), .B(KEYINPUT0), .ZN(n1162) );
NAND2_X1 U831 ( .A1(KEYINPUT17), .A2(n1163), .ZN(n1161) );
XOR2_X1 U832 ( .A(n1164), .B(n1165), .Z(n1159) );
XOR2_X1 U833 ( .A(n1166), .B(n1167), .Z(G69) );
XOR2_X1 U834 ( .A(n1168), .B(n1169), .Z(n1167) );
AND2_X1 U835 ( .A1(n1170), .A2(n1096), .ZN(n1169) );
NOR2_X1 U836 ( .A1(n1171), .A2(n1172), .ZN(n1168) );
XNOR2_X1 U837 ( .A(n1173), .B(n1174), .ZN(n1172) );
NAND2_X1 U838 ( .A1(KEYINPUT61), .A2(n1175), .ZN(n1173) );
NOR2_X1 U839 ( .A1(n1096), .A2(n1176), .ZN(n1171) );
XOR2_X1 U840 ( .A(KEYINPUT57), .B(G898), .Z(n1176) );
NOR3_X1 U841 ( .A1(n1096), .A2(KEYINPUT19), .A3(n1177), .ZN(n1166) );
AND2_X1 U842 ( .A1(G898), .A2(G224), .ZN(n1177) );
NOR2_X1 U843 ( .A1(n1178), .A2(n1179), .ZN(G66) );
NOR3_X1 U844 ( .A1(n1143), .A2(n1180), .A3(n1181), .ZN(n1179) );
AND4_X1 U845 ( .A1(n1182), .A2(KEYINPUT16), .A3(n1183), .A4(n1184), .ZN(n1181) );
INV_X1 U846 ( .A(n1145), .ZN(n1183) );
NOR2_X1 U847 ( .A1(n1185), .A2(n1182), .ZN(n1180) );
NOR3_X1 U848 ( .A1(n1186), .A2(n1093), .A3(n1145), .ZN(n1185) );
INV_X1 U849 ( .A(KEYINPUT16), .ZN(n1186) );
NOR2_X1 U850 ( .A1(n1178), .A2(n1187), .ZN(G63) );
XOR2_X1 U851 ( .A(n1188), .B(n1189), .Z(n1187) );
NOR2_X1 U852 ( .A1(KEYINPUT27), .A2(n1190), .ZN(n1189) );
XNOR2_X1 U853 ( .A(n1191), .B(KEYINPUT15), .ZN(n1190) );
NAND2_X1 U854 ( .A1(n1184), .A2(G478), .ZN(n1188) );
NOR2_X1 U855 ( .A1(n1178), .A2(n1192), .ZN(G60) );
XOR2_X1 U856 ( .A(n1193), .B(n1194), .Z(n1192) );
AND2_X1 U857 ( .A1(G475), .A2(n1184), .ZN(n1193) );
NAND2_X1 U858 ( .A1(n1195), .A2(n1196), .ZN(G6) );
OR2_X1 U859 ( .A1(n1197), .A2(G104), .ZN(n1196) );
NAND2_X1 U860 ( .A1(n1198), .A2(G104), .ZN(n1195) );
NAND2_X1 U861 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND2_X1 U862 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
INV_X1 U863 ( .A(KEYINPUT21), .ZN(n1202) );
NAND2_X1 U864 ( .A1(KEYINPUT21), .A2(n1197), .ZN(n1199) );
NAND2_X1 U865 ( .A1(KEYINPUT35), .A2(n1201), .ZN(n1197) );
NOR2_X1 U866 ( .A1(n1178), .A2(n1203), .ZN(G57) );
XOR2_X1 U867 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U868 ( .A(n1206), .B(n1207), .Z(n1205) );
AND2_X1 U869 ( .A1(G472), .A2(n1184), .ZN(n1206) );
NAND2_X1 U870 ( .A1(n1208), .A2(n1209), .ZN(n1204) );
NAND2_X1 U871 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND2_X1 U872 ( .A1(n1212), .A2(n1213), .ZN(n1208) );
XOR2_X1 U873 ( .A(n1214), .B(n1215), .Z(n1212) );
XOR2_X1 U874 ( .A(n1216), .B(n1217), .Z(n1215) );
NOR2_X1 U875 ( .A1(n1178), .A2(n1218), .ZN(G54) );
XOR2_X1 U876 ( .A(n1219), .B(n1220), .Z(n1218) );
NOR2_X1 U877 ( .A1(KEYINPUT49), .A2(n1221), .ZN(n1220) );
XOR2_X1 U878 ( .A(n1222), .B(n1223), .Z(n1221) );
XNOR2_X1 U879 ( .A(n1224), .B(n1225), .ZN(n1223) );
XOR2_X1 U880 ( .A(n1226), .B(n1227), .Z(n1222) );
XOR2_X1 U881 ( .A(KEYINPUT3), .B(G140), .Z(n1227) );
NAND2_X1 U882 ( .A1(n1184), .A2(G469), .ZN(n1219) );
NOR2_X1 U883 ( .A1(n1178), .A2(n1228), .ZN(G51) );
XOR2_X1 U884 ( .A(n1229), .B(n1230), .Z(n1228) );
NAND2_X1 U885 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND2_X1 U886 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
XOR2_X1 U887 ( .A(KEYINPUT1), .B(n1235), .Z(n1231) );
NOR2_X1 U888 ( .A1(n1233), .A2(n1234), .ZN(n1235) );
AND3_X1 U889 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1233) );
NAND2_X1 U890 ( .A1(n1239), .A2(n1240), .ZN(n1237) );
XOR2_X1 U891 ( .A(n1241), .B(n1242), .Z(n1239) );
NAND2_X1 U892 ( .A1(KEYINPUT41), .A2(n1243), .ZN(n1241) );
NAND3_X1 U893 ( .A1(n1244), .A2(n1243), .A3(n1245), .ZN(n1236) );
XOR2_X1 U894 ( .A(KEYINPUT41), .B(n1242), .Z(n1244) );
NAND3_X1 U895 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1229) );
OR2_X1 U896 ( .A1(n1184), .A2(KEYINPUT28), .ZN(n1247) );
NOR2_X1 U897 ( .A1(n1249), .A2(n1093), .ZN(n1184) );
NAND2_X1 U898 ( .A1(KEYINPUT28), .A2(n1250), .ZN(n1246) );
NAND2_X1 U899 ( .A1(n1093), .A2(G902), .ZN(n1250) );
NOR2_X1 U900 ( .A1(n1170), .A2(n1157), .ZN(n1093) );
NAND4_X1 U901 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1157) );
NOR4_X1 U902 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1254) );
NOR3_X1 U903 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1253) );
NOR4_X1 U904 ( .A1(n1262), .A2(n1263), .A3(n1134), .A4(n1117), .ZN(n1261) );
AND2_X1 U905 ( .A1(n1262), .A2(n1264), .ZN(n1260) );
INV_X1 U906 ( .A(KEYINPUT4), .ZN(n1262) );
INV_X1 U907 ( .A(n1265), .ZN(n1259) );
NAND4_X1 U908 ( .A1(n1266), .A2(n1267), .A3(n1268), .A4(n1269), .ZN(n1170) );
NOR4_X1 U909 ( .A1(n1270), .A2(n1201), .A3(n1271), .A4(n1272), .ZN(n1269) );
INV_X1 U910 ( .A(n1273), .ZN(n1272) );
INV_X1 U911 ( .A(n1092), .ZN(n1271) );
NAND4_X1 U912 ( .A1(n1118), .A2(n1274), .A3(n1098), .A4(n1275), .ZN(n1092) );
AND4_X1 U913 ( .A1(n1276), .A2(n1274), .A3(n1098), .A4(n1275), .ZN(n1201) );
NAND2_X1 U914 ( .A1(n1276), .A2(n1277), .ZN(n1268) );
NAND4_X1 U915 ( .A1(n1278), .A2(n1279), .A3(n1280), .A4(n1098), .ZN(n1267) );
NAND2_X1 U916 ( .A1(n1281), .A2(n1282), .ZN(n1266) );
NAND2_X1 U917 ( .A1(n1283), .A2(n1133), .ZN(n1282) );
INV_X1 U918 ( .A(n1284), .ZN(n1281) );
NOR2_X1 U919 ( .A1(n1096), .A2(G952), .ZN(n1178) );
XOR2_X1 U920 ( .A(n1285), .B(n1265), .Z(G48) );
NAND2_X1 U921 ( .A1(n1286), .A2(n1276), .ZN(n1265) );
XOR2_X1 U922 ( .A(n1287), .B(n1251), .Z(G45) );
NAND3_X1 U923 ( .A1(n1274), .A2(n1288), .A3(n1289), .ZN(n1251) );
NOR3_X1 U924 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1289) );
XOR2_X1 U925 ( .A(n1293), .B(n1264), .Z(G42) );
NOR3_X1 U926 ( .A1(n1283), .A2(n1117), .A3(n1263), .ZN(n1264) );
XOR2_X1 U927 ( .A(n1294), .B(KEYINPUT32), .Z(n1293) );
XNOR2_X1 U928 ( .A(G137), .B(n1252), .ZN(G39) );
NAND3_X1 U929 ( .A1(n1105), .A2(n1295), .A3(n1296), .ZN(n1252) );
XOR2_X1 U930 ( .A(G134), .B(n1258), .Z(G36) );
AND3_X1 U931 ( .A1(n1118), .A2(n1288), .A3(n1296), .ZN(n1258) );
INV_X1 U932 ( .A(n1263), .ZN(n1296) );
XOR2_X1 U933 ( .A(G131), .B(n1257), .Z(G33) );
NOR3_X1 U934 ( .A1(n1117), .A2(n1133), .A3(n1263), .ZN(n1257) );
NAND3_X1 U935 ( .A1(n1103), .A2(n1297), .A3(n1108), .ZN(n1263) );
INV_X1 U936 ( .A(n1102), .ZN(n1108) );
NAND2_X1 U937 ( .A1(n1130), .A2(n1298), .ZN(n1102) );
XOR2_X1 U938 ( .A(G128), .B(n1256), .Z(G30) );
AND2_X1 U939 ( .A1(n1286), .A2(n1118), .ZN(n1256) );
AND3_X1 U940 ( .A1(n1295), .A2(n1297), .A3(n1274), .ZN(n1286) );
XOR2_X1 U941 ( .A(n1299), .B(n1300), .Z(G3) );
XOR2_X1 U942 ( .A(KEYINPUT34), .B(G101), .Z(n1300) );
NOR2_X1 U943 ( .A1(n1301), .A2(n1284), .ZN(n1299) );
XOR2_X1 U944 ( .A(n1133), .B(KEYINPUT9), .Z(n1301) );
XOR2_X1 U945 ( .A(G125), .B(n1255), .Z(G27) );
AND4_X1 U946 ( .A1(n1134), .A2(n1276), .A3(n1302), .A4(n1114), .ZN(n1255) );
NOR2_X1 U947 ( .A1(n1291), .A2(n1127), .ZN(n1302) );
INV_X1 U948 ( .A(n1303), .ZN(n1127) );
INV_X1 U949 ( .A(n1297), .ZN(n1291) );
NAND2_X1 U950 ( .A1(n1123), .A2(n1304), .ZN(n1297) );
NAND4_X1 U951 ( .A1(G953), .A2(G902), .A3(n1305), .A4(n1151), .ZN(n1304) );
INV_X1 U952 ( .A(G900), .ZN(n1151) );
NAND2_X1 U953 ( .A1(n1306), .A2(n1307), .ZN(G24) );
NAND2_X1 U954 ( .A1(G122), .A2(n1308), .ZN(n1307) );
XOR2_X1 U955 ( .A(n1309), .B(KEYINPUT5), .Z(n1306) );
OR2_X1 U956 ( .A1(n1308), .A2(G122), .ZN(n1309) );
NAND2_X1 U957 ( .A1(n1303), .A2(n1310), .ZN(n1308) );
XOR2_X1 U958 ( .A(KEYINPUT37), .B(n1311), .Z(n1310) );
NOR3_X1 U959 ( .A1(n1312), .A2(n1290), .A3(n1313), .ZN(n1311) );
XNOR2_X1 U960 ( .A(n1114), .B(KEYINPUT40), .ZN(n1313) );
NAND3_X1 U961 ( .A1(n1098), .A2(n1275), .A3(n1280), .ZN(n1312) );
NAND2_X1 U962 ( .A1(n1314), .A2(n1315), .ZN(n1098) );
OR2_X1 U963 ( .A1(n1133), .A2(KEYINPUT55), .ZN(n1315) );
NAND3_X1 U964 ( .A1(n1146), .A2(n1316), .A3(KEYINPUT55), .ZN(n1314) );
XOR2_X1 U965 ( .A(n1317), .B(n1273), .Z(G21) );
NAND3_X1 U966 ( .A1(n1278), .A2(n1295), .A3(n1105), .ZN(n1273) );
NAND2_X1 U967 ( .A1(n1318), .A2(n1319), .ZN(n1295) );
OR3_X1 U968 ( .A1(n1316), .A2(n1146), .A3(KEYINPUT20), .ZN(n1319) );
NAND2_X1 U969 ( .A1(KEYINPUT20), .A2(n1288), .ZN(n1318) );
XOR2_X1 U970 ( .A(n1320), .B(n1270), .Z(G18) );
AND2_X1 U971 ( .A1(n1277), .A2(n1118), .ZN(n1270) );
NOR2_X1 U972 ( .A1(n1279), .A2(n1292), .ZN(n1118) );
NAND2_X1 U973 ( .A1(KEYINPUT24), .A2(n1321), .ZN(n1320) );
NAND2_X1 U974 ( .A1(n1322), .A2(n1323), .ZN(G15) );
OR2_X1 U975 ( .A1(n1324), .A2(G113), .ZN(n1323) );
NAND2_X1 U976 ( .A1(G113), .A2(n1325), .ZN(n1322) );
NAND2_X1 U977 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
NAND2_X1 U978 ( .A1(KEYINPUT7), .A2(n1324), .ZN(n1327) );
NAND3_X1 U979 ( .A1(n1277), .A2(n1328), .A3(n1276), .ZN(n1324) );
XOR2_X1 U980 ( .A(KEYINPUT8), .B(KEYINPUT23), .Z(n1328) );
NAND3_X1 U981 ( .A1(n1276), .A2(n1277), .A3(n1329), .ZN(n1326) );
INV_X1 U982 ( .A(KEYINPUT7), .ZN(n1329) );
AND2_X1 U983 ( .A1(n1278), .A2(n1288), .ZN(n1277) );
INV_X1 U984 ( .A(n1133), .ZN(n1288) );
NAND2_X1 U985 ( .A1(n1316), .A2(n1330), .ZN(n1133) );
INV_X1 U986 ( .A(n1146), .ZN(n1330) );
AND3_X1 U987 ( .A1(n1303), .A2(n1275), .A3(n1114), .ZN(n1278) );
AND2_X1 U988 ( .A1(n1113), .A2(n1331), .ZN(n1114) );
INV_X1 U989 ( .A(n1117), .ZN(n1276) );
NAND2_X1 U990 ( .A1(n1292), .A2(n1279), .ZN(n1117) );
XOR2_X1 U991 ( .A(G110), .B(n1332), .Z(G12) );
NOR2_X1 U992 ( .A1(n1284), .A2(n1283), .ZN(n1332) );
INV_X1 U993 ( .A(n1134), .ZN(n1283) );
NOR2_X1 U994 ( .A1(n1333), .A2(n1316), .ZN(n1134) );
XOR2_X1 U995 ( .A(n1145), .B(n1143), .Z(n1316) );
NOR2_X1 U996 ( .A1(n1182), .A2(G902), .ZN(n1143) );
NAND3_X1 U997 ( .A1(n1334), .A2(n1335), .A3(n1336), .ZN(n1182) );
NAND2_X1 U998 ( .A1(KEYINPUT2), .A2(n1337), .ZN(n1336) );
OR3_X1 U999 ( .A1(n1338), .A2(KEYINPUT2), .A3(n1339), .ZN(n1335) );
NAND2_X1 U1000 ( .A1(n1339), .A2(n1338), .ZN(n1334) );
NAND2_X1 U1001 ( .A1(KEYINPUT30), .A2(n1340), .ZN(n1338) );
INV_X1 U1002 ( .A(n1337), .ZN(n1340) );
XOR2_X1 U1003 ( .A(n1341), .B(n1342), .Z(n1337) );
NOR2_X1 U1004 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
XOR2_X1 U1005 ( .A(n1345), .B(KEYINPUT59), .Z(n1344) );
NAND2_X1 U1006 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
NOR2_X1 U1007 ( .A1(n1346), .A2(n1347), .ZN(n1343) );
XOR2_X1 U1008 ( .A(n1317), .B(G128), .Z(n1346) );
NAND2_X1 U1009 ( .A1(n1348), .A2(n1349), .ZN(n1341) );
NAND2_X1 U1010 ( .A1(n1163), .A2(n1285), .ZN(n1349) );
XOR2_X1 U1011 ( .A(n1350), .B(KEYINPUT22), .Z(n1348) );
OR2_X1 U1012 ( .A1(n1163), .A2(n1285), .ZN(n1350) );
XNOR2_X1 U1013 ( .A(n1351), .B(n1352), .ZN(n1339) );
XOR2_X1 U1014 ( .A(KEYINPUT36), .B(G137), .Z(n1352) );
NAND2_X1 U1015 ( .A1(G221), .A2(n1353), .ZN(n1351) );
NAND2_X1 U1016 ( .A1(G217), .A2(n1354), .ZN(n1145) );
XOR2_X1 U1017 ( .A(KEYINPUT55), .B(n1146), .Z(n1333) );
XOR2_X1 U1018 ( .A(n1355), .B(G472), .Z(n1146) );
NAND2_X1 U1019 ( .A1(n1356), .A2(n1249), .ZN(n1355) );
XNOR2_X1 U1020 ( .A(n1357), .B(n1207), .ZN(n1356) );
XNOR2_X1 U1021 ( .A(n1358), .B(G101), .ZN(n1207) );
NAND2_X1 U1022 ( .A1(G210), .A2(n1359), .ZN(n1358) );
NAND2_X1 U1023 ( .A1(n1360), .A2(n1361), .ZN(n1357) );
NAND2_X1 U1024 ( .A1(n1211), .A2(n1362), .ZN(n1361) );
NAND2_X1 U1025 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
OR2_X1 U1026 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
XOR2_X1 U1027 ( .A(n1367), .B(KEYINPUT52), .Z(n1363) );
NAND2_X1 U1028 ( .A1(n1365), .A2(n1366), .ZN(n1367) );
NAND2_X1 U1029 ( .A1(n1213), .A2(n1368), .ZN(n1360) );
NAND2_X1 U1030 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
OR2_X1 U1031 ( .A1(n1210), .A2(KEYINPUT52), .ZN(n1370) );
XOR2_X1 U1032 ( .A(n1242), .B(n1365), .Z(n1210) );
NAND3_X1 U1033 ( .A1(n1365), .A2(n1366), .A3(KEYINPUT52), .ZN(n1369) );
XOR2_X1 U1034 ( .A(n1371), .B(n1217), .Z(n1365) );
INV_X1 U1035 ( .A(n1211), .ZN(n1213) );
XOR2_X1 U1036 ( .A(n1372), .B(n1373), .Z(n1211) );
NOR2_X1 U1037 ( .A1(KEYINPUT47), .A2(n1321), .ZN(n1373) );
XOR2_X1 U1038 ( .A(n1317), .B(G113), .Z(n1372) );
NAND3_X1 U1039 ( .A1(n1274), .A2(n1275), .A3(n1105), .ZN(n1284) );
NOR2_X1 U1040 ( .A1(n1280), .A2(n1279), .ZN(n1105) );
INV_X1 U1041 ( .A(n1290), .ZN(n1279) );
XOR2_X1 U1042 ( .A(n1374), .B(G475), .Z(n1290) );
OR2_X1 U1043 ( .A1(n1194), .A2(G902), .ZN(n1374) );
XNOR2_X1 U1044 ( .A(n1375), .B(n1376), .ZN(n1194) );
XOR2_X1 U1045 ( .A(n1377), .B(n1378), .Z(n1376) );
XOR2_X1 U1046 ( .A(n1216), .B(n1163), .Z(n1378) );
XOR2_X1 U1047 ( .A(n1294), .B(n1243), .Z(n1163) );
INV_X1 U1048 ( .A(G140), .ZN(n1294) );
INV_X1 U1049 ( .A(n1379), .ZN(n1216) );
XOR2_X1 U1050 ( .A(n1380), .B(n1381), .Z(n1377) );
AND2_X1 U1051 ( .A1(n1359), .A2(G214), .ZN(n1381) );
NOR2_X1 U1052 ( .A1(G953), .A2(G237), .ZN(n1359) );
NAND2_X1 U1053 ( .A1(KEYINPUT43), .A2(n1382), .ZN(n1380) );
XOR2_X1 U1054 ( .A(n1383), .B(n1384), .Z(n1375) );
XOR2_X1 U1055 ( .A(G122), .B(G113), .Z(n1384) );
XNOR2_X1 U1056 ( .A(G131), .B(KEYINPUT45), .ZN(n1383) );
INV_X1 U1057 ( .A(n1292), .ZN(n1280) );
XOR2_X1 U1058 ( .A(n1385), .B(G478), .Z(n1292) );
NAND2_X1 U1059 ( .A1(n1191), .A2(n1249), .ZN(n1385) );
XNOR2_X1 U1060 ( .A(n1386), .B(n1387), .ZN(n1191) );
XOR2_X1 U1061 ( .A(n1214), .B(n1388), .Z(n1387) );
XOR2_X1 U1062 ( .A(n1389), .B(n1390), .Z(n1388) );
NOR2_X1 U1063 ( .A1(KEYINPUT38), .A2(n1391), .ZN(n1390) );
XOR2_X1 U1064 ( .A(G122), .B(G116), .Z(n1391) );
NAND2_X1 U1065 ( .A1(G217), .A2(n1353), .ZN(n1389) );
AND2_X1 U1066 ( .A1(G234), .A2(n1096), .ZN(n1353) );
INV_X1 U1067 ( .A(n1392), .ZN(n1214) );
XOR2_X1 U1068 ( .A(n1091), .B(n1393), .Z(n1386) );
XOR2_X1 U1069 ( .A(KEYINPUT63), .B(G143), .Z(n1393) );
NAND2_X1 U1070 ( .A1(n1394), .A2(n1123), .ZN(n1275) );
NAND3_X1 U1071 ( .A1(n1305), .A2(n1096), .A3(G952), .ZN(n1123) );
NAND4_X1 U1072 ( .A1(n1395), .A2(G953), .A3(G902), .A4(n1305), .ZN(n1394) );
NAND2_X1 U1073 ( .A1(G237), .A2(G234), .ZN(n1305) );
XNOR2_X1 U1074 ( .A(G898), .B(KEYINPUT57), .ZN(n1395) );
AND2_X1 U1075 ( .A1(n1103), .A2(n1303), .ZN(n1274) );
NOR2_X1 U1076 ( .A1(n1130), .A2(n1129), .ZN(n1303) );
INV_X1 U1077 ( .A(n1298), .ZN(n1129) );
NAND2_X1 U1078 ( .A1(G214), .A2(n1396), .ZN(n1298) );
XNOR2_X1 U1079 ( .A(n1397), .B(n1248), .ZN(n1130) );
INV_X1 U1080 ( .A(n1139), .ZN(n1248) );
NAND2_X1 U1081 ( .A1(G210), .A2(n1396), .ZN(n1139) );
NAND2_X1 U1082 ( .A1(n1398), .A2(n1249), .ZN(n1396) );
INV_X1 U1083 ( .A(G237), .ZN(n1398) );
NAND2_X1 U1084 ( .A1(KEYINPUT48), .A2(n1142), .ZN(n1397) );
NAND2_X1 U1085 ( .A1(n1399), .A2(n1249), .ZN(n1142) );
XOR2_X1 U1086 ( .A(n1234), .B(n1400), .Z(n1399) );
XOR2_X1 U1087 ( .A(KEYINPUT62), .B(n1401), .Z(n1400) );
NOR3_X1 U1088 ( .A1(n1402), .A2(n1403), .A3(n1404), .ZN(n1401) );
NOR3_X1 U1089 ( .A1(n1366), .A2(n1405), .A3(n1245), .ZN(n1404) );
INV_X1 U1090 ( .A(n1242), .ZN(n1366) );
NOR2_X1 U1091 ( .A1(n1242), .A2(n1406), .ZN(n1403) );
XOR2_X1 U1092 ( .A(n1240), .B(n1405), .Z(n1406) );
INV_X1 U1093 ( .A(n1245), .ZN(n1240) );
INV_X1 U1094 ( .A(n1238), .ZN(n1402) );
NAND3_X1 U1095 ( .A1(n1405), .A2(n1245), .A3(n1242), .ZN(n1238) );
XOR2_X1 U1096 ( .A(G128), .B(n1379), .Z(n1242) );
XNOR2_X1 U1097 ( .A(n1287), .B(G146), .ZN(n1379) );
INV_X1 U1098 ( .A(G143), .ZN(n1287) );
NAND2_X1 U1099 ( .A1(G224), .A2(n1096), .ZN(n1245) );
INV_X1 U1100 ( .A(G953), .ZN(n1096) );
INV_X1 U1101 ( .A(n1243), .ZN(n1405) );
XNOR2_X1 U1102 ( .A(G125), .B(KEYINPUT58), .ZN(n1243) );
XOR2_X1 U1103 ( .A(n1175), .B(n1174), .Z(n1234) );
XNOR2_X1 U1104 ( .A(n1407), .B(n1408), .ZN(n1174) );
XOR2_X1 U1105 ( .A(n1409), .B(n1225), .Z(n1408) );
XOR2_X1 U1106 ( .A(G101), .B(G110), .Z(n1225) );
NOR3_X1 U1107 ( .A1(n1410), .A2(KEYINPUT12), .A3(n1411), .ZN(n1409) );
XOR2_X1 U1108 ( .A(KEYINPUT39), .B(n1412), .Z(n1410) );
NOR2_X1 U1109 ( .A1(G104), .A2(n1091), .ZN(n1412) );
INV_X1 U1110 ( .A(G107), .ZN(n1091) );
XNOR2_X1 U1111 ( .A(G122), .B(KEYINPUT6), .ZN(n1407) );
AND2_X1 U1112 ( .A1(n1413), .A2(n1414), .ZN(n1175) );
NAND2_X1 U1113 ( .A1(n1415), .A2(n1416), .ZN(n1414) );
NAND2_X1 U1114 ( .A1(n1417), .A2(n1418), .ZN(n1416) );
NAND2_X1 U1115 ( .A1(n1419), .A2(n1420), .ZN(n1417) );
XOR2_X1 U1116 ( .A(KEYINPUT33), .B(G113), .Z(n1419) );
XOR2_X1 U1117 ( .A(n1321), .B(n1421), .Z(n1415) );
INV_X1 U1118 ( .A(G116), .ZN(n1321) );
NAND2_X1 U1119 ( .A1(n1422), .A2(n1423), .ZN(n1413) );
NAND2_X1 U1120 ( .A1(n1424), .A2(n1420), .ZN(n1423) );
INV_X1 U1121 ( .A(KEYINPUT44), .ZN(n1420) );
NAND2_X1 U1122 ( .A1(n1425), .A2(n1418), .ZN(n1424) );
INV_X1 U1123 ( .A(KEYINPUT26), .ZN(n1418) );
XOR2_X1 U1124 ( .A(n1421), .B(G116), .Z(n1425) );
NAND2_X1 U1125 ( .A1(KEYINPUT31), .A2(n1317), .ZN(n1421) );
INV_X1 U1126 ( .A(G119), .ZN(n1317) );
XOR2_X1 U1127 ( .A(KEYINPUT33), .B(n1426), .Z(n1422) );
INV_X1 U1128 ( .A(G113), .ZN(n1426) );
NOR2_X1 U1129 ( .A1(n1113), .A2(n1112), .ZN(n1103) );
INV_X1 U1130 ( .A(n1331), .ZN(n1112) );
NAND2_X1 U1131 ( .A1(G221), .A2(n1354), .ZN(n1331) );
NAND2_X1 U1132 ( .A1(G234), .A2(n1249), .ZN(n1354) );
XNOR2_X1 U1133 ( .A(n1427), .B(n1428), .ZN(n1113) );
XOR2_X1 U1134 ( .A(KEYINPUT11), .B(G469), .Z(n1428) );
NAND2_X1 U1135 ( .A1(n1429), .A2(n1249), .ZN(n1427) );
INV_X1 U1136 ( .A(G902), .ZN(n1249) );
XOR2_X1 U1137 ( .A(n1430), .B(n1431), .Z(n1429) );
XNOR2_X1 U1138 ( .A(G101), .B(n1224), .ZN(n1431) );
NAND3_X1 U1139 ( .A1(n1432), .A2(n1433), .A3(n1434), .ZN(n1224) );
NAND2_X1 U1140 ( .A1(n1411), .A2(n1435), .ZN(n1434) );
NOR2_X1 U1141 ( .A1(n1382), .A2(G107), .ZN(n1411) );
INV_X1 U1142 ( .A(G104), .ZN(n1382) );
OR3_X1 U1143 ( .A1(n1435), .A2(G104), .A3(G107), .ZN(n1433) );
NAND2_X1 U1144 ( .A1(n1436), .A2(G107), .ZN(n1432) );
XOR2_X1 U1145 ( .A(n1435), .B(G104), .Z(n1436) );
XOR2_X1 U1146 ( .A(n1164), .B(n1217), .Z(n1435) );
XOR2_X1 U1147 ( .A(n1165), .B(KEYINPUT14), .Z(n1217) );
XOR2_X1 U1148 ( .A(G131), .B(G137), .Z(n1165) );
XOR2_X1 U1149 ( .A(n1437), .B(n1438), .Z(n1164) );
XOR2_X1 U1150 ( .A(KEYINPUT13), .B(G143), .Z(n1438) );
XOR2_X1 U1151 ( .A(n1439), .B(n1392), .Z(n1437) );
XOR2_X1 U1152 ( .A(G128), .B(n1440), .Z(n1392) );
INV_X1 U1153 ( .A(n1371), .ZN(n1440) );
XNOR2_X1 U1154 ( .A(G134), .B(KEYINPUT50), .ZN(n1371) );
NAND2_X1 U1155 ( .A1(KEYINPUT29), .A2(n1285), .ZN(n1439) );
INV_X1 U1156 ( .A(G146), .ZN(n1285) );
NAND2_X1 U1157 ( .A1(n1441), .A2(KEYINPUT51), .ZN(n1430) );
XOR2_X1 U1158 ( .A(n1442), .B(n1443), .Z(n1441) );
NOR2_X1 U1159 ( .A1(KEYINPUT18), .A2(G140), .ZN(n1443) );
XOR2_X1 U1160 ( .A(n1347), .B(n1226), .Z(n1442) );
NOR2_X1 U1161 ( .A1(n1150), .A2(G953), .ZN(n1226) );
INV_X1 U1162 ( .A(G227), .ZN(n1150) );
INV_X1 U1163 ( .A(G110), .ZN(n1347) );
endmodule


