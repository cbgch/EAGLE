//Key = 0011101000100000100010000101101011010000010101001100001010011101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370;

XNOR2_X1 U752 ( .A(G107), .B(n1045), .ZN(G9) );
NOR2_X1 U753 ( .A1(n1046), .A2(n1047), .ZN(G75) );
NOR4_X1 U754 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
NOR2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
INV_X1 U756 ( .A(n1054), .ZN(n1053) );
NOR2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1052) );
NOR2_X1 U758 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
AND4_X1 U760 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(KEYINPUT49), .ZN(n1055) );
OR2_X1 U761 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U762 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
INV_X1 U763 ( .A(n1068), .ZN(n1067) );
NOR2_X1 U764 ( .A1(n1069), .A2(n1070), .ZN(n1066) );
NOR2_X1 U765 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR2_X1 U766 ( .A1(n1073), .A2(n1074), .ZN(n1064) );
INV_X1 U767 ( .A(n1075), .ZN(n1074) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1073) );
AND3_X1 U769 ( .A1(n1078), .A2(n1079), .A3(n1063), .ZN(n1050) );
NAND3_X1 U770 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1048) );
NAND4_X1 U771 ( .A1(n1083), .A2(n1078), .A3(n1063), .A4(n1084), .ZN(n1082) );
XNOR2_X1 U772 ( .A(KEYINPUT51), .B(n1085), .ZN(n1084) );
INV_X1 U773 ( .A(n1058), .ZN(n1078) );
NAND4_X1 U774 ( .A1(KEYINPUT49), .A2(n1068), .A3(n1075), .A4(n1061), .ZN(n1058) );
XNOR2_X1 U775 ( .A(n1086), .B(KEYINPUT31), .ZN(n1083) );
NOR3_X1 U776 ( .A1(n1087), .A2(G953), .A3(G952), .ZN(n1046) );
INV_X1 U777 ( .A(n1080), .ZN(n1087) );
NAND4_X1 U778 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1080) );
NOR4_X1 U779 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1071), .ZN(n1091) );
XNOR2_X1 U780 ( .A(n1095), .B(n1096), .ZN(n1092) );
INV_X1 U781 ( .A(n1086), .ZN(n1096) );
XNOR2_X1 U782 ( .A(KEYINPUT7), .B(KEYINPUT30), .ZN(n1095) );
NOR3_X1 U783 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1090) );
NAND2_X1 U784 ( .A1(n1100), .A2(n1101), .ZN(n1089) );
XOR2_X1 U785 ( .A(KEYINPUT14), .B(n1102), .Z(n1100) );
XOR2_X1 U786 ( .A(n1103), .B(n1104), .Z(n1088) );
NOR2_X1 U787 ( .A1(G475), .A2(KEYINPUT19), .ZN(n1104) );
XOR2_X1 U788 ( .A(n1105), .B(n1106), .Z(G72) );
XOR2_X1 U789 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U790 ( .A1(n1081), .A2(n1109), .ZN(n1108) );
XOR2_X1 U791 ( .A(KEYINPUT34), .B(n1110), .Z(n1109) );
NOR2_X1 U792 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U793 ( .A1(n1113), .A2(n1114), .ZN(n1107) );
NAND2_X1 U794 ( .A1(G953), .A2(n1112), .ZN(n1114) );
XOR2_X1 U795 ( .A(n1115), .B(n1116), .Z(n1113) );
XNOR2_X1 U796 ( .A(n1117), .B(n1118), .ZN(n1116) );
NAND2_X1 U797 ( .A1(KEYINPUT63), .A2(n1119), .ZN(n1117) );
XOR2_X1 U798 ( .A(n1120), .B(n1121), .Z(n1115) );
NOR2_X1 U799 ( .A1(KEYINPUT1), .A2(n1122), .ZN(n1121) );
XNOR2_X1 U800 ( .A(G125), .B(n1123), .ZN(n1120) );
NOR2_X1 U801 ( .A1(KEYINPUT29), .A2(n1124), .ZN(n1123) );
INV_X1 U802 ( .A(G140), .ZN(n1124) );
NAND2_X1 U803 ( .A1(n1081), .A2(n1125), .ZN(n1105) );
NAND2_X1 U804 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XNOR2_X1 U805 ( .A(KEYINPUT3), .B(n1128), .ZN(n1127) );
NAND3_X1 U806 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(G69) );
XOR2_X1 U807 ( .A(n1132), .B(KEYINPUT17), .Z(n1131) );
NAND3_X1 U808 ( .A1(n1133), .A2(n1134), .A3(G953), .ZN(n1132) );
NAND2_X1 U809 ( .A1(G898), .A2(G224), .ZN(n1133) );
NAND2_X1 U810 ( .A1(n1135), .A2(n1081), .ZN(n1130) );
XNOR2_X1 U811 ( .A(n1136), .B(n1134), .ZN(n1135) );
NAND2_X1 U812 ( .A1(n1137), .A2(n1045), .ZN(n1136) );
NAND3_X1 U813 ( .A1(n1138), .A2(G224), .A3(G953), .ZN(n1129) );
INV_X1 U814 ( .A(n1134), .ZN(n1138) );
NAND2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(n1134) );
NAND2_X1 U816 ( .A1(G953), .A2(n1141), .ZN(n1140) );
XOR2_X1 U817 ( .A(n1142), .B(n1143), .Z(n1139) );
NOR2_X1 U818 ( .A1(KEYINPUT50), .A2(n1144), .ZN(n1143) );
XOR2_X1 U819 ( .A(KEYINPUT56), .B(n1145), .Z(n1144) );
XOR2_X1 U820 ( .A(n1146), .B(KEYINPUT62), .Z(n1142) );
NOR2_X1 U821 ( .A1(n1147), .A2(n1148), .ZN(G66) );
XOR2_X1 U822 ( .A(n1149), .B(n1150), .Z(n1148) );
NAND3_X1 U823 ( .A1(n1151), .A2(n1152), .A3(KEYINPUT48), .ZN(n1149) );
XOR2_X1 U824 ( .A(KEYINPUT9), .B(G217), .Z(n1152) );
NOR2_X1 U825 ( .A1(n1147), .A2(n1153), .ZN(G63) );
XOR2_X1 U826 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U827 ( .A1(n1156), .A2(KEYINPUT5), .ZN(n1154) );
AND2_X1 U828 ( .A1(G478), .A2(n1151), .ZN(n1156) );
NOR2_X1 U829 ( .A1(n1147), .A2(n1157), .ZN(G60) );
NOR3_X1 U830 ( .A1(n1103), .A2(n1158), .A3(n1159), .ZN(n1157) );
NOR2_X1 U831 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
AND2_X1 U832 ( .A1(n1049), .A2(G475), .ZN(n1160) );
AND3_X1 U833 ( .A1(n1161), .A2(G475), .A3(n1151), .ZN(n1158) );
XNOR2_X1 U834 ( .A(G104), .B(n1162), .ZN(G6) );
NOR2_X1 U835 ( .A1(n1147), .A2(n1163), .ZN(G57) );
XOR2_X1 U836 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U837 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U838 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U839 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
INV_X1 U840 ( .A(KEYINPUT54), .ZN(n1171) );
NOR3_X1 U841 ( .A1(KEYINPUT54), .A2(n1172), .A3(n1173), .ZN(n1168) );
NOR2_X1 U842 ( .A1(KEYINPUT46), .A2(n1174), .ZN(n1166) );
XOR2_X1 U843 ( .A(n1175), .B(n1176), .Z(n1164) );
AND2_X1 U844 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
AND2_X1 U845 ( .A1(G472), .A2(n1151), .ZN(n1175) );
NOR2_X1 U846 ( .A1(n1147), .A2(n1179), .ZN(G54) );
XOR2_X1 U847 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U848 ( .A(n1182), .B(n1183), .Z(n1181) );
AND2_X1 U849 ( .A1(G469), .A2(n1151), .ZN(n1183) );
INV_X1 U850 ( .A(n1184), .ZN(n1151) );
NAND3_X1 U851 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1182) );
NAND2_X1 U852 ( .A1(KEYINPUT12), .A2(n1188), .ZN(n1187) );
OR3_X1 U853 ( .A1(n1188), .A2(KEYINPUT12), .A3(n1122), .ZN(n1186) );
NAND2_X1 U854 ( .A1(n1122), .A2(n1189), .ZN(n1185) );
NAND2_X1 U855 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
INV_X1 U856 ( .A(KEYINPUT12), .ZN(n1191) );
XNOR2_X1 U857 ( .A(n1192), .B(KEYINPUT32), .ZN(n1190) );
NOR2_X1 U858 ( .A1(n1193), .A2(n1194), .ZN(G51) );
XOR2_X1 U859 ( .A(KEYINPUT38), .B(n1147), .Z(n1194) );
NOR2_X1 U860 ( .A1(n1081), .A2(G952), .ZN(n1147) );
XOR2_X1 U861 ( .A(n1195), .B(n1196), .Z(n1193) );
NOR2_X1 U862 ( .A1(n1197), .A2(n1184), .ZN(n1196) );
NAND2_X1 U863 ( .A1(G902), .A2(n1049), .ZN(n1184) );
NAND4_X1 U864 ( .A1(n1198), .A2(n1137), .A3(n1126), .A4(n1128), .ZN(n1049) );
OR2_X1 U865 ( .A1(n1199), .A2(n1200), .ZN(n1128) );
AND4_X1 U866 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1126) );
AND4_X1 U867 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
NAND2_X1 U868 ( .A1(n1209), .A2(n1077), .ZN(n1203) );
AND4_X1 U869 ( .A1(n1162), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1137) );
AND4_X1 U870 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1212) );
NAND2_X1 U871 ( .A1(n1217), .A2(n1218), .ZN(n1211) );
NAND3_X1 U872 ( .A1(n1219), .A2(n1068), .A3(n1060), .ZN(n1162) );
XOR2_X1 U873 ( .A(n1045), .B(KEYINPUT11), .Z(n1198) );
NAND3_X1 U874 ( .A1(n1059), .A2(n1068), .A3(n1219), .ZN(n1045) );
NOR2_X1 U875 ( .A1(n1220), .A2(n1221), .ZN(n1195) );
XOR2_X1 U876 ( .A(n1222), .B(KEYINPUT35), .Z(n1221) );
NAND2_X1 U877 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
NOR2_X1 U878 ( .A1(n1223), .A2(n1224), .ZN(n1220) );
XOR2_X1 U879 ( .A(n1225), .B(n1226), .Z(n1224) );
XNOR2_X1 U880 ( .A(G146), .B(n1201), .ZN(G48) );
NAND3_X1 U881 ( .A1(n1060), .A2(n1070), .A3(n1227), .ZN(n1201) );
XNOR2_X1 U882 ( .A(n1228), .B(n1229), .ZN(G45) );
NOR2_X1 U883 ( .A1(n1199), .A2(n1230), .ZN(n1229) );
XNOR2_X1 U884 ( .A(KEYINPUT10), .B(n1200), .ZN(n1230) );
INV_X1 U885 ( .A(n1077), .ZN(n1200) );
NAND4_X1 U886 ( .A1(n1231), .A2(n1070), .A3(n1232), .A4(n1094), .ZN(n1199) );
XNOR2_X1 U887 ( .A(G140), .B(n1202), .ZN(G42) );
NAND2_X1 U888 ( .A1(n1209), .A2(n1076), .ZN(n1202) );
XNOR2_X1 U889 ( .A(G137), .B(n1206), .ZN(G39) );
NAND3_X1 U890 ( .A1(n1063), .A2(n1075), .A3(n1227), .ZN(n1206) );
NAND2_X1 U891 ( .A1(n1233), .A2(n1234), .ZN(G36) );
OR2_X1 U892 ( .A1(n1208), .A2(G134), .ZN(n1234) );
XOR2_X1 U893 ( .A(n1235), .B(KEYINPUT23), .Z(n1233) );
NAND2_X1 U894 ( .A1(G134), .A2(n1208), .ZN(n1235) );
NAND4_X1 U895 ( .A1(n1231), .A2(n1077), .A3(n1059), .A4(n1075), .ZN(n1208) );
XNOR2_X1 U896 ( .A(G131), .B(n1236), .ZN(G33) );
NAND2_X1 U897 ( .A1(n1237), .A2(n1209), .ZN(n1236) );
AND3_X1 U898 ( .A1(n1060), .A2(n1075), .A3(n1231), .ZN(n1209) );
NAND2_X1 U899 ( .A1(n1238), .A2(n1239), .ZN(n1075) );
NAND2_X1 U900 ( .A1(n1070), .A2(n1240), .ZN(n1239) );
INV_X1 U901 ( .A(KEYINPUT25), .ZN(n1240) );
NAND3_X1 U902 ( .A1(n1241), .A2(n1072), .A3(KEYINPUT25), .ZN(n1238) );
XNOR2_X1 U903 ( .A(n1077), .B(KEYINPUT6), .ZN(n1237) );
XNOR2_X1 U904 ( .A(G128), .B(n1205), .ZN(G30) );
NAND3_X1 U905 ( .A1(n1059), .A2(n1070), .A3(n1227), .ZN(n1205) );
AND3_X1 U906 ( .A1(n1093), .A2(n1242), .A3(n1231), .ZN(n1227) );
NOR2_X1 U907 ( .A1(n1243), .A2(n1244), .ZN(n1231) );
XNOR2_X1 U908 ( .A(G101), .B(n1210), .ZN(G3) );
NAND3_X1 U909 ( .A1(n1063), .A2(n1219), .A3(n1077), .ZN(n1210) );
XNOR2_X1 U910 ( .A(G125), .B(n1207), .ZN(G27) );
NAND4_X1 U911 ( .A1(n1076), .A2(n1070), .A3(n1054), .A4(n1245), .ZN(n1207) );
NOR2_X1 U912 ( .A1(n1246), .A2(n1243), .ZN(n1245) );
NAND2_X1 U913 ( .A1(n1247), .A2(n1061), .ZN(n1243) );
NAND2_X1 U914 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND3_X1 U915 ( .A1(G953), .A2(n1112), .A3(G902), .ZN(n1249) );
INV_X1 U916 ( .A(G900), .ZN(n1112) );
XNOR2_X1 U917 ( .A(G122), .B(n1216), .ZN(G24) );
NAND4_X1 U918 ( .A1(n1218), .A2(n1068), .A3(n1232), .A4(n1094), .ZN(n1216) );
NOR2_X1 U919 ( .A1(n1242), .A2(n1093), .ZN(n1068) );
XOR2_X1 U920 ( .A(n1250), .B(n1251), .Z(G21) );
NAND2_X1 U921 ( .A1(KEYINPUT45), .A2(n1252), .ZN(n1251) );
XOR2_X1 U922 ( .A(KEYINPUT0), .B(G119), .Z(n1252) );
NAND4_X1 U923 ( .A1(n1217), .A2(n1054), .A3(n1253), .A4(n1254), .ZN(n1250) );
XOR2_X1 U924 ( .A(KEYINPUT22), .B(n1070), .Z(n1254) );
AND3_X1 U925 ( .A1(n1093), .A2(n1242), .A3(n1063), .ZN(n1217) );
INV_X1 U926 ( .A(n1255), .ZN(n1242) );
XNOR2_X1 U927 ( .A(G116), .B(n1215), .ZN(G18) );
NAND3_X1 U928 ( .A1(n1218), .A2(n1059), .A3(n1077), .ZN(n1215) );
NOR2_X1 U929 ( .A1(n1232), .A2(n1256), .ZN(n1059) );
XNOR2_X1 U930 ( .A(G113), .B(n1214), .ZN(G15) );
NAND3_X1 U931 ( .A1(n1060), .A2(n1218), .A3(n1077), .ZN(n1214) );
NOR2_X1 U932 ( .A1(n1093), .A2(n1255), .ZN(n1077) );
AND3_X1 U933 ( .A1(n1253), .A2(n1070), .A3(n1054), .ZN(n1218) );
NOR2_X1 U934 ( .A1(n1086), .A2(n1099), .ZN(n1054) );
INV_X1 U935 ( .A(n1246), .ZN(n1060) );
NAND2_X1 U936 ( .A1(n1256), .A2(n1232), .ZN(n1246) );
INV_X1 U937 ( .A(n1094), .ZN(n1256) );
XNOR2_X1 U938 ( .A(G110), .B(n1213), .ZN(G12) );
NAND3_X1 U939 ( .A1(n1076), .A2(n1219), .A3(n1063), .ZN(n1213) );
NOR2_X1 U940 ( .A1(n1094), .A2(n1232), .ZN(n1063) );
XOR2_X1 U941 ( .A(n1103), .B(G475), .Z(n1232) );
NOR2_X1 U942 ( .A1(n1161), .A2(G902), .ZN(n1103) );
XOR2_X1 U943 ( .A(n1257), .B(n1258), .Z(n1161) );
XOR2_X1 U944 ( .A(n1259), .B(n1260), .Z(n1258) );
NOR2_X1 U945 ( .A1(G104), .A2(KEYINPUT8), .ZN(n1260) );
NOR2_X1 U946 ( .A1(n1261), .A2(n1262), .ZN(n1259) );
XOR2_X1 U947 ( .A(KEYINPUT15), .B(n1263), .Z(n1262) );
NOR2_X1 U948 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
AND2_X1 U949 ( .A1(n1264), .A2(n1265), .ZN(n1261) );
XOR2_X1 U950 ( .A(G113), .B(KEYINPUT36), .Z(n1265) );
INV_X1 U951 ( .A(G122), .ZN(n1264) );
NAND2_X1 U952 ( .A1(n1266), .A2(n1267), .ZN(n1257) );
NAND2_X1 U953 ( .A1(n1268), .A2(n1119), .ZN(n1267) );
INV_X1 U954 ( .A(G131), .ZN(n1119) );
XNOR2_X1 U955 ( .A(n1269), .B(KEYINPUT52), .ZN(n1268) );
NAND2_X1 U956 ( .A1(n1270), .A2(G131), .ZN(n1266) );
XNOR2_X1 U957 ( .A(KEYINPUT57), .B(n1271), .ZN(n1270) );
INV_X1 U958 ( .A(n1269), .ZN(n1271) );
XNOR2_X1 U959 ( .A(n1272), .B(n1273), .ZN(n1269) );
NOR2_X1 U960 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XOR2_X1 U961 ( .A(KEYINPUT18), .B(n1276), .Z(n1275) );
NOR2_X1 U962 ( .A1(G146), .A2(n1277), .ZN(n1276) );
AND2_X1 U963 ( .A1(n1277), .A2(G146), .ZN(n1274) );
XNOR2_X1 U964 ( .A(n1278), .B(n1228), .ZN(n1272) );
NAND2_X1 U965 ( .A1(n1279), .A2(G214), .ZN(n1278) );
XNOR2_X1 U966 ( .A(n1280), .B(G478), .ZN(n1094) );
NAND2_X1 U967 ( .A1(n1155), .A2(n1281), .ZN(n1280) );
XNOR2_X1 U968 ( .A(n1282), .B(n1283), .ZN(n1155) );
XOR2_X1 U969 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U970 ( .A(n1286), .B(G122), .ZN(n1285) );
XNOR2_X1 U971 ( .A(n1228), .B(G134), .ZN(n1284) );
INV_X1 U972 ( .A(G143), .ZN(n1228) );
XOR2_X1 U973 ( .A(n1287), .B(n1288), .Z(n1282) );
XOR2_X1 U974 ( .A(G116), .B(G107), .Z(n1288) );
NAND2_X1 U975 ( .A1(G217), .A2(n1289), .ZN(n1287) );
AND3_X1 U976 ( .A1(n1253), .A2(n1070), .A3(n1079), .ZN(n1219) );
INV_X1 U977 ( .A(n1244), .ZN(n1079) );
NAND2_X1 U978 ( .A1(n1290), .A2(n1086), .ZN(n1244) );
XNOR2_X1 U979 ( .A(n1291), .B(G469), .ZN(n1086) );
NAND2_X1 U980 ( .A1(n1292), .A2(n1281), .ZN(n1291) );
XOR2_X1 U981 ( .A(n1293), .B(n1294), .Z(n1292) );
XNOR2_X1 U982 ( .A(n1180), .B(n1188), .ZN(n1294) );
INV_X1 U983 ( .A(n1192), .ZN(n1188) );
XOR2_X1 U984 ( .A(n1295), .B(n1296), .Z(n1192) );
XOR2_X1 U985 ( .A(n1297), .B(n1298), .Z(n1180) );
XNOR2_X1 U986 ( .A(n1299), .B(n1300), .ZN(n1298) );
XNOR2_X1 U987 ( .A(G140), .B(n1301), .ZN(n1297) );
NOR2_X1 U988 ( .A1(G953), .A2(n1111), .ZN(n1301) );
INV_X1 U989 ( .A(G227), .ZN(n1111) );
XNOR2_X1 U990 ( .A(n1122), .B(KEYINPUT26), .ZN(n1293) );
XNOR2_X1 U991 ( .A(n1099), .B(KEYINPUT39), .ZN(n1290) );
INV_X1 U992 ( .A(n1085), .ZN(n1099) );
NAND2_X1 U993 ( .A1(G221), .A2(n1302), .ZN(n1085) );
NAND2_X1 U994 ( .A1(G234), .A2(n1281), .ZN(n1302) );
NOR2_X1 U995 ( .A1(n1241), .A2(n1097), .ZN(n1070) );
INV_X1 U996 ( .A(n1072), .ZN(n1097) );
NAND2_X1 U997 ( .A1(G214), .A2(n1303), .ZN(n1072) );
INV_X1 U998 ( .A(n1071), .ZN(n1241) );
XOR2_X1 U999 ( .A(n1304), .B(n1197), .Z(n1071) );
NAND2_X1 U1000 ( .A1(G210), .A2(n1303), .ZN(n1197) );
NAND2_X1 U1001 ( .A1(n1305), .A2(n1306), .ZN(n1303) );
INV_X1 U1002 ( .A(G237), .ZN(n1306) );
XNOR2_X1 U1003 ( .A(G902), .B(KEYINPUT44), .ZN(n1305) );
NAND2_X1 U1004 ( .A1(n1307), .A2(n1281), .ZN(n1304) );
XOR2_X1 U1005 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U1006 ( .A(n1225), .B(n1223), .Z(n1309) );
XOR2_X1 U1007 ( .A(n1146), .B(n1145), .Z(n1223) );
XNOR2_X1 U1008 ( .A(n1310), .B(n1311), .ZN(n1145) );
XNOR2_X1 U1009 ( .A(n1312), .B(n1296), .ZN(n1311) );
XNOR2_X1 U1010 ( .A(n1313), .B(KEYINPUT33), .ZN(n1296) );
XNOR2_X1 U1011 ( .A(n1314), .B(n1315), .ZN(n1310) );
INV_X1 U1012 ( .A(G113), .ZN(n1315) );
NAND2_X1 U1013 ( .A1(KEYINPUT27), .A2(n1295), .ZN(n1314) );
XOR2_X1 U1014 ( .A(G104), .B(G107), .Z(n1295) );
NAND2_X1 U1015 ( .A1(n1316), .A2(n1317), .ZN(n1146) );
NAND2_X1 U1016 ( .A1(G122), .A2(n1299), .ZN(n1317) );
XOR2_X1 U1017 ( .A(KEYINPUT43), .B(n1318), .Z(n1316) );
NOR2_X1 U1018 ( .A1(n1299), .A2(n1319), .ZN(n1318) );
XNOR2_X1 U1019 ( .A(G122), .B(KEYINPUT2), .ZN(n1319) );
NAND2_X1 U1020 ( .A1(G224), .A2(n1081), .ZN(n1225) );
XNOR2_X1 U1021 ( .A(KEYINPUT16), .B(n1320), .ZN(n1308) );
NOR3_X1 U1022 ( .A1(KEYINPUT37), .A2(n1321), .A3(n1322), .ZN(n1320) );
NOR3_X1 U1023 ( .A1(KEYINPUT41), .A2(n1172), .A3(n1323), .ZN(n1322) );
AND2_X1 U1024 ( .A1(n1226), .A2(KEYINPUT41), .ZN(n1321) );
XOR2_X1 U1025 ( .A(n1172), .B(n1323), .Z(n1226) );
INV_X1 U1026 ( .A(G125), .ZN(n1323) );
AND2_X1 U1027 ( .A1(n1061), .A2(n1324), .ZN(n1253) );
NAND2_X1 U1028 ( .A1(n1325), .A2(n1248), .ZN(n1324) );
NAND2_X1 U1029 ( .A1(G952), .A2(n1326), .ZN(n1248) );
XNOR2_X1 U1030 ( .A(KEYINPUT59), .B(n1081), .ZN(n1326) );
INV_X1 U1031 ( .A(G953), .ZN(n1081) );
NAND3_X1 U1032 ( .A1(G953), .A2(n1141), .A3(G902), .ZN(n1325) );
INV_X1 U1033 ( .A(G898), .ZN(n1141) );
NAND2_X1 U1034 ( .A1(G237), .A2(G234), .ZN(n1061) );
AND2_X1 U1035 ( .A1(n1255), .A2(n1093), .ZN(n1076) );
NAND3_X1 U1036 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1093) );
NAND2_X1 U1037 ( .A1(G217), .A2(G902), .ZN(n1329) );
NAND3_X1 U1038 ( .A1(n1150), .A2(n1281), .A3(n1330), .ZN(n1328) );
OR2_X1 U1039 ( .A1(n1330), .A2(n1150), .ZN(n1327) );
XNOR2_X1 U1040 ( .A(n1331), .B(n1332), .ZN(n1150) );
XNOR2_X1 U1041 ( .A(n1333), .B(n1277), .ZN(n1332) );
XOR2_X1 U1042 ( .A(G125), .B(G140), .Z(n1277) );
NAND2_X1 U1043 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NAND2_X1 U1044 ( .A1(G137), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1045 ( .A(n1337), .B(n1338), .Z(n1334) );
NOR2_X1 U1046 ( .A1(G137), .A2(n1336), .ZN(n1338) );
INV_X1 U1047 ( .A(KEYINPUT60), .ZN(n1336) );
NAND2_X1 U1048 ( .A1(n1289), .A2(G221), .ZN(n1337) );
NOR2_X1 U1049 ( .A1(n1339), .A2(G953), .ZN(n1289) );
XNOR2_X1 U1050 ( .A(n1340), .B(n1341), .ZN(n1331) );
NAND2_X1 U1051 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
NAND2_X1 U1052 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
XNOR2_X1 U1053 ( .A(KEYINPUT40), .B(n1299), .ZN(n1345) );
XNOR2_X1 U1054 ( .A(n1286), .B(G119), .ZN(n1344) );
INV_X1 U1055 ( .A(G128), .ZN(n1286) );
NAND2_X1 U1056 ( .A1(n1346), .A2(n1347), .ZN(n1342) );
XNOR2_X1 U1057 ( .A(KEYINPUT61), .B(n1299), .ZN(n1347) );
XNOR2_X1 U1058 ( .A(G110), .B(KEYINPUT55), .ZN(n1299) );
XNOR2_X1 U1059 ( .A(G119), .B(G128), .ZN(n1346) );
NAND2_X1 U1060 ( .A1(G217), .A2(n1339), .ZN(n1330) );
INV_X1 U1061 ( .A(G234), .ZN(n1339) );
NOR2_X1 U1062 ( .A1(n1348), .A2(n1098), .ZN(n1255) );
NOR2_X1 U1063 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
AND2_X1 U1064 ( .A1(n1349), .A2(n1101), .ZN(n1348) );
NAND3_X1 U1065 ( .A1(n1350), .A2(n1351), .A3(n1281), .ZN(n1101) );
INV_X1 U1066 ( .A(G902), .ZN(n1281) );
NAND2_X1 U1067 ( .A1(KEYINPUT28), .A2(n1352), .ZN(n1351) );
XOR2_X1 U1068 ( .A(n1353), .B(n1354), .Z(n1352) );
NOR2_X1 U1069 ( .A1(KEYINPUT58), .A2(n1355), .ZN(n1354) );
OR3_X1 U1070 ( .A1(n1353), .A2(n1356), .A3(KEYINPUT28), .ZN(n1350) );
INV_X1 U1071 ( .A(n1355), .ZN(n1356) );
NAND2_X1 U1072 ( .A1(n1357), .A2(n1178), .ZN(n1355) );
NAND2_X1 U1073 ( .A1(n1313), .A2(n1358), .ZN(n1178) );
NAND2_X1 U1074 ( .A1(n1279), .A2(G210), .ZN(n1358) );
INV_X1 U1075 ( .A(G101), .ZN(n1313) );
XOR2_X1 U1076 ( .A(n1177), .B(KEYINPUT21), .Z(n1357) );
NAND3_X1 U1077 ( .A1(G210), .A2(G101), .A3(n1279), .ZN(n1177) );
NOR2_X1 U1078 ( .A1(G953), .A2(G237), .ZN(n1279) );
NAND2_X1 U1079 ( .A1(n1359), .A2(n1360), .ZN(n1353) );
OR2_X1 U1080 ( .A1(n1174), .A2(n1170), .ZN(n1360) );
XOR2_X1 U1081 ( .A(n1361), .B(KEYINPUT42), .Z(n1359) );
NAND2_X1 U1082 ( .A1(n1170), .A2(n1174), .ZN(n1361) );
XNOR2_X1 U1083 ( .A(G113), .B(n1362), .ZN(n1174) );
NOR2_X1 U1084 ( .A1(KEYINPUT47), .A2(n1312), .ZN(n1362) );
XNOR2_X1 U1085 ( .A(G116), .B(G119), .ZN(n1312) );
XNOR2_X1 U1086 ( .A(n1172), .B(n1173), .ZN(n1170) );
INV_X1 U1087 ( .A(n1300), .ZN(n1173) );
XOR2_X1 U1088 ( .A(G131), .B(n1363), .Z(n1300) );
NOR2_X1 U1089 ( .A1(n1364), .A2(n1365), .ZN(n1363) );
NOR2_X1 U1090 ( .A1(KEYINPUT4), .A2(n1118), .ZN(n1365) );
INV_X1 U1091 ( .A(n1366), .ZN(n1118) );
NOR2_X1 U1092 ( .A1(KEYINPUT13), .A2(n1366), .ZN(n1364) );
XNOR2_X1 U1093 ( .A(G134), .B(G137), .ZN(n1366) );
NAND2_X1 U1094 ( .A1(n1367), .A2(n1368), .ZN(n1172) );
NAND2_X1 U1095 ( .A1(n1122), .A2(n1369), .ZN(n1368) );
XOR2_X1 U1096 ( .A(G128), .B(n1370), .Z(n1122) );
OR3_X1 U1097 ( .A1(n1370), .A2(G128), .A3(n1369), .ZN(n1367) );
INV_X1 U1098 ( .A(KEYINPUT53), .ZN(n1369) );
XNOR2_X1 U1099 ( .A(G143), .B(n1341), .ZN(n1370) );
INV_X1 U1100 ( .A(G146), .ZN(n1341) );
XNOR2_X1 U1101 ( .A(n1102), .B(KEYINPUT20), .ZN(n1349) );
XOR2_X1 U1102 ( .A(G472), .B(KEYINPUT24), .Z(n1102) );
endmodule


