//Key = 0010111000011101010011110100100010011101111111000000000111011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322;

XNOR2_X1 U729 ( .A(G107), .B(n1007), .ZN(G9) );
NOR2_X1 U730 ( .A1(n1008), .A2(n1009), .ZN(G75) );
NOR4_X1 U731 ( .A1(n1010), .A2(n1011), .A3(G953), .A4(n1012), .ZN(n1009) );
NOR3_X1 U732 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1011) );
NOR2_X1 U733 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
AND2_X1 U734 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NAND3_X1 U735 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1010) );
NAND3_X1 U736 ( .A1(n1023), .A2(n1024), .A3(n1018), .ZN(n1021) );
NAND3_X1 U737 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1023) );
NAND2_X1 U738 ( .A1(KEYINPUT24), .A2(n1028), .ZN(n1027) );
NAND4_X1 U739 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1028) );
NAND3_X1 U740 ( .A1(n1030), .A2(n1033), .A3(n1029), .ZN(n1026) );
NAND2_X1 U741 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U742 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
XOR2_X1 U743 ( .A(n1038), .B(n1039), .Z(n1036) );
NOR2_X1 U744 ( .A1(KEYINPUT34), .A2(n1040), .ZN(n1039) );
NAND2_X1 U745 ( .A1(n1032), .A2(n1041), .ZN(n1034) );
NAND2_X1 U746 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
OR2_X1 U747 ( .A1(n1044), .A2(KEYINPUT24), .ZN(n1043) );
NAND2_X1 U748 ( .A1(n1045), .A2(n1046), .ZN(n1025) );
OR2_X1 U749 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
INV_X1 U750 ( .A(n1013), .ZN(n1045) );
NAND3_X1 U751 ( .A1(n1032), .A2(n1037), .A3(n1029), .ZN(n1013) );
INV_X1 U752 ( .A(n1049), .ZN(n1029) );
NOR3_X1 U753 ( .A1(n1012), .A2(G953), .A3(G952), .ZN(n1008) );
AND4_X1 U754 ( .A1(n1050), .A2(n1037), .A3(n1051), .A4(n1052), .ZN(n1012) );
NOR4_X1 U755 ( .A1(n1053), .A2(n1019), .A3(n1054), .A4(n1055), .ZN(n1052) );
XOR2_X1 U756 ( .A(n1056), .B(KEYINPUT13), .Z(n1055) );
XOR2_X1 U757 ( .A(n1018), .B(KEYINPUT43), .Z(n1054) );
XOR2_X1 U758 ( .A(n1057), .B(n1058), .Z(n1051) );
XOR2_X1 U759 ( .A(KEYINPUT3), .B(G475), .Z(n1058) );
NAND2_X1 U760 ( .A1(n1059), .A2(n1060), .ZN(G72) );
NAND2_X1 U761 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U762 ( .A1(G953), .A2(n1063), .ZN(n1062) );
NAND2_X1 U763 ( .A1(G900), .A2(G227), .ZN(n1063) );
NAND2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(n1059) );
INV_X1 U765 ( .A(n1061), .ZN(n1065) );
NOR2_X1 U766 ( .A1(KEYINPUT9), .A2(n1066), .ZN(n1061) );
XOR2_X1 U767 ( .A(n1067), .B(n1068), .Z(n1066) );
NOR2_X1 U768 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XOR2_X1 U769 ( .A(n1071), .B(n1072), .Z(n1070) );
XNOR2_X1 U770 ( .A(n1073), .B(n1074), .ZN(n1072) );
NAND2_X1 U771 ( .A1(KEYINPUT35), .A2(n1075), .ZN(n1073) );
NAND2_X1 U772 ( .A1(n1076), .A2(n1077), .ZN(n1067) );
XOR2_X1 U773 ( .A(n1078), .B(KEYINPUT18), .Z(n1076) );
NAND2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1064) );
OR2_X1 U775 ( .A1(n1078), .A2(G227), .ZN(n1080) );
INV_X1 U776 ( .A(n1069), .ZN(n1079) );
XOR2_X1 U777 ( .A(n1081), .B(n1082), .Z(G69) );
XOR2_X1 U778 ( .A(n1083), .B(n1084), .Z(n1082) );
NOR2_X1 U779 ( .A1(n1020), .A2(G953), .ZN(n1084) );
NAND3_X1 U780 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1083) );
INV_X1 U781 ( .A(n1088), .ZN(n1087) );
NAND2_X1 U782 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NAND2_X1 U783 ( .A1(n1091), .A2(n1092), .ZN(n1085) );
XOR2_X1 U784 ( .A(n1089), .B(KEYINPUT5), .Z(n1092) );
XOR2_X1 U785 ( .A(n1093), .B(n1094), .Z(n1089) );
NAND2_X1 U786 ( .A1(G953), .A2(n1095), .ZN(n1081) );
NAND2_X1 U787 ( .A1(G898), .A2(G224), .ZN(n1095) );
NOR2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(G66) );
XNOR2_X1 U789 ( .A(n1098), .B(n1099), .ZN(n1097) );
NOR2_X1 U790 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U791 ( .A1(n1096), .A2(n1102), .ZN(G63) );
XOR2_X1 U792 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR2_X1 U793 ( .A1(n1105), .A2(n1101), .ZN(n1103) );
INV_X1 U794 ( .A(G478), .ZN(n1105) );
NOR2_X1 U795 ( .A1(n1096), .A2(n1106), .ZN(G60) );
NOR2_X1 U796 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XOR2_X1 U797 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U798 ( .A1(KEYINPUT50), .A2(n1111), .ZN(n1110) );
NOR2_X1 U799 ( .A1(n1112), .A2(n1101), .ZN(n1109) );
INV_X1 U800 ( .A(G475), .ZN(n1112) );
AND2_X1 U801 ( .A1(n1111), .A2(KEYINPUT50), .ZN(n1107) );
XOR2_X1 U802 ( .A(G104), .B(n1113), .Z(G6) );
NOR3_X1 U803 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1113) );
NOR2_X1 U804 ( .A1(n1096), .A2(n1117), .ZN(G57) );
XOR2_X1 U805 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND2_X1 U806 ( .A1(KEYINPUT6), .A2(n1120), .ZN(n1119) );
NAND3_X1 U807 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1118) );
NAND2_X1 U808 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
INV_X1 U809 ( .A(n1126), .ZN(n1125) );
NAND3_X1 U810 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1122) );
INV_X1 U811 ( .A(n1129), .ZN(n1128) );
NAND2_X1 U812 ( .A1(n1130), .A2(n1129), .ZN(n1121) );
XOR2_X1 U813 ( .A(n1127), .B(n1126), .Z(n1130) );
NOR3_X1 U814 ( .A1(KEYINPUT10), .A2(n1131), .A3(n1101), .ZN(n1126) );
INV_X1 U815 ( .A(G472), .ZN(n1131) );
NOR2_X1 U816 ( .A1(n1096), .A2(n1132), .ZN(G54) );
XOR2_X1 U817 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U818 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U819 ( .A1(n1137), .A2(n1101), .ZN(n1136) );
INV_X1 U820 ( .A(G469), .ZN(n1137) );
NOR2_X1 U821 ( .A1(n1096), .A2(n1138), .ZN(G51) );
XOR2_X1 U822 ( .A(n1139), .B(n1140), .Z(n1138) );
XNOR2_X1 U823 ( .A(n1141), .B(n1142), .ZN(n1140) );
NOR2_X1 U824 ( .A1(KEYINPUT51), .A2(n1143), .ZN(n1141) );
XNOR2_X1 U825 ( .A(n1144), .B(n1145), .ZN(n1143) );
XNOR2_X1 U826 ( .A(KEYINPUT28), .B(n1146), .ZN(n1145) );
NOR2_X1 U827 ( .A1(n1147), .A2(n1101), .ZN(n1139) );
NAND2_X1 U828 ( .A1(G902), .A2(n1148), .ZN(n1101) );
NAND2_X1 U829 ( .A1(n1022), .A2(n1020), .ZN(n1148) );
AND4_X1 U830 ( .A1(n1149), .A2(n1007), .A3(n1150), .A4(n1151), .ZN(n1020) );
NOR3_X1 U831 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
NOR2_X1 U832 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR3_X1 U833 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1155) );
NOR2_X1 U834 ( .A1(n1160), .A2(n1015), .ZN(n1159) );
XOR2_X1 U835 ( .A(n1161), .B(KEYINPUT8), .Z(n1160) );
AND3_X1 U836 ( .A1(n1162), .A2(n1163), .A3(n1037), .ZN(n1158) );
NOR2_X1 U837 ( .A1(n1164), .A2(n1165), .ZN(n1157) );
INV_X1 U838 ( .A(KEYINPUT41), .ZN(n1165) );
NOR4_X1 U839 ( .A1(KEYINPUT41), .A2(n1032), .A3(n1166), .A4(n1164), .ZN(n1153) );
NOR2_X1 U840 ( .A1(n1167), .A2(n1115), .ZN(n1152) );
NOR2_X1 U841 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U842 ( .A1(n1170), .A2(n1044), .ZN(n1169) );
XOR2_X1 U843 ( .A(n1015), .B(KEYINPUT7), .Z(n1170) );
INV_X1 U844 ( .A(n1030), .ZN(n1015) );
NOR2_X1 U845 ( .A1(n1171), .A2(n1114), .ZN(n1168) );
XOR2_X1 U846 ( .A(n1116), .B(KEYINPUT33), .Z(n1171) );
NAND3_X1 U847 ( .A1(n1172), .A2(n1048), .A3(n1037), .ZN(n1007) );
INV_X1 U848 ( .A(n1077), .ZN(n1022) );
NAND4_X1 U849 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1077) );
AND3_X1 U850 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1176) );
NAND2_X1 U851 ( .A1(n1180), .A2(n1181), .ZN(n1175) );
NAND4_X1 U852 ( .A1(n1182), .A2(n1164), .A3(n1183), .A4(n1184), .ZN(n1181) );
OR2_X1 U853 ( .A1(n1185), .A2(KEYINPUT30), .ZN(n1184) );
NAND3_X1 U854 ( .A1(n1047), .A2(n1042), .A3(KEYINPUT30), .ZN(n1183) );
INV_X1 U855 ( .A(n1186), .ZN(n1042) );
NAND2_X1 U856 ( .A1(n1187), .A2(n1030), .ZN(n1182) );
XOR2_X1 U857 ( .A(n1161), .B(KEYINPUT60), .Z(n1187) );
NOR2_X1 U858 ( .A1(n1188), .A2(G952), .ZN(n1096) );
XOR2_X1 U859 ( .A(KEYINPUT38), .B(n1078), .Z(n1188) );
XNOR2_X1 U860 ( .A(G146), .B(n1189), .ZN(G48) );
NAND2_X1 U861 ( .A1(KEYINPUT62), .A2(n1190), .ZN(n1189) );
INV_X1 U862 ( .A(n1173), .ZN(n1190) );
NAND3_X1 U863 ( .A1(n1191), .A2(n1047), .A3(n1192), .ZN(n1173) );
XOR2_X1 U864 ( .A(n1193), .B(n1174), .Z(G45) );
NAND4_X1 U865 ( .A1(n1031), .A2(n1191), .A3(n1162), .A4(n1163), .ZN(n1174) );
XOR2_X1 U866 ( .A(G140), .B(n1194), .Z(G42) );
NOR2_X1 U867 ( .A1(n1185), .A2(n1195), .ZN(n1194) );
XOR2_X1 U868 ( .A(G137), .B(n1196), .Z(G39) );
NOR3_X1 U869 ( .A1(n1197), .A2(n1161), .A3(n1195), .ZN(n1196) );
XOR2_X1 U870 ( .A(KEYINPUT23), .B(n1030), .Z(n1197) );
XOR2_X1 U871 ( .A(G134), .B(n1198), .Z(G36) );
NOR2_X1 U872 ( .A1(n1195), .A2(n1164), .ZN(n1198) );
XOR2_X1 U873 ( .A(n1177), .B(n1199), .Z(G33) );
NAND2_X1 U874 ( .A1(KEYINPUT37), .A2(G131), .ZN(n1199) );
NAND3_X1 U875 ( .A1(n1180), .A2(n1047), .A3(n1031), .ZN(n1177) );
INV_X1 U876 ( .A(n1195), .ZN(n1180) );
NAND3_X1 U877 ( .A1(n1018), .A2(n1038), .A3(n1200), .ZN(n1195) );
AND3_X1 U878 ( .A1(n1024), .A2(n1201), .A3(n1040), .ZN(n1200) );
NAND2_X1 U879 ( .A1(n1202), .A2(n1203), .ZN(G30) );
NAND2_X1 U880 ( .A1(G128), .A2(n1179), .ZN(n1203) );
XOR2_X1 U881 ( .A(n1204), .B(KEYINPUT46), .Z(n1202) );
OR2_X1 U882 ( .A1(n1179), .A2(G128), .ZN(n1204) );
NAND3_X1 U883 ( .A1(n1191), .A2(n1048), .A3(n1192), .ZN(n1179) );
AND4_X1 U884 ( .A1(n1038), .A2(n1017), .A3(n1040), .A4(n1201), .ZN(n1191) );
NAND2_X1 U885 ( .A1(n1205), .A2(n1206), .ZN(G3) );
NAND2_X1 U886 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U887 ( .A(n1209), .B(n1210), .Z(n1205) );
NOR2_X1 U888 ( .A1(n1208), .A2(n1207), .ZN(n1210) );
XOR2_X1 U889 ( .A(KEYINPUT11), .B(G101), .Z(n1207) );
INV_X1 U890 ( .A(KEYINPUT15), .ZN(n1208) );
NAND3_X1 U891 ( .A1(n1031), .A2(n1172), .A3(n1030), .ZN(n1209) );
XOR2_X1 U892 ( .A(n1211), .B(n1178), .Z(G27) );
NAND4_X1 U893 ( .A1(n1032), .A2(n1212), .A3(n1017), .A4(n1201), .ZN(n1178) );
NAND2_X1 U894 ( .A1(n1213), .A2(n1049), .ZN(n1201) );
NAND3_X1 U895 ( .A1(G902), .A2(n1214), .A3(n1069), .ZN(n1213) );
NOR2_X1 U896 ( .A1(n1078), .A2(G900), .ZN(n1069) );
INV_X1 U897 ( .A(n1185), .ZN(n1212) );
NAND2_X1 U898 ( .A1(n1186), .A2(n1047), .ZN(n1185) );
XOR2_X1 U899 ( .A(n1215), .B(n1216), .Z(G24) );
XOR2_X1 U900 ( .A(KEYINPUT32), .B(G122), .Z(n1216) );
NAND4_X1 U901 ( .A1(n1217), .A2(n1218), .A3(n1162), .A4(n1163), .ZN(n1215) );
XNOR2_X1 U902 ( .A(n1050), .B(KEYINPUT1), .ZN(n1163) );
XOR2_X1 U903 ( .A(n1116), .B(KEYINPUT61), .Z(n1217) );
INV_X1 U904 ( .A(n1037), .ZN(n1116) );
NOR2_X1 U905 ( .A1(n1219), .A2(n1220), .ZN(n1037) );
XOR2_X1 U906 ( .A(n1221), .B(n1222), .Z(G21) );
NAND3_X1 U907 ( .A1(n1030), .A2(n1192), .A3(n1218), .ZN(n1222) );
INV_X1 U908 ( .A(n1161), .ZN(n1192) );
NAND2_X1 U909 ( .A1(n1220), .A2(n1219), .ZN(n1161) );
INV_X1 U910 ( .A(n1223), .ZN(n1220) );
XOR2_X1 U911 ( .A(G116), .B(n1224), .Z(G18) );
NOR2_X1 U912 ( .A1(n1156), .A2(n1164), .ZN(n1224) );
NAND2_X1 U913 ( .A1(n1031), .A2(n1048), .ZN(n1164) );
NOR2_X1 U914 ( .A1(n1050), .A2(n1162), .ZN(n1048) );
XNOR2_X1 U915 ( .A(G113), .B(n1150), .ZN(G15) );
NAND3_X1 U916 ( .A1(n1031), .A2(n1047), .A3(n1218), .ZN(n1150) );
INV_X1 U917 ( .A(n1156), .ZN(n1218) );
NAND2_X1 U918 ( .A1(n1032), .A2(n1225), .ZN(n1156) );
NOR2_X1 U919 ( .A1(n1038), .A2(n1053), .ZN(n1032) );
INV_X1 U920 ( .A(n1040), .ZN(n1053) );
INV_X1 U921 ( .A(n1114), .ZN(n1047) );
NAND2_X1 U922 ( .A1(n1226), .A2(n1162), .ZN(n1114) );
XOR2_X1 U923 ( .A(n1050), .B(KEYINPUT54), .Z(n1226) );
INV_X1 U924 ( .A(n1044), .ZN(n1031) );
NAND2_X1 U925 ( .A1(n1223), .A2(n1219), .ZN(n1044) );
XOR2_X1 U926 ( .A(n1227), .B(n1149), .Z(G12) );
NAND3_X1 U927 ( .A1(n1186), .A2(n1172), .A3(n1030), .ZN(n1149) );
NOR2_X1 U928 ( .A1(n1228), .A2(n1162), .ZN(n1030) );
XOR2_X1 U929 ( .A(n1057), .B(n1229), .Z(n1162) );
NOR2_X1 U930 ( .A1(G475), .A2(KEYINPUT0), .ZN(n1229) );
NAND2_X1 U931 ( .A1(n1230), .A2(n1231), .ZN(n1057) );
XOR2_X1 U932 ( .A(KEYINPUT20), .B(n1111), .Z(n1230) );
XNOR2_X1 U933 ( .A(n1232), .B(n1233), .ZN(n1111) );
XOR2_X1 U934 ( .A(G104), .B(n1234), .Z(n1233) );
XOR2_X1 U935 ( .A(G122), .B(G113), .Z(n1234) );
XOR2_X1 U936 ( .A(n1235), .B(n1236), .Z(n1232) );
XOR2_X1 U937 ( .A(n1237), .B(n1238), .Z(n1236) );
NAND2_X1 U938 ( .A1(G214), .A2(n1239), .ZN(n1238) );
NAND2_X1 U939 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
OR2_X1 U940 ( .A1(n1211), .A2(G140), .ZN(n1241) );
XOR2_X1 U941 ( .A(n1242), .B(KEYINPUT52), .Z(n1240) );
NAND2_X1 U942 ( .A1(G140), .A2(n1211), .ZN(n1242) );
INV_X1 U943 ( .A(n1050), .ZN(n1228) );
XOR2_X1 U944 ( .A(n1243), .B(G478), .Z(n1050) );
OR2_X1 U945 ( .A1(n1104), .A2(G902), .ZN(n1243) );
XNOR2_X1 U946 ( .A(n1244), .B(n1245), .ZN(n1104) );
XOR2_X1 U947 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U948 ( .A(G122), .B(G116), .Z(n1247) );
XOR2_X1 U949 ( .A(G134), .B(G128), .Z(n1246) );
XOR2_X1 U950 ( .A(n1248), .B(n1249), .Z(n1244) );
XNOR2_X1 U951 ( .A(G107), .B(n1250), .ZN(n1249) );
NAND2_X1 U952 ( .A1(n1251), .A2(G217), .ZN(n1250) );
NAND2_X1 U953 ( .A1(KEYINPUT12), .A2(n1193), .ZN(n1248) );
INV_X1 U954 ( .A(n1115), .ZN(n1172) );
NAND3_X1 U955 ( .A1(n1038), .A2(n1040), .A3(n1225), .ZN(n1115) );
INV_X1 U956 ( .A(n1166), .ZN(n1225) );
NAND2_X1 U957 ( .A1(n1017), .A2(n1252), .ZN(n1166) );
NAND2_X1 U958 ( .A1(n1049), .A2(n1253), .ZN(n1252) );
NAND3_X1 U959 ( .A1(n1088), .A2(n1214), .A3(G902), .ZN(n1253) );
NOR2_X1 U960 ( .A1(n1078), .A2(G898), .ZN(n1088) );
NAND3_X1 U961 ( .A1(n1214), .A2(n1078), .A3(G952), .ZN(n1049) );
NAND2_X1 U962 ( .A1(G237), .A2(G234), .ZN(n1214) );
NOR2_X1 U963 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
INV_X1 U964 ( .A(n1024), .ZN(n1019) );
NAND2_X1 U965 ( .A1(G214), .A2(n1254), .ZN(n1024) );
XNOR2_X1 U966 ( .A(n1255), .B(n1147), .ZN(n1018) );
NAND2_X1 U967 ( .A1(G210), .A2(n1254), .ZN(n1147) );
NAND2_X1 U968 ( .A1(n1256), .A2(n1231), .ZN(n1254) );
INV_X1 U969 ( .A(G237), .ZN(n1256) );
NAND2_X1 U970 ( .A1(n1257), .A2(n1231), .ZN(n1255) );
XOR2_X1 U971 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U972 ( .A(n1142), .B(n1260), .Z(n1259) );
NOR2_X1 U973 ( .A1(KEYINPUT31), .A2(n1144), .ZN(n1260) );
XOR2_X1 U974 ( .A(n1211), .B(n1261), .Z(n1144) );
INV_X1 U975 ( .A(G125), .ZN(n1211) );
NAND2_X1 U976 ( .A1(n1262), .A2(n1263), .ZN(n1142) );
NAND2_X1 U977 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
XOR2_X1 U978 ( .A(n1266), .B(KEYINPUT55), .Z(n1265) );
XOR2_X1 U979 ( .A(n1093), .B(KEYINPUT42), .Z(n1264) );
NAND2_X1 U980 ( .A1(n1267), .A2(n1268), .ZN(n1262) );
XOR2_X1 U981 ( .A(KEYINPUT25), .B(n1269), .Z(n1268) );
INV_X1 U982 ( .A(n1266), .ZN(n1269) );
XOR2_X1 U983 ( .A(n1270), .B(n1271), .Z(n1266) );
XOR2_X1 U984 ( .A(KEYINPUT2), .B(n1091), .Z(n1271) );
INV_X1 U985 ( .A(n1090), .ZN(n1091) );
NAND2_X1 U986 ( .A1(n1272), .A2(n1273), .ZN(n1090) );
NAND2_X1 U987 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XNOR2_X1 U988 ( .A(G101), .B(KEYINPUT45), .ZN(n1274) );
XNOR2_X1 U989 ( .A(n1276), .B(KEYINPUT49), .ZN(n1272) );
NAND2_X1 U990 ( .A1(n1277), .A2(KEYINPUT17), .ZN(n1270) );
XNOR2_X1 U991 ( .A(n1094), .B(KEYINPUT29), .ZN(n1277) );
XNOR2_X1 U992 ( .A(n1278), .B(n1279), .ZN(n1094) );
XOR2_X1 U993 ( .A(KEYINPUT57), .B(G110), .Z(n1279) );
NAND2_X1 U994 ( .A1(n1280), .A2(KEYINPUT4), .ZN(n1278) );
XNOR2_X1 U995 ( .A(G122), .B(KEYINPUT16), .ZN(n1280) );
XNOR2_X1 U996 ( .A(KEYINPUT42), .B(n1093), .ZN(n1267) );
XOR2_X1 U997 ( .A(n1281), .B(n1282), .Z(n1093) );
XOR2_X1 U998 ( .A(KEYINPUT63), .B(G116), .Z(n1282) );
XOR2_X1 U999 ( .A(n1283), .B(G113), .Z(n1281) );
NAND2_X1 U1000 ( .A1(KEYINPUT36), .A2(n1221), .ZN(n1283) );
INV_X1 U1001 ( .A(G119), .ZN(n1221) );
XOR2_X1 U1002 ( .A(n1146), .B(KEYINPUT39), .Z(n1258) );
NAND2_X1 U1003 ( .A1(n1284), .A2(n1078), .ZN(n1146) );
XOR2_X1 U1004 ( .A(KEYINPUT26), .B(G224), .Z(n1284) );
NAND2_X1 U1005 ( .A1(G221), .A2(n1285), .ZN(n1040) );
XOR2_X1 U1006 ( .A(n1056), .B(KEYINPUT56), .Z(n1038) );
XOR2_X1 U1007 ( .A(n1286), .B(G469), .Z(n1056) );
NAND2_X1 U1008 ( .A1(n1287), .A2(n1231), .ZN(n1286) );
XOR2_X1 U1009 ( .A(n1288), .B(n1289), .Z(n1287) );
NOR2_X1 U1010 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NOR2_X1 U1011 ( .A1(KEYINPUT22), .A2(n1135), .ZN(n1291) );
INV_X1 U1012 ( .A(n1292), .ZN(n1135) );
NOR2_X1 U1013 ( .A1(KEYINPUT48), .A2(n1292), .ZN(n1290) );
NAND2_X1 U1014 ( .A1(G227), .A2(n1078), .ZN(n1292) );
XOR2_X1 U1015 ( .A(n1133), .B(KEYINPUT58), .Z(n1288) );
XOR2_X1 U1016 ( .A(n1293), .B(n1294), .Z(n1133) );
XOR2_X1 U1017 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1018 ( .A(n1227), .B(G140), .Z(n1296) );
NAND2_X1 U1019 ( .A1(n1297), .A2(n1298), .ZN(n1295) );
NAND2_X1 U1020 ( .A1(G101), .A2(n1275), .ZN(n1298) );
XOR2_X1 U1021 ( .A(KEYINPUT21), .B(n1276), .Z(n1297) );
NOR2_X1 U1022 ( .A1(n1275), .A2(G101), .ZN(n1276) );
XOR2_X1 U1023 ( .A(G104), .B(G107), .Z(n1275) );
XOR2_X1 U1024 ( .A(n1071), .B(n1299), .Z(n1293) );
XOR2_X1 U1025 ( .A(n1235), .B(n1300), .Z(n1071) );
XNOR2_X1 U1026 ( .A(n1301), .B(KEYINPUT19), .ZN(n1300) );
NAND2_X1 U1027 ( .A1(KEYINPUT44), .A2(n1302), .ZN(n1301) );
XOR2_X1 U1028 ( .A(KEYINPUT14), .B(G128), .Z(n1302) );
XNOR2_X1 U1029 ( .A(G131), .B(n1303), .ZN(n1235) );
XOR2_X1 U1030 ( .A(G146), .B(G143), .Z(n1303) );
NOR2_X1 U1031 ( .A1(n1219), .A2(n1223), .ZN(n1186) );
XNOR2_X1 U1032 ( .A(n1304), .B(n1100), .ZN(n1223) );
NAND2_X1 U1033 ( .A1(G217), .A2(n1285), .ZN(n1100) );
NAND2_X1 U1034 ( .A1(G234), .A2(n1231), .ZN(n1285) );
NAND2_X1 U1035 ( .A1(n1098), .A2(n1231), .ZN(n1304) );
XNOR2_X1 U1036 ( .A(n1305), .B(n1306), .ZN(n1098) );
XOR2_X1 U1037 ( .A(n1307), .B(n1308), .Z(n1306) );
XOR2_X1 U1038 ( .A(G128), .B(G119), .Z(n1308) );
XOR2_X1 U1039 ( .A(G146), .B(G137), .Z(n1307) );
XNOR2_X1 U1040 ( .A(n1309), .B(n1075), .ZN(n1305) );
XNOR2_X1 U1041 ( .A(G125), .B(G140), .ZN(n1075) );
XOR2_X1 U1042 ( .A(n1310), .B(G110), .Z(n1309) );
NAND2_X1 U1043 ( .A1(G221), .A2(n1251), .ZN(n1310) );
AND2_X1 U1044 ( .A1(G234), .A2(n1078), .ZN(n1251) );
INV_X1 U1045 ( .A(G953), .ZN(n1078) );
XNOR2_X1 U1046 ( .A(n1311), .B(G472), .ZN(n1219) );
NAND2_X1 U1047 ( .A1(n1312), .A2(n1231), .ZN(n1311) );
INV_X1 U1048 ( .A(G902), .ZN(n1231) );
XNOR2_X1 U1049 ( .A(n1313), .B(n1120), .ZN(n1312) );
XOR2_X1 U1050 ( .A(n1314), .B(G101), .Z(n1120) );
NAND2_X1 U1051 ( .A1(G210), .A2(n1239), .ZN(n1314) );
NOR2_X1 U1052 ( .A1(G953), .A2(G237), .ZN(n1239) );
NOR2_X1 U1053 ( .A1(n1124), .A2(n1315), .ZN(n1313) );
XOR2_X1 U1054 ( .A(n1316), .B(KEYINPUT40), .Z(n1315) );
NAND2_X1 U1055 ( .A1(n1317), .A2(n1129), .ZN(n1316) );
XOR2_X1 U1056 ( .A(n1127), .B(KEYINPUT53), .Z(n1317) );
NOR2_X1 U1057 ( .A1(n1129), .A2(n1127), .ZN(n1124) );
XOR2_X1 U1058 ( .A(n1261), .B(n1318), .Z(n1127) );
XOR2_X1 U1059 ( .A(G131), .B(n1299), .Z(n1318) );
XNOR2_X1 U1060 ( .A(n1319), .B(KEYINPUT27), .ZN(n1299) );
NAND2_X1 U1061 ( .A1(KEYINPUT59), .A2(n1074), .ZN(n1319) );
XOR2_X1 U1062 ( .A(G134), .B(G137), .Z(n1074) );
XOR2_X1 U1063 ( .A(n1320), .B(n1321), .Z(n1261) );
NOR2_X1 U1064 ( .A1(G146), .A2(KEYINPUT47), .ZN(n1321) );
XOR2_X1 U1065 ( .A(n1193), .B(G128), .Z(n1320) );
INV_X1 U1066 ( .A(G143), .ZN(n1193) );
XOR2_X1 U1067 ( .A(G113), .B(n1322), .Z(n1129) );
XOR2_X1 U1068 ( .A(G119), .B(G116), .Z(n1322) );
INV_X1 U1069 ( .A(G110), .ZN(n1227) );
endmodule


