//Key = 1100010100101110011110000101110000001011000000100011111001111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429;

XOR2_X1 U787 ( .A(n1090), .B(n1091), .Z(G9) );
NAND4_X1 U788 ( .A1(KEYINPUT39), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1091) );
NOR2_X1 U789 ( .A1(n1095), .A2(n1096), .ZN(G75) );
XOR2_X1 U790 ( .A(KEYINPUT24), .B(n1097), .Z(n1096) );
NOR3_X1 U791 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1097) );
NOR2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NOR2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
INV_X1 U795 ( .A(n1107), .ZN(n1106) );
NOR2_X1 U796 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
NOR2_X1 U797 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR2_X1 U798 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NOR2_X1 U799 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U800 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NOR2_X1 U801 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NOR2_X1 U802 ( .A1(n1120), .A2(n1121), .ZN(n1112) );
NOR2_X1 U803 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
NOR2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
XOR2_X1 U805 ( .A(n1126), .B(KEYINPUT49), .Z(n1124) );
NOR3_X1 U806 ( .A1(n1121), .A2(n1127), .A3(n1115), .ZN(n1108) );
NOR2_X1 U807 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR4_X1 U808 ( .A1(n1130), .A2(n1111), .A3(n1115), .A4(n1121), .ZN(n1103) );
NOR2_X1 U809 ( .A1(G952), .A2(n1100), .ZN(n1095) );
NAND2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1100) );
NAND4_X1 U811 ( .A1(n1133), .A2(n1125), .A3(n1134), .A4(n1135), .ZN(n1132) );
NOR4_X1 U812 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1135) );
XOR2_X1 U813 ( .A(n1140), .B(n1141), .Z(n1138) );
NOR2_X1 U814 ( .A1(G472), .A2(KEYINPUT34), .ZN(n1141) );
NAND3_X1 U815 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1136) );
XNOR2_X1 U816 ( .A(n1145), .B(n1146), .ZN(n1144) );
NAND3_X1 U817 ( .A1(G475), .A2(n1147), .A3(n1148), .ZN(n1143) );
OR2_X1 U818 ( .A1(n1148), .A2(G475), .ZN(n1142) );
INV_X1 U819 ( .A(KEYINPUT23), .ZN(n1148) );
NOR3_X1 U820 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1134) );
INV_X1 U821 ( .A(n1119), .ZN(n1149) );
NAND2_X1 U822 ( .A1(G469), .A2(n1152), .ZN(n1133) );
XOR2_X1 U823 ( .A(n1153), .B(n1154), .Z(G72) );
XOR2_X1 U824 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U825 ( .A1(n1157), .A2(G953), .ZN(n1156) );
NAND4_X1 U826 ( .A1(KEYINPUT5), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1155) );
NAND2_X1 U827 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U828 ( .A1(G953), .A2(n1163), .ZN(n1159) );
XOR2_X1 U829 ( .A(KEYINPUT28), .B(n1164), .Z(n1158) );
NOR2_X1 U830 ( .A1(n1161), .A2(n1162), .ZN(n1164) );
NAND2_X1 U831 ( .A1(n1165), .A2(n1166), .ZN(n1162) );
NAND2_X1 U832 ( .A1(G140), .A2(n1167), .ZN(n1166) );
XOR2_X1 U833 ( .A(n1168), .B(KEYINPUT56), .Z(n1165) );
NAND2_X1 U834 ( .A1(G125), .A2(n1169), .ZN(n1168) );
XOR2_X1 U835 ( .A(n1170), .B(n1171), .Z(n1161) );
XOR2_X1 U836 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U837 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XOR2_X1 U838 ( .A(n1176), .B(KEYINPUT52), .Z(n1175) );
NAND2_X1 U839 ( .A1(G131), .A2(n1177), .ZN(n1176) );
NOR2_X1 U840 ( .A1(G131), .A2(n1177), .ZN(n1174) );
XOR2_X1 U841 ( .A(G137), .B(G134), .Z(n1177) );
XOR2_X1 U842 ( .A(n1178), .B(G143), .Z(n1170) );
NAND2_X1 U843 ( .A1(G953), .A2(n1179), .ZN(n1153) );
NAND2_X1 U844 ( .A1(G900), .A2(G227), .ZN(n1179) );
XOR2_X1 U845 ( .A(n1180), .B(n1181), .Z(G69) );
NOR3_X1 U846 ( .A1(n1131), .A2(KEYINPUT35), .A3(n1182), .ZN(n1181) );
AND2_X1 U847 ( .A1(G224), .A2(G898), .ZN(n1182) );
NAND2_X1 U848 ( .A1(n1183), .A2(n1184), .ZN(n1180) );
NAND2_X1 U849 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U850 ( .A(n1187), .B(KEYINPUT16), .Z(n1183) );
OR2_X1 U851 ( .A1(n1186), .A2(n1185), .ZN(n1187) );
AND3_X1 U852 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1185) );
XOR2_X1 U853 ( .A(KEYINPUT51), .B(n1191), .Z(n1190) );
NOR2_X1 U854 ( .A1(G898), .A2(n1131), .ZN(n1191) );
NAND2_X1 U855 ( .A1(n1192), .A2(n1193), .ZN(n1189) );
NAND2_X1 U856 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NAND3_X1 U857 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1188) );
INV_X1 U858 ( .A(n1192), .ZN(n1196) );
XNOR2_X1 U859 ( .A(KEYINPUT53), .B(n1197), .ZN(n1194) );
NAND2_X1 U860 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U861 ( .A(KEYINPUT46), .B(n1200), .Z(n1199) );
NAND2_X1 U862 ( .A1(n1131), .A2(n1201), .ZN(n1186) );
NAND2_X1 U863 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NOR2_X1 U864 ( .A1(n1204), .A2(n1205), .ZN(G66) );
XOR2_X1 U865 ( .A(n1206), .B(n1207), .Z(n1205) );
NAND3_X1 U866 ( .A1(n1208), .A2(G217), .A3(KEYINPUT0), .ZN(n1206) );
NOR2_X1 U867 ( .A1(n1204), .A2(n1209), .ZN(G63) );
XOR2_X1 U868 ( .A(n1210), .B(n1211), .Z(n1209) );
NAND3_X1 U869 ( .A1(n1212), .A2(n1213), .A3(G478), .ZN(n1210) );
OR2_X1 U870 ( .A1(n1214), .A2(n1208), .ZN(n1213) );
NAND2_X1 U871 ( .A1(n1215), .A2(n1214), .ZN(n1212) );
INV_X1 U872 ( .A(KEYINPUT59), .ZN(n1214) );
NAND2_X1 U873 ( .A1(n1216), .A2(G902), .ZN(n1215) );
NOR2_X1 U874 ( .A1(n1204), .A2(n1217), .ZN(G60) );
XOR2_X1 U875 ( .A(n1218), .B(n1219), .Z(n1217) );
NAND2_X1 U876 ( .A1(n1208), .A2(G475), .ZN(n1218) );
NAND3_X1 U877 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(G6) );
OR2_X1 U878 ( .A1(n1203), .A2(G104), .ZN(n1222) );
NAND2_X1 U879 ( .A1(KEYINPUT43), .A2(n1223), .ZN(n1221) );
NAND2_X1 U880 ( .A1(G104), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U881 ( .A(KEYINPUT27), .B(n1203), .ZN(n1224) );
NAND2_X1 U882 ( .A1(n1225), .A2(n1226), .ZN(n1220) );
INV_X1 U883 ( .A(KEYINPUT43), .ZN(n1226) );
NAND2_X1 U884 ( .A1(n1227), .A2(n1228), .ZN(n1225) );
NAND3_X1 U885 ( .A1(KEYINPUT27), .A2(G104), .A3(n1203), .ZN(n1228) );
OR2_X1 U886 ( .A1(n1203), .A2(KEYINPUT27), .ZN(n1227) );
NOR2_X1 U887 ( .A1(n1204), .A2(n1229), .ZN(G57) );
NOR2_X1 U888 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U889 ( .A(n1232), .B(KEYINPUT18), .Z(n1231) );
NAND2_X1 U890 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NOR2_X1 U891 ( .A1(n1233), .A2(n1234), .ZN(n1230) );
XOR2_X1 U892 ( .A(G101), .B(n1235), .Z(n1234) );
NOR2_X1 U893 ( .A1(n1236), .A2(KEYINPUT15), .ZN(n1235) );
INV_X1 U894 ( .A(n1237), .ZN(n1236) );
XOR2_X1 U895 ( .A(n1238), .B(n1198), .Z(n1233) );
XOR2_X1 U896 ( .A(n1239), .B(n1240), .Z(n1238) );
NOR2_X1 U897 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
XOR2_X1 U898 ( .A(n1243), .B(KEYINPUT60), .Z(n1242) );
NAND2_X1 U899 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
NOR2_X1 U900 ( .A1(n1244), .A2(n1245), .ZN(n1241) );
NAND2_X1 U901 ( .A1(n1208), .A2(G472), .ZN(n1239) );
NOR2_X1 U902 ( .A1(n1246), .A2(n1247), .ZN(G54) );
XOR2_X1 U903 ( .A(KEYINPUT6), .B(n1204), .Z(n1247) );
XOR2_X1 U904 ( .A(n1248), .B(n1249), .Z(n1246) );
XOR2_X1 U905 ( .A(n1250), .B(n1251), .Z(n1248) );
NOR2_X1 U906 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
XOR2_X1 U907 ( .A(KEYINPUT21), .B(n1254), .Z(n1253) );
NOR2_X1 U908 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
AND2_X1 U909 ( .A1(n1255), .A2(n1256), .ZN(n1252) );
XNOR2_X1 U910 ( .A(n1169), .B(KEYINPUT48), .ZN(n1256) );
NAND2_X1 U911 ( .A1(n1208), .A2(G469), .ZN(n1250) );
NOR3_X1 U912 ( .A1(n1204), .A2(n1257), .A3(n1258), .ZN(G51) );
NOR2_X1 U913 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
XOR2_X1 U914 ( .A(n1261), .B(n1262), .Z(n1260) );
NOR2_X1 U915 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
INV_X1 U916 ( .A(KEYINPUT50), .ZN(n1259) );
NOR2_X1 U917 ( .A1(KEYINPUT50), .A2(n1265), .ZN(n1257) );
XOR2_X1 U918 ( .A(n1261), .B(n1266), .Z(n1265) );
NOR2_X1 U919 ( .A1(n1267), .A2(n1264), .ZN(n1266) );
INV_X1 U920 ( .A(KEYINPUT54), .ZN(n1264) );
XOR2_X1 U921 ( .A(n1268), .B(n1269), .Z(n1261) );
AND2_X1 U922 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U923 ( .A1(n1208), .A2(n1146), .ZN(n1268) );
NOR2_X1 U924 ( .A1(n1272), .A2(n1216), .ZN(n1208) );
INV_X1 U925 ( .A(n1098), .ZN(n1216) );
NAND3_X1 U926 ( .A1(n1202), .A2(n1273), .A3(n1157), .ZN(n1098) );
AND4_X1 U927 ( .A1(n1274), .A2(n1275), .A3(n1276), .A4(n1277), .ZN(n1157) );
NOR2_X1 U928 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NOR2_X1 U929 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NOR2_X1 U930 ( .A1(n1282), .A2(n1283), .ZN(n1280) );
NOR2_X1 U931 ( .A1(n1121), .A2(n1284), .ZN(n1283) );
NOR2_X1 U932 ( .A1(n1285), .A2(n1286), .ZN(n1282) );
NOR2_X1 U933 ( .A1(n1287), .A2(n1288), .ZN(n1285) );
NOR2_X1 U934 ( .A1(n1130), .A2(n1121), .ZN(n1288) );
NOR2_X1 U935 ( .A1(n1289), .A2(n1092), .ZN(n1130) );
NOR3_X1 U936 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1287) );
XNOR2_X1 U937 ( .A(KEYINPUT10), .B(n1203), .ZN(n1273) );
NAND3_X1 U938 ( .A1(n1093), .A2(n1094), .A3(n1289), .ZN(n1203) );
AND4_X1 U939 ( .A1(n1293), .A2(n1294), .A3(n1295), .A4(n1296), .ZN(n1202) );
AND4_X1 U940 ( .A1(n1297), .A2(n1298), .A3(n1299), .A4(n1300), .ZN(n1296) );
OR2_X1 U941 ( .A1(n1301), .A2(n1290), .ZN(n1295) );
NAND3_X1 U942 ( .A1(n1302), .A2(n1303), .A3(KEYINPUT57), .ZN(n1294) );
NAND2_X1 U943 ( .A1(n1304), .A2(n1305), .ZN(n1293) );
NAND2_X1 U944 ( .A1(n1306), .A2(n1307), .ZN(n1304) );
NAND4_X1 U945 ( .A1(n1308), .A2(n1092), .A3(n1093), .A4(n1123), .ZN(n1307) );
XOR2_X1 U946 ( .A(n1290), .B(KEYINPUT19), .Z(n1308) );
OR4_X1 U947 ( .A1(n1284), .A2(n1290), .A3(n1309), .A4(KEYINPUT57), .ZN(n1306) );
NOR2_X1 U948 ( .A1(n1131), .A2(G952), .ZN(n1204) );
XOR2_X1 U949 ( .A(G146), .B(n1278), .Z(G48) );
AND2_X1 U950 ( .A1(n1310), .A2(n1289), .ZN(n1278) );
XNOR2_X1 U951 ( .A(G143), .B(n1311), .ZN(G45) );
NAND4_X1 U952 ( .A1(n1128), .A2(n1117), .A3(n1312), .A4(n1313), .ZN(n1311) );
NOR3_X1 U953 ( .A1(n1314), .A2(n1291), .A3(n1292), .ZN(n1313) );
XNOR2_X1 U954 ( .A(n1315), .B(KEYINPUT44), .ZN(n1312) );
XOR2_X1 U955 ( .A(n1169), .B(n1276), .Z(G42) );
NAND4_X1 U956 ( .A1(n1316), .A2(n1317), .A3(n1129), .A4(n1289), .ZN(n1276) );
INV_X1 U957 ( .A(n1121), .ZN(n1316) );
XOR2_X1 U958 ( .A(G137), .B(n1318), .Z(G39) );
NOR3_X1 U959 ( .A1(n1284), .A2(n1319), .A3(n1281), .ZN(n1318) );
XOR2_X1 U960 ( .A(n1121), .B(KEYINPUT26), .Z(n1319) );
XNOR2_X1 U961 ( .A(G134), .B(n1320), .ZN(G36) );
NAND2_X1 U962 ( .A1(n1321), .A2(n1092), .ZN(n1320) );
XOR2_X1 U963 ( .A(n1322), .B(n1323), .Z(G33) );
NAND2_X1 U964 ( .A1(KEYINPUT14), .A2(G131), .ZN(n1323) );
NAND2_X1 U965 ( .A1(n1321), .A2(n1324), .ZN(n1322) );
XOR2_X1 U966 ( .A(KEYINPUT40), .B(n1289), .Z(n1324) );
NOR3_X1 U967 ( .A1(n1121), .A2(n1281), .A3(n1286), .ZN(n1321) );
INV_X1 U968 ( .A(n1317), .ZN(n1281) );
NAND2_X1 U969 ( .A1(n1325), .A2(n1119), .ZN(n1121) );
XOR2_X1 U970 ( .A(n1326), .B(G128), .Z(G30) );
NAND2_X1 U971 ( .A1(KEYINPUT12), .A2(n1274), .ZN(n1326) );
NAND2_X1 U972 ( .A1(n1310), .A2(n1092), .ZN(n1274) );
AND4_X1 U973 ( .A1(n1317), .A2(n1117), .A3(n1327), .A4(n1137), .ZN(n1310) );
NOR2_X1 U974 ( .A1(n1314), .A2(n1315), .ZN(n1317) );
XOR2_X1 U975 ( .A(n1328), .B(n1329), .Z(G3) );
NAND2_X1 U976 ( .A1(n1330), .A2(n1117), .ZN(n1329) );
XOR2_X1 U977 ( .A(n1301), .B(KEYINPUT58), .Z(n1330) );
NAND4_X1 U978 ( .A1(n1107), .A2(n1128), .A3(n1123), .A4(n1305), .ZN(n1301) );
XOR2_X1 U979 ( .A(n1331), .B(G125), .Z(G27) );
NAND2_X1 U980 ( .A1(KEYINPUT29), .A2(n1275), .ZN(n1331) );
NAND4_X1 U981 ( .A1(n1129), .A2(n1289), .A3(n1332), .A4(n1309), .ZN(n1275) );
NOR2_X1 U982 ( .A1(n1315), .A2(n1290), .ZN(n1332) );
AND2_X1 U983 ( .A1(n1333), .A2(n1102), .ZN(n1315) );
NAND4_X1 U984 ( .A1(G953), .A2(G902), .A3(n1334), .A4(n1163), .ZN(n1333) );
INV_X1 U985 ( .A(G900), .ZN(n1163) );
XOR2_X1 U986 ( .A(n1335), .B(n1298), .Z(G24) );
NAND4_X1 U987 ( .A1(n1302), .A2(n1093), .A3(n1336), .A4(n1337), .ZN(n1298) );
INV_X1 U988 ( .A(n1292), .ZN(n1336) );
INV_X1 U989 ( .A(n1111), .ZN(n1093) );
NAND2_X1 U990 ( .A1(n1338), .A2(n1339), .ZN(n1111) );
XNOR2_X1 U991 ( .A(G119), .B(n1340), .ZN(G21) );
NAND2_X1 U992 ( .A1(n1302), .A2(n1303), .ZN(n1340) );
INV_X1 U993 ( .A(n1284), .ZN(n1303) );
NAND3_X1 U994 ( .A1(n1327), .A2(n1137), .A3(n1107), .ZN(n1284) );
XOR2_X1 U995 ( .A(n1297), .B(n1341), .Z(G18) );
NAND2_X1 U996 ( .A1(KEYINPUT62), .A2(G116), .ZN(n1341) );
NAND3_X1 U997 ( .A1(n1128), .A2(n1092), .A3(n1302), .ZN(n1297) );
NOR2_X1 U998 ( .A1(n1337), .A2(n1292), .ZN(n1092) );
XNOR2_X1 U999 ( .A(n1139), .B(KEYINPUT22), .ZN(n1292) );
INV_X1 U1000 ( .A(n1291), .ZN(n1337) );
XNOR2_X1 U1001 ( .A(G113), .B(n1300), .ZN(G15) );
NAND3_X1 U1002 ( .A1(n1128), .A2(n1289), .A3(n1302), .ZN(n1300) );
AND3_X1 U1003 ( .A1(n1117), .A2(n1305), .A3(n1309), .ZN(n1302) );
INV_X1 U1004 ( .A(n1115), .ZN(n1309) );
NAND2_X1 U1005 ( .A1(n1342), .A2(n1125), .ZN(n1115) );
NOR2_X1 U1006 ( .A1(n1139), .A2(n1291), .ZN(n1289) );
INV_X1 U1007 ( .A(n1286), .ZN(n1128) );
NAND2_X1 U1008 ( .A1(n1339), .A2(n1327), .ZN(n1286) );
INV_X1 U1009 ( .A(n1338), .ZN(n1327) );
XNOR2_X1 U1010 ( .A(KEYINPUT9), .B(n1137), .ZN(n1339) );
XOR2_X1 U1011 ( .A(n1255), .B(n1299), .Z(G12) );
NAND3_X1 U1012 ( .A1(n1129), .A2(n1094), .A3(n1107), .ZN(n1299) );
NOR2_X1 U1013 ( .A1(n1343), .A2(n1139), .ZN(n1107) );
XOR2_X1 U1014 ( .A(G478), .B(n1344), .Z(n1139) );
AND2_X1 U1015 ( .A1(n1272), .A2(n1211), .ZN(n1344) );
XNOR2_X1 U1016 ( .A(n1345), .B(n1346), .ZN(n1211) );
NOR2_X1 U1017 ( .A1(KEYINPUT4), .A2(n1347), .ZN(n1346) );
XOR2_X1 U1018 ( .A(n1348), .B(n1349), .Z(n1347) );
XOR2_X1 U1019 ( .A(n1350), .B(n1351), .Z(n1349) );
NOR2_X1 U1020 ( .A1(KEYINPUT33), .A2(n1090), .ZN(n1350) );
INV_X1 U1021 ( .A(G107), .ZN(n1090) );
XNOR2_X1 U1022 ( .A(G116), .B(n1352), .ZN(n1348) );
XOR2_X1 U1023 ( .A(G143), .B(G122), .Z(n1352) );
NAND2_X1 U1024 ( .A1(G217), .A2(n1353), .ZN(n1345) );
XOR2_X1 U1025 ( .A(n1291), .B(KEYINPUT20), .Z(n1343) );
NOR2_X1 U1026 ( .A1(n1354), .A2(n1151), .ZN(n1291) );
NOR2_X1 U1027 ( .A1(n1147), .A2(G475), .ZN(n1151) );
AND2_X1 U1028 ( .A1(G475), .A2(n1147), .ZN(n1354) );
NAND2_X1 U1029 ( .A1(n1219), .A2(n1272), .ZN(n1147) );
XOR2_X1 U1030 ( .A(n1355), .B(n1356), .Z(n1219) );
XNOR2_X1 U1031 ( .A(n1357), .B(n1358), .ZN(n1356) );
NOR2_X1 U1032 ( .A1(KEYINPUT8), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1033 ( .A(n1360), .B(n1361), .Z(n1359) );
XNOR2_X1 U1034 ( .A(G113), .B(G104), .ZN(n1361) );
NAND2_X1 U1035 ( .A1(KEYINPUT38), .A2(n1335), .ZN(n1360) );
NAND4_X1 U1036 ( .A1(KEYINPUT13), .A2(G214), .A3(n1362), .A4(n1131), .ZN(n1357) );
XOR2_X1 U1037 ( .A(n1363), .B(n1364), .Z(n1355) );
NAND2_X1 U1038 ( .A1(n1365), .A2(KEYINPUT25), .ZN(n1363) );
XOR2_X1 U1039 ( .A(n1366), .B(n1367), .Z(n1365) );
AND3_X1 U1040 ( .A1(n1123), .A2(n1305), .A3(n1117), .ZN(n1094) );
INV_X1 U1041 ( .A(n1290), .ZN(n1117) );
NAND2_X1 U1042 ( .A1(n1118), .A2(n1119), .ZN(n1290) );
NAND2_X1 U1043 ( .A1(G214), .A2(n1368), .ZN(n1119) );
INV_X1 U1044 ( .A(n1325), .ZN(n1118) );
XOR2_X1 U1045 ( .A(n1369), .B(n1146), .Z(n1325) );
AND2_X1 U1046 ( .A1(G210), .A2(n1368), .ZN(n1146) );
NAND2_X1 U1047 ( .A1(n1362), .A2(n1272), .ZN(n1368) );
NAND2_X1 U1048 ( .A1(KEYINPUT1), .A2(n1145), .ZN(n1369) );
AND2_X1 U1049 ( .A1(n1370), .A2(n1272), .ZN(n1145) );
XOR2_X1 U1050 ( .A(n1371), .B(n1267), .Z(n1370) );
INV_X1 U1051 ( .A(n1263), .ZN(n1267) );
XOR2_X1 U1052 ( .A(n1372), .B(n1192), .Z(n1263) );
XNOR2_X1 U1053 ( .A(n1335), .B(G110), .ZN(n1192) );
INV_X1 U1054 ( .A(G122), .ZN(n1335) );
NAND2_X1 U1055 ( .A1(n1373), .A2(n1195), .ZN(n1372) );
NAND2_X1 U1056 ( .A1(n1200), .A2(n1374), .ZN(n1195) );
XOR2_X1 U1057 ( .A(n1375), .B(KEYINPUT41), .Z(n1373) );
OR2_X1 U1058 ( .A1(n1200), .A2(n1374), .ZN(n1375) );
INV_X1 U1059 ( .A(n1198), .ZN(n1374) );
XNOR2_X1 U1060 ( .A(n1328), .B(n1376), .ZN(n1200) );
INV_X1 U1061 ( .A(G101), .ZN(n1328) );
NAND2_X1 U1062 ( .A1(n1377), .A2(n1270), .ZN(n1371) );
NAND2_X1 U1063 ( .A1(n1378), .A2(n1379), .ZN(n1270) );
NAND2_X1 U1064 ( .A1(G224), .A2(n1131), .ZN(n1379) );
XOR2_X1 U1065 ( .A(n1167), .B(n1245), .Z(n1378) );
INV_X1 U1066 ( .A(G125), .ZN(n1167) );
XOR2_X1 U1067 ( .A(n1271), .B(KEYINPUT32), .Z(n1377) );
NAND3_X1 U1068 ( .A1(G224), .A2(n1131), .A3(n1380), .ZN(n1271) );
XOR2_X1 U1069 ( .A(n1245), .B(G125), .Z(n1380) );
NAND2_X1 U1070 ( .A1(n1102), .A2(n1381), .ZN(n1305) );
NAND4_X1 U1071 ( .A1(G953), .A2(G902), .A3(n1334), .A4(n1382), .ZN(n1381) );
INV_X1 U1072 ( .A(G898), .ZN(n1382) );
NAND3_X1 U1073 ( .A1(n1334), .A2(n1131), .A3(G952), .ZN(n1102) );
NAND2_X1 U1074 ( .A1(G237), .A2(G234), .ZN(n1334) );
INV_X1 U1075 ( .A(n1314), .ZN(n1123) );
NAND2_X1 U1076 ( .A1(n1125), .A2(n1126), .ZN(n1314) );
INV_X1 U1077 ( .A(n1342), .ZN(n1126) );
NOR2_X1 U1078 ( .A1(n1383), .A2(n1150), .ZN(n1342) );
NOR2_X1 U1079 ( .A1(n1152), .A2(G469), .ZN(n1150) );
AND2_X1 U1080 ( .A1(n1384), .A2(G469), .ZN(n1383) );
XOR2_X1 U1081 ( .A(n1152), .B(KEYINPUT37), .Z(n1384) );
NAND2_X1 U1082 ( .A1(n1385), .A2(n1272), .ZN(n1152) );
XOR2_X1 U1083 ( .A(n1386), .B(n1387), .Z(n1385) );
XOR2_X1 U1084 ( .A(n1169), .B(n1388), .Z(n1387) );
XNOR2_X1 U1085 ( .A(KEYINPUT45), .B(KEYINPUT3), .ZN(n1388) );
INV_X1 U1086 ( .A(G140), .ZN(n1169) );
XOR2_X1 U1087 ( .A(n1249), .B(n1255), .Z(n1386) );
XNOR2_X1 U1088 ( .A(n1389), .B(n1390), .ZN(n1249) );
XOR2_X1 U1089 ( .A(n1391), .B(n1392), .Z(n1390) );
XOR2_X1 U1090 ( .A(n1393), .B(n1394), .Z(n1392) );
AND2_X1 U1091 ( .A1(n1131), .A2(G227), .ZN(n1394) );
NOR2_X1 U1092 ( .A1(G101), .A2(KEYINPUT55), .ZN(n1393) );
XOR2_X1 U1093 ( .A(n1395), .B(n1172), .Z(n1391) );
NOR2_X1 U1094 ( .A1(KEYINPUT11), .A2(n1366), .ZN(n1172) );
XNOR2_X1 U1095 ( .A(n1364), .B(n1396), .ZN(n1389) );
XOR2_X1 U1096 ( .A(n1351), .B(n1376), .Z(n1396) );
XOR2_X1 U1097 ( .A(G107), .B(G104), .Z(n1376) );
XOR2_X1 U1098 ( .A(G134), .B(G128), .Z(n1351) );
XOR2_X1 U1099 ( .A(G131), .B(G143), .Z(n1364) );
NAND2_X1 U1100 ( .A1(G221), .A2(n1397), .ZN(n1125) );
NAND2_X1 U1101 ( .A1(G234), .A2(n1272), .ZN(n1397) );
AND2_X1 U1102 ( .A1(n1338), .A2(n1137), .ZN(n1129) );
NAND3_X1 U1103 ( .A1(n1398), .A2(n1399), .A3(n1400), .ZN(n1137) );
OR2_X1 U1104 ( .A1(n1401), .A2(n1207), .ZN(n1400) );
NAND3_X1 U1105 ( .A1(n1207), .A2(n1401), .A3(n1272), .ZN(n1399) );
NAND2_X1 U1106 ( .A1(G217), .A2(n1402), .ZN(n1401) );
XOR2_X1 U1107 ( .A(n1403), .B(n1404), .Z(n1207) );
XOR2_X1 U1108 ( .A(n1405), .B(n1406), .Z(n1404) );
XOR2_X1 U1109 ( .A(n1407), .B(n1408), .Z(n1406) );
AND2_X1 U1110 ( .A1(n1353), .A2(G221), .ZN(n1408) );
NOR2_X1 U1111 ( .A1(n1402), .A2(G953), .ZN(n1353) );
INV_X1 U1112 ( .A(G234), .ZN(n1402) );
NOR2_X1 U1113 ( .A1(KEYINPUT61), .A2(n1409), .ZN(n1407) );
NOR2_X1 U1114 ( .A1(KEYINPUT31), .A2(n1367), .ZN(n1405) );
XOR2_X1 U1115 ( .A(G125), .B(G140), .Z(n1367) );
XOR2_X1 U1116 ( .A(n1410), .B(n1411), .Z(n1403) );
XOR2_X1 U1117 ( .A(KEYINPUT36), .B(G146), .Z(n1411) );
XOR2_X1 U1118 ( .A(n1412), .B(G110), .Z(n1410) );
NAND2_X1 U1119 ( .A1(n1413), .A2(KEYINPUT63), .ZN(n1412) );
XNOR2_X1 U1120 ( .A(G119), .B(n1414), .ZN(n1413) );
NOR2_X1 U1121 ( .A1(KEYINPUT47), .A2(n1178), .ZN(n1414) );
INV_X1 U1122 ( .A(G128), .ZN(n1178) );
NAND2_X1 U1123 ( .A1(G902), .A2(G217), .ZN(n1398) );
XOR2_X1 U1124 ( .A(n1140), .B(G472), .Z(n1338) );
NAND2_X1 U1125 ( .A1(n1415), .A2(n1272), .ZN(n1140) );
INV_X1 U1126 ( .A(G902), .ZN(n1272) );
XOR2_X1 U1127 ( .A(n1416), .B(n1417), .Z(n1415) );
XOR2_X1 U1128 ( .A(n1418), .B(n1198), .Z(n1417) );
XNOR2_X1 U1129 ( .A(G113), .B(n1419), .ZN(n1198) );
XOR2_X1 U1130 ( .A(G119), .B(G116), .Z(n1419) );
NAND2_X1 U1131 ( .A1(KEYINPUT7), .A2(n1420), .ZN(n1418) );
XOR2_X1 U1132 ( .A(n1245), .B(n1244), .Z(n1420) );
XNOR2_X1 U1133 ( .A(n1395), .B(n1421), .ZN(n1244) );
XOR2_X1 U1134 ( .A(G134), .B(G131), .Z(n1421) );
NOR2_X1 U1135 ( .A1(KEYINPUT42), .A2(n1409), .ZN(n1395) );
INV_X1 U1136 ( .A(G137), .ZN(n1409) );
NAND2_X1 U1137 ( .A1(n1422), .A2(n1423), .ZN(n1245) );
OR2_X1 U1138 ( .A1(n1424), .A2(G128), .ZN(n1423) );
XOR2_X1 U1139 ( .A(n1425), .B(KEYINPUT30), .Z(n1422) );
NAND2_X1 U1140 ( .A1(G128), .A2(n1424), .ZN(n1425) );
NAND2_X1 U1141 ( .A1(n1426), .A2(n1427), .ZN(n1424) );
NAND2_X1 U1142 ( .A1(G143), .A2(n1366), .ZN(n1427) );
XOR2_X1 U1143 ( .A(KEYINPUT17), .B(n1428), .Z(n1426) );
NOR2_X1 U1144 ( .A1(G143), .A2(n1366), .ZN(n1428) );
INV_X1 U1145 ( .A(G146), .ZN(n1366) );
XOR2_X1 U1146 ( .A(G101), .B(n1429), .Z(n1416) );
NOR2_X1 U1147 ( .A1(KEYINPUT2), .A2(n1237), .ZN(n1429) );
NAND3_X1 U1148 ( .A1(n1362), .A2(n1131), .A3(G210), .ZN(n1237) );
INV_X1 U1149 ( .A(G953), .ZN(n1131) );
INV_X1 U1150 ( .A(G237), .ZN(n1362) );
INV_X1 U1151 ( .A(G110), .ZN(n1255) );
endmodule


