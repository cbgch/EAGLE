//Key = 1001000000101000111010100101100011110010111001011010000100001010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267;

XNOR2_X1 U698 ( .A(G107), .B(n956), .ZN(G9) );
NOR2_X1 U699 ( .A1(n957), .A2(n958), .ZN(G75) );
NOR4_X1 U700 ( .A1(n959), .A2(n960), .A3(G953), .A4(n961), .ZN(n958) );
NOR4_X1 U701 ( .A1(n962), .A2(n963), .A3(n964), .A4(n965), .ZN(n960) );
NOR2_X1 U702 ( .A1(n966), .A2(n967), .ZN(n964) );
NAND4_X1 U703 ( .A1(n968), .A2(n969), .A3(n970), .A4(n971), .ZN(n962) );
NAND3_X1 U704 ( .A1(n972), .A2(n973), .A3(n974), .ZN(n971) );
NAND2_X1 U705 ( .A1(n967), .A2(n975), .ZN(n974) );
NAND4_X1 U706 ( .A1(n976), .A2(n966), .A3(n977), .A4(n978), .ZN(n975) );
NAND2_X1 U707 ( .A1(n979), .A2(n980), .ZN(n970) );
NAND2_X1 U708 ( .A1(n981), .A2(n976), .ZN(n980) );
NAND2_X1 U709 ( .A1(n982), .A2(n983), .ZN(n969) );
NAND3_X1 U710 ( .A1(n967), .A2(n978), .A3(n966), .ZN(n983) );
INV_X1 U711 ( .A(KEYINPUT59), .ZN(n978) );
OR2_X1 U712 ( .A1(n976), .A2(n981), .ZN(n968) );
NAND3_X1 U713 ( .A1(n984), .A2(n985), .A3(n986), .ZN(n959) );
NAND3_X1 U714 ( .A1(n976), .A2(n981), .A3(n987), .ZN(n985) );
NOR3_X1 U715 ( .A1(n965), .A2(n979), .A3(n988), .ZN(n987) );
NOR2_X1 U716 ( .A1(n989), .A2(n990), .ZN(n988) );
AND3_X1 U717 ( .A1(n967), .A2(n991), .A3(n966), .ZN(n981) );
NOR3_X1 U718 ( .A1(n961), .A2(G953), .A3(G952), .ZN(n957) );
AND4_X1 U719 ( .A1(n992), .A2(n993), .A3(n994), .A4(n995), .ZN(n961) );
NOR4_X1 U720 ( .A1(n996), .A2(n997), .A3(n963), .A4(n998), .ZN(n995) );
XNOR2_X1 U721 ( .A(n999), .B(n1000), .ZN(n998) );
XOR2_X1 U722 ( .A(n1001), .B(KEYINPUT49), .Z(n1000) );
INV_X1 U723 ( .A(n1002), .ZN(n963) );
NOR2_X1 U724 ( .A1(n1003), .A2(n1004), .ZN(n996) );
XNOR2_X1 U725 ( .A(n1005), .B(n1006), .ZN(n994) );
XOR2_X1 U726 ( .A(n1007), .B(KEYINPUT30), .Z(n993) );
XNOR2_X1 U727 ( .A(n1008), .B(KEYINPUT15), .ZN(n992) );
XOR2_X1 U728 ( .A(n1009), .B(n1010), .Z(G72) );
XOR2_X1 U729 ( .A(n1011), .B(n1012), .Z(n1010) );
NOR2_X1 U730 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
AND2_X1 U731 ( .A1(G227), .A2(G900), .ZN(n1013) );
NAND2_X1 U732 ( .A1(n1015), .A2(n1016), .ZN(n1011) );
NAND2_X1 U733 ( .A1(n1017), .A2(G953), .ZN(n1016) );
XNOR2_X1 U734 ( .A(n1018), .B(n1019), .ZN(n1015) );
XNOR2_X1 U735 ( .A(n1020), .B(n1021), .ZN(n1019) );
NOR4_X1 U736 ( .A1(n1022), .A2(n1023), .A3(KEYINPUT37), .A4(n1024), .ZN(n1021) );
AND2_X1 U737 ( .A1(n1025), .A2(KEYINPUT57), .ZN(n1024) );
NOR2_X1 U738 ( .A1(n1026), .A2(n1027), .ZN(n1023) );
NOR2_X1 U739 ( .A1(KEYINPUT54), .A2(n1025), .ZN(n1026) );
NOR4_X1 U740 ( .A1(n1028), .A2(n1025), .A3(KEYINPUT57), .A4(KEYINPUT54), .ZN(n1022) );
NAND2_X1 U741 ( .A1(n1014), .A2(n1029), .ZN(n1009) );
XOR2_X1 U742 ( .A(n1030), .B(n1031), .Z(G69) );
XOR2_X1 U743 ( .A(n1032), .B(n1033), .Z(n1031) );
NOR2_X1 U744 ( .A1(KEYINPUT6), .A2(n1034), .ZN(n1033) );
NOR3_X1 U745 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NOR2_X1 U746 ( .A1(G898), .A2(n1014), .ZN(n1037) );
NOR2_X1 U747 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
XNOR2_X1 U748 ( .A(n1040), .B(n1041), .ZN(n1039) );
XOR2_X1 U749 ( .A(KEYINPUT56), .B(n1042), .Z(n1035) );
NOR2_X1 U750 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
XNOR2_X1 U751 ( .A(n1041), .B(n1045), .ZN(n1044) );
NOR2_X1 U752 ( .A1(n984), .A2(n1046), .ZN(n1032) );
XNOR2_X1 U753 ( .A(KEYINPUT31), .B(n1014), .ZN(n1046) );
NAND2_X1 U754 ( .A1(G953), .A2(n1047), .ZN(n1030) );
NAND2_X1 U755 ( .A1(n1048), .A2(G224), .ZN(n1047) );
XNOR2_X1 U756 ( .A(G898), .B(KEYINPUT45), .ZN(n1048) );
NOR2_X1 U757 ( .A1(n1049), .A2(n1050), .ZN(G66) );
XOR2_X1 U758 ( .A(n1051), .B(n1052), .Z(n1050) );
NAND3_X1 U759 ( .A1(n1053), .A2(n999), .A3(KEYINPUT62), .ZN(n1051) );
INV_X1 U760 ( .A(n1054), .ZN(n999) );
NOR3_X1 U761 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(G63) );
AND2_X1 U762 ( .A1(KEYINPUT10), .A2(n1049), .ZN(n1057) );
NOR3_X1 U763 ( .A1(KEYINPUT10), .A2(n1014), .A3(n1058), .ZN(n1056) );
INV_X1 U764 ( .A(G952), .ZN(n1058) );
XOR2_X1 U765 ( .A(n1059), .B(n1060), .Z(n1055) );
NOR2_X1 U766 ( .A1(KEYINPUT29), .A2(n1061), .ZN(n1060) );
NAND2_X1 U767 ( .A1(n1053), .A2(G478), .ZN(n1059) );
NOR2_X1 U768 ( .A1(n1049), .A2(n1062), .ZN(G60) );
NOR2_X1 U769 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U770 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U771 ( .A1(n1067), .A2(n1068), .ZN(n1063) );
XOR2_X1 U772 ( .A(KEYINPUT34), .B(n1066), .Z(n1068) );
XNOR2_X1 U773 ( .A(n1069), .B(KEYINPUT52), .ZN(n1066) );
XNOR2_X1 U774 ( .A(n1065), .B(KEYINPUT46), .ZN(n1067) );
AND2_X1 U775 ( .A1(n1053), .A2(G475), .ZN(n1065) );
XNOR2_X1 U776 ( .A(n1070), .B(n1071), .ZN(G6) );
XNOR2_X1 U777 ( .A(G104), .B(KEYINPUT8), .ZN(n1071) );
NOR2_X1 U778 ( .A1(n1049), .A2(n1072), .ZN(G57) );
XOR2_X1 U779 ( .A(n1073), .B(n1074), .Z(n1072) );
NOR2_X1 U780 ( .A1(KEYINPUT11), .A2(n1075), .ZN(n1074) );
XOR2_X1 U781 ( .A(n1076), .B(KEYINPUT20), .Z(n1075) );
XNOR2_X1 U782 ( .A(G101), .B(n1077), .ZN(n1073) );
NOR2_X1 U783 ( .A1(KEYINPUT24), .A2(n1078), .ZN(n1077) );
XOR2_X1 U784 ( .A(n1079), .B(n1080), .Z(n1078) );
AND2_X1 U785 ( .A1(G472), .A2(n1053), .ZN(n1080) );
NOR3_X1 U786 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1079) );
NOR2_X1 U787 ( .A1(n1049), .A2(n1084), .ZN(G54) );
XOR2_X1 U788 ( .A(n1085), .B(n1086), .Z(n1084) );
XOR2_X1 U789 ( .A(n1087), .B(n1088), .Z(n1086) );
NOR2_X1 U790 ( .A1(n1004), .A2(n1089), .ZN(n1087) );
XOR2_X1 U791 ( .A(n1090), .B(KEYINPUT42), .Z(n1085) );
NAND2_X1 U792 ( .A1(KEYINPUT32), .A2(n1091), .ZN(n1090) );
NOR3_X1 U793 ( .A1(n1049), .A2(n1092), .A3(n1093), .ZN(G51) );
NOR2_X1 U794 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
XOR2_X1 U795 ( .A(n1096), .B(KEYINPUT18), .Z(n1095) );
NOR2_X1 U796 ( .A1(n1097), .A2(n1098), .ZN(n1092) );
XOR2_X1 U797 ( .A(n1096), .B(KEYINPUT2), .Z(n1098) );
NAND2_X1 U798 ( .A1(n1053), .A2(n1099), .ZN(n1096) );
INV_X1 U799 ( .A(n1089), .ZN(n1053) );
NAND2_X1 U800 ( .A1(n1100), .A2(n1101), .ZN(n1089) );
NAND2_X1 U801 ( .A1(n986), .A2(n984), .ZN(n1101) );
AND4_X1 U802 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n984) );
AND4_X1 U803 ( .A1(n1106), .A2(n1107), .A3(n956), .A4(n1108), .ZN(n1105) );
NAND3_X1 U804 ( .A1(n989), .A2(n967), .A3(n1109), .ZN(n956) );
NOR2_X1 U805 ( .A1(n1110), .A2(n1070), .ZN(n1104) );
AND3_X1 U806 ( .A1(n1109), .A2(n967), .A3(n990), .ZN(n1070) );
NAND2_X1 U807 ( .A1(n1111), .A2(n1112), .ZN(n1103) );
NAND2_X1 U808 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND3_X1 U809 ( .A1(n1115), .A2(n1116), .A3(n967), .ZN(n1114) );
INV_X1 U810 ( .A(KEYINPUT33), .ZN(n1116) );
NAND2_X1 U811 ( .A1(KEYINPUT33), .A2(n1117), .ZN(n1102) );
INV_X1 U812 ( .A(n1029), .ZN(n986) );
NAND2_X1 U813 ( .A1(n1118), .A2(n1119), .ZN(n1029) );
NOR4_X1 U814 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1119) );
AND4_X1 U815 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1118) );
XNOR2_X1 U816 ( .A(KEYINPUT21), .B(n1128), .ZN(n1100) );
INV_X1 U817 ( .A(n1094), .ZN(n1097) );
NAND2_X1 U818 ( .A1(n1129), .A2(n1130), .ZN(n1094) );
NAND2_X1 U819 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U820 ( .A(n1133), .B(KEYINPUT26), .Z(n1129) );
OR2_X1 U821 ( .A1(n1132), .A2(n1131), .ZN(n1133) );
NAND2_X1 U822 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
XOR2_X1 U823 ( .A(KEYINPUT60), .B(n1136), .Z(n1134) );
NOR2_X1 U824 ( .A1(n1014), .A2(G952), .ZN(n1049) );
XNOR2_X1 U825 ( .A(G146), .B(n1125), .ZN(G48) );
NAND2_X1 U826 ( .A1(n1137), .A2(n990), .ZN(n1125) );
XNOR2_X1 U827 ( .A(G143), .B(n1124), .ZN(G45) );
NAND4_X1 U828 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1124) );
XOR2_X1 U829 ( .A(G140), .B(n1123), .Z(G42) );
AND3_X1 U830 ( .A1(n990), .A2(n1142), .A3(n1143), .ZN(n1123) );
XNOR2_X1 U831 ( .A(G137), .B(n1144), .ZN(G39) );
NOR2_X1 U832 ( .A1(n1122), .A2(KEYINPUT39), .ZN(n1144) );
NOR2_X1 U833 ( .A1(n1113), .A2(n1145), .ZN(n1122) );
XOR2_X1 U834 ( .A(G134), .B(n1121), .Z(G36) );
AND3_X1 U835 ( .A1(n1142), .A2(n989), .A3(n1139), .ZN(n1121) );
XOR2_X1 U836 ( .A(G131), .B(n1120), .Z(G33) );
AND3_X1 U837 ( .A1(n990), .A2(n1142), .A3(n1139), .ZN(n1120) );
INV_X1 U838 ( .A(n1145), .ZN(n1142) );
NAND4_X1 U839 ( .A1(n976), .A2(n977), .A3(n1141), .A4(n1146), .ZN(n1145) );
XOR2_X1 U840 ( .A(n1127), .B(n1147), .Z(G30) );
NOR2_X1 U841 ( .A1(G128), .A2(KEYINPUT5), .ZN(n1147) );
NAND2_X1 U842 ( .A1(n1137), .A2(n989), .ZN(n1127) );
AND4_X1 U843 ( .A1(n1148), .A2(n1140), .A3(n1008), .A4(n1141), .ZN(n1137) );
XNOR2_X1 U844 ( .A(G101), .B(n1106), .ZN(G3) );
NAND3_X1 U845 ( .A1(n1002), .A2(n1109), .A3(n1139), .ZN(n1106) );
XNOR2_X1 U846 ( .A(G125), .B(n1126), .ZN(G27) );
NAND4_X1 U847 ( .A1(n1149), .A2(n1141), .A3(n990), .A4(n1150), .ZN(n1126) );
NOR2_X1 U848 ( .A1(n972), .A2(n1146), .ZN(n1150) );
NAND2_X1 U849 ( .A1(n965), .A2(n1151), .ZN(n1141) );
NAND4_X1 U850 ( .A1(n1017), .A2(G902), .A3(G953), .A4(n1152), .ZN(n1151) );
XNOR2_X1 U851 ( .A(G900), .B(KEYINPUT1), .ZN(n1017) );
XNOR2_X1 U852 ( .A(n1153), .B(n1117), .ZN(G24) );
AND3_X1 U853 ( .A1(n1138), .A2(n967), .A3(n1111), .ZN(n1117) );
AND2_X1 U854 ( .A1(n1154), .A2(n1155), .ZN(n967) );
XNOR2_X1 U855 ( .A(n1156), .B(KEYINPUT28), .ZN(n1154) );
INV_X1 U856 ( .A(n1115), .ZN(n1138) );
NAND2_X1 U857 ( .A1(n1157), .A2(n1158), .ZN(n1115) );
XOR2_X1 U858 ( .A(n1159), .B(n1160), .Z(G21) );
NOR3_X1 U859 ( .A1(n1161), .A2(KEYINPUT44), .A3(n1113), .ZN(n1160) );
NAND3_X1 U860 ( .A1(n1002), .A2(n1008), .A3(n1148), .ZN(n1113) );
XNOR2_X1 U861 ( .A(G119), .B(KEYINPUT0), .ZN(n1159) );
XNOR2_X1 U862 ( .A(G116), .B(n1162), .ZN(G18) );
NOR2_X1 U863 ( .A1(n1163), .A2(KEYINPUT36), .ZN(n1162) );
INV_X1 U864 ( .A(n1107), .ZN(n1163) );
NAND3_X1 U865 ( .A1(n1139), .A2(n989), .A3(n1111), .ZN(n1107) );
NOR2_X1 U866 ( .A1(n1158), .A2(n1164), .ZN(n989) );
XNOR2_X1 U867 ( .A(n1165), .B(n1110), .ZN(G15) );
AND3_X1 U868 ( .A1(n1139), .A2(n990), .A3(n1111), .ZN(n1110) );
INV_X1 U869 ( .A(n1161), .ZN(n1111) );
NAND3_X1 U870 ( .A1(n1149), .A2(n1166), .A3(n966), .ZN(n1161) );
INV_X1 U871 ( .A(n1146), .ZN(n966) );
AND2_X1 U872 ( .A1(n1164), .A2(n1158), .ZN(n990) );
INV_X1 U873 ( .A(n1157), .ZN(n1164) );
INV_X1 U874 ( .A(n973), .ZN(n1139) );
NAND2_X1 U875 ( .A1(n1008), .A2(n1155), .ZN(n973) );
XNOR2_X1 U876 ( .A(G110), .B(n1108), .ZN(G12) );
NAND3_X1 U877 ( .A1(n1002), .A2(n1109), .A3(n1143), .ZN(n1108) );
INV_X1 U878 ( .A(n972), .ZN(n1143) );
NAND2_X1 U879 ( .A1(n1148), .A2(n1156), .ZN(n972) );
XOR2_X1 U880 ( .A(n1008), .B(KEYINPUT17), .Z(n1156) );
XNOR2_X1 U881 ( .A(n1167), .B(G472), .ZN(n1008) );
NAND2_X1 U882 ( .A1(n1168), .A2(n1128), .ZN(n1167) );
XOR2_X1 U883 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U884 ( .A(G101), .B(n1171), .Z(n1170) );
NOR2_X1 U885 ( .A1(KEYINPUT14), .A2(n1172), .ZN(n1171) );
XOR2_X1 U886 ( .A(n1076), .B(KEYINPUT22), .Z(n1172) );
NAND2_X1 U887 ( .A1(n1173), .A2(G210), .ZN(n1076) );
NAND3_X1 U888 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1169) );
INV_X1 U889 ( .A(n1082), .ZN(n1176) );
NOR3_X1 U890 ( .A1(n1177), .A2(n1178), .A3(n1018), .ZN(n1082) );
NAND2_X1 U891 ( .A1(n1179), .A2(n1180), .ZN(n1175) );
INV_X1 U892 ( .A(KEYINPUT51), .ZN(n1180) );
OR2_X1 U893 ( .A1(n1081), .A2(n1083), .ZN(n1179) );
NOR3_X1 U894 ( .A1(n1177), .A2(n1181), .A3(n1182), .ZN(n1083) );
NAND2_X1 U895 ( .A1(n1183), .A2(n1184), .ZN(n1081) );
NAND2_X1 U896 ( .A1(n1185), .A2(n1182), .ZN(n1184) );
NAND3_X1 U897 ( .A1(n1177), .A2(n1181), .A3(n1178), .ZN(n1183) );
NAND2_X1 U898 ( .A1(KEYINPUT51), .A2(n1186), .ZN(n1174) );
XNOR2_X1 U899 ( .A(n1178), .B(n1185), .ZN(n1186) );
INV_X1 U900 ( .A(n1182), .ZN(n1178) );
NAND3_X1 U901 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1182) );
OR2_X1 U902 ( .A1(G113), .A2(KEYINPUT16), .ZN(n1188) );
NAND2_X1 U903 ( .A1(n1190), .A2(KEYINPUT16), .ZN(n1187) );
XNOR2_X1 U904 ( .A(n1155), .B(KEYINPUT23), .ZN(n1148) );
XOR2_X1 U905 ( .A(n1191), .B(n1001), .Z(n1155) );
NAND2_X1 U906 ( .A1(n1052), .A2(n1128), .ZN(n1001) );
XNOR2_X1 U907 ( .A(n1192), .B(n1193), .ZN(n1052) );
XOR2_X1 U908 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U909 ( .A(G137), .B(G119), .Z(n1195) );
AND3_X1 U910 ( .A1(n1196), .A2(G234), .A3(G221), .ZN(n1194) );
XNOR2_X1 U911 ( .A(KEYINPUT19), .B(G953), .ZN(n1196) );
XNOR2_X1 U912 ( .A(n1197), .B(n1198), .ZN(n1192) );
XOR2_X1 U913 ( .A(n1199), .B(n1200), .Z(n1197) );
NAND2_X1 U914 ( .A1(KEYINPUT48), .A2(G110), .ZN(n1199) );
NAND2_X1 U915 ( .A1(KEYINPUT27), .A2(n1054), .ZN(n1191) );
NAND2_X1 U916 ( .A1(G217), .A2(n1201), .ZN(n1054) );
AND2_X1 U917 ( .A1(n1140), .A2(n1166), .ZN(n1109) );
NAND2_X1 U918 ( .A1(n1202), .A2(n1203), .ZN(n1166) );
NAND4_X1 U919 ( .A1(G902), .A2(G953), .A3(n1152), .A4(n1204), .ZN(n1203) );
INV_X1 U920 ( .A(G898), .ZN(n1204) );
XOR2_X1 U921 ( .A(n965), .B(KEYINPUT53), .Z(n1202) );
NAND3_X1 U922 ( .A1(n1152), .A2(n1014), .A3(G952), .ZN(n965) );
NAND2_X1 U923 ( .A1(G237), .A2(G234), .ZN(n1152) );
AND2_X1 U924 ( .A1(n1149), .A2(n1146), .ZN(n1140) );
NAND2_X1 U925 ( .A1(n1205), .A2(n1007), .ZN(n1146) );
NAND2_X1 U926 ( .A1(n1003), .A2(n1004), .ZN(n1007) );
INV_X1 U927 ( .A(G469), .ZN(n1004) );
INV_X1 U928 ( .A(n1206), .ZN(n1003) );
NAND2_X1 U929 ( .A1(G469), .A2(n1206), .ZN(n1205) );
NAND3_X1 U930 ( .A1(n1207), .A2(n1208), .A3(n1128), .ZN(n1206) );
NAND2_X1 U931 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
INV_X1 U932 ( .A(KEYINPUT4), .ZN(n1210) );
XOR2_X1 U933 ( .A(n1091), .B(n1088), .Z(n1209) );
NAND3_X1 U934 ( .A1(n1088), .A2(n1091), .A3(KEYINPUT4), .ZN(n1207) );
NAND2_X1 U935 ( .A1(n1211), .A2(n1212), .ZN(n1091) );
NAND2_X1 U936 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND2_X1 U937 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND2_X1 U938 ( .A1(n1181), .A2(n1217), .ZN(n1216) );
INV_X1 U939 ( .A(n1185), .ZN(n1215) );
NOR2_X1 U940 ( .A1(n1217), .A2(n1181), .ZN(n1185) );
INV_X1 U941 ( .A(n1218), .ZN(n1213) );
NAND2_X1 U942 ( .A1(n1219), .A2(n1218), .ZN(n1211) );
XNOR2_X1 U943 ( .A(n1177), .B(n1181), .ZN(n1219) );
INV_X1 U944 ( .A(n1217), .ZN(n1177) );
XOR2_X1 U945 ( .A(n1027), .B(n1025), .Z(n1217) );
INV_X1 U946 ( .A(n1028), .ZN(n1027) );
XNOR2_X1 U947 ( .A(G134), .B(G137), .ZN(n1028) );
XNOR2_X1 U948 ( .A(n1220), .B(n1221), .ZN(n1088) );
XOR2_X1 U949 ( .A(G140), .B(G110), .Z(n1221) );
NAND2_X1 U950 ( .A1(G227), .A2(n1014), .ZN(n1220) );
NOR2_X1 U951 ( .A1(n997), .A2(n976), .ZN(n1149) );
XNOR2_X1 U952 ( .A(n1099), .B(n1222), .ZN(n976) );
NOR2_X1 U953 ( .A1(KEYINPUT13), .A2(n1006), .ZN(n1222) );
NAND2_X1 U954 ( .A1(n1223), .A2(n1128), .ZN(n1006) );
XOR2_X1 U955 ( .A(n1224), .B(n1131), .Z(n1223) );
AND2_X1 U956 ( .A1(n1225), .A2(n1226), .ZN(n1131) );
NAND2_X1 U957 ( .A1(n1227), .A2(n1045), .ZN(n1226) );
INV_X1 U958 ( .A(n1040), .ZN(n1045) );
XOR2_X1 U959 ( .A(KEYINPUT12), .B(n1228), .Z(n1227) );
NAND2_X1 U960 ( .A1(n1228), .A2(n1040), .ZN(n1225) );
XOR2_X1 U961 ( .A(n1218), .B(KEYINPUT38), .Z(n1040) );
XOR2_X1 U962 ( .A(G101), .B(n1229), .Z(n1218) );
XNOR2_X1 U963 ( .A(n1230), .B(G104), .ZN(n1229) );
XNOR2_X1 U964 ( .A(n1041), .B(n1038), .ZN(n1228) );
INV_X1 U965 ( .A(n1043), .ZN(n1038) );
XOR2_X1 U966 ( .A(n1231), .B(n1153), .Z(n1043) );
NAND2_X1 U967 ( .A1(KEYINPUT35), .A2(G110), .ZN(n1231) );
NOR2_X1 U968 ( .A1(n1232), .A2(n1190), .ZN(n1041) );
NOR2_X1 U969 ( .A1(n1165), .A2(n1233), .ZN(n1190) );
XNOR2_X1 U970 ( .A(n1189), .B(KEYINPUT63), .ZN(n1232) );
NAND2_X1 U971 ( .A1(n1233), .A2(n1165), .ZN(n1189) );
INV_X1 U972 ( .A(G113), .ZN(n1165) );
XNOR2_X1 U973 ( .A(G116), .B(G119), .ZN(n1233) );
NOR2_X1 U974 ( .A1(n1136), .A2(n1234), .ZN(n1224) );
XOR2_X1 U975 ( .A(n1135), .B(KEYINPUT40), .Z(n1234) );
NAND3_X1 U976 ( .A1(G224), .A2(n1235), .A3(n1236), .ZN(n1135) );
XNOR2_X1 U977 ( .A(n1237), .B(n1018), .ZN(n1236) );
AND2_X1 U978 ( .A1(n1238), .A2(n1239), .ZN(n1136) );
NAND2_X1 U979 ( .A1(G224), .A2(n1235), .ZN(n1239) );
XNOR2_X1 U980 ( .A(KEYINPUT50), .B(n1014), .ZN(n1235) );
XNOR2_X1 U981 ( .A(n1237), .B(n1181), .ZN(n1238) );
INV_X1 U982 ( .A(n1018), .ZN(n1181) );
XOR2_X1 U983 ( .A(G143), .B(n1200), .Z(n1018) );
XOR2_X1 U984 ( .A(G146), .B(n1240), .Z(n1200) );
INV_X1 U985 ( .A(n1005), .ZN(n1099) );
NAND2_X1 U986 ( .A1(G210), .A2(n1241), .ZN(n1005) );
INV_X1 U987 ( .A(n977), .ZN(n997) );
NOR2_X1 U988 ( .A1(n979), .A2(n982), .ZN(n977) );
INV_X1 U989 ( .A(n991), .ZN(n982) );
NAND2_X1 U990 ( .A1(G221), .A2(n1201), .ZN(n991) );
NAND2_X1 U991 ( .A1(G234), .A2(n1128), .ZN(n1201) );
AND2_X1 U992 ( .A1(G214), .A2(n1241), .ZN(n979) );
NAND2_X1 U993 ( .A1(n1242), .A2(n1128), .ZN(n1241) );
INV_X1 U994 ( .A(G237), .ZN(n1242) );
NOR2_X1 U995 ( .A1(n1157), .A2(n1158), .ZN(n1002) );
XNOR2_X1 U996 ( .A(n1243), .B(G475), .ZN(n1158) );
NAND2_X1 U997 ( .A1(n1069), .A2(n1128), .ZN(n1243) );
INV_X1 U998 ( .A(G902), .ZN(n1128) );
XOR2_X1 U999 ( .A(n1244), .B(n1245), .Z(n1069) );
XNOR2_X1 U1000 ( .A(n1020), .B(n1246), .ZN(n1245) );
XNOR2_X1 U1001 ( .A(n1247), .B(n1248), .ZN(n1246) );
NOR2_X1 U1002 ( .A1(G104), .A2(KEYINPUT58), .ZN(n1248) );
NOR2_X1 U1003 ( .A1(KEYINPUT7), .A2(n1249), .ZN(n1247) );
XOR2_X1 U1004 ( .A(n1025), .B(n1250), .Z(n1249) );
XOR2_X1 U1005 ( .A(n1251), .B(G143), .Z(n1250) );
NAND2_X1 U1006 ( .A1(n1173), .A2(G214), .ZN(n1251) );
NOR2_X1 U1007 ( .A1(G953), .A2(G237), .ZN(n1173) );
XNOR2_X1 U1008 ( .A(G131), .B(KEYINPUT3), .ZN(n1025) );
INV_X1 U1009 ( .A(n1198), .ZN(n1020) );
XOR2_X1 U1010 ( .A(G140), .B(n1252), .Z(n1198) );
INV_X1 U1011 ( .A(n1237), .ZN(n1252) );
XOR2_X1 U1012 ( .A(G125), .B(KEYINPUT55), .Z(n1237) );
XOR2_X1 U1013 ( .A(n1253), .B(n1254), .Z(n1244) );
XNOR2_X1 U1014 ( .A(n1153), .B(G113), .ZN(n1254) );
INV_X1 U1015 ( .A(G122), .ZN(n1153) );
XNOR2_X1 U1016 ( .A(G146), .B(KEYINPUT25), .ZN(n1253) );
XNOR2_X1 U1017 ( .A(n1255), .B(G478), .ZN(n1157) );
OR2_X1 U1018 ( .A1(n1061), .A2(G902), .ZN(n1255) );
XNOR2_X1 U1019 ( .A(n1256), .B(n1257), .ZN(n1061) );
XNOR2_X1 U1020 ( .A(n1258), .B(n1240), .ZN(n1257) );
XOR2_X1 U1021 ( .A(G128), .B(KEYINPUT41), .Z(n1240) );
NAND2_X1 U1022 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
OR2_X1 U1023 ( .A1(n1261), .A2(n1230), .ZN(n1260) );
XOR2_X1 U1024 ( .A(n1262), .B(KEYINPUT61), .Z(n1259) );
NAND2_X1 U1025 ( .A1(n1261), .A2(n1230), .ZN(n1262) );
INV_X1 U1026 ( .A(G107), .ZN(n1230) );
XNOR2_X1 U1027 ( .A(n1263), .B(n1264), .ZN(n1261) );
NOR2_X1 U1028 ( .A1(KEYINPUT9), .A2(n1265), .ZN(n1264) );
XNOR2_X1 U1029 ( .A(G116), .B(KEYINPUT47), .ZN(n1265) );
XNOR2_X1 U1030 ( .A(G122), .B(KEYINPUT43), .ZN(n1263) );
XOR2_X1 U1031 ( .A(n1266), .B(n1267), .Z(n1256) );
AND3_X1 U1032 ( .A1(G217), .A2(n1014), .A3(G234), .ZN(n1267) );
INV_X1 U1033 ( .A(G953), .ZN(n1014) );
XNOR2_X1 U1034 ( .A(G134), .B(G143), .ZN(n1266) );
endmodule


