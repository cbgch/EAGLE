//Key = 1011000101011001110111001101010010000000100101010110110101010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404;

XNOR2_X1 U775 ( .A(G107), .B(n1076), .ZN(G9) );
NOR2_X1 U776 ( .A1(n1077), .A2(n1078), .ZN(G75) );
NOR4_X1 U777 ( .A1(n1079), .A2(n1080), .A3(G953), .A4(n1081), .ZN(n1078) );
NOR3_X1 U778 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1080) );
NOR4_X1 U779 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1084) );
NOR2_X1 U780 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR3_X1 U781 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1089) );
NOR2_X1 U782 ( .A1(KEYINPUT39), .A2(n1094), .ZN(n1093) );
NOR2_X1 U783 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
NOR2_X1 U784 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
AND2_X1 U785 ( .A1(n1099), .A2(KEYINPUT17), .ZN(n1097) );
NOR2_X1 U786 ( .A1(n1100), .A2(n1101), .ZN(n1091) );
NOR3_X1 U787 ( .A1(n1102), .A2(n1096), .A3(n1103), .ZN(n1087) );
XNOR2_X1 U788 ( .A(KEYINPUT63), .B(n1101), .ZN(n1102) );
NOR2_X1 U789 ( .A1(n1101), .A2(n1104), .ZN(n1086) );
NOR2_X1 U790 ( .A1(n1105), .A2(n1106), .ZN(n1083) );
NOR2_X1 U791 ( .A1(n1107), .A2(n1090), .ZN(n1106) );
NOR2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U793 ( .A1(n1094), .A2(n1110), .ZN(n1109) );
INV_X1 U794 ( .A(KEYINPUT39), .ZN(n1110) );
NAND3_X1 U795 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1094) );
NOR3_X1 U796 ( .A1(n1114), .A2(KEYINPUT17), .A3(n1096), .ZN(n1108) );
NAND3_X1 U797 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1079) );
NAND3_X1 U798 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1116) );
NAND2_X1 U799 ( .A1(n1121), .A2(n1122), .ZN(n1115) );
XOR2_X1 U800 ( .A(KEYINPUT51), .B(n1120), .Z(n1122) );
NOR4_X1 U801 ( .A1(n1082), .A2(n1090), .A3(n1101), .A4(n1096), .ZN(n1120) );
INV_X1 U802 ( .A(n1112), .ZN(n1101) );
INV_X1 U803 ( .A(n1123), .ZN(n1090) );
NOR3_X1 U804 ( .A1(n1081), .A2(G953), .A3(G952), .ZN(n1077) );
AND4_X1 U805 ( .A1(n1111), .A2(n1124), .A3(n1105), .A4(n1125), .ZN(n1081) );
NOR4_X1 U806 ( .A1(n1113), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1125) );
XOR2_X1 U807 ( .A(n1129), .B(n1130), .Z(n1127) );
NAND2_X1 U808 ( .A1(KEYINPUT59), .A2(n1131), .ZN(n1129) );
XOR2_X1 U809 ( .A(n1132), .B(n1133), .Z(n1126) );
XNOR2_X1 U810 ( .A(KEYINPUT0), .B(n1134), .ZN(n1133) );
XOR2_X1 U811 ( .A(n1135), .B(n1136), .Z(G72) );
NOR2_X1 U812 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U813 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
NAND2_X1 U814 ( .A1(n1141), .A2(n1142), .ZN(n1135) );
NAND2_X1 U815 ( .A1(n1143), .A2(n1138), .ZN(n1142) );
XOR2_X1 U816 ( .A(n1144), .B(n1145), .Z(n1143) );
NAND3_X1 U817 ( .A1(G900), .A2(n1145), .A3(G953), .ZN(n1141) );
XNOR2_X1 U818 ( .A(n1146), .B(n1147), .ZN(n1145) );
NAND3_X1 U819 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1146) );
NAND2_X1 U820 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
OR3_X1 U821 ( .A1(n1152), .A2(n1151), .A3(KEYINPUT10), .ZN(n1149) );
NAND2_X1 U822 ( .A1(KEYINPUT29), .A2(n1153), .ZN(n1152) );
INV_X1 U823 ( .A(n1154), .ZN(n1153) );
NAND2_X1 U824 ( .A1(n1154), .A2(KEYINPUT10), .ZN(n1148) );
XOR2_X1 U825 ( .A(n1155), .B(n1156), .Z(n1154) );
XNOR2_X1 U826 ( .A(KEYINPUT58), .B(KEYINPUT46), .ZN(n1155) );
XOR2_X1 U827 ( .A(n1157), .B(n1158), .Z(G69) );
NOR2_X1 U828 ( .A1(n1159), .A2(n1138), .ZN(n1158) );
NOR2_X1 U829 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR2_X1 U830 ( .A1(KEYINPUT42), .A2(n1162), .ZN(n1157) );
XOR2_X1 U831 ( .A(n1163), .B(n1164), .Z(n1162) );
NAND2_X1 U832 ( .A1(KEYINPUT9), .A2(n1165), .ZN(n1164) );
NAND2_X1 U833 ( .A1(n1166), .A2(n1138), .ZN(n1165) );
NAND2_X1 U834 ( .A1(n1167), .A2(n1168), .ZN(n1163) );
NAND2_X1 U835 ( .A1(G953), .A2(n1161), .ZN(n1168) );
XOR2_X1 U836 ( .A(n1169), .B(n1170), .Z(n1167) );
XNOR2_X1 U837 ( .A(G122), .B(G110), .ZN(n1170) );
NAND2_X1 U838 ( .A1(n1171), .A2(KEYINPUT55), .ZN(n1169) );
XNOR2_X1 U839 ( .A(n1172), .B(n1173), .ZN(n1171) );
NOR2_X1 U840 ( .A1(n1174), .A2(n1175), .ZN(G66) );
XOR2_X1 U841 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U842 ( .A1(n1178), .A2(G217), .ZN(n1176) );
NOR2_X1 U843 ( .A1(n1174), .A2(n1179), .ZN(G63) );
NOR3_X1 U844 ( .A1(n1130), .A2(n1180), .A3(n1181), .ZN(n1179) );
AND3_X1 U845 ( .A1(n1182), .A2(G478), .A3(n1178), .ZN(n1181) );
NOR2_X1 U846 ( .A1(n1183), .A2(n1182), .ZN(n1180) );
NOR2_X1 U847 ( .A1(n1117), .A2(n1131), .ZN(n1183) );
NOR2_X1 U848 ( .A1(n1174), .A2(n1184), .ZN(G60) );
XOR2_X1 U849 ( .A(n1185), .B(n1186), .Z(n1184) );
NAND2_X1 U850 ( .A1(n1178), .A2(G475), .ZN(n1185) );
XOR2_X1 U851 ( .A(n1187), .B(n1188), .Z(G6) );
NOR2_X1 U852 ( .A1(KEYINPUT48), .A2(n1173), .ZN(n1188) );
NOR3_X1 U853 ( .A1(n1174), .A2(n1189), .A3(n1190), .ZN(G57) );
NOR2_X1 U854 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NOR2_X1 U855 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
AND2_X1 U856 ( .A1(KEYINPUT13), .A2(n1195), .ZN(n1194) );
NOR3_X1 U857 ( .A1(KEYINPUT13), .A2(n1195), .A3(n1196), .ZN(n1193) );
NOR2_X1 U858 ( .A1(n1197), .A2(n1198), .ZN(n1189) );
INV_X1 U859 ( .A(n1191), .ZN(n1198) );
XNOR2_X1 U860 ( .A(n1199), .B(n1200), .ZN(n1191) );
XOR2_X1 U861 ( .A(n1201), .B(n1202), .Z(n1200) );
XNOR2_X1 U862 ( .A(n1203), .B(n1156), .ZN(n1199) );
XOR2_X1 U863 ( .A(n1204), .B(KEYINPUT34), .Z(n1203) );
NAND2_X1 U864 ( .A1(n1178), .A2(G472), .ZN(n1204) );
NOR2_X1 U865 ( .A1(n1195), .A2(n1196), .ZN(n1197) );
INV_X1 U866 ( .A(KEYINPUT19), .ZN(n1196) );
XNOR2_X1 U867 ( .A(n1205), .B(n1206), .ZN(n1195) );
NAND2_X1 U868 ( .A1(KEYINPUT16), .A2(G101), .ZN(n1205) );
NOR2_X1 U869 ( .A1(n1174), .A2(n1207), .ZN(G54) );
XOR2_X1 U870 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U871 ( .A(n1210), .B(n1211), .Z(n1209) );
XNOR2_X1 U872 ( .A(n1212), .B(n1213), .ZN(n1211) );
NOR2_X1 U873 ( .A1(KEYINPUT60), .A2(n1214), .ZN(n1213) );
XOR2_X1 U874 ( .A(n1215), .B(n1216), .Z(n1208) );
XOR2_X1 U875 ( .A(KEYINPUT22), .B(n1217), .Z(n1216) );
NOR2_X1 U876 ( .A1(KEYINPUT14), .A2(n1218), .ZN(n1217) );
XNOR2_X1 U877 ( .A(n1219), .B(n1220), .ZN(n1218) );
NOR2_X1 U878 ( .A1(G140), .A2(KEYINPUT23), .ZN(n1220) );
XOR2_X1 U879 ( .A(n1221), .B(n1222), .Z(n1215) );
NAND2_X1 U880 ( .A1(n1178), .A2(G469), .ZN(n1221) );
NOR2_X1 U881 ( .A1(n1174), .A2(n1223), .ZN(G51) );
XOR2_X1 U882 ( .A(n1224), .B(n1225), .Z(n1223) );
XNOR2_X1 U883 ( .A(n1226), .B(n1227), .ZN(n1225) );
XOR2_X1 U884 ( .A(n1228), .B(n1229), .Z(n1224) );
XNOR2_X1 U885 ( .A(KEYINPUT8), .B(KEYINPUT27), .ZN(n1229) );
NAND2_X1 U886 ( .A1(n1178), .A2(n1230), .ZN(n1228) );
NOR2_X1 U887 ( .A1(n1231), .A2(n1117), .ZN(n1178) );
NOR2_X1 U888 ( .A1(n1166), .A2(n1144), .ZN(n1117) );
NAND4_X1 U889 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1144) );
NOR4_X1 U890 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235) );
NOR4_X1 U891 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1085), .ZN(n1239) );
NOR2_X1 U892 ( .A1(n1243), .A2(n1244), .ZN(n1241) );
INV_X1 U893 ( .A(KEYINPUT5), .ZN(n1244) );
NOR3_X1 U894 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1243) );
NOR2_X1 U895 ( .A1(KEYINPUT5), .A2(n1248), .ZN(n1240) );
INV_X1 U896 ( .A(n1249), .ZN(n1238) );
NAND2_X1 U897 ( .A1(n1250), .A2(n1251), .ZN(n1234) );
INV_X1 U898 ( .A(KEYINPUT41), .ZN(n1251) );
NAND2_X1 U899 ( .A1(n1248), .A2(n1252), .ZN(n1233) );
NAND2_X1 U900 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NAND3_X1 U901 ( .A1(n1255), .A2(n1085), .A3(KEYINPUT41), .ZN(n1254) );
NAND3_X1 U902 ( .A1(n1256), .A2(n1257), .A3(KEYINPUT6), .ZN(n1253) );
NAND2_X1 U903 ( .A1(n1121), .A2(n1258), .ZN(n1232) );
NAND3_X1 U904 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1258) );
XOR2_X1 U905 ( .A(KEYINPUT32), .B(n1262), .Z(n1261) );
NAND3_X1 U906 ( .A1(n1099), .A2(n1263), .A3(n1264), .ZN(n1260) );
XNOR2_X1 U907 ( .A(KEYINPUT50), .B(n1265), .ZN(n1263) );
OR3_X1 U908 ( .A1(n1266), .A2(KEYINPUT6), .A3(n1267), .ZN(n1259) );
NAND4_X1 U909 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1166) );
NOR4_X1 U910 ( .A1(n1187), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1271) );
INV_X1 U911 ( .A(n1275), .ZN(n1273) );
INV_X1 U912 ( .A(n1076), .ZN(n1272) );
NAND3_X1 U913 ( .A1(n1255), .A2(n1112), .A3(n1276), .ZN(n1076) );
AND3_X1 U914 ( .A1(n1112), .A2(n1277), .A3(n1276), .ZN(n1187) );
NOR2_X1 U915 ( .A1(n1278), .A2(n1279), .ZN(n1270) );
NOR4_X1 U916 ( .A1(n1280), .A2(n1257), .A3(n1245), .A4(n1104), .ZN(n1279) );
INV_X1 U917 ( .A(n1264), .ZN(n1104) );
INV_X1 U918 ( .A(n1281), .ZN(n1278) );
NOR2_X1 U919 ( .A1(n1138), .A2(G952), .ZN(n1174) );
XNOR2_X1 U920 ( .A(G146), .B(n1282), .ZN(G48) );
NAND2_X1 U921 ( .A1(n1262), .A2(n1121), .ZN(n1282) );
AND2_X1 U922 ( .A1(n1283), .A2(n1277), .ZN(n1262) );
XOR2_X1 U923 ( .A(G143), .B(n1284), .Z(G45) );
NOR3_X1 U924 ( .A1(n1267), .A2(n1266), .A3(n1257), .ZN(n1284) );
INV_X1 U925 ( .A(n1256), .ZN(n1266) );
XNOR2_X1 U926 ( .A(G140), .B(n1249), .ZN(G42) );
NAND4_X1 U927 ( .A1(n1277), .A2(n1265), .A3(n1246), .A4(n1285), .ZN(n1249) );
NOR2_X1 U928 ( .A1(n1085), .A2(n1114), .ZN(n1285) );
INV_X1 U929 ( .A(n1099), .ZN(n1114) );
XOR2_X1 U930 ( .A(G137), .B(n1237), .Z(G39) );
AND3_X1 U931 ( .A1(n1123), .A2(n1105), .A3(n1283), .ZN(n1237) );
XOR2_X1 U932 ( .A(n1286), .B(n1250), .Z(G36) );
NOR3_X1 U933 ( .A1(n1085), .A2(n1103), .A3(n1267), .ZN(n1250) );
INV_X1 U934 ( .A(n1248), .ZN(n1267) );
INV_X1 U935 ( .A(n1255), .ZN(n1103) );
XNOR2_X1 U936 ( .A(G134), .B(KEYINPUT7), .ZN(n1286) );
XOR2_X1 U937 ( .A(n1287), .B(G131), .Z(G33) );
NAND2_X1 U938 ( .A1(KEYINPUT15), .A2(n1288), .ZN(n1287) );
NAND3_X1 U939 ( .A1(n1105), .A2(n1277), .A3(n1248), .ZN(n1288) );
NOR3_X1 U940 ( .A1(n1100), .A2(n1247), .A3(n1245), .ZN(n1248) );
INV_X1 U941 ( .A(n1098), .ZN(n1245) );
INV_X1 U942 ( .A(n1085), .ZN(n1105) );
NAND2_X1 U943 ( .A1(n1118), .A2(n1289), .ZN(n1085) );
XNOR2_X1 U944 ( .A(n1290), .B(n1236), .ZN(G30) );
AND3_X1 U945 ( .A1(n1255), .A2(n1121), .A3(n1283), .ZN(n1236) );
NOR4_X1 U946 ( .A1(n1291), .A2(n1100), .A3(n1247), .A4(n1124), .ZN(n1283) );
XNOR2_X1 U947 ( .A(G101), .B(n1281), .ZN(G3) );
NAND3_X1 U948 ( .A1(n1123), .A2(n1276), .A3(n1098), .ZN(n1281) );
XNOR2_X1 U949 ( .A(G125), .B(n1292), .ZN(G27) );
NAND4_X1 U950 ( .A1(n1264), .A2(n1099), .A3(n1293), .A4(n1294), .ZN(n1292) );
XNOR2_X1 U951 ( .A(KEYINPUT35), .B(n1257), .ZN(n1294) );
NOR2_X1 U952 ( .A1(KEYINPUT37), .A2(n1247), .ZN(n1293) );
INV_X1 U953 ( .A(n1265), .ZN(n1247) );
NAND2_X1 U954 ( .A1(n1295), .A2(n1082), .ZN(n1265) );
XOR2_X1 U955 ( .A(n1296), .B(KEYINPUT4), .Z(n1295) );
NAND4_X1 U956 ( .A1(G953), .A2(G902), .A3(n1297), .A4(n1140), .ZN(n1296) );
INV_X1 U957 ( .A(G900), .ZN(n1140) );
XNOR2_X1 U958 ( .A(G122), .B(n1268), .ZN(G24) );
NAND3_X1 U959 ( .A1(n1112), .A2(n1256), .A3(n1298), .ZN(n1268) );
NAND2_X1 U960 ( .A1(n1299), .A2(n1300), .ZN(n1256) );
NAND3_X1 U961 ( .A1(n1128), .A2(n1301), .A3(n1302), .ZN(n1300) );
NAND2_X1 U962 ( .A1(KEYINPUT33), .A2(n1255), .ZN(n1299) );
NOR2_X1 U963 ( .A1(n1303), .A2(n1304), .ZN(n1112) );
NAND3_X1 U964 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(G21) );
NAND2_X1 U965 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND2_X1 U966 ( .A1(n1310), .A2(KEYINPUT52), .ZN(n1308) );
XOR2_X1 U967 ( .A(n1269), .B(KEYINPUT26), .Z(n1310) );
NAND3_X1 U968 ( .A1(KEYINPUT52), .A2(G119), .A3(n1269), .ZN(n1306) );
OR2_X1 U969 ( .A1(n1269), .A2(KEYINPUT52), .ZN(n1305) );
NAND4_X1 U970 ( .A1(n1304), .A2(n1298), .A3(n1123), .A4(n1303), .ZN(n1269) );
XOR2_X1 U971 ( .A(G116), .B(n1274), .Z(G18) );
AND3_X1 U972 ( .A1(n1298), .A2(n1255), .A3(n1098), .ZN(n1274) );
NOR2_X1 U973 ( .A1(n1128), .A2(n1311), .ZN(n1255) );
NOR3_X1 U974 ( .A1(n1096), .A2(n1280), .A3(n1257), .ZN(n1298) );
XNOR2_X1 U975 ( .A(G113), .B(n1312), .ZN(G15) );
NAND4_X1 U976 ( .A1(KEYINPUT21), .A2(n1264), .A3(n1313), .A4(n1098), .ZN(n1312) );
NOR2_X1 U977 ( .A1(n1291), .A2(n1303), .ZN(n1098) );
NOR2_X1 U978 ( .A1(n1280), .A2(n1314), .ZN(n1313) );
XNOR2_X1 U979 ( .A(n1121), .B(KEYINPUT62), .ZN(n1314) );
NOR2_X1 U980 ( .A1(n1242), .A2(n1096), .ZN(n1264) );
AND2_X1 U981 ( .A1(n1315), .A2(n1316), .ZN(n1096) );
OR2_X1 U982 ( .A1(n1100), .A2(KEYINPUT47), .ZN(n1316) );
NAND3_X1 U983 ( .A1(n1111), .A2(n1317), .A3(KEYINPUT47), .ZN(n1315) );
INV_X1 U984 ( .A(n1277), .ZN(n1242) );
NAND2_X1 U985 ( .A1(n1318), .A2(n1319), .ZN(n1277) );
NAND3_X1 U986 ( .A1(n1128), .A2(n1311), .A3(n1302), .ZN(n1319) );
INV_X1 U987 ( .A(KEYINPUT33), .ZN(n1302) );
NAND2_X1 U988 ( .A1(KEYINPUT33), .A2(n1123), .ZN(n1318) );
XNOR2_X1 U989 ( .A(G110), .B(n1275), .ZN(G12) );
NAND3_X1 U990 ( .A1(n1123), .A2(n1276), .A3(n1099), .ZN(n1275) );
NOR2_X1 U991 ( .A1(n1304), .A2(n1124), .ZN(n1099) );
INV_X1 U992 ( .A(n1303), .ZN(n1124) );
NAND3_X1 U993 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1303) );
OR2_X1 U994 ( .A1(n1323), .A2(n1177), .ZN(n1322) );
NAND3_X1 U995 ( .A1(n1177), .A2(n1323), .A3(n1231), .ZN(n1321) );
NAND2_X1 U996 ( .A1(G217), .A2(n1324), .ZN(n1323) );
XOR2_X1 U997 ( .A(n1325), .B(n1326), .Z(n1177) );
XNOR2_X1 U998 ( .A(G137), .B(n1327), .ZN(n1326) );
NAND2_X1 U999 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NAND2_X1 U1000 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
XOR2_X1 U1001 ( .A(n1332), .B(KEYINPUT56), .Z(n1328) );
OR2_X1 U1002 ( .A1(n1331), .A2(n1330), .ZN(n1332) );
XOR2_X1 U1003 ( .A(n1333), .B(n1334), .Z(n1330) );
XNOR2_X1 U1004 ( .A(G128), .B(G110), .ZN(n1333) );
XOR2_X1 U1005 ( .A(n1147), .B(n1335), .Z(n1331) );
NOR2_X1 U1006 ( .A1(KEYINPUT28), .A2(n1336), .ZN(n1335) );
XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(G146), .ZN(n1336) );
XNOR2_X1 U1008 ( .A(G125), .B(n1337), .ZN(n1147) );
NAND2_X1 U1009 ( .A1(n1338), .A2(G221), .ZN(n1325) );
NAND2_X1 U1010 ( .A1(G217), .A2(G902), .ZN(n1320) );
INV_X1 U1011 ( .A(n1291), .ZN(n1304) );
XOR2_X1 U1012 ( .A(n1339), .B(n1132), .Z(n1291) );
NAND2_X1 U1013 ( .A1(n1340), .A2(n1231), .ZN(n1132) );
XOR2_X1 U1014 ( .A(n1341), .B(n1342), .Z(n1340) );
XNOR2_X1 U1015 ( .A(n1343), .B(n1202), .ZN(n1342) );
XOR2_X1 U1016 ( .A(n1344), .B(n1345), .Z(n1202) );
INV_X1 U1017 ( .A(n1346), .ZN(n1345) );
NAND2_X1 U1018 ( .A1(KEYINPUT25), .A2(n1334), .ZN(n1344) );
NAND2_X1 U1019 ( .A1(KEYINPUT45), .A2(n1347), .ZN(n1343) );
INV_X1 U1020 ( .A(G101), .ZN(n1347) );
XOR2_X1 U1021 ( .A(n1348), .B(n1206), .Z(n1341) );
AND3_X1 U1022 ( .A1(n1349), .A2(n1138), .A3(G210), .ZN(n1206) );
NAND2_X1 U1023 ( .A1(n1350), .A2(n1351), .ZN(n1348) );
NAND2_X1 U1024 ( .A1(n1352), .A2(n1212), .ZN(n1351) );
XOR2_X1 U1025 ( .A(n1353), .B(KEYINPUT18), .Z(n1350) );
OR2_X1 U1026 ( .A1(n1352), .A2(n1212), .ZN(n1353) );
XOR2_X1 U1027 ( .A(n1201), .B(KEYINPUT31), .Z(n1352) );
NAND2_X1 U1028 ( .A1(KEYINPUT20), .A2(n1134), .ZN(n1339) );
INV_X1 U1029 ( .A(G472), .ZN(n1134) );
NOR3_X1 U1030 ( .A1(n1100), .A2(n1280), .A3(n1257), .ZN(n1276) );
INV_X1 U1031 ( .A(n1121), .ZN(n1257) );
NOR2_X1 U1032 ( .A1(n1118), .A2(n1119), .ZN(n1121) );
INV_X1 U1033 ( .A(n1289), .ZN(n1119) );
NAND2_X1 U1034 ( .A1(G214), .A2(n1354), .ZN(n1289) );
XOR2_X1 U1035 ( .A(n1355), .B(n1230), .Z(n1118) );
AND2_X1 U1036 ( .A1(G210), .A2(n1354), .ZN(n1230) );
NAND2_X1 U1037 ( .A1(n1349), .A2(n1231), .ZN(n1354) );
NAND2_X1 U1038 ( .A1(n1356), .A2(n1231), .ZN(n1355) );
XOR2_X1 U1039 ( .A(n1226), .B(n1357), .Z(n1356) );
XNOR2_X1 U1040 ( .A(n1358), .B(KEYINPUT11), .ZN(n1357) );
NAND2_X1 U1041 ( .A1(KEYINPUT2), .A2(n1227), .ZN(n1358) );
XOR2_X1 U1042 ( .A(G125), .B(n1201), .Z(n1227) );
XOR2_X1 U1043 ( .A(n1359), .B(n1290), .Z(n1201) );
NAND2_X1 U1044 ( .A1(KEYINPUT40), .A2(n1360), .ZN(n1359) );
XOR2_X1 U1045 ( .A(n1361), .B(n1362), .Z(n1226) );
XNOR2_X1 U1046 ( .A(n1219), .B(n1363), .ZN(n1362) );
NOR2_X1 U1047 ( .A1(G953), .A2(n1160), .ZN(n1363) );
INV_X1 U1048 ( .A(G224), .ZN(n1160) );
INV_X1 U1049 ( .A(G110), .ZN(n1219) );
XOR2_X1 U1050 ( .A(n1172), .B(n1364), .Z(n1361) );
XOR2_X1 U1051 ( .A(n1365), .B(n1366), .Z(n1172) );
XOR2_X1 U1052 ( .A(n1334), .B(n1367), .Z(n1366) );
XNOR2_X1 U1053 ( .A(n1309), .B(KEYINPUT57), .ZN(n1334) );
INV_X1 U1054 ( .A(G119), .ZN(n1309) );
XNOR2_X1 U1055 ( .A(n1346), .B(KEYINPUT30), .ZN(n1365) );
XOR2_X1 U1056 ( .A(G113), .B(n1368), .Z(n1346) );
XOR2_X1 U1057 ( .A(KEYINPUT43), .B(G116), .Z(n1368) );
AND2_X1 U1058 ( .A1(n1082), .A2(n1369), .ZN(n1280) );
NAND4_X1 U1059 ( .A1(G953), .A2(G902), .A3(n1297), .A4(n1161), .ZN(n1369) );
INV_X1 U1060 ( .A(G898), .ZN(n1161) );
NAND3_X1 U1061 ( .A1(n1297), .A2(n1138), .A3(G952), .ZN(n1082) );
NAND2_X1 U1062 ( .A1(G237), .A2(G234), .ZN(n1297) );
INV_X1 U1063 ( .A(n1246), .ZN(n1100) );
NOR2_X1 U1064 ( .A1(n1111), .A2(n1113), .ZN(n1246) );
INV_X1 U1065 ( .A(n1317), .ZN(n1113) );
NAND2_X1 U1066 ( .A1(G221), .A2(n1370), .ZN(n1317) );
NAND2_X1 U1067 ( .A1(G234), .A2(n1231), .ZN(n1370) );
XOR2_X1 U1068 ( .A(n1371), .B(G469), .Z(n1111) );
NAND2_X1 U1069 ( .A1(n1372), .A2(n1231), .ZN(n1371) );
XOR2_X1 U1070 ( .A(n1373), .B(n1374), .Z(n1372) );
XNOR2_X1 U1071 ( .A(n1222), .B(n1156), .ZN(n1374) );
INV_X1 U1072 ( .A(n1212), .ZN(n1156) );
XOR2_X1 U1073 ( .A(G131), .B(n1375), .Z(n1212) );
XOR2_X1 U1074 ( .A(G137), .B(G134), .Z(n1375) );
NOR2_X1 U1075 ( .A1(n1139), .A2(G953), .ZN(n1222) );
INV_X1 U1076 ( .A(G227), .ZN(n1139) );
XOR2_X1 U1077 ( .A(n1376), .B(n1377), .Z(n1373) );
NOR2_X1 U1078 ( .A1(KEYINPUT38), .A2(n1378), .ZN(n1377) );
XNOR2_X1 U1079 ( .A(G140), .B(n1379), .ZN(n1378) );
NOR2_X1 U1080 ( .A1(G110), .A2(KEYINPUT44), .ZN(n1379) );
NAND2_X1 U1081 ( .A1(n1380), .A2(n1381), .ZN(n1376) );
NAND2_X1 U1082 ( .A1(n1214), .A2(n1210), .ZN(n1381) );
XOR2_X1 U1083 ( .A(KEYINPUT3), .B(n1382), .Z(n1380) );
NOR2_X1 U1084 ( .A1(n1214), .A2(n1210), .ZN(n1382) );
XNOR2_X1 U1085 ( .A(n1151), .B(KEYINPUT12), .ZN(n1210) );
XNOR2_X1 U1086 ( .A(n1383), .B(n1360), .ZN(n1151) );
XOR2_X1 U1087 ( .A(G143), .B(G146), .Z(n1360) );
NAND2_X1 U1088 ( .A1(KEYINPUT53), .A2(n1290), .ZN(n1383) );
XNOR2_X1 U1089 ( .A(G104), .B(n1367), .ZN(n1214) );
XNOR2_X1 U1090 ( .A(n1384), .B(G101), .ZN(n1367) );
INV_X1 U1091 ( .A(G107), .ZN(n1384) );
NOR2_X1 U1092 ( .A1(n1301), .A2(n1128), .ZN(n1123) );
XNOR2_X1 U1093 ( .A(n1385), .B(G475), .ZN(n1128) );
NAND2_X1 U1094 ( .A1(n1186), .A2(n1231), .ZN(n1385) );
INV_X1 U1095 ( .A(G902), .ZN(n1231) );
XNOR2_X1 U1096 ( .A(n1386), .B(n1387), .ZN(n1186) );
XNOR2_X1 U1097 ( .A(n1364), .B(n1388), .ZN(n1387) );
XNOR2_X1 U1098 ( .A(n1389), .B(n1390), .ZN(n1388) );
NOR2_X1 U1099 ( .A1(n1391), .A2(KEYINPUT54), .ZN(n1390) );
AND3_X1 U1100 ( .A1(G214), .A2(n1138), .A3(n1349), .ZN(n1391) );
INV_X1 U1101 ( .A(G237), .ZN(n1349) );
INV_X1 U1102 ( .A(G953), .ZN(n1138) );
NOR2_X1 U1103 ( .A1(KEYINPUT36), .A2(n1392), .ZN(n1389) );
XOR2_X1 U1104 ( .A(n1393), .B(n1394), .Z(n1392) );
XOR2_X1 U1105 ( .A(G125), .B(n1395), .Z(n1394) );
NOR2_X1 U1106 ( .A1(KEYINPUT61), .A2(n1396), .ZN(n1395) );
XOR2_X1 U1107 ( .A(KEYINPUT49), .B(G146), .Z(n1396) );
NAND2_X1 U1108 ( .A1(KEYINPUT24), .A2(n1337), .ZN(n1393) );
INV_X1 U1109 ( .A(G140), .ZN(n1337) );
XNOR2_X1 U1110 ( .A(n1173), .B(G122), .ZN(n1364) );
INV_X1 U1111 ( .A(G104), .ZN(n1173) );
XNOR2_X1 U1112 ( .A(G113), .B(n1397), .ZN(n1386) );
XOR2_X1 U1113 ( .A(G143), .B(G131), .Z(n1397) );
INV_X1 U1114 ( .A(n1311), .ZN(n1301) );
XOR2_X1 U1115 ( .A(n1130), .B(n1131), .Z(n1311) );
INV_X1 U1116 ( .A(G478), .ZN(n1131) );
NOR2_X1 U1117 ( .A1(n1182), .A2(G902), .ZN(n1130) );
XNOR2_X1 U1118 ( .A(n1398), .B(n1399), .ZN(n1182) );
XOR2_X1 U1119 ( .A(n1400), .B(n1401), .Z(n1399) );
XNOR2_X1 U1120 ( .A(G107), .B(n1402), .ZN(n1401) );
NOR2_X1 U1121 ( .A1(G143), .A2(KEYINPUT1), .ZN(n1402) );
NAND2_X1 U1122 ( .A1(G217), .A2(n1338), .ZN(n1400) );
NOR2_X1 U1123 ( .A1(n1324), .A2(G953), .ZN(n1338) );
INV_X1 U1124 ( .A(G234), .ZN(n1324) );
XOR2_X1 U1125 ( .A(n1403), .B(n1404), .Z(n1398) );
XNOR2_X1 U1126 ( .A(G134), .B(n1290), .ZN(n1404) );
INV_X1 U1127 ( .A(G128), .ZN(n1290) );
XNOR2_X1 U1128 ( .A(G116), .B(G122), .ZN(n1403) );
endmodule


