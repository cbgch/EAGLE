//Key = 0011101101110110111011101111111101101010111110010101101110101101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341;

XOR2_X1 U731 ( .A(n1016), .B(n1017), .Z(G9) );
XOR2_X1 U732 ( .A(KEYINPUT28), .B(G107), .Z(n1017) );
NOR2_X1 U733 ( .A1(n1018), .A2(n1019), .ZN(G75) );
NOR4_X1 U734 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1019) );
XOR2_X1 U735 ( .A(n1024), .B(KEYINPUT63), .Z(n1023) );
NAND4_X1 U736 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
XOR2_X1 U737 ( .A(KEYINPUT50), .B(n1029), .Z(n1028) );
NOR3_X1 U738 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1022) );
NOR2_X1 U739 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U740 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR3_X1 U741 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1035) );
NOR2_X1 U742 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U743 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U744 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U745 ( .A1(n1046), .A2(n1047), .ZN(n1037) );
AND3_X1 U746 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1033) );
NAND3_X1 U747 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1020) );
NAND3_X1 U748 ( .A1(n1054), .A2(n1055), .A3(n1025), .ZN(n1053) );
NOR3_X1 U749 ( .A1(n1032), .A2(n1041), .A3(n1047), .ZN(n1025) );
INV_X1 U750 ( .A(n1049), .ZN(n1041) );
NAND2_X1 U751 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR3_X1 U752 ( .A1(n1058), .A2(G953), .A3(G952), .ZN(n1018) );
INV_X1 U753 ( .A(n1051), .ZN(n1058) );
NAND4_X1 U754 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1051) );
NOR4_X1 U755 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1062) );
XOR2_X1 U756 ( .A(n1027), .B(KEYINPUT4), .Z(n1064) );
XOR2_X1 U757 ( .A(n1067), .B(KEYINPUT49), .Z(n1063) );
NOR3_X1 U758 ( .A1(n1068), .A2(n1069), .A3(n1029), .ZN(n1061) );
INV_X1 U759 ( .A(n1045), .ZN(n1068) );
NAND2_X1 U760 ( .A1(G478), .A2(n1070), .ZN(n1060) );
XNOR2_X1 U761 ( .A(n1071), .B(n1072), .ZN(n1059) );
NAND2_X1 U762 ( .A1(KEYINPUT40), .A2(n1073), .ZN(n1072) );
NAND2_X1 U763 ( .A1(n1074), .A2(n1075), .ZN(G72) );
NAND2_X1 U764 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U765 ( .A(KEYINPUT24), .B(n1078), .Z(n1074) );
NOR2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1078) );
AND2_X1 U767 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NAND2_X1 U768 ( .A1(n1081), .A2(n1052), .ZN(n1080) );
XOR2_X1 U769 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U770 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NOR2_X1 U771 ( .A1(n1056), .A2(n1086), .ZN(n1084) );
OR3_X1 U772 ( .A1(n1087), .A2(n1083), .A3(n1052), .ZN(n1079) );
XNOR2_X1 U773 ( .A(n1088), .B(n1089), .ZN(n1083) );
XNOR2_X1 U774 ( .A(n1090), .B(n1091), .ZN(n1089) );
NOR2_X1 U775 ( .A1(KEYINPUT5), .A2(n1092), .ZN(n1091) );
XOR2_X1 U776 ( .A(G140), .B(G125), .Z(n1092) );
NAND2_X1 U777 ( .A1(n1093), .A2(KEYINPUT56), .ZN(n1090) );
XOR2_X1 U778 ( .A(n1094), .B(n1095), .Z(n1093) );
XOR2_X1 U779 ( .A(n1096), .B(KEYINPUT48), .Z(n1094) );
NAND2_X1 U780 ( .A1(KEYINPUT42), .A2(G137), .ZN(n1096) );
NOR2_X1 U781 ( .A1(n1097), .A2(n1098), .ZN(n1076) );
AND2_X1 U782 ( .A1(G900), .A2(G227), .ZN(n1098) );
XOR2_X1 U783 ( .A(n1099), .B(n1100), .Z(G69) );
XOR2_X1 U784 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U785 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XOR2_X1 U786 ( .A(KEYINPUT39), .B(G953), .Z(n1104) );
NOR2_X1 U787 ( .A1(n1105), .A2(n1106), .ZN(n1101) );
XOR2_X1 U788 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U789 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND2_X1 U790 ( .A1(KEYINPUT34), .A2(n1111), .ZN(n1109) );
XNOR2_X1 U791 ( .A(n1112), .B(KEYINPUT14), .ZN(n1107) );
NAND2_X1 U792 ( .A1(KEYINPUT52), .A2(n1113), .ZN(n1112) );
NOR2_X1 U793 ( .A1(n1114), .A2(n1097), .ZN(n1099) );
XNOR2_X1 U794 ( .A(n1052), .B(KEYINPUT54), .ZN(n1097) );
AND2_X1 U795 ( .A1(G224), .A2(G898), .ZN(n1114) );
NOR2_X1 U796 ( .A1(n1115), .A2(n1116), .ZN(G66) );
XNOR2_X1 U797 ( .A(n1117), .B(n1118), .ZN(n1116) );
NOR2_X1 U798 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NOR2_X1 U799 ( .A1(n1115), .A2(n1121), .ZN(G63) );
XOR2_X1 U800 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U801 ( .A(KEYINPUT25), .B(n1124), .Z(n1123) );
NOR2_X1 U802 ( .A1(n1125), .A2(n1120), .ZN(n1124) );
INV_X1 U803 ( .A(G478), .ZN(n1125) );
NOR2_X1 U804 ( .A1(n1115), .A2(n1126), .ZN(G60) );
NOR3_X1 U805 ( .A1(n1071), .A2(n1127), .A3(n1128), .ZN(n1126) );
NOR4_X1 U806 ( .A1(n1129), .A2(n1120), .A3(KEYINPUT0), .A4(n1073), .ZN(n1128) );
NOR2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1127) );
NOR3_X1 U808 ( .A1(n1073), .A2(KEYINPUT0), .A3(n1132), .ZN(n1130) );
INV_X1 U809 ( .A(n1021), .ZN(n1132) );
INV_X1 U810 ( .A(G475), .ZN(n1073) );
XOR2_X1 U811 ( .A(G104), .B(n1133), .Z(G6) );
NOR2_X1 U812 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NOR2_X1 U813 ( .A1(n1115), .A2(n1136), .ZN(G57) );
XOR2_X1 U814 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
NAND2_X1 U816 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XOR2_X1 U817 ( .A(n1143), .B(n1144), .Z(n1139) );
NOR2_X1 U818 ( .A1(n1145), .A2(n1120), .ZN(n1144) );
INV_X1 U819 ( .A(G472), .ZN(n1145) );
OR2_X1 U820 ( .A1(n1142), .A2(n1141), .ZN(n1143) );
XNOR2_X1 U821 ( .A(n1146), .B(n1147), .ZN(n1141) );
XOR2_X1 U822 ( .A(n1148), .B(n1149), .Z(n1146) );
NAND2_X1 U823 ( .A1(KEYINPUT7), .A2(n1150), .ZN(n1148) );
INV_X1 U824 ( .A(KEYINPUT13), .ZN(n1142) );
NOR2_X1 U825 ( .A1(n1115), .A2(n1151), .ZN(G54) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U827 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND2_X1 U828 ( .A1(KEYINPUT2), .A2(n1156), .ZN(n1155) );
XNOR2_X1 U829 ( .A(n1157), .B(n1158), .ZN(n1156) );
NAND2_X1 U830 ( .A1(n1159), .A2(KEYINPUT55), .ZN(n1157) );
XOR2_X1 U831 ( .A(n1160), .B(KEYINPUT21), .Z(n1159) );
NAND2_X1 U832 ( .A1(n1161), .A2(n1162), .ZN(n1154) );
NAND2_X1 U833 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
INV_X1 U834 ( .A(n1165), .ZN(n1161) );
NOR2_X1 U835 ( .A1(n1166), .A2(n1120), .ZN(n1152) );
INV_X1 U836 ( .A(G469), .ZN(n1166) );
NOR2_X1 U837 ( .A1(n1115), .A2(n1167), .ZN(G51) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U839 ( .A1(n1170), .A2(n1120), .ZN(n1169) );
NAND2_X1 U840 ( .A1(G902), .A2(n1021), .ZN(n1120) );
NAND3_X1 U841 ( .A1(n1103), .A2(n1171), .A3(n1172), .ZN(n1021) );
XOR2_X1 U842 ( .A(n1173), .B(KEYINPUT8), .Z(n1172) );
NAND2_X1 U843 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
INV_X1 U844 ( .A(n1085), .ZN(n1171) );
NAND4_X1 U845 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1085) );
NOR3_X1 U846 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1179) );
NOR2_X1 U847 ( .A1(n1047), .A2(n1183), .ZN(n1182) );
NOR3_X1 U848 ( .A1(n1184), .A2(n1185), .A3(n1056), .ZN(n1181) );
NOR2_X1 U849 ( .A1(n1186), .A2(n1038), .ZN(n1185) );
NOR2_X1 U850 ( .A1(n1134), .A2(n1187), .ZN(n1186) );
AND4_X1 U851 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1103) );
AND4_X1 U852 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
OR2_X1 U853 ( .A1(n1016), .A2(KEYINPUT15), .ZN(n1190) );
NAND3_X1 U854 ( .A1(n1196), .A2(n1049), .A3(n1197), .ZN(n1016) );
NAND2_X1 U855 ( .A1(n1198), .A2(n1199), .ZN(n1189) );
NAND3_X1 U856 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1199) );
NAND2_X1 U857 ( .A1(n1203), .A2(n1197), .ZN(n1202) );
XOR2_X1 U858 ( .A(KEYINPUT22), .B(n1046), .Z(n1203) );
OR3_X1 U859 ( .A1(n1187), .A2(n1026), .A3(KEYINPUT9), .ZN(n1201) );
NAND2_X1 U860 ( .A1(KEYINPUT9), .A2(n1204), .ZN(n1200) );
NAND2_X1 U861 ( .A1(n1043), .A2(n1205), .ZN(n1188) );
NAND2_X1 U862 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U863 ( .A1(KEYINPUT15), .A2(n1208), .ZN(n1207) );
NAND4_X1 U864 ( .A1(n1197), .A2(n1050), .A3(n1049), .A4(n1209), .ZN(n1208) );
XOR2_X1 U865 ( .A(n1135), .B(KEYINPUT12), .Z(n1206) );
NAND4_X1 U866 ( .A1(n1175), .A2(n1050), .A3(n1049), .A4(n1209), .ZN(n1135) );
NOR2_X1 U867 ( .A1(n1052), .A2(G952), .ZN(n1115) );
XOR2_X1 U868 ( .A(n1210), .B(n1211), .Z(G48) );
NAND4_X1 U869 ( .A1(n1212), .A2(n1175), .A3(n1043), .A4(n1213), .ZN(n1211) );
XOR2_X1 U870 ( .A(KEYINPUT45), .B(n1214), .Z(n1213) );
XOR2_X1 U871 ( .A(n1215), .B(n1178), .Z(G45) );
NAND3_X1 U872 ( .A1(n1212), .A2(n1043), .A3(n1216), .ZN(n1178) );
NOR3_X1 U873 ( .A1(n1046), .A2(n1217), .A3(n1218), .ZN(n1216) );
INV_X1 U874 ( .A(n1219), .ZN(n1046) );
XOR2_X1 U875 ( .A(n1220), .B(n1221), .Z(G42) );
NAND3_X1 U876 ( .A1(n1038), .A2(n1212), .A3(n1222), .ZN(n1221) );
XOR2_X1 U877 ( .A(n1056), .B(KEYINPUT11), .Z(n1222) );
AND2_X1 U878 ( .A1(n1048), .A2(n1223), .ZN(n1038) );
XOR2_X1 U879 ( .A(G137), .B(n1224), .Z(G39) );
NOR2_X1 U880 ( .A1(n1225), .A2(n1047), .ZN(n1224) );
XOR2_X1 U881 ( .A(n1183), .B(KEYINPUT53), .Z(n1225) );
NAND2_X1 U882 ( .A1(n1212), .A2(n1204), .ZN(n1183) );
XOR2_X1 U883 ( .A(G134), .B(n1180), .Z(G36) );
NOR2_X1 U884 ( .A1(n1057), .A2(n1086), .ZN(n1180) );
NAND2_X1 U885 ( .A1(n1226), .A2(n1227), .ZN(G33) );
NAND2_X1 U886 ( .A1(G131), .A2(n1228), .ZN(n1227) );
XOR2_X1 U887 ( .A(KEYINPUT31), .B(n1229), .Z(n1226) );
NOR2_X1 U888 ( .A1(G131), .A2(n1228), .ZN(n1229) );
NAND2_X1 U889 ( .A1(n1174), .A2(n1230), .ZN(n1228) );
XOR2_X1 U890 ( .A(KEYINPUT1), .B(n1175), .Z(n1230) );
INV_X1 U891 ( .A(n1086), .ZN(n1174) );
NAND3_X1 U892 ( .A1(n1212), .A2(n1219), .A3(n1048), .ZN(n1086) );
INV_X1 U893 ( .A(n1047), .ZN(n1048) );
NAND2_X1 U894 ( .A1(n1067), .A2(n1045), .ZN(n1047) );
XNOR2_X1 U895 ( .A(G128), .B(n1176), .ZN(G30) );
NAND4_X1 U896 ( .A1(n1212), .A2(n1214), .A3(n1197), .A4(n1043), .ZN(n1176) );
INV_X1 U897 ( .A(n1184), .ZN(n1212) );
NAND2_X1 U898 ( .A1(n1050), .A2(n1231), .ZN(n1184) );
XOR2_X1 U899 ( .A(n1232), .B(n1195), .Z(G3) );
NAND3_X1 U900 ( .A1(n1196), .A2(n1219), .A3(n1026), .ZN(n1195) );
XOR2_X1 U901 ( .A(n1177), .B(n1233), .Z(G27) );
XOR2_X1 U902 ( .A(KEYINPUT3), .B(G125), .Z(n1233) );
NAND4_X1 U903 ( .A1(n1043), .A2(n1231), .A3(n1223), .A4(n1234), .ZN(n1177) );
NOR2_X1 U904 ( .A1(n1036), .A2(n1056), .ZN(n1234) );
NAND2_X1 U905 ( .A1(n1032), .A2(n1235), .ZN(n1231) );
NAND4_X1 U906 ( .A1(G902), .A2(G953), .A3(n1236), .A4(n1087), .ZN(n1235) );
INV_X1 U907 ( .A(G900), .ZN(n1087) );
XOR2_X1 U908 ( .A(n1194), .B(n1237), .Z(G24) );
NAND2_X1 U909 ( .A1(KEYINPUT6), .A2(G122), .ZN(n1237) );
NAND4_X1 U910 ( .A1(n1198), .A2(n1049), .A3(n1238), .A4(n1239), .ZN(n1194) );
NAND2_X1 U911 ( .A1(n1240), .A2(n1241), .ZN(n1049) );
OR3_X1 U912 ( .A1(n1066), .A2(n1065), .A3(KEYINPUT59), .ZN(n1241) );
NAND2_X1 U913 ( .A1(KEYINPUT59), .A2(n1223), .ZN(n1240) );
XOR2_X1 U914 ( .A(n1242), .B(n1243), .Z(G21) );
NAND2_X1 U915 ( .A1(n1204), .A2(n1198), .ZN(n1243) );
NOR2_X1 U916 ( .A1(n1187), .A2(n1030), .ZN(n1204) );
NAND2_X1 U917 ( .A1(KEYINPUT47), .A2(G119), .ZN(n1242) );
XNOR2_X1 U918 ( .A(G116), .B(n1244), .ZN(G18) );
NAND2_X1 U919 ( .A1(n1245), .A2(n1197), .ZN(n1244) );
INV_X1 U920 ( .A(n1057), .ZN(n1197) );
NAND2_X1 U921 ( .A1(n1218), .A2(n1239), .ZN(n1057) );
XNOR2_X1 U922 ( .A(G113), .B(n1193), .ZN(G15) );
NAND2_X1 U923 ( .A1(n1175), .A2(n1245), .ZN(n1193) );
AND2_X1 U924 ( .A1(n1198), .A2(n1219), .ZN(n1245) );
NAND2_X1 U925 ( .A1(n1246), .A2(n1247), .ZN(n1219) );
NAND3_X1 U926 ( .A1(n1066), .A2(n1248), .A3(n1249), .ZN(n1247) );
INV_X1 U927 ( .A(KEYINPUT59), .ZN(n1249) );
NAND2_X1 U928 ( .A1(KEYINPUT59), .A2(n1214), .ZN(n1246) );
INV_X1 U929 ( .A(n1187), .ZN(n1214) );
NAND2_X1 U930 ( .A1(n1065), .A2(n1066), .ZN(n1187) );
INV_X1 U931 ( .A(n1248), .ZN(n1065) );
AND3_X1 U932 ( .A1(n1043), .A2(n1209), .A3(n1054), .ZN(n1198) );
INV_X1 U933 ( .A(n1036), .ZN(n1054) );
NAND2_X1 U934 ( .A1(n1027), .A2(n1250), .ZN(n1036) );
INV_X1 U935 ( .A(n1056), .ZN(n1175) );
NAND2_X1 U936 ( .A1(n1217), .A2(n1238), .ZN(n1056) );
XNOR2_X1 U937 ( .A(G110), .B(n1192), .ZN(G12) );
NAND3_X1 U938 ( .A1(n1196), .A2(n1223), .A3(n1026), .ZN(n1192) );
INV_X1 U939 ( .A(n1030), .ZN(n1026) );
NAND2_X1 U940 ( .A1(n1217), .A2(n1218), .ZN(n1030) );
INV_X1 U941 ( .A(n1238), .ZN(n1218) );
XOR2_X1 U942 ( .A(n1071), .B(G475), .Z(n1238) );
NOR2_X1 U943 ( .A1(n1131), .A2(G902), .ZN(n1071) );
INV_X1 U944 ( .A(n1129), .ZN(n1131) );
XOR2_X1 U945 ( .A(n1251), .B(n1252), .Z(n1129) );
XOR2_X1 U946 ( .A(G104), .B(n1253), .Z(n1252) );
NOR2_X1 U947 ( .A1(KEYINPUT46), .A2(n1254), .ZN(n1253) );
XOR2_X1 U948 ( .A(n1255), .B(n1256), .Z(n1254) );
XOR2_X1 U949 ( .A(n1257), .B(n1258), .Z(n1256) );
AND2_X1 U950 ( .A1(n1259), .A2(G214), .ZN(n1258) );
XOR2_X1 U951 ( .A(G131), .B(n1215), .Z(n1255) );
XNOR2_X1 U952 ( .A(G113), .B(G122), .ZN(n1251) );
INV_X1 U953 ( .A(n1239), .ZN(n1217) );
NAND3_X1 U954 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1239) );
INV_X1 U955 ( .A(n1069), .ZN(n1262) );
NOR2_X1 U956 ( .A1(n1070), .A2(G478), .ZN(n1069) );
OR2_X1 U957 ( .A1(G478), .A2(KEYINPUT61), .ZN(n1261) );
NAND3_X1 U958 ( .A1(G478), .A2(n1070), .A3(KEYINPUT61), .ZN(n1260) );
NAND2_X1 U959 ( .A1(n1122), .A2(n1263), .ZN(n1070) );
XOR2_X1 U960 ( .A(n1264), .B(n1265), .Z(n1122) );
XOR2_X1 U961 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U962 ( .A(G134), .B(G128), .Z(n1267) );
XOR2_X1 U963 ( .A(KEYINPUT20), .B(G143), .Z(n1266) );
XOR2_X1 U964 ( .A(n1268), .B(n1269), .Z(n1264) );
XOR2_X1 U965 ( .A(G122), .B(G116), .Z(n1269) );
XOR2_X1 U966 ( .A(n1270), .B(G107), .Z(n1268) );
NAND2_X1 U967 ( .A1(G217), .A2(n1271), .ZN(n1270) );
INV_X1 U968 ( .A(n1272), .ZN(n1271) );
NOR2_X1 U969 ( .A1(n1066), .A2(n1248), .ZN(n1223) );
XNOR2_X1 U970 ( .A(n1273), .B(n1119), .ZN(n1248) );
NAND2_X1 U971 ( .A1(G217), .A2(n1274), .ZN(n1119) );
NAND2_X1 U972 ( .A1(n1117), .A2(n1263), .ZN(n1273) );
XNOR2_X1 U973 ( .A(n1275), .B(n1276), .ZN(n1117) );
NOR2_X1 U974 ( .A1(n1277), .A2(n1272), .ZN(n1276) );
NAND2_X1 U975 ( .A1(G234), .A2(n1052), .ZN(n1272) );
XNOR2_X1 U976 ( .A(G221), .B(KEYINPUT37), .ZN(n1277) );
XOR2_X1 U977 ( .A(n1278), .B(G137), .Z(n1275) );
NAND3_X1 U978 ( .A1(n1279), .A2(n1280), .A3(KEYINPUT33), .ZN(n1278) );
NAND2_X1 U979 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
INV_X1 U980 ( .A(KEYINPUT32), .ZN(n1282) );
XOR2_X1 U981 ( .A(n1283), .B(n1284), .Z(n1281) );
NAND2_X1 U982 ( .A1(KEYINPUT16), .A2(n1285), .ZN(n1283) );
INV_X1 U983 ( .A(n1257), .ZN(n1285) );
NAND3_X1 U984 ( .A1(n1284), .A2(n1257), .A3(KEYINPUT32), .ZN(n1279) );
XOR2_X1 U985 ( .A(n1220), .B(n1286), .Z(n1257) );
XOR2_X1 U986 ( .A(n1287), .B(n1288), .Z(n1284) );
XOR2_X1 U987 ( .A(G119), .B(n1289), .Z(n1288) );
NOR2_X1 U988 ( .A1(G128), .A2(KEYINPUT35), .ZN(n1289) );
NAND2_X1 U989 ( .A1(KEYINPUT36), .A2(G110), .ZN(n1287) );
XNOR2_X1 U990 ( .A(n1290), .B(G472), .ZN(n1066) );
NAND2_X1 U991 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XOR2_X1 U992 ( .A(KEYINPUT26), .B(G902), .Z(n1292) );
XOR2_X1 U993 ( .A(n1138), .B(n1293), .Z(n1291) );
XNOR2_X1 U994 ( .A(n1294), .B(n1149), .ZN(n1293) );
XOR2_X1 U995 ( .A(G113), .B(n1295), .Z(n1149) );
NOR2_X1 U996 ( .A1(KEYINPUT57), .A2(n1296), .ZN(n1295) );
NAND2_X1 U997 ( .A1(n1297), .A2(KEYINPUT51), .ZN(n1294) );
XOR2_X1 U998 ( .A(n1147), .B(n1150), .Z(n1297) );
XOR2_X1 U999 ( .A(n1210), .B(n1298), .Z(n1150) );
AND2_X1 U1000 ( .A1(n1299), .A2(n1300), .ZN(n1138) );
NAND2_X1 U1001 ( .A1(n1301), .A2(n1232), .ZN(n1300) );
NAND2_X1 U1002 ( .A1(G210), .A2(n1259), .ZN(n1301) );
NAND3_X1 U1003 ( .A1(G210), .A2(n1259), .A3(G101), .ZN(n1299) );
AND2_X1 U1004 ( .A1(n1302), .A2(n1052), .ZN(n1259) );
XOR2_X1 U1005 ( .A(n1303), .B(KEYINPUT23), .Z(n1302) );
AND3_X1 U1006 ( .A1(n1043), .A2(n1209), .A3(n1050), .ZN(n1196) );
NOR2_X1 U1007 ( .A1(n1027), .A2(n1029), .ZN(n1050) );
INV_X1 U1008 ( .A(n1250), .ZN(n1029) );
NAND2_X1 U1009 ( .A1(G221), .A2(n1274), .ZN(n1250) );
NAND2_X1 U1010 ( .A1(G234), .A2(n1263), .ZN(n1274) );
XOR2_X1 U1011 ( .A(n1304), .B(G469), .Z(n1027) );
NAND2_X1 U1012 ( .A1(n1305), .A2(n1263), .ZN(n1304) );
XOR2_X1 U1013 ( .A(n1306), .B(n1307), .Z(n1305) );
NOR3_X1 U1014 ( .A1(n1165), .A2(n1308), .A3(n1309), .ZN(n1307) );
AND3_X1 U1015 ( .A1(KEYINPUT38), .A2(n1164), .A3(n1163), .ZN(n1309) );
NOR2_X1 U1016 ( .A1(KEYINPUT38), .A2(n1164), .ZN(n1308) );
NOR2_X1 U1017 ( .A1(n1164), .A2(n1163), .ZN(n1165) );
AND2_X1 U1018 ( .A1(G227), .A2(n1052), .ZN(n1163) );
XOR2_X1 U1019 ( .A(G110), .B(n1220), .Z(n1164) );
INV_X1 U1020 ( .A(G140), .ZN(n1220) );
NAND2_X1 U1021 ( .A1(KEYINPUT17), .A2(n1310), .ZN(n1306) );
XOR2_X1 U1022 ( .A(n1311), .B(n1147), .Z(n1310) );
INV_X1 U1023 ( .A(n1160), .ZN(n1147) );
XNOR2_X1 U1024 ( .A(G137), .B(n1095), .ZN(n1160) );
XOR2_X1 U1025 ( .A(G134), .B(G131), .Z(n1095) );
NAND2_X1 U1026 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NAND3_X1 U1027 ( .A1(n1314), .A2(n1088), .A3(n1315), .ZN(n1313) );
INV_X1 U1028 ( .A(KEYINPUT10), .ZN(n1315) );
NAND2_X1 U1029 ( .A1(n1158), .A2(KEYINPUT10), .ZN(n1312) );
XOR2_X1 U1030 ( .A(n1088), .B(n1314), .Z(n1158) );
XOR2_X1 U1031 ( .A(n1110), .B(KEYINPUT60), .Z(n1314) );
XOR2_X1 U1032 ( .A(n1316), .B(G128), .Z(n1088) );
NAND2_X1 U1033 ( .A1(n1317), .A2(KEYINPUT41), .ZN(n1316) );
XOR2_X1 U1034 ( .A(n1318), .B(G143), .Z(n1317) );
NAND2_X1 U1035 ( .A1(KEYINPUT18), .A2(n1210), .ZN(n1318) );
INV_X1 U1036 ( .A(G146), .ZN(n1210) );
NAND2_X1 U1037 ( .A1(n1319), .A2(n1320), .ZN(n1209) );
NAND3_X1 U1038 ( .A1(n1105), .A2(n1236), .A3(G902), .ZN(n1320) );
NOR2_X1 U1039 ( .A1(n1052), .A2(G898), .ZN(n1105) );
XNOR2_X1 U1040 ( .A(KEYINPUT43), .B(n1032), .ZN(n1319) );
NAND3_X1 U1041 ( .A1(n1236), .A2(n1052), .A3(G952), .ZN(n1032) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1236) );
INV_X1 U1043 ( .A(n1134), .ZN(n1043) );
NAND2_X1 U1044 ( .A1(n1044), .A2(n1045), .ZN(n1134) );
NAND2_X1 U1045 ( .A1(G214), .A2(n1321), .ZN(n1045) );
INV_X1 U1046 ( .A(n1067), .ZN(n1044) );
XNOR2_X1 U1047 ( .A(n1322), .B(n1170), .ZN(n1067) );
NAND2_X1 U1048 ( .A1(G210), .A2(n1321), .ZN(n1170) );
NAND2_X1 U1049 ( .A1(n1303), .A2(n1263), .ZN(n1321) );
INV_X1 U1050 ( .A(G237), .ZN(n1303) );
NAND2_X1 U1051 ( .A1(n1323), .A2(n1263), .ZN(n1322) );
INV_X1 U1052 ( .A(G902), .ZN(n1263) );
XOR2_X1 U1053 ( .A(n1168), .B(KEYINPUT44), .Z(n1323) );
XOR2_X1 U1054 ( .A(n1324), .B(n1325), .Z(n1168) );
XOR2_X1 U1055 ( .A(n1286), .B(n1298), .Z(n1325) );
XNOR2_X1 U1056 ( .A(n1215), .B(n1326), .ZN(n1298) );
NOR2_X1 U1057 ( .A1(G128), .A2(KEYINPUT19), .ZN(n1326) );
INV_X1 U1058 ( .A(G143), .ZN(n1215) );
XOR2_X1 U1059 ( .A(G125), .B(G146), .Z(n1286) );
XOR2_X1 U1060 ( .A(n1327), .B(n1328), .Z(n1324) );
AND2_X1 U1061 ( .A1(n1052), .A2(G224), .ZN(n1328) );
INV_X1 U1062 ( .A(G953), .ZN(n1052) );
NAND2_X1 U1063 ( .A1(n1329), .A2(n1330), .ZN(n1327) );
NAND2_X1 U1064 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U1065 ( .A(n1111), .B(KEYINPUT27), .Z(n1332) );
XOR2_X1 U1066 ( .A(n1333), .B(KEYINPUT62), .Z(n1331) );
XOR2_X1 U1067 ( .A(KEYINPUT30), .B(n1334), .Z(n1329) );
NOR2_X1 U1068 ( .A1(n1335), .A2(n1333), .ZN(n1334) );
NAND2_X1 U1069 ( .A1(n1336), .A2(n1337), .ZN(n1333) );
NAND2_X1 U1070 ( .A1(n1110), .A2(n1338), .ZN(n1337) );
XOR2_X1 U1071 ( .A(KEYINPUT58), .B(n1339), .Z(n1336) );
NOR2_X1 U1072 ( .A1(n1110), .A2(n1338), .ZN(n1339) );
INV_X1 U1073 ( .A(n1113), .ZN(n1338) );
XOR2_X1 U1074 ( .A(G113), .B(n1296), .Z(n1113) );
XNOR2_X1 U1075 ( .A(G116), .B(G119), .ZN(n1296) );
XOR2_X1 U1076 ( .A(n1340), .B(n1341), .Z(n1110) );
XOR2_X1 U1077 ( .A(KEYINPUT29), .B(G107), .Z(n1341) );
XOR2_X1 U1078 ( .A(G104), .B(n1232), .Z(n1340) );
INV_X1 U1079 ( .A(G101), .ZN(n1232) );
INV_X1 U1080 ( .A(n1111), .ZN(n1335) );
XNOR2_X1 U1081 ( .A(G110), .B(G122), .ZN(n1111) );
endmodule


