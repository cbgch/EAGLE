//Key = 0010110010010111111110010110010101110101100110010110110101100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330;

XOR2_X1 U736 ( .A(n1016), .B(n1017), .Z(G9) );
NAND2_X1 U737 ( .A1(KEYINPUT15), .A2(G107), .ZN(n1017) );
NAND2_X1 U738 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
XNOR2_X1 U739 ( .A(KEYINPUT54), .B(n1020), .ZN(n1019) );
NAND2_X1 U740 ( .A1(n1021), .A2(n1022), .ZN(G75) );
NAND2_X1 U741 ( .A1(G952), .A2(n1023), .ZN(n1022) );
NAND4_X1 U742 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1023) );
XNOR2_X1 U743 ( .A(KEYINPUT49), .B(n1028), .ZN(n1027) );
NOR2_X1 U744 ( .A1(n1029), .A2(n1030), .ZN(n1026) );
INV_X1 U745 ( .A(n1031), .ZN(n1030) );
NOR2_X1 U746 ( .A1(n1032), .A2(n1033), .ZN(n1029) );
NOR2_X1 U747 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR3_X1 U748 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NOR2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U750 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR2_X1 U752 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U753 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U754 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1043) );
NOR2_X1 U756 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR3_X1 U757 ( .A1(n1052), .A2(n1055), .A3(n1046), .ZN(n1039) );
NOR4_X1 U758 ( .A1(n1056), .A2(n1042), .A3(n1046), .A4(n1052), .ZN(n1034) );
NOR2_X1 U759 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U760 ( .A1(n1055), .A2(n1036), .ZN(n1057) );
NOR3_X1 U761 ( .A1(n1059), .A2(n1060), .A3(n1037), .ZN(n1055) );
XOR2_X1 U762 ( .A(KEYINPUT28), .B(n1061), .Z(n1025) );
NAND2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1021) );
INV_X1 U764 ( .A(G952), .ZN(n1063) );
NAND2_X1 U765 ( .A1(n1031), .A2(n1028), .ZN(n1062) );
NAND4_X1 U766 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1028) );
NOR4_X1 U767 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1067) );
XNOR2_X1 U768 ( .A(KEYINPUT62), .B(n1072), .ZN(n1071) );
XNOR2_X1 U769 ( .A(KEYINPUT30), .B(n1073), .ZN(n1070) );
XNOR2_X1 U770 ( .A(n1074), .B(KEYINPUT23), .ZN(n1068) );
AND3_X1 U771 ( .A1(n1075), .A2(n1076), .A3(n1050), .ZN(n1066) );
XOR2_X1 U772 ( .A(n1077), .B(n1078), .Z(n1064) );
NOR2_X1 U773 ( .A1(KEYINPUT7), .A2(n1079), .ZN(n1077) );
XOR2_X1 U774 ( .A(n1080), .B(n1081), .Z(G72) );
NAND2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U776 ( .A1(G900), .A2(G227), .ZN(n1083) );
NAND2_X1 U777 ( .A1(KEYINPUT52), .A2(n1084), .ZN(n1080) );
XOR2_X1 U778 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U779 ( .A1(n1024), .A2(G953), .ZN(n1086) );
NOR2_X1 U780 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
XOR2_X1 U781 ( .A(n1089), .B(n1090), .Z(n1088) );
XOR2_X1 U782 ( .A(n1091), .B(n1092), .Z(n1090) );
XOR2_X1 U783 ( .A(n1093), .B(n1094), .Z(n1089) );
NOR2_X1 U784 ( .A1(KEYINPUT6), .A2(n1095), .ZN(n1094) );
XNOR2_X1 U785 ( .A(G125), .B(KEYINPUT29), .ZN(n1093) );
NOR2_X1 U786 ( .A1(G900), .A2(n1096), .ZN(n1087) );
NAND2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(G69) );
NAND2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U789 ( .A(KEYINPUT13), .B(n1101), .Z(n1097) );
NOR2_X1 U790 ( .A1(n1099), .A2(n1100), .ZN(n1101) );
NAND2_X1 U791 ( .A1(n1082), .A2(n1102), .ZN(n1100) );
NAND2_X1 U792 ( .A1(G898), .A2(G224), .ZN(n1102) );
XNOR2_X1 U793 ( .A(n1096), .B(KEYINPUT59), .ZN(n1082) );
XNOR2_X1 U794 ( .A(n1103), .B(n1104), .ZN(n1099) );
NOR3_X1 U795 ( .A1(n1061), .A2(KEYINPUT9), .A3(G953), .ZN(n1104) );
NAND2_X1 U796 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
XOR2_X1 U797 ( .A(KEYINPUT25), .B(n1107), .Z(n1106) );
NOR2_X1 U798 ( .A1(G898), .A2(n1108), .ZN(n1107) );
XNOR2_X1 U799 ( .A(KEYINPUT43), .B(n1096), .ZN(n1108) );
XNOR2_X1 U800 ( .A(n1109), .B(n1110), .ZN(n1105) );
NOR2_X1 U801 ( .A1(n1111), .A2(n1112), .ZN(G66) );
XNOR2_X1 U802 ( .A(n1113), .B(n1114), .ZN(n1112) );
NOR2_X1 U803 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NOR2_X1 U804 ( .A1(n1111), .A2(n1117), .ZN(G63) );
XNOR2_X1 U805 ( .A(n1118), .B(n1119), .ZN(n1117) );
AND2_X1 U806 ( .A1(G478), .A2(n1120), .ZN(n1119) );
NOR2_X1 U807 ( .A1(n1111), .A2(n1121), .ZN(G60) );
XOR2_X1 U808 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U809 ( .A(KEYINPUT40), .B(n1124), .Z(n1123) );
AND2_X1 U810 ( .A1(G475), .A2(n1120), .ZN(n1124) );
XNOR2_X1 U811 ( .A(n1125), .B(n1126), .ZN(G6) );
NAND2_X1 U812 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
OR3_X1 U813 ( .A1(n1129), .A2(n1054), .A3(KEYINPUT11), .ZN(n1128) );
NAND2_X1 U814 ( .A1(n1130), .A2(KEYINPUT11), .ZN(n1127) );
NOR2_X1 U815 ( .A1(n1111), .A2(n1131), .ZN(G57) );
XOR2_X1 U816 ( .A(n1132), .B(n1133), .Z(n1131) );
XNOR2_X1 U817 ( .A(n1134), .B(n1135), .ZN(n1133) );
NOR2_X1 U818 ( .A1(KEYINPUT32), .A2(n1136), .ZN(n1135) );
XOR2_X1 U819 ( .A(n1137), .B(n1138), .Z(n1136) );
XNOR2_X1 U820 ( .A(n1139), .B(n1140), .ZN(n1138) );
XNOR2_X1 U821 ( .A(n1141), .B(n1142), .ZN(n1137) );
NOR2_X1 U822 ( .A1(n1143), .A2(n1116), .ZN(n1141) );
NOR3_X1 U823 ( .A1(n1111), .A2(n1144), .A3(n1145), .ZN(G54) );
NOR2_X1 U824 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U825 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U826 ( .A1(KEYINPUT0), .A2(n1150), .ZN(n1149) );
NOR2_X1 U827 ( .A1(n1151), .A2(n1152), .ZN(n1144) );
XOR2_X1 U828 ( .A(n1148), .B(n1153), .Z(n1152) );
NOR2_X1 U829 ( .A1(KEYINPUT0), .A2(n1154), .ZN(n1153) );
INV_X1 U830 ( .A(n1150), .ZN(n1154) );
XNOR2_X1 U831 ( .A(n1155), .B(G110), .ZN(n1150) );
NAND2_X1 U832 ( .A1(KEYINPUT17), .A2(n1095), .ZN(n1155) );
XOR2_X1 U833 ( .A(n1156), .B(n1139), .Z(n1148) );
XOR2_X1 U834 ( .A(n1157), .B(n1158), .Z(n1156) );
AND2_X1 U835 ( .A1(G469), .A2(n1120), .ZN(n1158) );
NAND2_X1 U836 ( .A1(KEYINPUT19), .A2(n1159), .ZN(n1157) );
XOR2_X1 U837 ( .A(n1160), .B(n1161), .Z(n1159) );
XNOR2_X1 U838 ( .A(G101), .B(KEYINPUT61), .ZN(n1161) );
INV_X1 U839 ( .A(n1146), .ZN(n1151) );
NOR2_X1 U840 ( .A1(n1111), .A2(n1162), .ZN(G51) );
NOR2_X1 U841 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U842 ( .A(KEYINPUT51), .B(n1165), .Z(n1164) );
NOR2_X1 U843 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
AND2_X1 U844 ( .A1(n1167), .A2(n1166), .ZN(n1163) );
XOR2_X1 U845 ( .A(n1168), .B(n1169), .Z(n1166) );
XOR2_X1 U846 ( .A(n1142), .B(n1170), .Z(n1169) );
XNOR2_X1 U847 ( .A(G125), .B(n1171), .ZN(n1168) );
NAND2_X1 U848 ( .A1(n1120), .A2(n1172), .ZN(n1167) );
INV_X1 U849 ( .A(n1116), .ZN(n1120) );
NAND2_X1 U850 ( .A1(G902), .A2(n1173), .ZN(n1116) );
NAND2_X1 U851 ( .A1(n1024), .A2(n1061), .ZN(n1173) );
AND2_X1 U852 ( .A1(n1174), .A2(n1175), .ZN(n1061) );
NOR4_X1 U853 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1175) );
NOR4_X1 U854 ( .A1(n1180), .A2(n1130), .A3(n1181), .A4(n1182), .ZN(n1174) );
NOR2_X1 U855 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XNOR2_X1 U856 ( .A(KEYINPUT18), .B(n1052), .ZN(n1184) );
INV_X1 U857 ( .A(n1185), .ZN(n1183) );
NOR2_X1 U858 ( .A1(n1020), .A2(n1129), .ZN(n1181) );
NOR2_X1 U859 ( .A1(n1186), .A2(n1129), .ZN(n1130) );
INV_X1 U860 ( .A(n1018), .ZN(n1129) );
NOR3_X1 U861 ( .A1(n1187), .A2(n1042), .A3(n1188), .ZN(n1018) );
AND4_X1 U862 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1024) );
AND4_X1 U863 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
NOR3_X1 U864 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1191) );
NOR2_X1 U865 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
INV_X1 U866 ( .A(KEYINPUT5), .ZN(n1200) );
NOR4_X1 U867 ( .A1(KEYINPUT5), .A2(n1202), .A3(n1048), .A4(n1186), .ZN(n1198) );
NOR2_X1 U868 ( .A1(n1096), .A2(G952), .ZN(n1111) );
XNOR2_X1 U869 ( .A(G146), .B(n1201), .ZN(G48) );
NAND2_X1 U870 ( .A1(n1203), .A2(n1054), .ZN(n1201) );
XOR2_X1 U871 ( .A(n1204), .B(G143), .Z(G45) );
NAND2_X1 U872 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
OR2_X1 U873 ( .A1(n1189), .A2(KEYINPUT56), .ZN(n1206) );
NAND2_X1 U874 ( .A1(n1207), .A2(n1048), .ZN(n1189) );
NAND3_X1 U875 ( .A1(n1207), .A2(n1187), .A3(KEYINPUT56), .ZN(n1205) );
AND4_X1 U876 ( .A1(n1059), .A2(n1208), .A3(n1074), .A4(n1209), .ZN(n1207) );
XOR2_X1 U877 ( .A(n1194), .B(n1210), .Z(G42) );
NAND2_X1 U878 ( .A1(KEYINPUT16), .A2(G140), .ZN(n1210) );
NAND3_X1 U879 ( .A1(n1054), .A2(n1211), .A3(n1060), .ZN(n1194) );
XNOR2_X1 U880 ( .A(G137), .B(n1193), .ZN(G39) );
NAND4_X1 U881 ( .A1(n1212), .A2(n1211), .A3(n1069), .A4(n1213), .ZN(n1193) );
XNOR2_X1 U882 ( .A(G134), .B(n1190), .ZN(G36) );
NAND3_X1 U883 ( .A1(n1211), .A2(n1053), .A3(n1059), .ZN(n1190) );
XNOR2_X1 U884 ( .A(G131), .B(n1196), .ZN(G33) );
NAND3_X1 U885 ( .A1(n1054), .A2(n1211), .A3(n1059), .ZN(n1196) );
INV_X1 U886 ( .A(n1214), .ZN(n1059) );
AND4_X1 U887 ( .A1(n1073), .A2(n1048), .A3(n1215), .A4(n1075), .ZN(n1211) );
INV_X1 U888 ( .A(n1187), .ZN(n1048) );
XNOR2_X1 U889 ( .A(n1216), .B(n1217), .ZN(G30) );
NAND2_X1 U890 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
NAND2_X1 U891 ( .A1(n1197), .A2(n1220), .ZN(n1219) );
INV_X1 U892 ( .A(KEYINPUT63), .ZN(n1220) );
AND2_X1 U893 ( .A1(n1203), .A2(n1053), .ZN(n1197) );
NAND3_X1 U894 ( .A1(n1203), .A2(n1020), .A3(KEYINPUT63), .ZN(n1218) );
NOR2_X1 U895 ( .A1(n1202), .A2(n1187), .ZN(n1203) );
NAND3_X1 U896 ( .A1(n1069), .A2(n1213), .A3(n1208), .ZN(n1202) );
XNOR2_X1 U897 ( .A(n1134), .B(n1177), .ZN(G3) );
NOR4_X1 U898 ( .A1(n1214), .A2(n1046), .A3(n1188), .A4(n1187), .ZN(n1177) );
XNOR2_X1 U899 ( .A(G125), .B(n1195), .ZN(G27) );
NAND4_X1 U900 ( .A1(n1221), .A2(n1208), .A3(n1060), .A4(n1054), .ZN(n1195) );
INV_X1 U901 ( .A(n1222), .ZN(n1060) );
AND2_X1 U902 ( .A1(n1058), .A2(n1215), .ZN(n1208) );
NAND2_X1 U903 ( .A1(n1033), .A2(n1223), .ZN(n1215) );
NAND4_X1 U904 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1225), .ZN(n1223) );
INV_X1 U905 ( .A(G900), .ZN(n1225) );
XNOR2_X1 U906 ( .A(n1180), .B(n1226), .ZN(G24) );
XOR2_X1 U907 ( .A(KEYINPUT31), .B(G122), .Z(n1226) );
NOR4_X1 U908 ( .A1(n1227), .A2(n1072), .A3(n1042), .A4(n1228), .ZN(n1180) );
OR2_X1 U909 ( .A1(n1188), .A2(n1052), .ZN(n1228) );
NAND2_X1 U910 ( .A1(n1229), .A2(n1230), .ZN(n1042) );
NAND2_X1 U911 ( .A1(n1231), .A2(n1232), .ZN(G21) );
OR2_X1 U912 ( .A1(n1233), .A2(n1179), .ZN(n1232) );
XOR2_X1 U913 ( .A(n1234), .B(KEYINPUT48), .Z(n1231) );
NAND2_X1 U914 ( .A1(n1179), .A2(n1233), .ZN(n1234) );
INV_X1 U915 ( .A(G119), .ZN(n1233) );
NOR4_X1 U916 ( .A1(n1052), .A2(n1046), .A3(n1235), .A4(n1188), .ZN(n1179) );
NAND2_X1 U917 ( .A1(n1213), .A2(n1069), .ZN(n1235) );
XNOR2_X1 U918 ( .A(G116), .B(n1236), .ZN(G18) );
NAND2_X1 U919 ( .A1(n1185), .A2(n1221), .ZN(n1236) );
INV_X1 U920 ( .A(n1052), .ZN(n1221) );
NOR3_X1 U921 ( .A1(n1020), .A2(n1188), .A3(n1214), .ZN(n1185) );
INV_X1 U922 ( .A(n1053), .ZN(n1020) );
NOR2_X1 U923 ( .A1(n1209), .A2(n1227), .ZN(n1053) );
INV_X1 U924 ( .A(n1074), .ZN(n1227) );
XNOR2_X1 U925 ( .A(n1237), .B(n1176), .ZN(G15) );
NOR4_X1 U926 ( .A1(n1214), .A2(n1052), .A3(n1186), .A4(n1188), .ZN(n1176) );
INV_X1 U927 ( .A(n1054), .ZN(n1186) );
NOR2_X1 U928 ( .A1(n1074), .A2(n1072), .ZN(n1054) );
INV_X1 U929 ( .A(n1209), .ZN(n1072) );
NAND2_X1 U930 ( .A1(n1238), .A2(n1050), .ZN(n1052) );
NAND2_X1 U931 ( .A1(n1229), .A2(n1213), .ZN(n1214) );
XNOR2_X1 U932 ( .A(n1069), .B(KEYINPUT1), .ZN(n1229) );
XOR2_X1 U933 ( .A(G110), .B(n1178), .Z(G12) );
NOR4_X1 U934 ( .A1(n1222), .A2(n1046), .A3(n1188), .A4(n1187), .ZN(n1178) );
NAND2_X1 U935 ( .A1(n1049), .A2(n1050), .ZN(n1187) );
NAND2_X1 U936 ( .A1(G221), .A2(n1239), .ZN(n1050) );
INV_X1 U937 ( .A(n1238), .ZN(n1049) );
XNOR2_X1 U938 ( .A(n1078), .B(n1240), .ZN(n1238) );
NOR2_X1 U939 ( .A1(n1241), .A2(KEYINPUT42), .ZN(n1240) );
INV_X1 U940 ( .A(n1079), .ZN(n1241) );
NAND2_X1 U941 ( .A1(n1242), .A2(n1243), .ZN(n1079) );
XOR2_X1 U942 ( .A(n1244), .B(n1245), .Z(n1242) );
XOR2_X1 U943 ( .A(n1246), .B(n1160), .Z(n1245) );
XOR2_X1 U944 ( .A(n1091), .B(n1247), .Z(n1160) );
NOR2_X1 U945 ( .A1(KEYINPUT36), .A2(n1248), .ZN(n1247) );
XOR2_X1 U946 ( .A(n1249), .B(n1250), .Z(n1091) );
NAND2_X1 U947 ( .A1(KEYINPUT44), .A2(n1217), .ZN(n1249) );
XNOR2_X1 U948 ( .A(n1146), .B(n1251), .ZN(n1244) );
XNOR2_X1 U949 ( .A(n1095), .B(G110), .ZN(n1251) );
NAND2_X1 U950 ( .A1(G227), .A2(n1096), .ZN(n1146) );
XOR2_X1 U951 ( .A(G469), .B(KEYINPUT55), .Z(n1078) );
NAND2_X1 U952 ( .A1(n1058), .A2(n1252), .ZN(n1188) );
NAND2_X1 U953 ( .A1(n1033), .A2(n1253), .ZN(n1252) );
NAND4_X1 U954 ( .A1(G953), .A2(n1254), .A3(n1224), .A4(n1255), .ZN(n1253) );
INV_X1 U955 ( .A(G898), .ZN(n1255) );
XNOR2_X1 U956 ( .A(KEYINPUT22), .B(n1256), .ZN(n1254) );
NAND3_X1 U957 ( .A1(n1031), .A2(n1224), .A3(G952), .ZN(n1033) );
NAND2_X1 U958 ( .A1(G237), .A2(G234), .ZN(n1224) );
XOR2_X1 U959 ( .A(G953), .B(KEYINPUT8), .Z(n1031) );
NOR2_X1 U960 ( .A1(n1073), .A2(n1037), .ZN(n1058) );
INV_X1 U961 ( .A(n1075), .ZN(n1037) );
NAND2_X1 U962 ( .A1(G214), .A2(n1257), .ZN(n1075) );
INV_X1 U963 ( .A(n1036), .ZN(n1073) );
XNOR2_X1 U964 ( .A(n1258), .B(n1172), .ZN(n1036) );
AND2_X1 U965 ( .A1(G210), .A2(n1257), .ZN(n1172) );
NAND2_X1 U966 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
NAND3_X1 U967 ( .A1(n1243), .A2(n1261), .A3(n1262), .ZN(n1258) );
XOR2_X1 U968 ( .A(n1263), .B(KEYINPUT27), .Z(n1262) );
NAND2_X1 U969 ( .A1(n1170), .A2(n1264), .ZN(n1263) );
OR2_X1 U970 ( .A1(n1264), .A2(n1170), .ZN(n1261) );
XOR2_X1 U971 ( .A(n1265), .B(n1110), .Z(n1170) );
XOR2_X1 U972 ( .A(G110), .B(n1266), .Z(n1110) );
XOR2_X1 U973 ( .A(KEYINPUT33), .B(G122), .Z(n1266) );
NAND2_X1 U974 ( .A1(KEYINPUT50), .A2(n1109), .ZN(n1265) );
XNOR2_X1 U975 ( .A(n1267), .B(n1268), .ZN(n1109) );
XNOR2_X1 U976 ( .A(n1134), .B(n1269), .ZN(n1268) );
XNOR2_X1 U977 ( .A(KEYINPUT3), .B(n1237), .ZN(n1269) );
INV_X1 U978 ( .A(G101), .ZN(n1134) );
XOR2_X1 U979 ( .A(n1270), .B(n1248), .Z(n1267) );
XNOR2_X1 U980 ( .A(n1126), .B(G107), .ZN(n1248) );
INV_X1 U981 ( .A(G104), .ZN(n1126) );
NAND2_X1 U982 ( .A1(KEYINPUT34), .A2(n1271), .ZN(n1270) );
XNOR2_X1 U983 ( .A(n1272), .B(n1273), .ZN(n1264) );
XNOR2_X1 U984 ( .A(n1274), .B(KEYINPUT2), .ZN(n1273) );
NAND2_X1 U985 ( .A1(KEYINPUT57), .A2(n1275), .ZN(n1274) );
INV_X1 U986 ( .A(G125), .ZN(n1275) );
XOR2_X1 U987 ( .A(n1171), .B(n1142), .Z(n1272) );
AND2_X1 U988 ( .A1(G224), .A2(n1096), .ZN(n1171) );
INV_X1 U989 ( .A(n1212), .ZN(n1046) );
NOR2_X1 U990 ( .A1(n1074), .A2(n1209), .ZN(n1212) );
XNOR2_X1 U991 ( .A(n1276), .B(G475), .ZN(n1209) );
NAND2_X1 U992 ( .A1(n1243), .A2(n1122), .ZN(n1276) );
NAND2_X1 U993 ( .A1(n1277), .A2(n1278), .ZN(n1122) );
NAND2_X1 U994 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
XOR2_X1 U995 ( .A(KEYINPUT37), .B(n1281), .Z(n1277) );
NOR2_X1 U996 ( .A1(n1279), .A2(n1280), .ZN(n1281) );
NAND2_X1 U997 ( .A1(n1282), .A2(n1283), .ZN(n1280) );
NAND2_X1 U998 ( .A1(n1284), .A2(n1237), .ZN(n1283) );
XNOR2_X1 U999 ( .A(n1285), .B(KEYINPUT20), .ZN(n1284) );
NAND2_X1 U1000 ( .A1(n1286), .A2(G113), .ZN(n1282) );
XNOR2_X1 U1001 ( .A(KEYINPUT58), .B(n1287), .ZN(n1286) );
INV_X1 U1002 ( .A(n1285), .ZN(n1287) );
XOR2_X1 U1003 ( .A(G104), .B(G122), .Z(n1285) );
XOR2_X1 U1004 ( .A(n1288), .B(n1289), .Z(n1279) );
XNOR2_X1 U1005 ( .A(n1290), .B(n1291), .ZN(n1289) );
NOR4_X1 U1006 ( .A1(KEYINPUT12), .A2(G953), .A3(G237), .A4(n1292), .ZN(n1291) );
INV_X1 U1007 ( .A(G214), .ZN(n1292) );
XNOR2_X1 U1008 ( .A(G131), .B(G143), .ZN(n1290) );
NAND2_X1 U1009 ( .A1(n1293), .A2(KEYINPUT39), .ZN(n1288) );
XOR2_X1 U1010 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U1011 ( .A(G125), .B(KEYINPUT4), .ZN(n1294) );
XNOR2_X1 U1012 ( .A(n1296), .B(G478), .ZN(n1074) );
NAND2_X1 U1013 ( .A1(n1118), .A2(n1243), .ZN(n1296) );
XNOR2_X1 U1014 ( .A(n1297), .B(n1298), .ZN(n1118) );
NOR2_X1 U1015 ( .A1(KEYINPUT46), .A2(n1299), .ZN(n1298) );
XOR2_X1 U1016 ( .A(n1300), .B(n1301), .Z(n1299) );
NAND2_X1 U1017 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NAND2_X1 U1018 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
INV_X1 U1019 ( .A(G107), .ZN(n1305) );
XOR2_X1 U1020 ( .A(KEYINPUT38), .B(n1306), .Z(n1304) );
NAND2_X1 U1021 ( .A1(n1307), .A2(G107), .ZN(n1302) );
XNOR2_X1 U1022 ( .A(n1306), .B(KEYINPUT41), .ZN(n1307) );
XOR2_X1 U1023 ( .A(G116), .B(G122), .Z(n1306) );
NAND2_X1 U1024 ( .A1(KEYINPUT26), .A2(n1308), .ZN(n1300) );
XNOR2_X1 U1025 ( .A(n1217), .B(n1309), .ZN(n1308) );
XOR2_X1 U1026 ( .A(G143), .B(G134), .Z(n1309) );
NAND2_X1 U1027 ( .A1(n1310), .A2(G217), .ZN(n1297) );
NAND2_X1 U1028 ( .A1(n1230), .A2(n1069), .ZN(n1222) );
XOR2_X1 U1029 ( .A(n1311), .B(n1115), .Z(n1069) );
NAND2_X1 U1030 ( .A1(G217), .A2(n1239), .ZN(n1115) );
NAND2_X1 U1031 ( .A1(G234), .A2(n1259), .ZN(n1239) );
XNOR2_X1 U1032 ( .A(G902), .B(KEYINPUT45), .ZN(n1259) );
NAND2_X1 U1033 ( .A1(n1114), .A2(n1243), .ZN(n1311) );
XOR2_X1 U1034 ( .A(n1312), .B(n1313), .Z(n1114) );
XOR2_X1 U1035 ( .A(n1314), .B(n1315), .Z(n1313) );
NOR2_X1 U1036 ( .A1(G125), .A2(KEYINPUT10), .ZN(n1315) );
NOR2_X1 U1037 ( .A1(n1316), .A2(n1317), .ZN(n1314) );
XOR2_X1 U1038 ( .A(n1318), .B(KEYINPUT35), .Z(n1317) );
NAND2_X1 U1039 ( .A1(G110), .A2(n1319), .ZN(n1318) );
NOR2_X1 U1040 ( .A1(G110), .A2(n1319), .ZN(n1316) );
XNOR2_X1 U1041 ( .A(n1217), .B(G119), .ZN(n1319) );
INV_X1 U1042 ( .A(G128), .ZN(n1217) );
XOR2_X1 U1043 ( .A(n1320), .B(n1295), .Z(n1312) );
XNOR2_X1 U1044 ( .A(G146), .B(n1095), .ZN(n1295) );
INV_X1 U1045 ( .A(G140), .ZN(n1095) );
NAND2_X1 U1046 ( .A1(KEYINPUT53), .A2(n1321), .ZN(n1320) );
XNOR2_X1 U1047 ( .A(G137), .B(n1322), .ZN(n1321) );
NAND2_X1 U1048 ( .A1(n1310), .A2(G221), .ZN(n1322) );
AND2_X1 U1049 ( .A1(G234), .A2(n1096), .ZN(n1310) );
INV_X1 U1050 ( .A(n1213), .ZN(n1230) );
NAND2_X1 U1051 ( .A1(n1323), .A2(n1076), .ZN(n1213) );
NAND3_X1 U1052 ( .A1(n1243), .A2(n1143), .A3(n1324), .ZN(n1076) );
INV_X1 U1053 ( .A(G472), .ZN(n1143) );
XOR2_X1 U1054 ( .A(n1065), .B(KEYINPUT21), .Z(n1323) );
NAND2_X1 U1055 ( .A1(G472), .A2(n1325), .ZN(n1065) );
NAND2_X1 U1056 ( .A1(n1324), .A2(n1243), .ZN(n1325) );
XNOR2_X1 U1057 ( .A(n1256), .B(KEYINPUT47), .ZN(n1243) );
INV_X1 U1058 ( .A(G902), .ZN(n1256) );
XOR2_X1 U1059 ( .A(n1326), .B(n1327), .Z(n1324) );
XNOR2_X1 U1060 ( .A(n1132), .B(n1328), .ZN(n1327) );
NOR2_X1 U1061 ( .A1(KEYINPUT60), .A2(n1142), .ZN(n1328) );
XOR2_X1 U1062 ( .A(n1329), .B(n1250), .Z(n1142) );
XOR2_X1 U1063 ( .A(G146), .B(G143), .Z(n1250) );
XNOR2_X1 U1064 ( .A(G128), .B(KEYINPUT14), .ZN(n1329) );
NAND3_X1 U1065 ( .A1(n1260), .A2(n1096), .A3(G210), .ZN(n1132) );
INV_X1 U1066 ( .A(G953), .ZN(n1096) );
INV_X1 U1067 ( .A(G237), .ZN(n1260) );
XNOR2_X1 U1068 ( .A(n1246), .B(n1140), .ZN(n1326) );
XNOR2_X1 U1069 ( .A(n1237), .B(n1271), .ZN(n1140) );
XNOR2_X1 U1070 ( .A(G116), .B(G119), .ZN(n1271) );
INV_X1 U1071 ( .A(G113), .ZN(n1237) );
XNOR2_X1 U1072 ( .A(n1139), .B(G101), .ZN(n1246) );
XOR2_X1 U1073 ( .A(n1092), .B(KEYINPUT24), .Z(n1139) );
XOR2_X1 U1074 ( .A(G131), .B(n1330), .Z(n1092) );
XOR2_X1 U1075 ( .A(G137), .B(G134), .Z(n1330) );
endmodule


