//Key = 1111111011111001000000100000001101111000000010100000101000001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266;

XOR2_X1 U713 ( .A(n976), .B(n977), .Z(G9) );
NOR2_X1 U714 ( .A1(KEYINPUT27), .A2(n978), .ZN(n977) );
NAND4_X1 U715 ( .A1(n979), .A2(n980), .A3(n981), .A4(n982), .ZN(G75) );
NAND3_X1 U716 ( .A1(KEYINPUT38), .A2(n983), .A3(n984), .ZN(n982) );
NAND2_X1 U717 ( .A1(G952), .A2(n985), .ZN(n981) );
NAND4_X1 U718 ( .A1(n986), .A2(n987), .A3(n988), .A4(n983), .ZN(n985) );
NAND2_X1 U719 ( .A1(n989), .A2(n990), .ZN(n988) );
NAND2_X1 U720 ( .A1(n991), .A2(n992), .ZN(n990) );
NAND3_X1 U721 ( .A1(n993), .A2(n994), .A3(n995), .ZN(n992) );
NAND3_X1 U722 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n994) );
NAND2_X1 U723 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND2_X1 U724 ( .A1(n1001), .A2(n1002), .ZN(n997) );
XNOR2_X1 U725 ( .A(n999), .B(KEYINPUT46), .ZN(n1001) );
NAND2_X1 U726 ( .A1(n1003), .A2(n1004), .ZN(n996) );
NAND2_X1 U727 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND3_X1 U728 ( .A1(n999), .A2(n1007), .A3(n1003), .ZN(n991) );
NAND3_X1 U729 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1007) );
NAND2_X1 U730 ( .A1(n1011), .A2(n993), .ZN(n1010) );
NAND2_X1 U731 ( .A1(n995), .A2(n1012), .ZN(n1009) );
OR2_X1 U732 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U733 ( .A1(n1015), .A2(n1016), .ZN(n1008) );
XOR2_X1 U734 ( .A(KEYINPUT58), .B(n993), .Z(n1016) );
OR2_X1 U735 ( .A1(n983), .A2(KEYINPUT38), .ZN(n979) );
NAND4_X1 U736 ( .A1(n1003), .A2(n999), .A3(n995), .A4(n993), .ZN(n983) );
XOR2_X1 U737 ( .A(n1017), .B(n1018), .Z(G72) );
NOR2_X1 U738 ( .A1(KEYINPUT20), .A2(n1019), .ZN(n1018) );
XOR2_X1 U739 ( .A(n1020), .B(n1021), .Z(n1019) );
NOR2_X1 U740 ( .A1(n986), .A2(G953), .ZN(n1021) );
NOR3_X1 U741 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1020) );
NOR2_X1 U742 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
XOR2_X1 U743 ( .A(KEYINPUT42), .B(n1027), .Z(n1022) );
AND2_X1 U744 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
XNOR2_X1 U745 ( .A(n1028), .B(n1029), .ZN(n1025) );
XOR2_X1 U746 ( .A(KEYINPUT44), .B(KEYINPUT29), .Z(n1029) );
XOR2_X1 U747 ( .A(n1030), .B(n1031), .Z(n1028) );
NAND2_X1 U748 ( .A1(KEYINPUT1), .A2(G140), .ZN(n1030) );
NAND2_X1 U749 ( .A1(n1032), .A2(n1033), .ZN(n1026) );
NAND2_X1 U750 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
XOR2_X1 U751 ( .A(n1036), .B(KEYINPUT61), .Z(n1032) );
OR2_X1 U752 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
XOR2_X1 U753 ( .A(n1037), .B(n1038), .Z(n1034) );
XNOR2_X1 U754 ( .A(n1039), .B(n1040), .ZN(n1038) );
NOR2_X1 U755 ( .A1(KEYINPUT51), .A2(n1041), .ZN(n1040) );
NAND2_X1 U756 ( .A1(KEYINPUT0), .A2(G137), .ZN(n1039) );
NAND2_X1 U757 ( .A1(n1042), .A2(n1043), .ZN(n1017) );
NAND2_X1 U758 ( .A1(G900), .A2(G227), .ZN(n1043) );
XOR2_X1 U759 ( .A(n1044), .B(n1045), .Z(G69) );
XOR2_X1 U760 ( .A(n1046), .B(n1047), .Z(n1045) );
NOR2_X1 U761 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XNOR2_X1 U762 ( .A(n1050), .B(n1051), .ZN(n1049) );
NAND2_X1 U763 ( .A1(KEYINPUT33), .A2(n1052), .ZN(n1050) );
XOR2_X1 U764 ( .A(n1053), .B(n1054), .Z(n1052) );
XOR2_X1 U765 ( .A(n1055), .B(G104), .Z(n1054) );
NAND2_X1 U766 ( .A1(n1056), .A2(KEYINPUT4), .ZN(n1055) );
XOR2_X1 U767 ( .A(n1057), .B(G113), .Z(n1056) );
NAND2_X1 U768 ( .A1(n1042), .A2(n1058), .ZN(n1046) );
NAND2_X1 U769 ( .A1(G898), .A2(G224), .ZN(n1058) );
XOR2_X1 U770 ( .A(G953), .B(KEYINPUT37), .Z(n1042) );
NAND2_X1 U771 ( .A1(n980), .A2(n1059), .ZN(n1044) );
NOR3_X1 U772 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(G66) );
NOR3_X1 U773 ( .A1(n1063), .A2(n1064), .A3(n980), .ZN(n1062) );
INV_X1 U774 ( .A(KEYINPUT45), .ZN(n1063) );
NOR2_X1 U775 ( .A1(KEYINPUT45), .A2(n1065), .ZN(n1061) );
XOR2_X1 U776 ( .A(n1066), .B(n1067), .Z(n1060) );
NOR2_X1 U777 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U778 ( .A1(n1070), .A2(n1071), .ZN(G63) );
XOR2_X1 U779 ( .A(n1072), .B(n1073), .Z(n1071) );
NOR2_X1 U780 ( .A1(n1074), .A2(n1069), .ZN(n1073) );
NOR2_X1 U781 ( .A1(n1070), .A2(n1075), .ZN(G60) );
XOR2_X1 U782 ( .A(n1076), .B(n1077), .Z(n1075) );
XOR2_X1 U783 ( .A(KEYINPUT9), .B(n1078), .Z(n1077) );
NOR2_X1 U784 ( .A1(n1079), .A2(n1069), .ZN(n1078) );
INV_X1 U785 ( .A(G475), .ZN(n1079) );
XOR2_X1 U786 ( .A(n1080), .B(n1081), .Z(G6) );
NAND4_X1 U787 ( .A1(n1000), .A2(n993), .A3(n1082), .A4(n1083), .ZN(n1081) );
XNOR2_X1 U788 ( .A(KEYINPUT54), .B(n1084), .ZN(n1083) );
NOR3_X1 U789 ( .A1(n1070), .A2(n1085), .A3(n1086), .ZN(G57) );
NOR2_X1 U790 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U791 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR3_X1 U792 ( .A1(n1091), .A2(KEYINPUT25), .A3(n1092), .ZN(n1090) );
AND2_X1 U793 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
INV_X1 U794 ( .A(KEYINPUT52), .ZN(n1091) );
NOR2_X1 U795 ( .A1(n1093), .A2(n1094), .ZN(n1085) );
NOR2_X1 U796 ( .A1(KEYINPUT25), .A2(n1092), .ZN(n1093) );
XOR2_X1 U797 ( .A(n1095), .B(n1096), .Z(n1092) );
XOR2_X1 U798 ( .A(KEYINPUT53), .B(n1097), .Z(n1096) );
NOR2_X1 U799 ( .A1(n1098), .A2(n1069), .ZN(n1097) );
INV_X1 U800 ( .A(G472), .ZN(n1098) );
NOR2_X1 U801 ( .A1(n1070), .A2(n1099), .ZN(G54) );
XOR2_X1 U802 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR3_X1 U803 ( .A1(n1069), .A2(KEYINPUT43), .A3(n1102), .ZN(n1101) );
INV_X1 U804 ( .A(G469), .ZN(n1102) );
NOR2_X1 U805 ( .A1(n1070), .A2(n1103), .ZN(G51) );
XOR2_X1 U806 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U807 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U808 ( .A1(n1108), .A2(n1069), .ZN(n1107) );
NAND2_X1 U809 ( .A1(G902), .A2(n1109), .ZN(n1069) );
NAND2_X1 U810 ( .A1(n986), .A2(n987), .ZN(n1109) );
INV_X1 U811 ( .A(n1059), .ZN(n987) );
NAND4_X1 U812 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1059) );
NOR4_X1 U813 ( .A1(n1114), .A2(n1115), .A3(n976), .A4(n1116), .ZN(n1113) );
AND3_X1 U814 ( .A1(n1117), .A2(n1002), .A3(n993), .ZN(n976) );
AND2_X1 U815 ( .A1(n1118), .A2(n1119), .ZN(n1112) );
NAND3_X1 U816 ( .A1(n993), .A2(n1117), .A3(n1000), .ZN(n1111) );
NAND2_X1 U817 ( .A1(n1120), .A2(n1121), .ZN(n1110) );
XOR2_X1 U818 ( .A(KEYINPUT56), .B(n1122), .Z(n1121) );
AND4_X1 U819 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n986) );
NOR4_X1 U820 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1126) );
AND3_X1 U821 ( .A1(n1014), .A2(n1002), .A3(n1131), .ZN(n1127) );
NOR2_X1 U822 ( .A1(n1132), .A2(n1133), .ZN(n1125) );
NOR2_X1 U823 ( .A1(KEYINPUT50), .A2(n1134), .ZN(n1106) );
XNOR2_X1 U824 ( .A(n1135), .B(n1136), .ZN(n1134) );
INV_X1 U825 ( .A(n1065), .ZN(n1070) );
NAND2_X1 U826 ( .A1(n1064), .A2(G953), .ZN(n1065) );
XOR2_X1 U827 ( .A(n984), .B(KEYINPUT47), .Z(n1064) );
INV_X1 U828 ( .A(G952), .ZN(n984) );
XNOR2_X1 U829 ( .A(n1123), .B(n1137), .ZN(G48) );
NOR2_X1 U830 ( .A1(KEYINPUT23), .A2(n1138), .ZN(n1137) );
NAND4_X1 U831 ( .A1(n1139), .A2(n1000), .A3(n1082), .A4(n1140), .ZN(n1123) );
XOR2_X1 U832 ( .A(G143), .B(n1130), .Z(G45) );
AND3_X1 U833 ( .A1(n1014), .A2(n1141), .A3(n1142), .ZN(n1130) );
XNOR2_X1 U834 ( .A(G140), .B(n1124), .ZN(G42) );
NAND2_X1 U835 ( .A1(n1131), .A2(n1143), .ZN(n1124) );
XOR2_X1 U836 ( .A(n1133), .B(n1144), .Z(G39) );
NOR2_X1 U837 ( .A1(KEYINPUT40), .A2(n1145), .ZN(n1144) );
AND3_X1 U838 ( .A1(n1131), .A2(n1139), .A3(n1003), .ZN(n1133) );
XOR2_X1 U839 ( .A(n1146), .B(n1147), .Z(G36) );
XOR2_X1 U840 ( .A(n1148), .B(KEYINPUT16), .Z(n1147) );
NAND3_X1 U841 ( .A1(n1149), .A2(n1014), .A3(n1150), .ZN(n1146) );
AND3_X1 U842 ( .A1(n1002), .A2(n1140), .A3(n1015), .ZN(n1150) );
AND2_X1 U843 ( .A1(n1151), .A2(n1152), .ZN(n1002) );
XNOR2_X1 U844 ( .A(n999), .B(KEYINPUT36), .ZN(n1149) );
XNOR2_X1 U845 ( .A(n1129), .B(n1153), .ZN(G33) );
NOR2_X1 U846 ( .A1(G131), .A2(KEYINPUT59), .ZN(n1153) );
AND3_X1 U847 ( .A1(n1131), .A2(n1000), .A3(n1014), .ZN(n1129) );
AND3_X1 U848 ( .A1(n1015), .A2(n1140), .A3(n999), .ZN(n1131) );
NOR2_X1 U849 ( .A1(n1005), .A2(n1154), .ZN(n999) );
AND2_X1 U850 ( .A1(G214), .A2(n1155), .ZN(n1154) );
XOR2_X1 U851 ( .A(G128), .B(n1128), .Z(G30) );
AND3_X1 U852 ( .A1(n1151), .A2(n1139), .A3(n1142), .ZN(n1128) );
AND3_X1 U853 ( .A1(n1152), .A2(n1140), .A3(n1082), .ZN(n1142) );
NAND2_X1 U854 ( .A1(n1156), .A2(n1157), .ZN(G3) );
NAND2_X1 U855 ( .A1(G101), .A2(n1119), .ZN(n1157) );
XOR2_X1 U856 ( .A(KEYINPUT60), .B(n1158), .Z(n1156) );
NOR2_X1 U857 ( .A1(G101), .A2(n1119), .ZN(n1158) );
NAND3_X1 U858 ( .A1(n1003), .A2(n1117), .A3(n1014), .ZN(n1119) );
XOR2_X1 U859 ( .A(G125), .B(n1132), .Z(G27) );
AND4_X1 U860 ( .A1(n995), .A2(n1143), .A3(n1120), .A4(n1140), .ZN(n1132) );
NAND2_X1 U861 ( .A1(n1159), .A2(n1160), .ZN(n1140) );
NAND3_X1 U862 ( .A1(G902), .A2(n1161), .A3(n1023), .ZN(n1160) );
NOR2_X1 U863 ( .A1(n980), .A2(G900), .ZN(n1023) );
XOR2_X1 U864 ( .A(KEYINPUT35), .B(n989), .Z(n1159) );
INV_X1 U865 ( .A(n1162), .ZN(n989) );
AND3_X1 U866 ( .A1(n1013), .A2(n1163), .A3(n1000), .ZN(n1143) );
XOR2_X1 U867 ( .A(G122), .B(n1115), .Z(G24) );
AND3_X1 U868 ( .A1(n993), .A2(n1141), .A3(n1164), .ZN(n1115) );
AND2_X1 U869 ( .A1(n1013), .A2(n1165), .ZN(n993) );
XOR2_X1 U870 ( .A(n1166), .B(G119), .Z(G21) );
NAND2_X1 U871 ( .A1(KEYINPUT15), .A2(n1167), .ZN(n1166) );
NAND2_X1 U872 ( .A1(n1122), .A2(n1120), .ZN(n1167) );
AND4_X1 U873 ( .A1(n1003), .A2(n1139), .A3(n995), .A4(n1084), .ZN(n1122) );
NOR2_X1 U874 ( .A1(n1165), .A2(n1013), .ZN(n1139) );
XOR2_X1 U875 ( .A(G116), .B(n1114), .Z(G18) );
AND3_X1 U876 ( .A1(n1151), .A2(n1014), .A3(n1164), .ZN(n1114) );
AND4_X1 U877 ( .A1(n995), .A2(n1120), .A3(n1152), .A4(n1084), .ZN(n1164) );
XOR2_X1 U878 ( .A(n1118), .B(n1168), .Z(G15) );
NOR2_X1 U879 ( .A1(G113), .A2(KEYINPUT14), .ZN(n1168) );
NAND4_X1 U880 ( .A1(n1014), .A2(n995), .A3(n1169), .A4(n1000), .ZN(n1118) );
NOR2_X1 U881 ( .A1(n1152), .A2(n1151), .ZN(n1000) );
AND2_X1 U882 ( .A1(n1084), .A2(n1120), .ZN(n1169) );
AND2_X1 U883 ( .A1(n1011), .A2(n1170), .ZN(n995) );
NOR2_X1 U884 ( .A1(n1163), .A2(n1013), .ZN(n1014) );
XOR2_X1 U885 ( .A(G110), .B(n1116), .Z(G12) );
AND4_X1 U886 ( .A1(n1003), .A2(n1117), .A3(n1013), .A4(n1163), .ZN(n1116) );
INV_X1 U887 ( .A(n1165), .ZN(n1163) );
XOR2_X1 U888 ( .A(n1068), .B(n1171), .Z(n1165) );
NOR2_X1 U889 ( .A1(n1066), .A2(n1172), .ZN(n1171) );
XOR2_X1 U890 ( .A(n1173), .B(n1174), .Z(n1066) );
XOR2_X1 U891 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U892 ( .A(G128), .B(n1177), .Z(n1176) );
NOR2_X1 U893 ( .A1(KEYINPUT18), .A2(n1178), .ZN(n1177) );
XOR2_X1 U894 ( .A(n1179), .B(G137), .Z(n1178) );
NAND2_X1 U895 ( .A1(G221), .A2(n1180), .ZN(n1179) );
NOR2_X1 U896 ( .A1(KEYINPUT17), .A2(n1181), .ZN(n1175) );
XOR2_X1 U897 ( .A(n1182), .B(n1183), .Z(n1173) );
XOR2_X1 U898 ( .A(n1184), .B(n1031), .Z(n1182) );
NAND2_X1 U899 ( .A1(KEYINPUT11), .A2(n1185), .ZN(n1184) );
INV_X1 U900 ( .A(G119), .ZN(n1185) );
NAND2_X1 U901 ( .A1(G217), .A2(n1186), .ZN(n1068) );
XOR2_X1 U902 ( .A(n1187), .B(G472), .Z(n1013) );
NAND2_X1 U903 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U904 ( .A(n1095), .B(n1087), .Z(n1188) );
INV_X1 U905 ( .A(n1094), .ZN(n1087) );
XOR2_X1 U906 ( .A(n1190), .B(G101), .Z(n1094) );
NAND2_X1 U907 ( .A1(G210), .A2(n1191), .ZN(n1190) );
XOR2_X1 U908 ( .A(n1192), .B(n1193), .Z(n1095) );
XOR2_X1 U909 ( .A(G116), .B(n1194), .Z(n1193) );
XOR2_X1 U910 ( .A(KEYINPUT24), .B(G119), .Z(n1194) );
XOR2_X1 U911 ( .A(n1195), .B(n1196), .Z(n1192) );
XOR2_X1 U912 ( .A(n1197), .B(n1198), .Z(n1195) );
NAND2_X1 U913 ( .A1(KEYINPUT6), .A2(G113), .ZN(n1197) );
AND2_X1 U914 ( .A1(n1082), .A2(n1084), .ZN(n1117) );
NAND2_X1 U915 ( .A1(n1162), .A2(n1199), .ZN(n1084) );
NAND3_X1 U916 ( .A1(G902), .A2(n1161), .A3(n1048), .ZN(n1199) );
NOR2_X1 U917 ( .A1(n980), .A2(G898), .ZN(n1048) );
NAND3_X1 U918 ( .A1(n1161), .A2(n980), .A3(G952), .ZN(n1162) );
NAND2_X1 U919 ( .A1(G237), .A2(G234), .ZN(n1161) );
AND2_X1 U920 ( .A1(n1015), .A2(n1120), .ZN(n1082) );
INV_X1 U921 ( .A(n1006), .ZN(n1120) );
NAND2_X1 U922 ( .A1(n1005), .A2(n1200), .ZN(n1006) );
NAND2_X1 U923 ( .A1(G214), .A2(n1155), .ZN(n1200) );
XOR2_X1 U924 ( .A(n1201), .B(n1108), .Z(n1005) );
NAND2_X1 U925 ( .A1(G210), .A2(n1155), .ZN(n1108) );
NAND2_X1 U926 ( .A1(n1202), .A2(n1203), .ZN(n1155) );
INV_X1 U927 ( .A(G237), .ZN(n1203) );
NAND2_X1 U928 ( .A1(n1189), .A2(n1204), .ZN(n1201) );
XOR2_X1 U929 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U930 ( .A(n1136), .B(n1207), .Z(n1206) );
NOR3_X1 U931 ( .A1(KEYINPUT19), .A2(n1208), .A3(n1209), .ZN(n1207) );
AND3_X1 U932 ( .A1(KEYINPUT41), .A2(n1210), .A3(n1198), .ZN(n1209) );
NOR2_X1 U933 ( .A1(KEYINPUT41), .A2(n1135), .ZN(n1208) );
XNOR2_X1 U934 ( .A(n1198), .B(n1210), .ZN(n1135) );
INV_X1 U935 ( .A(n1031), .ZN(n1210) );
XNOR2_X1 U936 ( .A(n1211), .B(n1212), .ZN(n1198) );
XNOR2_X1 U937 ( .A(n1181), .B(n1213), .ZN(n1212) );
XNOR2_X1 U938 ( .A(G143), .B(KEYINPUT63), .ZN(n1211) );
AND2_X1 U939 ( .A1(G224), .A2(n980), .ZN(n1136) );
NOR2_X1 U940 ( .A1(KEYINPUT26), .A2(n1104), .ZN(n1205) );
XNOR2_X1 U941 ( .A(n1214), .B(n1215), .ZN(n1104) );
XOR2_X1 U942 ( .A(n1057), .B(n1216), .Z(n1215) );
NAND3_X1 U943 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1057) );
NAND2_X1 U944 ( .A1(G116), .A2(n1220), .ZN(n1219) );
OR3_X1 U945 ( .A1(n1220), .A2(n1221), .A3(G119), .ZN(n1218) );
INV_X1 U946 ( .A(KEYINPUT10), .ZN(n1220) );
NAND2_X1 U947 ( .A1(G119), .A2(n1221), .ZN(n1217) );
NAND2_X1 U948 ( .A1(KEYINPUT12), .A2(n1222), .ZN(n1221) );
XOR2_X1 U949 ( .A(n1053), .B(n1051), .Z(n1214) );
XOR2_X1 U950 ( .A(G110), .B(G122), .Z(n1051) );
XOR2_X1 U951 ( .A(n1223), .B(G101), .Z(n1053) );
NAND2_X1 U952 ( .A1(n1224), .A2(KEYINPUT8), .ZN(n1223) );
XOR2_X1 U953 ( .A(n978), .B(KEYINPUT57), .Z(n1224) );
NOR2_X1 U954 ( .A1(n1011), .A2(n1225), .ZN(n1015) );
INV_X1 U955 ( .A(n1170), .ZN(n1225) );
NAND2_X1 U956 ( .A1(G221), .A2(n1186), .ZN(n1170) );
NAND2_X1 U957 ( .A1(G234), .A2(n1202), .ZN(n1186) );
XNOR2_X1 U958 ( .A(G902), .B(KEYINPUT39), .ZN(n1202) );
XOR2_X1 U959 ( .A(n1226), .B(G469), .Z(n1011) );
NAND3_X1 U960 ( .A1(n1227), .A2(n1228), .A3(n1189), .ZN(n1226) );
NAND2_X1 U961 ( .A1(KEYINPUT30), .A2(n1100), .ZN(n1228) );
XOR2_X1 U962 ( .A(n1229), .B(n1230), .Z(n1100) );
OR3_X1 U963 ( .A1(n1229), .A2(n1230), .A3(KEYINPUT30), .ZN(n1227) );
XNOR2_X1 U964 ( .A(n1231), .B(n1232), .ZN(n1230) );
XOR2_X1 U965 ( .A(n1233), .B(n1234), .Z(n1232) );
XOR2_X1 U966 ( .A(n1080), .B(G107), .Z(n1234) );
NAND2_X1 U967 ( .A1(KEYINPUT31), .A2(n1235), .ZN(n1233) );
INV_X1 U968 ( .A(G101), .ZN(n1235) );
XNOR2_X1 U969 ( .A(n1196), .B(n1035), .ZN(n1231) );
XOR2_X1 U970 ( .A(n1181), .B(n1236), .Z(n1035) );
XNOR2_X1 U971 ( .A(n1237), .B(n1238), .ZN(n1236) );
NOR2_X1 U972 ( .A1(G143), .A2(KEYINPUT21), .ZN(n1238) );
NAND2_X1 U973 ( .A1(KEYINPUT2), .A2(n1213), .ZN(n1237) );
XNOR2_X1 U974 ( .A(G128), .B(KEYINPUT62), .ZN(n1213) );
XOR2_X1 U975 ( .A(n1239), .B(n1041), .Z(n1196) );
XOR2_X1 U976 ( .A(n1145), .B(n1240), .Z(n1239) );
NOR2_X1 U977 ( .A1(KEYINPUT49), .A2(n1037), .ZN(n1240) );
XOR2_X1 U978 ( .A(n1148), .B(KEYINPUT5), .Z(n1037) );
INV_X1 U979 ( .A(G134), .ZN(n1148) );
INV_X1 U980 ( .A(G137), .ZN(n1145) );
XOR2_X1 U981 ( .A(n1241), .B(n1183), .Z(n1229) );
XOR2_X1 U982 ( .A(G110), .B(G140), .Z(n1183) );
NAND2_X1 U983 ( .A1(G227), .A2(n980), .ZN(n1241) );
NOR2_X1 U984 ( .A1(n1152), .A2(n1141), .ZN(n1003) );
INV_X1 U985 ( .A(n1151), .ZN(n1141) );
XOR2_X1 U986 ( .A(n1242), .B(G475), .Z(n1151) );
NAND2_X1 U987 ( .A1(n1189), .A2(n1076), .ZN(n1242) );
XNOR2_X1 U988 ( .A(n1243), .B(n1244), .ZN(n1076) );
XOR2_X1 U989 ( .A(n1216), .B(n1245), .Z(n1244) );
XNOR2_X1 U990 ( .A(n1246), .B(n1041), .ZN(n1245) );
XNOR2_X1 U991 ( .A(G131), .B(KEYINPUT3), .ZN(n1041) );
NAND2_X1 U992 ( .A1(G214), .A2(n1191), .ZN(n1246) );
NOR2_X1 U993 ( .A1(G953), .A2(G237), .ZN(n1191) );
XOR2_X1 U994 ( .A(n1080), .B(G113), .Z(n1216) );
INV_X1 U995 ( .A(G104), .ZN(n1080) );
XOR2_X1 U996 ( .A(n1247), .B(n1248), .Z(n1243) );
NOR2_X1 U997 ( .A1(G122), .A2(KEYINPUT13), .ZN(n1248) );
XOR2_X1 U998 ( .A(n1249), .B(G143), .Z(n1247) );
NAND2_X1 U999 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
OR2_X1 U1000 ( .A1(n1252), .A2(n1181), .ZN(n1251) );
XOR2_X1 U1001 ( .A(n1253), .B(KEYINPUT28), .Z(n1250) );
NAND2_X1 U1002 ( .A1(n1252), .A2(n1181), .ZN(n1253) );
XNOR2_X1 U1003 ( .A(n1138), .B(KEYINPUT34), .ZN(n1181) );
INV_X1 U1004 ( .A(G146), .ZN(n1138) );
XOR2_X1 U1005 ( .A(G140), .B(n1031), .Z(n1252) );
XOR2_X1 U1006 ( .A(G125), .B(KEYINPUT22), .Z(n1031) );
XNOR2_X1 U1007 ( .A(n1074), .B(n1254), .ZN(n1152) );
NOR2_X1 U1008 ( .A1(n1072), .A2(n1172), .ZN(n1254) );
INV_X1 U1009 ( .A(n1189), .ZN(n1172) );
XNOR2_X1 U1010 ( .A(G902), .B(KEYINPUT7), .ZN(n1189) );
XOR2_X1 U1011 ( .A(n1255), .B(n1256), .Z(n1072) );
XOR2_X1 U1012 ( .A(n1257), .B(n1258), .Z(n1256) );
NAND2_X1 U1013 ( .A1(n1180), .A2(G217), .ZN(n1258) );
AND2_X1 U1014 ( .A1(G234), .A2(n980), .ZN(n1180) );
INV_X1 U1015 ( .A(G953), .ZN(n980) );
NAND2_X1 U1016 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
NAND2_X1 U1017 ( .A1(G116), .A2(n1261), .ZN(n1260) );
INV_X1 U1018 ( .A(G122), .ZN(n1261) );
XOR2_X1 U1019 ( .A(n1262), .B(KEYINPUT55), .Z(n1259) );
NAND2_X1 U1020 ( .A1(G122), .A2(n1222), .ZN(n1262) );
INV_X1 U1021 ( .A(G116), .ZN(n1222) );
XOR2_X1 U1022 ( .A(n1263), .B(n1264), .Z(n1255) );
NOR2_X1 U1023 ( .A1(KEYINPUT32), .A2(n1265), .ZN(n1264) );
XOR2_X1 U1024 ( .A(G128), .B(n1266), .Z(n1265) );
XOR2_X1 U1025 ( .A(G143), .B(G134), .Z(n1266) );
XOR2_X1 U1026 ( .A(n978), .B(KEYINPUT48), .Z(n1263) );
INV_X1 U1027 ( .A(G107), .ZN(n978) );
INV_X1 U1028 ( .A(G478), .ZN(n1074) );
endmodule


