//Key = 1001111110111101111010101101110011101000000110101101110011111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257;

XOR2_X1 U705 ( .A(G107), .B(n964), .Z(G9) );
NAND4_X1 U706 ( .A1(n965), .A2(n966), .A3(n967), .A4(n968), .ZN(G75) );
NAND3_X1 U707 ( .A1(KEYINPUT42), .A2(n969), .A3(n970), .ZN(n968) );
INV_X1 U708 ( .A(G952), .ZN(n970) );
NAND2_X1 U709 ( .A1(G952), .A2(n971), .ZN(n967) );
NAND3_X1 U710 ( .A1(n972), .A2(n969), .A3(n973), .ZN(n971) );
NAND2_X1 U711 ( .A1(n974), .A2(n975), .ZN(n972) );
NAND2_X1 U712 ( .A1(n976), .A2(n977), .ZN(n975) );
NAND3_X1 U713 ( .A1(n978), .A2(n979), .A3(n980), .ZN(n977) );
NAND2_X1 U714 ( .A1(n981), .A2(n982), .ZN(n979) );
NAND2_X1 U715 ( .A1(n983), .A2(n984), .ZN(n982) );
OR2_X1 U716 ( .A1(n985), .A2(n986), .ZN(n984) );
NAND2_X1 U717 ( .A1(n987), .A2(n988), .ZN(n981) );
XOR2_X1 U718 ( .A(n989), .B(n990), .Z(n987) );
NAND2_X1 U719 ( .A1(n991), .A2(KEYINPUT22), .ZN(n989) );
NAND3_X1 U720 ( .A1(n983), .A2(n992), .A3(n988), .ZN(n976) );
NAND2_X1 U721 ( .A1(n993), .A2(n994), .ZN(n992) );
NAND2_X1 U722 ( .A1(n978), .A2(n995), .ZN(n994) );
NAND2_X1 U723 ( .A1(n996), .A2(n997), .ZN(n995) );
NAND2_X1 U724 ( .A1(n980), .A2(n998), .ZN(n993) );
NAND2_X1 U725 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND2_X1 U726 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
XOR2_X1 U727 ( .A(KEYINPUT57), .B(n1003), .Z(n1002) );
INV_X1 U728 ( .A(n1004), .ZN(n974) );
OR2_X1 U729 ( .A1(n969), .A2(KEYINPUT42), .ZN(n965) );
NAND4_X1 U730 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n969) );
NOR3_X1 U731 ( .A1(n1009), .A2(n991), .A3(n1010), .ZN(n1008) );
NOR2_X1 U732 ( .A1(G469), .A2(n1011), .ZN(n1010) );
NAND3_X1 U733 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1009) );
NOR3_X1 U734 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1007) );
XOR2_X1 U735 ( .A(n1018), .B(KEYINPUT27), .Z(n1017) );
NAND2_X1 U736 ( .A1(n1019), .A2(n1011), .ZN(n1018) );
XNOR2_X1 U737 ( .A(G469), .B(KEYINPUT32), .ZN(n1019) );
XNOR2_X1 U738 ( .A(n1020), .B(n1021), .ZN(n1016) );
NOR2_X1 U739 ( .A1(G478), .A2(KEYINPUT41), .ZN(n1021) );
XOR2_X1 U740 ( .A(n1022), .B(G472), .Z(n1005) );
XOR2_X1 U741 ( .A(n1023), .B(n1024), .Z(G72) );
XOR2_X1 U742 ( .A(n1025), .B(n1026), .Z(n1024) );
NOR3_X1 U743 ( .A1(n1027), .A2(KEYINPUT21), .A3(n1028), .ZN(n1026) );
XNOR2_X1 U744 ( .A(G953), .B(n1029), .ZN(n1027) );
XNOR2_X1 U745 ( .A(KEYINPUT44), .B(KEYINPUT0), .ZN(n1029) );
NAND2_X1 U746 ( .A1(n1030), .A2(n1031), .ZN(n1025) );
NAND2_X1 U747 ( .A1(G953), .A2(n1032), .ZN(n1031) );
XOR2_X1 U748 ( .A(n1033), .B(n1034), .Z(n1030) );
XOR2_X1 U749 ( .A(n1035), .B(n1036), .Z(n1034) );
NAND2_X1 U750 ( .A1(KEYINPUT49), .A2(G140), .ZN(n1035) );
XOR2_X1 U751 ( .A(n1037), .B(n1038), .Z(n1033) );
XNOR2_X1 U752 ( .A(G125), .B(n1039), .ZN(n1038) );
NAND2_X1 U753 ( .A1(KEYINPUT20), .A2(n1040), .ZN(n1037) );
NAND2_X1 U754 ( .A1(G953), .A2(n1041), .ZN(n1023) );
NAND2_X1 U755 ( .A1(G900), .A2(G227), .ZN(n1041) );
XOR2_X1 U756 ( .A(n1042), .B(n1043), .Z(G69) );
XOR2_X1 U757 ( .A(n1044), .B(n1045), .Z(n1043) );
NAND2_X1 U758 ( .A1(G953), .A2(n1046), .ZN(n1045) );
NAND2_X1 U759 ( .A1(G898), .A2(G224), .ZN(n1046) );
NAND2_X1 U760 ( .A1(n1047), .A2(n1048), .ZN(n1044) );
NAND2_X1 U761 ( .A1(G953), .A2(n1049), .ZN(n1048) );
XOR2_X1 U762 ( .A(n1050), .B(n1051), .Z(n1047) );
XOR2_X1 U763 ( .A(n1052), .B(n1053), .Z(n1051) );
NOR2_X1 U764 ( .A1(KEYINPUT39), .A2(n1054), .ZN(n1053) );
XNOR2_X1 U765 ( .A(G122), .B(G110), .ZN(n1054) );
XNOR2_X1 U766 ( .A(G113), .B(KEYINPUT30), .ZN(n1050) );
NOR2_X1 U767 ( .A1(n1055), .A2(G953), .ZN(n1042) );
NOR2_X1 U768 ( .A1(n1056), .A2(n1057), .ZN(G66) );
XOR2_X1 U769 ( .A(n1058), .B(n1059), .Z(n1057) );
NAND2_X1 U770 ( .A1(KEYINPUT11), .A2(n1060), .ZN(n1059) );
INV_X1 U771 ( .A(n1061), .ZN(n1060) );
NAND2_X1 U772 ( .A1(n1062), .A2(G217), .ZN(n1058) );
NOR2_X1 U773 ( .A1(n1063), .A2(n1064), .ZN(G63) );
XOR2_X1 U774 ( .A(KEYINPUT37), .B(n1056), .Z(n1064) );
NOR3_X1 U775 ( .A1(n1020), .A2(n1065), .A3(n1066), .ZN(n1063) );
AND3_X1 U776 ( .A1(n1067), .A2(G478), .A3(n1062), .ZN(n1066) );
NOR2_X1 U777 ( .A1(n1068), .A2(n1067), .ZN(n1065) );
NOR2_X1 U778 ( .A1(n973), .A2(n1069), .ZN(n1068) );
NOR2_X1 U779 ( .A1(n1056), .A2(n1070), .ZN(G60) );
XOR2_X1 U780 ( .A(n1071), .B(n1072), .Z(n1070) );
NAND2_X1 U781 ( .A1(n1062), .A2(G475), .ZN(n1071) );
XOR2_X1 U782 ( .A(n1073), .B(n1074), .Z(G6) );
XNOR2_X1 U783 ( .A(KEYINPUT4), .B(n1075), .ZN(n1074) );
NOR2_X1 U784 ( .A1(n1056), .A2(n1076), .ZN(G57) );
XOR2_X1 U785 ( .A(n1077), .B(n1078), .Z(n1076) );
XOR2_X1 U786 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND3_X1 U787 ( .A1(n1081), .A2(n1082), .A3(KEYINPUT3), .ZN(n1079) );
OR3_X1 U788 ( .A1(n1083), .A2(n1084), .A3(KEYINPUT43), .ZN(n1082) );
NAND2_X1 U789 ( .A1(n1085), .A2(KEYINPUT43), .ZN(n1081) );
XOR2_X1 U790 ( .A(n1084), .B(n1083), .Z(n1085) );
XOR2_X1 U791 ( .A(n1086), .B(KEYINPUT17), .Z(n1083) );
XOR2_X1 U792 ( .A(n1087), .B(KEYINPUT40), .Z(n1077) );
NAND2_X1 U793 ( .A1(n1062), .A2(G472), .ZN(n1087) );
NOR2_X1 U794 ( .A1(n1056), .A2(n1088), .ZN(G54) );
XOR2_X1 U795 ( .A(n1089), .B(n1090), .Z(n1088) );
XOR2_X1 U796 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U797 ( .A1(KEYINPUT62), .A2(n1093), .ZN(n1092) );
NOR2_X1 U798 ( .A1(n1094), .A2(n1095), .ZN(n1091) );
XOR2_X1 U799 ( .A(KEYINPUT1), .B(n1096), .Z(n1095) );
AND2_X1 U800 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U801 ( .A1(n1098), .A2(n1097), .ZN(n1094) );
NAND2_X1 U802 ( .A1(G227), .A2(n966), .ZN(n1097) );
XNOR2_X1 U803 ( .A(G140), .B(n1099), .ZN(n1098) );
NAND3_X1 U804 ( .A1(n1062), .A2(G469), .A3(KEYINPUT29), .ZN(n1089) );
NOR2_X1 U805 ( .A1(n1056), .A2(n1100), .ZN(G51) );
XOR2_X1 U806 ( .A(n1101), .B(n1102), .Z(n1100) );
XNOR2_X1 U807 ( .A(n1103), .B(n1104), .ZN(n1102) );
XOR2_X1 U808 ( .A(n1105), .B(n1106), .Z(n1101) );
XNOR2_X1 U809 ( .A(n1107), .B(n1108), .ZN(n1105) );
NAND2_X1 U810 ( .A1(n1062), .A2(G210), .ZN(n1107) );
NOR2_X1 U811 ( .A1(n1109), .A2(n973), .ZN(n1062) );
AND2_X1 U812 ( .A1(n1055), .A2(n1028), .ZN(n973) );
AND4_X1 U813 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1028) );
NOR4_X1 U814 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1113) );
NOR3_X1 U815 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1112) );
NOR2_X1 U816 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
INV_X1 U817 ( .A(KEYINPUT58), .ZN(n1121) );
NOR3_X1 U818 ( .A1(KEYINPUT58), .A2(n985), .A3(n1123), .ZN(n1119) );
AND2_X1 U819 ( .A1(n1124), .A2(n1125), .ZN(n1055) );
NOR4_X1 U820 ( .A1(n1126), .A2(n964), .A3(n1127), .A4(n1128), .ZN(n1125) );
INV_X1 U821 ( .A(n1129), .ZN(n1127) );
AND3_X1 U822 ( .A1(n1130), .A2(n988), .A3(n1131), .ZN(n964) );
AND4_X1 U823 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1073), .ZN(n1124) );
NAND3_X1 U824 ( .A1(n1131), .A2(n988), .A3(n1135), .ZN(n1073) );
NOR2_X1 U825 ( .A1(n966), .A2(G952), .ZN(n1056) );
XNOR2_X1 U826 ( .A(G146), .B(n1111), .ZN(G48) );
NAND2_X1 U827 ( .A1(n1136), .A2(n1135), .ZN(n1111) );
XOR2_X1 U828 ( .A(n1122), .B(n1137), .Z(G45) );
NAND2_X1 U829 ( .A1(KEYINPUT16), .A2(G143), .ZN(n1137) );
OR2_X1 U830 ( .A1(n1123), .A2(n1138), .ZN(n1122) );
NAND4_X1 U831 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1015), .ZN(n1123) );
XOR2_X1 U832 ( .A(n1142), .B(n1117), .Z(G42) );
AND3_X1 U833 ( .A1(n1135), .A2(n986), .A3(n1143), .ZN(n1117) );
XNOR2_X1 U834 ( .A(G140), .B(KEYINPUT51), .ZN(n1142) );
XOR2_X1 U835 ( .A(G137), .B(n1116), .Z(G39) );
AND4_X1 U836 ( .A1(n1143), .A2(n980), .A3(n1144), .A4(n1145), .ZN(n1116) );
XNOR2_X1 U837 ( .A(n1040), .B(n1115), .ZN(G36) );
AND3_X1 U838 ( .A1(n985), .A2(n1130), .A3(n1143), .ZN(n1115) );
XNOR2_X1 U839 ( .A(n1118), .B(n1146), .ZN(G33) );
NAND2_X1 U840 ( .A1(n1147), .A2(KEYINPUT56), .ZN(n1146) );
XNOR2_X1 U841 ( .A(G131), .B(KEYINPUT5), .ZN(n1147) );
AND3_X1 U842 ( .A1(n1135), .A2(n985), .A3(n1143), .ZN(n1118) );
AND3_X1 U843 ( .A1(n983), .A2(n1148), .A3(n1141), .ZN(n1143) );
NAND2_X1 U844 ( .A1(n1149), .A2(n1150), .ZN(n983) );
NAND2_X1 U845 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
INV_X1 U846 ( .A(KEYINPUT22), .ZN(n1152) );
NAND3_X1 U847 ( .A1(n990), .A2(n1153), .A3(KEYINPUT22), .ZN(n1149) );
XOR2_X1 U848 ( .A(n1110), .B(n1154), .Z(G30) );
NAND2_X1 U849 ( .A1(KEYINPUT25), .A2(G128), .ZN(n1154) );
NAND2_X1 U850 ( .A1(n1136), .A2(n1130), .ZN(n1110) );
AND4_X1 U851 ( .A1(n1144), .A2(n1140), .A3(n1141), .A4(n1145), .ZN(n1136) );
XOR2_X1 U852 ( .A(n1134), .B(n1155), .Z(G3) );
XOR2_X1 U853 ( .A(KEYINPUT24), .B(G101), .Z(n1155) );
NAND2_X1 U854 ( .A1(n1156), .A2(n985), .ZN(n1134) );
XOR2_X1 U855 ( .A(G125), .B(n1114), .Z(G27) );
AND4_X1 U856 ( .A1(n1140), .A2(n1135), .A3(n986), .A4(n978), .ZN(n1114) );
AND2_X1 U857 ( .A1(n1151), .A2(n1148), .ZN(n1140) );
NAND2_X1 U858 ( .A1(n1004), .A2(n1157), .ZN(n1148) );
NAND4_X1 U859 ( .A1(G902), .A2(G953), .A3(n1158), .A4(n1032), .ZN(n1157) );
INV_X1 U860 ( .A(G900), .ZN(n1032) );
XNOR2_X1 U861 ( .A(G122), .B(n1133), .ZN(G24) );
NAND4_X1 U862 ( .A1(n1159), .A2(n988), .A3(n1139), .A4(n1015), .ZN(n1133) );
NOR2_X1 U863 ( .A1(n1145), .A2(n1144), .ZN(n988) );
NAND2_X1 U864 ( .A1(n1160), .A2(n1161), .ZN(G21) );
NAND2_X1 U865 ( .A1(G119), .A2(n1132), .ZN(n1161) );
XOR2_X1 U866 ( .A(KEYINPUT48), .B(n1162), .Z(n1160) );
NOR2_X1 U867 ( .A1(G119), .A2(n1132), .ZN(n1162) );
NAND4_X1 U868 ( .A1(n980), .A2(n1159), .A3(n1144), .A4(n1145), .ZN(n1132) );
XOR2_X1 U869 ( .A(G116), .B(n1126), .Z(G18) );
AND3_X1 U870 ( .A1(n985), .A2(n1130), .A3(n1159), .ZN(n1126) );
INV_X1 U871 ( .A(n997), .ZN(n1130) );
NAND2_X1 U872 ( .A1(n1163), .A2(n1139), .ZN(n997) );
XOR2_X1 U873 ( .A(n1164), .B(KEYINPUT8), .Z(n1139) );
XNOR2_X1 U874 ( .A(n1128), .B(n1165), .ZN(G15) );
NAND2_X1 U875 ( .A1(KEYINPUT15), .A2(G113), .ZN(n1165) );
AND3_X1 U876 ( .A1(n1159), .A2(n985), .A3(n1135), .ZN(n1128) );
INV_X1 U877 ( .A(n996), .ZN(n1135) );
NAND2_X1 U878 ( .A1(n1164), .A2(n1015), .ZN(n996) );
INV_X1 U879 ( .A(n1138), .ZN(n985) );
NAND2_X1 U880 ( .A1(n1144), .A2(n1166), .ZN(n1138) );
XNOR2_X1 U881 ( .A(KEYINPUT45), .B(n1145), .ZN(n1166) );
AND3_X1 U882 ( .A1(n1151), .A2(n1167), .A3(n978), .ZN(n1159) );
NOR2_X1 U883 ( .A1(n1003), .A2(n1001), .ZN(n978) );
XNOR2_X1 U884 ( .A(G110), .B(n1129), .ZN(G12) );
NAND2_X1 U885 ( .A1(n986), .A2(n1156), .ZN(n1129) );
AND2_X1 U886 ( .A1(n980), .A2(n1131), .ZN(n1156) );
AND3_X1 U887 ( .A1(n1141), .A2(n1167), .A3(n1151), .ZN(n1131) );
NOR2_X1 U888 ( .A1(n991), .A2(n990), .ZN(n1151) );
AND2_X1 U889 ( .A1(n1168), .A2(n1014), .ZN(n990) );
NAND2_X1 U890 ( .A1(n1169), .A2(n1170), .ZN(n1014) );
NAND2_X1 U891 ( .A1(G210), .A2(n1171), .ZN(n1170) );
INV_X1 U892 ( .A(n1172), .ZN(n1169) );
XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n1013), .ZN(n1168) );
NAND3_X1 U894 ( .A1(n1172), .A2(n1171), .A3(G210), .ZN(n1013) );
NAND2_X1 U895 ( .A1(n1173), .A2(n1109), .ZN(n1172) );
XOR2_X1 U896 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U897 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U898 ( .A1(KEYINPUT50), .A2(n1103), .ZN(n1177) );
XOR2_X1 U899 ( .A(n1052), .B(n1178), .Z(n1103) );
XNOR2_X1 U900 ( .A(n1099), .B(n1179), .ZN(n1178) );
XOR2_X1 U901 ( .A(n1180), .B(n1181), .Z(n1052) );
XOR2_X1 U902 ( .A(G119), .B(G101), .Z(n1181) );
XOR2_X1 U903 ( .A(n1182), .B(n1183), .Z(n1180) );
NAND2_X1 U904 ( .A1(KEYINPUT28), .A2(n1075), .ZN(n1182) );
NAND2_X1 U905 ( .A1(n1184), .A2(n1185), .ZN(n1176) );
NAND2_X1 U906 ( .A1(n1106), .A2(n1104), .ZN(n1185) );
INV_X1 U907 ( .A(n1186), .ZN(n1104) );
NAND2_X1 U908 ( .A1(n1187), .A2(n1186), .ZN(n1184) );
XOR2_X1 U909 ( .A(G128), .B(n1188), .Z(n1186) );
XOR2_X1 U910 ( .A(KEYINPUT63), .B(n1106), .Z(n1187) );
XOR2_X1 U911 ( .A(G125), .B(KEYINPUT13), .Z(n1106) );
XOR2_X1 U912 ( .A(n1108), .B(KEYINPUT61), .Z(n1174) );
NAND2_X1 U913 ( .A1(n1189), .A2(G224), .ZN(n1108) );
XNOR2_X1 U914 ( .A(G953), .B(KEYINPUT26), .ZN(n1189) );
INV_X1 U915 ( .A(n1153), .ZN(n991) );
NAND2_X1 U916 ( .A1(G214), .A2(n1171), .ZN(n1153) );
NAND2_X1 U917 ( .A1(n1190), .A2(n1109), .ZN(n1171) );
XNOR2_X1 U918 ( .A(G237), .B(KEYINPUT47), .ZN(n1190) );
NAND2_X1 U919 ( .A1(n1004), .A2(n1191), .ZN(n1167) );
NAND4_X1 U920 ( .A1(G902), .A2(G953), .A3(n1158), .A4(n1049), .ZN(n1191) );
INV_X1 U921 ( .A(G898), .ZN(n1049) );
NAND3_X1 U922 ( .A1(n1158), .A2(n966), .A3(G952), .ZN(n1004) );
INV_X1 U923 ( .A(G953), .ZN(n966) );
NAND2_X1 U924 ( .A1(G234), .A2(G237), .ZN(n1158) );
INV_X1 U925 ( .A(n999), .ZN(n1141) );
NAND2_X1 U926 ( .A1(n1192), .A2(n1003), .ZN(n999) );
XNOR2_X1 U927 ( .A(n1011), .B(G469), .ZN(n1003) );
NAND2_X1 U928 ( .A1(n1193), .A2(n1109), .ZN(n1011) );
XOR2_X1 U929 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U930 ( .A(n1093), .B(n1196), .Z(n1195) );
XOR2_X1 U931 ( .A(n1197), .B(n1198), .Z(n1196) );
NOR2_X1 U932 ( .A1(G140), .A2(n1199), .ZN(n1198) );
XOR2_X1 U933 ( .A(KEYINPUT2), .B(KEYINPUT19), .Z(n1199) );
NAND2_X1 U934 ( .A1(KEYINPUT12), .A2(G227), .ZN(n1197) );
XOR2_X1 U935 ( .A(n1200), .B(n1201), .Z(n1093) );
XNOR2_X1 U936 ( .A(n1202), .B(n1039), .ZN(n1200) );
NAND2_X1 U937 ( .A1(KEYINPUT6), .A2(n1203), .ZN(n1039) );
XNOR2_X1 U938 ( .A(G146), .B(n1204), .ZN(n1203) );
NAND2_X1 U939 ( .A1(KEYINPUT46), .A2(n1205), .ZN(n1204) );
NAND2_X1 U940 ( .A1(n1206), .A2(n1207), .ZN(n1202) );
NAND2_X1 U941 ( .A1(G101), .A2(n1208), .ZN(n1207) );
XOR2_X1 U942 ( .A(KEYINPUT34), .B(n1209), .Z(n1206) );
NOR2_X1 U943 ( .A1(G101), .A2(n1208), .ZN(n1209) );
XNOR2_X1 U944 ( .A(G107), .B(n1075), .ZN(n1208) );
XNOR2_X1 U945 ( .A(G110), .B(n1210), .ZN(n1194) );
XNOR2_X1 U946 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n1210) );
XNOR2_X1 U947 ( .A(n1001), .B(KEYINPUT9), .ZN(n1192) );
INV_X1 U948 ( .A(n1012), .ZN(n1001) );
NAND2_X1 U949 ( .A1(G221), .A2(n1211), .ZN(n1012) );
NAND2_X1 U950 ( .A1(G234), .A2(n1109), .ZN(n1211) );
AND2_X1 U951 ( .A1(n1163), .A2(n1164), .ZN(n980) );
XNOR2_X1 U952 ( .A(n1020), .B(n1212), .ZN(n1164) );
NOR2_X1 U953 ( .A1(KEYINPUT35), .A2(n1069), .ZN(n1212) );
INV_X1 U954 ( .A(G478), .ZN(n1069) );
NOR2_X1 U955 ( .A1(n1067), .A2(G902), .ZN(n1020) );
XNOR2_X1 U956 ( .A(n1213), .B(n1214), .ZN(n1067) );
XOR2_X1 U957 ( .A(G122), .B(n1215), .Z(n1214) );
XNOR2_X1 U958 ( .A(KEYINPUT52), .B(n1040), .ZN(n1215) );
XNOR2_X1 U959 ( .A(n1183), .B(n1216), .ZN(n1213) );
XNOR2_X1 U960 ( .A(n1217), .B(n1218), .ZN(n1216) );
AND3_X1 U961 ( .A1(G217), .A2(n1219), .A3(n1220), .ZN(n1218) );
INV_X1 U962 ( .A(KEYINPUT23), .ZN(n1219) );
NAND2_X1 U963 ( .A1(n1221), .A2(KEYINPUT60), .ZN(n1217) );
XNOR2_X1 U964 ( .A(G128), .B(n1222), .ZN(n1221) );
NOR2_X1 U965 ( .A1(KEYINPUT38), .A2(n1223), .ZN(n1222) );
XNOR2_X1 U966 ( .A(G143), .B(KEYINPUT33), .ZN(n1223) );
XOR2_X1 U967 ( .A(G116), .B(G107), .Z(n1183) );
INV_X1 U968 ( .A(n1015), .ZN(n1163) );
XNOR2_X1 U969 ( .A(n1224), .B(G475), .ZN(n1015) );
NAND2_X1 U970 ( .A1(n1072), .A2(n1109), .ZN(n1224) );
XOR2_X1 U971 ( .A(n1225), .B(n1226), .Z(n1072) );
XOR2_X1 U972 ( .A(n1227), .B(n1228), .Z(n1226) );
XNOR2_X1 U973 ( .A(n1229), .B(n1075), .ZN(n1228) );
INV_X1 U974 ( .A(G104), .ZN(n1075) );
NAND2_X1 U975 ( .A1(KEYINPUT53), .A2(n1230), .ZN(n1229) );
INV_X1 U976 ( .A(G131), .ZN(n1230) );
NAND2_X1 U977 ( .A1(n1231), .A2(G214), .ZN(n1227) );
XNOR2_X1 U978 ( .A(n1179), .B(n1232), .ZN(n1225) );
XNOR2_X1 U979 ( .A(n1233), .B(n1234), .ZN(n1232) );
XOR2_X1 U980 ( .A(G113), .B(G122), .Z(n1179) );
NOR2_X1 U981 ( .A1(n1144), .A2(n1006), .ZN(n986) );
INV_X1 U982 ( .A(n1145), .ZN(n1006) );
NAND3_X1 U983 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1145) );
NAND2_X1 U984 ( .A1(G217), .A2(G902), .ZN(n1237) );
NAND3_X1 U985 ( .A1(n1061), .A2(n1109), .A3(n1238), .ZN(n1236) );
OR2_X1 U986 ( .A1(n1238), .A2(n1061), .ZN(n1235) );
XNOR2_X1 U987 ( .A(n1239), .B(n1240), .ZN(n1061) );
XNOR2_X1 U988 ( .A(n1099), .B(n1241), .ZN(n1240) );
XNOR2_X1 U989 ( .A(n1242), .B(G119), .ZN(n1241) );
INV_X1 U990 ( .A(G110), .ZN(n1099) );
XOR2_X1 U991 ( .A(n1243), .B(n1234), .Z(n1239) );
XOR2_X1 U992 ( .A(G125), .B(G140), .Z(n1234) );
XOR2_X1 U993 ( .A(n1244), .B(n1245), .Z(n1243) );
NAND2_X1 U994 ( .A1(n1220), .A2(G221), .ZN(n1244) );
NOR2_X1 U995 ( .A1(n1246), .A2(G953), .ZN(n1220) );
NAND2_X1 U996 ( .A1(G217), .A2(n1246), .ZN(n1238) );
INV_X1 U997 ( .A(G234), .ZN(n1246) );
XOR2_X1 U998 ( .A(n1247), .B(G472), .Z(n1144) );
NAND2_X1 U999 ( .A1(KEYINPUT10), .A2(n1022), .ZN(n1247) );
NAND4_X1 U1000 ( .A1(n1248), .A2(n1109), .A3(n1249), .A4(n1250), .ZN(n1022) );
NAND3_X1 U1001 ( .A1(KEYINPUT59), .A2(n1251), .A3(n1080), .ZN(n1250) );
OR2_X1 U1002 ( .A1(n1080), .A2(n1251), .ZN(n1249) );
NOR2_X1 U1003 ( .A1(KEYINPUT14), .A2(n1252), .ZN(n1251) );
XNOR2_X1 U1004 ( .A(n1253), .B(G101), .ZN(n1080) );
NAND2_X1 U1005 ( .A1(n1231), .A2(G210), .ZN(n1253) );
NOR2_X1 U1006 ( .A1(G953), .A2(G237), .ZN(n1231) );
INV_X1 U1007 ( .A(G902), .ZN(n1109) );
NAND2_X1 U1008 ( .A1(n1252), .A2(n1254), .ZN(n1248) );
INV_X1 U1009 ( .A(KEYINPUT59), .ZN(n1254) );
XNOR2_X1 U1010 ( .A(n1255), .B(n1086), .ZN(n1252) );
XOR2_X1 U1011 ( .A(n1201), .B(n1188), .Z(n1086) );
XNOR2_X1 U1012 ( .A(n1233), .B(KEYINPUT18), .ZN(n1188) );
XNOR2_X1 U1013 ( .A(n1205), .B(n1242), .ZN(n1233) );
INV_X1 U1014 ( .A(G146), .ZN(n1242) );
INV_X1 U1015 ( .A(G143), .ZN(n1205) );
XOR2_X1 U1016 ( .A(n1036), .B(n1040), .Z(n1201) );
INV_X1 U1017 ( .A(G134), .ZN(n1040) );
XNOR2_X1 U1018 ( .A(G131), .B(n1245), .ZN(n1036) );
XOR2_X1 U1019 ( .A(G137), .B(G128), .Z(n1245) );
NAND2_X1 U1020 ( .A1(n1256), .A2(n1084), .ZN(n1255) );
XOR2_X1 U1021 ( .A(G113), .B(n1257), .Z(n1084) );
XOR2_X1 U1022 ( .A(G119), .B(G116), .Z(n1257) );
XOR2_X1 U1023 ( .A(KEYINPUT7), .B(KEYINPUT31), .Z(n1256) );
endmodule


