//Key = 0011011111001100111101110011101010001001110110111110101100001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295;

XNOR2_X1 U716 ( .A(G107), .B(n985), .ZN(G9) );
NAND2_X1 U717 ( .A1(KEYINPUT50), .A2(n986), .ZN(n985) );
NOR2_X1 U718 ( .A1(n987), .A2(n988), .ZN(G75) );
NOR4_X1 U719 ( .A1(G953), .A2(n989), .A3(n990), .A4(n991), .ZN(n988) );
NOR2_X1 U720 ( .A1(n992), .A2(n993), .ZN(n990) );
NOR2_X1 U721 ( .A1(n994), .A2(n995), .ZN(n992) );
NOR3_X1 U722 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n995) );
NOR2_X1 U723 ( .A1(n999), .A2(n1000), .ZN(n997) );
NOR2_X1 U724 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
NOR2_X1 U725 ( .A1(n1003), .A2(n1004), .ZN(n999) );
NOR2_X1 U726 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
NOR2_X1 U727 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NOR2_X1 U728 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NOR3_X1 U729 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1009) );
NOR2_X1 U730 ( .A1(n1014), .A2(n1002), .ZN(n1005) );
NOR2_X1 U731 ( .A1(n1007), .A2(n1012), .ZN(n1014) );
INV_X1 U732 ( .A(KEYINPUT36), .ZN(n1012) );
NOR4_X1 U733 ( .A1(n1007), .A2(n1015), .A3(n1002), .A4(n1004), .ZN(n994) );
INV_X1 U734 ( .A(n1016), .ZN(n1002) );
NOR2_X1 U735 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NOR2_X1 U736 ( .A1(n1019), .A2(n996), .ZN(n1018) );
NOR2_X1 U737 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NOR2_X1 U738 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U739 ( .A1(n1024), .A2(n998), .ZN(n1017) );
NOR2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NOR3_X1 U741 ( .A1(n989), .A2(G953), .A3(G952), .ZN(n987) );
AND4_X1 U742 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n989) );
NOR3_X1 U743 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
NOR2_X1 U744 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR2_X1 U745 ( .A1(n1036), .A2(n1037), .ZN(n1032) );
INV_X1 U746 ( .A(n1038), .ZN(n1037) );
XOR2_X1 U747 ( .A(n1039), .B(KEYINPUT55), .Z(n1036) );
NAND3_X1 U748 ( .A1(n1040), .A2(n1011), .A3(n1041), .ZN(n1031) );
NOR3_X1 U749 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1029) );
XOR2_X1 U750 ( .A(n1045), .B(n1046), .Z(n1044) );
XOR2_X1 U751 ( .A(KEYINPUT60), .B(G475), .Z(n1046) );
XOR2_X1 U752 ( .A(n1047), .B(KEYINPUT52), .Z(n1043) );
NAND2_X1 U753 ( .A1(n1035), .A2(n1034), .ZN(n1047) );
XNOR2_X1 U754 ( .A(KEYINPUT31), .B(n1048), .ZN(n1035) );
XNOR2_X1 U755 ( .A(n1013), .B(KEYINPUT8), .ZN(n1042) );
XOR2_X1 U756 ( .A(n1049), .B(KEYINPUT10), .Z(n1027) );
XOR2_X1 U757 ( .A(n1050), .B(n1051), .Z(G72) );
XOR2_X1 U758 ( .A(n1052), .B(n1053), .Z(n1051) );
NAND2_X1 U759 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U760 ( .A1(G953), .A2(n1056), .ZN(n1055) );
XNOR2_X1 U761 ( .A(n1057), .B(n1058), .ZN(n1054) );
NOR2_X1 U762 ( .A1(KEYINPUT38), .A2(n1059), .ZN(n1058) );
XOR2_X1 U763 ( .A(n1060), .B(n1061), .Z(n1059) );
XOR2_X1 U764 ( .A(KEYINPUT30), .B(n1062), .Z(n1061) );
XOR2_X1 U765 ( .A(n1063), .B(n1064), .Z(n1060) );
NAND2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1052) );
NAND2_X1 U767 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XOR2_X1 U768 ( .A(KEYINPUT48), .B(n1069), .Z(n1068) );
NOR2_X1 U769 ( .A1(n1070), .A2(n1065), .ZN(n1050) );
NOR2_X1 U770 ( .A1(n1071), .A2(n1056), .ZN(n1070) );
XOR2_X1 U771 ( .A(n1072), .B(n1073), .Z(G69) );
XOR2_X1 U772 ( .A(n1074), .B(n1075), .Z(n1073) );
NAND2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
INV_X1 U774 ( .A(n1078), .ZN(n1077) );
XNOR2_X1 U775 ( .A(n1079), .B(n1080), .ZN(n1076) );
NOR2_X1 U776 ( .A1(KEYINPUT34), .A2(n1081), .ZN(n1080) );
NAND2_X1 U777 ( .A1(n1082), .A2(n1065), .ZN(n1074) );
NAND4_X1 U778 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1082) );
XOR2_X1 U779 ( .A(KEYINPUT2), .B(n986), .Z(n1085) );
XOR2_X1 U780 ( .A(n1087), .B(KEYINPUT53), .Z(n1083) );
NOR2_X1 U781 ( .A1(n1088), .A2(n1065), .ZN(n1072) );
AND2_X1 U782 ( .A1(G224), .A2(G898), .ZN(n1088) );
NOR2_X1 U783 ( .A1(n1089), .A2(n1090), .ZN(G66) );
XOR2_X1 U784 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U785 ( .A1(n1039), .A2(n1093), .ZN(n1091) );
NOR2_X1 U786 ( .A1(n1089), .A2(n1094), .ZN(G63) );
XOR2_X1 U787 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U788 ( .A1(n1097), .A2(n1093), .ZN(n1095) );
XNOR2_X1 U789 ( .A(G478), .B(KEYINPUT57), .ZN(n1097) );
NOR2_X1 U790 ( .A1(n1089), .A2(n1098), .ZN(G60) );
NOR3_X1 U791 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
NOR3_X1 U792 ( .A1(n1102), .A2(n1103), .A3(n1093), .ZN(n1101) );
NOR2_X1 U793 ( .A1(n1104), .A2(n1105), .ZN(n1100) );
AND2_X1 U794 ( .A1(n991), .A2(G475), .ZN(n1104) );
XOR2_X1 U795 ( .A(G104), .B(n1106), .Z(G6) );
NOR4_X1 U796 ( .A1(KEYINPUT61), .A2(n998), .A3(n1107), .A4(n1108), .ZN(n1106) );
NOR2_X1 U797 ( .A1(n1089), .A2(n1109), .ZN(G57) );
XOR2_X1 U798 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U799 ( .A(G101), .B(n1112), .Z(n1111) );
NOR2_X1 U800 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
INV_X1 U801 ( .A(n1115), .ZN(n1113) );
XOR2_X1 U802 ( .A(n1116), .B(n1117), .Z(n1110) );
NOR2_X1 U803 ( .A1(n1034), .A2(n1093), .ZN(n1117) );
INV_X1 U804 ( .A(G472), .ZN(n1034) );
NAND2_X1 U805 ( .A1(KEYINPUT12), .A2(n1118), .ZN(n1116) );
NOR2_X1 U806 ( .A1(n1089), .A2(n1119), .ZN(G54) );
XOR2_X1 U807 ( .A(n1120), .B(n1121), .Z(n1119) );
XOR2_X1 U808 ( .A(n1122), .B(n1123), .Z(n1121) );
NAND3_X1 U809 ( .A1(n1124), .A2(n1125), .A3(KEYINPUT54), .ZN(n1122) );
XOR2_X1 U810 ( .A(KEYINPUT20), .B(G469), .Z(n1125) );
INV_X1 U811 ( .A(n1093), .ZN(n1124) );
XOR2_X1 U812 ( .A(KEYINPUT27), .B(n1126), .Z(n1120) );
NOR2_X1 U813 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U814 ( .A(n1129), .B(KEYINPUT39), .Z(n1128) );
NAND2_X1 U815 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U816 ( .A1(n1131), .A2(n1130), .ZN(n1127) );
XOR2_X1 U817 ( .A(n1132), .B(G140), .Z(n1130) );
NAND2_X1 U818 ( .A1(KEYINPUT21), .A2(G110), .ZN(n1132) );
NOR2_X1 U819 ( .A1(n1089), .A2(n1133), .ZN(G51) );
XOR2_X1 U820 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U821 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U822 ( .A1(KEYINPUT43), .A2(n1138), .ZN(n1136) );
XOR2_X1 U823 ( .A(n1139), .B(n1140), .Z(n1134) );
NOR2_X1 U824 ( .A1(n1141), .A2(n1093), .ZN(n1140) );
NAND2_X1 U825 ( .A1(G902), .A2(n991), .ZN(n1093) );
NAND4_X1 U826 ( .A1(n1067), .A2(n1084), .A3(n1142), .A4(n1143), .ZN(n991) );
NOR3_X1 U827 ( .A1(n1144), .A2(n1069), .A3(n986), .ZN(n1143) );
AND3_X1 U828 ( .A1(n1025), .A2(n1145), .A3(n1146), .ZN(n986) );
XOR2_X1 U829 ( .A(n1086), .B(KEYINPUT45), .Z(n1142) );
NAND4_X1 U830 ( .A1(n1147), .A2(n1026), .A3(n1148), .A4(n1145), .ZN(n1086) );
NOR2_X1 U831 ( .A1(n1149), .A2(n1001), .ZN(n1148) );
XOR2_X1 U832 ( .A(n1150), .B(KEYINPUT32), .Z(n1147) );
AND4_X1 U833 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1084) );
NOR2_X1 U834 ( .A1(n1155), .A2(n1156), .ZN(n1153) );
AND4_X1 U835 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1067) );
AND4_X1 U836 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1160) );
XOR2_X1 U837 ( .A(n1165), .B(n1166), .Z(n1139) );
NOR2_X1 U838 ( .A1(n1065), .A2(G952), .ZN(n1089) );
XOR2_X1 U839 ( .A(G146), .B(n1069), .Z(G48) );
AND3_X1 U840 ( .A1(n1167), .A2(n1010), .A3(n1026), .ZN(n1069) );
XOR2_X1 U841 ( .A(n1168), .B(n1169), .Z(G45) );
NAND2_X1 U842 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NAND2_X1 U843 ( .A1(KEYINPUT16), .A2(n1159), .ZN(n1171) );
NAND2_X1 U844 ( .A1(KEYINPUT14), .A2(n1172), .ZN(n1170) );
INV_X1 U845 ( .A(n1159), .ZN(n1172) );
NAND4_X1 U846 ( .A1(n1173), .A2(n1174), .A3(n1010), .A4(n1175), .ZN(n1159) );
XNOR2_X1 U847 ( .A(G140), .B(n1157), .ZN(G42) );
NAND3_X1 U848 ( .A1(n1176), .A2(n1177), .A3(n1016), .ZN(n1157) );
XNOR2_X1 U849 ( .A(G137), .B(n1158), .ZN(G39) );
NAND3_X1 U850 ( .A1(n1016), .A2(n1167), .A3(n1178), .ZN(n1158) );
XNOR2_X1 U851 ( .A(G134), .B(n1164), .ZN(G36) );
NAND3_X1 U852 ( .A1(n1174), .A2(n1025), .A3(n1016), .ZN(n1164) );
XNOR2_X1 U853 ( .A(G131), .B(n1163), .ZN(G33) );
NAND3_X1 U854 ( .A1(n1174), .A2(n1026), .A3(n1016), .ZN(n1163) );
NOR2_X1 U855 ( .A1(n1013), .A2(n1179), .ZN(n1016) );
INV_X1 U856 ( .A(n1011), .ZN(n1179) );
AND3_X1 U857 ( .A1(n1177), .A2(n1180), .A3(n1021), .ZN(n1174) );
XOR2_X1 U858 ( .A(n1162), .B(n1181), .Z(G30) );
NAND2_X1 U859 ( .A1(KEYINPUT9), .A2(G128), .ZN(n1181) );
NAND3_X1 U860 ( .A1(n1025), .A2(n1010), .A3(n1167), .ZN(n1162) );
AND4_X1 U861 ( .A1(n1177), .A2(n1023), .A3(n1180), .A4(n1182), .ZN(n1167) );
INV_X1 U862 ( .A(n1001), .ZN(n1177) );
XNOR2_X1 U863 ( .A(G101), .B(n1151), .ZN(G3) );
NAND3_X1 U864 ( .A1(n1021), .A2(n1146), .A3(n1178), .ZN(n1151) );
XOR2_X1 U865 ( .A(n1165), .B(n1161), .Z(G27) );
NAND4_X1 U866 ( .A1(n1049), .A2(n1176), .A3(n1010), .A4(n1041), .ZN(n1161) );
INV_X1 U867 ( .A(n1150), .ZN(n1010) );
AND4_X1 U868 ( .A1(n1183), .A2(n1026), .A3(n1180), .A4(n1182), .ZN(n1176) );
NAND2_X1 U869 ( .A1(n993), .A2(n1184), .ZN(n1180) );
NAND4_X1 U870 ( .A1(G902), .A2(G953), .A3(n1185), .A4(n1056), .ZN(n1184) );
INV_X1 U871 ( .A(G900), .ZN(n1056) );
XOR2_X1 U872 ( .A(n1186), .B(n1152), .Z(G24) );
NAND4_X1 U873 ( .A1(n1173), .A2(n1187), .A3(n1145), .A4(n1175), .ZN(n1152) );
INV_X1 U874 ( .A(n998), .ZN(n1145) );
NAND2_X1 U875 ( .A1(n1022), .A2(n1183), .ZN(n998) );
XNOR2_X1 U876 ( .A(G119), .B(n1154), .ZN(G21) );
NAND4_X1 U877 ( .A1(n1187), .A2(n1178), .A3(n1023), .A4(n1182), .ZN(n1154) );
XOR2_X1 U878 ( .A(G116), .B(n1144), .Z(G18) );
INV_X1 U879 ( .A(n1087), .ZN(n1144) );
NAND3_X1 U880 ( .A1(n1021), .A2(n1025), .A3(n1187), .ZN(n1087) );
NOR2_X1 U881 ( .A1(n1028), .A2(n1173), .ZN(n1025) );
XOR2_X1 U882 ( .A(G113), .B(n1156), .Z(G15) );
AND3_X1 U883 ( .A1(n1021), .A2(n1026), .A3(n1187), .ZN(n1156) );
NOR4_X1 U884 ( .A1(n1004), .A2(n1150), .A3(n1149), .A4(n1007), .ZN(n1187) );
INV_X1 U885 ( .A(n1041), .ZN(n1007) );
INV_X1 U886 ( .A(n1108), .ZN(n1026) );
NAND2_X1 U887 ( .A1(n1173), .A2(n1028), .ZN(n1108) );
NOR2_X1 U888 ( .A1(n1182), .A2(n1183), .ZN(n1021) );
XOR2_X1 U889 ( .A(n1155), .B(n1188), .Z(G12) );
NOR2_X1 U890 ( .A1(KEYINPUT29), .A2(n1189), .ZN(n1188) );
NOR4_X1 U891 ( .A1(n996), .A2(n1107), .A3(n1023), .A4(n1022), .ZN(n1155) );
INV_X1 U892 ( .A(n1182), .ZN(n1022) );
NAND2_X1 U893 ( .A1(n1190), .A2(n1040), .ZN(n1182) );
OR2_X1 U894 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
NAND2_X1 U895 ( .A1(n1038), .A2(n1039), .ZN(n1190) );
NAND2_X1 U896 ( .A1(G217), .A2(n1191), .ZN(n1039) );
NOR2_X1 U897 ( .A1(n1092), .A2(G902), .ZN(n1038) );
XNOR2_X1 U898 ( .A(n1192), .B(n1193), .ZN(n1092) );
XNOR2_X1 U899 ( .A(n1057), .B(n1194), .ZN(n1193) );
XOR2_X1 U900 ( .A(n1195), .B(n1196), .Z(n1194) );
NOR2_X1 U901 ( .A1(KEYINPUT63), .A2(G146), .ZN(n1196) );
NAND2_X1 U902 ( .A1(n1197), .A2(G221), .ZN(n1195) );
XOR2_X1 U903 ( .A(n1198), .B(n1199), .Z(n1192) );
NOR2_X1 U904 ( .A1(KEYINPUT4), .A2(n1200), .ZN(n1199) );
XOR2_X1 U905 ( .A(n1201), .B(n1202), .Z(n1200) );
XOR2_X1 U906 ( .A(G128), .B(G110), .Z(n1202) );
XNOR2_X1 U907 ( .A(G137), .B(KEYINPUT56), .ZN(n1198) );
INV_X1 U908 ( .A(n1183), .ZN(n1023) );
XOR2_X1 U909 ( .A(n1048), .B(G472), .Z(n1183) );
NAND3_X1 U910 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1048) );
NAND3_X1 U911 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1204) );
INV_X1 U912 ( .A(KEYINPUT23), .ZN(n1208) );
NAND2_X1 U913 ( .A1(n1209), .A2(KEYINPUT23), .ZN(n1203) );
XOR2_X1 U914 ( .A(n1207), .B(n1206), .Z(n1209) );
XOR2_X1 U915 ( .A(n1210), .B(KEYINPUT1), .Z(n1206) );
NAND3_X1 U916 ( .A1(n1211), .A2(n1212), .A3(n1115), .ZN(n1210) );
NAND3_X1 U917 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1115) );
NAND2_X1 U918 ( .A1(n1216), .A2(n1217), .ZN(n1212) );
INV_X1 U919 ( .A(KEYINPUT41), .ZN(n1217) );
XOR2_X1 U920 ( .A(n1215), .B(n1218), .Z(n1216) );
NOR2_X1 U921 ( .A1(n1214), .A2(n1213), .ZN(n1218) );
NAND2_X1 U922 ( .A1(KEYINPUT41), .A2(n1114), .ZN(n1211) );
NAND2_X1 U923 ( .A1(n1219), .A2(n1220), .ZN(n1114) );
NAND3_X1 U924 ( .A1(n1221), .A2(n1138), .A3(n1214), .ZN(n1220) );
INV_X1 U925 ( .A(n1215), .ZN(n1221) );
NAND2_X1 U926 ( .A1(n1222), .A2(n1223), .ZN(n1219) );
INV_X1 U927 ( .A(n1214), .ZN(n1223) );
XOR2_X1 U928 ( .A(n1213), .B(n1215), .Z(n1222) );
XOR2_X1 U929 ( .A(n1224), .B(KEYINPUT15), .Z(n1215) );
XNOR2_X1 U930 ( .A(n1118), .B(n1225), .ZN(n1207) );
XOR2_X1 U931 ( .A(KEYINPUT47), .B(G101), .Z(n1225) );
AND3_X1 U932 ( .A1(n1226), .A2(n1065), .A3(n1227), .ZN(n1118) );
XOR2_X1 U933 ( .A(n1141), .B(KEYINPUT26), .Z(n1227) );
INV_X1 U934 ( .A(G210), .ZN(n1141) );
INV_X1 U935 ( .A(n1146), .ZN(n1107) );
NOR3_X1 U936 ( .A1(n1150), .A2(n1149), .A3(n1001), .ZN(n1146) );
NAND2_X1 U937 ( .A1(n1004), .A2(n1041), .ZN(n1001) );
NAND2_X1 U938 ( .A1(G221), .A2(n1191), .ZN(n1041) );
NAND2_X1 U939 ( .A1(n1228), .A2(n1205), .ZN(n1191) );
XOR2_X1 U940 ( .A(KEYINPUT37), .B(G234), .Z(n1228) );
INV_X1 U941 ( .A(n1049), .ZN(n1004) );
XOR2_X1 U942 ( .A(n1229), .B(G469), .Z(n1049) );
NAND2_X1 U943 ( .A1(n1230), .A2(n1205), .ZN(n1229) );
XOR2_X1 U944 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U945 ( .A(n1123), .B(n1131), .Z(n1232) );
NOR2_X1 U946 ( .A1(n1071), .A2(G953), .ZN(n1131) );
INV_X1 U947 ( .A(G227), .ZN(n1071) );
XOR2_X1 U948 ( .A(n1233), .B(n1234), .Z(n1123) );
XOR2_X1 U949 ( .A(n1214), .B(n1235), .Z(n1234) );
XNOR2_X1 U950 ( .A(KEYINPUT19), .B(n1236), .ZN(n1235) );
NOR2_X1 U951 ( .A1(KEYINPUT62), .A2(n1237), .ZN(n1236) );
XOR2_X1 U952 ( .A(n1238), .B(n1239), .Z(n1214) );
NOR2_X1 U953 ( .A1(KEYINPUT35), .A2(n1064), .ZN(n1239) );
XOR2_X1 U954 ( .A(G134), .B(G137), .Z(n1064) );
XOR2_X1 U955 ( .A(n1063), .B(n1240), .Z(n1233) );
XOR2_X1 U956 ( .A(n1241), .B(KEYINPUT17), .Z(n1063) );
NAND2_X1 U957 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
OR2_X1 U958 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XOR2_X1 U959 ( .A(n1246), .B(KEYINPUT58), .Z(n1242) );
NAND2_X1 U960 ( .A1(n1245), .A2(n1244), .ZN(n1246) );
INV_X1 U961 ( .A(G128), .ZN(n1244) );
XNOR2_X1 U962 ( .A(n1247), .B(G146), .ZN(n1245) );
NAND2_X1 U963 ( .A1(KEYINPUT22), .A2(n1168), .ZN(n1247) );
INV_X1 U964 ( .A(G143), .ZN(n1168) );
XOR2_X1 U965 ( .A(n1189), .B(n1248), .Z(n1231) );
XOR2_X1 U966 ( .A(KEYINPUT3), .B(G140), .Z(n1248) );
AND2_X1 U967 ( .A1(n993), .A2(n1249), .ZN(n1149) );
NAND3_X1 U968 ( .A1(n1078), .A2(n1185), .A3(G902), .ZN(n1249) );
NOR2_X1 U969 ( .A1(n1065), .A2(G898), .ZN(n1078) );
NAND3_X1 U970 ( .A1(n1185), .A2(n1065), .A3(G952), .ZN(n993) );
NAND2_X1 U971 ( .A1(G237), .A2(G234), .ZN(n1185) );
NAND2_X1 U972 ( .A1(n1013), .A2(n1011), .ZN(n1150) );
NAND2_X1 U973 ( .A1(G214), .A2(n1250), .ZN(n1011) );
XNOR2_X1 U974 ( .A(n1251), .B(n1252), .ZN(n1013) );
NOR2_X1 U975 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
XOR2_X1 U976 ( .A(KEYINPUT7), .B(G210), .Z(n1254) );
INV_X1 U977 ( .A(n1250), .ZN(n1253) );
NAND2_X1 U978 ( .A1(n1205), .A2(n1226), .ZN(n1250) );
NAND3_X1 U979 ( .A1(n1255), .A2(n1256), .A3(n1205), .ZN(n1251) );
NAND2_X1 U980 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XOR2_X1 U981 ( .A(KEYINPUT24), .B(n1259), .Z(n1257) );
NAND2_X1 U982 ( .A1(n1260), .A2(n1261), .ZN(n1255) );
INV_X1 U983 ( .A(n1258), .ZN(n1261) );
XOR2_X1 U984 ( .A(n1262), .B(n1138), .Z(n1258) );
INV_X1 U985 ( .A(n1213), .ZN(n1138) );
XOR2_X1 U986 ( .A(n1263), .B(n1264), .Z(n1213) );
NOR2_X1 U987 ( .A1(KEYINPUT33), .A2(G143), .ZN(n1264) );
XOR2_X1 U988 ( .A(n1265), .B(G128), .Z(n1263) );
INV_X1 U989 ( .A(G146), .ZN(n1265) );
XOR2_X1 U990 ( .A(n1266), .B(n1166), .Z(n1262) );
AND2_X1 U991 ( .A1(G224), .A2(n1065), .ZN(n1166) );
NAND2_X1 U992 ( .A1(KEYINPUT44), .A2(n1165), .ZN(n1266) );
XOR2_X1 U993 ( .A(KEYINPUT18), .B(n1259), .Z(n1260) );
INV_X1 U994 ( .A(n1137), .ZN(n1259) );
XOR2_X1 U995 ( .A(n1267), .B(n1079), .Z(n1137) );
XNOR2_X1 U996 ( .A(n1189), .B(G122), .ZN(n1079) );
INV_X1 U997 ( .A(G110), .ZN(n1189) );
NAND2_X1 U998 ( .A1(KEYINPUT6), .A2(n1081), .ZN(n1267) );
XOR2_X1 U999 ( .A(n1268), .B(n1237), .Z(n1081) );
XOR2_X1 U1000 ( .A(G101), .B(KEYINPUT25), .Z(n1237) );
XOR2_X1 U1001 ( .A(n1224), .B(n1269), .Z(n1268) );
NOR2_X1 U1002 ( .A1(KEYINPUT59), .A2(n1270), .ZN(n1269) );
XNOR2_X1 U1003 ( .A(n1240), .B(KEYINPUT13), .ZN(n1270) );
XOR2_X1 U1004 ( .A(n1271), .B(n1272), .Z(n1240) );
INV_X1 U1005 ( .A(G104), .ZN(n1271) );
XOR2_X1 U1006 ( .A(n1273), .B(n1274), .Z(n1224) );
XOR2_X1 U1007 ( .A(KEYINPUT5), .B(G116), .Z(n1274) );
XNOR2_X1 U1008 ( .A(G113), .B(n1201), .ZN(n1273) );
XOR2_X1 U1009 ( .A(G119), .B(KEYINPUT46), .Z(n1201) );
INV_X1 U1010 ( .A(n1178), .ZN(n996) );
NOR2_X1 U1011 ( .A1(n1175), .A2(n1173), .ZN(n1178) );
XOR2_X1 U1012 ( .A(n1275), .B(n1099), .Z(n1173) );
INV_X1 U1013 ( .A(n1045), .ZN(n1099) );
NAND2_X1 U1014 ( .A1(n1102), .A2(n1205), .ZN(n1045) );
INV_X1 U1015 ( .A(G902), .ZN(n1205) );
INV_X1 U1016 ( .A(n1105), .ZN(n1102) );
XOR2_X1 U1017 ( .A(n1276), .B(n1277), .Z(n1105) );
XOR2_X1 U1018 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U1019 ( .A(G122), .B(G113), .Z(n1279) );
XOR2_X1 U1020 ( .A(KEYINPUT40), .B(G143), .Z(n1278) );
XOR2_X1 U1021 ( .A(n1280), .B(n1281), .Z(n1276) );
XOR2_X1 U1022 ( .A(G104), .B(n1282), .Z(n1281) );
NOR2_X1 U1023 ( .A1(KEYINPUT11), .A2(n1283), .ZN(n1282) );
XOR2_X1 U1024 ( .A(G146), .B(n1057), .Z(n1283) );
XNOR2_X1 U1025 ( .A(n1165), .B(G140), .ZN(n1057) );
INV_X1 U1026 ( .A(G125), .ZN(n1165) );
XOR2_X1 U1027 ( .A(n1284), .B(n1062), .Z(n1280) );
INV_X1 U1028 ( .A(n1238), .ZN(n1062) );
XNOR2_X1 U1029 ( .A(G131), .B(KEYINPUT42), .ZN(n1238) );
NAND3_X1 U1030 ( .A1(n1226), .A2(n1065), .A3(G214), .ZN(n1284) );
INV_X1 U1031 ( .A(G237), .ZN(n1226) );
NAND2_X1 U1032 ( .A1(KEYINPUT28), .A2(n1103), .ZN(n1275) );
INV_X1 U1033 ( .A(G475), .ZN(n1103) );
INV_X1 U1034 ( .A(n1028), .ZN(n1175) );
XOR2_X1 U1035 ( .A(n1285), .B(G478), .Z(n1028) );
OR2_X1 U1036 ( .A1(n1096), .A2(G902), .ZN(n1285) );
XNOR2_X1 U1037 ( .A(n1286), .B(n1287), .ZN(n1096) );
XOR2_X1 U1038 ( .A(G128), .B(n1288), .Z(n1287) );
XOR2_X1 U1039 ( .A(G143), .B(G134), .Z(n1288) );
XOR2_X1 U1040 ( .A(n1289), .B(n1290), .Z(n1286) );
AND2_X1 U1041 ( .A1(n1197), .A2(G217), .ZN(n1290) );
AND2_X1 U1042 ( .A1(G234), .A2(n1065), .ZN(n1197) );
INV_X1 U1043 ( .A(G953), .ZN(n1065) );
NAND3_X1 U1044 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n1289) );
NAND2_X1 U1045 ( .A1(n1272), .A2(n1294), .ZN(n1293) );
OR3_X1 U1046 ( .A1(n1294), .A2(n1272), .A3(KEYINPUT0), .ZN(n1292) );
XNOR2_X1 U1047 ( .A(G107), .B(KEYINPUT49), .ZN(n1272) );
OR2_X1 U1048 ( .A1(KEYINPUT51), .A2(n1295), .ZN(n1294) );
NAND2_X1 U1049 ( .A1(KEYINPUT0), .A2(n1295), .ZN(n1291) );
XOR2_X1 U1050 ( .A(G116), .B(n1186), .Z(n1295) );
INV_X1 U1051 ( .A(G122), .ZN(n1186) );
endmodule


