//Key = 1011001000011011111000001100100101101110101110100110011111111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340;

XNOR2_X1 U739 ( .A(n1019), .B(n1020), .ZN(G9) );
NOR2_X1 U740 ( .A1(G107), .A2(KEYINPUT26), .ZN(n1020) );
NOR2_X1 U741 ( .A1(n1021), .A2(n1022), .ZN(G75) );
NOR4_X1 U742 ( .A1(n1023), .A2(n1024), .A3(G953), .A4(n1025), .ZN(n1022) );
NOR2_X1 U743 ( .A1(KEYINPUT57), .A2(n1026), .ZN(n1024) );
AND2_X1 U744 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND3_X1 U745 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1023) );
NAND2_X1 U746 ( .A1(n1028), .A2(n1032), .ZN(n1030) );
NAND3_X1 U747 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1032) );
NAND2_X1 U748 ( .A1(KEYINPUT57), .A2(n1027), .ZN(n1035) );
NAND2_X1 U749 ( .A1(n1036), .A2(n1037), .ZN(n1027) );
NAND2_X1 U750 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U751 ( .A1(n1040), .A2(n1041), .ZN(n1036) );
NAND2_X1 U752 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND3_X1 U753 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NAND2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1042) );
NAND2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U756 ( .A1(n1046), .A2(n1051), .ZN(n1050) );
NAND2_X1 U757 ( .A1(n1040), .A2(n1052), .ZN(n1034) );
NAND2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND4_X1 U759 ( .A1(KEYINPUT11), .A2(n1055), .A3(n1056), .A4(n1046), .ZN(n1054) );
NOR2_X1 U760 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U761 ( .A1(n1045), .A2(n1059), .ZN(n1053) );
NAND2_X1 U762 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND3_X1 U763 ( .A1(n1062), .A2(n1047), .A3(n1063), .ZN(n1061) );
NAND2_X1 U764 ( .A1(n1046), .A2(n1064), .ZN(n1060) );
NAND2_X1 U765 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
OR2_X1 U766 ( .A1(n1057), .A2(KEYINPUT11), .ZN(n1066) );
XOR2_X1 U767 ( .A(n1067), .B(KEYINPUT41), .Z(n1057) );
NAND2_X1 U768 ( .A1(n1038), .A2(n1068), .ZN(n1033) );
AND3_X1 U769 ( .A1(n1045), .A2(n1047), .A3(n1046), .ZN(n1038) );
INV_X1 U770 ( .A(n1069), .ZN(n1028) );
NOR3_X1 U771 ( .A1(n1025), .A2(G953), .A3(G952), .ZN(n1021) );
AND4_X1 U772 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1025) );
NOR4_X1 U773 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1073) );
XNOR2_X1 U774 ( .A(KEYINPUT22), .B(n1078), .ZN(n1077) );
XOR2_X1 U775 ( .A(KEYINPUT58), .B(n1079), .Z(n1076) );
NOR3_X1 U776 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
XNOR2_X1 U777 ( .A(G472), .B(n1083), .ZN(n1080) );
NOR2_X1 U778 ( .A1(n1084), .A2(n1085), .ZN(n1075) );
NOR2_X1 U779 ( .A1(G469), .A2(n1086), .ZN(n1074) );
NOR2_X1 U780 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
AND2_X1 U781 ( .A1(n1085), .A2(KEYINPUT38), .ZN(n1088) );
NAND2_X1 U782 ( .A1(KEYINPUT17), .A2(n1089), .ZN(n1085) );
NOR2_X1 U783 ( .A1(KEYINPUT38), .A2(n1090), .ZN(n1087) );
XOR2_X1 U784 ( .A(n1091), .B(KEYINPUT30), .Z(n1072) );
OR2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U786 ( .A1(n1093), .A2(n1092), .ZN(n1070) );
XOR2_X1 U787 ( .A(n1094), .B(n1095), .Z(G72) );
XOR2_X1 U788 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
AND2_X1 U790 ( .A1(G227), .A2(G900), .ZN(n1098) );
NAND2_X1 U791 ( .A1(n1100), .A2(n1101), .ZN(n1096) );
NAND2_X1 U792 ( .A1(G953), .A2(n1102), .ZN(n1101) );
XOR2_X1 U793 ( .A(n1103), .B(n1104), .Z(n1100) );
XOR2_X1 U794 ( .A(n1105), .B(n1106), .Z(n1104) );
XNOR2_X1 U795 ( .A(n1107), .B(G134), .ZN(n1106) );
NOR2_X1 U796 ( .A1(G131), .A2(KEYINPUT1), .ZN(n1105) );
XOR2_X1 U797 ( .A(n1108), .B(n1109), .Z(n1103) );
NAND2_X1 U798 ( .A1(n1099), .A2(n1110), .ZN(n1094) );
XOR2_X1 U799 ( .A(n1111), .B(n1112), .Z(G69) );
XOR2_X1 U800 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U801 ( .A1(n1099), .A2(n1115), .ZN(n1114) );
XOR2_X1 U802 ( .A(KEYINPUT62), .B(n1116), .Z(n1115) );
AND2_X1 U803 ( .A1(G224), .A2(G898), .ZN(n1116) );
NAND2_X1 U804 ( .A1(n1117), .A2(n1118), .ZN(n1113) );
NAND2_X1 U805 ( .A1(G953), .A2(n1119), .ZN(n1118) );
XNOR2_X1 U806 ( .A(n1120), .B(n1121), .ZN(n1117) );
NAND2_X1 U807 ( .A1(n1099), .A2(n1122), .ZN(n1111) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1124), .ZN(G66) );
XOR2_X1 U809 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR3_X1 U810 ( .A1(n1127), .A2(KEYINPUT39), .A3(n1128), .ZN(n1125) );
NOR2_X1 U811 ( .A1(n1123), .A2(n1129), .ZN(G63) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1129) );
AND2_X1 U813 ( .A1(G478), .A2(n1132), .ZN(n1130) );
NOR2_X1 U814 ( .A1(n1123), .A2(n1133), .ZN(G60) );
XNOR2_X1 U815 ( .A(n1134), .B(n1135), .ZN(n1133) );
AND2_X1 U816 ( .A1(G475), .A2(n1132), .ZN(n1134) );
XNOR2_X1 U817 ( .A(n1136), .B(n1137), .ZN(G6) );
NOR4_X1 U818 ( .A1(KEYINPUT52), .A2(n1138), .A3(n1067), .A4(n1139), .ZN(n1137) );
NOR2_X1 U819 ( .A1(n1140), .A2(n1141), .ZN(G57) );
XOR2_X1 U820 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U821 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U822 ( .A(KEYINPUT4), .B(n1146), .Z(n1145) );
AND2_X1 U823 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NOR2_X1 U824 ( .A1(KEYINPUT9), .A2(n1149), .ZN(n1142) );
XOR2_X1 U825 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U827 ( .A1(KEYINPUT19), .A2(n1154), .ZN(n1153) );
NAND3_X1 U828 ( .A1(n1132), .A2(G472), .A3(KEYINPUT40), .ZN(n1150) );
INV_X1 U829 ( .A(n1127), .ZN(n1132) );
XNOR2_X1 U830 ( .A(n1123), .B(KEYINPUT2), .ZN(n1140) );
NOR2_X1 U831 ( .A1(n1123), .A2(n1155), .ZN(G54) );
NOR2_X1 U832 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U833 ( .A(KEYINPUT61), .B(n1158), .Z(n1157) );
AND2_X1 U834 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U835 ( .A1(n1160), .A2(n1159), .ZN(n1156) );
XNOR2_X1 U836 ( .A(n1161), .B(n1162), .ZN(n1159) );
XOR2_X1 U837 ( .A(n1163), .B(n1164), .Z(n1162) );
NAND2_X1 U838 ( .A1(KEYINPUT36), .A2(n1165), .ZN(n1164) );
NAND3_X1 U839 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1163) );
OR2_X1 U840 ( .A1(n1169), .A2(KEYINPUT8), .ZN(n1167) );
NAND2_X1 U841 ( .A1(KEYINPUT8), .A2(n1170), .ZN(n1166) );
INV_X1 U842 ( .A(n1171), .ZN(n1170) );
NOR2_X1 U843 ( .A1(n1127), .A2(n1084), .ZN(n1160) );
INV_X1 U844 ( .A(G469), .ZN(n1084) );
NOR2_X1 U845 ( .A1(n1123), .A2(n1172), .ZN(G51) );
XOR2_X1 U846 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U847 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR3_X1 U848 ( .A1(n1127), .A2(KEYINPUT23), .A3(n1092), .ZN(n1175) );
NAND2_X1 U849 ( .A1(G902), .A2(n1177), .ZN(n1127) );
NAND2_X1 U850 ( .A1(n1031), .A2(n1029), .ZN(n1177) );
INV_X1 U851 ( .A(n1110), .ZN(n1029) );
NAND4_X1 U852 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1110) );
NOR4_X1 U853 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181) );
NOR2_X1 U854 ( .A1(n1186), .A2(n1187), .ZN(n1180) );
NOR3_X1 U855 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
INV_X1 U856 ( .A(n1122), .ZN(n1031) );
NAND4_X1 U857 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1122) );
NOR4_X1 U858 ( .A1(n1195), .A2(n1019), .A3(n1196), .A4(n1197), .ZN(n1194) );
NOR3_X1 U859 ( .A1(n1067), .A2(n1138), .A3(n1190), .ZN(n1019) );
INV_X1 U860 ( .A(n1047), .ZN(n1067) );
NOR2_X1 U861 ( .A1(n1198), .A2(n1199), .ZN(n1193) );
NOR3_X1 U862 ( .A1(n1200), .A2(n1139), .A3(n1201), .ZN(n1199) );
XNOR2_X1 U863 ( .A(KEYINPUT31), .B(n1202), .ZN(n1201) );
NAND3_X1 U864 ( .A1(n1203), .A2(n1204), .A3(n1047), .ZN(n1200) );
XOR2_X1 U865 ( .A(n1205), .B(KEYINPUT24), .Z(n1173) );
NAND3_X1 U866 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1205) );
NAND2_X1 U867 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
OR3_X1 U868 ( .A1(n1210), .A2(n1209), .A3(KEYINPUT21), .ZN(n1207) );
OR2_X1 U869 ( .A1(KEYINPUT35), .A2(n1211), .ZN(n1210) );
NAND2_X1 U870 ( .A1(KEYINPUT21), .A2(n1211), .ZN(n1206) );
NOR2_X1 U871 ( .A1(n1099), .A2(G952), .ZN(n1123) );
XNOR2_X1 U872 ( .A(n1212), .B(n1186), .ZN(G48) );
NOR3_X1 U873 ( .A1(n1139), .A2(n1189), .A3(n1188), .ZN(n1186) );
XOR2_X1 U874 ( .A(n1213), .B(G143), .Z(G45) );
NAND2_X1 U875 ( .A1(KEYINPUT43), .A2(n1179), .ZN(n1213) );
NAND4_X1 U876 ( .A1(n1214), .A2(n1203), .A3(n1215), .A4(n1216), .ZN(n1179) );
XNOR2_X1 U877 ( .A(G140), .B(n1217), .ZN(G42) );
NOR2_X1 U878 ( .A1(n1185), .A2(KEYINPUT51), .ZN(n1217) );
NOR3_X1 U879 ( .A1(n1218), .A2(n1202), .A3(n1219), .ZN(n1185) );
XNOR2_X1 U880 ( .A(n1107), .B(n1184), .ZN(G39) );
NOR3_X1 U881 ( .A1(n1219), .A2(n1081), .A3(n1188), .ZN(n1184) );
INV_X1 U882 ( .A(n1046), .ZN(n1219) );
XNOR2_X1 U883 ( .A(G134), .B(n1220), .ZN(G36) );
NAND2_X1 U884 ( .A1(KEYINPUT49), .A2(n1183), .ZN(n1220) );
AND3_X1 U885 ( .A1(n1214), .A2(n1068), .A3(n1046), .ZN(n1183) );
XNOR2_X1 U886 ( .A(G131), .B(n1178), .ZN(G33) );
NAND3_X1 U887 ( .A1(n1214), .A2(n1039), .A3(n1046), .ZN(n1178) );
NOR2_X1 U888 ( .A1(n1221), .A2(n1062), .ZN(n1046) );
AND3_X1 U889 ( .A1(n1051), .A2(n1222), .A3(n1044), .ZN(n1214) );
XOR2_X1 U890 ( .A(G128), .B(n1223), .Z(G30) );
NOR3_X1 U891 ( .A1(n1224), .A2(n1190), .A3(n1188), .ZN(n1223) );
NAND4_X1 U892 ( .A1(n1051), .A2(n1082), .A3(n1225), .A4(n1222), .ZN(n1188) );
INV_X1 U893 ( .A(n1068), .ZN(n1190) );
XNOR2_X1 U894 ( .A(KEYINPUT50), .B(n1189), .ZN(n1224) );
INV_X1 U895 ( .A(n1203), .ZN(n1189) );
XNOR2_X1 U896 ( .A(n1198), .B(n1226), .ZN(G3) );
NAND2_X1 U897 ( .A1(KEYINPUT44), .A2(G101), .ZN(n1226) );
NOR3_X1 U898 ( .A1(n1081), .A2(n1138), .A3(n1227), .ZN(n1198) );
INV_X1 U899 ( .A(n1044), .ZN(n1227) );
XNOR2_X1 U900 ( .A(n1182), .B(n1228), .ZN(G27) );
NAND2_X1 U901 ( .A1(KEYINPUT54), .A2(G125), .ZN(n1228) );
NOR2_X1 U902 ( .A1(n1218), .A2(n1049), .ZN(n1182) );
NAND3_X1 U903 ( .A1(n1229), .A2(n1222), .A3(n1039), .ZN(n1218) );
NAND2_X1 U904 ( .A1(n1069), .A2(n1230), .ZN(n1222) );
NAND4_X1 U905 ( .A1(G953), .A2(G902), .A3(n1231), .A4(n1102), .ZN(n1230) );
INV_X1 U906 ( .A(G900), .ZN(n1102) );
XNOR2_X1 U907 ( .A(G122), .B(n1191), .ZN(G24) );
NAND4_X1 U908 ( .A1(n1232), .A2(n1047), .A3(n1215), .A4(n1216), .ZN(n1191) );
NOR2_X1 U909 ( .A1(n1225), .A2(n1082), .ZN(n1047) );
XNOR2_X1 U910 ( .A(G119), .B(n1192), .ZN(G21) );
NAND4_X1 U911 ( .A1(n1232), .A2(n1040), .A3(n1082), .A4(n1225), .ZN(n1192) );
XOR2_X1 U912 ( .A(n1233), .B(n1197), .Z(G18) );
AND3_X1 U913 ( .A1(n1044), .A2(n1068), .A3(n1232), .ZN(n1197) );
NOR2_X1 U914 ( .A1(n1216), .A2(n1234), .ZN(n1068) );
XNOR2_X1 U915 ( .A(G116), .B(KEYINPUT6), .ZN(n1233) );
XNOR2_X1 U916 ( .A(n1235), .B(n1196), .ZN(G15) );
AND3_X1 U917 ( .A1(n1044), .A2(n1039), .A3(n1232), .ZN(n1196) );
NOR2_X1 U918 ( .A1(n1049), .A2(n1236), .ZN(n1232) );
NAND2_X1 U919 ( .A1(n1045), .A2(n1203), .ZN(n1049) );
NOR2_X1 U920 ( .A1(n1058), .A2(n1055), .ZN(n1045) );
INV_X1 U921 ( .A(n1071), .ZN(n1055) );
INV_X1 U922 ( .A(n1139), .ZN(n1039) );
NAND2_X1 U923 ( .A1(n1234), .A2(n1216), .ZN(n1139) );
INV_X1 U924 ( .A(n1215), .ZN(n1234) );
NOR2_X1 U925 ( .A1(n1082), .A2(n1237), .ZN(n1044) );
NAND2_X1 U926 ( .A1(n1238), .A2(n1239), .ZN(G12) );
NAND2_X1 U927 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
XOR2_X1 U928 ( .A(KEYINPUT53), .B(n1242), .Z(n1238) );
NOR2_X1 U929 ( .A1(n1241), .A2(n1240), .ZN(n1242) );
NAND2_X1 U930 ( .A1(n1243), .A2(n1244), .ZN(n1240) );
NAND2_X1 U931 ( .A1(n1195), .A2(n1245), .ZN(n1244) );
INV_X1 U932 ( .A(KEYINPUT10), .ZN(n1245) );
NOR3_X1 U933 ( .A1(n1081), .A2(n1138), .A3(n1065), .ZN(n1195) );
NAND3_X1 U934 ( .A1(n1203), .A2(n1204), .A3(n1051), .ZN(n1138) );
INV_X1 U935 ( .A(n1202), .ZN(n1051) );
INV_X1 U936 ( .A(n1040), .ZN(n1081) );
NAND4_X1 U937 ( .A1(n1229), .A2(n1040), .A3(n1246), .A4(KEYINPUT10), .ZN(n1243) );
NOR3_X1 U938 ( .A1(n1202), .A2(n1203), .A3(n1236), .ZN(n1246) );
INV_X1 U939 ( .A(n1204), .ZN(n1236) );
NAND2_X1 U940 ( .A1(n1247), .A2(n1069), .ZN(n1204) );
NAND3_X1 U941 ( .A1(n1231), .A2(n1099), .A3(G952), .ZN(n1069) );
XOR2_X1 U942 ( .A(n1248), .B(KEYINPUT47), .Z(n1247) );
NAND4_X1 U943 ( .A1(G953), .A2(G902), .A3(n1119), .A4(n1231), .ZN(n1248) );
NAND2_X1 U944 ( .A1(G237), .A2(G234), .ZN(n1231) );
XOR2_X1 U945 ( .A(KEYINPUT25), .B(G898), .Z(n1119) );
NOR2_X1 U946 ( .A1(n1063), .A2(n1062), .ZN(n1203) );
INV_X1 U947 ( .A(n1078), .ZN(n1062) );
NAND2_X1 U948 ( .A1(G214), .A2(n1249), .ZN(n1078) );
INV_X1 U949 ( .A(n1221), .ZN(n1063) );
XNOR2_X1 U950 ( .A(n1093), .B(n1092), .ZN(n1221) );
NAND2_X1 U951 ( .A1(G210), .A2(n1249), .ZN(n1092) );
NAND2_X1 U952 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
AND3_X1 U953 ( .A1(n1252), .A2(n1251), .A3(n1253), .ZN(n1093) );
XOR2_X1 U954 ( .A(KEYINPUT16), .B(n1254), .Z(n1253) );
NOR2_X1 U955 ( .A1(n1255), .A2(n1176), .ZN(n1254) );
NAND2_X1 U956 ( .A1(n1255), .A2(n1176), .ZN(n1252) );
XOR2_X1 U957 ( .A(n1121), .B(n1256), .Z(n1176) );
NOR2_X1 U958 ( .A1(KEYINPUT5), .A2(n1120), .ZN(n1256) );
AND2_X1 U959 ( .A1(n1257), .A2(n1258), .ZN(n1120) );
NAND2_X1 U960 ( .A1(n1259), .A2(n1235), .ZN(n1258) );
INV_X1 U961 ( .A(G113), .ZN(n1235) );
NAND2_X1 U962 ( .A1(n1260), .A2(G113), .ZN(n1257) );
XOR2_X1 U963 ( .A(n1259), .B(KEYINPUT60), .Z(n1260) );
XOR2_X1 U964 ( .A(n1261), .B(n1262), .Z(n1259) );
NAND2_X1 U965 ( .A1(n1263), .A2(n1264), .ZN(n1261) );
NAND2_X1 U966 ( .A1(G101), .A2(n1265), .ZN(n1264) );
XOR2_X1 U967 ( .A(KEYINPUT14), .B(n1266), .Z(n1263) );
NOR2_X1 U968 ( .A1(G101), .A2(n1265), .ZN(n1266) );
XNOR2_X1 U969 ( .A(G107), .B(n1136), .ZN(n1265) );
INV_X1 U970 ( .A(G104), .ZN(n1136) );
XNOR2_X1 U971 ( .A(G110), .B(n1267), .ZN(n1121) );
XOR2_X1 U972 ( .A(n1209), .B(n1268), .Z(n1255) );
XNOR2_X1 U973 ( .A(n1269), .B(KEYINPUT7), .ZN(n1268) );
NAND2_X1 U974 ( .A1(KEYINPUT59), .A2(n1270), .ZN(n1269) );
INV_X1 U975 ( .A(n1211), .ZN(n1270) );
NAND2_X1 U976 ( .A1(G224), .A2(n1099), .ZN(n1211) );
XOR2_X1 U977 ( .A(n1271), .B(n1272), .Z(n1209) );
XOR2_X1 U978 ( .A(KEYINPUT63), .B(G125), .Z(n1272) );
NAND2_X1 U979 ( .A1(n1058), .A2(n1071), .ZN(n1202) );
NAND2_X1 U980 ( .A1(G221), .A2(n1273), .ZN(n1071) );
XNOR2_X1 U981 ( .A(n1274), .B(G469), .ZN(n1058) );
NAND2_X1 U982 ( .A1(KEYINPUT15), .A2(n1090), .ZN(n1274) );
INV_X1 U983 ( .A(n1089), .ZN(n1090) );
NAND2_X1 U984 ( .A1(n1251), .A2(n1275), .ZN(n1089) );
NAND2_X1 U985 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND3_X1 U986 ( .A1(n1169), .A2(n1168), .A3(n1278), .ZN(n1277) );
XOR2_X1 U987 ( .A(KEYINPUT55), .B(n1279), .Z(n1276) );
NOR2_X1 U988 ( .A1(n1280), .A2(n1278), .ZN(n1279) );
XNOR2_X1 U989 ( .A(n1161), .B(n1165), .ZN(n1278) );
XOR2_X1 U990 ( .A(n1108), .B(G146), .Z(n1165) );
XOR2_X1 U991 ( .A(n1281), .B(n1282), .Z(n1108) );
XOR2_X1 U992 ( .A(KEYINPUT28), .B(G143), .Z(n1282) );
NAND2_X1 U993 ( .A1(KEYINPUT33), .A2(G128), .ZN(n1281) );
XOR2_X1 U994 ( .A(n1283), .B(n1284), .Z(n1161) );
XNOR2_X1 U995 ( .A(n1285), .B(n1148), .ZN(n1283) );
NAND3_X1 U996 ( .A1(n1286), .A2(n1287), .A3(KEYINPUT56), .ZN(n1285) );
NAND2_X1 U997 ( .A1(KEYINPUT37), .A2(n1288), .ZN(n1287) );
XOR2_X1 U998 ( .A(G107), .B(n1289), .Z(n1288) );
OR3_X1 U999 ( .A1(n1289), .A2(G107), .A3(KEYINPUT37), .ZN(n1286) );
XNOR2_X1 U1000 ( .A(G104), .B(KEYINPUT29), .ZN(n1289) );
AND2_X1 U1001 ( .A1(n1168), .A2(n1169), .ZN(n1280) );
NAND2_X1 U1002 ( .A1(n1290), .A2(n1171), .ZN(n1169) );
OR2_X1 U1003 ( .A1(n1171), .A2(n1290), .ZN(n1168) );
XNOR2_X1 U1004 ( .A(G140), .B(n1241), .ZN(n1290) );
NAND2_X1 U1005 ( .A1(G227), .A2(n1099), .ZN(n1171) );
NOR2_X1 U1006 ( .A1(n1215), .A2(n1216), .ZN(n1040) );
XNOR2_X1 U1007 ( .A(n1291), .B(G475), .ZN(n1216) );
NAND2_X1 U1008 ( .A1(n1135), .A2(n1292), .ZN(n1291) );
XNOR2_X1 U1009 ( .A(KEYINPUT18), .B(n1251), .ZN(n1292) );
XOR2_X1 U1010 ( .A(n1293), .B(n1294), .Z(n1135) );
XOR2_X1 U1011 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1012 ( .A(n1297), .B(n1298), .Z(n1296) );
NOR2_X1 U1013 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XOR2_X1 U1014 ( .A(n1301), .B(KEYINPUT46), .Z(n1300) );
NAND2_X1 U1015 ( .A1(n1302), .A2(G146), .ZN(n1301) );
NOR2_X1 U1016 ( .A1(G146), .A2(n1302), .ZN(n1299) );
XNOR2_X1 U1017 ( .A(KEYINPUT3), .B(n1303), .ZN(n1302) );
NAND2_X1 U1018 ( .A1(KEYINPUT42), .A2(n1304), .ZN(n1297) );
INV_X1 U1019 ( .A(G131), .ZN(n1304) );
NAND3_X1 U1020 ( .A1(n1250), .A2(n1099), .A3(G214), .ZN(n1295) );
XOR2_X1 U1021 ( .A(n1305), .B(n1306), .Z(n1293) );
XNOR2_X1 U1022 ( .A(G143), .B(n1267), .ZN(n1306) );
INV_X1 U1023 ( .A(G122), .ZN(n1267) );
XNOR2_X1 U1024 ( .A(G104), .B(G113), .ZN(n1305) );
XNOR2_X1 U1025 ( .A(n1307), .B(G478), .ZN(n1215) );
OR2_X1 U1026 ( .A1(n1131), .A2(G902), .ZN(n1307) );
XNOR2_X1 U1027 ( .A(n1308), .B(n1309), .ZN(n1131) );
XOR2_X1 U1028 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U1029 ( .A(G107), .B(n1312), .ZN(n1311) );
NOR2_X1 U1030 ( .A1(G143), .A2(KEYINPUT32), .ZN(n1312) );
NAND2_X1 U1031 ( .A1(G217), .A2(n1313), .ZN(n1310) );
XOR2_X1 U1032 ( .A(n1314), .B(n1315), .Z(n1308) );
XOR2_X1 U1033 ( .A(G134), .B(G128), .Z(n1315) );
XNOR2_X1 U1034 ( .A(G116), .B(G122), .ZN(n1314) );
INV_X1 U1035 ( .A(n1065), .ZN(n1229) );
NAND2_X1 U1036 ( .A1(n1237), .A2(n1082), .ZN(n1065) );
XOR2_X1 U1037 ( .A(n1316), .B(n1128), .Z(n1082) );
NAND2_X1 U1038 ( .A1(G217), .A2(n1273), .ZN(n1128) );
NAND2_X1 U1039 ( .A1(G234), .A2(n1251), .ZN(n1273) );
OR2_X1 U1040 ( .A1(n1126), .A2(G902), .ZN(n1316) );
XNOR2_X1 U1041 ( .A(n1317), .B(n1318), .ZN(n1126) );
XOR2_X1 U1042 ( .A(n1319), .B(n1109), .Z(n1318) );
XNOR2_X1 U1043 ( .A(n1212), .B(n1303), .ZN(n1109) );
XOR2_X1 U1044 ( .A(G125), .B(G140), .Z(n1303) );
AND2_X1 U1045 ( .A1(n1313), .A2(G221), .ZN(n1319) );
AND2_X1 U1046 ( .A1(G234), .A2(n1099), .ZN(n1313) );
XOR2_X1 U1047 ( .A(n1320), .B(n1321), .Z(n1317) );
NOR2_X1 U1048 ( .A1(KEYINPUT48), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1049 ( .A(G119), .B(n1323), .Z(n1322) );
XOR2_X1 U1050 ( .A(KEYINPUT27), .B(G128), .Z(n1323) );
XNOR2_X1 U1051 ( .A(G110), .B(G137), .ZN(n1320) );
INV_X1 U1052 ( .A(n1225), .ZN(n1237) );
XOR2_X1 U1053 ( .A(G472), .B(n1324), .Z(n1225) );
NOR2_X1 U1054 ( .A1(KEYINPUT20), .A2(n1083), .ZN(n1324) );
NAND2_X1 U1055 ( .A1(n1325), .A2(n1251), .ZN(n1083) );
INV_X1 U1056 ( .A(G902), .ZN(n1251) );
XOR2_X1 U1057 ( .A(n1326), .B(n1327), .Z(n1325) );
NAND3_X1 U1058 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1327) );
INV_X1 U1059 ( .A(n1144), .ZN(n1330) );
NOR2_X1 U1060 ( .A1(n1148), .A2(n1147), .ZN(n1144) );
NAND3_X1 U1061 ( .A1(KEYINPUT34), .A2(n1147), .A3(n1148), .ZN(n1329) );
NAND3_X1 U1062 ( .A1(n1250), .A2(n1099), .A3(G210), .ZN(n1147) );
INV_X1 U1063 ( .A(G953), .ZN(n1099) );
INV_X1 U1064 ( .A(G237), .ZN(n1250) );
OR2_X1 U1065 ( .A1(n1148), .A2(KEYINPUT34), .ZN(n1328) );
INV_X1 U1066 ( .A(G101), .ZN(n1148) );
NAND2_X1 U1067 ( .A1(n1331), .A2(n1332), .ZN(n1326) );
OR2_X1 U1068 ( .A1(n1152), .A2(n1154), .ZN(n1332) );
XOR2_X1 U1069 ( .A(n1333), .B(KEYINPUT13), .Z(n1331) );
NAND2_X1 U1070 ( .A1(n1154), .A2(n1152), .ZN(n1333) );
NAND2_X1 U1071 ( .A1(n1334), .A2(n1335), .ZN(n1152) );
OR2_X1 U1072 ( .A1(n1262), .A2(G113), .ZN(n1335) );
XOR2_X1 U1073 ( .A(n1336), .B(KEYINPUT45), .Z(n1334) );
NAND2_X1 U1074 ( .A1(G113), .A2(n1262), .ZN(n1336) );
XOR2_X1 U1075 ( .A(G116), .B(G119), .Z(n1262) );
XOR2_X1 U1076 ( .A(n1271), .B(n1284), .Z(n1154) );
XNOR2_X1 U1077 ( .A(n1337), .B(G131), .ZN(n1284) );
NAND2_X1 U1078 ( .A1(n1338), .A2(KEYINPUT12), .ZN(n1337) );
XOR2_X1 U1079 ( .A(n1339), .B(G134), .Z(n1338) );
NAND2_X1 U1080 ( .A1(KEYINPUT0), .A2(n1107), .ZN(n1339) );
INV_X1 U1081 ( .A(G137), .ZN(n1107) );
XNOR2_X1 U1082 ( .A(G128), .B(n1340), .ZN(n1271) );
XNOR2_X1 U1083 ( .A(n1212), .B(G143), .ZN(n1340) );
INV_X1 U1084 ( .A(G146), .ZN(n1212) );
INV_X1 U1085 ( .A(G110), .ZN(n1241) );
endmodule


