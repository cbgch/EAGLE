//Key = 0010100010100100100101111001010000111010100000001110001000011011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375;

XOR2_X1 U764 ( .A(n1046), .B(n1047), .Z(G9) );
NOR2_X1 U765 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR4_X1 U766 ( .A1(G953), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1049) );
NOR2_X1 U767 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U768 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U769 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U770 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U771 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U772 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U773 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U774 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR2_X1 U775 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR2_X1 U776 ( .A1(n1071), .A2(n1072), .ZN(n1063) );
NOR2_X1 U777 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR3_X1 U778 ( .A1(n1072), .A2(n1075), .A3(n1066), .ZN(n1059) );
XOR2_X1 U779 ( .A(n1076), .B(n1077), .Z(n1075) );
NOR4_X1 U780 ( .A1(n1078), .A2(n1066), .A3(n1062), .A4(n1072), .ZN(n1055) );
NOR2_X1 U781 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR3_X1 U782 ( .A1(n1050), .A2(G953), .A3(G952), .ZN(n1048) );
AND4_X1 U783 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1050) );
NOR3_X1 U784 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
XOR2_X1 U785 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U786 ( .A1(n1090), .A2(KEYINPUT41), .ZN(n1089) );
XOR2_X1 U787 ( .A(n1091), .B(n1092), .Z(n1086) );
NAND2_X1 U788 ( .A1(KEYINPUT13), .A2(n1093), .ZN(n1091) );
NAND3_X1 U789 ( .A1(n1094), .A2(n1070), .A3(n1095), .ZN(n1085) );
NAND2_X1 U790 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR3_X1 U791 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1083) );
NOR2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U793 ( .A(n1103), .B(KEYINPUT40), .Z(n1102) );
NOR2_X1 U794 ( .A1(G472), .A2(n1104), .ZN(n1099) );
XOR2_X1 U795 ( .A(n1103), .B(n1105), .Z(n1104) );
XNOR2_X1 U796 ( .A(KEYINPUT62), .B(KEYINPUT37), .ZN(n1105) );
XOR2_X1 U797 ( .A(KEYINPUT56), .B(n1106), .Z(n1098) );
NOR2_X1 U798 ( .A1(n1097), .A2(n1096), .ZN(n1106) );
XOR2_X1 U799 ( .A(n1107), .B(KEYINPUT34), .Z(n1096) );
XOR2_X1 U800 ( .A(n1108), .B(n1109), .Z(n1081) );
XOR2_X1 U801 ( .A(n1110), .B(n1111), .Z(G72) );
XOR2_X1 U802 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND2_X1 U803 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U804 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND3_X1 U805 ( .A1(KEYINPUT16), .A2(n1118), .A3(n1119), .ZN(n1112) );
XOR2_X1 U806 ( .A(n1120), .B(n1121), .Z(n1119) );
XNOR2_X1 U807 ( .A(G125), .B(n1122), .ZN(n1121) );
NAND2_X1 U808 ( .A1(KEYINPUT23), .A2(n1123), .ZN(n1122) );
NAND2_X1 U809 ( .A1(n1124), .A2(n1125), .ZN(n1118) );
NOR2_X1 U810 ( .A1(n1126), .A2(n1114), .ZN(n1110) );
AND2_X1 U811 ( .A1(G227), .A2(G900), .ZN(n1126) );
XOR2_X1 U812 ( .A(n1127), .B(n1128), .Z(G69) );
NOR2_X1 U813 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U814 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U815 ( .A(n1133), .B(KEYINPUT18), .Z(n1132) );
AND2_X1 U816 ( .A1(n1133), .A2(n1131), .ZN(n1129) );
AND2_X1 U817 ( .A1(n1134), .A2(n1135), .ZN(n1131) );
NAND2_X1 U818 ( .A1(n1124), .A2(n1136), .ZN(n1135) );
XOR2_X1 U819 ( .A(n1137), .B(n1138), .Z(n1134) );
NAND2_X1 U820 ( .A1(n1114), .A2(n1139), .ZN(n1133) );
NAND3_X1 U821 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
XOR2_X1 U822 ( .A(n1143), .B(KEYINPUT52), .Z(n1142) );
OR2_X1 U823 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U824 ( .A(n1146), .B(KEYINPUT55), .Z(n1140) );
NAND2_X1 U825 ( .A1(G953), .A2(n1147), .ZN(n1127) );
NAND2_X1 U826 ( .A1(G898), .A2(G224), .ZN(n1147) );
NOR2_X1 U827 ( .A1(n1148), .A2(n1149), .ZN(G66) );
NOR3_X1 U828 ( .A1(n1092), .A2(n1150), .A3(n1151), .ZN(n1149) );
NOR3_X1 U829 ( .A1(n1152), .A2(n1093), .A3(n1153), .ZN(n1151) );
NOR2_X1 U830 ( .A1(n1154), .A2(n1155), .ZN(n1150) );
NOR2_X1 U831 ( .A1(n1156), .A2(n1093), .ZN(n1154) );
NOR2_X1 U832 ( .A1(n1148), .A2(n1157), .ZN(G63) );
XOR2_X1 U833 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND3_X1 U834 ( .A1(G478), .A2(n1052), .A3(n1160), .ZN(n1158) );
XOR2_X1 U835 ( .A(n1161), .B(KEYINPUT19), .Z(n1160) );
NOR3_X1 U836 ( .A1(n1148), .A2(n1162), .A3(n1163), .ZN(G60) );
NOR2_X1 U837 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NOR2_X1 U838 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NOR3_X1 U839 ( .A1(n1168), .A2(KEYINPUT25), .A3(n1169), .ZN(n1167) );
AND2_X1 U840 ( .A1(n1168), .A2(n1169), .ZN(n1166) );
INV_X1 U841 ( .A(KEYINPUT38), .ZN(n1168) );
INV_X1 U842 ( .A(n1170), .ZN(n1164) );
NOR2_X1 U843 ( .A1(n1171), .A2(n1170), .ZN(n1162) );
NOR2_X1 U844 ( .A1(KEYINPUT25), .A2(n1169), .ZN(n1171) );
NAND3_X1 U845 ( .A1(G902), .A2(n1172), .A3(G475), .ZN(n1169) );
XOR2_X1 U846 ( .A(KEYINPUT36), .B(n1156), .Z(n1172) );
INV_X1 U847 ( .A(n1052), .ZN(n1156) );
XOR2_X1 U848 ( .A(G104), .B(n1173), .Z(G6) );
NOR2_X1 U849 ( .A1(n1145), .A2(n1174), .ZN(n1173) );
XNOR2_X1 U850 ( .A(KEYINPUT59), .B(n1175), .ZN(n1174) );
NOR2_X1 U851 ( .A1(n1148), .A2(n1176), .ZN(G57) );
XOR2_X1 U852 ( .A(n1177), .B(n1178), .Z(n1176) );
XNOR2_X1 U853 ( .A(n1179), .B(n1120), .ZN(n1178) );
XOR2_X1 U854 ( .A(n1180), .B(n1181), .Z(n1177) );
NOR2_X1 U855 ( .A1(n1101), .A2(n1153), .ZN(n1181) );
INV_X1 U856 ( .A(G472), .ZN(n1101) );
NAND2_X1 U857 ( .A1(n1182), .A2(KEYINPUT60), .ZN(n1180) );
XOR2_X1 U858 ( .A(n1183), .B(G101), .Z(n1182) );
NOR2_X1 U859 ( .A1(n1148), .A2(n1184), .ZN(G54) );
XOR2_X1 U860 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U861 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U862 ( .A(G143), .B(n1189), .Z(n1188) );
NOR2_X1 U863 ( .A1(KEYINPUT0), .A2(n1190), .ZN(n1189) );
XOR2_X1 U864 ( .A(G131), .B(n1191), .Z(n1190) );
NOR3_X1 U865 ( .A1(n1153), .A2(KEYINPUT9), .A3(n1088), .ZN(n1187) );
XNOR2_X1 U866 ( .A(n1192), .B(n1193), .ZN(n1185) );
XOR2_X1 U867 ( .A(n1194), .B(n1195), .Z(n1193) );
NAND2_X1 U868 ( .A1(KEYINPUT54), .A2(n1138), .ZN(n1195) );
NAND3_X1 U869 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1194) );
NAND2_X1 U870 ( .A1(n1199), .A2(n1200), .ZN(n1197) );
XOR2_X1 U871 ( .A(n1201), .B(n1123), .Z(n1199) );
NAND3_X1 U872 ( .A1(n1201), .A2(n1123), .A3(G110), .ZN(n1196) );
NOR2_X1 U873 ( .A1(n1148), .A2(n1202), .ZN(G51) );
XOR2_X1 U874 ( .A(n1203), .B(n1204), .Z(n1202) );
NOR2_X1 U875 ( .A1(KEYINPUT6), .A2(n1205), .ZN(n1204) );
XOR2_X1 U876 ( .A(n1206), .B(n1207), .Z(n1205) );
NAND2_X1 U877 ( .A1(n1208), .A2(n1209), .ZN(n1206) );
OR2_X1 U878 ( .A1(n1153), .A2(n1210), .ZN(n1203) );
NAND2_X1 U879 ( .A1(G902), .A2(n1052), .ZN(n1153) );
NAND3_X1 U880 ( .A1(n1116), .A2(n1141), .A3(n1211), .ZN(n1052) );
NOR3_X1 U881 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1211) );
NOR2_X1 U882 ( .A1(n1145), .A2(n1144), .ZN(n1214) );
INV_X1 U883 ( .A(n1146), .ZN(n1213) );
XOR2_X1 U884 ( .A(n1117), .B(KEYINPUT29), .Z(n1212) );
AND4_X1 U885 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1047), .ZN(n1141) );
NAND3_X1 U886 ( .A1(n1079), .A2(n1218), .A3(n1219), .ZN(n1047) );
NAND2_X1 U887 ( .A1(n1068), .A2(n1220), .ZN(n1215) );
NAND3_X1 U888 ( .A1(n1175), .A2(n1221), .A3(n1222), .ZN(n1220) );
XNOR2_X1 U889 ( .A(KEYINPUT35), .B(n1223), .ZN(n1222) );
NAND3_X1 U890 ( .A1(n1080), .A2(n1218), .A3(n1224), .ZN(n1175) );
NOR3_X1 U891 ( .A1(n1076), .A2(n1225), .A3(n1077), .ZN(n1224) );
AND4_X1 U892 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1116) );
NOR4_X1 U893 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1229) );
INV_X1 U894 ( .A(n1234), .ZN(n1231) );
NAND3_X1 U895 ( .A1(n1079), .A2(n1068), .A3(n1235), .ZN(n1228) );
NOR2_X1 U896 ( .A1(n1236), .A2(G952), .ZN(n1148) );
XOR2_X1 U897 ( .A(G953), .B(KEYINPUT22), .Z(n1236) );
XOR2_X1 U898 ( .A(G146), .B(n1233), .Z(G48) );
AND3_X1 U899 ( .A1(n1080), .A2(n1068), .A3(n1235), .ZN(n1233) );
INV_X1 U900 ( .A(n1237), .ZN(n1235) );
XOR2_X1 U901 ( .A(n1238), .B(n1226), .Z(G45) );
NAND3_X1 U902 ( .A1(n1239), .A2(n1074), .A3(n1240), .ZN(n1226) );
NOR3_X1 U903 ( .A1(n1145), .A2(n1082), .A3(n1241), .ZN(n1240) );
XNOR2_X1 U904 ( .A(n1117), .B(n1242), .ZN(G42) );
NOR2_X1 U905 ( .A1(KEYINPUT61), .A2(n1243), .ZN(n1242) );
NAND4_X1 U906 ( .A1(n1244), .A2(n1239), .A3(n1080), .A4(n1073), .ZN(n1117) );
XOR2_X1 U907 ( .A(n1232), .B(n1245), .Z(G39) );
NOR2_X1 U908 ( .A1(KEYINPUT42), .A2(n1246), .ZN(n1245) );
XNOR2_X1 U909 ( .A(G137), .B(KEYINPUT46), .ZN(n1246) );
NOR3_X1 U910 ( .A1(n1072), .A2(n1058), .A3(n1237), .ZN(n1232) );
XNOR2_X1 U911 ( .A(G134), .B(n1227), .ZN(G36) );
NAND4_X1 U912 ( .A1(n1244), .A2(n1239), .A3(n1074), .A4(n1079), .ZN(n1227) );
XOR2_X1 U913 ( .A(n1247), .B(n1234), .Z(G33) );
NAND4_X1 U914 ( .A1(n1244), .A2(n1239), .A3(n1074), .A4(n1080), .ZN(n1234) );
INV_X1 U915 ( .A(n1072), .ZN(n1244) );
NAND2_X1 U916 ( .A1(n1248), .A2(n1070), .ZN(n1072) );
INV_X1 U917 ( .A(n1069), .ZN(n1248) );
XOR2_X1 U918 ( .A(G128), .B(n1249), .Z(G30) );
NOR3_X1 U919 ( .A1(n1237), .A2(n1250), .A3(n1251), .ZN(n1249) );
XOR2_X1 U920 ( .A(n1145), .B(KEYINPUT30), .Z(n1250) );
NAND3_X1 U921 ( .A1(n1252), .A2(n1253), .A3(n1239), .ZN(n1237) );
NOR3_X1 U922 ( .A1(n1254), .A2(n1077), .A3(n1076), .ZN(n1239) );
XOR2_X1 U923 ( .A(n1255), .B(n1216), .Z(G3) );
NAND3_X1 U924 ( .A1(n1256), .A2(n1219), .A3(n1074), .ZN(n1216) );
XNOR2_X1 U925 ( .A(n1230), .B(n1257), .ZN(G27) );
NAND2_X1 U926 ( .A1(KEYINPUT50), .A2(G125), .ZN(n1257) );
AND4_X1 U927 ( .A1(n1080), .A2(n1258), .A3(n1259), .A4(n1073), .ZN(n1230) );
NOR2_X1 U928 ( .A1(n1254), .A2(n1145), .ZN(n1259) );
AND2_X1 U929 ( .A1(n1260), .A2(n1261), .ZN(n1254) );
NAND4_X1 U930 ( .A1(G902), .A2(n1124), .A3(n1262), .A4(n1125), .ZN(n1261) );
INV_X1 U931 ( .A(G900), .ZN(n1125) );
INV_X1 U932 ( .A(n1062), .ZN(n1258) );
XOR2_X1 U933 ( .A(n1263), .B(n1264), .Z(G24) );
NOR2_X1 U934 ( .A1(G122), .A2(KEYINPUT51), .ZN(n1264) );
NAND2_X1 U935 ( .A1(n1068), .A2(n1265), .ZN(n1263) );
XNOR2_X1 U936 ( .A(KEYINPUT11), .B(n1144), .ZN(n1265) );
NAND4_X1 U937 ( .A1(n1266), .A2(n1218), .A3(n1267), .A4(n1268), .ZN(n1144) );
INV_X1 U938 ( .A(n1066), .ZN(n1218) );
NAND2_X1 U939 ( .A1(n1269), .A2(n1270), .ZN(n1066) );
XOR2_X1 U940 ( .A(G119), .B(n1271), .Z(G21) );
NOR2_X1 U941 ( .A1(n1145), .A2(n1223), .ZN(n1271) );
NAND4_X1 U942 ( .A1(n1266), .A2(n1256), .A3(n1252), .A4(n1253), .ZN(n1223) );
XOR2_X1 U943 ( .A(G116), .B(n1272), .Z(G18) );
NOR2_X1 U944 ( .A1(n1273), .A2(n1221), .ZN(n1272) );
NAND3_X1 U945 ( .A1(n1074), .A2(n1079), .A3(n1266), .ZN(n1221) );
INV_X1 U946 ( .A(n1251), .ZN(n1079) );
NAND2_X1 U947 ( .A1(n1274), .A2(n1268), .ZN(n1251) );
XOR2_X1 U948 ( .A(n1275), .B(KEYINPUT5), .Z(n1274) );
XOR2_X1 U949 ( .A(n1145), .B(KEYINPUT39), .Z(n1273) );
XNOR2_X1 U950 ( .A(G113), .B(n1217), .ZN(G15) );
NAND4_X1 U951 ( .A1(n1266), .A2(n1074), .A3(n1080), .A4(n1068), .ZN(n1217) );
INV_X1 U952 ( .A(n1145), .ZN(n1068) );
NOR2_X1 U953 ( .A1(n1268), .A2(n1241), .ZN(n1080) );
INV_X1 U954 ( .A(n1267), .ZN(n1241) );
XNOR2_X1 U955 ( .A(n1275), .B(KEYINPUT7), .ZN(n1267) );
INV_X1 U956 ( .A(n1082), .ZN(n1268) );
AND2_X1 U957 ( .A1(n1269), .A2(n1252), .ZN(n1074) );
NOR2_X1 U958 ( .A1(n1062), .A2(n1225), .ZN(n1266) );
NAND2_X1 U959 ( .A1(n1076), .A2(n1094), .ZN(n1062) );
XOR2_X1 U960 ( .A(n1200), .B(n1146), .Z(G12) );
NAND3_X1 U961 ( .A1(n1073), .A2(n1219), .A3(n1256), .ZN(n1146) );
INV_X1 U962 ( .A(n1058), .ZN(n1256) );
NAND2_X1 U963 ( .A1(n1082), .A2(n1275), .ZN(n1058) );
XNOR2_X1 U964 ( .A(n1107), .B(n1097), .ZN(n1275) );
XNOR2_X1 U965 ( .A(G475), .B(KEYINPUT47), .ZN(n1097) );
NAND2_X1 U966 ( .A1(n1170), .A2(n1161), .ZN(n1107) );
XOR2_X1 U967 ( .A(n1276), .B(n1277), .Z(n1170) );
XOR2_X1 U968 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U969 ( .A(n1280), .B(G104), .Z(n1279) );
NAND2_X1 U970 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND2_X1 U971 ( .A1(G113), .A2(n1283), .ZN(n1282) );
XOR2_X1 U972 ( .A(KEYINPUT49), .B(n1284), .Z(n1281) );
NOR2_X1 U973 ( .A1(G113), .A2(n1283), .ZN(n1284) );
INV_X1 U974 ( .A(G122), .ZN(n1283) );
NAND2_X1 U975 ( .A1(n1285), .A2(n1286), .ZN(n1278) );
OR2_X1 U976 ( .A1(n1287), .A2(G146), .ZN(n1286) );
XOR2_X1 U977 ( .A(n1288), .B(KEYINPUT44), .Z(n1285) );
NAND2_X1 U978 ( .A1(n1289), .A2(n1287), .ZN(n1288) );
XOR2_X1 U979 ( .A(G125), .B(n1123), .Z(n1287) );
XOR2_X1 U980 ( .A(KEYINPUT45), .B(G146), .Z(n1289) );
XOR2_X1 U981 ( .A(n1290), .B(n1291), .Z(n1276) );
NAND2_X1 U982 ( .A1(n1292), .A2(G214), .ZN(n1290) );
XOR2_X1 U983 ( .A(n1293), .B(G478), .Z(n1082) );
NAND2_X1 U984 ( .A1(n1159), .A2(n1161), .ZN(n1293) );
XOR2_X1 U985 ( .A(n1294), .B(n1295), .Z(n1159) );
AND2_X1 U986 ( .A1(n1296), .A2(G217), .ZN(n1295) );
NAND2_X1 U987 ( .A1(n1297), .A2(n1298), .ZN(n1294) );
NAND3_X1 U988 ( .A1(KEYINPUT21), .A2(n1046), .A3(n1299), .ZN(n1298) );
XOR2_X1 U989 ( .A(n1300), .B(n1301), .Z(n1299) );
NOR2_X1 U990 ( .A1(KEYINPUT3), .A2(n1302), .ZN(n1301) );
NAND2_X1 U991 ( .A1(n1303), .A2(n1304), .ZN(n1297) );
NAND2_X1 U992 ( .A1(KEYINPUT21), .A2(n1046), .ZN(n1304) );
INV_X1 U993 ( .A(G107), .ZN(n1046) );
XOR2_X1 U994 ( .A(n1300), .B(n1305), .Z(n1303) );
NOR2_X1 U995 ( .A1(KEYINPUT3), .A2(n1306), .ZN(n1305) );
INV_X1 U996 ( .A(n1302), .ZN(n1306) );
XOR2_X1 U997 ( .A(G116), .B(G122), .Z(n1302) );
XOR2_X1 U998 ( .A(n1307), .B(G134), .Z(n1300) );
NAND3_X1 U999 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1307) );
XNOR2_X1 U1000 ( .A(KEYINPUT27), .B(KEYINPUT2), .ZN(n1310) );
NAND2_X1 U1001 ( .A1(n1311), .A2(n1238), .ZN(n1309) );
INV_X1 U1002 ( .A(G143), .ZN(n1238) );
XOR2_X1 U1003 ( .A(KEYINPUT48), .B(G128), .Z(n1311) );
NAND2_X1 U1004 ( .A1(n1312), .A2(G143), .ZN(n1308) );
XOR2_X1 U1005 ( .A(KEYINPUT15), .B(G128), .Z(n1312) );
NOR4_X1 U1006 ( .A1(n1145), .A2(n1076), .A3(n1077), .A4(n1225), .ZN(n1219) );
AND2_X1 U1007 ( .A1(n1313), .A2(n1260), .ZN(n1225) );
NAND2_X1 U1008 ( .A1(n1314), .A2(n1114), .ZN(n1260) );
INV_X1 U1009 ( .A(n1054), .ZN(n1314) );
NAND2_X1 U1010 ( .A1(G952), .A2(n1262), .ZN(n1054) );
XOR2_X1 U1011 ( .A(KEYINPUT10), .B(n1315), .Z(n1313) );
AND4_X1 U1012 ( .A1(n1136), .A2(n1262), .A3(n1124), .A4(G902), .ZN(n1315) );
XNOR2_X1 U1013 ( .A(n1114), .B(KEYINPUT31), .ZN(n1124) );
NAND2_X1 U1014 ( .A1(n1316), .A2(G237), .ZN(n1262) );
XNOR2_X1 U1015 ( .A(G234), .B(KEYINPUT4), .ZN(n1316) );
INV_X1 U1016 ( .A(G898), .ZN(n1136) );
INV_X1 U1017 ( .A(n1094), .ZN(n1077) );
NAND2_X1 U1018 ( .A1(G221), .A2(n1317), .ZN(n1094) );
XOR2_X1 U1019 ( .A(n1090), .B(n1088), .Z(n1076) );
INV_X1 U1020 ( .A(G469), .ZN(n1088) );
AND3_X1 U1021 ( .A1(n1318), .A2(n1319), .A3(n1161), .ZN(n1090) );
NAND2_X1 U1022 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
INV_X1 U1023 ( .A(KEYINPUT33), .ZN(n1321) );
XOR2_X1 U1024 ( .A(n1322), .B(n1323), .Z(n1320) );
NAND3_X1 U1025 ( .A1(n1322), .A2(n1323), .A3(KEYINPUT33), .ZN(n1318) );
XNOR2_X1 U1026 ( .A(n1120), .B(n1138), .ZN(n1323) );
AND3_X1 U1027 ( .A1(n1324), .A2(n1325), .A3(n1198), .ZN(n1322) );
NAND3_X1 U1028 ( .A1(G110), .A2(n1326), .A3(n1327), .ZN(n1198) );
NAND3_X1 U1029 ( .A1(n1328), .A2(n1200), .A3(n1326), .ZN(n1325) );
XOR2_X1 U1030 ( .A(KEYINPUT17), .B(n1123), .Z(n1328) );
NAND2_X1 U1031 ( .A1(n1329), .A2(n1201), .ZN(n1324) );
INV_X1 U1032 ( .A(n1326), .ZN(n1201) );
NAND2_X1 U1033 ( .A1(G227), .A2(n1114), .ZN(n1326) );
XOR2_X1 U1034 ( .A(n1330), .B(n1123), .Z(n1329) );
NOR2_X1 U1035 ( .A1(G110), .A2(KEYINPUT17), .ZN(n1330) );
NAND2_X1 U1036 ( .A1(n1069), .A2(n1070), .ZN(n1145) );
NAND2_X1 U1037 ( .A1(G214), .A2(n1331), .ZN(n1070) );
NAND3_X1 U1038 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1069) );
NAND2_X1 U1039 ( .A1(n1109), .A2(n1108), .ZN(n1334) );
NAND2_X1 U1040 ( .A1(KEYINPUT1), .A2(n1335), .ZN(n1333) );
NAND2_X1 U1041 ( .A1(n1336), .A2(n1210), .ZN(n1335) );
XOR2_X1 U1042 ( .A(n1108), .B(KEYINPUT63), .Z(n1336) );
NAND2_X1 U1043 ( .A1(n1337), .A2(n1338), .ZN(n1332) );
INV_X1 U1044 ( .A(KEYINPUT1), .ZN(n1338) );
NAND2_X1 U1045 ( .A1(n1339), .A2(n1340), .ZN(n1337) );
NAND2_X1 U1046 ( .A1(n1108), .A2(n1341), .ZN(n1340) );
OR3_X1 U1047 ( .A1(n1108), .A2(n1109), .A3(n1341), .ZN(n1339) );
INV_X1 U1048 ( .A(KEYINPUT63), .ZN(n1341) );
INV_X1 U1049 ( .A(n1210), .ZN(n1109) );
NAND2_X1 U1050 ( .A1(G210), .A2(n1331), .ZN(n1210) );
NAND2_X1 U1051 ( .A1(n1342), .A2(n1161), .ZN(n1331) );
INV_X1 U1052 ( .A(G237), .ZN(n1342) );
NAND2_X1 U1053 ( .A1(n1343), .A2(n1161), .ZN(n1108) );
XOR2_X1 U1054 ( .A(n1207), .B(n1344), .Z(n1343) );
XOR2_X1 U1055 ( .A(KEYINPUT43), .B(n1345), .Z(n1344) );
NOR3_X1 U1056 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1345) );
AND2_X1 U1057 ( .A1(n1349), .A2(KEYINPUT28), .ZN(n1348) );
NOR2_X1 U1058 ( .A1(KEYINPUT28), .A2(n1209), .ZN(n1347) );
NAND3_X1 U1059 ( .A1(G224), .A2(n1114), .A3(n1350), .ZN(n1209) );
INV_X1 U1060 ( .A(n1349), .ZN(n1350) );
INV_X1 U1061 ( .A(n1208), .ZN(n1346) );
NAND2_X1 U1062 ( .A1(n1349), .A2(n1351), .ZN(n1208) );
NAND2_X1 U1063 ( .A1(G224), .A2(n1114), .ZN(n1351) );
XOR2_X1 U1064 ( .A(n1352), .B(G143), .Z(n1349) );
XOR2_X1 U1065 ( .A(n1353), .B(n1354), .Z(n1207) );
INV_X1 U1066 ( .A(n1137), .ZN(n1354) );
XOR2_X1 U1067 ( .A(n1355), .B(n1356), .Z(n1137) );
XOR2_X1 U1068 ( .A(G122), .B(G113), .Z(n1356) );
XOR2_X1 U1069 ( .A(n1200), .B(n1357), .Z(n1355) );
NAND2_X1 U1070 ( .A1(KEYINPUT24), .A2(n1138), .ZN(n1353) );
XOR2_X1 U1071 ( .A(G101), .B(n1358), .Z(n1138) );
XOR2_X1 U1072 ( .A(G107), .B(G104), .Z(n1358) );
AND2_X1 U1073 ( .A1(n1270), .A2(n1253), .ZN(n1073) );
INV_X1 U1074 ( .A(n1269), .ZN(n1253) );
XNOR2_X1 U1075 ( .A(n1359), .B(n1093), .ZN(n1269) );
NAND2_X1 U1076 ( .A1(G217), .A2(n1317), .ZN(n1093) );
NAND2_X1 U1077 ( .A1(G234), .A2(n1161), .ZN(n1317) );
XNOR2_X1 U1078 ( .A(n1092), .B(KEYINPUT14), .ZN(n1359) );
NOR2_X1 U1079 ( .A1(n1155), .A2(G902), .ZN(n1092) );
INV_X1 U1080 ( .A(n1152), .ZN(n1155) );
XOR2_X1 U1081 ( .A(n1360), .B(n1361), .Z(n1152) );
XOR2_X1 U1082 ( .A(n1352), .B(n1123), .Z(n1361) );
INV_X1 U1083 ( .A(n1327), .ZN(n1123) );
XOR2_X1 U1084 ( .A(n1243), .B(KEYINPUT12), .Z(n1327) );
INV_X1 U1085 ( .A(G140), .ZN(n1243) );
XOR2_X1 U1086 ( .A(G125), .B(n1192), .Z(n1352) );
XOR2_X1 U1087 ( .A(n1362), .B(n1363), .Z(n1360) );
NOR2_X1 U1088 ( .A1(KEYINPUT57), .A2(n1364), .ZN(n1363) );
XNOR2_X1 U1089 ( .A(G137), .B(n1365), .ZN(n1364) );
NAND2_X1 U1090 ( .A1(n1296), .A2(G221), .ZN(n1365) );
AND2_X1 U1091 ( .A1(G234), .A2(n1114), .ZN(n1296) );
INV_X1 U1092 ( .A(G953), .ZN(n1114) );
XOR2_X1 U1093 ( .A(G119), .B(n1200), .Z(n1362) );
XOR2_X1 U1094 ( .A(n1252), .B(KEYINPUT8), .Z(n1270) );
XNOR2_X1 U1095 ( .A(n1103), .B(G472), .ZN(n1252) );
NAND2_X1 U1096 ( .A1(n1366), .A2(n1161), .ZN(n1103) );
INV_X1 U1097 ( .A(G902), .ZN(n1161) );
XOR2_X1 U1098 ( .A(n1367), .B(n1368), .Z(n1366) );
XOR2_X1 U1099 ( .A(n1120), .B(n1369), .Z(n1368) );
XOR2_X1 U1100 ( .A(n1183), .B(n1370), .Z(n1369) );
NOR2_X1 U1101 ( .A1(KEYINPUT20), .A2(n1255), .ZN(n1370) );
INV_X1 U1102 ( .A(G101), .ZN(n1255) );
NAND2_X1 U1103 ( .A1(n1292), .A2(G210), .ZN(n1183) );
NOR2_X1 U1104 ( .A1(G953), .A2(G237), .ZN(n1292) );
XNOR2_X1 U1105 ( .A(n1291), .B(n1371), .ZN(n1120) );
XOR2_X1 U1106 ( .A(n1191), .B(n1192), .Z(n1371) );
XNOR2_X1 U1107 ( .A(n1372), .B(G146), .ZN(n1192) );
INV_X1 U1108 ( .A(G128), .ZN(n1372) );
XOR2_X1 U1109 ( .A(G134), .B(G137), .Z(n1191) );
XNOR2_X1 U1110 ( .A(n1247), .B(G143), .ZN(n1291) );
INV_X1 U1111 ( .A(G131), .ZN(n1247) );
XOR2_X1 U1112 ( .A(n1373), .B(n1374), .Z(n1367) );
XOR2_X1 U1113 ( .A(KEYINPUT53), .B(KEYINPUT26), .Z(n1374) );
NOR2_X1 U1114 ( .A1(KEYINPUT32), .A2(n1179), .ZN(n1373) );
XOR2_X1 U1115 ( .A(n1357), .B(n1375), .Z(n1179) );
NOR2_X1 U1116 ( .A1(G113), .A2(KEYINPUT58), .ZN(n1375) );
XOR2_X1 U1117 ( .A(G116), .B(G119), .Z(n1357) );
INV_X1 U1118 ( .A(G110), .ZN(n1200) );
endmodule


