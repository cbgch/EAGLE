//Key = 1111000110100001001010111001101011100100001001110110011101010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306;

XOR2_X1 U724 ( .A(n991), .B(n992), .Z(G9) );
XNOR2_X1 U725 ( .A(G107), .B(KEYINPUT16), .ZN(n992) );
NOR2_X1 U726 ( .A1(n993), .A2(n994), .ZN(G75) );
NOR4_X1 U727 ( .A1(n995), .A2(n996), .A3(n997), .A4(n998), .ZN(n994) );
NOR2_X1 U728 ( .A1(n999), .A2(n1000), .ZN(n998) );
XNOR2_X1 U729 ( .A(KEYINPUT33), .B(n1001), .ZN(n1000) );
NOR3_X1 U730 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n997) );
NAND4_X1 U731 ( .A1(n1004), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n1001) );
NAND3_X1 U732 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n995) );
NAND3_X1 U733 ( .A1(n1011), .A2(n1012), .A3(n1004), .ZN(n1010) );
INV_X1 U734 ( .A(n1013), .ZN(n1004) );
NAND2_X1 U735 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NAND3_X1 U736 ( .A1(n1007), .A2(n1016), .A3(n1005), .ZN(n1015) );
OR2_X1 U737 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND2_X1 U738 ( .A1(n1006), .A2(n1019), .ZN(n1014) );
NAND2_X1 U739 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U740 ( .A1(n1007), .A2(n1022), .ZN(n1021) );
NAND2_X1 U741 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U742 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U743 ( .A1(n1005), .A2(n1027), .ZN(n1020) );
OR2_X1 U744 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR3_X1 U745 ( .A1(n1030), .A2(G953), .A3(G952), .ZN(n993) );
INV_X1 U746 ( .A(n1008), .ZN(n1030) );
NAND4_X1 U747 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1008) );
NOR4_X1 U748 ( .A1(n1025), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1034) );
XOR2_X1 U749 ( .A(n1038), .B(KEYINPUT62), .Z(n1037) );
NOR2_X1 U750 ( .A1(n1039), .A2(n1040), .ZN(n1033) );
XNOR2_X1 U751 ( .A(KEYINPUT9), .B(n1041), .ZN(n1040) );
INV_X1 U752 ( .A(n1007), .ZN(n1039) );
XOR2_X1 U753 ( .A(n1042), .B(G469), .Z(n1032) );
XOR2_X1 U754 ( .A(n1043), .B(n1044), .Z(n1031) );
NAND2_X1 U755 ( .A1(n1045), .A2(n1046), .ZN(G72) );
NAND2_X1 U756 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U757 ( .A1(n1049), .A2(n1050), .ZN(n1045) );
NAND2_X1 U758 ( .A1(n1051), .A2(n1048), .ZN(n1050) );
NAND2_X1 U759 ( .A1(G953), .A2(n1052), .ZN(n1048) );
INV_X1 U760 ( .A(G227), .ZN(n1052) );
INV_X1 U761 ( .A(n1047), .ZN(n1049) );
XNOR2_X1 U762 ( .A(n1053), .B(n1054), .ZN(n1047) );
NOR2_X1 U763 ( .A1(n1055), .A2(G953), .ZN(n1054) );
NOR2_X1 U764 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U765 ( .A1(n1058), .A2(n1051), .ZN(n1053) );
INV_X1 U766 ( .A(n1059), .ZN(n1051) );
XOR2_X1 U767 ( .A(n1060), .B(n1061), .Z(n1058) );
NAND2_X1 U768 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
XNOR2_X1 U769 ( .A(n1064), .B(n1065), .ZN(n1063) );
NAND2_X1 U770 ( .A1(KEYINPUT22), .A2(n1066), .ZN(n1064) );
XNOR2_X1 U771 ( .A(KEYINPUT61), .B(KEYINPUT39), .ZN(n1062) );
XOR2_X1 U772 ( .A(n1067), .B(n1068), .Z(G69) );
XOR2_X1 U773 ( .A(n1069), .B(n1070), .Z(n1068) );
NOR2_X1 U774 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XOR2_X1 U775 ( .A(KEYINPUT36), .B(n1073), .Z(n1072) );
NOR3_X1 U776 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
XNOR2_X1 U777 ( .A(n1077), .B(KEYINPUT0), .ZN(n1075) );
XNOR2_X1 U778 ( .A(G953), .B(KEYINPUT49), .ZN(n1071) );
NOR2_X1 U779 ( .A1(KEYINPUT4), .A2(n1078), .ZN(n1069) );
NOR2_X1 U780 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U781 ( .A(KEYINPUT40), .B(n1081), .Z(n1080) );
NOR3_X1 U782 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NOR2_X1 U783 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U784 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR4_X1 U785 ( .A1(n1089), .A2(n1088), .A3(KEYINPUT13), .A4(n1087), .ZN(n1083) );
INV_X1 U786 ( .A(KEYINPUT37), .ZN(n1088) );
INV_X1 U787 ( .A(n1086), .ZN(n1089) );
AND2_X1 U788 ( .A1(n1087), .A2(KEYINPUT13), .ZN(n1082) );
XNOR2_X1 U789 ( .A(n1090), .B(n1091), .ZN(n1087) );
NAND2_X1 U790 ( .A1(KEYINPUT59), .A2(n1092), .ZN(n1090) );
NOR2_X1 U791 ( .A1(G898), .A2(n1093), .ZN(n1079) );
XNOR2_X1 U792 ( .A(KEYINPUT32), .B(n1009), .ZN(n1093) );
NAND2_X1 U793 ( .A1(G953), .A2(n1094), .ZN(n1067) );
NAND2_X1 U794 ( .A1(G898), .A2(G224), .ZN(n1094) );
NOR2_X1 U795 ( .A1(n1095), .A2(n1096), .ZN(G66) );
XOR2_X1 U796 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U797 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NOR2_X1 U798 ( .A1(n1095), .A2(n1101), .ZN(G63) );
XOR2_X1 U799 ( .A(n1102), .B(n1103), .Z(n1101) );
AND2_X1 U800 ( .A1(G478), .A2(n1104), .ZN(n1102) );
NOR3_X1 U801 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(G60) );
NOR3_X1 U802 ( .A1(n1108), .A2(G953), .A3(G952), .ZN(n1107) );
AND2_X1 U803 ( .A1(n1108), .A2(n1095), .ZN(n1106) );
INV_X1 U804 ( .A(KEYINPUT48), .ZN(n1108) );
XOR2_X1 U805 ( .A(n1109), .B(n1110), .Z(n1105) );
NOR2_X1 U806 ( .A1(KEYINPUT11), .A2(n1111), .ZN(n1110) );
AND2_X1 U807 ( .A1(G475), .A2(n1104), .ZN(n1109) );
XNOR2_X1 U808 ( .A(G104), .B(n1112), .ZN(G6) );
NOR2_X1 U809 ( .A1(n1095), .A2(n1113), .ZN(G57) );
NOR2_X1 U810 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U811 ( .A(KEYINPUT14), .B(n1116), .Z(n1115) );
NOR2_X1 U812 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XNOR2_X1 U813 ( .A(n1119), .B(n1120), .ZN(n1118) );
INV_X1 U814 ( .A(n1121), .ZN(n1117) );
NOR2_X1 U815 ( .A1(n1122), .A2(n1121), .ZN(n1114) );
XOR2_X1 U816 ( .A(G101), .B(n1123), .Z(n1121) );
NOR2_X1 U817 ( .A1(KEYINPUT21), .A2(n1124), .ZN(n1123) );
XNOR2_X1 U818 ( .A(n1125), .B(n1120), .ZN(n1122) );
XNOR2_X1 U819 ( .A(n1126), .B(n1127), .ZN(n1120) );
NOR2_X1 U820 ( .A1(KEYINPUT6), .A2(n1128), .ZN(n1127) );
NAND2_X1 U821 ( .A1(n1104), .A2(G472), .ZN(n1126) );
NOR2_X1 U822 ( .A1(n1095), .A2(n1129), .ZN(G54) );
XOR2_X1 U823 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U824 ( .A(n1132), .B(n1133), .Z(n1131) );
XNOR2_X1 U825 ( .A(n1134), .B(n1135), .ZN(n1130) );
XOR2_X1 U826 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U827 ( .A1(n1138), .A2(KEYINPUT3), .ZN(n1137) );
XNOR2_X1 U828 ( .A(G134), .B(n1139), .ZN(n1138) );
NAND3_X1 U829 ( .A1(n1140), .A2(n996), .A3(G469), .ZN(n1136) );
XNOR2_X1 U830 ( .A(KEYINPUT58), .B(n1141), .ZN(n1140) );
NOR2_X1 U831 ( .A1(n1009), .A2(G952), .ZN(n1095) );
NOR2_X1 U832 ( .A1(n1142), .A2(n1143), .ZN(G51) );
XOR2_X1 U833 ( .A(n1144), .B(n1145), .Z(n1143) );
NOR2_X1 U834 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U835 ( .A(n1148), .B(KEYINPUT45), .Z(n1147) );
NAND2_X1 U836 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U837 ( .A1(n1149), .A2(n1150), .ZN(n1146) );
XNOR2_X1 U838 ( .A(n1134), .B(n1151), .ZN(n1150) );
NAND2_X1 U839 ( .A1(KEYINPUT34), .A2(n1152), .ZN(n1144) );
NAND2_X1 U840 ( .A1(n1104), .A2(n1044), .ZN(n1152) );
INV_X1 U841 ( .A(n1100), .ZN(n1104) );
NAND2_X1 U842 ( .A1(G902), .A2(n996), .ZN(n1100) );
NAND4_X1 U843 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n996) );
INV_X1 U844 ( .A(n1074), .ZN(n1156) );
NAND3_X1 U845 ( .A1(n1112), .A2(n991), .A3(n1157), .ZN(n1074) );
NAND4_X1 U846 ( .A1(n1028), .A2(n1006), .A3(n1158), .A4(n1159), .ZN(n1157) );
OR2_X1 U847 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U848 ( .A1(n1162), .A2(n1160), .ZN(n1158) );
INV_X1 U849 ( .A(KEYINPUT8), .ZN(n1160) );
NAND3_X1 U850 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1162) );
NAND3_X1 U851 ( .A1(n1018), .A2(n1007), .A3(n1161), .ZN(n991) );
NAND3_X1 U852 ( .A1(n1161), .A2(n1007), .A3(n1017), .ZN(n1112) );
NOR2_X1 U853 ( .A1(n1077), .A2(n1057), .ZN(n1155) );
NAND4_X1 U854 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1057) );
AND4_X1 U855 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1169) );
NAND4_X1 U856 ( .A1(n1174), .A2(n1175), .A3(n1165), .A4(n1176), .ZN(n1168) );
XNOR2_X1 U857 ( .A(n1011), .B(KEYINPUT20), .ZN(n1174) );
NAND2_X1 U858 ( .A1(n1177), .A2(n1178), .ZN(n1166) );
INV_X1 U859 ( .A(n1179), .ZN(n1178) );
XNOR2_X1 U860 ( .A(n1029), .B(KEYINPUT42), .ZN(n1177) );
INV_X1 U861 ( .A(n1180), .ZN(n1077) );
XOR2_X1 U862 ( .A(n1076), .B(KEYINPUT53), .Z(n1154) );
NAND4_X1 U863 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1076) );
XNOR2_X1 U864 ( .A(n1056), .B(KEYINPUT17), .ZN(n1153) );
INV_X1 U865 ( .A(n1185), .ZN(n1056) );
NOR2_X1 U866 ( .A1(G952), .A2(n1186), .ZN(n1142) );
XNOR2_X1 U867 ( .A(G953), .B(KEYINPUT12), .ZN(n1186) );
XNOR2_X1 U868 ( .A(n1187), .B(n1188), .ZN(G48) );
NAND2_X1 U869 ( .A1(n1189), .A2(n1190), .ZN(n1187) );
OR2_X1 U870 ( .A1(n1185), .A2(KEYINPUT19), .ZN(n1190) );
NAND3_X1 U871 ( .A1(n1191), .A2(n1017), .A3(n1192), .ZN(n1185) );
NAND4_X1 U872 ( .A1(n1017), .A2(n1193), .A3(n1192), .A4(KEYINPUT19), .ZN(n1189) );
XOR2_X1 U873 ( .A(G143), .B(n1194), .Z(G45) );
NOR2_X1 U874 ( .A1(n1195), .A2(n1179), .ZN(n1194) );
NAND3_X1 U875 ( .A1(n1196), .A2(n1197), .A3(n1192), .ZN(n1179) );
XNOR2_X1 U876 ( .A(G140), .B(n1167), .ZN(G42) );
NAND3_X1 U877 ( .A1(n1028), .A2(n1017), .A3(n1198), .ZN(n1167) );
XOR2_X1 U878 ( .A(n1199), .B(n1200), .Z(G39) );
NAND2_X1 U879 ( .A1(n1175), .A2(n1198), .ZN(n1200) );
NAND2_X1 U880 ( .A1(KEYINPUT2), .A2(G137), .ZN(n1199) );
XOR2_X1 U881 ( .A(n1173), .B(n1201), .Z(G36) );
XNOR2_X1 U882 ( .A(G134), .B(KEYINPUT41), .ZN(n1201) );
NAND3_X1 U883 ( .A1(n1029), .A2(n1018), .A3(n1198), .ZN(n1173) );
XNOR2_X1 U884 ( .A(G131), .B(n1172), .ZN(G33) );
NAND3_X1 U885 ( .A1(n1017), .A2(n1029), .A3(n1198), .ZN(n1172) );
AND3_X1 U886 ( .A1(n1165), .A2(n1176), .A3(n1011), .ZN(n1198) );
NOR2_X1 U887 ( .A1(n1002), .A2(n1036), .ZN(n1011) );
INV_X1 U888 ( .A(n1003), .ZN(n1036) );
XNOR2_X1 U889 ( .A(G128), .B(n1171), .ZN(G30) );
NAND3_X1 U890 ( .A1(n1191), .A2(n1018), .A3(n1192), .ZN(n1171) );
NOR3_X1 U891 ( .A1(n999), .A2(n1202), .A3(n1023), .ZN(n1192) );
XNOR2_X1 U892 ( .A(G101), .B(n1180), .ZN(G3) );
NAND3_X1 U893 ( .A1(n1029), .A2(n1161), .A3(n1006), .ZN(n1180) );
XNOR2_X1 U894 ( .A(G125), .B(n1170), .ZN(G27) );
NAND4_X1 U895 ( .A1(n1005), .A2(n1028), .A3(n1203), .A4(n1017), .ZN(n1170) );
NOR2_X1 U896 ( .A1(n1202), .A2(n999), .ZN(n1203) );
INV_X1 U897 ( .A(n1176), .ZN(n1202) );
NAND2_X1 U898 ( .A1(n1013), .A2(n1204), .ZN(n1176) );
NAND3_X1 U899 ( .A1(G902), .A2(n1205), .A3(n1059), .ZN(n1204) );
NOR2_X1 U900 ( .A1(G900), .A2(n1009), .ZN(n1059) );
NAND2_X1 U901 ( .A1(n1206), .A2(n1207), .ZN(G24) );
NAND2_X1 U902 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XOR2_X1 U903 ( .A(KEYINPUT7), .B(n1210), .Z(n1206) );
NOR2_X1 U904 ( .A1(n1208), .A2(n1209), .ZN(n1210) );
INV_X1 U905 ( .A(n1181), .ZN(n1208) );
NAND4_X1 U906 ( .A1(n1211), .A2(n1007), .A3(n1196), .A4(n1197), .ZN(n1181) );
NOR2_X1 U907 ( .A1(n1212), .A2(n1213), .ZN(n1007) );
XNOR2_X1 U908 ( .A(G119), .B(n1182), .ZN(G21) );
NAND2_X1 U909 ( .A1(n1211), .A2(n1175), .ZN(n1182) );
AND2_X1 U910 ( .A1(n1191), .A2(n1006), .ZN(n1175) );
INV_X1 U911 ( .A(n1193), .ZN(n1191) );
NAND2_X1 U912 ( .A1(n1213), .A2(n1212), .ZN(n1193) );
XOR2_X1 U913 ( .A(n1183), .B(n1214), .Z(G18) );
XOR2_X1 U914 ( .A(KEYINPUT57), .B(G116), .Z(n1214) );
NAND3_X1 U915 ( .A1(n1029), .A2(n1018), .A3(n1211), .ZN(n1183) );
NOR3_X1 U916 ( .A1(n999), .A2(n1215), .A3(n1216), .ZN(n1211) );
XOR2_X1 U917 ( .A(n1164), .B(KEYINPUT56), .Z(n999) );
AND2_X1 U918 ( .A1(n1041), .A2(n1197), .ZN(n1018) );
XNOR2_X1 U919 ( .A(G113), .B(n1184), .ZN(G15) );
NAND4_X1 U920 ( .A1(n1005), .A2(n1017), .A3(n1217), .A4(n1029), .ZN(n1184) );
INV_X1 U921 ( .A(n1195), .ZN(n1029) );
NAND2_X1 U922 ( .A1(n1218), .A2(n1212), .ZN(n1195) );
NOR2_X1 U923 ( .A1(n1215), .A2(n1164), .ZN(n1217) );
NOR2_X1 U924 ( .A1(n1197), .A2(n1041), .ZN(n1017) );
INV_X1 U925 ( .A(n1196), .ZN(n1041) );
INV_X1 U926 ( .A(n1216), .ZN(n1005) );
NAND2_X1 U927 ( .A1(n1219), .A2(n1026), .ZN(n1216) );
XOR2_X1 U928 ( .A(KEYINPUT46), .B(n1025), .Z(n1219) );
XNOR2_X1 U929 ( .A(G110), .B(n1220), .ZN(G12) );
NAND3_X1 U930 ( .A1(n1006), .A2(n1161), .A3(n1028), .ZN(n1220) );
NOR2_X1 U931 ( .A1(n1212), .A2(n1218), .ZN(n1028) );
INV_X1 U932 ( .A(n1213), .ZN(n1218) );
XOR2_X1 U933 ( .A(n1221), .B(n1099), .Z(n1213) );
NAND2_X1 U934 ( .A1(G217), .A2(n1222), .ZN(n1099) );
OR2_X1 U935 ( .A1(n1098), .A2(G902), .ZN(n1221) );
XNOR2_X1 U936 ( .A(n1223), .B(n1224), .ZN(n1098) );
XOR2_X1 U937 ( .A(n1225), .B(n1226), .Z(n1224) );
XNOR2_X1 U938 ( .A(n1227), .B(n1228), .ZN(n1226) );
NAND2_X1 U939 ( .A1(KEYINPUT23), .A2(n1188), .ZN(n1228) );
NAND2_X1 U940 ( .A1(KEYINPUT18), .A2(G140), .ZN(n1227) );
NAND2_X1 U941 ( .A1(n1229), .A2(G221), .ZN(n1225) );
XOR2_X1 U942 ( .A(n1230), .B(n1231), .Z(n1223) );
XNOR2_X1 U943 ( .A(G137), .B(n1232), .ZN(n1231) );
XOR2_X1 U944 ( .A(n1233), .B(G110), .Z(n1230) );
NAND2_X1 U945 ( .A1(KEYINPUT1), .A2(n1234), .ZN(n1233) );
XOR2_X1 U946 ( .A(G128), .B(G119), .Z(n1234) );
XNOR2_X1 U947 ( .A(n1235), .B(G472), .ZN(n1212) );
NAND2_X1 U948 ( .A1(n1236), .A2(n1141), .ZN(n1235) );
XOR2_X1 U949 ( .A(n1237), .B(n1238), .Z(n1236) );
XNOR2_X1 U950 ( .A(n1119), .B(n1128), .ZN(n1238) );
XOR2_X1 U951 ( .A(n1239), .B(n1240), .Z(n1128) );
NOR2_X1 U952 ( .A1(G113), .A2(KEYINPUT51), .ZN(n1240) );
INV_X1 U953 ( .A(n1125), .ZN(n1119) );
XOR2_X1 U954 ( .A(n1124), .B(n1241), .Z(n1237) );
XNOR2_X1 U955 ( .A(KEYINPUT43), .B(n1242), .ZN(n1241) );
NAND2_X1 U956 ( .A1(n1243), .A2(G210), .ZN(n1124) );
NOR3_X1 U957 ( .A1(n1023), .A2(n1215), .A3(n1164), .ZN(n1161) );
NAND2_X1 U958 ( .A1(n1002), .A2(n1003), .ZN(n1164) );
NAND2_X1 U959 ( .A1(G214), .A2(n1244), .ZN(n1003) );
XOR2_X1 U960 ( .A(n1245), .B(n1246), .Z(n1002) );
XOR2_X1 U961 ( .A(KEYINPUT35), .B(n1044), .Z(n1246) );
AND2_X1 U962 ( .A1(G210), .A2(n1244), .ZN(n1044) );
NAND2_X1 U963 ( .A1(n1247), .A2(n1141), .ZN(n1244) );
INV_X1 U964 ( .A(G237), .ZN(n1247) );
NAND2_X1 U965 ( .A1(KEYINPUT30), .A2(n1043), .ZN(n1245) );
NAND2_X1 U966 ( .A1(n1248), .A2(n1141), .ZN(n1043) );
XOR2_X1 U967 ( .A(n1149), .B(n1249), .Z(n1248) );
XOR2_X1 U968 ( .A(KEYINPUT31), .B(n1250), .Z(n1249) );
NOR3_X1 U969 ( .A1(KEYINPUT44), .A2(n1251), .A3(n1252), .ZN(n1250) );
NOR2_X1 U970 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
XOR2_X1 U971 ( .A(KEYINPUT28), .B(n1151), .Z(n1254) );
INV_X1 U972 ( .A(n1134), .ZN(n1253) );
NOR2_X1 U973 ( .A1(n1151), .A2(n1134), .ZN(n1251) );
XNOR2_X1 U974 ( .A(n1232), .B(n1255), .ZN(n1151) );
AND2_X1 U975 ( .A1(n1009), .A2(G224), .ZN(n1255) );
INV_X1 U976 ( .A(G125), .ZN(n1232) );
XNOR2_X1 U977 ( .A(n1256), .B(n1086), .ZN(n1149) );
XOR2_X1 U978 ( .A(G110), .B(n1209), .Z(n1086) );
XNOR2_X1 U979 ( .A(n1092), .B(n1091), .ZN(n1256) );
XOR2_X1 U980 ( .A(G113), .B(n1239), .Z(n1091) );
XOR2_X1 U981 ( .A(G116), .B(G119), .Z(n1239) );
XOR2_X1 U982 ( .A(n1257), .B(n1242), .Z(n1092) );
INV_X1 U983 ( .A(G101), .ZN(n1242) );
NAND3_X1 U984 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1257) );
OR2_X1 U985 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
NAND3_X1 U986 ( .A1(n1262), .A2(n1261), .A3(KEYINPUT47), .ZN(n1259) );
NOR2_X1 U987 ( .A1(KEYINPUT38), .A2(n1263), .ZN(n1262) );
NAND2_X1 U988 ( .A1(n1263), .A2(n1264), .ZN(n1258) );
INV_X1 U989 ( .A(KEYINPUT47), .ZN(n1264) );
INV_X1 U990 ( .A(n1163), .ZN(n1215) );
NAND2_X1 U991 ( .A1(n1013), .A2(n1265), .ZN(n1163) );
NAND4_X1 U992 ( .A1(G953), .A2(G902), .A3(n1205), .A4(n1266), .ZN(n1265) );
INV_X1 U993 ( .A(G898), .ZN(n1266) );
NAND3_X1 U994 ( .A1(n1205), .A2(n1009), .A3(G952), .ZN(n1013) );
NAND2_X1 U995 ( .A1(G237), .A2(G234), .ZN(n1205) );
INV_X1 U996 ( .A(n1165), .ZN(n1023) );
NOR2_X1 U997 ( .A1(n1026), .A2(n1267), .ZN(n1165) );
XNOR2_X1 U998 ( .A(KEYINPUT46), .B(n1025), .ZN(n1267) );
AND2_X1 U999 ( .A1(G221), .A2(n1222), .ZN(n1025) );
NAND2_X1 U1000 ( .A1(G234), .A2(n1141), .ZN(n1222) );
XNOR2_X1 U1001 ( .A(n1042), .B(n1268), .ZN(n1026) );
NOR2_X1 U1002 ( .A1(G469), .A2(KEYINPUT52), .ZN(n1268) );
NAND2_X1 U1003 ( .A1(n1269), .A2(n1141), .ZN(n1042) );
XOR2_X1 U1004 ( .A(n1132), .B(n1270), .Z(n1269) );
XNOR2_X1 U1005 ( .A(n1271), .B(n1125), .ZN(n1270) );
XOR2_X1 U1006 ( .A(G134), .B(n1065), .Z(n1125) );
XNOR2_X1 U1007 ( .A(n1139), .B(n1134), .ZN(n1065) );
XOR2_X1 U1008 ( .A(G146), .B(n1272), .Z(n1134) );
XOR2_X1 U1009 ( .A(G131), .B(G137), .Z(n1139) );
NAND2_X1 U1010 ( .A1(KEYINPUT24), .A2(n1133), .ZN(n1271) );
XNOR2_X1 U1011 ( .A(n1273), .B(n1274), .ZN(n1133) );
XOR2_X1 U1012 ( .A(G140), .B(G110), .Z(n1274) );
NAND2_X1 U1013 ( .A1(G227), .A2(n1009), .ZN(n1273) );
XNOR2_X1 U1014 ( .A(n1275), .B(G101), .ZN(n1132) );
NAND2_X1 U1015 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND2_X1 U1016 ( .A1(KEYINPUT27), .A2(n1278), .ZN(n1277) );
NAND2_X1 U1017 ( .A1(KEYINPUT29), .A2(n1279), .ZN(n1276) );
INV_X1 U1018 ( .A(n1278), .ZN(n1279) );
NAND3_X1 U1019 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1278) );
OR2_X1 U1020 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NAND3_X1 U1021 ( .A1(n1284), .A2(n1283), .A3(KEYINPUT10), .ZN(n1281) );
XNOR2_X1 U1022 ( .A(n1263), .B(KEYINPUT25), .ZN(n1283) );
NOR2_X1 U1023 ( .A1(G104), .A2(KEYINPUT5), .ZN(n1284) );
OR2_X1 U1024 ( .A1(n1261), .A2(KEYINPUT10), .ZN(n1280) );
INV_X1 U1025 ( .A(G104), .ZN(n1261) );
NOR2_X1 U1026 ( .A1(n1197), .A2(n1196), .ZN(n1006) );
XNOR2_X1 U1027 ( .A(n1285), .B(G475), .ZN(n1196) );
NAND2_X1 U1028 ( .A1(n1111), .A2(n1141), .ZN(n1285) );
INV_X1 U1029 ( .A(G902), .ZN(n1141) );
XNOR2_X1 U1030 ( .A(n1286), .B(n1287), .ZN(n1111) );
XOR2_X1 U1031 ( .A(n1288), .B(n1061), .Z(n1287) );
XNOR2_X1 U1032 ( .A(G125), .B(G140), .ZN(n1061) );
NAND2_X1 U1033 ( .A1(n1289), .A2(KEYINPUT50), .ZN(n1288) );
XOR2_X1 U1034 ( .A(n1290), .B(n1291), .Z(n1289) );
NOR2_X1 U1035 ( .A1(G143), .A2(KEYINPUT60), .ZN(n1291) );
XOR2_X1 U1036 ( .A(n1292), .B(G131), .Z(n1290) );
NAND2_X1 U1037 ( .A1(n1243), .A2(G214), .ZN(n1292) );
NOR2_X1 U1038 ( .A1(G953), .A2(G237), .ZN(n1243) );
XOR2_X1 U1039 ( .A(n1293), .B(n1294), .Z(n1286) );
XNOR2_X1 U1040 ( .A(n1188), .B(G104), .ZN(n1294) );
INV_X1 U1041 ( .A(G146), .ZN(n1188) );
NAND2_X1 U1042 ( .A1(n1295), .A2(KEYINPUT55), .ZN(n1293) );
XNOR2_X1 U1043 ( .A(G122), .B(n1296), .ZN(n1295) );
NOR2_X1 U1044 ( .A1(G113), .A2(KEYINPUT26), .ZN(n1296) );
NAND2_X1 U1045 ( .A1(n1297), .A2(n1038), .ZN(n1197) );
NAND2_X1 U1046 ( .A1(G478), .A2(n1298), .ZN(n1038) );
OR2_X1 U1047 ( .A1(n1103), .A2(G902), .ZN(n1298) );
XNOR2_X1 U1048 ( .A(n1035), .B(KEYINPUT63), .ZN(n1297) );
NOR3_X1 U1049 ( .A1(G478), .A2(G902), .A3(n1103), .ZN(n1035) );
XNOR2_X1 U1050 ( .A(n1299), .B(n1300), .ZN(n1103) );
XOR2_X1 U1051 ( .A(n1301), .B(n1263), .Z(n1300) );
XNOR2_X1 U1052 ( .A(G107), .B(KEYINPUT54), .ZN(n1263) );
NAND2_X1 U1053 ( .A1(G217), .A2(n1229), .ZN(n1301) );
AND2_X1 U1054 ( .A1(G234), .A2(n1009), .ZN(n1229) );
INV_X1 U1055 ( .A(G953), .ZN(n1009) );
XOR2_X1 U1056 ( .A(n1302), .B(n1303), .Z(n1299) );
XNOR2_X1 U1057 ( .A(n1209), .B(G116), .ZN(n1303) );
INV_X1 U1058 ( .A(G122), .ZN(n1209) );
NAND2_X1 U1059 ( .A1(n1304), .A2(n1305), .ZN(n1302) );
NAND2_X1 U1060 ( .A1(n1272), .A2(n1066), .ZN(n1305) );
XOR2_X1 U1061 ( .A(KEYINPUT15), .B(n1306), .Z(n1304) );
NOR2_X1 U1062 ( .A1(n1272), .A2(n1066), .ZN(n1306) );
INV_X1 U1063 ( .A(G134), .ZN(n1066) );
XNOR2_X1 U1064 ( .A(G128), .B(G143), .ZN(n1272) );
endmodule


