//Key = 1110110010011100101100010011000011100000100011101011010010100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336;

XOR2_X1 U735 ( .A(G107), .B(n1015), .Z(G9) );
NOR2_X1 U736 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U737 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
XOR2_X1 U738 ( .A(KEYINPUT27), .B(n1022), .Z(n1019) );
NOR3_X1 U739 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NOR3_X1 U740 ( .A1(n1026), .A2(KEYINPUT0), .A3(n1027), .ZN(n1025) );
AND4_X1 U741 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1027) );
NOR3_X1 U742 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1024) );
NOR2_X1 U743 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U744 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U745 ( .A1(n1039), .A2(n1026), .ZN(n1035) );
NOR2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
AND2_X1 U747 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
AND3_X1 U748 ( .A1(KEYINPUT0), .A2(n1028), .A3(n1030), .ZN(n1040) );
AND2_X1 U749 ( .A1(n1044), .A2(n1045), .ZN(n1023) );
NAND4_X1 U750 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1018) );
NAND3_X1 U751 ( .A1(n1029), .A2(n1050), .A3(n1031), .ZN(n1047) );
NAND3_X1 U752 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1050) );
NAND3_X1 U753 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NAND4_X1 U754 ( .A1(n1057), .A2(n1042), .A3(n1058), .A4(n1059), .ZN(n1052) );
XOR2_X1 U755 ( .A(KEYINPUT42), .B(n1060), .Z(n1058) );
NAND4_X1 U756 ( .A1(n1061), .A2(n1060), .A3(n1062), .A4(n1030), .ZN(n1051) );
NAND2_X1 U757 ( .A1(n1045), .A2(n1063), .ZN(n1046) );
NOR3_X1 U758 ( .A1(n1026), .A2(n1038), .A3(n1032), .ZN(n1045) );
INV_X1 U759 ( .A(n1031), .ZN(n1032) );
NOR2_X1 U760 ( .A1(KEYINPUT60), .A2(n1064), .ZN(n1031) );
INV_X1 U761 ( .A(n1060), .ZN(n1026) );
NOR3_X1 U762 ( .A1(n1065), .A2(G953), .A3(G952), .ZN(n1016) );
INV_X1 U763 ( .A(n1048), .ZN(n1065) );
NAND4_X1 U764 ( .A1(n1066), .A2(n1042), .A3(n1067), .A4(n1068), .ZN(n1048) );
NOR4_X1 U765 ( .A1(n1056), .A2(n1069), .A3(n1070), .A4(n1059), .ZN(n1068) );
NOR2_X1 U766 ( .A1(KEYINPUT63), .A2(n1071), .ZN(n1070) );
NOR2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1069) );
NOR2_X1 U768 ( .A1(KEYINPUT63), .A2(n1074), .ZN(n1072) );
NOR2_X1 U769 ( .A1(n1075), .A2(n1076), .ZN(n1067) );
XNOR2_X1 U770 ( .A(n1077), .B(n1078), .ZN(n1066) );
NAND2_X1 U771 ( .A1(KEYINPUT34), .A2(G472), .ZN(n1077) );
XOR2_X1 U772 ( .A(n1079), .B(n1080), .Z(G72) );
NOR2_X1 U773 ( .A1(n1081), .A2(n1049), .ZN(n1080) );
NOR2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XOR2_X1 U775 ( .A(KEYINPUT12), .B(G900), .Z(n1083) );
INV_X1 U776 ( .A(G227), .ZN(n1082) );
NAND2_X1 U777 ( .A1(n1084), .A2(n1085), .ZN(n1079) );
OR3_X1 U778 ( .A1(n1086), .A2(G953), .A3(n1087), .ZN(n1085) );
NAND3_X1 U779 ( .A1(n1088), .A2(n1089), .A3(n1087), .ZN(n1084) );
XNOR2_X1 U780 ( .A(n1090), .B(n1091), .ZN(n1087) );
XOR2_X1 U781 ( .A(G125), .B(n1092), .Z(n1091) );
NAND2_X1 U782 ( .A1(G953), .A2(n1093), .ZN(n1089) );
XOR2_X1 U783 ( .A(KEYINPUT52), .B(n1086), .Z(n1088) );
XOR2_X1 U784 ( .A(n1094), .B(n1095), .Z(G69) );
NOR2_X1 U785 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U786 ( .A1(KEYINPUT55), .A2(n1098), .ZN(n1097) );
INV_X1 U787 ( .A(n1099), .ZN(n1098) );
NOR2_X1 U788 ( .A1(KEYINPUT44), .A2(n1099), .ZN(n1096) );
XOR2_X1 U789 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR3_X1 U790 ( .A1(n1102), .A2(KEYINPUT17), .A3(G953), .ZN(n1101) );
NAND2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(n1100) );
NAND2_X1 U792 ( .A1(G953), .A2(n1105), .ZN(n1104) );
XOR2_X1 U793 ( .A(n1106), .B(n1107), .Z(n1103) );
XOR2_X1 U794 ( .A(G122), .B(n1108), .Z(n1107) );
NOR2_X1 U795 ( .A1(n1109), .A2(n1049), .ZN(n1094) );
NOR2_X1 U796 ( .A1(n1110), .A2(n1105), .ZN(n1109) );
NOR2_X1 U797 ( .A1(n1111), .A2(n1112), .ZN(G66) );
XOR2_X1 U798 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U799 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U800 ( .A1(n1111), .A2(n1117), .ZN(G63) );
XOR2_X1 U801 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR3_X1 U802 ( .A1(n1116), .A2(KEYINPUT54), .A3(n1120), .ZN(n1118) );
INV_X1 U803 ( .A(G478), .ZN(n1120) );
NOR2_X1 U804 ( .A1(n1111), .A2(n1121), .ZN(G60) );
XNOR2_X1 U805 ( .A(n1122), .B(n1123), .ZN(n1121) );
XOR2_X1 U806 ( .A(KEYINPUT7), .B(n1124), .Z(n1123) );
NOR2_X1 U807 ( .A1(n1125), .A2(n1116), .ZN(n1124) );
INV_X1 U808 ( .A(G475), .ZN(n1125) );
XOR2_X1 U809 ( .A(G104), .B(n1126), .Z(G6) );
NOR2_X1 U810 ( .A1(n1111), .A2(n1127), .ZN(G57) );
XOR2_X1 U811 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U813 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U814 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U815 ( .A(KEYINPUT56), .B(KEYINPUT53), .Z(n1135) );
NOR2_X1 U816 ( .A1(n1136), .A2(n1116), .ZN(n1130) );
XNOR2_X1 U817 ( .A(n1137), .B(n1138), .ZN(n1128) );
NOR2_X1 U818 ( .A1(n1111), .A2(n1139), .ZN(G54) );
XNOR2_X1 U819 ( .A(n1140), .B(n1141), .ZN(n1139) );
NOR2_X1 U820 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NOR2_X1 U821 ( .A1(KEYINPUT31), .A2(n1144), .ZN(n1143) );
AND2_X1 U822 ( .A1(KEYINPUT41), .A2(n1144), .ZN(n1142) );
NOR2_X1 U823 ( .A1(n1116), .A2(n1145), .ZN(n1144) );
NOR2_X1 U824 ( .A1(n1111), .A2(n1146), .ZN(G51) );
XOR2_X1 U825 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U826 ( .A(n1149), .B(n1150), .Z(n1147) );
NOR2_X1 U827 ( .A1(n1074), .A2(n1116), .ZN(n1150) );
NAND2_X1 U828 ( .A1(G902), .A2(n1151), .ZN(n1116) );
NAND2_X1 U829 ( .A1(n1102), .A2(n1086), .ZN(n1151) );
INV_X1 U830 ( .A(n1020), .ZN(n1086) );
NAND4_X1 U831 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1020) );
NOR4_X1 U832 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
NOR2_X1 U833 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR2_X1 U834 ( .A1(n1037), .A2(n1162), .ZN(n1158) );
NOR2_X1 U835 ( .A1(n1163), .A2(n1164), .ZN(n1154) );
INV_X1 U836 ( .A(n1021), .ZN(n1102) );
NAND4_X1 U837 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1021) );
NOR4_X1 U838 ( .A1(n1169), .A2(n1170), .A3(n1126), .A4(n1015), .ZN(n1168) );
AND3_X1 U839 ( .A1(n1030), .A2(n1063), .A3(n1171), .ZN(n1015) );
AND3_X1 U840 ( .A1(n1171), .A2(n1030), .A3(n1044), .ZN(n1126) );
NOR2_X1 U841 ( .A1(n1172), .A2(n1173), .ZN(n1167) );
NOR2_X1 U842 ( .A1(n1174), .A2(n1037), .ZN(n1173) );
XOR2_X1 U843 ( .A(n1175), .B(KEYINPUT22), .Z(n1174) );
INV_X1 U844 ( .A(n1176), .ZN(n1172) );
NAND2_X1 U845 ( .A1(n1177), .A2(n1178), .ZN(n1149) );
NAND2_X1 U846 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XOR2_X1 U847 ( .A(n1181), .B(KEYINPUT59), .Z(n1179) );
NOR2_X1 U848 ( .A1(n1049), .A2(G952), .ZN(n1111) );
XOR2_X1 U849 ( .A(n1153), .B(n1182), .Z(G48) );
XOR2_X1 U850 ( .A(KEYINPUT40), .B(G146), .Z(n1182) );
NAND4_X1 U851 ( .A1(n1028), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1153) );
AND2_X1 U852 ( .A1(n1044), .A2(n1186), .ZN(n1185) );
XOR2_X1 U853 ( .A(n1187), .B(G143), .Z(G45) );
NAND2_X1 U854 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
OR3_X1 U855 ( .A1(n1190), .A2(n1028), .A3(KEYINPUT5), .ZN(n1189) );
NAND2_X1 U856 ( .A1(n1157), .A2(KEYINPUT5), .ZN(n1188) );
NOR2_X1 U857 ( .A1(n1190), .A2(n1191), .ZN(n1157) );
INV_X1 U858 ( .A(n1028), .ZN(n1191) );
NAND3_X1 U859 ( .A1(n1192), .A2(n1043), .A3(n1193), .ZN(n1190) );
AND3_X1 U860 ( .A1(n1184), .A2(n1183), .A3(n1076), .ZN(n1193) );
XOR2_X1 U861 ( .A(G140), .B(n1194), .Z(G42) );
NOR3_X1 U862 ( .A1(n1161), .A2(KEYINPUT3), .A3(n1160), .ZN(n1194) );
XOR2_X1 U863 ( .A(G137), .B(n1156), .Z(G39) );
NOR3_X1 U864 ( .A1(n1195), .A2(n1034), .A3(n1161), .ZN(n1156) );
INV_X1 U865 ( .A(n1029), .ZN(n1034) );
XOR2_X1 U866 ( .A(G134), .B(n1164), .Z(G36) );
AND3_X1 U867 ( .A1(n1043), .A2(n1063), .A3(n1196), .ZN(n1164) );
XOR2_X1 U868 ( .A(n1197), .B(n1163), .Z(G33) );
AND3_X1 U869 ( .A1(n1044), .A2(n1043), .A3(n1196), .ZN(n1163) );
INV_X1 U870 ( .A(n1161), .ZN(n1196) );
NAND3_X1 U871 ( .A1(n1028), .A2(n1183), .A3(n1060), .ZN(n1161) );
NOR2_X1 U872 ( .A1(n1198), .A2(n1056), .ZN(n1060) );
NOR2_X1 U873 ( .A1(n1199), .A2(n1200), .ZN(n1197) );
XOR2_X1 U874 ( .A(KEYINPUT48), .B(KEYINPUT33), .Z(n1200) );
INV_X1 U875 ( .A(G131), .ZN(n1199) );
XNOR2_X1 U876 ( .A(G128), .B(n1201), .ZN(G30) );
NAND2_X1 U877 ( .A1(n1202), .A2(n1184), .ZN(n1201) );
XOR2_X1 U878 ( .A(n1162), .B(KEYINPUT11), .Z(n1202) );
NAND4_X1 U879 ( .A1(n1203), .A2(n1186), .A3(n1063), .A4(n1183), .ZN(n1162) );
XOR2_X1 U880 ( .A(n1170), .B(n1204), .Z(G3) );
XOR2_X1 U881 ( .A(KEYINPUT49), .B(G101), .Z(n1204) );
AND3_X1 U882 ( .A1(n1171), .A2(n1029), .A3(n1043), .ZN(n1170) );
NAND2_X1 U883 ( .A1(n1205), .A2(n1206), .ZN(G27) );
NAND2_X1 U884 ( .A1(G125), .A2(n1152), .ZN(n1206) );
XOR2_X1 U885 ( .A(KEYINPUT4), .B(n1207), .Z(n1205) );
NOR2_X1 U886 ( .A1(G125), .A2(n1152), .ZN(n1207) );
NAND4_X1 U887 ( .A1(n1208), .A2(n1042), .A3(n1184), .A4(n1183), .ZN(n1152) );
NAND2_X1 U888 ( .A1(n1209), .A2(n1210), .ZN(n1183) );
NAND4_X1 U889 ( .A1(G953), .A2(G902), .A3(n1211), .A4(n1093), .ZN(n1210) );
INV_X1 U890 ( .A(G900), .ZN(n1093) );
INV_X1 U891 ( .A(n1160), .ZN(n1208) );
NAND3_X1 U892 ( .A1(n1057), .A2(n1059), .A3(n1044), .ZN(n1160) );
XOR2_X1 U893 ( .A(G122), .B(n1212), .Z(G24) );
NOR2_X1 U894 ( .A1(n1037), .A2(n1175), .ZN(n1212) );
NAND4_X1 U895 ( .A1(n1192), .A2(n1055), .A3(n1076), .A4(n1213), .ZN(n1175) );
INV_X1 U896 ( .A(n1038), .ZN(n1055) );
NAND2_X1 U897 ( .A1(n1042), .A2(n1030), .ZN(n1038) );
NOR2_X1 U898 ( .A1(n1059), .A2(n1214), .ZN(n1030) );
INV_X1 U899 ( .A(n1184), .ZN(n1037) );
XOR2_X1 U900 ( .A(n1215), .B(n1176), .Z(G21) );
NAND3_X1 U901 ( .A1(n1216), .A2(n1029), .A3(n1186), .ZN(n1176) );
INV_X1 U902 ( .A(n1195), .ZN(n1186) );
NAND2_X1 U903 ( .A1(n1214), .A2(n1059), .ZN(n1195) );
INV_X1 U904 ( .A(n1057), .ZN(n1214) );
XOR2_X1 U905 ( .A(n1217), .B(n1165), .Z(G18) );
NAND3_X1 U906 ( .A1(n1043), .A2(n1063), .A3(n1216), .ZN(n1165) );
NAND2_X1 U907 ( .A1(n1218), .A2(n1219), .ZN(n1063) );
NAND3_X1 U908 ( .A1(n1220), .A2(n1076), .A3(n1221), .ZN(n1219) );
INV_X1 U909 ( .A(KEYINPUT21), .ZN(n1221) );
NAND2_X1 U910 ( .A1(KEYINPUT21), .A2(n1029), .ZN(n1218) );
XNOR2_X1 U911 ( .A(G113), .B(n1166), .ZN(G15) );
NAND3_X1 U912 ( .A1(n1044), .A2(n1043), .A3(n1216), .ZN(n1166) );
AND3_X1 U913 ( .A1(n1184), .A2(n1213), .A3(n1042), .ZN(n1216) );
NOR2_X1 U914 ( .A1(n1222), .A2(n1061), .ZN(n1042) );
NOR2_X1 U915 ( .A1(n1059), .A2(n1057), .ZN(n1043) );
NOR2_X1 U916 ( .A1(n1220), .A2(n1076), .ZN(n1044) );
INV_X1 U917 ( .A(n1192), .ZN(n1220) );
XNOR2_X1 U918 ( .A(n1169), .B(n1223), .ZN(G12) );
NAND2_X1 U919 ( .A1(KEYINPUT45), .A2(G110), .ZN(n1223) );
AND4_X1 U920 ( .A1(n1171), .A2(n1029), .A3(n1057), .A4(n1059), .ZN(n1169) );
NAND3_X1 U921 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1059) );
NAND2_X1 U922 ( .A1(G217), .A2(G902), .ZN(n1226) );
OR3_X1 U923 ( .A1(n1113), .A2(G902), .A3(n1227), .ZN(n1225) );
NAND2_X1 U924 ( .A1(n1113), .A2(n1227), .ZN(n1224) );
NOR2_X1 U925 ( .A1(n1115), .A2(G234), .ZN(n1227) );
XOR2_X1 U926 ( .A(n1228), .B(n1229), .Z(n1113) );
XOR2_X1 U927 ( .A(G110), .B(n1230), .Z(n1229) );
XOR2_X1 U928 ( .A(G146), .B(G137), .Z(n1230) );
XOR2_X1 U929 ( .A(n1231), .B(n1232), .Z(n1228) );
XOR2_X1 U930 ( .A(n1233), .B(n1234), .Z(n1232) );
NAND3_X1 U931 ( .A1(G234), .A2(n1049), .A3(G221), .ZN(n1234) );
NAND3_X1 U932 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1233) );
NAND2_X1 U933 ( .A1(KEYINPUT14), .A2(n1215), .ZN(n1237) );
NAND3_X1 U934 ( .A1(n1238), .A2(n1239), .A3(G128), .ZN(n1236) );
INV_X1 U935 ( .A(KEYINPUT14), .ZN(n1239) );
OR2_X1 U936 ( .A1(n1238), .A2(G128), .ZN(n1235) );
NOR2_X1 U937 ( .A1(KEYINPUT28), .A2(n1215), .ZN(n1238) );
NAND2_X1 U938 ( .A1(n1240), .A2(n1241), .ZN(n1231) );
NAND2_X1 U939 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XNOR2_X1 U940 ( .A(n1244), .B(KEYINPUT13), .ZN(n1242) );
NAND2_X1 U941 ( .A1(n1245), .A2(G125), .ZN(n1240) );
XNOR2_X1 U942 ( .A(n1244), .B(KEYINPUT35), .ZN(n1245) );
XOR2_X1 U943 ( .A(n1078), .B(n1246), .Z(n1057) );
NOR2_X1 U944 ( .A1(KEYINPUT20), .A2(n1136), .ZN(n1246) );
INV_X1 U945 ( .A(G472), .ZN(n1136) );
NAND2_X1 U946 ( .A1(n1247), .A2(n1248), .ZN(n1078) );
XOR2_X1 U947 ( .A(n1249), .B(n1250), .Z(n1247) );
XOR2_X1 U948 ( .A(n1138), .B(n1134), .Z(n1250) );
XNOR2_X1 U949 ( .A(n1251), .B(n1252), .ZN(n1134) );
XNOR2_X1 U950 ( .A(n1253), .B(G101), .ZN(n1138) );
NAND2_X1 U951 ( .A1(n1254), .A2(G210), .ZN(n1253) );
XNOR2_X1 U952 ( .A(n1255), .B(n1256), .ZN(n1249) );
NAND2_X1 U953 ( .A1(KEYINPUT8), .A2(n1137), .ZN(n1256) );
NAND2_X1 U954 ( .A1(KEYINPUT19), .A2(n1132), .ZN(n1255) );
AND3_X1 U955 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1132) );
NAND2_X1 U956 ( .A1(n1260), .A2(n1215), .ZN(n1259) );
XOR2_X1 U957 ( .A(n1217), .B(n1261), .Z(n1260) );
INV_X1 U958 ( .A(n1262), .ZN(n1257) );
NOR2_X1 U959 ( .A1(n1076), .A2(n1192), .ZN(n1029) );
XNOR2_X1 U960 ( .A(n1075), .B(KEYINPUT51), .ZN(n1192) );
XNOR2_X1 U961 ( .A(n1263), .B(G475), .ZN(n1075) );
NAND2_X1 U962 ( .A1(n1122), .A2(n1248), .ZN(n1263) );
XNOR2_X1 U963 ( .A(n1264), .B(n1265), .ZN(n1122) );
XOR2_X1 U964 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U965 ( .A(n1243), .B(n1268), .Z(n1267) );
NOR2_X1 U966 ( .A1(KEYINPUT36), .A2(n1269), .ZN(n1268) );
XOR2_X1 U967 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U968 ( .A(G104), .B(n1261), .Z(n1271) );
XOR2_X1 U969 ( .A(KEYINPUT47), .B(G122), .Z(n1270) );
NAND2_X1 U970 ( .A1(KEYINPUT61), .A2(n1272), .ZN(n1266) );
XOR2_X1 U971 ( .A(n1273), .B(n1274), .Z(n1264) );
AND2_X1 U972 ( .A1(G214), .A2(n1254), .ZN(n1274) );
NOR2_X1 U973 ( .A1(G953), .A2(G237), .ZN(n1254) );
XNOR2_X1 U974 ( .A(n1275), .B(G478), .ZN(n1076) );
OR2_X1 U975 ( .A1(n1119), .A2(G902), .ZN(n1275) );
XNOR2_X1 U976 ( .A(n1276), .B(n1277), .ZN(n1119) );
XOR2_X1 U977 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U978 ( .A(n1280), .B(n1281), .Z(n1279) );
NOR3_X1 U979 ( .A1(n1282), .A2(n1283), .A3(n1115), .ZN(n1281) );
INV_X1 U980 ( .A(G217), .ZN(n1115) );
INV_X1 U981 ( .A(G234), .ZN(n1283) );
XOR2_X1 U982 ( .A(KEYINPUT43), .B(G953), .Z(n1282) );
NAND2_X1 U983 ( .A1(n1284), .A2(n1285), .ZN(n1280) );
NAND2_X1 U984 ( .A1(G116), .A2(n1286), .ZN(n1285) );
INV_X1 U985 ( .A(G122), .ZN(n1286) );
XOR2_X1 U986 ( .A(n1287), .B(KEYINPUT57), .Z(n1284) );
NAND2_X1 U987 ( .A1(n1288), .A2(n1217), .ZN(n1287) );
XOR2_X1 U988 ( .A(KEYINPUT25), .B(G122), .Z(n1288) );
NAND2_X1 U989 ( .A1(KEYINPUT50), .A2(G128), .ZN(n1278) );
XOR2_X1 U990 ( .A(n1289), .B(n1290), .Z(n1276) );
XOR2_X1 U991 ( .A(KEYINPUT39), .B(G143), .Z(n1290) );
XOR2_X1 U992 ( .A(G134), .B(n1291), .Z(n1289) );
AND3_X1 U993 ( .A1(n1203), .A2(n1213), .A3(n1184), .ZN(n1171) );
NOR2_X1 U994 ( .A1(n1056), .A2(n1054), .ZN(n1184) );
INV_X1 U995 ( .A(n1198), .ZN(n1054) );
NAND2_X1 U996 ( .A1(n1292), .A2(n1071), .ZN(n1198) );
NAND2_X1 U997 ( .A1(n1293), .A2(n1073), .ZN(n1071) );
OR2_X1 U998 ( .A1(n1073), .A2(n1293), .ZN(n1292) );
INV_X1 U999 ( .A(n1074), .ZN(n1293) );
NAND2_X1 U1000 ( .A1(G210), .A2(n1294), .ZN(n1074) );
NAND2_X1 U1001 ( .A1(n1295), .A2(n1248), .ZN(n1073) );
XOR2_X1 U1002 ( .A(n1296), .B(n1297), .Z(n1295) );
NOR2_X1 U1003 ( .A1(KEYINPUT24), .A2(n1148), .ZN(n1297) );
XNOR2_X1 U1004 ( .A(n1106), .B(n1298), .ZN(n1148) );
XOR2_X1 U1005 ( .A(G101), .B(n1299), .Z(n1298) );
NOR2_X1 U1006 ( .A1(KEYINPUT30), .A2(n1300), .ZN(n1299) );
XOR2_X1 U1007 ( .A(G122), .B(G110), .Z(n1300) );
XOR2_X1 U1008 ( .A(n1301), .B(n1302), .Z(n1106) );
NOR2_X1 U1009 ( .A1(KEYINPUT9), .A2(n1303), .ZN(n1302) );
NOR2_X1 U1010 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NOR2_X1 U1011 ( .A1(G104), .A2(n1291), .ZN(n1304) );
INV_X1 U1012 ( .A(G107), .ZN(n1291) );
NAND4_X1 U1013 ( .A1(n1306), .A2(n1258), .A3(n1307), .A4(n1308), .ZN(n1301) );
NAND3_X1 U1014 ( .A1(KEYINPUT15), .A2(n1261), .A3(G119), .ZN(n1308) );
NAND2_X1 U1015 ( .A1(n1309), .A2(n1215), .ZN(n1307) );
XOR2_X1 U1016 ( .A(n1310), .B(n1261), .Z(n1309) );
NAND2_X1 U1017 ( .A1(G116), .A2(n1311), .ZN(n1310) );
NAND3_X1 U1018 ( .A1(n1261), .A2(n1217), .A3(G119), .ZN(n1258) );
NAND2_X1 U1019 ( .A1(n1262), .A2(n1311), .ZN(n1306) );
INV_X1 U1020 ( .A(KEYINPUT15), .ZN(n1311) );
NOR3_X1 U1021 ( .A1(n1217), .A2(n1215), .A3(n1261), .ZN(n1262) );
XOR2_X1 U1022 ( .A(G113), .B(KEYINPUT6), .Z(n1261) );
INV_X1 U1023 ( .A(G119), .ZN(n1215) );
INV_X1 U1024 ( .A(G116), .ZN(n1217) );
NAND2_X1 U1025 ( .A1(n1312), .A2(n1313), .ZN(n1296) );
NAND2_X1 U1026 ( .A1(n1180), .A2(n1181), .ZN(n1313) );
XNOR2_X1 U1027 ( .A(KEYINPUT1), .B(n1177), .ZN(n1312) );
OR2_X1 U1028 ( .A1(n1181), .A2(n1180), .ZN(n1177) );
NOR2_X1 U1029 ( .A1(n1110), .A2(G953), .ZN(n1180) );
INV_X1 U1030 ( .A(G224), .ZN(n1110) );
XOR2_X1 U1031 ( .A(n1137), .B(n1243), .Z(n1181) );
INV_X1 U1032 ( .A(G125), .ZN(n1243) );
XNOR2_X1 U1033 ( .A(n1314), .B(n1315), .ZN(n1137) );
XOR2_X1 U1034 ( .A(G146), .B(G143), .Z(n1315) );
NAND2_X1 U1035 ( .A1(KEYINPUT2), .A2(G128), .ZN(n1314) );
AND2_X1 U1036 ( .A1(G214), .A2(n1294), .ZN(n1056) );
NAND2_X1 U1037 ( .A1(n1316), .A2(n1248), .ZN(n1294) );
XOR2_X1 U1038 ( .A(KEYINPUT26), .B(G237), .Z(n1316) );
NAND2_X1 U1039 ( .A1(n1317), .A2(n1209), .ZN(n1213) );
OR2_X1 U1040 ( .A1(n1064), .A2(G953), .ZN(n1209) );
NAND2_X1 U1041 ( .A1(n1318), .A2(n1211), .ZN(n1064) );
XNOR2_X1 U1042 ( .A(G952), .B(KEYINPUT62), .ZN(n1318) );
NAND4_X1 U1043 ( .A1(n1319), .A2(G953), .A3(G902), .A4(n1105), .ZN(n1317) );
INV_X1 U1044 ( .A(G898), .ZN(n1105) );
XOR2_X1 U1045 ( .A(n1211), .B(KEYINPUT37), .Z(n1319) );
NAND2_X1 U1046 ( .A1(G237), .A2(G234), .ZN(n1211) );
XNOR2_X1 U1047 ( .A(n1028), .B(KEYINPUT18), .ZN(n1203) );
NOR2_X1 U1048 ( .A1(n1062), .A2(n1061), .ZN(n1028) );
AND2_X1 U1049 ( .A1(G221), .A2(n1320), .ZN(n1061) );
NAND2_X1 U1050 ( .A1(G234), .A2(n1248), .ZN(n1320) );
INV_X1 U1051 ( .A(n1222), .ZN(n1062) );
XOR2_X1 U1052 ( .A(n1321), .B(n1145), .Z(n1222) );
INV_X1 U1053 ( .A(G469), .ZN(n1145) );
NAND2_X1 U1054 ( .A1(n1140), .A2(n1248), .ZN(n1321) );
INV_X1 U1055 ( .A(G902), .ZN(n1248) );
XNOR2_X1 U1056 ( .A(n1322), .B(n1323), .ZN(n1140) );
XOR2_X1 U1057 ( .A(n1324), .B(n1325), .Z(n1323) );
XOR2_X1 U1058 ( .A(n1251), .B(n1326), .Z(n1325) );
NOR2_X1 U1059 ( .A1(n1305), .A2(n1327), .ZN(n1326) );
XOR2_X1 U1060 ( .A(n1328), .B(KEYINPUT23), .Z(n1327) );
NAND2_X1 U1061 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XOR2_X1 U1062 ( .A(KEYINPUT10), .B(G107), .Z(n1329) );
NOR2_X1 U1063 ( .A1(n1330), .A2(G107), .ZN(n1305) );
INV_X1 U1064 ( .A(G104), .ZN(n1330) );
NAND2_X1 U1065 ( .A1(KEYINPUT58), .A2(n1092), .ZN(n1251) );
XOR2_X1 U1066 ( .A(G134), .B(n1331), .Z(n1092) );
XOR2_X1 U1067 ( .A(KEYINPUT29), .B(G137), .Z(n1331) );
NAND2_X1 U1068 ( .A1(G227), .A2(n1049), .ZN(n1324) );
INV_X1 U1069 ( .A(G953), .ZN(n1049) );
XOR2_X1 U1070 ( .A(n1090), .B(n1108), .Z(n1322) );
XOR2_X1 U1071 ( .A(G101), .B(G110), .Z(n1108) );
XOR2_X1 U1072 ( .A(n1332), .B(n1333), .Z(n1090) );
XOR2_X1 U1073 ( .A(n1334), .B(n1273), .Z(n1333) );
XOR2_X1 U1074 ( .A(n1335), .B(n1252), .Z(n1273) );
XOR2_X1 U1075 ( .A(G131), .B(KEYINPUT16), .Z(n1252) );
XOR2_X1 U1076 ( .A(n1336), .B(n1244), .Z(n1335) );
XOR2_X1 U1077 ( .A(G140), .B(KEYINPUT46), .Z(n1244) );
INV_X1 U1078 ( .A(G146), .ZN(n1336) );
NAND2_X1 U1079 ( .A1(KEYINPUT32), .A2(n1272), .ZN(n1334) );
INV_X1 U1080 ( .A(G143), .ZN(n1272) );
XNOR2_X1 U1081 ( .A(G128), .B(KEYINPUT38), .ZN(n1332) );
endmodule


