//Key = 0011000011100100100011111101010111101100000000010111001110100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363;

XNOR2_X1 U752 ( .A(n1033), .B(n1034), .ZN(G9) );
NOR2_X1 U753 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND4_X1 U754 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(G75) );
NAND3_X1 U755 ( .A1(KEYINPUT41), .A2(n1041), .A3(n1042), .ZN(n1040) );
NAND2_X1 U756 ( .A1(G952), .A2(n1043), .ZN(n1039) );
NAND3_X1 U757 ( .A1(n1044), .A2(n1041), .A3(n1045), .ZN(n1043) );
NAND2_X1 U758 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NAND2_X1 U759 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND3_X1 U760 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
NAND2_X1 U761 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NAND2_X1 U762 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U763 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U764 ( .A1(n1059), .A2(n1060), .ZN(n1053) );
NAND2_X1 U765 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U766 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
INV_X1 U767 ( .A(n1065), .ZN(n1061) );
NAND3_X1 U768 ( .A1(n1055), .A2(n1066), .A3(n1059), .ZN(n1048) );
NAND2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U770 ( .A1(n1052), .A2(n1069), .ZN(n1068) );
NAND2_X1 U771 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U772 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
INV_X1 U773 ( .A(n1074), .ZN(n1070) );
NAND2_X1 U774 ( .A1(n1050), .A2(n1075), .ZN(n1067) );
NAND2_X1 U775 ( .A1(n1036), .A2(n1076), .ZN(n1075) );
NAND2_X1 U776 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
INV_X1 U777 ( .A(n1079), .ZN(n1046) );
OR2_X1 U778 ( .A1(n1041), .A2(KEYINPUT41), .ZN(n1038) );
NAND4_X1 U779 ( .A1(n1055), .A2(n1052), .A3(n1080), .A4(n1081), .ZN(n1041) );
NOR4_X1 U780 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1081) );
XOR2_X1 U781 ( .A(n1086), .B(n1087), .Z(n1083) );
NAND2_X1 U782 ( .A1(KEYINPUT55), .A2(n1088), .ZN(n1086) );
AND2_X1 U783 ( .A1(n1089), .A2(n1090), .ZN(n1082) );
NOR2_X1 U784 ( .A1(n1091), .A2(n1092), .ZN(n1080) );
NOR2_X1 U785 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
INV_X1 U786 ( .A(KEYINPUT10), .ZN(n1094) );
NOR2_X1 U787 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NOR3_X1 U788 ( .A1(n1089), .A2(KEYINPUT11), .A3(n1090), .ZN(n1096) );
AND2_X1 U789 ( .A1(n1089), .A2(KEYINPUT11), .ZN(n1095) );
INV_X1 U790 ( .A(G478), .ZN(n1089) );
NOR2_X1 U791 ( .A1(KEYINPUT10), .A2(n1097), .ZN(n1091) );
NOR2_X1 U792 ( .A1(n1090), .A2(n1098), .ZN(n1097) );
XNOR2_X1 U793 ( .A(KEYINPUT11), .B(G478), .ZN(n1098) );
XOR2_X1 U794 ( .A(n1099), .B(n1100), .Z(G72) );
XOR2_X1 U795 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U796 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
AND2_X1 U797 ( .A1(G227), .A2(G900), .ZN(n1103) );
NAND2_X1 U798 ( .A1(n1105), .A2(n1106), .ZN(n1101) );
NAND2_X1 U799 ( .A1(G953), .A2(n1107), .ZN(n1106) );
XOR2_X1 U800 ( .A(n1108), .B(n1109), .Z(n1105) );
XNOR2_X1 U801 ( .A(n1110), .B(n1111), .ZN(n1109) );
XNOR2_X1 U802 ( .A(n1112), .B(n1113), .ZN(n1108) );
NAND2_X1 U803 ( .A1(n1104), .A2(n1114), .ZN(n1099) );
NAND2_X1 U804 ( .A1(n1115), .A2(n1116), .ZN(G69) );
NAND2_X1 U805 ( .A1(n1117), .A2(n1104), .ZN(n1116) );
XNOR2_X1 U806 ( .A(n1118), .B(n1119), .ZN(n1117) );
NAND2_X1 U807 ( .A1(n1120), .A2(G953), .ZN(n1115) );
NAND2_X1 U808 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U809 ( .A1(n1119), .A2(n1123), .ZN(n1122) );
INV_X1 U810 ( .A(G224), .ZN(n1123) );
NAND2_X1 U811 ( .A1(G224), .A2(n1124), .ZN(n1121) );
NAND2_X1 U812 ( .A1(G898), .A2(n1119), .ZN(n1124) );
NAND2_X1 U813 ( .A1(n1125), .A2(n1126), .ZN(n1119) );
NAND2_X1 U814 ( .A1(G953), .A2(n1127), .ZN(n1126) );
XNOR2_X1 U815 ( .A(n1128), .B(n1129), .ZN(n1125) );
NOR2_X1 U816 ( .A1(n1130), .A2(n1131), .ZN(G66) );
XOR2_X1 U817 ( .A(n1132), .B(KEYINPUT20), .Z(n1131) );
NAND2_X1 U818 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U819 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U820 ( .A(KEYINPUT56), .B(n1137), .Z(n1133) );
NOR2_X1 U821 ( .A1(n1135), .A2(n1136), .ZN(n1137) );
NAND3_X1 U822 ( .A1(G217), .A2(n1138), .A3(n1139), .ZN(n1136) );
NOR2_X1 U823 ( .A1(n1130), .A2(n1140), .ZN(G63) );
XOR2_X1 U824 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U825 ( .A(n1143), .B(KEYINPUT33), .Z(n1142) );
NAND2_X1 U826 ( .A1(n1139), .A2(G478), .ZN(n1143) );
NOR2_X1 U827 ( .A1(n1130), .A2(n1144), .ZN(G60) );
XOR2_X1 U828 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND2_X1 U829 ( .A1(n1139), .A2(G475), .ZN(n1145) );
XNOR2_X1 U830 ( .A(G104), .B(n1147), .ZN(G6) );
NOR2_X1 U831 ( .A1(n1130), .A2(n1148), .ZN(G57) );
XOR2_X1 U832 ( .A(n1149), .B(n1150), .Z(n1148) );
XNOR2_X1 U833 ( .A(G101), .B(n1151), .ZN(n1150) );
NAND2_X1 U834 ( .A1(KEYINPUT8), .A2(n1152), .ZN(n1151) );
NAND2_X1 U835 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND2_X1 U836 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XNOR2_X1 U837 ( .A(n1157), .B(n1158), .ZN(n1156) );
XOR2_X1 U838 ( .A(n1159), .B(KEYINPUT50), .Z(n1155) );
NAND2_X1 U839 ( .A1(n1160), .A2(n1159), .ZN(n1153) );
NAND2_X1 U840 ( .A1(n1139), .A2(G472), .ZN(n1159) );
XOR2_X1 U841 ( .A(n1158), .B(n1157), .Z(n1160) );
NOR2_X1 U842 ( .A1(KEYINPUT30), .A2(n1161), .ZN(n1157) );
NAND2_X1 U843 ( .A1(n1162), .A2(n1163), .ZN(n1158) );
NAND2_X1 U844 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XOR2_X1 U845 ( .A(n1166), .B(KEYINPUT18), .Z(n1162) );
NAND2_X1 U846 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NOR2_X1 U847 ( .A1(KEYINPUT60), .A2(n1169), .ZN(n1149) );
NOR2_X1 U848 ( .A1(n1130), .A2(n1170), .ZN(G54) );
XOR2_X1 U849 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U850 ( .A(n1173), .B(n1174), .Z(n1172) );
XNOR2_X1 U851 ( .A(n1175), .B(n1176), .ZN(n1174) );
NAND2_X1 U852 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
NAND2_X1 U853 ( .A1(KEYINPUT27), .A2(n1179), .ZN(n1178) );
OR3_X1 U854 ( .A1(n1180), .A2(G110), .A3(KEYINPUT27), .ZN(n1177) );
XOR2_X1 U855 ( .A(n1181), .B(n1182), .Z(n1173) );
NOR2_X1 U856 ( .A1(KEYINPUT45), .A2(n1183), .ZN(n1182) );
NAND2_X1 U857 ( .A1(n1139), .A2(G469), .ZN(n1181) );
XOR2_X1 U858 ( .A(n1184), .B(n1185), .Z(n1171) );
XNOR2_X1 U859 ( .A(n1164), .B(n1186), .ZN(n1185) );
XOR2_X1 U860 ( .A(KEYINPUT49), .B(KEYINPUT44), .Z(n1184) );
NOR2_X1 U861 ( .A1(n1187), .A2(G952), .ZN(n1130) );
NOR2_X1 U862 ( .A1(n1188), .A2(n1189), .ZN(G51) );
NOR2_X1 U863 ( .A1(n1187), .A2(n1190), .ZN(n1189) );
XNOR2_X1 U864 ( .A(KEYINPUT59), .B(n1042), .ZN(n1190) );
INV_X1 U865 ( .A(G952), .ZN(n1042) );
XOR2_X1 U866 ( .A(n1104), .B(KEYINPUT7), .Z(n1187) );
NOR2_X1 U867 ( .A1(n1191), .A2(n1192), .ZN(n1188) );
XOR2_X1 U868 ( .A(n1193), .B(KEYINPUT24), .Z(n1192) );
NAND2_X1 U869 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
XNOR2_X1 U870 ( .A(n1196), .B(n1197), .ZN(n1195) );
NOR2_X1 U871 ( .A1(KEYINPUT6), .A2(n1198), .ZN(n1196) );
NOR3_X1 U872 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1191) );
NOR2_X1 U873 ( .A1(n1198), .A2(n1202), .ZN(n1201) );
XNOR2_X1 U874 ( .A(KEYINPUT6), .B(n1197), .ZN(n1202) );
NOR2_X1 U875 ( .A1(n1203), .A2(n1197), .ZN(n1200) );
XOR2_X1 U876 ( .A(n1204), .B(n1205), .Z(n1197) );
XNOR2_X1 U877 ( .A(n1194), .B(KEYINPUT47), .ZN(n1199) );
AND2_X1 U878 ( .A1(n1139), .A2(n1206), .ZN(n1194) );
NOR2_X1 U879 ( .A1(n1207), .A2(n1045), .ZN(n1139) );
NOR2_X1 U880 ( .A1(n1114), .A2(n1118), .ZN(n1045) );
NAND4_X1 U881 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1118) );
AND4_X1 U882 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1211) );
NOR2_X1 U883 ( .A1(n1216), .A2(n1217), .ZN(n1210) );
NOR2_X1 U884 ( .A1(n1218), .A2(n1036), .ZN(n1217) );
INV_X1 U885 ( .A(n1219), .ZN(n1036) );
XOR2_X1 U886 ( .A(n1035), .B(KEYINPUT5), .Z(n1218) );
NAND4_X1 U887 ( .A1(n1065), .A2(n1220), .A3(n1050), .A4(n1221), .ZN(n1035) );
INV_X1 U888 ( .A(n1147), .ZN(n1216) );
NAND3_X1 U889 ( .A1(n1222), .A2(n1050), .A3(n1223), .ZN(n1147) );
NAND4_X1 U890 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1114) );
NOR4_X1 U891 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1227) );
AND2_X1 U892 ( .A1(n1232), .A2(n1233), .ZN(n1226) );
XNOR2_X1 U893 ( .A(G146), .B(n1224), .ZN(G48) );
NAND3_X1 U894 ( .A1(n1222), .A2(n1219), .A3(n1234), .ZN(n1224) );
XNOR2_X1 U895 ( .A(G143), .B(n1225), .ZN(G45) );
NAND4_X1 U896 ( .A1(n1235), .A2(n1219), .A3(n1236), .A4(n1085), .ZN(n1225) );
XNOR2_X1 U897 ( .A(n1180), .B(n1231), .ZN(G42) );
AND3_X1 U898 ( .A1(n1052), .A2(n1065), .A3(n1237), .ZN(n1231) );
INV_X1 U899 ( .A(G140), .ZN(n1180) );
XOR2_X1 U900 ( .A(G137), .B(n1230), .Z(G39) );
AND3_X1 U901 ( .A1(n1234), .A2(n1052), .A3(n1059), .ZN(n1230) );
XNOR2_X1 U902 ( .A(G134), .B(n1233), .ZN(G36) );
NAND3_X1 U903 ( .A1(n1052), .A2(n1220), .A3(n1235), .ZN(n1233) );
XNOR2_X1 U904 ( .A(G131), .B(n1232), .ZN(G33) );
NAND3_X1 U905 ( .A1(n1222), .A2(n1052), .A3(n1235), .ZN(n1232) );
AND3_X1 U906 ( .A1(n1074), .A2(n1238), .A3(n1065), .ZN(n1235) );
NOR2_X1 U907 ( .A1(n1239), .A2(n1077), .ZN(n1052) );
XOR2_X1 U908 ( .A(G128), .B(n1229), .Z(G30) );
AND3_X1 U909 ( .A1(n1219), .A2(n1220), .A3(n1234), .ZN(n1229) );
AND4_X1 U910 ( .A1(n1065), .A2(n1073), .A3(n1084), .A4(n1238), .ZN(n1234) );
XNOR2_X1 U911 ( .A(G101), .B(n1208), .ZN(G3) );
NAND3_X1 U912 ( .A1(n1059), .A2(n1074), .A3(n1223), .ZN(n1208) );
XOR2_X1 U913 ( .A(n1240), .B(n1228), .Z(G27) );
AND3_X1 U914 ( .A1(n1055), .A2(n1219), .A3(n1237), .ZN(n1228) );
AND4_X1 U915 ( .A1(n1072), .A2(n1222), .A3(n1073), .A4(n1238), .ZN(n1237) );
NAND2_X1 U916 ( .A1(n1079), .A2(n1241), .ZN(n1238) );
NAND4_X1 U917 ( .A1(G953), .A2(G902), .A3(n1242), .A4(n1107), .ZN(n1241) );
INV_X1 U918 ( .A(G900), .ZN(n1107) );
XNOR2_X1 U919 ( .A(G125), .B(KEYINPUT31), .ZN(n1240) );
XNOR2_X1 U920 ( .A(G122), .B(n1209), .ZN(G24) );
NAND4_X1 U921 ( .A1(n1236), .A2(n1243), .A3(n1050), .A4(n1085), .ZN(n1209) );
NAND2_X1 U922 ( .A1(n1244), .A2(n1245), .ZN(n1050) );
OR3_X1 U923 ( .A1(n1073), .A2(n1084), .A3(KEYINPUT26), .ZN(n1245) );
NAND2_X1 U924 ( .A1(KEYINPUT26), .A2(n1074), .ZN(n1244) );
XNOR2_X1 U925 ( .A(G119), .B(n1215), .ZN(G21) );
NAND4_X1 U926 ( .A1(n1243), .A2(n1059), .A3(n1073), .A4(n1084), .ZN(n1215) );
XNOR2_X1 U927 ( .A(G116), .B(n1214), .ZN(G18) );
NAND3_X1 U928 ( .A1(n1220), .A2(n1074), .A3(n1243), .ZN(n1214) );
INV_X1 U929 ( .A(n1058), .ZN(n1220) );
NAND2_X1 U930 ( .A1(n1236), .A2(n1246), .ZN(n1058) );
XOR2_X1 U931 ( .A(KEYINPUT37), .B(n1085), .Z(n1246) );
XNOR2_X1 U932 ( .A(G113), .B(n1213), .ZN(G15) );
NAND3_X1 U933 ( .A1(n1222), .A2(n1074), .A3(n1243), .ZN(n1213) );
AND3_X1 U934 ( .A1(n1219), .A2(n1221), .A3(n1055), .ZN(n1243) );
NOR2_X1 U935 ( .A1(n1247), .A2(n1063), .ZN(n1055) );
NOR2_X1 U936 ( .A1(n1073), .A2(n1072), .ZN(n1074) );
INV_X1 U937 ( .A(n1057), .ZN(n1222) );
NAND2_X1 U938 ( .A1(n1248), .A2(n1085), .ZN(n1057) );
XNOR2_X1 U939 ( .A(KEYINPUT17), .B(n1236), .ZN(n1248) );
XOR2_X1 U940 ( .A(n1212), .B(n1249), .Z(G12) );
XOR2_X1 U941 ( .A(KEYINPUT23), .B(G110), .Z(n1249) );
NAND4_X1 U942 ( .A1(n1223), .A2(n1059), .A3(n1072), .A4(n1073), .ZN(n1212) );
XNOR2_X1 U943 ( .A(n1088), .B(n1087), .ZN(n1073) );
AND2_X1 U944 ( .A1(G217), .A2(n1250), .ZN(n1087) );
XNOR2_X1 U945 ( .A(KEYINPUT34), .B(n1138), .ZN(n1250) );
NAND2_X1 U946 ( .A1(n1251), .A2(n1135), .ZN(n1088) );
XNOR2_X1 U947 ( .A(n1252), .B(n1253), .ZN(n1135) );
NOR2_X1 U948 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
XOR2_X1 U949 ( .A(KEYINPUT35), .B(n1256), .Z(n1255) );
NOR2_X1 U950 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NOR2_X1 U951 ( .A1(n1259), .A2(n1260), .ZN(n1254) );
XOR2_X1 U952 ( .A(n1257), .B(KEYINPUT22), .Z(n1260) );
XNOR2_X1 U953 ( .A(G146), .B(n1261), .ZN(n1257) );
NOR2_X1 U954 ( .A1(KEYINPUT19), .A2(n1112), .ZN(n1261) );
INV_X1 U955 ( .A(n1258), .ZN(n1259) );
XOR2_X1 U956 ( .A(G110), .B(n1262), .Z(n1258) );
XNOR2_X1 U957 ( .A(G128), .B(n1263), .ZN(n1262) );
NAND2_X1 U958 ( .A1(n1264), .A2(KEYINPUT2), .ZN(n1252) );
XOR2_X1 U959 ( .A(n1265), .B(G137), .Z(n1264) );
NAND2_X1 U960 ( .A1(n1266), .A2(G221), .ZN(n1265) );
XNOR2_X1 U961 ( .A(G902), .B(KEYINPUT15), .ZN(n1251) );
INV_X1 U962 ( .A(n1084), .ZN(n1072) );
XNOR2_X1 U963 ( .A(n1267), .B(G472), .ZN(n1084) );
NAND2_X1 U964 ( .A1(n1268), .A2(n1207), .ZN(n1267) );
XOR2_X1 U965 ( .A(n1269), .B(n1270), .Z(n1268) );
XNOR2_X1 U966 ( .A(n1271), .B(n1161), .ZN(n1270) );
XNOR2_X1 U967 ( .A(n1272), .B(n1273), .ZN(n1161) );
XNOR2_X1 U968 ( .A(KEYINPUT28), .B(n1274), .ZN(n1273) );
INV_X1 U969 ( .A(G116), .ZN(n1274) );
XOR2_X1 U970 ( .A(n1275), .B(G113), .Z(n1272) );
NAND2_X1 U971 ( .A1(KEYINPUT58), .A2(n1263), .ZN(n1275) );
NAND3_X1 U972 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1271) );
NAND2_X1 U973 ( .A1(KEYINPUT43), .A2(n1165), .ZN(n1278) );
NAND3_X1 U974 ( .A1(n1279), .A2(n1280), .A3(n1164), .ZN(n1277) );
INV_X1 U975 ( .A(KEYINPUT43), .ZN(n1280) );
OR2_X1 U976 ( .A1(n1279), .A2(n1164), .ZN(n1276) );
NOR2_X1 U977 ( .A1(KEYINPUT0), .A2(n1165), .ZN(n1279) );
XNOR2_X1 U978 ( .A(G101), .B(n1169), .ZN(n1269) );
NAND2_X1 U979 ( .A1(n1281), .A2(G210), .ZN(n1169) );
NOR2_X1 U980 ( .A1(n1282), .A2(n1236), .ZN(n1059) );
XNOR2_X1 U981 ( .A(n1090), .B(n1283), .ZN(n1236) );
NOR2_X1 U982 ( .A1(G478), .A2(KEYINPUT62), .ZN(n1283) );
NOR2_X1 U983 ( .A1(n1141), .A2(G902), .ZN(n1090) );
XOR2_X1 U984 ( .A(n1284), .B(n1285), .Z(n1141) );
XOR2_X1 U985 ( .A(n1286), .B(n1287), .Z(n1285) );
NAND2_X1 U986 ( .A1(G217), .A2(n1266), .ZN(n1287) );
AND2_X1 U987 ( .A1(G234), .A2(n1104), .ZN(n1266) );
NAND2_X1 U988 ( .A1(KEYINPUT3), .A2(n1288), .ZN(n1286) );
XNOR2_X1 U989 ( .A(n1289), .B(G128), .ZN(n1288) );
XOR2_X1 U990 ( .A(n1290), .B(n1291), .Z(n1284) );
NOR2_X1 U991 ( .A1(KEYINPUT52), .A2(n1292), .ZN(n1291) );
XNOR2_X1 U992 ( .A(G116), .B(G122), .ZN(n1292) );
XNOR2_X1 U993 ( .A(G134), .B(G107), .ZN(n1290) );
XNOR2_X1 U994 ( .A(KEYINPUT21), .B(n1085), .ZN(n1282) );
XNOR2_X1 U995 ( .A(n1293), .B(G475), .ZN(n1085) );
NAND2_X1 U996 ( .A1(n1146), .A2(n1207), .ZN(n1293) );
XOR2_X1 U997 ( .A(n1294), .B(n1295), .Z(n1146) );
XOR2_X1 U998 ( .A(KEYINPUT16), .B(G122), .Z(n1295) );
XOR2_X1 U999 ( .A(n1296), .B(n1297), .Z(n1294) );
NAND2_X1 U1000 ( .A1(n1298), .A2(n1299), .ZN(n1296) );
NAND2_X1 U1001 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
XOR2_X1 U1002 ( .A(KEYINPUT51), .B(n1302), .Z(n1298) );
NOR2_X1 U1003 ( .A1(n1300), .A2(n1301), .ZN(n1302) );
XOR2_X1 U1004 ( .A(n1303), .B(n1304), .Z(n1301) );
XNOR2_X1 U1005 ( .A(n1289), .B(G131), .ZN(n1304) );
NAND2_X1 U1006 ( .A1(n1281), .A2(G214), .ZN(n1303) );
NOR2_X1 U1007 ( .A1(G953), .A2(G237), .ZN(n1281) );
XOR2_X1 U1008 ( .A(n1305), .B(n1112), .Z(n1300) );
XOR2_X1 U1009 ( .A(G140), .B(n1306), .Z(n1112) );
NAND2_X1 U1010 ( .A1(KEYINPUT13), .A2(n1307), .ZN(n1305) );
INV_X1 U1011 ( .A(G146), .ZN(n1307) );
AND3_X1 U1012 ( .A1(n1065), .A2(n1221), .A3(n1219), .ZN(n1223) );
NOR2_X1 U1013 ( .A1(n1078), .A2(n1077), .ZN(n1219) );
AND2_X1 U1014 ( .A1(G214), .A2(n1308), .ZN(n1077) );
INV_X1 U1015 ( .A(n1239), .ZN(n1078) );
XNOR2_X1 U1016 ( .A(n1309), .B(n1206), .ZN(n1239) );
AND2_X1 U1017 ( .A1(G210), .A2(n1308), .ZN(n1206) );
OR2_X1 U1018 ( .A1(G902), .A2(G237), .ZN(n1308) );
NAND2_X1 U1019 ( .A1(n1310), .A2(n1207), .ZN(n1309) );
INV_X1 U1020 ( .A(G902), .ZN(n1207) );
XNOR2_X1 U1021 ( .A(n1311), .B(n1203), .ZN(n1310) );
INV_X1 U1022 ( .A(n1198), .ZN(n1203) );
XOR2_X1 U1023 ( .A(n1129), .B(n1312), .Z(n1198) );
NOR2_X1 U1024 ( .A1(KEYINPUT53), .A2(n1128), .ZN(n1312) );
XNOR2_X1 U1025 ( .A(n1313), .B(n1314), .ZN(n1128) );
XNOR2_X1 U1026 ( .A(n1033), .B(n1315), .ZN(n1314) );
XNOR2_X1 U1027 ( .A(n1263), .B(G116), .ZN(n1315) );
INV_X1 U1028 ( .A(G119), .ZN(n1263) );
XNOR2_X1 U1029 ( .A(G101), .B(n1297), .ZN(n1313) );
XNOR2_X1 U1030 ( .A(n1316), .B(G113), .ZN(n1297) );
INV_X1 U1031 ( .A(G104), .ZN(n1316) );
XOR2_X1 U1032 ( .A(G110), .B(n1317), .Z(n1129) );
XOR2_X1 U1033 ( .A(KEYINPUT12), .B(G122), .Z(n1317) );
XOR2_X1 U1034 ( .A(n1318), .B(KEYINPUT32), .Z(n1311) );
NAND2_X1 U1035 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
NAND2_X1 U1036 ( .A1(n1321), .A2(n1205), .ZN(n1320) );
XOR2_X1 U1037 ( .A(n1322), .B(KEYINPUT57), .Z(n1319) );
OR2_X1 U1038 ( .A1(n1205), .A2(n1321), .ZN(n1322) );
XNOR2_X1 U1039 ( .A(n1204), .B(KEYINPUT48), .ZN(n1321) );
NAND2_X1 U1040 ( .A1(G224), .A2(n1104), .ZN(n1204) );
XNOR2_X1 U1041 ( .A(n1306), .B(n1167), .ZN(n1205) );
INV_X1 U1042 ( .A(n1165), .ZN(n1167) );
XOR2_X1 U1043 ( .A(G143), .B(n1323), .Z(n1165) );
XOR2_X1 U1044 ( .A(G125), .B(KEYINPUT29), .Z(n1306) );
NAND2_X1 U1045 ( .A1(n1079), .A2(n1324), .ZN(n1221) );
NAND4_X1 U1046 ( .A1(G953), .A2(G902), .A3(n1242), .A4(n1127), .ZN(n1324) );
INV_X1 U1047 ( .A(G898), .ZN(n1127) );
NAND3_X1 U1048 ( .A1(n1037), .A2(n1242), .A3(G952), .ZN(n1079) );
NAND2_X1 U1049 ( .A1(G237), .A2(G234), .ZN(n1242) );
XNOR2_X1 U1050 ( .A(G953), .B(KEYINPUT14), .ZN(n1037) );
NOR2_X1 U1051 ( .A1(n1064), .A2(n1063), .ZN(n1065) );
AND2_X1 U1052 ( .A1(G221), .A2(n1138), .ZN(n1063) );
NAND2_X1 U1053 ( .A1(n1325), .A2(G234), .ZN(n1138) );
XNOR2_X1 U1054 ( .A(G902), .B(KEYINPUT63), .ZN(n1325) );
INV_X1 U1055 ( .A(n1247), .ZN(n1064) );
XOR2_X1 U1056 ( .A(G469), .B(n1326), .Z(n1247) );
NOR2_X1 U1057 ( .A1(n1327), .A2(G902), .ZN(n1326) );
NOR2_X1 U1058 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
XOR2_X1 U1059 ( .A(KEYINPUT42), .B(n1330), .Z(n1329) );
NOR2_X1 U1060 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NOR2_X1 U1061 ( .A1(n1333), .A2(n1334), .ZN(n1331) );
NOR3_X1 U1062 ( .A1(n1334), .A2(n1335), .A3(n1333), .ZN(n1328) );
AND2_X1 U1063 ( .A1(n1179), .A2(n1336), .ZN(n1333) );
XNOR2_X1 U1064 ( .A(KEYINPUT38), .B(n1186), .ZN(n1336) );
INV_X1 U1065 ( .A(n1332), .ZN(n1335) );
NAND2_X1 U1066 ( .A1(n1337), .A2(n1338), .ZN(n1332) );
NAND2_X1 U1067 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
NAND2_X1 U1068 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
NAND2_X1 U1069 ( .A1(KEYINPUT36), .A2(n1168), .ZN(n1342) );
INV_X1 U1070 ( .A(KEYINPUT1), .ZN(n1341) );
NAND2_X1 U1071 ( .A1(n1164), .A2(n1343), .ZN(n1337) );
NAND2_X1 U1072 ( .A1(KEYINPUT36), .A2(n1344), .ZN(n1343) );
OR2_X1 U1073 ( .A1(n1339), .A2(KEYINPUT1), .ZN(n1344) );
XNOR2_X1 U1074 ( .A(n1345), .B(n1183), .ZN(n1339) );
XOR2_X1 U1075 ( .A(n1346), .B(n1347), .Z(n1183) );
NOR2_X1 U1076 ( .A1(KEYINPUT46), .A2(n1033), .ZN(n1347) );
INV_X1 U1077 ( .A(G107), .ZN(n1033) );
XNOR2_X1 U1078 ( .A(G104), .B(n1348), .ZN(n1346) );
NOR2_X1 U1079 ( .A1(G101), .A2(KEYINPUT39), .ZN(n1348) );
NAND2_X1 U1080 ( .A1(n1349), .A2(n1350), .ZN(n1345) );
NAND2_X1 U1081 ( .A1(KEYINPUT4), .A2(n1176), .ZN(n1350) );
INV_X1 U1082 ( .A(n1113), .ZN(n1176) );
NAND2_X1 U1083 ( .A1(KEYINPUT9), .A2(n1113), .ZN(n1349) );
XNOR2_X1 U1084 ( .A(n1351), .B(n1323), .ZN(n1113) );
XOR2_X1 U1085 ( .A(G128), .B(G146), .Z(n1323) );
XOR2_X1 U1086 ( .A(n1352), .B(KEYINPUT40), .Z(n1351) );
NAND2_X1 U1087 ( .A1(KEYINPUT25), .A2(n1289), .ZN(n1352) );
INV_X1 U1088 ( .A(G143), .ZN(n1289) );
INV_X1 U1089 ( .A(n1168), .ZN(n1164) );
NAND3_X1 U1090 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1168) );
NAND2_X1 U1091 ( .A1(n1356), .A2(n1110), .ZN(n1355) );
NAND2_X1 U1092 ( .A1(n1357), .A2(n1358), .ZN(n1354) );
INV_X1 U1093 ( .A(KEYINPUT54), .ZN(n1358) );
NAND2_X1 U1094 ( .A1(n1359), .A2(n1111), .ZN(n1357) );
XNOR2_X1 U1095 ( .A(KEYINPUT61), .B(n1110), .ZN(n1359) );
NAND2_X1 U1096 ( .A1(KEYINPUT54), .A2(n1360), .ZN(n1353) );
NAND2_X1 U1097 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
NAND2_X1 U1098 ( .A1(KEYINPUT61), .A2(n1110), .ZN(n1362) );
OR3_X1 U1099 ( .A1(n1356), .A2(KEYINPUT61), .A3(n1110), .ZN(n1361) );
INV_X1 U1100 ( .A(G131), .ZN(n1110) );
INV_X1 U1101 ( .A(n1111), .ZN(n1356) );
XOR2_X1 U1102 ( .A(G134), .B(G137), .Z(n1111) );
NOR2_X1 U1103 ( .A1(n1179), .A2(n1363), .ZN(n1334) );
INV_X1 U1104 ( .A(n1186), .ZN(n1363) );
NAND2_X1 U1105 ( .A1(G227), .A2(n1104), .ZN(n1186) );
INV_X1 U1106 ( .A(G953), .ZN(n1104) );
XNOR2_X1 U1107 ( .A(G110), .B(G140), .ZN(n1179) );
endmodule


