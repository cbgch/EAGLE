//Key = 0101110000101001101111011100100101011001011001010010001110100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317;

XNOR2_X1 U707 ( .A(G107), .B(n990), .ZN(G9) );
NAND4_X1 U708 ( .A1(n991), .A2(n992), .A3(n993), .A4(n994), .ZN(n990) );
AND2_X1 U709 ( .A1(n995), .A2(n996), .ZN(n993) );
XOR2_X1 U710 ( .A(n997), .B(KEYINPUT23), .Z(n991) );
NOR2_X1 U711 ( .A1(n998), .A2(n999), .ZN(G75) );
NOR4_X1 U712 ( .A1(n1000), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(n999) );
INV_X1 U713 ( .A(G952), .ZN(n1002) );
NAND3_X1 U714 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1000) );
NAND2_X1 U715 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND2_X1 U716 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND3_X1 U717 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1010) );
NAND2_X1 U718 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NAND2_X1 U719 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U720 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND2_X1 U721 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U722 ( .A1(n996), .A2(n1022), .ZN(n1014) );
NAND2_X1 U723 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U724 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND4_X1 U725 ( .A1(n1016), .A2(n996), .A3(n1027), .A4(n1028), .ZN(n1009) );
NAND2_X1 U726 ( .A1(n1029), .A2(n997), .ZN(n1028) );
NAND2_X1 U727 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND3_X1 U728 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
OR2_X1 U729 ( .A1(n1011), .A2(n1013), .ZN(n1027) );
INV_X1 U730 ( .A(n1035), .ZN(n1007) );
NOR3_X1 U731 ( .A1(n1036), .A2(G953), .A3(n1037), .ZN(n998) );
INV_X1 U732 ( .A(n1004), .ZN(n1037) );
NAND2_X1 U733 ( .A1(n1038), .A2(n1039), .ZN(n1004) );
NOR4_X1 U734 ( .A1(n1040), .A2(n1025), .A3(n1041), .A4(n1020), .ZN(n1039) );
XNOR2_X1 U735 ( .A(n1042), .B(n1043), .ZN(n1041) );
NOR2_X1 U736 ( .A1(G475), .A2(KEYINPUT38), .ZN(n1043) );
INV_X1 U737 ( .A(n1044), .ZN(n1025) );
NOR4_X1 U738 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1038) );
XNOR2_X1 U739 ( .A(G472), .B(n1049), .ZN(n1048) );
XOR2_X1 U740 ( .A(n1050), .B(n1051), .Z(n1047) );
XNOR2_X1 U741 ( .A(G469), .B(KEYINPUT43), .ZN(n1051) );
XOR2_X1 U742 ( .A(KEYINPUT48), .B(G952), .Z(n1036) );
XOR2_X1 U743 ( .A(n1052), .B(n1053), .Z(G72) );
XOR2_X1 U744 ( .A(n1054), .B(n1055), .Z(n1053) );
NOR2_X1 U745 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
XOR2_X1 U746 ( .A(n1058), .B(n1059), .Z(n1057) );
XNOR2_X1 U747 ( .A(n1060), .B(n1061), .ZN(n1059) );
NOR2_X1 U748 ( .A1(G140), .A2(KEYINPUT17), .ZN(n1061) );
NAND2_X1 U749 ( .A1(n1062), .A2(KEYINPUT63), .ZN(n1060) );
XOR2_X1 U750 ( .A(n1063), .B(KEYINPUT12), .Z(n1062) );
XOR2_X1 U751 ( .A(n1064), .B(n1065), .Z(n1058) );
NOR2_X1 U752 ( .A1(G900), .A2(n1005), .ZN(n1056) );
NOR2_X1 U753 ( .A1(G953), .A2(n1066), .ZN(n1054) );
XOR2_X1 U754 ( .A(n1001), .B(KEYINPUT36), .Z(n1066) );
NOR2_X1 U755 ( .A1(n1067), .A2(n1005), .ZN(n1052) );
AND2_X1 U756 ( .A1(G227), .A2(G900), .ZN(n1067) );
XOR2_X1 U757 ( .A(n1068), .B(n1069), .Z(G69) );
NOR2_X1 U758 ( .A1(n1070), .A2(n1005), .ZN(n1069) );
NOR2_X1 U759 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XOR2_X1 U760 ( .A(n1073), .B(KEYINPUT7), .Z(n1071) );
NAND3_X1 U761 ( .A1(n1074), .A2(n1075), .A3(KEYINPUT10), .ZN(n1068) );
NAND3_X1 U762 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NAND2_X1 U763 ( .A1(G953), .A2(n1073), .ZN(n1077) );
XOR2_X1 U764 ( .A(n1079), .B(KEYINPUT6), .Z(n1076) );
NAND2_X1 U765 ( .A1(n1005), .A2(n1003), .ZN(n1079) );
NAND3_X1 U766 ( .A1(n1003), .A2(n1005), .A3(n1080), .ZN(n1074) );
INV_X1 U767 ( .A(n1078), .ZN(n1080) );
XOR2_X1 U768 ( .A(n1081), .B(n1082), .Z(n1078) );
NAND2_X1 U769 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
XOR2_X1 U770 ( .A(n1085), .B(KEYINPUT11), .Z(n1083) );
NOR2_X1 U771 ( .A1(n1086), .A2(n1087), .ZN(G66) );
XOR2_X1 U772 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U773 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR2_X1 U774 ( .A1(n1086), .A2(n1092), .ZN(G63) );
XOR2_X1 U775 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND2_X1 U776 ( .A1(n1090), .A2(G478), .ZN(n1093) );
NOR2_X1 U777 ( .A1(n1086), .A2(n1095), .ZN(G60) );
NOR3_X1 U778 ( .A1(n1042), .A2(n1096), .A3(n1097), .ZN(n1095) );
NOR3_X1 U779 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1097) );
NOR2_X1 U780 ( .A1(n1101), .A2(n1102), .ZN(n1096) );
NOR2_X1 U781 ( .A1(n1103), .A2(n1099), .ZN(n1102) );
INV_X1 U782 ( .A(G475), .ZN(n1099) );
NOR2_X1 U783 ( .A1(n1003), .A2(n1001), .ZN(n1103) );
XOR2_X1 U784 ( .A(n1104), .B(n1105), .Z(G6) );
NOR2_X1 U785 ( .A1(n1086), .A2(n1106), .ZN(G57) );
XOR2_X1 U786 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U787 ( .A(n1109), .B(n1110), .Z(n1107) );
NOR2_X1 U788 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U789 ( .A(KEYINPUT37), .B(n1113), .Z(n1112) );
NOR2_X1 U790 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U791 ( .A1(n1116), .A2(n1117), .ZN(n1111) );
XOR2_X1 U792 ( .A(KEYINPUT25), .B(n1114), .Z(n1117) );
XOR2_X1 U793 ( .A(n1115), .B(KEYINPUT15), .Z(n1116) );
NAND2_X1 U794 ( .A1(n1090), .A2(G472), .ZN(n1115) );
NOR2_X1 U795 ( .A1(n1086), .A2(n1118), .ZN(G54) );
XOR2_X1 U796 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U797 ( .A(n1121), .B(n1122), .Z(n1120) );
NAND2_X1 U798 ( .A1(n1090), .A2(G469), .ZN(n1121) );
XOR2_X1 U799 ( .A(n1123), .B(n1124), .Z(n1119) );
XNOR2_X1 U800 ( .A(KEYINPUT40), .B(n1125), .ZN(n1124) );
NOR2_X1 U801 ( .A1(KEYINPUT59), .A2(n1126), .ZN(n1125) );
XOR2_X1 U802 ( .A(n1063), .B(n1127), .Z(n1126) );
NAND3_X1 U803 ( .A1(n1128), .A2(n1129), .A3(KEYINPUT45), .ZN(n1123) );
NAND2_X1 U804 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U805 ( .A(KEYINPUT42), .B(n1132), .Z(n1128) );
NOR2_X1 U806 ( .A1(n1131), .A2(n1130), .ZN(n1132) );
XOR2_X1 U807 ( .A(KEYINPUT29), .B(n1133), .Z(n1130) );
NOR2_X1 U808 ( .A1(n1086), .A2(n1134), .ZN(G51) );
XOR2_X1 U809 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U810 ( .A(n1137), .B(n1138), .Z(n1136) );
XNOR2_X1 U811 ( .A(n1139), .B(KEYINPUT56), .ZN(n1135) );
NAND3_X1 U812 ( .A1(n1090), .A2(n1140), .A3(KEYINPUT50), .ZN(n1139) );
INV_X1 U813 ( .A(n1100), .ZN(n1090) );
NAND2_X1 U814 ( .A1(G902), .A2(n1141), .ZN(n1100) );
OR2_X1 U815 ( .A1(n1001), .A2(n1003), .ZN(n1141) );
NAND4_X1 U816 ( .A1(n1142), .A2(n1105), .A3(n1143), .A4(n1144), .ZN(n1003) );
AND4_X1 U817 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1144) );
NOR2_X1 U818 ( .A1(n1149), .A2(n1150), .ZN(n1143) );
NOR2_X1 U819 ( .A1(n1023), .A2(n1151), .ZN(n1150) );
NOR2_X1 U820 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
NAND4_X1 U821 ( .A1(n1154), .A2(n1155), .A3(n996), .A4(n995), .ZN(n1105) );
NAND3_X1 U822 ( .A1(n1156), .A2(n1157), .A3(n1154), .ZN(n1142) );
NAND2_X1 U823 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND3_X1 U824 ( .A1(n1160), .A2(n1153), .A3(n1013), .ZN(n1159) );
INV_X1 U825 ( .A(KEYINPUT58), .ZN(n1153) );
INV_X1 U826 ( .A(n995), .ZN(n1158) );
NAND2_X1 U827 ( .A1(n1161), .A2(n995), .ZN(n1156) );
NAND2_X1 U828 ( .A1(n994), .A2(n996), .ZN(n1161) );
NAND4_X1 U829 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1001) );
AND4_X1 U830 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
AND2_X1 U831 ( .A1(n1170), .A2(n1171), .ZN(n1164) );
NAND3_X1 U832 ( .A1(n1172), .A2(n1155), .A3(n1160), .ZN(n1163) );
NAND2_X1 U833 ( .A1(n1173), .A2(n992), .ZN(n1162) );
XOR2_X1 U834 ( .A(n1174), .B(KEYINPUT28), .Z(n1173) );
NOR2_X1 U835 ( .A1(n1005), .A2(G952), .ZN(n1086) );
XOR2_X1 U836 ( .A(n1175), .B(G146), .Z(G48) );
NAND2_X1 U837 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
OR3_X1 U838 ( .A1(n1174), .A2(n1023), .A3(KEYINPUT49), .ZN(n1177) );
NAND3_X1 U839 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1174) );
NAND4_X1 U840 ( .A1(n1180), .A2(n1154), .A3(n1181), .A4(KEYINPUT49), .ZN(n1176) );
NOR3_X1 U841 ( .A1(n1032), .A2(n1182), .A3(n1021), .ZN(n1180) );
XOR2_X1 U842 ( .A(n1183), .B(n1171), .Z(G45) );
NAND3_X1 U843 ( .A1(n1160), .A2(n1154), .A3(n1184), .ZN(n1171) );
NOR3_X1 U844 ( .A1(n1185), .A2(n1181), .A3(n1186), .ZN(n1184) );
XNOR2_X1 U845 ( .A(G140), .B(n1170), .ZN(G42) );
NAND2_X1 U846 ( .A1(n1172), .A2(n1187), .ZN(n1170) );
XNOR2_X1 U847 ( .A(G137), .B(n1169), .ZN(G39) );
NAND3_X1 U848 ( .A1(n1172), .A2(n1188), .A3(n1189), .ZN(n1169) );
XNOR2_X1 U849 ( .A(G134), .B(n1168), .ZN(G36) );
NAND3_X1 U850 ( .A1(n1172), .A2(n994), .A3(n1160), .ZN(n1168) );
AND3_X1 U851 ( .A1(n1178), .A2(n1179), .A3(n1016), .ZN(n1172) );
XOR2_X1 U852 ( .A(n1190), .B(n1191), .Z(G33) );
NAND4_X1 U853 ( .A1(n1192), .A2(n1160), .A3(n1193), .A4(n1016), .ZN(n1191) );
AND2_X1 U854 ( .A1(n1194), .A2(n1044), .ZN(n1016) );
XOR2_X1 U855 ( .A(KEYINPUT47), .B(n1046), .Z(n1194) );
NOR2_X1 U856 ( .A1(n1181), .A2(n1032), .ZN(n1193) );
XOR2_X1 U857 ( .A(n997), .B(KEYINPUT20), .Z(n1192) );
XNOR2_X1 U858 ( .A(G128), .B(n1167), .ZN(G30) );
NAND3_X1 U859 ( .A1(n1154), .A2(n1188), .A3(n1195), .ZN(n1167) );
NOR3_X1 U860 ( .A1(n1034), .A2(n1181), .A3(n1182), .ZN(n1195) );
INV_X1 U861 ( .A(n1179), .ZN(n1181) );
XNOR2_X1 U862 ( .A(G101), .B(n1152), .ZN(G3) );
NAND4_X1 U863 ( .A1(n1013), .A2(n1160), .A3(n1154), .A4(n995), .ZN(n1152) );
NOR2_X1 U864 ( .A1(n1023), .A2(n997), .ZN(n1154) );
NAND2_X1 U865 ( .A1(n1196), .A2(n1197), .ZN(G27) );
OR2_X1 U866 ( .A1(n1198), .A2(G125), .ZN(n1197) );
NAND2_X1 U867 ( .A1(G125), .A2(n1199), .ZN(n1196) );
NAND2_X1 U868 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
OR2_X1 U869 ( .A1(n1166), .A2(KEYINPUT1), .ZN(n1201) );
NAND2_X1 U870 ( .A1(KEYINPUT1), .A2(n1198), .ZN(n1200) );
OR2_X1 U871 ( .A1(KEYINPUT57), .A2(n1166), .ZN(n1198) );
NAND4_X1 U872 ( .A1(n1187), .A2(n1011), .A3(n992), .A4(n1179), .ZN(n1166) );
NAND2_X1 U873 ( .A1(n1035), .A2(n1202), .ZN(n1179) );
NAND4_X1 U874 ( .A1(G953), .A2(G902), .A3(n1203), .A4(n1204), .ZN(n1202) );
XOR2_X1 U875 ( .A(KEYINPUT33), .B(G900), .Z(n1203) );
NOR3_X1 U876 ( .A1(n1182), .A2(n1188), .A3(n1032), .ZN(n1187) );
XOR2_X1 U877 ( .A(n1148), .B(n1205), .Z(G24) );
XOR2_X1 U878 ( .A(n1206), .B(KEYINPUT61), .Z(n1205) );
NAND4_X1 U879 ( .A1(n1207), .A2(n996), .A3(n1208), .A4(n1045), .ZN(n1148) );
NOR2_X1 U880 ( .A1(n1020), .A2(n1188), .ZN(n996) );
XNOR2_X1 U881 ( .A(G119), .B(n1147), .ZN(G21) );
NAND3_X1 U882 ( .A1(n1189), .A2(n1188), .A3(n1207), .ZN(n1147) );
XOR2_X1 U883 ( .A(n1146), .B(n1209), .Z(G18) );
NOR2_X1 U884 ( .A1(G116), .A2(KEYINPUT14), .ZN(n1209) );
NAND3_X1 U885 ( .A1(n1160), .A2(n994), .A3(n1207), .ZN(n1146) );
INV_X1 U886 ( .A(n1034), .ZN(n994) );
NAND2_X1 U887 ( .A1(n1185), .A2(n1045), .ZN(n1034) );
INV_X1 U888 ( .A(n1208), .ZN(n1185) );
XOR2_X1 U889 ( .A(n1210), .B(n1145), .Z(G15) );
NAND3_X1 U890 ( .A1(n1160), .A2(n1155), .A3(n1207), .ZN(n1145) );
AND3_X1 U891 ( .A1(n992), .A2(n995), .A3(n1011), .ZN(n1207) );
NOR2_X1 U892 ( .A1(n1211), .A2(n1040), .ZN(n1011) );
INV_X1 U893 ( .A(n1033), .ZN(n1040) );
INV_X1 U894 ( .A(n1023), .ZN(n992) );
INV_X1 U895 ( .A(n1032), .ZN(n1155) );
NAND2_X1 U896 ( .A1(n1186), .A2(n1208), .ZN(n1032) );
INV_X1 U897 ( .A(n1018), .ZN(n1160) );
NAND2_X1 U898 ( .A1(n1188), .A2(n1182), .ZN(n1018) );
INV_X1 U899 ( .A(n1021), .ZN(n1188) );
XOR2_X1 U900 ( .A(G110), .B(n1212), .Z(G12) );
NOR2_X1 U901 ( .A1(n1213), .A2(n1023), .ZN(n1212) );
NAND2_X1 U902 ( .A1(n1046), .A2(n1044), .ZN(n1023) );
NAND2_X1 U903 ( .A1(G214), .A2(n1214), .ZN(n1044) );
INV_X1 U904 ( .A(n1026), .ZN(n1046) );
XOR2_X1 U905 ( .A(n1215), .B(n1140), .Z(n1026) );
AND2_X1 U906 ( .A1(G210), .A2(n1214), .ZN(n1140) );
NAND2_X1 U907 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
NAND3_X1 U908 ( .A1(n1218), .A2(n1219), .A3(n1217), .ZN(n1215) );
NAND2_X1 U909 ( .A1(n1138), .A2(n1137), .ZN(n1219) );
INV_X1 U910 ( .A(n1220), .ZN(n1137) );
NAND2_X1 U911 ( .A1(n1221), .A2(n1220), .ZN(n1218) );
XNOR2_X1 U912 ( .A(n1064), .B(n1222), .ZN(n1220) );
XNOR2_X1 U913 ( .A(KEYINPUT27), .B(n1138), .ZN(n1221) );
XOR2_X1 U914 ( .A(n1223), .B(n1082), .Z(n1138) );
XOR2_X1 U915 ( .A(G110), .B(G122), .Z(n1082) );
XOR2_X1 U916 ( .A(n1224), .B(n1225), .Z(n1223) );
NOR2_X1 U917 ( .A1(G953), .A2(n1072), .ZN(n1225) );
INV_X1 U918 ( .A(G224), .ZN(n1072) );
NAND2_X1 U919 ( .A1(n1084), .A2(n1085), .ZN(n1224) );
NAND2_X1 U920 ( .A1(n1226), .A2(n1227), .ZN(n1085) );
XOR2_X1 U921 ( .A(G113), .B(n1228), .Z(n1227) );
XNOR2_X1 U922 ( .A(KEYINPUT52), .B(n1229), .ZN(n1226) );
NAND2_X1 U923 ( .A1(n1230), .A2(n1231), .ZN(n1084) );
XOR2_X1 U924 ( .A(KEYINPUT52), .B(n1229), .Z(n1231) );
XOR2_X1 U925 ( .A(n1210), .B(n1228), .Z(n1230) );
NOR2_X1 U926 ( .A1(KEYINPUT60), .A2(n1232), .ZN(n1228) );
XOR2_X1 U927 ( .A(n1151), .B(KEYINPUT44), .Z(n1213) );
NAND4_X1 U928 ( .A1(n1189), .A2(n1178), .A3(n1021), .A4(n995), .ZN(n1151) );
NAND2_X1 U929 ( .A1(n1035), .A2(n1233), .ZN(n995) );
NAND4_X1 U930 ( .A1(G953), .A2(G902), .A3(n1204), .A4(n1073), .ZN(n1233) );
INV_X1 U931 ( .A(G898), .ZN(n1073) );
NAND3_X1 U932 ( .A1(n1204), .A2(n1005), .A3(G952), .ZN(n1035) );
NAND2_X1 U933 ( .A1(G237), .A2(G234), .ZN(n1204) );
NAND3_X1 U934 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1021) );
NAND2_X1 U935 ( .A1(G472), .A2(n1237), .ZN(n1236) );
NAND2_X1 U936 ( .A1(n1238), .A2(n1049), .ZN(n1237) );
INV_X1 U937 ( .A(n1239), .ZN(n1238) );
NAND3_X1 U938 ( .A1(n1239), .A2(n1049), .A3(n1240), .ZN(n1235) );
XOR2_X1 U939 ( .A(n1241), .B(G472), .Z(n1239) );
XNOR2_X1 U940 ( .A(KEYINPUT41), .B(KEYINPUT21), .ZN(n1241) );
OR2_X1 U941 ( .A1(n1049), .A2(n1240), .ZN(n1234) );
INV_X1 U942 ( .A(KEYINPUT51), .ZN(n1240) );
NAND2_X1 U943 ( .A1(n1242), .A2(n1217), .ZN(n1049) );
XOR2_X1 U944 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U945 ( .A(n1114), .B(n1109), .Z(n1244) );
NAND3_X1 U946 ( .A1(n1216), .A2(n1005), .A3(G210), .ZN(n1109) );
XNOR2_X1 U947 ( .A(n1245), .B(n1232), .ZN(n1114) );
XOR2_X1 U948 ( .A(G116), .B(G119), .Z(n1232) );
XOR2_X1 U949 ( .A(n1246), .B(n1247), .Z(n1245) );
NAND2_X1 U950 ( .A1(KEYINPUT16), .A2(n1210), .ZN(n1246) );
INV_X1 U951 ( .A(G113), .ZN(n1210) );
XNOR2_X1 U952 ( .A(KEYINPUT34), .B(n1248), .ZN(n1243) );
NOR2_X1 U953 ( .A1(KEYINPUT30), .A2(n1108), .ZN(n1248) );
INV_X1 U954 ( .A(n997), .ZN(n1178) );
NAND2_X1 U955 ( .A1(n1211), .A2(n1033), .ZN(n997) );
NAND2_X1 U956 ( .A1(G221), .A2(n1249), .ZN(n1033) );
INV_X1 U957 ( .A(n1030), .ZN(n1211) );
XNOR2_X1 U958 ( .A(n1250), .B(n1050), .ZN(n1030) );
NAND2_X1 U959 ( .A1(n1251), .A2(n1217), .ZN(n1050) );
XOR2_X1 U960 ( .A(n1252), .B(n1253), .Z(n1251) );
XNOR2_X1 U961 ( .A(n1127), .B(n1131), .ZN(n1253) );
XOR2_X1 U962 ( .A(G110), .B(n1254), .Z(n1131) );
XOR2_X1 U963 ( .A(KEYINPUT31), .B(G140), .Z(n1254) );
XNOR2_X1 U964 ( .A(n1229), .B(KEYINPUT18), .ZN(n1127) );
XNOR2_X1 U965 ( .A(n1255), .B(n1108), .ZN(n1229) );
XOR2_X1 U966 ( .A(G101), .B(KEYINPUT2), .Z(n1108) );
XOR2_X1 U967 ( .A(n1104), .B(G107), .Z(n1255) );
XOR2_X1 U968 ( .A(n1247), .B(n1256), .Z(n1252) );
XOR2_X1 U969 ( .A(KEYINPUT40), .B(n1133), .Z(n1256) );
AND2_X1 U970 ( .A1(G227), .A2(n1005), .ZN(n1133) );
XOR2_X1 U971 ( .A(n1065), .B(n1222), .Z(n1247) );
INV_X1 U972 ( .A(n1063), .ZN(n1222) );
XOR2_X1 U973 ( .A(n1257), .B(n1258), .Z(n1063) );
XOR2_X1 U974 ( .A(n1259), .B(G143), .Z(n1257) );
INV_X1 U975 ( .A(n1122), .ZN(n1065) );
XOR2_X1 U976 ( .A(n1260), .B(n1261), .Z(n1122) );
INV_X1 U977 ( .A(n1262), .ZN(n1261) );
XOR2_X1 U978 ( .A(n1190), .B(G134), .Z(n1260) );
INV_X1 U979 ( .A(G131), .ZN(n1190) );
NAND2_X1 U980 ( .A1(KEYINPUT39), .A2(G469), .ZN(n1250) );
AND2_X1 U981 ( .A1(n1013), .A2(n1020), .ZN(n1189) );
INV_X1 U982 ( .A(n1182), .ZN(n1020) );
XOR2_X1 U983 ( .A(n1263), .B(n1091), .Z(n1182) );
AND2_X1 U984 ( .A1(G217), .A2(n1249), .ZN(n1091) );
NAND2_X1 U985 ( .A1(G234), .A2(n1264), .ZN(n1249) );
XOR2_X1 U986 ( .A(KEYINPUT19), .B(G902), .Z(n1264) );
NAND2_X1 U987 ( .A1(n1089), .A2(n1217), .ZN(n1263) );
XNOR2_X1 U988 ( .A(n1265), .B(n1266), .ZN(n1089) );
XOR2_X1 U989 ( .A(n1262), .B(n1267), .Z(n1266) );
XOR2_X1 U990 ( .A(n1268), .B(n1269), .Z(n1267) );
AND2_X1 U991 ( .A1(n1270), .A2(G221), .ZN(n1269) );
NAND2_X1 U992 ( .A1(n1271), .A2(KEYINPUT5), .ZN(n1268) );
XOR2_X1 U993 ( .A(n1272), .B(KEYINPUT26), .Z(n1271) );
XNOR2_X1 U994 ( .A(G137), .B(KEYINPUT22), .ZN(n1262) );
XOR2_X1 U995 ( .A(n1273), .B(n1274), .Z(n1265) );
XOR2_X1 U996 ( .A(G146), .B(G119), .Z(n1274) );
XOR2_X1 U997 ( .A(n1275), .B(G110), .Z(n1273) );
NAND2_X1 U998 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XNOR2_X1 U999 ( .A(KEYINPUT24), .B(n1278), .ZN(n1276) );
NOR2_X1 U1000 ( .A1(n1045), .A2(n1208), .ZN(n1013) );
XOR2_X1 U1001 ( .A(n1042), .B(G475), .Z(n1208) );
NOR2_X1 U1002 ( .A1(n1101), .A2(G902), .ZN(n1042) );
INV_X1 U1003 ( .A(n1098), .ZN(n1101) );
NAND2_X1 U1004 ( .A1(n1279), .A2(n1280), .ZN(n1098) );
NAND2_X1 U1005 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XOR2_X1 U1006 ( .A(n1283), .B(KEYINPUT13), .Z(n1279) );
OR2_X1 U1007 ( .A1(n1282), .A2(n1281), .ZN(n1283) );
XOR2_X1 U1008 ( .A(n1284), .B(n1285), .Z(n1281) );
NOR2_X1 U1009 ( .A1(KEYINPUT8), .A2(n1104), .ZN(n1285) );
INV_X1 U1010 ( .A(G104), .ZN(n1104) );
XOR2_X1 U1011 ( .A(n1206), .B(n1286), .Z(n1284) );
NOR2_X1 U1012 ( .A1(G113), .A2(KEYINPUT0), .ZN(n1286) );
INV_X1 U1013 ( .A(G122), .ZN(n1206) );
NAND2_X1 U1014 ( .A1(n1287), .A2(n1288), .ZN(n1282) );
NAND3_X1 U1015 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1288) );
INV_X1 U1016 ( .A(n1292), .ZN(n1291) );
XOR2_X1 U1017 ( .A(n1293), .B(KEYINPUT32), .Z(n1287) );
NAND2_X1 U1018 ( .A1(n1292), .A2(n1294), .ZN(n1293) );
NAND2_X1 U1019 ( .A1(n1289), .A2(n1290), .ZN(n1294) );
NAND2_X1 U1020 ( .A1(n1295), .A2(n1259), .ZN(n1290) );
INV_X1 U1021 ( .A(G146), .ZN(n1259) );
XOR2_X1 U1022 ( .A(KEYINPUT53), .B(n1296), .Z(n1295) );
AND2_X1 U1023 ( .A1(n1278), .A2(n1277), .ZN(n1296) );
NAND2_X1 U1024 ( .A1(G146), .A2(n1297), .ZN(n1289) );
NAND2_X1 U1025 ( .A1(n1278), .A2(n1277), .ZN(n1297) );
NAND2_X1 U1026 ( .A1(n1298), .A2(n1064), .ZN(n1277) );
XNOR2_X1 U1027 ( .A(KEYINPUT4), .B(G140), .ZN(n1298) );
NAND2_X1 U1028 ( .A1(n1299), .A2(n1300), .ZN(n1278) );
INV_X1 U1029 ( .A(n1064), .ZN(n1300) );
XNOR2_X1 U1030 ( .A(G125), .B(KEYINPUT9), .ZN(n1064) );
XOR2_X1 U1031 ( .A(KEYINPUT4), .B(G140), .Z(n1299) );
XOR2_X1 U1032 ( .A(n1301), .B(n1302), .Z(n1292) );
XOR2_X1 U1033 ( .A(KEYINPUT62), .B(G131), .Z(n1302) );
NAND3_X1 U1034 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(n1301) );
NAND4_X1 U1035 ( .A1(G214), .A2(n1306), .A3(n1216), .A4(n1005), .ZN(n1305) );
NAND2_X1 U1036 ( .A1(KEYINPUT35), .A2(n1307), .ZN(n1306) );
NAND2_X1 U1037 ( .A1(KEYINPUT54), .A2(G143), .ZN(n1307) );
OR2_X1 U1038 ( .A1(n1183), .A2(KEYINPUT35), .ZN(n1304) );
NAND3_X1 U1039 ( .A1(n1308), .A2(n1183), .A3(KEYINPUT35), .ZN(n1303) );
INV_X1 U1040 ( .A(G143), .ZN(n1183) );
NAND4_X1 U1041 ( .A1(KEYINPUT54), .A2(G214), .A3(n1216), .A4(n1005), .ZN(n1308) );
INV_X1 U1042 ( .A(G237), .ZN(n1216) );
INV_X1 U1043 ( .A(n1186), .ZN(n1045) );
XOR2_X1 U1044 ( .A(n1309), .B(G478), .Z(n1186) );
NAND2_X1 U1045 ( .A1(n1094), .A2(n1217), .ZN(n1309) );
INV_X1 U1046 ( .A(G902), .ZN(n1217) );
XNOR2_X1 U1047 ( .A(n1310), .B(n1311), .ZN(n1094) );
XOR2_X1 U1048 ( .A(G107), .B(n1312), .Z(n1311) );
XOR2_X1 U1049 ( .A(G143), .B(G134), .Z(n1312) );
XOR2_X1 U1050 ( .A(n1313), .B(n1314), .Z(n1310) );
XOR2_X1 U1051 ( .A(n1315), .B(n1316), .Z(n1314) );
NAND2_X1 U1052 ( .A1(G217), .A2(n1270), .ZN(n1316) );
AND2_X1 U1053 ( .A1(G234), .A2(n1005), .ZN(n1270) );
INV_X1 U1054 ( .A(G953), .ZN(n1005) );
NAND2_X1 U1055 ( .A1(KEYINPUT55), .A2(n1317), .ZN(n1315) );
XOR2_X1 U1056 ( .A(G122), .B(G116), .Z(n1317) );
NAND2_X1 U1057 ( .A1(KEYINPUT3), .A2(n1258), .ZN(n1313) );
INV_X1 U1058 ( .A(n1272), .ZN(n1258) );
XNOR2_X1 U1059 ( .A(G128), .B(KEYINPUT46), .ZN(n1272) );
endmodule


