//Key = 0010000011000011001010111011000101011110001100010100111111010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342;

XNOR2_X1 U743 ( .A(G107), .B(n1028), .ZN(G9) );
NOR2_X1 U744 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U745 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
XOR2_X1 U746 ( .A(KEYINPUT34), .B(n1035), .Z(n1032) );
NOR4_X1 U747 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
NAND3_X1 U748 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1036) );
NAND4_X1 U749 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1031) );
NAND4_X1 U750 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1042), .ZN(n1044) );
NAND3_X1 U751 ( .A1(n1050), .A2(n1041), .A3(n1051), .ZN(n1043) );
NAND2_X1 U752 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NAND3_X1 U753 ( .A1(n1054), .A2(n1040), .A3(n1042), .ZN(n1053) );
NAND2_X1 U754 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U755 ( .A1(n1049), .A2(n1057), .ZN(n1056) );
XOR2_X1 U756 ( .A(n1058), .B(n1059), .Z(n1057) );
NOR2_X1 U757 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
INV_X1 U758 ( .A(KEYINPUT63), .ZN(n1060) );
NAND2_X1 U759 ( .A1(n1048), .A2(n1062), .ZN(n1055) );
NAND3_X1 U760 ( .A1(n1048), .A2(n1049), .A3(n1047), .ZN(n1052) );
AND3_X1 U761 ( .A1(n1063), .A2(n1064), .A3(n1040), .ZN(n1047) );
NAND4_X1 U762 ( .A1(n1065), .A2(n1066), .A3(n1051), .A4(n1041), .ZN(n1064) );
NAND2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1063) );
INV_X1 U764 ( .A(n1041), .ZN(n1068) );
XOR2_X1 U765 ( .A(KEYINPUT58), .B(n1039), .Z(n1067) );
AND3_X1 U766 ( .A1(n1045), .A2(n1046), .A3(n1069), .ZN(n1029) );
NAND4_X1 U767 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1045) );
NOR4_X1 U768 ( .A1(n1074), .A2(n1059), .A3(n1039), .A4(n1075), .ZN(n1073) );
XOR2_X1 U769 ( .A(n1076), .B(n1077), .Z(n1075) );
NAND2_X1 U770 ( .A1(KEYINPUT55), .A2(G475), .ZN(n1077) );
XOR2_X1 U771 ( .A(n1078), .B(G478), .Z(n1072) );
NAND2_X1 U772 ( .A1(KEYINPUT33), .A2(n1079), .ZN(n1078) );
XNOR2_X1 U773 ( .A(n1080), .B(KEYINPUT17), .ZN(n1071) );
XOR2_X1 U774 ( .A(n1081), .B(n1082), .Z(n1070) );
NOR2_X1 U775 ( .A1(KEYINPUT30), .A2(n1083), .ZN(n1082) );
XOR2_X1 U776 ( .A(n1084), .B(n1085), .Z(G72) );
XOR2_X1 U777 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND2_X1 U778 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NAND2_X1 U779 ( .A1(G900), .A2(G227), .ZN(n1088) );
NAND2_X1 U780 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NAND2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U782 ( .A(n1093), .B(n1094), .Z(n1089) );
XNOR2_X1 U783 ( .A(n1095), .B(n1096), .ZN(n1094) );
XOR2_X1 U784 ( .A(KEYINPUT22), .B(G140), .Z(n1093) );
AND2_X1 U785 ( .A1(n1034), .A2(n1046), .ZN(n1084) );
NAND2_X1 U786 ( .A1(n1097), .A2(n1098), .ZN(G69) );
NAND4_X1 U787 ( .A1(G953), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1098) );
INV_X1 U788 ( .A(KEYINPUT4), .ZN(n1101) );
NAND4_X1 U789 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1097) );
NAND3_X1 U790 ( .A1(n1106), .A2(n1033), .A3(n1046), .ZN(n1105) );
NAND2_X1 U791 ( .A1(G953), .A2(n1107), .ZN(n1104) );
NAND2_X1 U792 ( .A1(n1106), .A2(n1108), .ZN(n1107) );
NAND2_X1 U793 ( .A1(n1109), .A2(n1099), .ZN(n1108) );
INV_X1 U794 ( .A(n1100), .ZN(n1106) );
NAND2_X1 U795 ( .A1(KEYINPUT6), .A2(n1109), .ZN(n1103) );
NAND3_X1 U796 ( .A1(n1110), .A2(n1099), .A3(G953), .ZN(n1109) );
NAND2_X1 U797 ( .A1(G898), .A2(G224), .ZN(n1099) );
OR2_X1 U798 ( .A1(KEYINPUT4), .A2(KEYINPUT6), .ZN(n1110) );
NAND2_X1 U799 ( .A1(n1111), .A2(n1100), .ZN(n1102) );
NAND2_X1 U800 ( .A1(n1112), .A2(n1113), .ZN(n1100) );
NAND2_X1 U801 ( .A1(n1092), .A2(n1114), .ZN(n1113) );
XOR2_X1 U802 ( .A(n1115), .B(n1116), .Z(n1112) );
NAND2_X1 U803 ( .A1(KEYINPUT57), .A2(n1117), .ZN(n1115) );
NOR2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(G66) );
NOR2_X1 U805 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U806 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U807 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NOR2_X1 U808 ( .A1(n1126), .A2(n1127), .ZN(n1122) );
INV_X1 U809 ( .A(KEYINPUT59), .ZN(n1127) );
XOR2_X1 U810 ( .A(n1128), .B(KEYINPUT54), .Z(n1126) );
NOR2_X1 U811 ( .A1(KEYINPUT59), .A2(n1129), .ZN(n1120) );
XOR2_X1 U812 ( .A(KEYINPUT54), .B(n1130), .Z(n1129) );
INV_X1 U813 ( .A(n1128), .ZN(n1130) );
NOR2_X1 U814 ( .A1(n1118), .A2(n1131), .ZN(G63) );
XOR2_X1 U815 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U816 ( .A1(n1134), .A2(n1125), .ZN(n1132) );
INV_X1 U817 ( .A(G478), .ZN(n1134) );
NOR2_X1 U818 ( .A1(n1118), .A2(n1135), .ZN(G60) );
XNOR2_X1 U819 ( .A(n1136), .B(n1137), .ZN(n1135) );
NOR2_X1 U820 ( .A1(n1138), .A2(n1125), .ZN(n1137) );
INV_X1 U821 ( .A(G475), .ZN(n1138) );
XOR2_X1 U822 ( .A(G104), .B(n1139), .Z(G6) );
NOR3_X1 U823 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(G57) );
AND2_X1 U824 ( .A1(KEYINPUT14), .A2(n1118), .ZN(n1142) );
NOR3_X1 U825 ( .A1(KEYINPUT14), .A2(G952), .A3(n1143), .ZN(n1141) );
XOR2_X1 U826 ( .A(n1144), .B(n1145), .Z(n1140) );
XOR2_X1 U827 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U828 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U829 ( .A1(n1083), .A2(n1125), .ZN(n1149) );
INV_X1 U830 ( .A(G472), .ZN(n1083) );
NAND3_X1 U831 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1146) );
NAND2_X1 U832 ( .A1(KEYINPUT32), .A2(n1153), .ZN(n1152) );
NAND3_X1 U833 ( .A1(n1154), .A2(n1155), .A3(n1096), .ZN(n1151) );
INV_X1 U834 ( .A(KEYINPUT32), .ZN(n1155) );
OR2_X1 U835 ( .A1(n1096), .A2(n1154), .ZN(n1150) );
NOR2_X1 U836 ( .A1(KEYINPUT11), .A2(n1153), .ZN(n1154) );
XNOR2_X1 U837 ( .A(n1156), .B(n1157), .ZN(n1144) );
NOR2_X1 U838 ( .A1(KEYINPUT45), .A2(n1158), .ZN(n1157) );
NOR2_X1 U839 ( .A1(n1118), .A2(n1159), .ZN(G54) );
XOR2_X1 U840 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U841 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U842 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
OR2_X1 U843 ( .A1(n1166), .A2(n1096), .ZN(n1165) );
NAND2_X1 U844 ( .A1(n1096), .A2(n1167), .ZN(n1164) );
XOR2_X1 U845 ( .A(n1166), .B(n1168), .Z(n1167) );
XOR2_X1 U846 ( .A(KEYINPUT41), .B(KEYINPUT39), .Z(n1168) );
NAND2_X1 U847 ( .A1(n1169), .A2(n1170), .ZN(n1166) );
XNOR2_X1 U848 ( .A(KEYINPUT49), .B(n1171), .ZN(n1169) );
XOR2_X1 U849 ( .A(n1172), .B(n1173), .Z(n1160) );
NOR2_X1 U850 ( .A1(n1174), .A2(n1125), .ZN(n1173) );
NAND2_X1 U851 ( .A1(KEYINPUT8), .A2(n1175), .ZN(n1172) );
NOR2_X1 U852 ( .A1(n1118), .A2(n1176), .ZN(G51) );
XOR2_X1 U853 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U854 ( .A(n1179), .B(n1180), .Z(n1177) );
NOR2_X1 U855 ( .A1(n1181), .A2(n1125), .ZN(n1180) );
NAND2_X1 U856 ( .A1(G902), .A2(n1182), .ZN(n1125) );
NAND2_X1 U857 ( .A1(n1111), .A2(n1183), .ZN(n1182) );
XNOR2_X1 U858 ( .A(KEYINPUT50), .B(n1034), .ZN(n1183) );
NAND2_X1 U859 ( .A1(n1184), .A2(n1185), .ZN(n1034) );
NOR4_X1 U860 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1185) );
NOR2_X1 U861 ( .A1(KEYINPUT1), .A2(n1190), .ZN(n1186) );
NOR4_X1 U862 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1184) );
NOR2_X1 U863 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NOR2_X1 U864 ( .A1(n1197), .A2(n1198), .ZN(n1195) );
AND3_X1 U865 ( .A1(KEYINPUT1), .A2(n1038), .A3(n1199), .ZN(n1198) );
INV_X1 U866 ( .A(n1033), .ZN(n1111) );
NAND4_X1 U867 ( .A1(n1200), .A2(n1028), .A3(n1201), .A4(n1202), .ZN(n1033) );
NOR4_X1 U868 ( .A1(n1139), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1202) );
NOR2_X1 U869 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NOR2_X1 U870 ( .A1(n1208), .A2(n1209), .ZN(n1206) );
AND2_X1 U871 ( .A1(n1197), .A2(KEYINPUT56), .ZN(n1209) );
NOR2_X1 U872 ( .A1(n1210), .A2(n1211), .ZN(n1208) );
NOR3_X1 U873 ( .A1(n1065), .A2(n1212), .A3(n1213), .ZN(n1204) );
XNOR2_X1 U874 ( .A(n1049), .B(KEYINPUT19), .ZN(n1212) );
NOR4_X1 U875 ( .A1(KEYINPUT56), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1203) );
NOR3_X1 U876 ( .A1(n1210), .A2(n1213), .A3(n1038), .ZN(n1139) );
AND2_X1 U877 ( .A1(n1217), .A2(n1218), .ZN(n1201) );
NAND3_X1 U878 ( .A1(n1062), .A2(n1219), .A3(n1042), .ZN(n1028) );
NAND2_X1 U879 ( .A1(n1220), .A2(KEYINPUT42), .ZN(n1179) );
XOR2_X1 U880 ( .A(n1221), .B(n1222), .Z(n1220) );
XOR2_X1 U881 ( .A(n1223), .B(n1224), .Z(n1222) );
INV_X1 U882 ( .A(G125), .ZN(n1223) );
NAND2_X1 U883 ( .A1(KEYINPUT26), .A2(n1225), .ZN(n1221) );
AND2_X1 U884 ( .A1(n1143), .A2(n1069), .ZN(n1118) );
INV_X1 U885 ( .A(G952), .ZN(n1069) );
XOR2_X1 U886 ( .A(G953), .B(KEYINPUT28), .Z(n1143) );
XOR2_X1 U887 ( .A(G146), .B(n1192), .Z(G48) );
AND3_X1 U888 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1192) );
XOR2_X1 U889 ( .A(G143), .B(n1191), .Z(G45) );
NOR3_X1 U890 ( .A1(n1229), .A2(n1065), .A3(n1211), .ZN(n1191) );
INV_X1 U891 ( .A(n1199), .ZN(n1065) );
XOR2_X1 U892 ( .A(G140), .B(n1189), .Z(G42) );
NOR3_X1 U893 ( .A1(n1038), .A2(n1196), .A3(n1066), .ZN(n1189) );
XOR2_X1 U894 ( .A(n1188), .B(n1230), .Z(G39) );
XOR2_X1 U895 ( .A(KEYINPUT16), .B(G137), .Z(n1230) );
AND3_X1 U896 ( .A1(n1226), .A2(n1231), .A3(n1049), .ZN(n1188) );
XOR2_X1 U897 ( .A(G134), .B(n1232), .Z(G36) );
NOR2_X1 U898 ( .A1(n1196), .A2(n1216), .ZN(n1232) );
XOR2_X1 U899 ( .A(n1190), .B(n1233), .Z(G33) );
NAND2_X1 U900 ( .A1(n1234), .A2(KEYINPUT15), .ZN(n1233) );
XNOR2_X1 U901 ( .A(G131), .B(KEYINPUT37), .ZN(n1234) );
NAND3_X1 U902 ( .A1(n1199), .A2(n1231), .A3(n1227), .ZN(n1190) );
INV_X1 U903 ( .A(n1196), .ZN(n1231) );
NAND4_X1 U904 ( .A1(n1051), .A2(n1235), .A3(n1059), .A4(n1236), .ZN(n1196) );
XNOR2_X1 U905 ( .A(n1187), .B(n1237), .ZN(G30) );
NAND2_X1 U906 ( .A1(KEYINPUT35), .A2(G128), .ZN(n1237) );
AND3_X1 U907 ( .A1(n1226), .A2(n1062), .A3(n1228), .ZN(n1187) );
INV_X1 U908 ( .A(n1229), .ZN(n1228) );
NAND4_X1 U909 ( .A1(n1235), .A2(n1059), .A3(n1039), .A4(n1236), .ZN(n1229) );
XNOR2_X1 U910 ( .A(G101), .B(n1238), .ZN(G3) );
NAND2_X1 U911 ( .A1(n1239), .A2(n1199), .ZN(n1238) );
XOR2_X1 U912 ( .A(n1240), .B(n1241), .Z(G27) );
XOR2_X1 U913 ( .A(KEYINPUT27), .B(G125), .Z(n1241) );
NAND2_X1 U914 ( .A1(KEYINPUT43), .A2(n1193), .ZN(n1240) );
AND4_X1 U915 ( .A1(n1242), .A2(n1243), .A3(n1227), .A4(n1236), .ZN(n1193) );
NAND2_X1 U916 ( .A1(n1244), .A2(n1245), .ZN(n1236) );
NAND2_X1 U917 ( .A1(n1091), .A2(n1246), .ZN(n1245) );
XNOR2_X1 U918 ( .A(G900), .B(KEYINPUT25), .ZN(n1091) );
XOR2_X1 U919 ( .A(n1247), .B(n1248), .Z(G24) );
NOR3_X1 U920 ( .A1(n1207), .A2(n1249), .A3(n1210), .ZN(n1248) );
INV_X1 U921 ( .A(n1042), .ZN(n1210) );
NOR2_X1 U922 ( .A1(n1250), .A2(n1080), .ZN(n1042) );
XOR2_X1 U923 ( .A(n1211), .B(KEYINPUT12), .Z(n1249) );
NAND2_X1 U924 ( .A1(n1251), .A2(n1252), .ZN(n1211) );
XOR2_X1 U925 ( .A(n1253), .B(KEYINPUT38), .Z(n1247) );
XOR2_X1 U926 ( .A(n1254), .B(n1218), .Z(G21) );
NAND3_X1 U927 ( .A1(n1049), .A2(n1226), .A3(n1255), .ZN(n1218) );
AND2_X1 U928 ( .A1(n1080), .A2(n1250), .ZN(n1226) );
INV_X1 U929 ( .A(n1256), .ZN(n1250) );
XNOR2_X1 U930 ( .A(G116), .B(n1257), .ZN(G18) );
NAND3_X1 U931 ( .A1(n1197), .A2(n1255), .A3(KEYINPUT23), .ZN(n1257) );
INV_X1 U932 ( .A(n1216), .ZN(n1197) );
NAND2_X1 U933 ( .A1(n1199), .A2(n1062), .ZN(n1216) );
NOR2_X1 U934 ( .A1(n1252), .A2(n1258), .ZN(n1062) );
XOR2_X1 U935 ( .A(n1259), .B(n1217), .Z(G15) );
NAND3_X1 U936 ( .A1(n1227), .A2(n1199), .A3(n1255), .ZN(n1217) );
INV_X1 U937 ( .A(n1207), .ZN(n1255) );
NAND2_X1 U938 ( .A1(n1242), .A2(n1215), .ZN(n1207) );
INV_X1 U939 ( .A(n1214), .ZN(n1242) );
NAND3_X1 U940 ( .A1(n1039), .A2(n1041), .A3(n1048), .ZN(n1214) );
INV_X1 U941 ( .A(n1037), .ZN(n1048) );
NAND2_X1 U942 ( .A1(n1260), .A2(n1061), .ZN(n1037) );
XOR2_X1 U943 ( .A(KEYINPUT63), .B(n1059), .Z(n1260) );
NOR2_X1 U944 ( .A1(n1080), .A2(n1256), .ZN(n1199) );
INV_X1 U945 ( .A(n1038), .ZN(n1227) );
NAND2_X1 U946 ( .A1(n1258), .A2(n1252), .ZN(n1038) );
INV_X1 U947 ( .A(n1251), .ZN(n1258) );
XOR2_X1 U948 ( .A(n1200), .B(n1261), .Z(G12) );
NOR2_X1 U949 ( .A1(G110), .A2(KEYINPUT21), .ZN(n1261) );
NAND2_X1 U950 ( .A1(n1239), .A2(n1243), .ZN(n1200) );
INV_X1 U951 ( .A(n1066), .ZN(n1243) );
NAND2_X1 U952 ( .A1(n1256), .A2(n1080), .ZN(n1066) );
XOR2_X1 U953 ( .A(n1262), .B(n1124), .Z(n1080) );
NAND2_X1 U954 ( .A1(G217), .A2(n1263), .ZN(n1124) );
NAND2_X1 U955 ( .A1(n1128), .A2(n1264), .ZN(n1262) );
XOR2_X1 U956 ( .A(n1265), .B(n1266), .Z(n1128) );
XNOR2_X1 U957 ( .A(n1163), .B(n1267), .ZN(n1266) );
XOR2_X1 U958 ( .A(n1268), .B(n1269), .Z(n1267) );
NAND2_X1 U959 ( .A1(KEYINPUT53), .A2(n1270), .ZN(n1268) );
NAND3_X1 U960 ( .A1(G234), .A2(n1046), .A3(G221), .ZN(n1270) );
XOR2_X1 U961 ( .A(n1271), .B(n1272), .Z(n1265) );
XOR2_X1 U962 ( .A(G125), .B(G119), .Z(n1272) );
XOR2_X1 U963 ( .A(n1273), .B(KEYINPUT5), .Z(n1271) );
INV_X1 U964 ( .A(G137), .ZN(n1273) );
XOR2_X1 U965 ( .A(n1081), .B(G472), .Z(n1256) );
NAND2_X1 U966 ( .A1(n1274), .A2(n1264), .ZN(n1081) );
XOR2_X1 U967 ( .A(n1275), .B(n1276), .Z(n1274) );
XNOR2_X1 U968 ( .A(n1096), .B(n1153), .ZN(n1276) );
XOR2_X1 U969 ( .A(n1225), .B(KEYINPUT31), .Z(n1153) );
XOR2_X1 U970 ( .A(n1158), .B(n1277), .Z(n1275) );
XNOR2_X1 U971 ( .A(n1148), .B(n1278), .ZN(n1277) );
NOR2_X1 U972 ( .A1(KEYINPUT0), .A2(n1156), .ZN(n1278) );
XNOR2_X1 U973 ( .A(n1279), .B(n1280), .ZN(n1156) );
XOR2_X1 U974 ( .A(G116), .B(n1281), .Z(n1280) );
NOR2_X1 U975 ( .A1(KEYINPUT10), .A2(n1259), .ZN(n1281) );
INV_X1 U976 ( .A(G113), .ZN(n1259) );
NAND2_X1 U977 ( .A1(KEYINPUT52), .A2(n1254), .ZN(n1279) );
INV_X1 U978 ( .A(G119), .ZN(n1254) );
NAND2_X1 U979 ( .A1(G210), .A2(n1282), .ZN(n1148) );
AND2_X1 U980 ( .A1(n1049), .A2(n1219), .ZN(n1239) );
INV_X1 U981 ( .A(n1213), .ZN(n1219) );
NAND4_X1 U982 ( .A1(n1235), .A2(n1059), .A3(n1039), .A4(n1215), .ZN(n1213) );
NAND2_X1 U983 ( .A1(n1244), .A2(n1283), .ZN(n1215) );
NAND2_X1 U984 ( .A1(n1246), .A2(n1114), .ZN(n1283) );
INV_X1 U985 ( .A(G898), .ZN(n1114) );
AND3_X1 U986 ( .A1(n1092), .A2(n1040), .A3(G902), .ZN(n1246) );
XOR2_X1 U987 ( .A(n1046), .B(KEYINPUT24), .Z(n1092) );
NAND2_X1 U988 ( .A1(n1284), .A2(n1040), .ZN(n1244) );
NAND2_X1 U989 ( .A1(G237), .A2(G234), .ZN(n1040) );
AND2_X1 U990 ( .A1(n1285), .A2(G952), .ZN(n1284) );
XOR2_X1 U991 ( .A(n1046), .B(KEYINPUT60), .Z(n1285) );
INV_X1 U992 ( .A(n1051), .ZN(n1039) );
XNOR2_X1 U993 ( .A(n1286), .B(n1181), .ZN(n1051) );
NAND2_X1 U994 ( .A1(G210), .A2(n1287), .ZN(n1181) );
NAND3_X1 U995 ( .A1(n1288), .A2(n1264), .A3(n1289), .ZN(n1286) );
XOR2_X1 U996 ( .A(n1290), .B(KEYINPUT13), .Z(n1289) );
NAND2_X1 U997 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XNOR2_X1 U998 ( .A(n1224), .B(n1293), .ZN(n1292) );
XOR2_X1 U999 ( .A(KEYINPUT48), .B(n1178), .Z(n1291) );
NAND2_X1 U1000 ( .A1(n1294), .A2(n1295), .ZN(n1288) );
XOR2_X1 U1001 ( .A(n1224), .B(n1293), .Z(n1295) );
NOR2_X1 U1002 ( .A1(KEYINPUT44), .A2(n1095), .ZN(n1293) );
XOR2_X1 U1003 ( .A(G125), .B(n1225), .Z(n1095) );
NAND2_X1 U1004 ( .A1(n1296), .A2(n1046), .ZN(n1224) );
XNOR2_X1 U1005 ( .A(G224), .B(KEYINPUT2), .ZN(n1296) );
XNOR2_X1 U1006 ( .A(KEYINPUT48), .B(n1178), .ZN(n1294) );
XNOR2_X1 U1007 ( .A(n1117), .B(n1297), .ZN(n1178) );
NOR2_X1 U1008 ( .A1(KEYINPUT61), .A2(n1116), .ZN(n1297) );
NAND2_X1 U1009 ( .A1(n1298), .A2(n1299), .ZN(n1116) );
NAND2_X1 U1010 ( .A1(n1300), .A2(n1253), .ZN(n1299) );
INV_X1 U1011 ( .A(G122), .ZN(n1253) );
XOR2_X1 U1012 ( .A(KEYINPUT18), .B(G110), .Z(n1300) );
NAND2_X1 U1013 ( .A1(G122), .A2(n1301), .ZN(n1298) );
XNOR2_X1 U1014 ( .A(G110), .B(KEYINPUT47), .ZN(n1301) );
XOR2_X1 U1015 ( .A(n1302), .B(n1303), .Z(n1117) );
XOR2_X1 U1016 ( .A(G113), .B(n1304), .Z(n1303) );
XOR2_X1 U1017 ( .A(G119), .B(G116), .Z(n1304) );
XOR2_X1 U1018 ( .A(n1158), .B(n1305), .Z(n1302) );
NOR2_X1 U1019 ( .A1(KEYINPUT29), .A2(n1306), .ZN(n1305) );
XOR2_X1 U1020 ( .A(n1307), .B(n1174), .Z(n1059) );
INV_X1 U1021 ( .A(G469), .ZN(n1174) );
NAND2_X1 U1022 ( .A1(n1308), .A2(n1264), .ZN(n1307) );
XNOR2_X1 U1023 ( .A(n1096), .B(n1309), .ZN(n1308) );
XOR2_X1 U1024 ( .A(n1310), .B(n1311), .Z(n1309) );
NOR2_X1 U1025 ( .A1(KEYINPUT46), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U1026 ( .A(n1175), .B(n1163), .ZN(n1312) );
XOR2_X1 U1027 ( .A(G110), .B(G140), .Z(n1163) );
AND2_X1 U1028 ( .A1(G227), .A2(n1046), .ZN(n1175) );
NAND2_X1 U1029 ( .A1(n1171), .A2(n1170), .ZN(n1310) );
NAND2_X1 U1030 ( .A1(n1313), .A2(n1314), .ZN(n1170) );
XOR2_X1 U1031 ( .A(n1315), .B(n1158), .Z(n1314) );
XOR2_X1 U1032 ( .A(KEYINPUT22), .B(n1316), .Z(n1313) );
INV_X1 U1033 ( .A(n1225), .ZN(n1316) );
NAND2_X1 U1034 ( .A1(n1317), .A2(n1318), .ZN(n1171) );
XOR2_X1 U1035 ( .A(n1315), .B(n1319), .Z(n1318) );
INV_X1 U1036 ( .A(n1158), .ZN(n1319) );
XNOR2_X1 U1037 ( .A(G101), .B(KEYINPUT7), .ZN(n1158) );
NAND2_X1 U1038 ( .A1(n1320), .A2(KEYINPUT9), .ZN(n1315) );
XOR2_X1 U1039 ( .A(n1306), .B(KEYINPUT3), .Z(n1320) );
XNOR2_X1 U1040 ( .A(G104), .B(n1321), .ZN(n1306) );
XOR2_X1 U1041 ( .A(KEYINPUT51), .B(G107), .Z(n1321) );
XOR2_X1 U1042 ( .A(n1225), .B(KEYINPUT22), .Z(n1317) );
XOR2_X1 U1043 ( .A(n1322), .B(n1269), .Z(n1225) );
XOR2_X1 U1044 ( .A(G128), .B(G146), .Z(n1269) );
XOR2_X1 U1045 ( .A(G131), .B(n1323), .Z(n1096) );
XOR2_X1 U1046 ( .A(G137), .B(G134), .Z(n1323) );
INV_X1 U1047 ( .A(n1074), .ZN(n1235) );
NAND2_X1 U1048 ( .A1(n1061), .A2(n1041), .ZN(n1074) );
NAND2_X1 U1049 ( .A1(G214), .A2(n1287), .ZN(n1041) );
NAND2_X1 U1050 ( .A1(n1324), .A2(n1264), .ZN(n1287) );
INV_X1 U1051 ( .A(G237), .ZN(n1324) );
NAND2_X1 U1052 ( .A1(G221), .A2(n1263), .ZN(n1061) );
NAND2_X1 U1053 ( .A1(G234), .A2(n1264), .ZN(n1263) );
NOR2_X1 U1054 ( .A1(n1251), .A2(n1252), .ZN(n1049) );
XNOR2_X1 U1055 ( .A(n1076), .B(G475), .ZN(n1252) );
NAND2_X1 U1056 ( .A1(n1136), .A2(n1264), .ZN(n1076) );
INV_X1 U1057 ( .A(G902), .ZN(n1264) );
XNOR2_X1 U1058 ( .A(n1325), .B(n1326), .ZN(n1136) );
XOR2_X1 U1059 ( .A(G140), .B(G131), .Z(n1326) );
XOR2_X1 U1060 ( .A(n1327), .B(n1328), .Z(n1325) );
XOR2_X1 U1061 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1062 ( .A(G143), .B(G122), .Z(n1330) );
XOR2_X1 U1063 ( .A(KEYINPUT20), .B(G146), .Z(n1329) );
XOR2_X1 U1064 ( .A(n1331), .B(n1332), .Z(n1327) );
XOR2_X1 U1065 ( .A(G113), .B(G104), .Z(n1332) );
XOR2_X1 U1066 ( .A(n1333), .B(n1334), .Z(n1331) );
NOR2_X1 U1067 ( .A1(G125), .A2(KEYINPUT62), .ZN(n1334) );
NAND2_X1 U1068 ( .A1(G214), .A2(n1282), .ZN(n1333) );
NOR2_X1 U1069 ( .A1(G953), .A2(G237), .ZN(n1282) );
XOR2_X1 U1070 ( .A(n1079), .B(G478), .Z(n1251) );
NOR2_X1 U1071 ( .A1(n1133), .A2(G902), .ZN(n1079) );
XNOR2_X1 U1072 ( .A(n1335), .B(n1336), .ZN(n1133) );
XOR2_X1 U1073 ( .A(n1337), .B(n1338), .Z(n1336) );
XOR2_X1 U1074 ( .A(G107), .B(n1339), .Z(n1338) );
NOR2_X1 U1075 ( .A1(G128), .A2(n1340), .ZN(n1339) );
XNOR2_X1 U1076 ( .A(KEYINPUT40), .B(KEYINPUT36), .ZN(n1340) );
AND3_X1 U1077 ( .A1(G217), .A2(n1046), .A3(G234), .ZN(n1337) );
INV_X1 U1078 ( .A(G953), .ZN(n1046) );
XOR2_X1 U1079 ( .A(n1341), .B(n1342), .Z(n1335) );
XOR2_X1 U1080 ( .A(G122), .B(G116), .Z(n1342) );
XOR2_X1 U1081 ( .A(G134), .B(n1322), .Z(n1341) );
INV_X1 U1082 ( .A(G143), .ZN(n1322) );
endmodule


