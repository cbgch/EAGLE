//Key = 0110111110000010100111011110000010111001011100110111101101001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501;

XOR2_X1 U820 ( .A(G107), .B(n1153), .Z(G9) );
NOR3_X1 U821 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1153) );
XNOR2_X1 U822 ( .A(n1157), .B(KEYINPUT30), .ZN(n1155) );
NOR2_X1 U823 ( .A1(n1158), .A2(n1159), .ZN(G75) );
NOR4_X1 U824 ( .A1(G953), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1159) );
XOR2_X1 U825 ( .A(KEYINPUT39), .B(n1163), .Z(n1162) );
NOR3_X1 U826 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1163) );
NOR3_X1 U827 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1166) );
NOR2_X1 U828 ( .A1(n1170), .A2(n1171), .ZN(n1168) );
NOR2_X1 U829 ( .A1(n1172), .A2(n1156), .ZN(n1171) );
NOR2_X1 U830 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NOR2_X1 U831 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NOR2_X1 U832 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
NOR2_X1 U833 ( .A1(n1179), .A2(n1180), .ZN(n1177) );
NOR2_X1 U834 ( .A1(n1181), .A2(n1182), .ZN(n1173) );
NOR2_X1 U835 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
NOR2_X1 U836 ( .A1(n1185), .A2(n1186), .ZN(n1183) );
NOR3_X1 U837 ( .A1(n1182), .A2(n1187), .A3(n1176), .ZN(n1170) );
NOR2_X1 U838 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NOR3_X1 U839 ( .A1(n1190), .A2(n1191), .A3(n1182), .ZN(n1165) );
NOR2_X1 U840 ( .A1(n1192), .A2(n1157), .ZN(n1191) );
NOR2_X1 U841 ( .A1(KEYINPUT15), .A2(n1193), .ZN(n1192) );
NOR3_X1 U842 ( .A1(n1194), .A2(n1195), .A3(n1182), .ZN(n1164) );
NOR2_X1 U843 ( .A1(n1193), .A2(n1190), .ZN(n1195) );
OR3_X1 U844 ( .A1(n1176), .A2(n1156), .A3(n1167), .ZN(n1190) );
INV_X1 U845 ( .A(KEYINPUT15), .ZN(n1194) );
NOR3_X1 U846 ( .A1(n1160), .A2(G953), .A3(G952), .ZN(n1158) );
AND4_X1 U847 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1160) );
NOR4_X1 U848 ( .A1(n1200), .A2(n1156), .A3(n1201), .A4(n1202), .ZN(n1199) );
XOR2_X1 U849 ( .A(n1203), .B(n1204), .Z(n1202) );
XOR2_X1 U850 ( .A(G478), .B(n1205), .Z(n1201) );
INV_X1 U851 ( .A(n1206), .ZN(n1156) );
NOR2_X1 U852 ( .A1(n1207), .A2(n1208), .ZN(n1200) );
XOR2_X1 U853 ( .A(n1209), .B(KEYINPUT37), .Z(n1208) );
AND3_X1 U854 ( .A1(n1186), .A2(n1210), .A3(n1179), .ZN(n1198) );
XOR2_X1 U855 ( .A(n1211), .B(n1212), .Z(G72) );
NOR2_X1 U856 ( .A1(n1213), .A2(G953), .ZN(n1212) );
XOR2_X1 U857 ( .A(n1214), .B(n1215), .Z(n1211) );
NOR2_X1 U858 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
XOR2_X1 U859 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U860 ( .A(n1220), .B(n1221), .Z(n1219) );
NAND2_X1 U861 ( .A1(n1222), .A2(n1223), .ZN(n1218) );
NAND2_X1 U862 ( .A1(n1224), .A2(G137), .ZN(n1223) );
NAND2_X1 U863 ( .A1(n1225), .A2(n1226), .ZN(n1222) );
XNOR2_X1 U864 ( .A(n1224), .B(KEYINPUT28), .ZN(n1225) );
NOR2_X1 U865 ( .A1(G900), .A2(n1227), .ZN(n1216) );
XOR2_X1 U866 ( .A(n1228), .B(KEYINPUT40), .Z(n1227) );
NAND2_X1 U867 ( .A1(KEYINPUT57), .A2(n1229), .ZN(n1214) );
NAND2_X1 U868 ( .A1(G953), .A2(n1230), .ZN(n1229) );
NAND2_X1 U869 ( .A1(G900), .A2(G227), .ZN(n1230) );
NAND3_X1 U870 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(G69) );
OR2_X1 U871 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND3_X1 U872 ( .A1(n1235), .A2(n1234), .A3(G953), .ZN(n1232) );
NAND2_X1 U873 ( .A1(G898), .A2(G224), .ZN(n1235) );
NAND2_X1 U874 ( .A1(n1236), .A2(n1228), .ZN(n1231) );
NAND2_X1 U875 ( .A1(n1234), .A2(n1237), .ZN(n1236) );
NAND2_X1 U876 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
OR2_X1 U877 ( .A1(n1238), .A2(n1240), .ZN(n1234) );
XNOR2_X1 U878 ( .A(KEYINPUT49), .B(n1241), .ZN(n1240) );
NOR2_X1 U879 ( .A1(n1242), .A2(G953), .ZN(n1241) );
NAND2_X1 U880 ( .A1(n1243), .A2(n1244), .ZN(n1238) );
NAND2_X1 U881 ( .A1(G953), .A2(n1245), .ZN(n1244) );
XOR2_X1 U882 ( .A(n1246), .B(n1247), .Z(n1243) );
NOR2_X1 U883 ( .A1(KEYINPUT59), .A2(n1248), .ZN(n1246) );
NOR2_X1 U884 ( .A1(n1249), .A2(n1250), .ZN(G66) );
XOR2_X1 U885 ( .A(n1251), .B(n1252), .Z(n1250) );
XOR2_X1 U886 ( .A(KEYINPUT43), .B(n1253), .Z(n1252) );
NOR2_X1 U887 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NOR2_X1 U888 ( .A1(n1249), .A2(n1256), .ZN(G63) );
NOR3_X1 U889 ( .A1(n1205), .A2(n1257), .A3(n1258), .ZN(n1256) );
AND3_X1 U890 ( .A1(n1259), .A2(G478), .A3(n1260), .ZN(n1258) );
NOR2_X1 U891 ( .A1(n1261), .A2(n1259), .ZN(n1257) );
AND2_X1 U892 ( .A1(n1161), .A2(G478), .ZN(n1261) );
NOR2_X1 U893 ( .A1(n1249), .A2(n1262), .ZN(G60) );
NOR3_X1 U894 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1262) );
NOR3_X1 U895 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(n1265) );
AND2_X1 U896 ( .A1(n1266), .A2(n1268), .ZN(n1264) );
NAND2_X1 U897 ( .A1(n1269), .A2(G475), .ZN(n1268) );
XOR2_X1 U898 ( .A(n1161), .B(KEYINPUT0), .Z(n1269) );
XOR2_X1 U899 ( .A(G104), .B(n1270), .Z(G6) );
NOR2_X1 U900 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NOR2_X1 U901 ( .A1(n1273), .A2(n1274), .ZN(G57) );
XOR2_X1 U902 ( .A(n1275), .B(n1276), .Z(n1274) );
XOR2_X1 U903 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U904 ( .A(n1279), .B(n1280), .Z(n1275) );
XOR2_X1 U905 ( .A(n1281), .B(n1282), .Z(n1280) );
AND2_X1 U906 ( .A1(G472), .A2(n1260), .ZN(n1282) );
INV_X1 U907 ( .A(n1255), .ZN(n1260) );
NOR2_X1 U908 ( .A1(n1283), .A2(n1284), .ZN(n1281) );
XOR2_X1 U909 ( .A(n1285), .B(KEYINPUT55), .Z(n1284) );
NAND2_X1 U910 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U911 ( .A(n1288), .B(KEYINPUT13), .Z(n1286) );
NOR2_X1 U912 ( .A1(n1287), .A2(n1288), .ZN(n1283) );
XOR2_X1 U913 ( .A(n1289), .B(KEYINPUT11), .Z(n1287) );
NAND2_X1 U914 ( .A1(KEYINPUT20), .A2(n1290), .ZN(n1279) );
NOR2_X1 U915 ( .A1(n1291), .A2(n1228), .ZN(n1273) );
XNOR2_X1 U916 ( .A(G952), .B(KEYINPUT60), .ZN(n1291) );
NOR2_X1 U917 ( .A1(n1249), .A2(n1292), .ZN(G54) );
XOR2_X1 U918 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U919 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U920 ( .A(n1297), .B(n1220), .Z(n1296) );
XOR2_X1 U921 ( .A(n1298), .B(n1299), .Z(n1295) );
NOR2_X1 U922 ( .A1(n1203), .A2(n1255), .ZN(n1298) );
INV_X1 U923 ( .A(G469), .ZN(n1203) );
XOR2_X1 U924 ( .A(n1300), .B(n1301), .Z(n1293) );
XOR2_X1 U925 ( .A(G110), .B(n1302), .Z(n1301) );
XOR2_X1 U926 ( .A(KEYINPUT1), .B(G140), .Z(n1300) );
NOR2_X1 U927 ( .A1(n1249), .A2(n1303), .ZN(G51) );
XOR2_X1 U928 ( .A(n1304), .B(n1305), .Z(n1303) );
NOR2_X1 U929 ( .A1(n1209), .A2(n1255), .ZN(n1305) );
NAND2_X1 U930 ( .A1(G902), .A2(n1161), .ZN(n1255) );
NAND2_X1 U931 ( .A1(n1242), .A2(n1213), .ZN(n1161) );
AND4_X1 U932 ( .A1(n1306), .A2(n1307), .A3(n1308), .A4(n1309), .ZN(n1213) );
AND4_X1 U933 ( .A1(n1310), .A2(n1311), .A3(n1312), .A4(n1313), .ZN(n1309) );
INV_X1 U934 ( .A(n1314), .ZN(n1312) );
NOR2_X1 U935 ( .A1(n1315), .A2(n1316), .ZN(n1308) );
NOR2_X1 U936 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
INV_X1 U937 ( .A(KEYINPUT6), .ZN(n1317) );
NOR3_X1 U938 ( .A1(KEYINPUT6), .A2(n1319), .A3(n1182), .ZN(n1315) );
NAND2_X1 U939 ( .A1(n1320), .A2(n1321), .ZN(n1307) );
NAND3_X1 U940 ( .A1(n1322), .A2(n1323), .A3(n1324), .ZN(n1321) );
NAND3_X1 U941 ( .A1(n1325), .A2(n1326), .A3(n1327), .ZN(n1324) );
NAND3_X1 U942 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1323) );
XOR2_X1 U943 ( .A(KEYINPUT46), .B(n1331), .Z(n1330) );
XOR2_X1 U944 ( .A(KEYINPUT38), .B(n1327), .Z(n1329) );
NAND4_X1 U945 ( .A1(n1332), .A2(n1189), .A3(n1271), .A4(n1333), .ZN(n1322) );
OR2_X1 U946 ( .A1(n1333), .A2(n1334), .ZN(n1306) );
INV_X1 U947 ( .A(KEYINPUT19), .ZN(n1333) );
INV_X1 U948 ( .A(n1239), .ZN(n1242) );
NAND4_X1 U949 ( .A1(n1335), .A2(n1336), .A3(n1337), .A4(n1338), .ZN(n1239) );
NOR4_X1 U950 ( .A1(n1339), .A2(n1340), .A3(n1341), .A4(n1342), .ZN(n1338) );
NAND2_X1 U951 ( .A1(n1178), .A2(n1343), .ZN(n1337) );
XNOR2_X1 U952 ( .A(KEYINPUT22), .B(n1272), .ZN(n1343) );
NAND4_X1 U953 ( .A1(n1328), .A2(n1206), .A3(n1184), .A4(n1344), .ZN(n1272) );
NAND3_X1 U954 ( .A1(n1325), .A2(n1326), .A3(n1345), .ZN(n1336) );
NAND2_X1 U955 ( .A1(n1206), .A2(n1346), .ZN(n1335) );
NAND2_X1 U956 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
NAND2_X1 U957 ( .A1(n1332), .A2(n1345), .ZN(n1348) );
NAND2_X1 U958 ( .A1(n1349), .A2(n1157), .ZN(n1347) );
INV_X1 U959 ( .A(n1154), .ZN(n1349) );
NOR2_X1 U960 ( .A1(n1228), .A2(G952), .ZN(n1249) );
XOR2_X1 U961 ( .A(n1350), .B(n1313), .Z(G48) );
NAND3_X1 U962 ( .A1(n1328), .A2(n1326), .A3(n1351), .ZN(n1313) );
XNOR2_X1 U963 ( .A(G143), .B(n1334), .ZN(G45) );
NAND3_X1 U964 ( .A1(n1332), .A2(n1189), .A3(n1351), .ZN(n1334) );
INV_X1 U965 ( .A(n1352), .ZN(n1332) );
XOR2_X1 U966 ( .A(G140), .B(n1314), .Z(G42) );
NOR2_X1 U967 ( .A1(n1353), .A2(n1354), .ZN(n1314) );
XOR2_X1 U968 ( .A(n1226), .B(n1355), .Z(G39) );
NAND4_X1 U969 ( .A1(n1356), .A2(n1327), .A3(n1320), .A4(n1325), .ZN(n1355) );
XNOR2_X1 U970 ( .A(KEYINPUT42), .B(n1326), .ZN(n1356) );
XOR2_X1 U971 ( .A(n1318), .B(n1357), .Z(G36) );
XOR2_X1 U972 ( .A(KEYINPUT14), .B(G134), .Z(n1357) );
NAND2_X1 U973 ( .A1(n1319), .A2(n1327), .ZN(n1318) );
AND3_X1 U974 ( .A1(n1157), .A2(n1189), .A3(n1320), .ZN(n1319) );
XOR2_X1 U975 ( .A(G131), .B(n1358), .Z(G33) );
NOR2_X1 U976 ( .A1(n1331), .A2(n1353), .ZN(n1358) );
NAND3_X1 U977 ( .A1(n1320), .A2(n1328), .A3(n1327), .ZN(n1353) );
INV_X1 U978 ( .A(n1182), .ZN(n1327) );
NAND2_X1 U979 ( .A1(n1359), .A2(n1360), .ZN(n1182) );
INV_X1 U980 ( .A(n1180), .ZN(n1359) );
NAND2_X1 U981 ( .A1(n1361), .A2(n1362), .ZN(G30) );
NAND2_X1 U982 ( .A1(G128), .A2(n1311), .ZN(n1362) );
XOR2_X1 U983 ( .A(n1363), .B(KEYINPUT45), .Z(n1361) );
OR2_X1 U984 ( .A1(n1311), .A2(G128), .ZN(n1363) );
NAND3_X1 U985 ( .A1(n1157), .A2(n1326), .A3(n1351), .ZN(n1311) );
AND2_X1 U986 ( .A1(n1320), .A2(n1178), .ZN(n1351) );
AND2_X1 U987 ( .A1(n1184), .A2(n1364), .ZN(n1320) );
XOR2_X1 U988 ( .A(G101), .B(n1342), .Z(G3) );
NOR3_X1 U989 ( .A1(n1154), .A2(n1331), .A3(n1169), .ZN(n1342) );
INV_X1 U990 ( .A(n1189), .ZN(n1331) );
XNOR2_X1 U991 ( .A(G125), .B(n1310), .ZN(G27) );
NAND4_X1 U992 ( .A1(n1178), .A2(n1364), .A3(n1188), .A4(n1365), .ZN(n1310) );
NOR2_X1 U993 ( .A1(n1176), .A2(n1193), .ZN(n1365) );
NAND2_X1 U994 ( .A1(n1366), .A2(n1167), .ZN(n1364) );
NAND4_X1 U995 ( .A1(G953), .A2(G902), .A3(n1367), .A4(n1368), .ZN(n1366) );
INV_X1 U996 ( .A(G900), .ZN(n1368) );
XNOR2_X1 U997 ( .A(G122), .B(n1369), .ZN(G24) );
NAND4_X1 U998 ( .A1(n1178), .A2(n1370), .A3(n1206), .A4(n1371), .ZN(n1369) );
NOR2_X1 U999 ( .A1(n1176), .A2(n1352), .ZN(n1371) );
NAND2_X1 U1000 ( .A1(n1372), .A2(n1373), .ZN(n1352) );
XNOR2_X1 U1001 ( .A(KEYINPUT4), .B(n1344), .ZN(n1370) );
XOR2_X1 U1002 ( .A(n1374), .B(n1375), .Z(G21) );
XOR2_X1 U1003 ( .A(n1376), .B(KEYINPUT17), .Z(n1375) );
NAND4_X1 U1004 ( .A1(n1377), .A2(n1325), .A3(n1378), .A4(n1379), .ZN(n1374) );
XOR2_X1 U1005 ( .A(KEYINPUT29), .B(n1178), .Z(n1379) );
AND2_X1 U1006 ( .A1(n1344), .A2(n1326), .ZN(n1378) );
NAND2_X1 U1007 ( .A1(n1380), .A2(n1381), .ZN(n1326) );
NAND3_X1 U1008 ( .A1(n1382), .A2(n1383), .A3(n1384), .ZN(n1381) );
NAND2_X1 U1009 ( .A1(KEYINPUT10), .A2(n1188), .ZN(n1380) );
INV_X1 U1010 ( .A(n1169), .ZN(n1325) );
XOR2_X1 U1011 ( .A(G116), .B(n1341), .Z(G18) );
AND3_X1 U1012 ( .A1(n1157), .A2(n1189), .A3(n1345), .ZN(n1341) );
AND2_X1 U1013 ( .A1(n1385), .A2(n1372), .ZN(n1157) );
NAND2_X1 U1014 ( .A1(n1386), .A2(n1387), .ZN(G15) );
NAND2_X1 U1015 ( .A1(n1340), .A2(n1388), .ZN(n1387) );
XOR2_X1 U1016 ( .A(KEYINPUT7), .B(n1389), .Z(n1386) );
NOR2_X1 U1017 ( .A1(n1340), .A2(n1388), .ZN(n1389) );
AND3_X1 U1018 ( .A1(n1328), .A2(n1189), .A3(n1345), .ZN(n1340) );
AND3_X1 U1019 ( .A1(n1178), .A2(n1344), .A3(n1377), .ZN(n1345) );
INV_X1 U1020 ( .A(n1176), .ZN(n1377) );
NAND2_X1 U1021 ( .A1(n1390), .A2(n1186), .ZN(n1176) );
INV_X1 U1022 ( .A(n1185), .ZN(n1390) );
NAND2_X1 U1023 ( .A1(n1391), .A2(n1392), .ZN(n1189) );
NAND3_X1 U1024 ( .A1(n1383), .A2(n1393), .A3(n1384), .ZN(n1392) );
INV_X1 U1025 ( .A(KEYINPUT10), .ZN(n1384) );
NAND2_X1 U1026 ( .A1(KEYINPUT10), .A2(n1206), .ZN(n1391) );
NOR2_X1 U1027 ( .A1(n1383), .A2(n1382), .ZN(n1206) );
INV_X1 U1028 ( .A(n1393), .ZN(n1382) );
INV_X1 U1029 ( .A(n1193), .ZN(n1328) );
NAND2_X1 U1030 ( .A1(n1394), .A2(n1373), .ZN(n1193) );
XOR2_X1 U1031 ( .A(G110), .B(n1339), .Z(G12) );
NOR3_X1 U1032 ( .A1(n1169), .A2(n1154), .A3(n1354), .ZN(n1339) );
INV_X1 U1033 ( .A(n1188), .ZN(n1354) );
NOR2_X1 U1034 ( .A1(n1383), .A2(n1393), .ZN(n1188) );
XNOR2_X1 U1035 ( .A(n1395), .B(n1254), .ZN(n1393) );
NAND2_X1 U1036 ( .A1(G217), .A2(n1396), .ZN(n1254) );
NAND2_X1 U1037 ( .A1(n1251), .A2(n1267), .ZN(n1395) );
XNOR2_X1 U1038 ( .A(n1397), .B(n1398), .ZN(n1251) );
XOR2_X1 U1039 ( .A(n1399), .B(n1400), .Z(n1398) );
NAND2_X1 U1040 ( .A1(KEYINPUT47), .A2(n1376), .ZN(n1400) );
INV_X1 U1041 ( .A(G119), .ZN(n1376) );
NAND3_X1 U1042 ( .A1(n1401), .A2(n1402), .A3(n1403), .ZN(n1399) );
NAND2_X1 U1043 ( .A1(KEYINPUT33), .A2(n1404), .ZN(n1403) );
NAND3_X1 U1044 ( .A1(n1405), .A2(n1406), .A3(n1226), .ZN(n1402) );
INV_X1 U1045 ( .A(KEYINPUT33), .ZN(n1406) );
OR2_X1 U1046 ( .A1(n1226), .A2(n1405), .ZN(n1401) );
NOR2_X1 U1047 ( .A1(KEYINPUT3), .A2(n1404), .ZN(n1405) );
NAND3_X1 U1048 ( .A1(G234), .A2(n1228), .A3(G221), .ZN(n1404) );
XOR2_X1 U1049 ( .A(n1407), .B(n1408), .Z(n1397) );
NOR2_X1 U1050 ( .A1(KEYINPUT44), .A2(n1409), .ZN(n1408) );
XNOR2_X1 U1051 ( .A(n1221), .B(n1410), .ZN(n1409) );
NOR2_X1 U1052 ( .A1(KEYINPUT12), .A2(n1350), .ZN(n1410) );
INV_X1 U1053 ( .A(G146), .ZN(n1350) );
XOR2_X1 U1054 ( .A(G125), .B(G140), .Z(n1221) );
XOR2_X1 U1055 ( .A(G128), .B(n1411), .Z(n1407) );
XNOR2_X1 U1056 ( .A(n1412), .B(G472), .ZN(n1383) );
NAND2_X1 U1057 ( .A1(n1413), .A2(n1267), .ZN(n1412) );
XOR2_X1 U1058 ( .A(n1414), .B(n1415), .Z(n1413) );
XOR2_X1 U1059 ( .A(n1278), .B(n1290), .Z(n1415) );
XOR2_X1 U1060 ( .A(n1416), .B(G113), .Z(n1278) );
NAND2_X1 U1061 ( .A1(KEYINPUT21), .A2(n1417), .ZN(n1416) );
XOR2_X1 U1062 ( .A(n1418), .B(n1419), .Z(n1414) );
NOR2_X1 U1063 ( .A1(KEYINPUT9), .A2(n1277), .ZN(n1419) );
XOR2_X1 U1064 ( .A(n1289), .B(G101), .Z(n1418) );
NAND2_X1 U1065 ( .A1(n1420), .A2(G210), .ZN(n1289) );
NAND3_X1 U1066 ( .A1(n1178), .A2(n1344), .A3(n1184), .ZN(n1154) );
AND2_X1 U1067 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND2_X1 U1068 ( .A1(G221), .A2(n1396), .ZN(n1186) );
NAND2_X1 U1069 ( .A1(G234), .A2(n1267), .ZN(n1396) );
NAND2_X1 U1070 ( .A1(n1421), .A2(n1422), .ZN(n1185) );
NAND2_X1 U1071 ( .A1(G469), .A2(n1204), .ZN(n1422) );
XOR2_X1 U1072 ( .A(n1423), .B(KEYINPUT56), .Z(n1421) );
NAND2_X1 U1073 ( .A1(n1424), .A2(n1425), .ZN(n1423) );
XOR2_X1 U1074 ( .A(KEYINPUT32), .B(G469), .Z(n1425) );
INV_X1 U1075 ( .A(n1204), .ZN(n1424) );
NAND2_X1 U1076 ( .A1(n1426), .A2(n1267), .ZN(n1204) );
XOR2_X1 U1077 ( .A(n1427), .B(n1428), .Z(n1426) );
XOR2_X1 U1078 ( .A(n1429), .B(n1430), .Z(n1428) );
XNOR2_X1 U1079 ( .A(n1302), .B(KEYINPUT8), .ZN(n1430) );
AND2_X1 U1080 ( .A1(G227), .A2(n1228), .ZN(n1302) );
NAND2_X1 U1081 ( .A1(KEYINPUT24), .A2(n1297), .ZN(n1429) );
XOR2_X1 U1082 ( .A(n1288), .B(n1431), .Z(n1297) );
XOR2_X1 U1083 ( .A(G107), .B(G104), .Z(n1431) );
INV_X1 U1084 ( .A(G101), .ZN(n1288) );
XOR2_X1 U1085 ( .A(n1432), .B(n1433), .Z(n1427) );
INV_X1 U1086 ( .A(n1220), .ZN(n1433) );
XOR2_X1 U1087 ( .A(n1434), .B(n1435), .Z(n1220) );
XOR2_X1 U1088 ( .A(G146), .B(G128), .Z(n1435) );
NAND2_X1 U1089 ( .A1(KEYINPUT35), .A2(G143), .ZN(n1434) );
XOR2_X1 U1090 ( .A(n1436), .B(n1299), .Z(n1432) );
INV_X1 U1091 ( .A(n1277), .ZN(n1299) );
XOR2_X1 U1092 ( .A(n1226), .B(n1224), .Z(n1277) );
XOR2_X1 U1093 ( .A(G131), .B(G134), .Z(n1224) );
INV_X1 U1094 ( .A(G137), .ZN(n1226) );
NAND3_X1 U1095 ( .A1(n1437), .A2(n1438), .A3(KEYINPUT50), .ZN(n1436) );
NAND2_X1 U1096 ( .A1(G140), .A2(n1411), .ZN(n1438) );
XOR2_X1 U1097 ( .A(KEYINPUT51), .B(n1439), .Z(n1437) );
NOR2_X1 U1098 ( .A1(G140), .A2(n1411), .ZN(n1439) );
INV_X1 U1099 ( .A(G110), .ZN(n1411) );
NAND2_X1 U1100 ( .A1(n1167), .A2(n1440), .ZN(n1344) );
NAND4_X1 U1101 ( .A1(G953), .A2(G902), .A3(n1367), .A4(n1245), .ZN(n1440) );
INV_X1 U1102 ( .A(G898), .ZN(n1245) );
NAND3_X1 U1103 ( .A1(n1367), .A2(n1228), .A3(G952), .ZN(n1167) );
NAND2_X1 U1104 ( .A1(G237), .A2(G234), .ZN(n1367) );
INV_X1 U1105 ( .A(n1271), .ZN(n1178) );
NAND2_X1 U1106 ( .A1(n1360), .A2(n1180), .ZN(n1271) );
NAND2_X1 U1107 ( .A1(n1441), .A2(n1210), .ZN(n1180) );
NAND2_X1 U1108 ( .A1(n1207), .A2(n1209), .ZN(n1210) );
OR2_X1 U1109 ( .A1(n1209), .A2(n1207), .ZN(n1441) );
AND2_X1 U1110 ( .A1(n1442), .A2(n1267), .ZN(n1207) );
XOR2_X1 U1111 ( .A(n1304), .B(n1443), .Z(n1442) );
XOR2_X1 U1112 ( .A(KEYINPUT61), .B(KEYINPUT31), .Z(n1443) );
XOR2_X1 U1113 ( .A(n1444), .B(n1445), .Z(n1304) );
XOR2_X1 U1114 ( .A(n1290), .B(n1446), .Z(n1445) );
XOR2_X1 U1115 ( .A(G125), .B(n1447), .Z(n1446) );
AND2_X1 U1116 ( .A1(n1228), .A2(G224), .ZN(n1447) );
XOR2_X1 U1117 ( .A(G146), .B(n1448), .Z(n1290) );
XNOR2_X1 U1118 ( .A(n1247), .B(n1248), .ZN(n1444) );
XOR2_X1 U1119 ( .A(G122), .B(G110), .Z(n1248) );
XNOR2_X1 U1120 ( .A(n1449), .B(n1450), .ZN(n1247) );
XOR2_X1 U1121 ( .A(n1451), .B(n1417), .Z(n1450) );
XOR2_X1 U1122 ( .A(G116), .B(G119), .Z(n1417) );
NOR2_X1 U1123 ( .A1(n1452), .A2(n1453), .ZN(n1451) );
XOR2_X1 U1124 ( .A(KEYINPUT18), .B(n1454), .Z(n1453) );
NOR2_X1 U1125 ( .A1(n1455), .A2(n1456), .ZN(n1454) );
XOR2_X1 U1126 ( .A(KEYINPUT27), .B(G107), .Z(n1456) );
NOR2_X1 U1127 ( .A1(G104), .A2(n1457), .ZN(n1452) );
XOR2_X1 U1128 ( .A(KEYINPUT41), .B(G107), .Z(n1457) );
XOR2_X1 U1129 ( .A(n1458), .B(G101), .Z(n1449) );
NAND2_X1 U1130 ( .A1(KEYINPUT54), .A2(n1388), .ZN(n1458) );
INV_X1 U1131 ( .A(G113), .ZN(n1388) );
NAND2_X1 U1132 ( .A1(G210), .A2(n1459), .ZN(n1209) );
XNOR2_X1 U1133 ( .A(n1179), .B(KEYINPUT16), .ZN(n1360) );
NAND2_X1 U1134 ( .A1(G214), .A2(n1459), .ZN(n1179) );
NAND2_X1 U1135 ( .A1(n1267), .A2(n1460), .ZN(n1459) );
INV_X1 U1136 ( .A(G237), .ZN(n1460) );
NAND2_X1 U1137 ( .A1(n1394), .A2(n1385), .ZN(n1169) );
INV_X1 U1138 ( .A(n1373), .ZN(n1385) );
NAND3_X1 U1139 ( .A1(n1461), .A2(n1462), .A3(n1197), .ZN(n1373) );
NAND2_X1 U1140 ( .A1(n1263), .A2(n1463), .ZN(n1197) );
OR2_X1 U1141 ( .A1(n1196), .A2(KEYINPUT48), .ZN(n1462) );
OR2_X1 U1142 ( .A1(n1463), .A2(n1263), .ZN(n1196) );
INV_X1 U1143 ( .A(G475), .ZN(n1463) );
NAND2_X1 U1144 ( .A1(KEYINPUT48), .A2(n1263), .ZN(n1461) );
AND2_X1 U1145 ( .A1(n1266), .A2(n1267), .ZN(n1263) );
INV_X1 U1146 ( .A(G902), .ZN(n1267) );
NAND2_X1 U1147 ( .A1(n1464), .A2(n1465), .ZN(n1266) );
NAND4_X1 U1148 ( .A1(KEYINPUT23), .A2(n1466), .A3(n1467), .A4(n1468), .ZN(n1465) );
NAND2_X1 U1149 ( .A1(n1469), .A2(n1455), .ZN(n1468) );
NAND2_X1 U1150 ( .A1(n1470), .A2(G104), .ZN(n1467) );
NAND3_X1 U1151 ( .A1(n1471), .A2(n1472), .A3(n1473), .ZN(n1464) );
NAND2_X1 U1152 ( .A1(KEYINPUT23), .A2(n1466), .ZN(n1473) );
XOR2_X1 U1153 ( .A(G122), .B(G113), .Z(n1466) );
NAND2_X1 U1154 ( .A1(n1469), .A2(G104), .ZN(n1472) );
NAND2_X1 U1155 ( .A1(n1470), .A2(n1455), .ZN(n1471) );
INV_X1 U1156 ( .A(G104), .ZN(n1455) );
XNOR2_X1 U1157 ( .A(n1474), .B(n1469), .ZN(n1470) );
XOR2_X1 U1158 ( .A(n1475), .B(n1476), .Z(n1469) );
XOR2_X1 U1159 ( .A(G125), .B(n1477), .Z(n1476) );
XOR2_X1 U1160 ( .A(KEYINPUT2), .B(G146), .Z(n1477) );
XNOR2_X1 U1161 ( .A(n1478), .B(n1479), .ZN(n1475) );
NAND2_X1 U1162 ( .A1(KEYINPUT25), .A2(n1480), .ZN(n1479) );
INV_X1 U1163 ( .A(G140), .ZN(n1480) );
NAND2_X1 U1164 ( .A1(n1481), .A2(KEYINPUT36), .ZN(n1478) );
XOR2_X1 U1165 ( .A(n1482), .B(n1483), .Z(n1481) );
XOR2_X1 U1166 ( .A(G143), .B(G131), .Z(n1483) );
NAND2_X1 U1167 ( .A1(n1420), .A2(G214), .ZN(n1482) );
NOR2_X1 U1168 ( .A1(G953), .A2(G237), .ZN(n1420) );
XNOR2_X1 U1169 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n1474) );
XOR2_X1 U1170 ( .A(n1372), .B(KEYINPUT5), .Z(n1394) );
XNOR2_X1 U1171 ( .A(n1205), .B(n1484), .ZN(n1372) );
NOR2_X1 U1172 ( .A1(G478), .A2(KEYINPUT62), .ZN(n1484) );
NOR2_X1 U1173 ( .A1(n1259), .A2(G902), .ZN(n1205) );
XOR2_X1 U1174 ( .A(n1485), .B(n1486), .Z(n1259) );
XOR2_X1 U1175 ( .A(n1487), .B(n1488), .Z(n1486) );
NAND3_X1 U1176 ( .A1(G234), .A2(n1228), .A3(G217), .ZN(n1488) );
INV_X1 U1177 ( .A(G953), .ZN(n1228) );
NAND2_X1 U1178 ( .A1(n1489), .A2(n1490), .ZN(n1487) );
NAND2_X1 U1179 ( .A1(G107), .A2(n1491), .ZN(n1490) );
NAND2_X1 U1180 ( .A1(KEYINPUT34), .A2(n1492), .ZN(n1491) );
NAND2_X1 U1181 ( .A1(KEYINPUT26), .A2(n1493), .ZN(n1492) );
NAND2_X1 U1182 ( .A1(n1494), .A2(n1495), .ZN(n1489) );
NAND2_X1 U1183 ( .A1(KEYINPUT26), .A2(n1496), .ZN(n1495) );
NAND2_X1 U1184 ( .A1(KEYINPUT34), .A2(n1497), .ZN(n1496) );
INV_X1 U1185 ( .A(G107), .ZN(n1497) );
INV_X1 U1186 ( .A(n1493), .ZN(n1494) );
XOR2_X1 U1187 ( .A(n1498), .B(G122), .Z(n1493) );
INV_X1 U1188 ( .A(G116), .ZN(n1498) );
NAND2_X1 U1189 ( .A1(n1499), .A2(KEYINPUT63), .ZN(n1485) );
XOR2_X1 U1190 ( .A(n1500), .B(n1448), .Z(n1499) );
XOR2_X1 U1191 ( .A(G128), .B(G143), .Z(n1448) );
XOR2_X1 U1192 ( .A(n1501), .B(KEYINPUT58), .Z(n1500) );
INV_X1 U1193 ( .A(G134), .ZN(n1501) );
endmodule


