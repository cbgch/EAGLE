//Key = 0000000001011110010110011001001011100010111000011111011110010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297;

XNOR2_X1 U696 ( .A(n981), .B(n982), .ZN(G9) );
NOR2_X1 U697 ( .A1(n983), .A2(n984), .ZN(G75) );
NOR3_X1 U698 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n984) );
NOR2_X1 U699 ( .A1(n988), .A2(n989), .ZN(n986) );
INV_X1 U700 ( .A(n990), .ZN(n989) );
NOR2_X1 U701 ( .A1(n991), .A2(n992), .ZN(n988) );
NOR2_X1 U702 ( .A1(KEYINPUT33), .A2(n993), .ZN(n992) );
NOR4_X1 U703 ( .A1(n994), .A2(n995), .A3(n996), .A4(n997), .ZN(n993) );
OR2_X1 U704 ( .A1(n998), .A2(n999), .ZN(n995) );
NOR3_X1 U705 ( .A1(n994), .A2(n1000), .A3(n1001), .ZN(n991) );
NOR2_X1 U706 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
AND2_X1 U707 ( .A1(KEYINPUT20), .A2(n1004), .ZN(n1002) );
NOR2_X1 U708 ( .A1(n999), .A2(n1005), .ZN(n1000) );
NOR2_X1 U709 ( .A1(n1006), .A2(n998), .ZN(n1005) );
NOR2_X1 U710 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NOR2_X1 U711 ( .A1(n1009), .A2(n997), .ZN(n1008) );
NOR2_X1 U712 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
AND2_X1 U713 ( .A1(n1012), .A2(KEYINPUT33), .ZN(n1010) );
NOR2_X1 U714 ( .A1(n1013), .A2(n1014), .ZN(n1007) );
NOR2_X1 U715 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NAND3_X1 U716 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n985) );
NAND4_X1 U717 ( .A1(n1004), .A2(n1003), .A3(n1020), .A4(n1021), .ZN(n1019) );
NAND2_X1 U718 ( .A1(n1022), .A2(n994), .ZN(n1021) );
XNOR2_X1 U719 ( .A(n990), .B(KEYINPUT29), .ZN(n1022) );
NAND2_X1 U720 ( .A1(n1023), .A2(n1024), .ZN(n1020) );
NAND2_X1 U721 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U722 ( .A1(KEYINPUT20), .A2(n990), .ZN(n1026) );
NAND2_X1 U723 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR3_X1 U724 ( .A1(n998), .A2(n1014), .A3(n997), .ZN(n1004) );
INV_X1 U725 ( .A(n1029), .ZN(n997) );
NOR3_X1 U726 ( .A1(n1030), .A2(G953), .A3(G952), .ZN(n983) );
INV_X1 U727 ( .A(n1017), .ZN(n1030) );
NAND4_X1 U728 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1017) );
NOR4_X1 U729 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1034) );
XNOR2_X1 U730 ( .A(n1028), .B(KEYINPUT53), .ZN(n1036) );
XOR2_X1 U731 ( .A(n1039), .B(KEYINPUT51), .Z(n1035) );
NAND2_X1 U732 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
XNOR2_X1 U733 ( .A(KEYINPUT31), .B(n1042), .ZN(n1040) );
NOR3_X1 U734 ( .A1(n999), .A2(n1043), .A3(n1027), .ZN(n1033) );
INV_X1 U735 ( .A(n1003), .ZN(n999) );
XNOR2_X1 U736 ( .A(n1044), .B(n1045), .ZN(n1032) );
NOR2_X1 U737 ( .A1(n1046), .A2(KEYINPUT8), .ZN(n1045) );
XOR2_X1 U738 ( .A(n1047), .B(n1048), .Z(n1031) );
XNOR2_X1 U739 ( .A(KEYINPUT45), .B(KEYINPUT32), .ZN(n1048) );
NAND2_X1 U740 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
OR2_X1 U741 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U742 ( .A(n1053), .B(n1054), .Z(G72) );
XOR2_X1 U743 ( .A(n1055), .B(n1056), .Z(n1054) );
NOR2_X1 U744 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
XNOR2_X1 U745 ( .A(G953), .B(KEYINPUT14), .ZN(n1058) );
NAND3_X1 U746 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1055) );
NAND2_X1 U747 ( .A1(G953), .A2(n1062), .ZN(n1061) );
NAND2_X1 U748 ( .A1(n1063), .A2(n1064), .ZN(n1060) );
XNOR2_X1 U749 ( .A(G140), .B(n1065), .ZN(n1064) );
XOR2_X1 U750 ( .A(n1066), .B(KEYINPUT39), .Z(n1063) );
NAND2_X1 U751 ( .A1(n1067), .A2(n1068), .ZN(n1059) );
XOR2_X1 U752 ( .A(n1066), .B(KEYINPUT9), .Z(n1068) );
XNOR2_X1 U753 ( .A(n1069), .B(n1070), .ZN(n1066) );
XNOR2_X1 U754 ( .A(G125), .B(G140), .ZN(n1067) );
NAND2_X1 U755 ( .A1(G953), .A2(n1071), .ZN(n1053) );
NAND2_X1 U756 ( .A1(G900), .A2(G227), .ZN(n1071) );
XOR2_X1 U757 ( .A(n1072), .B(n1073), .Z(G69) );
NOR2_X1 U758 ( .A1(n1074), .A2(n1018), .ZN(n1073) );
NOR2_X1 U759 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U760 ( .A1(KEYINPUT37), .A2(n1077), .ZN(n1072) );
XOR2_X1 U761 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U762 ( .A1(G953), .A2(n1080), .ZN(n1079) );
NAND2_X1 U763 ( .A1(n1081), .A2(n1082), .ZN(n1078) );
NAND2_X1 U764 ( .A1(G953), .A2(n1076), .ZN(n1082) );
XOR2_X1 U765 ( .A(n1083), .B(KEYINPUT56), .Z(n1081) );
NAND2_X1 U766 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U767 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XNOR2_X1 U768 ( .A(n1088), .B(KEYINPUT35), .ZN(n1087) );
XNOR2_X1 U769 ( .A(n1089), .B(KEYINPUT58), .ZN(n1086) );
XOR2_X1 U770 ( .A(n1090), .B(KEYINPUT25), .Z(n1084) );
NAND2_X1 U771 ( .A1(n1088), .A2(n1089), .ZN(n1090) );
AND2_X1 U772 ( .A1(n1091), .A2(n1092), .ZN(n1088) );
NAND2_X1 U773 ( .A1(KEYINPUT55), .A2(n1093), .ZN(n1092) );
OR3_X1 U774 ( .A1(n1094), .A2(n1095), .A3(KEYINPUT55), .ZN(n1091) );
NOR3_X1 U775 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(G66) );
NOR3_X1 U776 ( .A1(n1099), .A2(G953), .A3(G952), .ZN(n1098) );
AND2_X1 U777 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
INV_X1 U778 ( .A(KEYINPUT57), .ZN(n1099) );
XOR2_X1 U779 ( .A(n1101), .B(n1102), .Z(n1096) );
NOR2_X1 U780 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U781 ( .A1(n1100), .A2(n1105), .ZN(G63) );
XNOR2_X1 U782 ( .A(n1106), .B(n1107), .ZN(n1105) );
NOR2_X1 U783 ( .A1(n1108), .A2(n1104), .ZN(n1107) );
NOR2_X1 U784 ( .A1(n1100), .A2(n1109), .ZN(G60) );
XOR2_X1 U785 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U786 ( .A1(n1042), .A2(n1104), .ZN(n1111) );
INV_X1 U787 ( .A(G475), .ZN(n1042) );
NAND2_X1 U788 ( .A1(KEYINPUT63), .A2(n1112), .ZN(n1110) );
XOR2_X1 U789 ( .A(G104), .B(n1113), .Z(G6) );
NOR2_X1 U790 ( .A1(n1100), .A2(n1114), .ZN(G57) );
XOR2_X1 U791 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U792 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U793 ( .A1(G101), .A2(KEYINPUT28), .ZN(n1118) );
NOR2_X1 U794 ( .A1(n1104), .A2(n1119), .ZN(n1117) );
XOR2_X1 U795 ( .A(KEYINPUT12), .B(G472), .Z(n1119) );
XOR2_X1 U796 ( .A(n1120), .B(n1121), .Z(n1115) );
NOR2_X1 U797 ( .A1(n1100), .A2(n1122), .ZN(G54) );
XOR2_X1 U798 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U799 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR3_X1 U800 ( .A1(n1104), .A2(KEYINPUT61), .A3(n1044), .ZN(n1125) );
NAND2_X1 U801 ( .A1(G902), .A2(n987), .ZN(n1104) );
NOR2_X1 U802 ( .A1(n1100), .A2(n1127), .ZN(G51) );
XNOR2_X1 U803 ( .A(n1128), .B(n1129), .ZN(n1127) );
XOR2_X1 U804 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U805 ( .A1(KEYINPUT17), .A2(n1132), .ZN(n1131) );
NAND3_X1 U806 ( .A1(n1133), .A2(G902), .A3(n1134), .ZN(n1130) );
XOR2_X1 U807 ( .A(n987), .B(KEYINPUT15), .Z(n1134) );
NAND2_X1 U808 ( .A1(n1057), .A2(n1080), .ZN(n987) );
AND4_X1 U809 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1080) );
NOR4_X1 U810 ( .A1(n1139), .A2(n982), .A3(n1140), .A4(n1141), .ZN(n1138) );
INV_X1 U811 ( .A(n1142), .ZN(n1141) );
AND3_X1 U812 ( .A1(n1015), .A2(n1143), .A3(n1144), .ZN(n982) );
NOR2_X1 U813 ( .A1(n1113), .A2(n1145), .ZN(n1137) );
AND3_X1 U814 ( .A1(n1146), .A2(n1147), .A3(n1029), .ZN(n1145) );
AND3_X1 U815 ( .A1(n1144), .A2(n1143), .A3(n1016), .ZN(n1113) );
AND4_X1 U816 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1057) );
NOR4_X1 U817 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1151) );
NOR2_X1 U818 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XNOR2_X1 U819 ( .A(n1016), .B(KEYINPUT3), .ZN(n1156) );
INV_X1 U820 ( .A(n1158), .ZN(n1154) );
AND2_X1 U821 ( .A1(n1159), .A2(n1160), .ZN(n1150) );
NOR2_X1 U822 ( .A1(n1018), .A2(G952), .ZN(n1100) );
XNOR2_X1 U823 ( .A(G146), .B(n1158), .ZN(G48) );
NAND3_X1 U824 ( .A1(n1016), .A2(n1147), .A3(n1161), .ZN(n1158) );
XNOR2_X1 U825 ( .A(n1153), .B(n1162), .ZN(G45) );
NAND2_X1 U826 ( .A1(KEYINPUT11), .A2(n1163), .ZN(n1162) );
XNOR2_X1 U827 ( .A(KEYINPUT26), .B(n1164), .ZN(n1163) );
AND4_X1 U828 ( .A1(n1161), .A2(n1012), .A3(n1038), .A4(n1165), .ZN(n1153) );
XOR2_X1 U829 ( .A(G140), .B(n1166), .Z(G42) );
NOR2_X1 U830 ( .A1(KEYINPUT2), .A2(n1159), .ZN(n1166) );
NAND3_X1 U831 ( .A1(n1011), .A2(n1167), .A3(n1016), .ZN(n1159) );
XOR2_X1 U832 ( .A(G137), .B(n1152), .Z(G39) );
AND3_X1 U833 ( .A1(n1167), .A2(n1147), .A3(n1029), .ZN(n1152) );
XNOR2_X1 U834 ( .A(G134), .B(n1148), .ZN(G36) );
NAND2_X1 U835 ( .A1(n1168), .A2(n1015), .ZN(n1148) );
XNOR2_X1 U836 ( .A(G131), .B(n1169), .ZN(G33) );
NAND2_X1 U837 ( .A1(n1168), .A2(n1016), .ZN(n1169) );
INV_X1 U838 ( .A(n1157), .ZN(n1168) );
NAND2_X1 U839 ( .A1(n1012), .A2(n1167), .ZN(n1157) );
AND4_X1 U840 ( .A1(n990), .A2(n994), .A3(n1170), .A4(n1003), .ZN(n1167) );
NOR2_X1 U841 ( .A1(n1028), .A2(n1027), .ZN(n990) );
INV_X1 U842 ( .A(n1171), .ZN(n1027) );
NAND2_X1 U843 ( .A1(n1172), .A2(n1173), .ZN(G30) );
NAND2_X1 U844 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XNOR2_X1 U845 ( .A(KEYINPUT36), .B(n1149), .ZN(n1174) );
NAND2_X1 U846 ( .A1(n1176), .A2(G128), .ZN(n1172) );
XNOR2_X1 U847 ( .A(KEYINPUT48), .B(n1149), .ZN(n1176) );
NAND3_X1 U848 ( .A1(n1015), .A2(n1147), .A3(n1161), .ZN(n1149) );
AND2_X1 U849 ( .A1(n1177), .A2(n994), .ZN(n1161) );
XNOR2_X1 U850 ( .A(G101), .B(n1135), .ZN(G3) );
NAND3_X1 U851 ( .A1(n1012), .A2(n1144), .A3(n1029), .ZN(n1135) );
XNOR2_X1 U852 ( .A(G125), .B(n1160), .ZN(G27) );
NAND4_X1 U853 ( .A1(n1023), .A2(n1177), .A3(n1016), .A4(n1011), .ZN(n1160) );
AND4_X1 U854 ( .A1(n1028), .A2(n1170), .A3(n1003), .A4(n1171), .ZN(n1177) );
NAND2_X1 U855 ( .A1(n1178), .A2(n1179), .ZN(n1170) );
NAND4_X1 U856 ( .A1(G953), .A2(G902), .A3(n1062), .A4(n1180), .ZN(n1179) );
XOR2_X1 U857 ( .A(KEYINPUT23), .B(G900), .Z(n1062) );
XOR2_X1 U858 ( .A(n998), .B(KEYINPUT16), .Z(n1178) );
XNOR2_X1 U859 ( .A(G122), .B(n1136), .ZN(G24) );
NAND4_X1 U860 ( .A1(n1146), .A2(n1143), .A3(n1038), .A4(n1165), .ZN(n1136) );
INV_X1 U861 ( .A(n1014), .ZN(n1143) );
NAND2_X1 U862 ( .A1(n1181), .A2(n1182), .ZN(n1014) );
XNOR2_X1 U863 ( .A(G119), .B(n1183), .ZN(G21) );
NAND4_X1 U864 ( .A1(KEYINPUT42), .A2(n1146), .A3(n1029), .A4(n1147), .ZN(n1183) );
NAND2_X1 U865 ( .A1(n1184), .A2(n1185), .ZN(n1147) );
OR3_X1 U866 ( .A1(n1182), .A2(n1181), .A3(KEYINPUT1), .ZN(n1185) );
INV_X1 U867 ( .A(n1037), .ZN(n1181) );
NAND2_X1 U868 ( .A1(KEYINPUT1), .A2(n1012), .ZN(n1184) );
XOR2_X1 U869 ( .A(G116), .B(n1186), .Z(G18) );
NOR2_X1 U870 ( .A1(KEYINPUT18), .A2(n1142), .ZN(n1186) );
NAND3_X1 U871 ( .A1(n1012), .A2(n1015), .A3(n1146), .ZN(n1142) );
NOR2_X1 U872 ( .A1(n1165), .A2(n1187), .ZN(n1015) );
INV_X1 U873 ( .A(n1038), .ZN(n1187) );
XOR2_X1 U874 ( .A(G113), .B(n1139), .Z(G15) );
AND3_X1 U875 ( .A1(n1012), .A2(n1016), .A3(n1146), .ZN(n1139) );
AND3_X1 U876 ( .A1(n1188), .A2(n1003), .A3(n1023), .ZN(n1146) );
NOR2_X1 U877 ( .A1(n1038), .A2(n1189), .ZN(n1016) );
INV_X1 U878 ( .A(n996), .ZN(n1012) );
NAND2_X1 U879 ( .A1(n1037), .A2(n1182), .ZN(n996) );
NAND2_X1 U880 ( .A1(n1190), .A2(n1191), .ZN(G12) );
NAND2_X1 U881 ( .A1(n1140), .A2(n1192), .ZN(n1191) );
INV_X1 U882 ( .A(n1193), .ZN(n1140) );
XOR2_X1 U883 ( .A(n1194), .B(KEYINPUT46), .Z(n1190) );
NAND2_X1 U884 ( .A1(G110), .A2(n1193), .ZN(n1194) );
NAND3_X1 U885 ( .A1(n1011), .A2(n1144), .A3(n1029), .ZN(n1193) );
NOR2_X1 U886 ( .A1(n1038), .A2(n1165), .ZN(n1029) );
INV_X1 U887 ( .A(n1189), .ZN(n1165) );
NOR2_X1 U888 ( .A1(n1195), .A2(n1043), .ZN(n1189) );
NOR2_X1 U889 ( .A1(n1041), .A2(G475), .ZN(n1043) );
AND2_X1 U890 ( .A1(G475), .A2(n1041), .ZN(n1195) );
NAND2_X1 U891 ( .A1(n1112), .A2(n1196), .ZN(n1041) );
XNOR2_X1 U892 ( .A(n1197), .B(n1198), .ZN(n1112) );
XOR2_X1 U893 ( .A(G104), .B(n1199), .Z(n1198) );
NOR2_X1 U894 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U895 ( .A(n1202), .B(KEYINPUT49), .Z(n1201) );
NAND2_X1 U896 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NOR2_X1 U897 ( .A1(n1203), .A2(n1204), .ZN(n1200) );
XNOR2_X1 U898 ( .A(n1205), .B(n1206), .ZN(n1204) );
XNOR2_X1 U899 ( .A(n1164), .B(G131), .ZN(n1206) );
NAND3_X1 U900 ( .A1(G214), .A2(n1018), .A3(n1207), .ZN(n1205) );
XOR2_X1 U901 ( .A(n1208), .B(n1209), .Z(n1203) );
XNOR2_X1 U902 ( .A(n1210), .B(G140), .ZN(n1209) );
NAND2_X1 U903 ( .A1(KEYINPUT19), .A2(n1211), .ZN(n1208) );
XNOR2_X1 U904 ( .A(KEYINPUT59), .B(n1065), .ZN(n1211) );
XNOR2_X1 U905 ( .A(G113), .B(G122), .ZN(n1197) );
XOR2_X1 U906 ( .A(n1212), .B(n1108), .Z(n1038) );
INV_X1 U907 ( .A(G478), .ZN(n1108) );
NAND2_X1 U908 ( .A1(n1106), .A2(n1196), .ZN(n1212) );
XNOR2_X1 U909 ( .A(n1213), .B(n1214), .ZN(n1106) );
NOR2_X1 U910 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
INV_X1 U911 ( .A(G217), .ZN(n1216) );
NAND4_X1 U912 ( .A1(KEYINPUT47), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1213) );
NAND3_X1 U913 ( .A1(n1220), .A2(n1221), .A3(KEYINPUT34), .ZN(n1219) );
NAND2_X1 U914 ( .A1(n1222), .A2(n1223), .ZN(n1218) );
INV_X1 U915 ( .A(KEYINPUT34), .ZN(n1223) );
OR2_X1 U916 ( .A1(n1221), .A2(n1220), .ZN(n1217) );
NOR2_X1 U917 ( .A1(KEYINPUT5), .A2(n1222), .ZN(n1220) );
XOR2_X1 U918 ( .A(n1224), .B(n1225), .Z(n1222) );
XNOR2_X1 U919 ( .A(n1070), .B(G128), .ZN(n1225) );
XNOR2_X1 U920 ( .A(n1226), .B(n1164), .ZN(n1224) );
INV_X1 U921 ( .A(G143), .ZN(n1164) );
XNOR2_X1 U922 ( .A(KEYINPUT7), .B(KEYINPUT24), .ZN(n1226) );
XOR2_X1 U923 ( .A(n1227), .B(n1228), .Z(n1221) );
XNOR2_X1 U924 ( .A(KEYINPUT0), .B(n1229), .ZN(n1228) );
INV_X1 U925 ( .A(G122), .ZN(n1229) );
XNOR2_X1 U926 ( .A(G116), .B(G107), .ZN(n1227) );
AND3_X1 U927 ( .A1(n994), .A2(n1003), .A3(n1188), .ZN(n1144) );
AND3_X1 U928 ( .A1(n1230), .A2(n1171), .A3(n1028), .ZN(n1188) );
XNOR2_X1 U929 ( .A(n1231), .B(n1133), .ZN(n1028) );
AND2_X1 U930 ( .A1(G210), .A2(n1232), .ZN(n1133) );
NAND2_X1 U931 ( .A1(n1233), .A2(n1196), .ZN(n1231) );
XNOR2_X1 U932 ( .A(n1234), .B(n1132), .ZN(n1233) );
XNOR2_X1 U933 ( .A(n1235), .B(n1093), .ZN(n1132) );
XOR2_X1 U934 ( .A(n1095), .B(n1094), .Z(n1093) );
NAND2_X1 U935 ( .A1(n1236), .A2(n1237), .ZN(n1095) );
NAND2_X1 U936 ( .A1(G101), .A2(n1238), .ZN(n1237) );
NAND2_X1 U937 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
XNOR2_X1 U938 ( .A(n1241), .B(KEYINPUT52), .ZN(n1239) );
NAND2_X1 U939 ( .A1(n1242), .A2(n1243), .ZN(n1236) );
NAND2_X1 U940 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
NAND3_X1 U941 ( .A1(n1240), .A2(n1246), .A3(n1247), .ZN(n1245) );
INV_X1 U942 ( .A(KEYINPUT52), .ZN(n1247) );
NAND2_X1 U943 ( .A1(n1241), .A2(KEYINPUT52), .ZN(n1244) );
NAND2_X1 U944 ( .A1(KEYINPUT41), .A2(n1089), .ZN(n1235) );
XOR2_X1 U945 ( .A(G110), .B(G122), .Z(n1089) );
INV_X1 U946 ( .A(n1128), .ZN(n1234) );
XNOR2_X1 U947 ( .A(n1248), .B(n1249), .ZN(n1128) );
XNOR2_X1 U948 ( .A(n1065), .B(n1250), .ZN(n1249) );
NOR2_X1 U949 ( .A1(G953), .A2(n1075), .ZN(n1250) );
INV_X1 U950 ( .A(G224), .ZN(n1075) );
INV_X1 U951 ( .A(G125), .ZN(n1065) );
NAND2_X1 U952 ( .A1(G214), .A2(n1232), .ZN(n1171) );
NAND2_X1 U953 ( .A1(n1251), .A2(n1252), .ZN(n1232) );
XNOR2_X1 U954 ( .A(KEYINPUT30), .B(n1196), .ZN(n1251) );
NAND2_X1 U955 ( .A1(n998), .A2(n1253), .ZN(n1230) );
NAND4_X1 U956 ( .A1(G953), .A2(G902), .A3(n1180), .A4(n1076), .ZN(n1253) );
INV_X1 U957 ( .A(G898), .ZN(n1076) );
NAND3_X1 U958 ( .A1(n1180), .A2(n1018), .A3(G952), .ZN(n998) );
NAND2_X1 U959 ( .A1(G237), .A2(G234), .ZN(n1180) );
NAND2_X1 U960 ( .A1(G221), .A2(n1254), .ZN(n1003) );
INV_X1 U961 ( .A(n1023), .ZN(n994) );
XOR2_X1 U962 ( .A(n1046), .B(n1044), .Z(n1023) );
INV_X1 U963 ( .A(G469), .ZN(n1044) );
AND2_X1 U964 ( .A1(n1255), .A2(n1196), .ZN(n1046) );
XOR2_X1 U965 ( .A(n1256), .B(n1126), .Z(n1255) );
XNOR2_X1 U966 ( .A(n1257), .B(n1258), .ZN(n1126) );
NOR2_X1 U967 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
XNOR2_X1 U968 ( .A(KEYINPUT62), .B(n1018), .ZN(n1260) );
INV_X1 U969 ( .A(G227), .ZN(n1259) );
XNOR2_X1 U970 ( .A(G110), .B(G140), .ZN(n1257) );
NOR2_X1 U971 ( .A1(KEYINPUT10), .A2(n1123), .ZN(n1256) );
XOR2_X1 U972 ( .A(n1261), .B(n1262), .Z(n1123) );
XOR2_X1 U973 ( .A(n1263), .B(n1069), .Z(n1262) );
XNOR2_X1 U974 ( .A(n1264), .B(n1265), .ZN(n1069) );
NOR2_X1 U975 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XOR2_X1 U976 ( .A(n1268), .B(KEYINPUT50), .Z(n1267) );
NAND2_X1 U977 ( .A1(n1269), .A2(n1175), .ZN(n1268) );
XOR2_X1 U978 ( .A(KEYINPUT44), .B(n1270), .Z(n1269) );
NOR2_X1 U979 ( .A1(n1175), .A2(n1270), .ZN(n1266) );
XOR2_X1 U980 ( .A(n1271), .B(KEYINPUT27), .Z(n1270) );
INV_X1 U981 ( .A(G128), .ZN(n1175) );
XNOR2_X1 U982 ( .A(n1272), .B(n1243), .ZN(n1261) );
INV_X1 U983 ( .A(G101), .ZN(n1243) );
NAND2_X1 U984 ( .A1(n1246), .A2(n1240), .ZN(n1272) );
NAND2_X1 U985 ( .A1(n1273), .A2(n981), .ZN(n1240) );
INV_X1 U986 ( .A(n1241), .ZN(n1246) );
NOR2_X1 U987 ( .A1(n981), .A2(n1273), .ZN(n1241) );
XNOR2_X1 U988 ( .A(G104), .B(KEYINPUT38), .ZN(n1273) );
INV_X1 U989 ( .A(G107), .ZN(n981) );
NOR2_X1 U990 ( .A1(n1182), .A2(n1037), .ZN(n1011) );
XNOR2_X1 U991 ( .A(n1274), .B(G472), .ZN(n1037) );
NAND2_X1 U992 ( .A1(n1275), .A2(n1196), .ZN(n1274) );
XOR2_X1 U993 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U994 ( .A(n1120), .B(n1278), .Z(n1277) );
NOR2_X1 U995 ( .A1(KEYINPUT22), .A2(n1121), .ZN(n1278) );
XNOR2_X1 U996 ( .A(n1263), .B(n1264), .ZN(n1121) );
XOR2_X1 U997 ( .A(G131), .B(G137), .Z(n1264) );
NAND2_X1 U998 ( .A1(KEYINPUT54), .A2(n1070), .ZN(n1263) );
INV_X1 U999 ( .A(G134), .ZN(n1070) );
XOR2_X1 U1000 ( .A(n1279), .B(n1280), .Z(n1120) );
XOR2_X1 U1001 ( .A(KEYINPUT43), .B(n1281), .Z(n1280) );
AND3_X1 U1002 ( .A1(n1207), .A2(n1018), .A3(G210), .ZN(n1281) );
XOR2_X1 U1003 ( .A(n1252), .B(KEYINPUT60), .Z(n1207) );
INV_X1 U1004 ( .A(G237), .ZN(n1252) );
XNOR2_X1 U1005 ( .A(n1248), .B(n1094), .ZN(n1279) );
XNOR2_X1 U1006 ( .A(G113), .B(n1282), .ZN(n1094) );
XOR2_X1 U1007 ( .A(G119), .B(G116), .Z(n1282) );
XNOR2_X1 U1008 ( .A(G128), .B(n1271), .ZN(n1248) );
XNOR2_X1 U1009 ( .A(G143), .B(n1210), .ZN(n1271) );
XNOR2_X1 U1010 ( .A(G101), .B(KEYINPUT6), .ZN(n1276) );
NAND3_X1 U1011 ( .A1(n1283), .A2(n1284), .A3(n1049), .ZN(n1182) );
NAND2_X1 U1012 ( .A1(n1052), .A2(n1051), .ZN(n1049) );
OR3_X1 U1013 ( .A1(n1051), .A2(n1052), .A3(KEYINPUT21), .ZN(n1284) );
NOR2_X1 U1014 ( .A1(n1101), .A2(G902), .ZN(n1051) );
XOR2_X1 U1015 ( .A(n1285), .B(n1286), .Z(n1101) );
NOR2_X1 U1016 ( .A1(n1287), .A2(n1215), .ZN(n1286) );
NAND2_X1 U1017 ( .A1(G234), .A2(n1018), .ZN(n1215) );
INV_X1 U1018 ( .A(G953), .ZN(n1018) );
INV_X1 U1019 ( .A(G221), .ZN(n1287) );
XOR2_X1 U1020 ( .A(n1288), .B(G137), .Z(n1285) );
NAND2_X1 U1021 ( .A1(KEYINPUT40), .A2(n1289), .ZN(n1288) );
XOR2_X1 U1022 ( .A(n1290), .B(n1291), .Z(n1289) );
XNOR2_X1 U1023 ( .A(n1292), .B(n1192), .ZN(n1291) );
INV_X1 U1024 ( .A(G110), .ZN(n1192) );
NAND2_X1 U1025 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
NAND2_X1 U1026 ( .A1(n1295), .A2(n1210), .ZN(n1294) );
XOR2_X1 U1027 ( .A(KEYINPUT13), .B(n1296), .Z(n1293) );
NOR2_X1 U1028 ( .A1(n1210), .A2(n1295), .ZN(n1296) );
XOR2_X1 U1029 ( .A(G140), .B(n1297), .Z(n1295) );
NOR2_X1 U1030 ( .A1(G125), .A2(KEYINPUT4), .ZN(n1297) );
INV_X1 U1031 ( .A(G146), .ZN(n1210) );
XNOR2_X1 U1032 ( .A(G119), .B(G128), .ZN(n1290) );
NAND2_X1 U1033 ( .A1(KEYINPUT21), .A2(n1052), .ZN(n1283) );
INV_X1 U1034 ( .A(n1103), .ZN(n1052) );
NAND2_X1 U1035 ( .A1(G217), .A2(n1254), .ZN(n1103) );
NAND2_X1 U1036 ( .A1(G234), .A2(n1196), .ZN(n1254) );
INV_X1 U1037 ( .A(G902), .ZN(n1196) );
endmodule


