//Key = 0110010110100111010001111100010100100111111101111011111000001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330;

XNOR2_X1 U719 ( .A(G107), .B(n997), .ZN(G9) );
NAND3_X1 U720 ( .A1(n998), .A2(n999), .A3(KEYINPUT23), .ZN(n997) );
NOR2_X1 U721 ( .A1(n1000), .A2(n1001), .ZN(G75) );
XOR2_X1 U722 ( .A(n1002), .B(KEYINPUT45), .Z(n1001) );
NAND3_X1 U723 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1002) );
NOR3_X1 U724 ( .A1(n1006), .A2(n1003), .A3(n1007), .ZN(n1000) );
NAND3_X1 U725 ( .A1(n1005), .A2(n1004), .A3(n1008), .ZN(n1006) );
NAND2_X1 U726 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND2_X1 U727 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND3_X1 U728 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
OR2_X1 U729 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NAND2_X1 U730 ( .A1(n1018), .A2(n1019), .ZN(n1011) );
NAND2_X1 U731 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U732 ( .A1(n1015), .A2(n1022), .ZN(n1021) );
NAND2_X1 U733 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U734 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U735 ( .A1(n1013), .A2(n1027), .ZN(n1020) );
NAND3_X1 U736 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
NAND2_X1 U737 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
XNOR2_X1 U738 ( .A(n1033), .B(KEYINPUT52), .ZN(n1031) );
NAND3_X1 U739 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1029) );
XOR2_X1 U740 ( .A(KEYINPUT62), .B(n1036), .Z(n1034) );
NAND2_X1 U741 ( .A1(n1037), .A2(n1038), .ZN(n1028) );
NAND2_X1 U742 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
INV_X1 U743 ( .A(n1041), .ZN(n1009) );
NAND4_X1 U744 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1018), .ZN(n1005) );
XNOR2_X1 U745 ( .A(n1045), .B(G478), .ZN(n1043) );
XOR2_X1 U746 ( .A(n1046), .B(KEYINPUT1), .Z(n1042) );
NAND3_X1 U747 ( .A1(n1047), .A2(n1048), .A3(n1013), .ZN(n1046) );
XOR2_X1 U748 ( .A(KEYINPUT14), .B(n1036), .Z(n1047) );
XOR2_X1 U749 ( .A(n1049), .B(n1050), .Z(G72) );
XOR2_X1 U750 ( .A(n1051), .B(n1052), .Z(n1050) );
NAND2_X1 U751 ( .A1(G953), .A2(n1053), .ZN(n1052) );
NAND2_X1 U752 ( .A1(n1054), .A2(G227), .ZN(n1053) );
XNOR2_X1 U753 ( .A(G900), .B(KEYINPUT41), .ZN(n1054) );
NAND2_X1 U754 ( .A1(n1055), .A2(n1056), .ZN(n1051) );
NAND2_X1 U755 ( .A1(G953), .A2(n1057), .ZN(n1056) );
XOR2_X1 U756 ( .A(n1058), .B(KEYINPUT36), .Z(n1055) );
NAND2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U758 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
XNOR2_X1 U759 ( .A(n1063), .B(n1064), .ZN(n1062) );
XNOR2_X1 U760 ( .A(n1065), .B(KEYINPUT24), .ZN(n1061) );
NAND2_X1 U761 ( .A1(n1066), .A2(n1067), .ZN(n1059) );
XNOR2_X1 U762 ( .A(n1068), .B(n1063), .ZN(n1067) );
XNOR2_X1 U763 ( .A(KEYINPUT34), .B(n1069), .ZN(n1066) );
AND2_X1 U764 ( .A1(n1070), .A2(n1004), .ZN(n1049) );
NAND2_X1 U765 ( .A1(n1071), .A2(n1072), .ZN(G69) );
NAND2_X1 U766 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U767 ( .A1(G953), .A2(n1075), .ZN(n1074) );
NAND2_X1 U768 ( .A1(G898), .A2(G224), .ZN(n1075) );
NAND2_X1 U769 ( .A1(n1076), .A2(n1077), .ZN(n1071) );
NAND2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
OR2_X1 U771 ( .A1(n1004), .A2(G224), .ZN(n1079) );
INV_X1 U772 ( .A(n1073), .ZN(n1076) );
NAND2_X1 U773 ( .A1(n1080), .A2(n1081), .ZN(n1073) );
NAND2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
INV_X1 U775 ( .A(n1084), .ZN(n1082) );
NAND2_X1 U776 ( .A1(n1085), .A2(n1084), .ZN(n1080) );
NAND2_X1 U777 ( .A1(n1086), .A2(n1078), .ZN(n1084) );
INV_X1 U778 ( .A(n1087), .ZN(n1078) );
XOR2_X1 U779 ( .A(n1088), .B(n1089), .Z(n1086) );
XNOR2_X1 U780 ( .A(KEYINPUT59), .B(n1083), .ZN(n1085) );
NAND2_X1 U781 ( .A1(n1004), .A2(n1090), .ZN(n1083) );
NOR2_X1 U782 ( .A1(n1091), .A2(n1092), .ZN(G66) );
XNOR2_X1 U783 ( .A(n1093), .B(n1094), .ZN(n1092) );
NOR2_X1 U784 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U785 ( .A1(n1091), .A2(n1097), .ZN(G63) );
NOR3_X1 U786 ( .A1(n1045), .A2(n1098), .A3(n1099), .ZN(n1097) );
NOR4_X1 U787 ( .A1(n1100), .A2(n1096), .A3(KEYINPUT0), .A4(n1101), .ZN(n1099) );
NOR2_X1 U788 ( .A1(n1102), .A2(n1103), .ZN(n1098) );
NOR3_X1 U789 ( .A1(n1101), .A2(KEYINPUT0), .A3(n1104), .ZN(n1103) );
INV_X1 U790 ( .A(G478), .ZN(n1101) );
NOR3_X1 U791 ( .A1(n1105), .A2(n1091), .A3(n1106), .ZN(G60) );
NOR3_X1 U792 ( .A1(n1096), .A2(n1107), .A3(n1108), .ZN(n1106) );
INV_X1 U793 ( .A(n1109), .ZN(n1107) );
NOR2_X1 U794 ( .A1(n1110), .A2(n1111), .ZN(n1105) );
XNOR2_X1 U795 ( .A(n1109), .B(KEYINPUT43), .ZN(n1111) );
NOR2_X1 U796 ( .A1(n1108), .A2(n1096), .ZN(n1110) );
XOR2_X1 U797 ( .A(n1112), .B(n1113), .Z(G6) );
XNOR2_X1 U798 ( .A(G104), .B(KEYINPUT11), .ZN(n1113) );
NAND2_X1 U799 ( .A1(n1114), .A2(n999), .ZN(n1112) );
INV_X1 U800 ( .A(n1115), .ZN(n999) );
NOR2_X1 U801 ( .A1(n1091), .A2(n1116), .ZN(G57) );
XOR2_X1 U802 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U803 ( .A(n1119), .B(n1120), .Z(n1118) );
NOR2_X1 U804 ( .A1(n1121), .A2(n1096), .ZN(n1120) );
XOR2_X1 U805 ( .A(n1122), .B(n1123), .Z(n1117) );
NOR2_X1 U806 ( .A1(KEYINPUT16), .A2(n1124), .ZN(n1123) );
XOR2_X1 U807 ( .A(n1125), .B(KEYINPUT4), .Z(n1122) );
NAND2_X1 U808 ( .A1(KEYINPUT63), .A2(n1126), .ZN(n1125) );
XNOR2_X1 U809 ( .A(n1063), .B(n1127), .ZN(n1126) );
XOR2_X1 U810 ( .A(n1128), .B(KEYINPUT25), .Z(n1127) );
XNOR2_X1 U811 ( .A(G128), .B(n1129), .ZN(n1063) );
NOR2_X1 U812 ( .A1(n1091), .A2(n1130), .ZN(G54) );
XOR2_X1 U813 ( .A(n1129), .B(n1131), .Z(n1130) );
XOR2_X1 U814 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U815 ( .A1(n1134), .A2(n1096), .ZN(n1133) );
NAND2_X1 U816 ( .A1(G902), .A2(n1007), .ZN(n1096) );
INV_X1 U817 ( .A(n1104), .ZN(n1007) );
INV_X1 U818 ( .A(G469), .ZN(n1134) );
NOR2_X1 U819 ( .A1(n1091), .A2(n1135), .ZN(G51) );
XOR2_X1 U820 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U821 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR3_X1 U822 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
XNOR2_X1 U823 ( .A(n1104), .B(KEYINPUT31), .ZN(n1141) );
NOR2_X1 U824 ( .A1(n1070), .A2(n1090), .ZN(n1104) );
NAND4_X1 U825 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1090) );
AND4_X1 U826 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1146) );
NOR2_X1 U827 ( .A1(n1151), .A2(n1152), .ZN(n1145) );
NOR2_X1 U828 ( .A1(n1023), .A2(n1153), .ZN(n1152) );
NOR2_X1 U829 ( .A1(n1154), .A2(n1115), .ZN(n1151) );
NAND2_X1 U830 ( .A1(n1018), .A2(n1155), .ZN(n1115) );
NOR2_X1 U831 ( .A1(n1114), .A2(n1156), .ZN(n1154) );
XNOR2_X1 U832 ( .A(n998), .B(KEYINPUT53), .ZN(n1156) );
OR2_X1 U833 ( .A1(n1157), .A2(KEYINPUT6), .ZN(n1144) );
NAND4_X1 U834 ( .A1(n1158), .A2(n1159), .A3(n1015), .A4(KEYINPUT6), .ZN(n1143) );
AND2_X1 U835 ( .A1(n1033), .A2(n1037), .ZN(n1015) );
NAND4_X1 U836 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1070) );
AND4_X1 U837 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1163) );
OR2_X1 U838 ( .A1(n1040), .A2(n1168), .ZN(n1164) );
AND2_X1 U839 ( .A1(n1169), .A2(n1170), .ZN(n1162) );
NAND4_X1 U840 ( .A1(n1159), .A2(n1114), .A3(n1171), .A4(n1172), .ZN(n1160) );
OR2_X1 U841 ( .A1(n1173), .A2(KEYINPUT3), .ZN(n1172) );
NAND2_X1 U842 ( .A1(KEYINPUT3), .A2(n1174), .ZN(n1171) );
NAND2_X1 U843 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XNOR2_X1 U844 ( .A(n1177), .B(n1178), .ZN(n1136) );
NAND2_X1 U845 ( .A1(n1179), .A2(n1180), .ZN(n1177) );
NAND2_X1 U846 ( .A1(n1181), .A2(G125), .ZN(n1180) );
XOR2_X1 U847 ( .A(n1182), .B(KEYINPUT30), .Z(n1179) );
OR2_X1 U848 ( .A1(n1181), .A2(G125), .ZN(n1182) );
NOR2_X1 U849 ( .A1(n1004), .A2(G952), .ZN(n1091) );
XNOR2_X1 U850 ( .A(G146), .B(n1183), .ZN(G48) );
NAND3_X1 U851 ( .A1(n1159), .A2(n1114), .A3(n1173), .ZN(n1183) );
XNOR2_X1 U852 ( .A(G143), .B(n1167), .ZN(G45) );
NAND4_X1 U853 ( .A1(n1017), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1167) );
NOR2_X1 U854 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XNOR2_X1 U855 ( .A(G140), .B(n1166), .ZN(G42) );
NAND4_X1 U856 ( .A1(n1173), .A2(n1114), .A3(n1013), .A4(n1016), .ZN(n1166) );
XNOR2_X1 U857 ( .A(G137), .B(n1165), .ZN(G39) );
NAND4_X1 U858 ( .A1(n1033), .A2(n1173), .A3(n1013), .A4(n1189), .ZN(n1165) );
XNOR2_X1 U859 ( .A(G134), .B(n1190), .ZN(G36) );
NAND4_X1 U860 ( .A1(n1191), .A2(n1173), .A3(n998), .A4(n1017), .ZN(n1190) );
XNOR2_X1 U861 ( .A(n1013), .B(KEYINPUT17), .ZN(n1191) );
NAND2_X1 U862 ( .A1(n1192), .A2(n1193), .ZN(G33) );
NAND2_X1 U863 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
XNOR2_X1 U864 ( .A(KEYINPUT27), .B(n1161), .ZN(n1194) );
NAND2_X1 U865 ( .A1(n1196), .A2(G131), .ZN(n1192) );
XNOR2_X1 U866 ( .A(KEYINPUT8), .B(n1161), .ZN(n1196) );
OR2_X1 U867 ( .A1(n1168), .A2(n1039), .ZN(n1161) );
INV_X1 U868 ( .A(n1114), .ZN(n1039) );
NAND3_X1 U869 ( .A1(n1013), .A2(n1017), .A3(n1173), .ZN(n1168) );
NOR2_X1 U870 ( .A1(n1197), .A2(n1025), .ZN(n1013) );
XNOR2_X1 U871 ( .A(G128), .B(n1170), .ZN(G30) );
NAND3_X1 U872 ( .A1(n1159), .A2(n998), .A3(n1173), .ZN(n1170) );
INV_X1 U873 ( .A(n1187), .ZN(n1173) );
NAND2_X1 U874 ( .A1(n1032), .A2(n1175), .ZN(n1187) );
AND2_X1 U875 ( .A1(n1185), .A2(n1189), .ZN(n1159) );
XNOR2_X1 U876 ( .A(n1150), .B(n1198), .ZN(G3) );
NOR2_X1 U877 ( .A1(KEYINPUT49), .A2(n1199), .ZN(n1198) );
NAND3_X1 U878 ( .A1(n1155), .A2(n1017), .A3(n1033), .ZN(n1150) );
XNOR2_X1 U879 ( .A(G125), .B(n1169), .ZN(G27) );
NAND4_X1 U880 ( .A1(n1016), .A2(n1175), .A3(n1185), .A4(n1200), .ZN(n1169) );
AND2_X1 U881 ( .A1(n1037), .A2(n1114), .ZN(n1200) );
NAND2_X1 U882 ( .A1(n1041), .A2(n1201), .ZN(n1175) );
NAND4_X1 U883 ( .A1(G902), .A2(G953), .A3(n1202), .A4(n1057), .ZN(n1201) );
INV_X1 U884 ( .A(G900), .ZN(n1057) );
XOR2_X1 U885 ( .A(n1149), .B(n1203), .Z(G24) );
NOR2_X1 U886 ( .A1(G122), .A2(KEYINPUT56), .ZN(n1203) );
NAND4_X1 U887 ( .A1(n1204), .A2(n1205), .A3(n1018), .A4(n1184), .ZN(n1149) );
XNOR2_X1 U888 ( .A(G119), .B(n1157), .ZN(G21) );
NAND3_X1 U889 ( .A1(n1033), .A2(n1189), .A3(n1205), .ZN(n1157) );
NAND2_X1 U890 ( .A1(n1206), .A2(n1207), .ZN(n1189) );
NAND2_X1 U891 ( .A1(n1017), .A2(n1208), .ZN(n1207) );
NAND3_X1 U892 ( .A1(n1209), .A2(n1210), .A3(KEYINPUT47), .ZN(n1206) );
XNOR2_X1 U893 ( .A(KEYINPUT15), .B(n1211), .ZN(n1209) );
XOR2_X1 U894 ( .A(G116), .B(n1212), .Z(G18) );
NOR2_X1 U895 ( .A1(n1213), .A2(n1023), .ZN(n1212) );
XOR2_X1 U896 ( .A(n1153), .B(KEYINPUT33), .Z(n1213) );
NAND4_X1 U897 ( .A1(n1037), .A2(n998), .A3(n1017), .A4(n1214), .ZN(n1153) );
INV_X1 U898 ( .A(n1040), .ZN(n998) );
NAND2_X1 U899 ( .A1(n1188), .A2(n1184), .ZN(n1040) );
XNOR2_X1 U900 ( .A(G113), .B(n1148), .ZN(G15) );
NAND3_X1 U901 ( .A1(n1114), .A2(n1017), .A3(n1205), .ZN(n1148) );
AND2_X1 U902 ( .A1(n1037), .A2(n1215), .ZN(n1205) );
NOR2_X1 U903 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
INV_X1 U904 ( .A(n1048), .ZN(n1035) );
NAND2_X1 U905 ( .A1(n1216), .A2(n1217), .ZN(n1017) );
NAND2_X1 U906 ( .A1(n1018), .A2(n1218), .ZN(n1217) );
OR3_X1 U907 ( .A1(n1210), .A2(n1219), .A3(n1218), .ZN(n1216) );
INV_X1 U908 ( .A(KEYINPUT15), .ZN(n1218) );
NOR2_X1 U909 ( .A1(n1184), .A2(n1188), .ZN(n1114) );
XOR2_X1 U910 ( .A(n1147), .B(n1220), .Z(G12) );
NAND2_X1 U911 ( .A1(n1221), .A2(KEYINPUT10), .ZN(n1220) );
XNOR2_X1 U912 ( .A(G110), .B(KEYINPUT46), .ZN(n1221) );
NAND3_X1 U913 ( .A1(n1155), .A2(n1016), .A3(n1033), .ZN(n1147) );
NOR2_X1 U914 ( .A1(n1184), .A2(n1204), .ZN(n1033) );
INV_X1 U915 ( .A(n1188), .ZN(n1204) );
XNOR2_X1 U916 ( .A(n1044), .B(KEYINPUT5), .ZN(n1188) );
XNOR2_X1 U917 ( .A(n1222), .B(n1108), .ZN(n1044) );
INV_X1 U918 ( .A(G475), .ZN(n1108) );
NAND2_X1 U919 ( .A1(n1109), .A2(n1140), .ZN(n1222) );
XNOR2_X1 U920 ( .A(n1223), .B(n1224), .ZN(n1109) );
XOR2_X1 U921 ( .A(n1225), .B(n1226), .Z(n1224) );
XNOR2_X1 U922 ( .A(n1227), .B(n1228), .ZN(n1226) );
NOR2_X1 U923 ( .A1(KEYINPUT57), .A2(n1229), .ZN(n1228) );
NAND3_X1 U924 ( .A1(n1230), .A2(n1231), .A3(KEYINPUT61), .ZN(n1227) );
NAND2_X1 U925 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
INV_X1 U926 ( .A(KEYINPUT35), .ZN(n1233) );
XOR2_X1 U927 ( .A(n1234), .B(n1235), .Z(n1232) );
NAND2_X1 U928 ( .A1(KEYINPUT21), .A2(n1236), .ZN(n1234) );
NAND3_X1 U929 ( .A1(n1237), .A2(n1236), .A3(KEYINPUT35), .ZN(n1230) );
XOR2_X1 U930 ( .A(KEYINPUT21), .B(n1235), .Z(n1237) );
NOR2_X1 U931 ( .A1(n1238), .A2(n1239), .ZN(n1235) );
INV_X1 U932 ( .A(G214), .ZN(n1238) );
XOR2_X1 U933 ( .A(n1240), .B(n1241), .Z(n1223) );
XNOR2_X1 U934 ( .A(n1195), .B(G122), .ZN(n1241) );
INV_X1 U935 ( .A(G131), .ZN(n1195) );
NAND2_X1 U936 ( .A1(n1242), .A2(n1243), .ZN(n1240) );
NAND2_X1 U937 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XNOR2_X1 U938 ( .A(G125), .B(KEYINPUT9), .ZN(n1245) );
XNOR2_X1 U939 ( .A(G140), .B(KEYINPUT51), .ZN(n1244) );
XOR2_X1 U940 ( .A(n1246), .B(KEYINPUT20), .Z(n1242) );
NAND2_X1 U941 ( .A1(G125), .A2(n1247), .ZN(n1246) );
NAND2_X1 U942 ( .A1(n1248), .A2(n1249), .ZN(n1184) );
NAND2_X1 U943 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
XNOR2_X1 U944 ( .A(KEYINPUT29), .B(n1252), .ZN(n1251) );
XNOR2_X1 U945 ( .A(G478), .B(KEYINPUT60), .ZN(n1250) );
XOR2_X1 U946 ( .A(KEYINPUT48), .B(n1253), .Z(n1248) );
NOR2_X1 U947 ( .A1(G478), .A2(n1252), .ZN(n1253) );
INV_X1 U948 ( .A(n1045), .ZN(n1252) );
NOR2_X1 U949 ( .A1(n1102), .A2(G902), .ZN(n1045) );
INV_X1 U950 ( .A(n1100), .ZN(n1102) );
NAND2_X1 U951 ( .A1(n1254), .A2(n1255), .ZN(n1100) );
NAND3_X1 U952 ( .A1(n1256), .A2(n1257), .A3(G217), .ZN(n1255) );
XOR2_X1 U953 ( .A(n1258), .B(n1259), .Z(n1257) );
NAND2_X1 U954 ( .A1(n1260), .A2(n1261), .ZN(n1254) );
NAND2_X1 U955 ( .A1(G217), .A2(n1256), .ZN(n1261) );
XNOR2_X1 U956 ( .A(n1259), .B(n1258), .ZN(n1260) );
XNOR2_X1 U957 ( .A(n1262), .B(n1263), .ZN(n1258) );
XNOR2_X1 U958 ( .A(G116), .B(G122), .ZN(n1262) );
XOR2_X1 U959 ( .A(G134), .B(n1264), .Z(n1259) );
XNOR2_X1 U960 ( .A(KEYINPUT37), .B(n1236), .ZN(n1264) );
NAND2_X1 U961 ( .A1(n1265), .A2(n1266), .ZN(n1016) );
NAND2_X1 U962 ( .A1(n1018), .A2(n1208), .ZN(n1266) );
INV_X1 U963 ( .A(KEYINPUT47), .ZN(n1208) );
NOR2_X1 U964 ( .A1(n1210), .A2(n1211), .ZN(n1018) );
INV_X1 U965 ( .A(n1219), .ZN(n1211) );
NAND3_X1 U966 ( .A1(n1210), .A2(n1219), .A3(KEYINPUT47), .ZN(n1265) );
XNOR2_X1 U967 ( .A(n1267), .B(n1268), .ZN(n1219) );
XNOR2_X1 U968 ( .A(KEYINPUT54), .B(n1121), .ZN(n1268) );
INV_X1 U969 ( .A(G472), .ZN(n1121) );
NAND2_X1 U970 ( .A1(n1269), .A2(n1140), .ZN(n1267) );
XOR2_X1 U971 ( .A(n1270), .B(n1271), .Z(n1269) );
XNOR2_X1 U972 ( .A(n1124), .B(n1119), .ZN(n1271) );
XNOR2_X1 U973 ( .A(G113), .B(n1272), .ZN(n1119) );
NOR2_X1 U974 ( .A1(KEYINPUT12), .A2(n1273), .ZN(n1272) );
XOR2_X1 U975 ( .A(G101), .B(n1274), .Z(n1124) );
NOR2_X1 U976 ( .A1(n1239), .A2(n1275), .ZN(n1274) );
INV_X1 U977 ( .A(G210), .ZN(n1275) );
NAND2_X1 U978 ( .A1(n1276), .A2(n1277), .ZN(n1239) );
XOR2_X1 U979 ( .A(n1129), .B(n1278), .Z(n1270) );
XNOR2_X1 U980 ( .A(n1279), .B(KEYINPUT22), .ZN(n1278) );
NAND2_X1 U981 ( .A1(KEYINPUT7), .A2(n1181), .ZN(n1279) );
XOR2_X1 U982 ( .A(n1280), .B(n1095), .Z(n1210) );
NAND2_X1 U983 ( .A1(G217), .A2(n1281), .ZN(n1095) );
NAND2_X1 U984 ( .A1(n1140), .A2(n1093), .ZN(n1280) );
NAND2_X1 U985 ( .A1(n1282), .A2(n1283), .ZN(n1093) );
NAND2_X1 U986 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U987 ( .A(n1286), .B(KEYINPUT44), .Z(n1282) );
OR2_X1 U988 ( .A1(n1285), .A2(n1284), .ZN(n1286) );
XNOR2_X1 U989 ( .A(G137), .B(n1287), .ZN(n1284) );
AND2_X1 U990 ( .A1(n1256), .A2(G221), .ZN(n1287) );
AND2_X1 U991 ( .A1(G234), .A2(n1276), .ZN(n1256) );
XNOR2_X1 U992 ( .A(n1288), .B(n1289), .ZN(n1285) );
XNOR2_X1 U993 ( .A(n1229), .B(n1290), .ZN(n1289) );
NOR2_X1 U994 ( .A1(KEYINPUT55), .A2(n1069), .ZN(n1290) );
INV_X1 U995 ( .A(n1065), .ZN(n1069) );
XNOR2_X1 U996 ( .A(G140), .B(n1291), .ZN(n1065) );
NAND2_X1 U997 ( .A1(n1292), .A2(n1293), .ZN(n1288) );
NAND2_X1 U998 ( .A1(G110), .A2(n1294), .ZN(n1293) );
XOR2_X1 U999 ( .A(n1295), .B(KEYINPUT28), .Z(n1292) );
OR2_X1 U1000 ( .A1(n1294), .A2(G110), .ZN(n1295) );
XNOR2_X1 U1001 ( .A(G119), .B(n1296), .ZN(n1294) );
AND2_X1 U1002 ( .A1(n1032), .A2(n1215), .ZN(n1155) );
NOR2_X1 U1003 ( .A1(n1023), .A2(n1158), .ZN(n1215) );
INV_X1 U1004 ( .A(n1214), .ZN(n1158) );
NAND2_X1 U1005 ( .A1(n1041), .A2(n1297), .ZN(n1214) );
NAND3_X1 U1006 ( .A1(n1087), .A2(n1202), .A3(G902), .ZN(n1297) );
NOR2_X1 U1007 ( .A1(n1004), .A2(G898), .ZN(n1087) );
NAND3_X1 U1008 ( .A1(n1202), .A2(n1004), .A3(n1298), .ZN(n1041) );
XNOR2_X1 U1009 ( .A(KEYINPUT18), .B(n1003), .ZN(n1298) );
INV_X1 U1010 ( .A(G952), .ZN(n1003) );
NAND2_X1 U1011 ( .A1(G237), .A2(G234), .ZN(n1202) );
INV_X1 U1012 ( .A(n1185), .ZN(n1023) );
NOR2_X1 U1013 ( .A1(n1026), .A2(n1025), .ZN(n1185) );
AND2_X1 U1014 ( .A1(G214), .A2(n1299), .ZN(n1025) );
INV_X1 U1015 ( .A(n1197), .ZN(n1026) );
XOR2_X1 U1016 ( .A(n1300), .B(n1142), .Z(n1197) );
NAND2_X1 U1017 ( .A1(G210), .A2(n1299), .ZN(n1142) );
NAND2_X1 U1018 ( .A1(n1277), .A2(n1140), .ZN(n1299) );
INV_X1 U1019 ( .A(G237), .ZN(n1277) );
NAND2_X1 U1020 ( .A1(n1301), .A2(n1140), .ZN(n1300) );
XOR2_X1 U1021 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U1022 ( .A(n1138), .B(n1181), .Z(n1303) );
XNOR2_X1 U1023 ( .A(n1128), .B(n1296), .ZN(n1181) );
NAND3_X1 U1024 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n1128) );
NAND2_X1 U1025 ( .A1(G146), .A2(n1307), .ZN(n1306) );
NAND2_X1 U1026 ( .A1(n1308), .A2(n1236), .ZN(n1307) );
INV_X1 U1027 ( .A(G143), .ZN(n1236) );
OR3_X1 U1028 ( .A1(n1308), .A2(G143), .A3(KEYINPUT58), .ZN(n1305) );
XOR2_X1 U1029 ( .A(n1309), .B(G146), .Z(n1308) );
XNOR2_X1 U1030 ( .A(KEYINPUT40), .B(KEYINPUT32), .ZN(n1309) );
NAND2_X1 U1031 ( .A1(KEYINPUT58), .A2(G143), .ZN(n1304) );
XNOR2_X1 U1032 ( .A(n1088), .B(n1310), .ZN(n1138) );
NOR2_X1 U1033 ( .A1(KEYINPUT26), .A2(n1089), .ZN(n1310) );
XNOR2_X1 U1034 ( .A(n1311), .B(n1312), .ZN(n1089) );
XOR2_X1 U1035 ( .A(n1273), .B(n1225), .Z(n1312) );
XOR2_X1 U1036 ( .A(G104), .B(G113), .Z(n1225) );
XOR2_X1 U1037 ( .A(G116), .B(G119), .Z(n1273) );
XNOR2_X1 U1038 ( .A(G101), .B(n1313), .ZN(n1311) );
XNOR2_X1 U1039 ( .A(KEYINPUT38), .B(n1314), .ZN(n1313) );
INV_X1 U1040 ( .A(G107), .ZN(n1314) );
XOR2_X1 U1041 ( .A(G110), .B(G122), .Z(n1088) );
XNOR2_X1 U1042 ( .A(n1315), .B(n1291), .ZN(n1302) );
INV_X1 U1043 ( .A(G125), .ZN(n1291) );
NAND2_X1 U1044 ( .A1(KEYINPUT42), .A2(n1178), .ZN(n1315) );
NAND2_X1 U1045 ( .A1(G224), .A2(n1276), .ZN(n1178) );
INV_X1 U1046 ( .A(n1176), .ZN(n1032) );
NAND2_X1 U1047 ( .A1(n1036), .A2(n1048), .ZN(n1176) );
NAND2_X1 U1048 ( .A1(G221), .A2(n1281), .ZN(n1048) );
NAND2_X1 U1049 ( .A1(G234), .A2(n1140), .ZN(n1281) );
XNOR2_X1 U1050 ( .A(n1316), .B(G469), .ZN(n1036) );
NAND2_X1 U1051 ( .A1(n1317), .A2(n1140), .ZN(n1316) );
INV_X1 U1052 ( .A(G902), .ZN(n1140) );
XOR2_X1 U1053 ( .A(n1132), .B(n1318), .Z(n1317) );
XNOR2_X1 U1054 ( .A(n1319), .B(KEYINPUT2), .ZN(n1318) );
NAND2_X1 U1055 ( .A1(KEYINPUT39), .A2(n1129), .ZN(n1319) );
XOR2_X1 U1056 ( .A(n1320), .B(n1321), .Z(n1129) );
XOR2_X1 U1057 ( .A(KEYINPUT19), .B(G137), .Z(n1321) );
XNOR2_X1 U1058 ( .A(G134), .B(G131), .ZN(n1320) );
XOR2_X1 U1059 ( .A(n1322), .B(n1323), .Z(n1132) );
XOR2_X1 U1060 ( .A(n1324), .B(n1325), .Z(n1323) );
XNOR2_X1 U1061 ( .A(G104), .B(n1199), .ZN(n1325) );
INV_X1 U1062 ( .A(G101), .ZN(n1199) );
XNOR2_X1 U1063 ( .A(n1247), .B(G110), .ZN(n1324) );
INV_X1 U1064 ( .A(G140), .ZN(n1247) );
XNOR2_X1 U1065 ( .A(n1263), .B(n1326), .ZN(n1322) );
XNOR2_X1 U1066 ( .A(n1064), .B(n1327), .ZN(n1326) );
NAND2_X1 U1067 ( .A1(G227), .A2(n1276), .ZN(n1327) );
XNOR2_X1 U1068 ( .A(n1004), .B(KEYINPUT13), .ZN(n1276) );
INV_X1 U1069 ( .A(G953), .ZN(n1004) );
INV_X1 U1070 ( .A(n1068), .ZN(n1064) );
NAND2_X1 U1071 ( .A1(n1328), .A2(n1329), .ZN(n1068) );
NAND2_X1 U1072 ( .A1(G143), .A2(n1229), .ZN(n1329) );
XOR2_X1 U1073 ( .A(KEYINPUT50), .B(n1330), .Z(n1328) );
NOR2_X1 U1074 ( .A1(G143), .A2(n1229), .ZN(n1330) );
INV_X1 U1075 ( .A(G146), .ZN(n1229) );
XNOR2_X1 U1076 ( .A(G107), .B(n1296), .ZN(n1263) );
INV_X1 U1077 ( .A(G128), .ZN(n1296) );
endmodule


