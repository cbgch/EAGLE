//Key = 1110001001000110101100100010001010101001100110111001111011110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
n1422, n1423, n1424;

XNOR2_X1 U772 ( .A(G107), .B(n1082), .ZN(G9) );
NOR2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(G75) );
NOR3_X1 U774 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
NAND3_X1 U775 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1085) );
NAND2_X1 U776 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U777 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND4_X1 U778 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1094) );
NAND3_X1 U779 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
INV_X1 U780 ( .A(n1102), .ZN(n1101) );
NAND3_X1 U781 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1100) );
INV_X1 U782 ( .A(KEYINPUT7), .ZN(n1105) );
NAND2_X1 U783 ( .A1(KEYINPUT7), .A2(n1106), .ZN(n1099) );
NAND3_X1 U784 ( .A1(n1106), .A2(n1104), .A3(n1107), .ZN(n1093) );
NAND2_X1 U785 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND3_X1 U786 ( .A1(n1096), .A2(n1110), .A3(n1095), .ZN(n1109) );
OR2_X1 U787 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U788 ( .A1(n1097), .A2(n1113), .ZN(n1108) );
NAND2_X1 U789 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U790 ( .A1(n1095), .A2(n1116), .ZN(n1115) );
NAND2_X1 U791 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U792 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U793 ( .A1(n1096), .A2(n1121), .ZN(n1114) );
NAND2_X1 U794 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U795 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
INV_X1 U796 ( .A(n1126), .ZN(n1091) );
AND3_X1 U797 ( .A1(n1088), .A2(n1089), .A3(n1127), .ZN(n1083) );
NAND4_X1 U798 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1088) );
NOR4_X1 U799 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1131) );
AND3_X1 U800 ( .A1(KEYINPUT34), .A2(n1136), .A3(G478), .ZN(n1135) );
NOR2_X1 U801 ( .A1(KEYINPUT34), .A2(G478), .ZN(n1134) );
XNOR2_X1 U802 ( .A(G469), .B(n1137), .ZN(n1133) );
NAND3_X1 U803 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1132) );
XOR2_X1 U804 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U805 ( .A1(n1143), .A2(KEYINPUT4), .ZN(n1142) );
XOR2_X1 U806 ( .A(n1144), .B(KEYINPUT43), .Z(n1141) );
XNOR2_X1 U807 ( .A(n1145), .B(KEYINPUT23), .ZN(n1138) );
NOR3_X1 U808 ( .A1(n1124), .A2(n1146), .A3(n1103), .ZN(n1130) );
NAND2_X1 U809 ( .A1(G475), .A2(n1147), .ZN(n1128) );
XOR2_X1 U810 ( .A(n1148), .B(n1149), .Z(G72) );
NOR2_X1 U811 ( .A1(n1089), .A2(n1150), .ZN(n1149) );
XOR2_X1 U812 ( .A(KEYINPUT3), .B(n1151), .Z(n1150) );
NOR2_X1 U813 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U814 ( .A1(n1154), .A2(n1155), .ZN(n1148) );
NAND2_X1 U815 ( .A1(n1156), .A2(n1089), .ZN(n1155) );
XOR2_X1 U816 ( .A(n1086), .B(n1157), .Z(n1156) );
NAND3_X1 U817 ( .A1(G900), .A2(n1157), .A3(G953), .ZN(n1154) );
XNOR2_X1 U818 ( .A(n1158), .B(n1159), .ZN(n1157) );
XOR2_X1 U819 ( .A(KEYINPUT33), .B(n1160), .Z(n1159) );
NOR2_X1 U820 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XOR2_X1 U821 ( .A(KEYINPUT35), .B(n1163), .Z(n1162) );
NOR2_X1 U822 ( .A1(G140), .A2(n1164), .ZN(n1163) );
AND2_X1 U823 ( .A1(n1164), .A2(G140), .ZN(n1161) );
XOR2_X1 U824 ( .A(n1165), .B(n1166), .Z(n1158) );
XOR2_X1 U825 ( .A(n1167), .B(n1168), .Z(G69) );
NAND2_X1 U826 ( .A1(G953), .A2(n1169), .ZN(n1168) );
NAND2_X1 U827 ( .A1(G898), .A2(G224), .ZN(n1169) );
NAND4_X1 U828 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1167) );
OR3_X1 U829 ( .A1(n1174), .A2(n1175), .A3(KEYINPUT12), .ZN(n1173) );
NAND2_X1 U830 ( .A1(KEYINPUT12), .A2(n1176), .ZN(n1172) );
NAND2_X1 U831 ( .A1(G953), .A2(n1177), .ZN(n1171) );
NAND2_X1 U832 ( .A1(n1175), .A2(n1174), .ZN(n1170) );
NAND2_X1 U833 ( .A1(KEYINPUT51), .A2(n1178), .ZN(n1174) );
INV_X1 U834 ( .A(n1176), .ZN(n1178) );
NAND2_X1 U835 ( .A1(n1089), .A2(n1087), .ZN(n1176) );
NOR2_X1 U836 ( .A1(n1179), .A2(n1180), .ZN(G66) );
XNOR2_X1 U837 ( .A(n1181), .B(n1182), .ZN(n1180) );
NOR2_X1 U838 ( .A1(n1144), .A2(n1183), .ZN(n1182) );
NOR2_X1 U839 ( .A1(n1179), .A2(n1184), .ZN(G63) );
XNOR2_X1 U840 ( .A(n1185), .B(n1186), .ZN(n1184) );
NOR2_X1 U841 ( .A1(n1187), .A2(n1183), .ZN(n1186) );
INV_X1 U842 ( .A(G478), .ZN(n1187) );
NOR2_X1 U843 ( .A1(n1179), .A2(n1188), .ZN(G60) );
XOR2_X1 U844 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U845 ( .A1(n1191), .A2(n1183), .ZN(n1190) );
NAND2_X1 U846 ( .A1(KEYINPUT14), .A2(n1192), .ZN(n1189) );
XNOR2_X1 U847 ( .A(G104), .B(n1193), .ZN(G6) );
NOR2_X1 U848 ( .A1(n1179), .A2(n1194), .ZN(G57) );
XOR2_X1 U849 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U850 ( .A(n1197), .B(n1198), .Z(n1196) );
NOR2_X1 U851 ( .A1(n1199), .A2(n1183), .ZN(n1198) );
NOR2_X1 U852 ( .A1(n1200), .A2(n1201), .ZN(n1197) );
XNOR2_X1 U853 ( .A(n1202), .B(KEYINPUT19), .ZN(n1201) );
XNOR2_X1 U854 ( .A(n1203), .B(n1204), .ZN(n1195) );
NOR3_X1 U855 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(G54) );
AND2_X1 U856 ( .A1(KEYINPUT13), .A2(n1179), .ZN(n1207) );
NOR3_X1 U857 ( .A1(KEYINPUT13), .A2(n1089), .A3(n1127), .ZN(n1206) );
INV_X1 U858 ( .A(G952), .ZN(n1127) );
XOR2_X1 U859 ( .A(n1208), .B(n1209), .Z(n1205) );
XOR2_X1 U860 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U861 ( .A(n1165), .B(n1212), .Z(n1211) );
XOR2_X1 U862 ( .A(n1213), .B(n1214), .Z(n1208) );
XOR2_X1 U863 ( .A(n1215), .B(n1216), .Z(n1214) );
NOR3_X1 U864 ( .A1(n1183), .A2(KEYINPUT11), .A3(n1217), .ZN(n1216) );
NOR3_X1 U865 ( .A1(n1179), .A2(n1218), .A3(n1219), .ZN(G51) );
NOR2_X1 U866 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
XOR2_X1 U867 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR2_X1 U868 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NOR2_X1 U869 ( .A1(n1226), .A2(n1227), .ZN(n1218) );
XOR2_X1 U870 ( .A(n1222), .B(n1228), .Z(n1227) );
NOR2_X1 U871 ( .A1(n1229), .A2(n1225), .ZN(n1228) );
INV_X1 U872 ( .A(KEYINPUT61), .ZN(n1225) );
XOR2_X1 U873 ( .A(n1175), .B(n1230), .Z(n1222) );
NOR2_X1 U874 ( .A1(n1231), .A2(n1183), .ZN(n1230) );
NAND2_X1 U875 ( .A1(G902), .A2(n1232), .ZN(n1183) );
OR2_X1 U876 ( .A1(n1087), .A2(n1086), .ZN(n1232) );
NAND4_X1 U877 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1086) );
NOR4_X1 U878 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1236) );
NOR2_X1 U879 ( .A1(n1241), .A2(n1242), .ZN(n1235) );
INV_X1 U880 ( .A(n1243), .ZN(n1241) );
NAND2_X1 U881 ( .A1(n1244), .A2(n1245), .ZN(n1234) );
NAND2_X1 U882 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
OR3_X1 U883 ( .A1(n1248), .A2(KEYINPUT30), .A3(n1249), .ZN(n1247) );
XOR2_X1 U884 ( .A(KEYINPUT18), .B(n1250), .Z(n1246) );
NAND2_X1 U885 ( .A1(KEYINPUT30), .A2(n1251), .ZN(n1233) );
NAND4_X1 U886 ( .A1(n1252), .A2(n1253), .A3(n1254), .A4(n1255), .ZN(n1087) );
NOR4_X1 U887 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1255) );
INV_X1 U888 ( .A(n1082), .ZN(n1256) );
NAND3_X1 U889 ( .A1(n1096), .A2(n1111), .A3(n1260), .ZN(n1082) );
AND2_X1 U890 ( .A1(n1261), .A2(n1193), .ZN(n1254) );
NAND3_X1 U891 ( .A1(n1260), .A2(n1096), .A3(n1112), .ZN(n1193) );
NAND2_X1 U892 ( .A1(n1244), .A2(n1262), .ZN(n1253) );
NAND2_X1 U893 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
NAND2_X1 U894 ( .A1(KEYINPUT27), .A2(n1265), .ZN(n1264) );
OR2_X1 U895 ( .A1(n1266), .A2(KEYINPUT27), .ZN(n1252) );
NOR2_X1 U896 ( .A1(n1089), .A2(G952), .ZN(n1179) );
XNOR2_X1 U897 ( .A(G146), .B(n1267), .ZN(G48) );
NAND2_X1 U898 ( .A1(n1250), .A2(n1244), .ZN(n1267) );
AND2_X1 U899 ( .A1(n1268), .A2(n1112), .ZN(n1250) );
XNOR2_X1 U900 ( .A(n1269), .B(n1251), .ZN(G45) );
AND3_X1 U901 ( .A1(n1248), .A2(n1244), .A3(n1270), .ZN(n1251) );
XOR2_X1 U902 ( .A(G140), .B(n1242), .Z(G42) );
AND3_X1 U903 ( .A1(n1095), .A2(n1102), .A3(n1271), .ZN(n1242) );
NAND2_X1 U904 ( .A1(n1272), .A2(n1273), .ZN(G39) );
NAND2_X1 U905 ( .A1(n1240), .A2(n1274), .ZN(n1273) );
XOR2_X1 U906 ( .A(KEYINPUT22), .B(n1275), .Z(n1272) );
NOR2_X1 U907 ( .A1(n1240), .A2(n1274), .ZN(n1275) );
AND3_X1 U908 ( .A1(n1268), .A2(n1097), .A3(n1095), .ZN(n1240) );
XOR2_X1 U909 ( .A(G134), .B(n1239), .Z(G36) );
AND3_X1 U910 ( .A1(n1095), .A2(n1111), .A3(n1270), .ZN(n1239) );
XOR2_X1 U911 ( .A(n1276), .B(n1277), .Z(G33) );
XOR2_X1 U912 ( .A(KEYINPUT26), .B(G131), .Z(n1277) );
NAND2_X1 U913 ( .A1(KEYINPUT56), .A2(n1238), .ZN(n1276) );
AND3_X1 U914 ( .A1(n1095), .A2(n1112), .A3(n1270), .ZN(n1238) );
INV_X1 U915 ( .A(n1249), .ZN(n1270) );
NAND3_X1 U916 ( .A1(n1102), .A2(n1278), .A3(n1279), .ZN(n1249) );
AND2_X1 U917 ( .A1(n1125), .A2(n1280), .ZN(n1095) );
XOR2_X1 U918 ( .A(G128), .B(n1237), .Z(G30) );
AND3_X1 U919 ( .A1(n1244), .A2(n1111), .A3(n1268), .ZN(n1237) );
AND4_X1 U920 ( .A1(n1102), .A2(n1120), .A3(n1145), .A4(n1278), .ZN(n1268) );
XNOR2_X1 U921 ( .A(G101), .B(n1261), .ZN(G3) );
NAND3_X1 U922 ( .A1(n1260), .A2(n1097), .A3(n1279), .ZN(n1261) );
XNOR2_X1 U923 ( .A(G125), .B(n1243), .ZN(G27) );
NAND4_X1 U924 ( .A1(n1271), .A2(n1244), .A3(n1106), .A4(n1104), .ZN(n1243) );
AND4_X1 U925 ( .A1(n1119), .A2(n1112), .A3(n1120), .A4(n1278), .ZN(n1271) );
NAND2_X1 U926 ( .A1(n1126), .A2(n1281), .ZN(n1278) );
NAND4_X1 U927 ( .A1(G953), .A2(G902), .A3(n1282), .A4(n1153), .ZN(n1281) );
INV_X1 U928 ( .A(G900), .ZN(n1153) );
NAND2_X1 U929 ( .A1(n1283), .A2(n1284), .ZN(G24) );
NAND2_X1 U930 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
XNOR2_X1 U931 ( .A(KEYINPUT38), .B(n1266), .ZN(n1285) );
INV_X1 U932 ( .A(n1287), .ZN(n1266) );
NAND2_X1 U933 ( .A1(G122), .A2(n1288), .ZN(n1283) );
XNOR2_X1 U934 ( .A(n1287), .B(KEYINPUT20), .ZN(n1288) );
NOR2_X1 U935 ( .A1(n1265), .A2(n1122), .ZN(n1287) );
NAND3_X1 U936 ( .A1(n1096), .A2(n1248), .A3(n1289), .ZN(n1265) );
NOR2_X1 U937 ( .A1(n1145), .A2(n1120), .ZN(n1096) );
XNOR2_X1 U938 ( .A(n1290), .B(n1259), .ZN(G21) );
AND4_X1 U939 ( .A1(n1120), .A2(n1145), .A3(n1097), .A4(n1291), .ZN(n1259) );
NOR2_X1 U940 ( .A1(n1122), .A2(n1292), .ZN(n1291) );
XOR2_X1 U941 ( .A(n1293), .B(n1294), .Z(G18) );
NOR2_X1 U942 ( .A1(n1295), .A2(n1122), .ZN(n1294) );
XOR2_X1 U943 ( .A(n1263), .B(KEYINPUT60), .Z(n1295) );
NAND3_X1 U944 ( .A1(n1289), .A2(n1111), .A3(n1279), .ZN(n1263) );
NAND2_X1 U945 ( .A1(n1296), .A2(n1297), .ZN(n1111) );
OR3_X1 U946 ( .A1(n1298), .A2(n1299), .A3(KEYINPUT8), .ZN(n1297) );
NAND2_X1 U947 ( .A1(KEYINPUT8), .A2(n1248), .ZN(n1296) );
NOR2_X1 U948 ( .A1(n1299), .A2(n1300), .ZN(n1248) );
INV_X1 U949 ( .A(n1292), .ZN(n1289) );
NAND2_X1 U950 ( .A1(KEYINPUT2), .A2(n1301), .ZN(n1293) );
XOR2_X1 U951 ( .A(G113), .B(n1258), .Z(G15) );
NOR4_X1 U952 ( .A1(n1117), .A2(n1292), .A3(n1302), .A4(n1122), .ZN(n1258) );
INV_X1 U953 ( .A(n1244), .ZN(n1122) );
NAND3_X1 U954 ( .A1(n1106), .A2(n1104), .A3(n1303), .ZN(n1292) );
INV_X1 U955 ( .A(n1279), .ZN(n1117) );
NOR2_X1 U956 ( .A1(n1120), .A2(n1119), .ZN(n1279) );
XNOR2_X1 U957 ( .A(G110), .B(n1304), .ZN(G12) );
NAND2_X1 U958 ( .A1(KEYINPUT47), .A2(n1257), .ZN(n1304) );
AND4_X1 U959 ( .A1(n1119), .A2(n1260), .A3(n1097), .A4(n1120), .ZN(n1257) );
XOR2_X1 U960 ( .A(n1305), .B(n1144), .Z(n1120) );
NAND2_X1 U961 ( .A1(G217), .A2(n1306), .ZN(n1144) );
XNOR2_X1 U962 ( .A(n1143), .B(KEYINPUT31), .ZN(n1305) );
AND2_X1 U963 ( .A1(n1307), .A2(n1181), .ZN(n1143) );
XNOR2_X1 U964 ( .A(n1308), .B(G110), .ZN(n1181) );
XOR2_X1 U965 ( .A(n1309), .B(n1310), .Z(n1308) );
XOR2_X1 U966 ( .A(n1311), .B(n1312), .Z(n1310) );
XNOR2_X1 U967 ( .A(n1274), .B(G125), .ZN(n1312) );
INV_X1 U968 ( .A(G137), .ZN(n1274) );
XOR2_X1 U969 ( .A(KEYINPUT59), .B(KEYINPUT45), .Z(n1311) );
XOR2_X1 U970 ( .A(n1313), .B(n1314), .Z(n1309) );
XOR2_X1 U971 ( .A(n1315), .B(n1316), .Z(n1314) );
NOR2_X1 U972 ( .A1(G146), .A2(KEYINPUT24), .ZN(n1315) );
XOR2_X1 U973 ( .A(n1317), .B(n1318), .Z(n1313) );
AND4_X1 U974 ( .A1(n1319), .A2(n1089), .A3(G234), .A4(G221), .ZN(n1318) );
INV_X1 U975 ( .A(KEYINPUT49), .ZN(n1319) );
NAND2_X1 U976 ( .A1(n1320), .A2(n1321), .ZN(n1317) );
NAND2_X1 U977 ( .A1(n1322), .A2(n1290), .ZN(n1321) );
XOR2_X1 U978 ( .A(KEYINPUT44), .B(n1323), .Z(n1320) );
NOR2_X1 U979 ( .A1(n1322), .A2(n1290), .ZN(n1323) );
NAND2_X1 U980 ( .A1(n1324), .A2(n1325), .ZN(n1097) );
NAND3_X1 U981 ( .A1(n1299), .A2(n1300), .A3(n1326), .ZN(n1325) );
INV_X1 U982 ( .A(KEYINPUT8), .ZN(n1326) );
INV_X1 U983 ( .A(n1298), .ZN(n1300) );
NAND2_X1 U984 ( .A1(KEYINPUT8), .A2(n1112), .ZN(n1324) );
INV_X1 U985 ( .A(n1302), .ZN(n1112) );
NAND2_X1 U986 ( .A1(n1299), .A2(n1298), .ZN(n1302) );
NAND3_X1 U987 ( .A1(n1327), .A2(n1328), .A3(n1129), .ZN(n1298) );
NAND2_X1 U988 ( .A1(n1329), .A2(n1191), .ZN(n1129) );
OR3_X1 U989 ( .A1(n1191), .A2(n1329), .A3(KEYINPUT15), .ZN(n1328) );
INV_X1 U990 ( .A(n1147), .ZN(n1329) );
NAND2_X1 U991 ( .A1(n1192), .A2(n1307), .ZN(n1147) );
XOR2_X1 U992 ( .A(n1330), .B(n1331), .Z(n1192) );
XOR2_X1 U993 ( .A(n1332), .B(n1333), .Z(n1331) );
XOR2_X1 U994 ( .A(G131), .B(G113), .Z(n1333) );
XNOR2_X1 U995 ( .A(G146), .B(n1269), .ZN(n1332) );
XOR2_X1 U996 ( .A(n1334), .B(n1335), .Z(n1330) );
XNOR2_X1 U997 ( .A(n1336), .B(n1337), .ZN(n1335) );
AND3_X1 U998 ( .A1(G214), .A2(n1089), .A3(n1338), .ZN(n1336) );
XNOR2_X1 U999 ( .A(n1339), .B(n1340), .ZN(n1334) );
NAND3_X1 U1000 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1339) );
NAND2_X1 U1001 ( .A1(G125), .A2(n1344), .ZN(n1343) );
NAND3_X1 U1002 ( .A1(n1345), .A2(n1164), .A3(KEYINPUT46), .ZN(n1342) );
INV_X1 U1003 ( .A(G125), .ZN(n1164) );
INV_X1 U1004 ( .A(n1344), .ZN(n1345) );
NAND2_X1 U1005 ( .A1(KEYINPUT48), .A2(n1316), .ZN(n1344) );
OR2_X1 U1006 ( .A1(n1316), .A2(KEYINPUT46), .ZN(n1341) );
XOR2_X1 U1007 ( .A(G140), .B(KEYINPUT40), .Z(n1316) );
NAND2_X1 U1008 ( .A1(KEYINPUT15), .A2(n1191), .ZN(n1327) );
INV_X1 U1009 ( .A(G475), .ZN(n1191) );
NOR2_X1 U1010 ( .A1(n1146), .A2(n1346), .ZN(n1299) );
AND2_X1 U1011 ( .A1(G478), .A2(n1136), .ZN(n1346) );
NOR2_X1 U1012 ( .A1(n1136), .A2(G478), .ZN(n1146) );
NAND2_X1 U1013 ( .A1(n1307), .A2(n1185), .ZN(n1136) );
NAND2_X1 U1014 ( .A1(n1347), .A2(n1348), .ZN(n1185) );
NAND4_X1 U1015 ( .A1(G217), .A2(G234), .A3(n1349), .A4(n1089), .ZN(n1348) );
XOR2_X1 U1016 ( .A(n1350), .B(KEYINPUT63), .Z(n1347) );
NAND2_X1 U1017 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
NAND3_X1 U1018 ( .A1(G234), .A2(n1089), .A3(G217), .ZN(n1352) );
INV_X1 U1019 ( .A(n1349), .ZN(n1351) );
XNOR2_X1 U1020 ( .A(n1353), .B(n1354), .ZN(n1349) );
XOR2_X1 U1021 ( .A(n1355), .B(n1356), .Z(n1354) );
XNOR2_X1 U1022 ( .A(n1301), .B(G107), .ZN(n1356) );
INV_X1 U1023 ( .A(G116), .ZN(n1301) );
XOR2_X1 U1024 ( .A(KEYINPUT37), .B(G134), .Z(n1355) );
XNOR2_X1 U1025 ( .A(n1357), .B(n1322), .ZN(n1353) );
XNOR2_X1 U1026 ( .A(n1358), .B(n1337), .ZN(n1357) );
NAND2_X1 U1027 ( .A1(KEYINPUT9), .A2(n1269), .ZN(n1358) );
AND3_X1 U1028 ( .A1(n1244), .A2(n1303), .A3(n1102), .ZN(n1260) );
NOR2_X1 U1029 ( .A1(n1104), .A2(n1103), .ZN(n1102) );
INV_X1 U1030 ( .A(n1106), .ZN(n1103) );
NAND2_X1 U1031 ( .A1(G221), .A2(n1306), .ZN(n1106) );
NAND2_X1 U1032 ( .A1(n1359), .A2(n1360), .ZN(n1306) );
XNOR2_X1 U1033 ( .A(G234), .B(KEYINPUT58), .ZN(n1359) );
NAND2_X1 U1034 ( .A1(n1361), .A2(n1362), .ZN(n1104) );
NAND2_X1 U1035 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
NAND2_X1 U1036 ( .A1(KEYINPUT32), .A2(n1365), .ZN(n1364) );
NAND2_X1 U1037 ( .A1(G469), .A2(n1366), .ZN(n1365) );
INV_X1 U1038 ( .A(n1137), .ZN(n1363) );
NAND2_X1 U1039 ( .A1(n1367), .A2(n1217), .ZN(n1361) );
INV_X1 U1040 ( .A(G469), .ZN(n1217) );
NAND2_X1 U1041 ( .A1(n1366), .A2(n1368), .ZN(n1367) );
NAND2_X1 U1042 ( .A1(KEYINPUT32), .A2(n1137), .ZN(n1368) );
NAND3_X1 U1043 ( .A1(n1369), .A2(n1370), .A3(n1307), .ZN(n1137) );
NAND2_X1 U1044 ( .A1(KEYINPUT52), .A2(n1371), .ZN(n1370) );
XOR2_X1 U1045 ( .A(n1372), .B(n1373), .Z(n1371) );
OR3_X1 U1046 ( .A1(n1372), .A2(n1373), .A3(KEYINPUT52), .ZN(n1369) );
XOR2_X1 U1047 ( .A(n1212), .B(n1374), .Z(n1373) );
XNOR2_X1 U1048 ( .A(n1375), .B(n1376), .ZN(n1374) );
NOR2_X1 U1049 ( .A1(KEYINPUT29), .A2(n1165), .ZN(n1376) );
XOR2_X1 U1050 ( .A(n1377), .B(n1378), .Z(n1165) );
XNOR2_X1 U1051 ( .A(n1379), .B(n1380), .ZN(n1377) );
NOR2_X1 U1052 ( .A1(KEYINPUT41), .A2(n1322), .ZN(n1380) );
NOR2_X1 U1053 ( .A1(G146), .A2(KEYINPUT21), .ZN(n1379) );
NAND2_X1 U1054 ( .A1(KEYINPUT0), .A2(n1210), .ZN(n1375) );
XOR2_X1 U1055 ( .A(G101), .B(n1381), .Z(n1212) );
XNOR2_X1 U1056 ( .A(n1382), .B(G104), .ZN(n1381) );
XOR2_X1 U1057 ( .A(n1383), .B(n1215), .Z(n1372) );
NOR2_X1 U1058 ( .A1(n1152), .A2(G953), .ZN(n1215) );
INV_X1 U1059 ( .A(G227), .ZN(n1152) );
NAND2_X1 U1060 ( .A1(KEYINPUT16), .A2(n1213), .ZN(n1383) );
XOR2_X1 U1061 ( .A(G110), .B(G140), .Z(n1213) );
INV_X1 U1062 ( .A(KEYINPUT10), .ZN(n1366) );
NAND2_X1 U1063 ( .A1(n1126), .A2(n1384), .ZN(n1303) );
NAND4_X1 U1064 ( .A1(G953), .A2(G902), .A3(n1282), .A4(n1177), .ZN(n1384) );
INV_X1 U1065 ( .A(G898), .ZN(n1177) );
NAND3_X1 U1066 ( .A1(n1282), .A2(n1089), .A3(G952), .ZN(n1126) );
NAND2_X1 U1067 ( .A1(G237), .A2(G234), .ZN(n1282) );
NOR2_X1 U1068 ( .A1(n1125), .A2(n1124), .ZN(n1244) );
INV_X1 U1069 ( .A(n1280), .ZN(n1124) );
NAND2_X1 U1070 ( .A1(G214), .A2(n1385), .ZN(n1280) );
XNOR2_X1 U1071 ( .A(n1139), .B(KEYINPUT39), .ZN(n1125) );
XNOR2_X1 U1072 ( .A(n1386), .B(n1231), .ZN(n1139) );
NAND2_X1 U1073 ( .A1(G210), .A2(n1385), .ZN(n1231) );
NAND2_X1 U1074 ( .A1(n1338), .A2(n1360), .ZN(n1385) );
INV_X1 U1075 ( .A(G902), .ZN(n1360) );
NAND2_X1 U1076 ( .A1(n1387), .A2(n1307), .ZN(n1386) );
XOR2_X1 U1077 ( .A(n1388), .B(n1175), .Z(n1387) );
XOR2_X1 U1078 ( .A(n1389), .B(n1390), .Z(n1175) );
XNOR2_X1 U1079 ( .A(n1391), .B(n1392), .ZN(n1390) );
XOR2_X1 U1080 ( .A(KEYINPUT6), .B(G110), .Z(n1392) );
XOR2_X1 U1081 ( .A(n1393), .B(n1394), .Z(n1389) );
XOR2_X1 U1082 ( .A(n1395), .B(n1396), .Z(n1393) );
NOR2_X1 U1083 ( .A1(KEYINPUT28), .A2(n1337), .ZN(n1396) );
XOR2_X1 U1084 ( .A(n1286), .B(KEYINPUT1), .Z(n1337) );
INV_X1 U1085 ( .A(G122), .ZN(n1286) );
NAND3_X1 U1086 ( .A1(n1397), .A2(n1398), .A3(n1399), .ZN(n1395) );
NAND2_X1 U1087 ( .A1(G104), .A2(n1382), .ZN(n1399) );
INV_X1 U1088 ( .A(G107), .ZN(n1382) );
NAND2_X1 U1089 ( .A1(n1400), .A2(n1401), .ZN(n1398) );
INV_X1 U1090 ( .A(KEYINPUT36), .ZN(n1401) );
NAND2_X1 U1091 ( .A1(n1402), .A2(n1340), .ZN(n1400) );
XNOR2_X1 U1092 ( .A(KEYINPUT54), .B(G107), .ZN(n1402) );
NAND2_X1 U1093 ( .A1(KEYINPUT36), .A2(n1403), .ZN(n1397) );
NAND2_X1 U1094 ( .A1(n1404), .A2(n1405), .ZN(n1403) );
OR2_X1 U1095 ( .A1(G107), .A2(KEYINPUT54), .ZN(n1405) );
NAND3_X1 U1096 ( .A1(G107), .A2(n1340), .A3(KEYINPUT54), .ZN(n1404) );
INV_X1 U1097 ( .A(G104), .ZN(n1340) );
NAND2_X1 U1098 ( .A1(n1406), .A2(n1407), .ZN(n1388) );
NAND2_X1 U1099 ( .A1(n1408), .A2(n1220), .ZN(n1407) );
XNOR2_X1 U1100 ( .A(n1229), .B(KEYINPUT17), .ZN(n1408) );
NAND2_X1 U1101 ( .A1(n1409), .A2(n1226), .ZN(n1406) );
INV_X1 U1102 ( .A(n1220), .ZN(n1226) );
NAND2_X1 U1103 ( .A1(G224), .A2(n1089), .ZN(n1220) );
XNOR2_X1 U1104 ( .A(n1224), .B(n1410), .ZN(n1409) );
XOR2_X1 U1105 ( .A(KEYINPUT62), .B(KEYINPUT53), .Z(n1410) );
INV_X1 U1106 ( .A(n1229), .ZN(n1224) );
XNOR2_X1 U1107 ( .A(G125), .B(n1411), .ZN(n1229) );
INV_X1 U1108 ( .A(n1145), .ZN(n1119) );
XOR2_X1 U1109 ( .A(n1412), .B(n1199), .Z(n1145) );
INV_X1 U1110 ( .A(G472), .ZN(n1199) );
NAND2_X1 U1111 ( .A1(n1307), .A2(n1413), .ZN(n1412) );
XOR2_X1 U1112 ( .A(n1414), .B(n1415), .Z(n1413) );
NOR2_X1 U1113 ( .A1(n1202), .A2(n1200), .ZN(n1415) );
NOR2_X1 U1114 ( .A1(n1391), .A2(n1416), .ZN(n1200) );
AND2_X1 U1115 ( .A1(n1416), .A2(n1391), .ZN(n1202) );
INV_X1 U1116 ( .A(G101), .ZN(n1391) );
NAND3_X1 U1117 ( .A1(n1338), .A2(n1089), .A3(G210), .ZN(n1416) );
INV_X1 U1118 ( .A(G953), .ZN(n1089) );
INV_X1 U1119 ( .A(G237), .ZN(n1338) );
NOR2_X1 U1120 ( .A1(KEYINPUT55), .A2(n1417), .ZN(n1414) );
XNOR2_X1 U1121 ( .A(n1204), .B(n1418), .ZN(n1417) );
NOR2_X1 U1122 ( .A1(KEYINPUT42), .A2(n1411), .ZN(n1418) );
INV_X1 U1123 ( .A(n1203), .ZN(n1411) );
XNOR2_X1 U1124 ( .A(n1419), .B(n1378), .ZN(n1203) );
XNOR2_X1 U1125 ( .A(n1269), .B(KEYINPUT50), .ZN(n1378) );
INV_X1 U1126 ( .A(G143), .ZN(n1269) );
XOR2_X1 U1127 ( .A(G146), .B(n1322), .Z(n1419) );
XNOR2_X1 U1128 ( .A(G128), .B(KEYINPUT57), .ZN(n1322) );
XNOR2_X1 U1129 ( .A(n1210), .B(n1394), .ZN(n1204) );
XOR2_X1 U1130 ( .A(G113), .B(n1420), .Z(n1394) );
XNOR2_X1 U1131 ( .A(n1290), .B(G116), .ZN(n1420) );
INV_X1 U1132 ( .A(G119), .ZN(n1290) );
NAND2_X1 U1133 ( .A1(n1421), .A2(n1422), .ZN(n1210) );
NAND2_X1 U1134 ( .A1(n1166), .A2(n1423), .ZN(n1422) );
INV_X1 U1135 ( .A(KEYINPUT5), .ZN(n1423) );
XOR2_X1 U1136 ( .A(G131), .B(n1424), .Z(n1166) );
NAND3_X1 U1137 ( .A1(G131), .A2(n1424), .A3(KEYINPUT5), .ZN(n1421) );
XOR2_X1 U1138 ( .A(G134), .B(G137), .Z(n1424) );
XNOR2_X1 U1139 ( .A(G902), .B(KEYINPUT25), .ZN(n1307) );
endmodule


