//Key = 0110111110011001111001110100101000001111011011100000010010011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410;

XNOR2_X1 U771 ( .A(G107), .B(n1063), .ZN(G9) );
NOR2_X1 U772 ( .A1(n1064), .A2(n1065), .ZN(G75) );
NOR3_X1 U773 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
NOR2_X1 U774 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR4_X1 U775 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1069) );
NAND2_X1 U776 ( .A1(n1075), .A2(n1076), .ZN(n1071) );
NAND3_X1 U777 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1066) );
NAND2_X1 U778 ( .A1(n1075), .A2(n1080), .ZN(n1079) );
NAND2_X1 U779 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND3_X1 U780 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
NAND2_X1 U781 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NAND2_X1 U782 ( .A1(n1076), .A2(n1088), .ZN(n1087) );
NAND2_X1 U783 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U784 ( .A1(n1091), .A2(n1070), .ZN(n1090) );
INV_X1 U785 ( .A(KEYINPUT29), .ZN(n1070) );
NAND2_X1 U786 ( .A1(n1092), .A2(n1093), .ZN(n1086) );
NAND2_X1 U787 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND3_X1 U789 ( .A1(n1092), .A2(n1098), .A3(n1076), .ZN(n1081) );
INV_X1 U790 ( .A(n1099), .ZN(n1076) );
NAND2_X1 U791 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NAND2_X1 U792 ( .A1(n1085), .A2(n1102), .ZN(n1101) );
NAND2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U795 ( .A1(n1083), .A2(n1107), .ZN(n1100) );
NAND2_X1 U796 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U797 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
INV_X1 U798 ( .A(n1112), .ZN(n1110) );
INV_X1 U799 ( .A(n1113), .ZN(n1075) );
NOR3_X1 U800 ( .A1(n1114), .A2(G953), .A3(G952), .ZN(n1064) );
INV_X1 U801 ( .A(n1077), .ZN(n1114) );
NAND4_X1 U802 ( .A1(n1115), .A2(n1116), .A3(n1117), .A4(n1118), .ZN(n1077) );
NOR3_X1 U803 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1118) );
XOR2_X1 U804 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U805 ( .A(n1124), .B(n1125), .Z(n1120) );
NOR2_X1 U806 ( .A1(KEYINPUT43), .A2(n1126), .ZN(n1125) );
NAND3_X1 U807 ( .A1(n1127), .A2(n1128), .A3(n1112), .ZN(n1119) );
NOR3_X1 U808 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1117) );
AND3_X1 U809 ( .A1(KEYINPUT44), .A2(n1132), .A3(G478), .ZN(n1131) );
NOR2_X1 U810 ( .A1(KEYINPUT44), .A2(G478), .ZN(n1130) );
XOR2_X1 U811 ( .A(n1133), .B(n1134), .Z(n1129) );
XOR2_X1 U812 ( .A(n1135), .B(G469), .Z(n1116) );
XOR2_X1 U813 ( .A(n1136), .B(G472), .Z(n1115) );
NAND3_X1 U814 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(G72) );
NAND2_X1 U815 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
OR3_X1 U816 ( .A1(n1141), .A2(n1140), .A3(n1142), .ZN(n1138) );
INV_X1 U817 ( .A(n1143), .ZN(n1140) );
INV_X1 U818 ( .A(KEYINPUT30), .ZN(n1141) );
NAND2_X1 U819 ( .A1(n1144), .A2(n1142), .ZN(n1137) );
NAND2_X1 U820 ( .A1(G953), .A2(n1145), .ZN(n1142) );
NAND2_X1 U821 ( .A1(G900), .A2(G227), .ZN(n1145) );
NAND3_X1 U822 ( .A1(n1146), .A2(n1143), .A3(KEYINPUT30), .ZN(n1144) );
NAND3_X1 U823 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1143) );
NAND2_X1 U824 ( .A1(G953), .A2(n1150), .ZN(n1148) );
OR2_X1 U825 ( .A1(n1147), .A2(n1149), .ZN(n1146) );
XNOR2_X1 U826 ( .A(n1151), .B(n1152), .ZN(n1147) );
XOR2_X1 U827 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1151) );
XOR2_X1 U829 ( .A(KEYINPUT12), .B(G137), .Z(n1156) );
NAND2_X1 U830 ( .A1(n1157), .A2(n1158), .ZN(G69) );
NAND3_X1 U831 ( .A1(n1159), .A2(n1160), .A3(G953), .ZN(n1158) );
XOR2_X1 U832 ( .A(n1161), .B(KEYINPUT58), .Z(n1157) );
NAND3_X1 U833 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1161) );
NAND2_X1 U834 ( .A1(n1165), .A2(n1160), .ZN(n1164) );
OR3_X1 U835 ( .A1(n1160), .A2(n1165), .A3(G953), .ZN(n1163) );
AND2_X1 U836 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U837 ( .A(n1168), .B(KEYINPUT40), .Z(n1166) );
NAND2_X1 U838 ( .A1(G953), .A2(n1169), .ZN(n1162) );
OR2_X1 U839 ( .A1(n1160), .A2(n1159), .ZN(n1169) );
NAND2_X1 U840 ( .A1(G898), .A2(G224), .ZN(n1159) );
NAND2_X1 U841 ( .A1(n1170), .A2(n1171), .ZN(n1160) );
NAND2_X1 U842 ( .A1(G953), .A2(n1172), .ZN(n1171) );
XOR2_X1 U843 ( .A(n1173), .B(n1174), .Z(n1170) );
XOR2_X1 U844 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n1177), .ZN(n1175) );
NOR2_X1 U846 ( .A1(n1178), .A2(n1179), .ZN(G66) );
NOR3_X1 U847 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1179) );
NOR3_X1 U848 ( .A1(n1183), .A2(n1134), .A3(n1184), .ZN(n1182) );
NOR2_X1 U849 ( .A1(n1185), .A2(n1186), .ZN(n1181) );
NOR2_X1 U850 ( .A1(n1187), .A2(n1134), .ZN(n1185) );
NOR2_X1 U851 ( .A1(n1178), .A2(n1188), .ZN(G63) );
XOR2_X1 U852 ( .A(n1189), .B(n1190), .Z(n1188) );
NAND3_X1 U853 ( .A1(n1191), .A2(G478), .A3(KEYINPUT21), .ZN(n1189) );
NOR2_X1 U854 ( .A1(n1178), .A2(n1192), .ZN(G60) );
NOR3_X1 U855 ( .A1(n1124), .A2(n1193), .A3(n1194), .ZN(n1192) );
AND3_X1 U856 ( .A1(n1195), .A2(G475), .A3(n1191), .ZN(n1194) );
NOR2_X1 U857 ( .A1(n1196), .A2(n1195), .ZN(n1193) );
NOR2_X1 U858 ( .A1(n1187), .A2(n1126), .ZN(n1196) );
INV_X1 U859 ( .A(n1068), .ZN(n1187) );
XNOR2_X1 U860 ( .A(G104), .B(n1197), .ZN(G6) );
NAND4_X1 U861 ( .A1(n1198), .A2(n1199), .A3(n1083), .A4(n1200), .ZN(n1197) );
NOR2_X1 U862 ( .A1(n1178), .A2(n1201), .ZN(G57) );
XOR2_X1 U863 ( .A(n1202), .B(n1203), .Z(n1201) );
XOR2_X1 U864 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U865 ( .A(n1206), .B(n1207), .Z(n1202) );
NOR2_X1 U866 ( .A1(n1208), .A2(n1184), .ZN(n1207) );
NOR2_X1 U867 ( .A1(n1178), .A2(n1209), .ZN(G54) );
XOR2_X1 U868 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U869 ( .A(n1212), .B(n1213), .Z(n1211) );
XOR2_X1 U870 ( .A(n1214), .B(n1215), .Z(n1210) );
XOR2_X1 U871 ( .A(n1216), .B(n1217), .Z(n1215) );
AND2_X1 U872 ( .A1(G469), .A2(n1191), .ZN(n1217) );
INV_X1 U873 ( .A(n1184), .ZN(n1191) );
NAND2_X1 U874 ( .A1(KEYINPUT8), .A2(n1218), .ZN(n1214) );
NOR2_X1 U875 ( .A1(n1178), .A2(n1219), .ZN(G51) );
XOR2_X1 U876 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U877 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR2_X1 U878 ( .A1(n1122), .A2(n1184), .ZN(n1223) );
NAND2_X1 U879 ( .A1(G902), .A2(n1068), .ZN(n1184) );
NAND3_X1 U880 ( .A1(n1167), .A2(n1168), .A3(n1149), .ZN(n1068) );
AND2_X1 U881 ( .A1(n1224), .A2(n1225), .ZN(n1149) );
NOR4_X1 U882 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1225) );
INV_X1 U883 ( .A(n1230), .ZN(n1227) );
NOR4_X1 U884 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1224) );
NOR3_X1 U885 ( .A1(n1235), .A2(n1073), .A3(n1072), .ZN(n1234) );
INV_X1 U886 ( .A(n1236), .ZN(n1233) );
NAND3_X1 U887 ( .A1(n1237), .A2(n1199), .A3(n1238), .ZN(n1168) );
NOR3_X1 U888 ( .A1(n1074), .A2(n1239), .A3(n1108), .ZN(n1238) );
XNOR2_X1 U889 ( .A(n1240), .B(KEYINPUT31), .ZN(n1237) );
AND4_X1 U890 ( .A1(n1241), .A2(n1242), .A3(n1063), .A4(n1243), .ZN(n1167) );
NOR3_X1 U891 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1243) );
NOR4_X1 U892 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1244) );
XOR2_X1 U893 ( .A(n1074), .B(KEYINPUT52), .Z(n1248) );
NAND3_X1 U894 ( .A1(n1251), .A2(n1252), .A3(n1083), .ZN(n1063) );
INV_X1 U895 ( .A(n1074), .ZN(n1083) );
NAND2_X1 U896 ( .A1(n1200), .A2(n1253), .ZN(n1241) );
NAND2_X1 U897 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND3_X1 U898 ( .A1(n1092), .A2(n1256), .A3(n1198), .ZN(n1255) );
XOR2_X1 U899 ( .A(n1257), .B(KEYINPUT49), .Z(n1220) );
NAND3_X1 U900 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1257) );
INV_X1 U901 ( .A(n1261), .ZN(n1260) );
OR2_X1 U902 ( .A1(n1262), .A2(n1263), .ZN(n1259) );
NAND3_X1 U903 ( .A1(n1264), .A2(n1262), .A3(n1263), .ZN(n1258) );
NAND2_X1 U904 ( .A1(n1265), .A2(n1266), .ZN(n1262) );
XOR2_X1 U905 ( .A(n1267), .B(KEYINPUT11), .Z(n1265) );
NOR2_X1 U906 ( .A1(n1078), .A2(G952), .ZN(n1178) );
XOR2_X1 U907 ( .A(n1231), .B(n1268), .Z(G48) );
NOR2_X1 U908 ( .A1(KEYINPUT51), .A2(n1269), .ZN(n1268) );
XNOR2_X1 U909 ( .A(G146), .B(KEYINPUT26), .ZN(n1269) );
AND4_X1 U910 ( .A1(n1270), .A2(n1199), .A3(n1271), .A4(n1200), .ZN(n1231) );
NAND2_X1 U911 ( .A1(n1272), .A2(n1273), .ZN(G45) );
NAND2_X1 U912 ( .A1(n1229), .A2(n1274), .ZN(n1273) );
XOR2_X1 U913 ( .A(KEYINPUT39), .B(n1275), .Z(n1272) );
NOR2_X1 U914 ( .A1(n1229), .A2(n1274), .ZN(n1275) );
NOR4_X1 U915 ( .A1(n1250), .A2(n1235), .A3(n1108), .A4(n1247), .ZN(n1229) );
INV_X1 U916 ( .A(n1276), .ZN(n1250) );
XOR2_X1 U917 ( .A(G140), .B(n1228), .Z(G42) );
AND4_X1 U918 ( .A1(n1270), .A2(n1199), .A3(n1085), .A4(n1106), .ZN(n1228) );
XOR2_X1 U919 ( .A(n1277), .B(n1230), .Z(G39) );
NAND4_X1 U920 ( .A1(n1092), .A2(n1270), .A3(n1085), .A4(n1271), .ZN(n1230) );
INV_X1 U921 ( .A(n1072), .ZN(n1085) );
AND3_X1 U922 ( .A1(n1278), .A2(n1279), .A3(n1105), .ZN(n1270) );
XOR2_X1 U923 ( .A(G134), .B(n1280), .Z(G36) );
NOR3_X1 U924 ( .A1(n1235), .A2(n1281), .A3(n1073), .ZN(n1280) );
XOR2_X1 U925 ( .A(n1072), .B(KEYINPUT27), .Z(n1281) );
XOR2_X1 U926 ( .A(G131), .B(n1226), .Z(G33) );
NOR3_X1 U927 ( .A1(n1235), .A2(n1072), .A3(n1089), .ZN(n1226) );
NAND2_X1 U928 ( .A1(n1111), .A2(n1112), .ZN(n1072) );
NAND3_X1 U929 ( .A1(n1278), .A2(n1279), .A3(n1256), .ZN(n1235) );
XOR2_X1 U930 ( .A(n1282), .B(n1236), .Z(G30) );
NAND4_X1 U931 ( .A1(n1105), .A2(n1271), .A3(n1251), .A4(n1279), .ZN(n1236) );
NOR3_X1 U932 ( .A1(n1073), .A2(n1239), .A3(n1108), .ZN(n1251) );
XNOR2_X1 U933 ( .A(G101), .B(n1283), .ZN(G3) );
NAND4_X1 U934 ( .A1(n1284), .A2(n1198), .A3(n1092), .A4(n1256), .ZN(n1283) );
INV_X1 U935 ( .A(n1103), .ZN(n1256) );
XOR2_X1 U936 ( .A(n1108), .B(KEYINPUT38), .Z(n1284) );
NAND2_X1 U937 ( .A1(n1285), .A2(n1286), .ZN(G27) );
NAND2_X1 U938 ( .A1(n1287), .A2(n1267), .ZN(n1286) );
XOR2_X1 U939 ( .A(n1288), .B(KEYINPUT48), .Z(n1285) );
OR2_X1 U940 ( .A1(n1287), .A2(n1267), .ZN(n1288) );
NAND2_X1 U941 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
NAND3_X1 U942 ( .A1(n1291), .A2(n1089), .A3(n1292), .ZN(n1290) );
INV_X1 U943 ( .A(KEYINPUT17), .ZN(n1292) );
NAND2_X1 U944 ( .A1(n1232), .A2(KEYINPUT17), .ZN(n1289) );
AND2_X1 U945 ( .A1(n1291), .A2(n1199), .ZN(n1232) );
INV_X1 U946 ( .A(n1089), .ZN(n1199) );
AND4_X1 U947 ( .A1(n1279), .A2(n1106), .A3(n1200), .A4(n1293), .ZN(n1291) );
NOR2_X1 U948 ( .A1(n1099), .A2(n1294), .ZN(n1293) );
NAND2_X1 U949 ( .A1(n1113), .A2(n1295), .ZN(n1279) );
NAND4_X1 U950 ( .A1(G902), .A2(G953), .A3(n1296), .A4(n1150), .ZN(n1295) );
INV_X1 U951 ( .A(G900), .ZN(n1150) );
XNOR2_X1 U952 ( .A(G122), .B(n1297), .ZN(G24) );
NAND3_X1 U953 ( .A1(n1276), .A2(n1298), .A3(n1299), .ZN(n1297) );
NOR3_X1 U954 ( .A1(n1074), .A2(KEYINPUT61), .A3(n1247), .ZN(n1299) );
NAND2_X1 U955 ( .A1(n1294), .A2(n1106), .ZN(n1074) );
XNOR2_X1 U956 ( .A(G119), .B(n1242), .ZN(G21) );
NAND4_X1 U957 ( .A1(n1298), .A2(n1092), .A3(n1105), .A4(n1271), .ZN(n1242) );
XOR2_X1 U958 ( .A(G116), .B(n1246), .Z(G18) );
NOR3_X1 U959 ( .A1(n1103), .A2(n1073), .A3(n1249), .ZN(n1246) );
INV_X1 U960 ( .A(n1091), .ZN(n1073) );
NOR2_X1 U961 ( .A1(n1276), .A2(n1247), .ZN(n1091) );
XOR2_X1 U962 ( .A(n1245), .B(n1300), .Z(G15) );
NOR2_X1 U963 ( .A1(KEYINPUT34), .A2(n1301), .ZN(n1300) );
NOR3_X1 U964 ( .A1(n1089), .A2(n1103), .A3(n1249), .ZN(n1245) );
INV_X1 U965 ( .A(n1298), .ZN(n1249) );
NOR3_X1 U966 ( .A1(n1108), .A2(n1240), .A3(n1099), .ZN(n1298) );
NAND2_X1 U967 ( .A1(n1097), .A2(n1127), .ZN(n1099) );
INV_X1 U968 ( .A(n1200), .ZN(n1108) );
NAND2_X1 U969 ( .A1(n1271), .A2(n1294), .ZN(n1103) );
INV_X1 U970 ( .A(n1105), .ZN(n1294) );
INV_X1 U971 ( .A(n1106), .ZN(n1271) );
NAND2_X1 U972 ( .A1(n1302), .A2(n1276), .ZN(n1089) );
XOR2_X1 U973 ( .A(n1303), .B(KEYINPUT15), .Z(n1302) );
XOR2_X1 U974 ( .A(n1304), .B(n1305), .Z(G12) );
NAND2_X1 U975 ( .A1(KEYINPUT23), .A2(G110), .ZN(n1305) );
NAND2_X1 U976 ( .A1(n1306), .A2(n1200), .ZN(n1304) );
NOR2_X1 U977 ( .A1(n1111), .A2(n1307), .ZN(n1200) );
XOR2_X1 U978 ( .A(KEYINPUT6), .B(n1112), .Z(n1307) );
NAND2_X1 U979 ( .A1(G214), .A2(n1308), .ZN(n1112) );
XNOR2_X1 U980 ( .A(n1309), .B(n1310), .ZN(n1111) );
XNOR2_X1 U981 ( .A(KEYINPUT13), .B(n1122), .ZN(n1310) );
NAND2_X1 U982 ( .A1(G210), .A2(n1308), .ZN(n1122) );
NAND2_X1 U983 ( .A1(n1311), .A2(n1312), .ZN(n1308) );
NAND2_X1 U984 ( .A1(KEYINPUT16), .A2(n1123), .ZN(n1309) );
NAND2_X1 U985 ( .A1(n1313), .A2(n1312), .ZN(n1123) );
XOR2_X1 U986 ( .A(n1222), .B(n1314), .Z(n1313) );
NOR3_X1 U987 ( .A1(n1261), .A2(n1315), .A3(n1316), .ZN(n1314) );
NOR3_X1 U988 ( .A1(G125), .A2(n1204), .A3(n1317), .ZN(n1316) );
NOR2_X1 U989 ( .A1(n1267), .A2(n1318), .ZN(n1315) );
XOR2_X1 U990 ( .A(n1263), .B(n1204), .Z(n1318) );
NOR2_X1 U991 ( .A1(n1264), .A2(n1263), .ZN(n1261) );
INV_X1 U992 ( .A(n1317), .ZN(n1263) );
NAND2_X1 U993 ( .A1(G224), .A2(n1319), .ZN(n1317) );
NAND2_X1 U994 ( .A1(n1204), .A2(n1267), .ZN(n1264) );
INV_X1 U995 ( .A(n1266), .ZN(n1204) );
XOR2_X1 U996 ( .A(n1320), .B(n1176), .Z(n1222) );
XNOR2_X1 U997 ( .A(n1321), .B(n1322), .ZN(n1176) );
XOR2_X1 U998 ( .A(KEYINPUT55), .B(G110), .Z(n1322) );
NAND2_X1 U999 ( .A1(KEYINPUT5), .A2(G122), .ZN(n1321) );
NAND2_X1 U1000 ( .A1(n1323), .A2(n1324), .ZN(n1320) );
NAND2_X1 U1001 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1002 ( .A(KEYINPUT53), .B(n1327), .Z(n1323) );
NOR2_X1 U1003 ( .A1(n1326), .A2(n1325), .ZN(n1327) );
INV_X1 U1004 ( .A(n1177), .ZN(n1325) );
XOR2_X1 U1005 ( .A(n1254), .B(KEYINPUT59), .Z(n1306) );
NAND4_X1 U1006 ( .A1(n1198), .A2(n1092), .A3(n1105), .A4(n1106), .ZN(n1254) );
NAND3_X1 U1007 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1106) );
NAND2_X1 U1008 ( .A1(KEYINPUT50), .A2(n1331), .ZN(n1330) );
NAND3_X1 U1009 ( .A1(n1332), .A2(n1333), .A3(n1136), .ZN(n1329) );
INV_X1 U1010 ( .A(KEYINPUT50), .ZN(n1333) );
OR2_X1 U1011 ( .A1(n1136), .A2(n1332), .ZN(n1328) );
NOR2_X1 U1012 ( .A1(KEYINPUT20), .A2(n1331), .ZN(n1332) );
XOR2_X1 U1013 ( .A(n1208), .B(KEYINPUT4), .Z(n1331) );
INV_X1 U1014 ( .A(G472), .ZN(n1208) );
NAND2_X1 U1015 ( .A1(n1334), .A2(n1312), .ZN(n1136) );
XNOR2_X1 U1016 ( .A(n1205), .B(n1335), .ZN(n1334) );
NOR2_X1 U1017 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XOR2_X1 U1018 ( .A(KEYINPUT9), .B(n1338), .Z(n1337) );
NOR2_X1 U1019 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
XOR2_X1 U1020 ( .A(KEYINPUT14), .B(n1341), .Z(n1340) );
AND2_X1 U1021 ( .A1(n1339), .A2(n1341), .ZN(n1336) );
XNOR2_X1 U1022 ( .A(n1266), .B(KEYINPUT22), .ZN(n1341) );
XNOR2_X1 U1023 ( .A(n1342), .B(n1343), .ZN(n1266) );
NOR2_X1 U1024 ( .A1(KEYINPUT62), .A2(n1282), .ZN(n1343) );
XNOR2_X1 U1025 ( .A(n1344), .B(n1345), .ZN(n1205) );
XOR2_X1 U1026 ( .A(n1346), .B(n1326), .Z(n1345) );
INV_X1 U1027 ( .A(n1173), .ZN(n1326) );
XOR2_X1 U1028 ( .A(n1301), .B(n1347), .Z(n1173) );
XOR2_X1 U1029 ( .A(G119), .B(G116), .Z(n1347) );
XOR2_X1 U1030 ( .A(n1348), .B(KEYINPUT60), .Z(n1344) );
NAND2_X1 U1031 ( .A1(G210), .A2(n1349), .ZN(n1348) );
XOR2_X1 U1032 ( .A(n1350), .B(n1180), .Z(n1105) );
INV_X1 U1033 ( .A(n1133), .ZN(n1180) );
NAND2_X1 U1034 ( .A1(n1183), .A2(n1312), .ZN(n1133) );
INV_X1 U1035 ( .A(n1186), .ZN(n1183) );
XOR2_X1 U1036 ( .A(n1351), .B(n1352), .Z(n1186) );
XOR2_X1 U1037 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1038 ( .A(n1355), .B(n1356), .Z(n1354) );
AND3_X1 U1039 ( .A1(G234), .A2(G221), .A3(n1319), .ZN(n1356) );
NAND2_X1 U1040 ( .A1(KEYINPUT46), .A2(n1357), .ZN(n1353) );
XNOR2_X1 U1041 ( .A(G146), .B(n1358), .ZN(n1357) );
NAND2_X1 U1042 ( .A1(KEYINPUT1), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1043 ( .A(n1360), .B(n1361), .Z(n1359) );
XNOR2_X1 U1044 ( .A(KEYINPUT28), .B(G140), .ZN(n1361) );
NAND2_X1 U1045 ( .A1(KEYINPUT37), .A2(n1267), .ZN(n1360) );
XNOR2_X1 U1046 ( .A(G119), .B(n1362), .ZN(n1351) );
XOR2_X1 U1047 ( .A(G137), .B(G128), .Z(n1362) );
NAND2_X1 U1048 ( .A1(KEYINPUT18), .A2(n1134), .ZN(n1350) );
NAND2_X1 U1049 ( .A1(G217), .A2(n1363), .ZN(n1134) );
NOR2_X1 U1050 ( .A1(n1303), .A2(n1276), .ZN(n1092) );
XOR2_X1 U1051 ( .A(n1364), .B(n1124), .Z(n1276) );
NOR2_X1 U1052 ( .A1(n1195), .A2(G902), .ZN(n1124) );
XOR2_X1 U1053 ( .A(n1365), .B(n1366), .Z(n1195) );
XOR2_X1 U1054 ( .A(n1367), .B(n1368), .Z(n1366) );
XOR2_X1 U1055 ( .A(n1154), .B(n1342), .Z(n1368) );
XOR2_X1 U1056 ( .A(n1267), .B(n1369), .Z(n1154) );
XOR2_X1 U1057 ( .A(G140), .B(G131), .Z(n1369) );
INV_X1 U1058 ( .A(G125), .ZN(n1267) );
XOR2_X1 U1059 ( .A(n1370), .B(G104), .Z(n1367) );
NAND2_X1 U1060 ( .A1(G214), .A2(n1349), .ZN(n1370) );
AND2_X1 U1061 ( .A1(n1319), .A2(n1311), .ZN(n1349) );
INV_X1 U1062 ( .A(G237), .ZN(n1311) );
XOR2_X1 U1063 ( .A(n1371), .B(n1372), .Z(n1365) );
XOR2_X1 U1064 ( .A(KEYINPUT41), .B(KEYINPUT28), .Z(n1372) );
XOR2_X1 U1065 ( .A(n1301), .B(G122), .Z(n1371) );
INV_X1 U1066 ( .A(G113), .ZN(n1301) );
NAND2_X1 U1067 ( .A1(KEYINPUT2), .A2(n1126), .ZN(n1364) );
INV_X1 U1068 ( .A(G475), .ZN(n1126) );
XNOR2_X1 U1069 ( .A(n1247), .B(KEYINPUT47), .ZN(n1303) );
AND2_X1 U1070 ( .A1(n1128), .A2(n1373), .ZN(n1247) );
NAND2_X1 U1071 ( .A1(G478), .A2(n1132), .ZN(n1373) );
OR2_X1 U1072 ( .A1(n1132), .A2(G478), .ZN(n1128) );
NAND2_X1 U1073 ( .A1(n1190), .A2(n1312), .ZN(n1132) );
XNOR2_X1 U1074 ( .A(n1374), .B(n1375), .ZN(n1190) );
XOR2_X1 U1075 ( .A(n1376), .B(n1377), .Z(n1375) );
XNOR2_X1 U1076 ( .A(n1378), .B(n1379), .ZN(n1377) );
AND4_X1 U1077 ( .A1(n1380), .A2(n1319), .A3(G234), .A4(G217), .ZN(n1379) );
INV_X1 U1078 ( .A(KEYINPUT10), .ZN(n1380) );
NAND2_X1 U1079 ( .A1(KEYINPUT25), .A2(n1155), .ZN(n1378) );
NOR2_X1 U1080 ( .A1(n1381), .A2(n1382), .ZN(n1376) );
XOR2_X1 U1081 ( .A(KEYINPUT3), .B(n1383), .Z(n1382) );
NOR2_X1 U1082 ( .A1(G143), .A2(n1282), .ZN(n1383) );
INV_X1 U1083 ( .A(G128), .ZN(n1282) );
NOR2_X1 U1084 ( .A1(G128), .A2(n1274), .ZN(n1381) );
INV_X1 U1085 ( .A(G143), .ZN(n1274) );
XOR2_X1 U1086 ( .A(n1384), .B(n1385), .Z(n1374) );
XOR2_X1 U1087 ( .A(KEYINPUT24), .B(G122), .Z(n1385) );
XNOR2_X1 U1088 ( .A(G107), .B(G116), .ZN(n1384) );
NOR2_X1 U1089 ( .A1(n1239), .A2(n1240), .ZN(n1198) );
INV_X1 U1090 ( .A(n1252), .ZN(n1240) );
NAND2_X1 U1091 ( .A1(n1113), .A2(n1386), .ZN(n1252) );
NAND4_X1 U1092 ( .A1(n1387), .A2(G902), .A3(n1296), .A4(n1172), .ZN(n1386) );
INV_X1 U1093 ( .A(G898), .ZN(n1172) );
XOR2_X1 U1094 ( .A(n1078), .B(KEYINPUT42), .Z(n1387) );
NAND3_X1 U1095 ( .A1(n1296), .A2(n1078), .A3(G952), .ZN(n1113) );
NAND2_X1 U1096 ( .A1(G237), .A2(G234), .ZN(n1296) );
XOR2_X1 U1097 ( .A(n1094), .B(KEYINPUT57), .Z(n1239) );
INV_X1 U1098 ( .A(n1278), .ZN(n1094) );
NOR2_X1 U1099 ( .A1(n1097), .A2(n1096), .ZN(n1278) );
INV_X1 U1100 ( .A(n1127), .ZN(n1096) );
NAND2_X1 U1101 ( .A1(G221), .A2(n1363), .ZN(n1127) );
NAND2_X1 U1102 ( .A1(G234), .A2(n1312), .ZN(n1363) );
XNOR2_X1 U1103 ( .A(n1135), .B(n1388), .ZN(n1097) );
NOR2_X1 U1104 ( .A1(G469), .A2(KEYINPUT35), .ZN(n1388) );
NAND2_X1 U1105 ( .A1(n1389), .A2(n1312), .ZN(n1135) );
INV_X1 U1106 ( .A(G902), .ZN(n1312) );
XOR2_X1 U1107 ( .A(n1390), .B(n1218), .Z(n1389) );
XOR2_X1 U1108 ( .A(n1339), .B(KEYINPUT7), .Z(n1218) );
INV_X1 U1109 ( .A(n1206), .ZN(n1339) );
XOR2_X1 U1110 ( .A(n1391), .B(G131), .Z(n1206) );
NAND3_X1 U1111 ( .A1(n1392), .A2(n1393), .A3(n1394), .ZN(n1391) );
NAND2_X1 U1112 ( .A1(G137), .A2(n1155), .ZN(n1394) );
NAND2_X1 U1113 ( .A1(n1395), .A2(n1396), .ZN(n1393) );
INV_X1 U1114 ( .A(KEYINPUT63), .ZN(n1396) );
NAND2_X1 U1115 ( .A1(n1397), .A2(n1277), .ZN(n1395) );
XOR2_X1 U1116 ( .A(KEYINPUT36), .B(n1155), .Z(n1397) );
INV_X1 U1117 ( .A(G134), .ZN(n1155) );
NAND2_X1 U1118 ( .A1(KEYINPUT63), .A2(n1398), .ZN(n1392) );
NAND2_X1 U1119 ( .A1(n1399), .A2(n1400), .ZN(n1398) );
OR2_X1 U1120 ( .A1(G134), .A2(KEYINPUT36), .ZN(n1400) );
NAND3_X1 U1121 ( .A1(G134), .A2(n1277), .A3(KEYINPUT36), .ZN(n1399) );
INV_X1 U1122 ( .A(G137), .ZN(n1277) );
XOR2_X1 U1123 ( .A(n1401), .B(n1212), .Z(n1390) );
XOR2_X1 U1124 ( .A(n1153), .B(n1177), .Z(n1212) );
XOR2_X1 U1125 ( .A(n1402), .B(n1346), .Z(n1177) );
XOR2_X1 U1126 ( .A(G101), .B(KEYINPUT0), .Z(n1346) );
XNOR2_X1 U1127 ( .A(G104), .B(G107), .ZN(n1402) );
NAND2_X1 U1128 ( .A1(n1403), .A2(n1404), .ZN(n1153) );
NAND2_X1 U1129 ( .A1(G128), .A2(n1342), .ZN(n1404) );
XOR2_X1 U1130 ( .A(n1405), .B(KEYINPUT32), .Z(n1403) );
OR2_X1 U1131 ( .A1(n1342), .A2(G128), .ZN(n1405) );
XOR2_X1 U1132 ( .A(G146), .B(G143), .Z(n1342) );
NAND2_X1 U1133 ( .A1(n1406), .A2(n1407), .ZN(n1401) );
OR2_X1 U1134 ( .A1(n1216), .A2(n1408), .ZN(n1407) );
XOR2_X1 U1135 ( .A(n1409), .B(KEYINPUT54), .Z(n1406) );
NAND2_X1 U1136 ( .A1(n1408), .A2(n1216), .ZN(n1409) );
NAND2_X1 U1137 ( .A1(G227), .A2(n1319), .ZN(n1216) );
XOR2_X1 U1138 ( .A(n1078), .B(KEYINPUT19), .Z(n1319) );
INV_X1 U1139 ( .A(G953), .ZN(n1078) );
XOR2_X1 U1140 ( .A(n1213), .B(KEYINPUT56), .Z(n1408) );
XNOR2_X1 U1141 ( .A(n1355), .B(n1410), .ZN(n1213) );
XOR2_X1 U1142 ( .A(KEYINPUT45), .B(G140), .Z(n1410) );
INV_X1 U1143 ( .A(G110), .ZN(n1355) );
endmodule


