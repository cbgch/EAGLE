//Key = 1000101110110001000010011110000001100101011010111010111101010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290;

XOR2_X1 U715 ( .A(n990), .B(n991), .Z(G9) );
NOR2_X1 U716 ( .A1(KEYINPUT21), .A2(n992), .ZN(n991) );
NOR2_X1 U717 ( .A1(n993), .A2(n994), .ZN(G75) );
NOR4_X1 U718 ( .A1(n995), .A2(n996), .A3(n997), .A4(n998), .ZN(n994) );
XOR2_X1 U719 ( .A(KEYINPUT3), .B(n999), .Z(n998) );
NOR2_X1 U720 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NOR2_X1 U721 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NOR4_X1 U722 ( .A1(n1004), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n1003) );
NOR2_X1 U723 ( .A1(n1008), .A2(n1009), .ZN(n1005) );
NOR2_X1 U724 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NOR3_X1 U725 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1011) );
NOR2_X1 U726 ( .A1(n1015), .A2(n1016), .ZN(n1010) );
NOR2_X1 U727 ( .A1(n1017), .A2(n1018), .ZN(n1004) );
NOR2_X1 U728 ( .A1(n1012), .A2(n1019), .ZN(n1017) );
NOR4_X1 U729 ( .A1(n1008), .A2(n1020), .A3(n1019), .A4(n1012), .ZN(n1002) );
NOR3_X1 U730 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NOR2_X1 U731 ( .A1(n1024), .A2(n1006), .ZN(n1023) );
NOR2_X1 U732 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NOR2_X1 U733 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
XOR2_X1 U734 ( .A(KEYINPUT14), .B(n1029), .Z(n1028) );
NOR3_X1 U735 ( .A1(n1007), .A2(n1030), .A3(n1031), .ZN(n1022) );
NOR2_X1 U736 ( .A1(n1032), .A2(n1033), .ZN(n1021) );
XNOR2_X1 U737 ( .A(n1034), .B(KEYINPUT12), .ZN(n1032) );
NOR3_X1 U738 ( .A1(n996), .A2(G952), .A3(n995), .ZN(n993) );
AND4_X1 U739 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n995) );
NOR4_X1 U740 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1006), .ZN(n1038) );
XOR2_X1 U741 ( .A(n1042), .B(KEYINPUT26), .Z(n1041) );
NAND2_X1 U742 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
XOR2_X1 U743 ( .A(n1045), .B(n1046), .Z(n1040) );
NOR2_X1 U744 ( .A1(n1047), .A2(KEYINPUT16), .ZN(n1046) );
INV_X1 U745 ( .A(n1048), .ZN(n1047) );
XNOR2_X1 U746 ( .A(n1049), .B(KEYINPUT25), .ZN(n1039) );
NOR3_X1 U747 ( .A1(n1008), .A2(n1050), .A3(n1051), .ZN(n1037) );
NAND2_X1 U748 ( .A1(n1052), .A2(n1053), .ZN(n1036) );
XNOR2_X1 U749 ( .A(KEYINPUT62), .B(n1043), .ZN(n1052) );
XNOR2_X1 U750 ( .A(G469), .B(KEYINPUT51), .ZN(n1043) );
XOR2_X1 U751 ( .A(n1054), .B(n1055), .Z(G72) );
NOR2_X1 U752 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
AND2_X1 U753 ( .A1(G227), .A2(G900), .ZN(n1056) );
NAND2_X1 U754 ( .A1(n1058), .A2(n1059), .ZN(n1054) );
NAND2_X1 U755 ( .A1(n1060), .A2(n1057), .ZN(n1059) );
XOR2_X1 U756 ( .A(n1061), .B(n1062), .Z(n1060) );
NAND2_X1 U757 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NAND3_X1 U758 ( .A1(G900), .A2(n1062), .A3(G953), .ZN(n1058) );
XNOR2_X1 U759 ( .A(n1065), .B(n1066), .ZN(n1062) );
XNOR2_X1 U760 ( .A(n1067), .B(n1068), .ZN(n1066) );
XNOR2_X1 U761 ( .A(KEYINPUT7), .B(n1069), .ZN(n1068) );
XNOR2_X1 U762 ( .A(n1070), .B(n1071), .ZN(n1065) );
INV_X1 U763 ( .A(n1072), .ZN(n1071) );
NAND2_X1 U764 ( .A1(KEYINPUT44), .A2(n1073), .ZN(n1070) );
XOR2_X1 U765 ( .A(G137), .B(n1074), .Z(n1073) );
NAND2_X1 U766 ( .A1(n1075), .A2(n1076), .ZN(G69) );
NAND2_X1 U767 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
OR2_X1 U768 ( .A1(n1057), .A2(G224), .ZN(n1078) );
NAND3_X1 U769 ( .A1(G953), .A2(n1079), .A3(n1080), .ZN(n1075) );
XNOR2_X1 U770 ( .A(n1077), .B(KEYINPUT17), .ZN(n1080) );
XNOR2_X1 U771 ( .A(n1081), .B(n1082), .ZN(n1077) );
NOR3_X1 U772 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
NOR2_X1 U773 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U774 ( .A(n1088), .B(n1089), .Z(n1086) );
NOR2_X1 U775 ( .A1(n1090), .A2(n1091), .ZN(n1084) );
XOR2_X1 U776 ( .A(KEYINPUT54), .B(n1087), .Z(n1091) );
XNOR2_X1 U777 ( .A(G110), .B(n1092), .ZN(n1087) );
XNOR2_X1 U778 ( .A(n1088), .B(n1089), .ZN(n1090) );
NAND2_X1 U779 ( .A1(n1093), .A2(KEYINPUT4), .ZN(n1088) );
XOR2_X1 U780 ( .A(n1094), .B(n1095), .Z(n1093) );
XNOR2_X1 U781 ( .A(G113), .B(KEYINPUT13), .ZN(n1094) );
NAND2_X1 U782 ( .A1(n1057), .A2(n1096), .ZN(n1081) );
NAND2_X1 U783 ( .A1(G898), .A2(G224), .ZN(n1079) );
NOR2_X1 U784 ( .A1(n1097), .A2(n1098), .ZN(G66) );
XOR2_X1 U785 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U786 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR2_X1 U787 ( .A1(n1097), .A2(n1103), .ZN(G63) );
XNOR2_X1 U788 ( .A(n1104), .B(n1105), .ZN(n1103) );
AND2_X1 U789 ( .A1(G478), .A2(n1106), .ZN(n1105) );
NOR2_X1 U790 ( .A1(n1097), .A2(n1107), .ZN(G60) );
XOR2_X1 U791 ( .A(n1108), .B(n1109), .Z(n1107) );
AND2_X1 U792 ( .A1(G475), .A2(n1106), .ZN(n1108) );
XNOR2_X1 U793 ( .A(n1110), .B(n1111), .ZN(G6) );
NOR2_X1 U794 ( .A1(G104), .A2(KEYINPUT58), .ZN(n1111) );
NOR2_X1 U795 ( .A1(n1097), .A2(n1112), .ZN(G57) );
XOR2_X1 U796 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U797 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U798 ( .A1(KEYINPUT30), .A2(n1117), .ZN(n1115) );
XOR2_X1 U799 ( .A(n1118), .B(KEYINPUT45), .Z(n1117) );
XNOR2_X1 U800 ( .A(n1119), .B(n1120), .ZN(n1113) );
NOR2_X1 U801 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NOR2_X1 U802 ( .A1(KEYINPUT52), .A2(n1123), .ZN(n1122) );
INV_X1 U803 ( .A(n1124), .ZN(n1123) );
NOR2_X1 U804 ( .A1(KEYINPUT40), .A2(n1124), .ZN(n1121) );
NAND2_X1 U805 ( .A1(n1106), .A2(G472), .ZN(n1124) );
NOR3_X1 U806 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(G54) );
AND2_X1 U807 ( .A1(KEYINPUT39), .A2(n1097), .ZN(n1127) );
NOR3_X1 U808 ( .A1(KEYINPUT39), .A2(n1057), .A3(n1128), .ZN(n1126) );
INV_X1 U809 ( .A(G952), .ZN(n1128) );
XOR2_X1 U810 ( .A(n1129), .B(n1130), .Z(n1125) );
NOR2_X1 U811 ( .A1(KEYINPUT1), .A2(n1131), .ZN(n1130) );
AND2_X1 U812 ( .A1(G469), .A2(n1106), .ZN(n1129) );
INV_X1 U813 ( .A(n1102), .ZN(n1106) );
NOR2_X1 U814 ( .A1(n1097), .A2(n1132), .ZN(G51) );
XOR2_X1 U815 ( .A(n1133), .B(n1134), .Z(n1132) );
XNOR2_X1 U816 ( .A(n1135), .B(n1072), .ZN(n1134) );
XOR2_X1 U817 ( .A(G125), .B(n1136), .Z(n1072) );
XOR2_X1 U818 ( .A(n1137), .B(n1138), .Z(n1133) );
NOR2_X1 U819 ( .A1(n1048), .A2(n1102), .ZN(n1138) );
NAND2_X1 U820 ( .A1(G902), .A2(n997), .ZN(n1102) );
NAND3_X1 U821 ( .A1(n1139), .A2(n1063), .A3(n1140), .ZN(n997) );
XOR2_X1 U822 ( .A(n1064), .B(KEYINPUT28), .Z(n1140) );
AND4_X1 U823 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1063) );
AND4_X1 U824 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1144) );
OR2_X1 U825 ( .A1(n1149), .A2(n1150), .ZN(n1143) );
NAND3_X1 U826 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1142) );
NAND2_X1 U827 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NAND3_X1 U828 ( .A1(n1007), .A2(n1149), .A3(n1013), .ZN(n1155) );
INV_X1 U829 ( .A(KEYINPUT41), .ZN(n1149) );
OR2_X1 U830 ( .A1(n1156), .A2(n1007), .ZN(n1141) );
INV_X1 U831 ( .A(n1096), .ZN(n1139) );
NAND4_X1 U832 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1096) );
NOR4_X1 U833 ( .A1(n990), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1160) );
AND3_X1 U834 ( .A1(n1164), .A2(n1165), .A3(n1014), .ZN(n990) );
NOR2_X1 U835 ( .A1(n1110), .A2(n1166), .ZN(n1159) );
NOR3_X1 U836 ( .A1(n1019), .A2(n1167), .A3(n1033), .ZN(n1166) );
AND3_X1 U837 ( .A1(n1164), .A2(n1165), .A3(n1013), .ZN(n1110) );
INV_X1 U838 ( .A(n1167), .ZN(n1165) );
NAND2_X1 U839 ( .A1(n1026), .A2(n1168), .ZN(n1158) );
NAND2_X1 U840 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
OR2_X1 U841 ( .A1(n1171), .A2(KEYINPUT19), .ZN(n1170) );
XOR2_X1 U842 ( .A(n1172), .B(KEYINPUT38), .Z(n1169) );
NAND3_X1 U843 ( .A1(KEYINPUT19), .A2(n1173), .A3(n1174), .ZN(n1157) );
INV_X1 U844 ( .A(n1171), .ZN(n1173) );
NOR2_X1 U845 ( .A1(n1057), .A2(G952), .ZN(n1097) );
XNOR2_X1 U846 ( .A(G146), .B(n1148), .ZN(G48) );
NAND3_X1 U847 ( .A1(n1175), .A2(n1013), .A3(n1153), .ZN(n1148) );
XNOR2_X1 U848 ( .A(G143), .B(n1176), .ZN(G45) );
NAND3_X1 U849 ( .A1(n1153), .A2(n1177), .A3(n1178), .ZN(n1176) );
XNOR2_X1 U850 ( .A(n1151), .B(KEYINPUT8), .ZN(n1178) );
XNOR2_X1 U851 ( .A(n1064), .B(n1179), .ZN(G42) );
NOR2_X1 U852 ( .A1(KEYINPUT43), .A2(n1069), .ZN(n1179) );
NAND3_X1 U853 ( .A1(n1180), .A2(n1013), .A3(n1181), .ZN(n1064) );
XNOR2_X1 U854 ( .A(G137), .B(n1147), .ZN(G39) );
NAND3_X1 U855 ( .A1(n1015), .A2(n1031), .A3(n1181), .ZN(n1147) );
NOR3_X1 U856 ( .A1(n1182), .A2(n1030), .A3(n1007), .ZN(n1181) );
INV_X1 U857 ( .A(n1153), .ZN(n1182) );
XOR2_X1 U858 ( .A(n1183), .B(n1184), .Z(G36) );
NOR3_X1 U859 ( .A1(n1007), .A2(KEYINPUT29), .A3(n1185), .ZN(n1184) );
XOR2_X1 U860 ( .A(n1156), .B(KEYINPUT63), .Z(n1185) );
NAND3_X1 U861 ( .A1(n1151), .A2(n1014), .A3(n1153), .ZN(n1156) );
INV_X1 U862 ( .A(n1034), .ZN(n1007) );
XNOR2_X1 U863 ( .A(G134), .B(KEYINPUT0), .ZN(n1183) );
NAND2_X1 U864 ( .A1(n1186), .A2(n1187), .ZN(G33) );
NAND2_X1 U865 ( .A1(G131), .A2(n1150), .ZN(n1187) );
XOR2_X1 U866 ( .A(KEYINPUT20), .B(n1188), .Z(n1186) );
NOR2_X1 U867 ( .A1(G131), .A2(n1150), .ZN(n1188) );
NAND4_X1 U868 ( .A1(n1034), .A2(n1153), .A3(n1013), .A4(n1151), .ZN(n1150) );
NOR2_X1 U869 ( .A1(n1029), .A2(n1051), .ZN(n1034) );
XNOR2_X1 U870 ( .A(G128), .B(n1146), .ZN(G30) );
NAND3_X1 U871 ( .A1(n1175), .A2(n1014), .A3(n1153), .ZN(n1146) );
NOR3_X1 U872 ( .A1(n1008), .A2(n1189), .A3(n1016), .ZN(n1153) );
XOR2_X1 U873 ( .A(G101), .B(n1190), .Z(G3) );
NOR3_X1 U874 ( .A1(n1019), .A2(n1191), .A3(n1167), .ZN(n1190) );
NAND4_X1 U875 ( .A1(n1026), .A2(n1012), .A3(n1192), .A4(n1018), .ZN(n1167) );
XNOR2_X1 U876 ( .A(n1151), .B(KEYINPUT18), .ZN(n1191) );
INV_X1 U877 ( .A(n1015), .ZN(n1019) );
XNOR2_X1 U878 ( .A(G125), .B(n1145), .ZN(G27) );
NAND3_X1 U879 ( .A1(n1193), .A2(n1013), .A3(n1194), .ZN(n1145) );
NOR3_X1 U880 ( .A1(n1012), .A2(n1189), .A3(n1174), .ZN(n1194) );
AND2_X1 U881 ( .A1(n1195), .A2(n1001), .ZN(n1189) );
NAND4_X1 U882 ( .A1(G953), .A2(G902), .A3(n1196), .A4(n1197), .ZN(n1195) );
INV_X1 U883 ( .A(G900), .ZN(n1197) );
NAND2_X1 U884 ( .A1(n1198), .A2(n1199), .ZN(G24) );
NAND2_X1 U885 ( .A1(n1200), .A2(n1092), .ZN(n1199) );
XOR2_X1 U886 ( .A(KEYINPUT31), .B(n1163), .Z(n1200) );
NAND2_X1 U887 ( .A1(n1201), .A2(G122), .ZN(n1198) );
XOR2_X1 U888 ( .A(KEYINPUT10), .B(n1163), .Z(n1201) );
AND3_X1 U889 ( .A1(n1202), .A2(n1164), .A3(n1177), .ZN(n1163) );
INV_X1 U890 ( .A(n1154), .ZN(n1177) );
NAND3_X1 U891 ( .A1(n1026), .A2(n1203), .A3(n1204), .ZN(n1154) );
XNOR2_X1 U892 ( .A(n1035), .B(KEYINPUT49), .ZN(n1204) );
INV_X1 U893 ( .A(n1006), .ZN(n1164) );
NAND2_X1 U894 ( .A1(n1180), .A2(n1030), .ZN(n1006) );
XOR2_X1 U895 ( .A(G119), .B(n1162), .Z(G21) );
AND3_X1 U896 ( .A1(n1175), .A2(n1202), .A3(n1015), .ZN(n1162) );
NOR3_X1 U897 ( .A1(n1030), .A2(n1180), .A3(n1174), .ZN(n1175) );
INV_X1 U898 ( .A(n1031), .ZN(n1180) );
XOR2_X1 U899 ( .A(G116), .B(n1205), .Z(G18) );
NOR2_X1 U900 ( .A1(n1174), .A2(n1172), .ZN(n1205) );
NAND3_X1 U901 ( .A1(n1151), .A2(n1014), .A3(n1202), .ZN(n1172) );
NOR2_X1 U902 ( .A1(n1203), .A2(n1035), .ZN(n1014) );
XOR2_X1 U903 ( .A(G113), .B(n1161), .Z(G15) );
AND4_X1 U904 ( .A1(n1202), .A2(n1013), .A3(n1151), .A4(n1026), .ZN(n1161) );
INV_X1 U905 ( .A(n1033), .ZN(n1151) );
NAND2_X1 U906 ( .A1(n1030), .A2(n1031), .ZN(n1033) );
NOR2_X1 U907 ( .A1(n1206), .A2(n1207), .ZN(n1013) );
AND3_X1 U908 ( .A1(n1192), .A2(n1018), .A3(n1016), .ZN(n1202) );
INV_X1 U909 ( .A(n1012), .ZN(n1016) );
XOR2_X1 U910 ( .A(G110), .B(n1208), .Z(G12) );
NOR2_X1 U911 ( .A1(n1209), .A2(n1171), .ZN(n1208) );
NAND4_X1 U912 ( .A1(n1193), .A2(n1015), .A3(n1012), .A4(n1192), .ZN(n1171) );
NAND2_X1 U913 ( .A1(n1001), .A2(n1210), .ZN(n1192) );
NAND3_X1 U914 ( .A1(G902), .A2(n1196), .A3(n1083), .ZN(n1210) );
NOR2_X1 U915 ( .A1(n1057), .A2(G898), .ZN(n1083) );
NAND3_X1 U916 ( .A1(n1211), .A2(n1196), .A3(G952), .ZN(n1001) );
NAND2_X1 U917 ( .A1(G237), .A2(G234), .ZN(n1196) );
INV_X1 U918 ( .A(n996), .ZN(n1211) );
XOR2_X1 U919 ( .A(G953), .B(KEYINPUT36), .Z(n996) );
XOR2_X1 U920 ( .A(n1044), .B(G469), .Z(n1012) );
INV_X1 U921 ( .A(n1053), .ZN(n1044) );
NAND2_X1 U922 ( .A1(n1212), .A2(n1213), .ZN(n1053) );
XNOR2_X1 U923 ( .A(KEYINPUT37), .B(n1131), .ZN(n1212) );
XOR2_X1 U924 ( .A(n1214), .B(n1215), .Z(n1131) );
XOR2_X1 U925 ( .A(n1216), .B(n1217), .Z(n1215) );
XNOR2_X1 U926 ( .A(n992), .B(G101), .ZN(n1217) );
XNOR2_X1 U927 ( .A(n1069), .B(G110), .ZN(n1216) );
XOR2_X1 U928 ( .A(n1118), .B(n1218), .Z(n1214) );
XOR2_X1 U929 ( .A(n1219), .B(n1220), .Z(n1218) );
NAND2_X1 U930 ( .A1(KEYINPUT34), .A2(G104), .ZN(n1220) );
NAND2_X1 U931 ( .A1(G227), .A2(n1057), .ZN(n1219) );
NOR2_X1 U932 ( .A1(n1203), .A2(n1206), .ZN(n1015) );
INV_X1 U933 ( .A(n1035), .ZN(n1206) );
XNOR2_X1 U934 ( .A(n1221), .B(n1222), .ZN(n1035) );
XOR2_X1 U935 ( .A(KEYINPUT23), .B(G478), .Z(n1222) );
NAND2_X1 U936 ( .A1(n1104), .A2(n1213), .ZN(n1221) );
XNOR2_X1 U937 ( .A(n1223), .B(n1224), .ZN(n1104) );
XOR2_X1 U938 ( .A(n1225), .B(n1226), .Z(n1224) );
XNOR2_X1 U939 ( .A(G107), .B(n1227), .ZN(n1226) );
AND4_X1 U940 ( .A1(n1228), .A2(n1057), .A3(G217), .A4(G234), .ZN(n1227) );
INV_X1 U941 ( .A(KEYINPUT5), .ZN(n1228) );
NAND2_X1 U942 ( .A1(KEYINPUT24), .A2(n1229), .ZN(n1225) );
XNOR2_X1 U943 ( .A(n1092), .B(G116), .ZN(n1229) );
XNOR2_X1 U944 ( .A(G128), .B(n1230), .ZN(n1223) );
XNOR2_X1 U945 ( .A(n1231), .B(G134), .ZN(n1230) );
INV_X1 U946 ( .A(n1207), .ZN(n1203) );
NOR2_X1 U947 ( .A1(n1050), .A2(n1049), .ZN(n1207) );
AND2_X1 U948 ( .A1(G475), .A2(n1232), .ZN(n1049) );
OR2_X1 U949 ( .A1(n1109), .A2(G902), .ZN(n1232) );
NOR3_X1 U950 ( .A1(G475), .A2(G902), .A3(n1109), .ZN(n1050) );
XNOR2_X1 U951 ( .A(n1233), .B(n1234), .ZN(n1109) );
XOR2_X1 U952 ( .A(n1235), .B(n1236), .Z(n1234) );
XNOR2_X1 U953 ( .A(n1237), .B(n1238), .ZN(n1236) );
NOR2_X1 U954 ( .A1(KEYINPUT27), .A2(n1239), .ZN(n1238) );
XNOR2_X1 U955 ( .A(n1240), .B(n1241), .ZN(n1239) );
XNOR2_X1 U956 ( .A(G146), .B(n1069), .ZN(n1241) );
INV_X1 U957 ( .A(G140), .ZN(n1069) );
NAND2_X1 U958 ( .A1(KEYINPUT42), .A2(n1231), .ZN(n1237) );
INV_X1 U959 ( .A(G143), .ZN(n1231) );
XOR2_X1 U960 ( .A(n1242), .B(n1243), .Z(n1233) );
XOR2_X1 U961 ( .A(G104), .B(n1244), .Z(n1243) );
AND3_X1 U962 ( .A1(G214), .A2(n1057), .A3(n1245), .ZN(n1244) );
XNOR2_X1 U963 ( .A(G131), .B(KEYINPUT15), .ZN(n1242) );
NOR3_X1 U964 ( .A1(n1030), .A2(n1008), .A3(n1031), .ZN(n1193) );
XNOR2_X1 U965 ( .A(n1246), .B(G472), .ZN(n1031) );
NAND3_X1 U966 ( .A1(n1247), .A2(n1248), .A3(n1213), .ZN(n1246) );
NAND2_X1 U967 ( .A1(KEYINPUT59), .A2(n1249), .ZN(n1248) );
XOR2_X1 U968 ( .A(n1250), .B(n1116), .Z(n1249) );
NAND2_X1 U969 ( .A1(n1251), .A2(KEYINPUT11), .ZN(n1250) );
NAND3_X1 U970 ( .A1(n1252), .A2(n1251), .A3(n1253), .ZN(n1247) );
INV_X1 U971 ( .A(KEYINPUT59), .ZN(n1253) );
XNOR2_X1 U972 ( .A(n1118), .B(n1254), .ZN(n1251) );
INV_X1 U973 ( .A(n1119), .ZN(n1254) );
XNOR2_X1 U974 ( .A(n1255), .B(n1095), .ZN(n1119) );
NAND2_X1 U975 ( .A1(KEYINPUT57), .A2(G113), .ZN(n1255) );
XOR2_X1 U976 ( .A(n1256), .B(n1257), .Z(n1118) );
XOR2_X1 U977 ( .A(n1258), .B(n1259), .Z(n1257) );
NAND2_X1 U978 ( .A1(KEYINPUT47), .A2(G137), .ZN(n1259) );
NAND2_X1 U979 ( .A1(KEYINPUT48), .A2(n1067), .ZN(n1258) );
INV_X1 U980 ( .A(G131), .ZN(n1067) );
XNOR2_X1 U981 ( .A(n1074), .B(n1136), .ZN(n1256) );
XOR2_X1 U982 ( .A(G134), .B(KEYINPUT33), .Z(n1074) );
XOR2_X1 U983 ( .A(KEYINPUT11), .B(n1116), .Z(n1252) );
XNOR2_X1 U984 ( .A(n1260), .B(G101), .ZN(n1116) );
NAND3_X1 U985 ( .A1(n1245), .A2(n1057), .A3(G210), .ZN(n1260) );
INV_X1 U986 ( .A(n1018), .ZN(n1008) );
NAND2_X1 U987 ( .A1(G221), .A2(n1261), .ZN(n1018) );
XNOR2_X1 U988 ( .A(n1262), .B(n1101), .ZN(n1030) );
NAND2_X1 U989 ( .A1(G217), .A2(n1261), .ZN(n1101) );
NAND2_X1 U990 ( .A1(n1263), .A2(n1213), .ZN(n1261) );
XOR2_X1 U991 ( .A(KEYINPUT60), .B(G234), .Z(n1263) );
OR2_X1 U992 ( .A1(n1100), .A2(G902), .ZN(n1262) );
XNOR2_X1 U993 ( .A(n1264), .B(n1265), .ZN(n1100) );
XNOR2_X1 U994 ( .A(n1266), .B(n1267), .ZN(n1265) );
XOR2_X1 U995 ( .A(n1268), .B(n1269), .Z(n1267) );
AND3_X1 U996 ( .A1(G221), .A2(n1057), .A3(G234), .ZN(n1269) );
NAND3_X1 U997 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1268) );
NAND2_X1 U998 ( .A1(KEYINPUT32), .A2(G125), .ZN(n1272) );
OR3_X1 U999 ( .A1(n1273), .A2(KEYINPUT32), .A3(G140), .ZN(n1271) );
NAND2_X1 U1000 ( .A1(G140), .A2(n1273), .ZN(n1270) );
NAND2_X1 U1001 ( .A1(KEYINPUT55), .A2(n1240), .ZN(n1273) );
INV_X1 U1002 ( .A(G125), .ZN(n1240) );
XOR2_X1 U1003 ( .A(n1274), .B(n1275), .Z(n1264) );
XOR2_X1 U1004 ( .A(KEYINPUT46), .B(G137), .Z(n1275) );
XNOR2_X1 U1005 ( .A(G119), .B(G110), .ZN(n1274) );
XNOR2_X1 U1006 ( .A(n1026), .B(KEYINPUT56), .ZN(n1209) );
INV_X1 U1007 ( .A(n1174), .ZN(n1026) );
NAND2_X1 U1008 ( .A1(n1276), .A2(n1029), .ZN(n1174) );
XOR2_X1 U1009 ( .A(n1045), .B(n1048), .Z(n1029) );
NAND2_X1 U1010 ( .A1(G210), .A2(n1277), .ZN(n1048) );
NAND2_X1 U1011 ( .A1(n1278), .A2(n1213), .ZN(n1045) );
INV_X1 U1012 ( .A(G902), .ZN(n1213) );
XOR2_X1 U1013 ( .A(n1279), .B(n1135), .Z(n1278) );
XOR2_X1 U1014 ( .A(n1280), .B(n1281), .Z(n1135) );
XOR2_X1 U1015 ( .A(n1095), .B(n1282), .Z(n1281) );
XOR2_X1 U1016 ( .A(KEYINPUT35), .B(G110), .Z(n1282) );
XOR2_X1 U1017 ( .A(G116), .B(G119), .Z(n1095) );
XNOR2_X1 U1018 ( .A(n1235), .B(n1089), .ZN(n1280) );
XNOR2_X1 U1019 ( .A(n1283), .B(n1284), .ZN(n1089) );
XNOR2_X1 U1020 ( .A(KEYINPUT50), .B(n992), .ZN(n1284) );
INV_X1 U1021 ( .A(G107), .ZN(n992) );
XNOR2_X1 U1022 ( .A(G101), .B(G104), .ZN(n1283) );
XNOR2_X1 U1023 ( .A(G113), .B(n1092), .ZN(n1235) );
INV_X1 U1024 ( .A(G122), .ZN(n1092) );
NAND2_X1 U1025 ( .A1(n1285), .A2(KEYINPUT6), .ZN(n1279) );
XOR2_X1 U1026 ( .A(n1286), .B(n1136), .Z(n1285) );
XNOR2_X1 U1027 ( .A(n1287), .B(n1266), .ZN(n1136) );
XOR2_X1 U1028 ( .A(G128), .B(G146), .Z(n1266) );
XNOR2_X1 U1029 ( .A(G143), .B(KEYINPUT61), .ZN(n1287) );
XOR2_X1 U1030 ( .A(n1137), .B(n1288), .Z(n1286) );
NOR2_X1 U1031 ( .A1(G125), .A2(KEYINPUT22), .ZN(n1288) );
NAND2_X1 U1032 ( .A1(G224), .A2(n1057), .ZN(n1137) );
INV_X1 U1033 ( .A(G953), .ZN(n1057) );
XNOR2_X1 U1034 ( .A(n1051), .B(KEYINPUT2), .ZN(n1276) );
INV_X1 U1035 ( .A(n1027), .ZN(n1051) );
NAND2_X1 U1036 ( .A1(G214), .A2(n1277), .ZN(n1027) );
NAND2_X1 U1037 ( .A1(n1289), .A2(n1290), .ZN(n1277) );
XNOR2_X1 U1038 ( .A(KEYINPUT53), .B(n1245), .ZN(n1290) );
INV_X1 U1039 ( .A(G237), .ZN(n1245) );
XNOR2_X1 U1040 ( .A(G902), .B(KEYINPUT9), .ZN(n1289) );
endmodule


