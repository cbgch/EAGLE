//Key = 0100000111101001100000011110000011011111111111001010011100110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
n1477, n1478, n1479, n1480;

XOR2_X1 U803 ( .A(G107), .B(n1117), .Z(G9) );
NOR2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(G75) );
NOR3_X1 U805 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
XOR2_X1 U806 ( .A(KEYINPUT27), .B(n1123), .Z(n1122) );
NOR2_X1 U807 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NOR2_X1 U808 ( .A1(n1126), .A2(n1127), .ZN(n1124) );
NOR2_X1 U809 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR2_X1 U810 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
NOR2_X1 U811 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NOR2_X1 U812 ( .A1(n1134), .A2(n1135), .ZN(n1130) );
NOR2_X1 U813 ( .A1(n1136), .A2(n1137), .ZN(n1134) );
NOR2_X1 U814 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR4_X1 U815 ( .A1(n1140), .A2(n1141), .A3(n1135), .A4(n1133), .ZN(n1126) );
INV_X1 U816 ( .A(n1142), .ZN(n1133) );
INV_X1 U817 ( .A(n1143), .ZN(n1121) );
NAND3_X1 U818 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1120) );
NAND2_X1 U819 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U820 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NAND4_X1 U821 ( .A1(n1151), .A2(n1142), .A3(n1152), .A4(n1153), .ZN(n1150) );
NAND2_X1 U822 ( .A1(n1154), .A2(n1155), .ZN(n1149) );
NAND3_X1 U823 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1155) );
NAND2_X1 U824 ( .A1(n1142), .A2(n1159), .ZN(n1158) );
NOR2_X1 U825 ( .A1(n1160), .A2(n1139), .ZN(n1142) );
NAND4_X1 U826 ( .A1(n1161), .A2(n1162), .A3(n1153), .A4(n1163), .ZN(n1157) );
NAND3_X1 U827 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1156) );
XNOR2_X1 U828 ( .A(KEYINPUT51), .B(n1129), .ZN(n1165) );
INV_X1 U829 ( .A(n1125), .ZN(n1147) );
NOR3_X1 U830 ( .A1(n1167), .A2(G953), .A3(G952), .ZN(n1118) );
INV_X1 U831 ( .A(n1144), .ZN(n1167) );
NAND4_X1 U832 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1144) );
NOR4_X1 U833 ( .A1(n1151), .A2(n1172), .A3(n1161), .A4(n1129), .ZN(n1171) );
NOR4_X1 U834 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1170) );
NOR2_X1 U835 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XNOR2_X1 U836 ( .A(n1179), .B(KEYINPUT54), .ZN(n1178) );
NOR2_X1 U837 ( .A1(G475), .A2(n1180), .ZN(n1175) );
XNOR2_X1 U838 ( .A(n1179), .B(KEYINPUT4), .ZN(n1180) );
NOR3_X1 U839 ( .A1(n1181), .A2(KEYINPUT52), .A3(n1182), .ZN(n1174) );
AND2_X1 U840 ( .A1(n1181), .A2(KEYINPUT52), .ZN(n1173) );
XNOR2_X1 U841 ( .A(n1183), .B(n1184), .ZN(n1169) );
NAND2_X1 U842 ( .A1(KEYINPUT53), .A2(G469), .ZN(n1183) );
XNOR2_X1 U843 ( .A(n1185), .B(n1186), .ZN(n1168) );
XOR2_X1 U844 ( .A(n1187), .B(n1188), .Z(G72) );
NOR2_X1 U845 ( .A1(n1189), .A2(n1145), .ZN(n1188) );
AND2_X1 U846 ( .A1(G227), .A2(G900), .ZN(n1189) );
NAND2_X1 U847 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
NAND3_X1 U848 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1191) );
INV_X1 U849 ( .A(n1195), .ZN(n1193) );
OR2_X1 U850 ( .A1(n1192), .A2(n1194), .ZN(n1190) );
XOR2_X1 U851 ( .A(n1196), .B(n1197), .Z(n1194) );
XOR2_X1 U852 ( .A(n1198), .B(n1199), .Z(n1197) );
NAND2_X1 U853 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND2_X1 U854 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
INV_X1 U855 ( .A(KEYINPUT61), .ZN(n1203) );
NAND2_X1 U856 ( .A1(n1204), .A2(n1205), .ZN(n1202) );
NAND2_X1 U857 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U858 ( .A1(KEYINPUT48), .A2(n1208), .ZN(n1204) );
NAND2_X1 U859 ( .A1(KEYINPUT61), .A2(n1209), .ZN(n1200) );
NAND2_X1 U860 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND2_X1 U861 ( .A1(KEYINPUT48), .A2(n1206), .ZN(n1211) );
NAND2_X1 U862 ( .A1(n1212), .A2(n1213), .ZN(n1206) );
NAND2_X1 U863 ( .A1(n1208), .A2(n1207), .ZN(n1210) );
INV_X1 U864 ( .A(KEYINPUT48), .ZN(n1207) );
XNOR2_X1 U865 ( .A(G125), .B(G140), .ZN(n1208) );
XNOR2_X1 U866 ( .A(n1214), .B(G137), .ZN(n1196) );
NAND2_X1 U867 ( .A1(n1145), .A2(n1215), .ZN(n1192) );
NAND2_X1 U868 ( .A1(n1216), .A2(n1217), .ZN(G69) );
NAND2_X1 U869 ( .A1(n1218), .A2(n1145), .ZN(n1217) );
XNOR2_X1 U870 ( .A(n1219), .B(n1220), .ZN(n1218) );
NAND2_X1 U871 ( .A1(n1221), .A2(G953), .ZN(n1216) );
NAND2_X1 U872 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NAND2_X1 U873 ( .A1(n1219), .A2(n1224), .ZN(n1223) );
NAND2_X1 U874 ( .A1(G224), .A2(n1225), .ZN(n1222) );
NAND2_X1 U875 ( .A1(G898), .A2(n1219), .ZN(n1225) );
NAND3_X1 U876 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1219) );
NAND2_X1 U877 ( .A1(G953), .A2(n1229), .ZN(n1228) );
NAND4_X1 U878 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1227) );
OR2_X1 U879 ( .A1(n1234), .A2(KEYINPUT20), .ZN(n1233) );
NAND2_X1 U880 ( .A1(KEYINPUT20), .A2(n1235), .ZN(n1232) );
NAND2_X1 U881 ( .A1(KEYINPUT55), .A2(n1236), .ZN(n1230) );
NAND3_X1 U882 ( .A1(n1236), .A2(n1237), .A3(KEYINPUT55), .ZN(n1226) );
NAND3_X1 U883 ( .A1(n1238), .A2(n1239), .A3(n1234), .ZN(n1237) );
OR2_X1 U884 ( .A1(n1231), .A2(KEYINPUT20), .ZN(n1239) );
NAND2_X1 U885 ( .A1(KEYINPUT20), .A2(n1240), .ZN(n1238) );
NOR2_X1 U886 ( .A1(n1241), .A2(n1242), .ZN(G66) );
NOR2_X1 U887 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XOR2_X1 U888 ( .A(KEYINPUT56), .B(n1245), .Z(n1244) );
NOR2_X1 U889 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
AND2_X1 U890 ( .A1(n1247), .A2(n1246), .ZN(n1243) );
XOR2_X1 U891 ( .A(n1248), .B(KEYINPUT46), .Z(n1246) );
NAND2_X1 U892 ( .A1(n1249), .A2(n1250), .ZN(n1247) );
NOR2_X1 U893 ( .A1(n1241), .A2(n1251), .ZN(G63) );
XOR2_X1 U894 ( .A(n1252), .B(n1253), .Z(n1251) );
NOR2_X1 U895 ( .A1(n1181), .A2(n1254), .ZN(n1252) );
NOR2_X1 U896 ( .A1(n1241), .A2(n1255), .ZN(G60) );
NOR3_X1 U897 ( .A1(n1179), .A2(n1256), .A3(n1257), .ZN(n1255) );
AND3_X1 U898 ( .A1(n1258), .A2(G475), .A3(n1249), .ZN(n1257) );
NOR2_X1 U899 ( .A1(n1259), .A2(n1258), .ZN(n1256) );
NOR2_X1 U900 ( .A1(n1143), .A2(n1177), .ZN(n1259) );
XOR2_X1 U901 ( .A(n1260), .B(n1261), .Z(G6) );
NOR2_X1 U902 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XNOR2_X1 U903 ( .A(KEYINPUT59), .B(KEYINPUT31), .ZN(n1262) );
NOR2_X1 U904 ( .A1(n1241), .A2(n1264), .ZN(G57) );
XOR2_X1 U905 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U906 ( .A(n1267), .B(n1268), .Z(n1266) );
AND2_X1 U907 ( .A1(G472), .A2(n1249), .ZN(n1268) );
NOR2_X1 U908 ( .A1(n1269), .A2(n1270), .ZN(n1267) );
XOR2_X1 U909 ( .A(n1271), .B(n1272), .Z(n1265) );
NOR2_X1 U910 ( .A1(KEYINPUT5), .A2(n1273), .ZN(n1272) );
NOR2_X1 U911 ( .A1(n1241), .A2(n1274), .ZN(G54) );
XOR2_X1 U912 ( .A(n1275), .B(n1276), .Z(n1274) );
NOR2_X1 U913 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NOR2_X1 U914 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NOR2_X1 U915 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
INV_X1 U916 ( .A(KEYINPUT9), .ZN(n1282) );
NOR2_X1 U917 ( .A1(n1283), .A2(n1284), .ZN(n1281) );
XOR2_X1 U918 ( .A(n1285), .B(KEYINPUT42), .Z(n1284) );
INV_X1 U919 ( .A(n1286), .ZN(n1283) );
AND2_X1 U920 ( .A1(KEYINPUT9), .A2(n1279), .ZN(n1277) );
NOR2_X1 U921 ( .A1(n1286), .A2(n1285), .ZN(n1279) );
XOR2_X1 U922 ( .A(G140), .B(n1287), .Z(n1286) );
NOR2_X1 U923 ( .A1(KEYINPUT62), .A2(n1288), .ZN(n1287) );
XOR2_X1 U924 ( .A(n1289), .B(n1290), .Z(n1275) );
AND2_X1 U925 ( .A1(G469), .A2(n1249), .ZN(n1290) );
NOR3_X1 U926 ( .A1(n1291), .A2(n1241), .A3(n1292), .ZN(G51) );
NOR3_X1 U927 ( .A1(n1293), .A2(KEYINPUT34), .A3(n1294), .ZN(n1292) );
XOR2_X1 U928 ( .A(n1295), .B(n1296), .Z(n1294) );
AND2_X1 U929 ( .A1(n1297), .A2(KEYINPUT37), .ZN(n1296) );
NOR2_X1 U930 ( .A1(n1145), .A2(G952), .ZN(n1241) );
NOR2_X1 U931 ( .A1(n1298), .A2(n1299), .ZN(n1291) );
XOR2_X1 U932 ( .A(n1295), .B(n1300), .Z(n1299) );
NOR2_X1 U933 ( .A1(n1297), .A2(n1301), .ZN(n1300) );
INV_X1 U934 ( .A(KEYINPUT37), .ZN(n1301) );
NAND3_X1 U935 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1295) );
INV_X1 U936 ( .A(n1186), .ZN(n1304) );
NAND2_X1 U937 ( .A1(KEYINPUT1), .A2(n1254), .ZN(n1303) );
INV_X1 U938 ( .A(n1249), .ZN(n1254) );
NOR2_X1 U939 ( .A1(n1305), .A2(n1143), .ZN(n1249) );
NAND2_X1 U940 ( .A1(n1306), .A2(n1307), .ZN(n1302) );
INV_X1 U941 ( .A(KEYINPUT1), .ZN(n1307) );
NAND2_X1 U942 ( .A1(n1143), .A2(G902), .ZN(n1306) );
NOR2_X1 U943 ( .A1(n1220), .A2(n1215), .ZN(n1143) );
NAND4_X1 U944 ( .A1(n1308), .A2(n1309), .A3(n1310), .A4(n1311), .ZN(n1215) );
NOR3_X1 U945 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(n1311) );
INV_X1 U946 ( .A(n1315), .ZN(n1312) );
NAND2_X1 U947 ( .A1(n1166), .A2(n1316), .ZN(n1310) );
NAND2_X1 U948 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND2_X1 U949 ( .A1(n1319), .A2(n1320), .ZN(n1317) );
NAND2_X1 U950 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NAND4_X1 U951 ( .A1(n1323), .A2(n1324), .A3(n1325), .A4(n1326), .ZN(n1220) );
NOR4_X1 U952 ( .A1(n1117), .A2(n1260), .A3(n1327), .A4(n1328), .ZN(n1326) );
NOR2_X1 U953 ( .A1(n1138), .A2(n1329), .ZN(n1328) );
NOR3_X1 U954 ( .A1(n1330), .A2(n1331), .A3(n1139), .ZN(n1327) );
AND2_X1 U955 ( .A1(n1332), .A2(n1333), .ZN(n1260) );
AND2_X1 U956 ( .A1(n1164), .A2(n1333), .ZN(n1117) );
AND3_X1 U957 ( .A1(n1334), .A2(n1153), .A3(n1335), .ZN(n1333) );
NOR2_X1 U958 ( .A1(n1336), .A2(n1337), .ZN(n1325) );
NOR2_X1 U959 ( .A1(KEYINPUT34), .A2(n1293), .ZN(n1298) );
XNOR2_X1 U960 ( .A(n1338), .B(n1339), .ZN(n1293) );
XNOR2_X1 U961 ( .A(n1340), .B(n1341), .ZN(n1338) );
NOR2_X1 U962 ( .A1(G125), .A2(KEYINPUT47), .ZN(n1341) );
XNOR2_X1 U963 ( .A(G146), .B(n1308), .ZN(G48) );
NAND3_X1 U964 ( .A1(n1332), .A2(n1342), .A3(n1343), .ZN(n1308) );
XNOR2_X1 U965 ( .A(n1309), .B(n1344), .ZN(G45) );
NOR2_X1 U966 ( .A1(KEYINPUT3), .A2(n1345), .ZN(n1344) );
INV_X1 U967 ( .A(G143), .ZN(n1345) );
NAND4_X1 U968 ( .A1(n1319), .A2(n1342), .A3(n1346), .A4(n1347), .ZN(n1309) );
NAND2_X1 U969 ( .A1(n1348), .A2(n1349), .ZN(G42) );
NAND2_X1 U970 ( .A1(n1314), .A2(n1350), .ZN(n1349) );
XOR2_X1 U971 ( .A(KEYINPUT50), .B(n1351), .Z(n1348) );
NOR2_X1 U972 ( .A1(n1314), .A2(n1350), .ZN(n1351) );
AND4_X1 U973 ( .A1(n1159), .A2(n1352), .A3(n1334), .A4(n1136), .ZN(n1314) );
NOR2_X1 U974 ( .A1(n1321), .A2(n1160), .ZN(n1136) );
XNOR2_X1 U975 ( .A(G137), .B(n1353), .ZN(G39) );
NAND2_X1 U976 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
XNOR2_X1 U977 ( .A(KEYINPUT29), .B(n1160), .ZN(n1355) );
INV_X1 U978 ( .A(n1318), .ZN(n1354) );
NAND2_X1 U979 ( .A1(n1343), .A2(n1162), .ZN(n1318) );
XOR2_X1 U980 ( .A(G134), .B(n1356), .Z(G36) );
NOR3_X1 U981 ( .A1(n1160), .A2(KEYINPUT11), .A3(n1357), .ZN(n1356) );
XOR2_X1 U982 ( .A(n1358), .B(KEYINPUT2), .Z(n1357) );
NAND2_X1 U983 ( .A1(n1319), .A2(n1164), .ZN(n1358) );
INV_X1 U984 ( .A(n1359), .ZN(n1319) );
XOR2_X1 U985 ( .A(n1360), .B(n1361), .Z(G33) );
NOR3_X1 U986 ( .A1(n1359), .A2(n1362), .A3(n1321), .ZN(n1361) );
XNOR2_X1 U987 ( .A(n1166), .B(KEYINPUT57), .ZN(n1362) );
INV_X1 U988 ( .A(n1160), .ZN(n1166) );
NAND2_X1 U989 ( .A1(n1163), .A2(n1363), .ZN(n1160) );
NAND2_X1 U990 ( .A1(n1364), .A2(n1352), .ZN(n1359) );
NAND2_X1 U991 ( .A1(KEYINPUT26), .A2(n1365), .ZN(n1360) );
INV_X1 U992 ( .A(G131), .ZN(n1365) );
XNOR2_X1 U993 ( .A(n1366), .B(n1313), .ZN(G30) );
AND3_X1 U994 ( .A1(n1164), .A2(n1342), .A3(n1343), .ZN(n1313) );
AND4_X1 U995 ( .A1(n1334), .A2(n1141), .A3(n1367), .A4(n1352), .ZN(n1343) );
XNOR2_X1 U996 ( .A(G101), .B(n1368), .ZN(G3) );
NAND2_X1 U997 ( .A1(n1369), .A2(n1342), .ZN(n1368) );
XOR2_X1 U998 ( .A(n1329), .B(KEYINPUT8), .Z(n1369) );
NAND3_X1 U999 ( .A1(n1162), .A2(n1370), .A3(n1364), .ZN(n1329) );
NOR3_X1 U1000 ( .A1(n1141), .A2(n1140), .A3(n1132), .ZN(n1364) );
INV_X1 U1001 ( .A(n1334), .ZN(n1132) );
XNOR2_X1 U1002 ( .A(G125), .B(n1315), .ZN(G27) );
NAND4_X1 U1003 ( .A1(n1159), .A2(n1352), .A3(n1342), .A4(n1371), .ZN(n1315) );
NOR2_X1 U1004 ( .A1(n1135), .A2(n1321), .ZN(n1371) );
NAND2_X1 U1005 ( .A1(n1125), .A2(n1372), .ZN(n1352) );
NAND3_X1 U1006 ( .A1(G902), .A2(n1373), .A3(n1195), .ZN(n1372) );
NOR2_X1 U1007 ( .A1(n1145), .A2(G900), .ZN(n1195) );
XNOR2_X1 U1008 ( .A(KEYINPUT36), .B(n1374), .ZN(n1373) );
XOR2_X1 U1009 ( .A(n1375), .B(n1337), .Z(G24) );
AND3_X1 U1010 ( .A1(n1154), .A2(n1335), .A3(n1376), .ZN(n1337) );
NOR3_X1 U1011 ( .A1(n1129), .A2(n1377), .A3(n1378), .ZN(n1376) );
NAND2_X1 U1012 ( .A1(KEYINPUT10), .A2(n1379), .ZN(n1375) );
XNOR2_X1 U1013 ( .A(G119), .B(n1380), .ZN(G21) );
NAND4_X1 U1014 ( .A1(KEYINPUT38), .A2(n1154), .A3(n1381), .A4(n1382), .ZN(n1380) );
NOR4_X1 U1015 ( .A1(n1383), .A2(n1140), .A3(n1331), .A4(n1139), .ZN(n1382) );
INV_X1 U1016 ( .A(n1162), .ZN(n1139) );
INV_X1 U1017 ( .A(n1141), .ZN(n1331) );
XNOR2_X1 U1018 ( .A(n1342), .B(KEYINPUT16), .ZN(n1381) );
XOR2_X1 U1019 ( .A(G116), .B(n1336), .Z(G18) );
NOR3_X1 U1020 ( .A1(n1141), .A2(n1322), .A3(n1330), .ZN(n1336) );
INV_X1 U1021 ( .A(n1164), .ZN(n1322) );
NOR2_X1 U1022 ( .A1(n1346), .A2(n1377), .ZN(n1164) );
XNOR2_X1 U1023 ( .A(G113), .B(n1323), .ZN(G15) );
OR3_X1 U1024 ( .A1(n1141), .A2(n1321), .A3(n1330), .ZN(n1323) );
NAND3_X1 U1025 ( .A1(n1335), .A2(n1367), .A3(n1154), .ZN(n1330) );
INV_X1 U1026 ( .A(n1135), .ZN(n1154) );
NAND2_X1 U1027 ( .A1(n1384), .A2(n1385), .ZN(n1135) );
XNOR2_X1 U1028 ( .A(KEYINPUT39), .B(n1152), .ZN(n1384) );
INV_X1 U1029 ( .A(n1332), .ZN(n1321) );
NOR2_X1 U1030 ( .A1(n1347), .A2(n1378), .ZN(n1332) );
XOR2_X1 U1031 ( .A(n1324), .B(n1386), .Z(G12) );
NOR2_X1 U1032 ( .A1(G110), .A2(KEYINPUT19), .ZN(n1386) );
NAND4_X1 U1033 ( .A1(n1162), .A2(n1335), .A3(n1334), .A4(n1159), .ZN(n1324) );
NAND2_X1 U1034 ( .A1(n1387), .A2(n1388), .ZN(n1159) );
OR2_X1 U1035 ( .A1(n1129), .A2(KEYINPUT23), .ZN(n1388) );
INV_X1 U1036 ( .A(n1153), .ZN(n1129) );
NOR2_X1 U1037 ( .A1(n1367), .A2(n1141), .ZN(n1153) );
NAND3_X1 U1038 ( .A1(n1141), .A2(n1140), .A3(KEYINPUT23), .ZN(n1387) );
INV_X1 U1039 ( .A(n1367), .ZN(n1140) );
XNOR2_X1 U1040 ( .A(n1389), .B(G472), .ZN(n1367) );
NAND2_X1 U1041 ( .A1(n1305), .A2(n1390), .ZN(n1389) );
NAND2_X1 U1042 ( .A1(n1391), .A2(n1392), .ZN(n1390) );
NAND2_X1 U1043 ( .A1(n1393), .A2(n1394), .ZN(n1392) );
XOR2_X1 U1044 ( .A(n1395), .B(n1396), .Z(n1391) );
NOR2_X1 U1045 ( .A1(n1269), .A2(n1397), .ZN(n1396) );
XNOR2_X1 U1046 ( .A(n1270), .B(KEYINPUT43), .ZN(n1397) );
AND2_X1 U1047 ( .A1(n1398), .A2(G101), .ZN(n1270) );
NOR2_X1 U1048 ( .A1(G101), .A2(n1398), .ZN(n1269) );
AND3_X1 U1049 ( .A1(n1399), .A2(n1145), .A3(G210), .ZN(n1398) );
OR2_X1 U1050 ( .A1(n1394), .A2(n1393), .ZN(n1395) );
XNOR2_X1 U1051 ( .A(n1271), .B(n1273), .ZN(n1393) );
XNOR2_X1 U1052 ( .A(n1400), .B(n1401), .ZN(n1273) );
XNOR2_X1 U1053 ( .A(n1402), .B(n1403), .ZN(n1271) );
INV_X1 U1054 ( .A(n1404), .ZN(n1403) );
NAND2_X1 U1055 ( .A1(KEYINPUT40), .A2(n1405), .ZN(n1402) );
INV_X1 U1056 ( .A(KEYINPUT41), .ZN(n1394) );
XNOR2_X1 U1057 ( .A(n1406), .B(n1250), .ZN(n1141) );
AND2_X1 U1058 ( .A1(G217), .A2(n1407), .ZN(n1250) );
NAND2_X1 U1059 ( .A1(n1248), .A2(n1305), .ZN(n1406) );
XNOR2_X1 U1060 ( .A(n1408), .B(n1409), .ZN(n1248) );
XOR2_X1 U1061 ( .A(G137), .B(n1410), .Z(n1409) );
NOR2_X1 U1062 ( .A1(KEYINPUT0), .A2(n1411), .ZN(n1410) );
XOR2_X1 U1063 ( .A(n1412), .B(n1413), .Z(n1411) );
XNOR2_X1 U1064 ( .A(n1288), .B(n1414), .ZN(n1413) );
XNOR2_X1 U1065 ( .A(n1366), .B(G119), .ZN(n1414) );
XNOR2_X1 U1066 ( .A(n1415), .B(n1416), .ZN(n1412) );
NAND2_X1 U1067 ( .A1(n1417), .A2(n1213), .ZN(n1415) );
XNOR2_X1 U1068 ( .A(KEYINPUT35), .B(n1212), .ZN(n1417) );
NAND2_X1 U1069 ( .A1(G221), .A2(n1418), .ZN(n1408) );
NOR2_X1 U1070 ( .A1(n1152), .A2(n1151), .ZN(n1334) );
INV_X1 U1071 ( .A(n1385), .ZN(n1151) );
NAND2_X1 U1072 ( .A1(G221), .A2(n1407), .ZN(n1385) );
NAND2_X1 U1073 ( .A1(G234), .A2(n1419), .ZN(n1407) );
XNOR2_X1 U1074 ( .A(KEYINPUT33), .B(n1305), .ZN(n1419) );
XOR2_X1 U1075 ( .A(n1184), .B(G469), .Z(n1152) );
NAND2_X1 U1076 ( .A1(n1420), .A2(n1305), .ZN(n1184) );
XOR2_X1 U1077 ( .A(n1421), .B(n1422), .Z(n1420) );
XNOR2_X1 U1078 ( .A(n1288), .B(n1423), .ZN(n1422) );
XNOR2_X1 U1079 ( .A(KEYINPUT6), .B(n1350), .ZN(n1423) );
INV_X1 U1080 ( .A(G110), .ZN(n1288) );
XNOR2_X1 U1081 ( .A(n1289), .B(n1285), .ZN(n1421) );
NAND2_X1 U1082 ( .A1(G227), .A2(n1145), .ZN(n1285) );
XOR2_X1 U1083 ( .A(n1424), .B(n1425), .Z(n1289) );
XNOR2_X1 U1084 ( .A(n1366), .B(n1426), .ZN(n1425) );
NOR2_X1 U1085 ( .A1(KEYINPUT13), .A2(n1427), .ZN(n1426) );
XNOR2_X1 U1086 ( .A(n1401), .B(n1428), .ZN(n1424) );
XOR2_X1 U1087 ( .A(n1429), .B(n1430), .Z(n1401) );
INV_X1 U1088 ( .A(n1214), .ZN(n1430) );
XOR2_X1 U1089 ( .A(G131), .B(n1431), .Z(n1214) );
XOR2_X1 U1090 ( .A(n1432), .B(KEYINPUT21), .Z(n1429) );
NAND2_X1 U1091 ( .A1(KEYINPUT44), .A2(n1433), .ZN(n1432) );
XOR2_X1 U1092 ( .A(G137), .B(n1434), .Z(n1433) );
NOR2_X1 U1093 ( .A1(G134), .A2(KEYINPUT18), .ZN(n1434) );
NOR2_X1 U1094 ( .A1(n1138), .A2(n1383), .ZN(n1335) );
INV_X1 U1095 ( .A(n1370), .ZN(n1383) );
NAND2_X1 U1096 ( .A1(n1435), .A2(n1125), .ZN(n1370) );
NAND3_X1 U1097 ( .A1(n1374), .A2(n1145), .A3(G952), .ZN(n1125) );
NAND4_X1 U1098 ( .A1(G953), .A2(G902), .A3(n1374), .A4(n1229), .ZN(n1435) );
INV_X1 U1099 ( .A(G898), .ZN(n1229) );
NAND2_X1 U1100 ( .A1(G234), .A2(n1436), .ZN(n1374) );
XNOR2_X1 U1101 ( .A(KEYINPUT28), .B(n1399), .ZN(n1436) );
INV_X1 U1102 ( .A(n1342), .ZN(n1138) );
NOR2_X1 U1103 ( .A1(n1163), .A2(n1161), .ZN(n1342) );
INV_X1 U1104 ( .A(n1363), .ZN(n1161) );
NAND2_X1 U1105 ( .A1(G214), .A2(n1437), .ZN(n1363) );
XOR2_X1 U1106 ( .A(n1438), .B(n1185), .Z(n1163) );
NAND2_X1 U1107 ( .A1(n1439), .A2(n1305), .ZN(n1185) );
XNOR2_X1 U1108 ( .A(n1440), .B(n1297), .ZN(n1439) );
NAND2_X1 U1109 ( .A1(n1441), .A2(n1442), .ZN(n1297) );
NAND2_X1 U1110 ( .A1(n1236), .A2(n1443), .ZN(n1442) );
NAND2_X1 U1111 ( .A1(n1234), .A2(n1231), .ZN(n1443) );
OR2_X1 U1112 ( .A1(n1444), .A2(n1240), .ZN(n1231) );
NAND2_X1 U1113 ( .A1(n1240), .A2(n1444), .ZN(n1234) );
INV_X1 U1114 ( .A(n1235), .ZN(n1240) );
INV_X1 U1115 ( .A(n1445), .ZN(n1236) );
NAND2_X1 U1116 ( .A1(n1445), .A2(n1446), .ZN(n1441) );
XNOR2_X1 U1117 ( .A(n1444), .B(n1235), .ZN(n1446) );
XOR2_X1 U1118 ( .A(G110), .B(n1447), .Z(n1235) );
XNOR2_X1 U1119 ( .A(n1404), .B(n1405), .ZN(n1444) );
INV_X1 U1120 ( .A(G119), .ZN(n1405) );
XOR2_X1 U1121 ( .A(G113), .B(n1448), .Z(n1404) );
XNOR2_X1 U1122 ( .A(n1449), .B(n1428), .ZN(n1445) );
XOR2_X1 U1123 ( .A(G101), .B(KEYINPUT24), .Z(n1428) );
NAND2_X1 U1124 ( .A1(KEYINPUT32), .A2(n1450), .ZN(n1449) );
XNOR2_X1 U1125 ( .A(KEYINPUT49), .B(n1427), .ZN(n1450) );
XOR2_X1 U1126 ( .A(n1263), .B(G107), .Z(n1427) );
NOR3_X1 U1127 ( .A1(n1451), .A2(KEYINPUT14), .A3(n1452), .ZN(n1440) );
NOR2_X1 U1128 ( .A1(n1340), .A2(n1453), .ZN(n1452) );
XOR2_X1 U1129 ( .A(n1454), .B(n1339), .Z(n1453) );
XOR2_X1 U1130 ( .A(KEYINPUT60), .B(n1455), .Z(n1451) );
NOR2_X1 U1131 ( .A1(n1456), .A2(n1457), .ZN(n1455) );
INV_X1 U1132 ( .A(n1340), .ZN(n1457) );
NOR2_X1 U1133 ( .A1(n1224), .A2(G953), .ZN(n1340) );
INV_X1 U1134 ( .A(G224), .ZN(n1224) );
XNOR2_X1 U1135 ( .A(n1339), .B(n1454), .ZN(n1456) );
AND2_X1 U1136 ( .A1(KEYINPUT58), .A2(n1458), .ZN(n1454) );
XNOR2_X1 U1137 ( .A(n1400), .B(n1431), .ZN(n1339) );
XNOR2_X1 U1138 ( .A(G143), .B(n1416), .ZN(n1431) );
NAND2_X1 U1139 ( .A1(KEYINPUT12), .A2(n1366), .ZN(n1400) );
INV_X1 U1140 ( .A(G128), .ZN(n1366) );
NAND2_X1 U1141 ( .A1(KEYINPUT45), .A2(n1186), .ZN(n1438) );
NAND2_X1 U1142 ( .A1(G210), .A2(n1437), .ZN(n1186) );
NAND2_X1 U1143 ( .A1(n1399), .A2(n1305), .ZN(n1437) );
INV_X1 U1144 ( .A(G902), .ZN(n1305) );
NOR2_X1 U1145 ( .A1(n1347), .A2(n1346), .ZN(n1162) );
INV_X1 U1146 ( .A(n1378), .ZN(n1346) );
XOR2_X1 U1147 ( .A(n1179), .B(n1177), .Z(n1378) );
INV_X1 U1148 ( .A(G475), .ZN(n1177) );
NOR2_X1 U1149 ( .A1(n1258), .A2(G902), .ZN(n1179) );
XOR2_X1 U1150 ( .A(n1459), .B(n1460), .Z(n1258) );
XOR2_X1 U1151 ( .A(n1461), .B(n1462), .Z(n1460) );
XNOR2_X1 U1152 ( .A(G113), .B(n1263), .ZN(n1462) );
INV_X1 U1153 ( .A(G104), .ZN(n1263) );
NOR2_X1 U1154 ( .A1(KEYINPUT63), .A2(n1463), .ZN(n1461) );
XOR2_X1 U1155 ( .A(n1464), .B(n1465), .Z(n1463) );
AND3_X1 U1156 ( .A1(G214), .A2(n1145), .A3(n1399), .ZN(n1465) );
INV_X1 U1157 ( .A(G237), .ZN(n1399) );
XNOR2_X1 U1158 ( .A(G131), .B(G143), .ZN(n1464) );
XOR2_X1 U1159 ( .A(n1466), .B(n1447), .Z(n1459) );
NAND3_X1 U1160 ( .A1(n1467), .A2(n1468), .A3(n1469), .ZN(n1466) );
NAND2_X1 U1161 ( .A1(KEYINPUT22), .A2(n1470), .ZN(n1469) );
OR3_X1 U1162 ( .A1(n1470), .A2(KEYINPUT22), .A3(n1416), .ZN(n1468) );
NAND2_X1 U1163 ( .A1(n1416), .A2(n1471), .ZN(n1467) );
NAND2_X1 U1164 ( .A1(n1472), .A2(n1473), .ZN(n1471) );
INV_X1 U1165 ( .A(KEYINPUT22), .ZN(n1473) );
XNOR2_X1 U1166 ( .A(KEYINPUT17), .B(n1470), .ZN(n1472) );
NAND2_X1 U1167 ( .A1(n1474), .A2(n1213), .ZN(n1470) );
NAND2_X1 U1168 ( .A1(G125), .A2(n1350), .ZN(n1213) );
INV_X1 U1169 ( .A(G140), .ZN(n1350) );
XNOR2_X1 U1170 ( .A(KEYINPUT25), .B(n1212), .ZN(n1474) );
NAND2_X1 U1171 ( .A1(G140), .A2(n1458), .ZN(n1212) );
INV_X1 U1172 ( .A(G125), .ZN(n1458) );
XNOR2_X1 U1173 ( .A(G146), .B(KEYINPUT15), .ZN(n1416) );
INV_X1 U1174 ( .A(n1377), .ZN(n1347) );
NOR2_X1 U1175 ( .A1(n1172), .A2(n1475), .ZN(n1377) );
NOR2_X1 U1176 ( .A1(n1181), .A2(n1182), .ZN(n1475) );
AND2_X1 U1177 ( .A1(n1182), .A2(n1181), .ZN(n1172) );
INV_X1 U1178 ( .A(G478), .ZN(n1181) );
NOR2_X1 U1179 ( .A1(n1253), .A2(G902), .ZN(n1182) );
XNOR2_X1 U1180 ( .A(n1476), .B(n1477), .ZN(n1253) );
XOR2_X1 U1181 ( .A(n1478), .B(n1479), .Z(n1477) );
XNOR2_X1 U1182 ( .A(G107), .B(G143), .ZN(n1479) );
NAND2_X1 U1183 ( .A1(G217), .A2(n1418), .ZN(n1478) );
AND2_X1 U1184 ( .A1(G234), .A2(n1145), .ZN(n1418) );
INV_X1 U1185 ( .A(G953), .ZN(n1145) );
XOR2_X1 U1186 ( .A(n1198), .B(n1480), .Z(n1476) );
XOR2_X1 U1187 ( .A(n1448), .B(n1447), .Z(n1480) );
XNOR2_X1 U1188 ( .A(n1379), .B(KEYINPUT30), .ZN(n1447) );
INV_X1 U1189 ( .A(G122), .ZN(n1379) );
XOR2_X1 U1190 ( .A(G116), .B(KEYINPUT7), .Z(n1448) );
XNOR2_X1 U1191 ( .A(G134), .B(G128), .ZN(n1198) );
endmodule


