//Key = 0011101110010111101101010011001001101011000100110100001111011111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360;

XNOR2_X1 U738 ( .A(G107), .B(n1029), .ZN(G9) );
NOR2_X1 U739 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U740 ( .A1(G953), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1031) );
NOR2_X1 U741 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U742 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR3_X1 U743 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NOR2_X1 U744 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR3_X1 U745 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NOR3_X1 U746 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NOR2_X1 U747 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U748 ( .A1(n1052), .A2(n1053), .ZN(n1045) );
AND2_X1 U749 ( .A1(n1054), .A2(n1052), .ZN(n1042) );
NOR4_X1 U750 ( .A1(n1047), .A2(n1055), .A3(n1056), .A4(n1044), .ZN(n1037) );
INV_X1 U751 ( .A(n1052), .ZN(n1056) );
NOR2_X1 U752 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U753 ( .A1(n1059), .A2(n1039), .ZN(n1058) );
NOR2_X1 U754 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U755 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
XNOR2_X1 U756 ( .A(n1064), .B(KEYINPUT50), .ZN(n1062) );
NOR2_X1 U757 ( .A1(n1065), .A2(n1041), .ZN(n1057) );
INV_X1 U758 ( .A(n1066), .ZN(n1041) );
NOR2_X1 U759 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR3_X1 U760 ( .A1(n1032), .A2(G953), .A3(G952), .ZN(n1030) );
AND4_X1 U761 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1032) );
NOR4_X1 U762 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1072) );
XOR2_X1 U763 ( .A(n1077), .B(G472), .Z(n1075) );
NAND2_X1 U764 ( .A1(KEYINPUT60), .A2(n1078), .ZN(n1077) );
XOR2_X1 U765 ( .A(n1079), .B(n1080), .Z(n1074) );
NOR2_X1 U766 ( .A1(G475), .A2(KEYINPUT0), .ZN(n1080) );
XNOR2_X1 U767 ( .A(n1081), .B(n1082), .ZN(n1073) );
NAND2_X1 U768 ( .A1(KEYINPUT6), .A2(n1083), .ZN(n1081) );
NOR3_X1 U769 ( .A1(n1047), .A2(n1084), .A3(n1085), .ZN(n1071) );
NAND2_X1 U770 ( .A1(n1086), .A2(n1087), .ZN(n1070) );
XOR2_X1 U771 ( .A(n1088), .B(n1089), .Z(n1069) );
NAND2_X1 U772 ( .A1(KEYINPUT13), .A2(n1090), .ZN(n1089) );
XOR2_X1 U773 ( .A(n1091), .B(n1092), .Z(G72) );
NAND2_X1 U774 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND4_X1 U775 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1094) );
XOR2_X1 U776 ( .A(n1099), .B(KEYINPUT28), .Z(n1095) );
NAND3_X1 U777 ( .A1(G900), .A2(G227), .A3(G953), .ZN(n1093) );
NAND2_X1 U778 ( .A1(n1100), .A2(n1101), .ZN(n1091) );
NAND2_X1 U779 ( .A1(G953), .A2(n1102), .ZN(n1101) );
XOR2_X1 U780 ( .A(n1103), .B(n1104), .Z(n1100) );
XOR2_X1 U781 ( .A(n1105), .B(n1106), .Z(n1103) );
NAND3_X1 U782 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1105) );
OR2_X1 U783 ( .A1(n1110), .A2(KEYINPUT26), .ZN(n1109) );
NAND3_X1 U784 ( .A1(KEYINPUT26), .A2(n1110), .A3(n1111), .ZN(n1108) );
INV_X1 U785 ( .A(G131), .ZN(n1111) );
NAND2_X1 U786 ( .A1(G131), .A2(n1112), .ZN(n1107) );
NAND2_X1 U787 ( .A1(n1113), .A2(KEYINPUT26), .ZN(n1112) );
XOR2_X1 U788 ( .A(n1110), .B(KEYINPUT22), .Z(n1113) );
NAND2_X1 U789 ( .A1(n1114), .A2(n1115), .ZN(G69) );
NAND2_X1 U790 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U791 ( .A1(n1118), .A2(n1119), .ZN(n1114) );
INV_X1 U792 ( .A(n1116), .ZN(n1119) );
NOR2_X1 U793 ( .A1(KEYINPUT10), .A2(n1120), .ZN(n1116) );
XOR2_X1 U794 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U795 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U796 ( .A(n1125), .B(n1126), .Z(n1124) );
XNOR2_X1 U797 ( .A(n1127), .B(KEYINPUT37), .ZN(n1126) );
NAND2_X1 U798 ( .A1(KEYINPUT21), .A2(n1128), .ZN(n1127) );
XNOR2_X1 U799 ( .A(n1129), .B(n1130), .ZN(n1125) );
NAND2_X1 U800 ( .A1(n1098), .A2(n1131), .ZN(n1121) );
NAND2_X1 U801 ( .A1(n1132), .A2(n1117), .ZN(n1118) );
NAND2_X1 U802 ( .A1(G953), .A2(n1133), .ZN(n1117) );
INV_X1 U803 ( .A(G224), .ZN(n1133) );
INV_X1 U804 ( .A(n1123), .ZN(n1132) );
NOR2_X1 U805 ( .A1(n1098), .A2(G898), .ZN(n1123) );
NOR2_X1 U806 ( .A1(n1134), .A2(n1135), .ZN(G66) );
XNOR2_X1 U807 ( .A(n1136), .B(n1137), .ZN(n1135) );
NOR2_X1 U808 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR2_X1 U809 ( .A1(n1134), .A2(n1140), .ZN(G63) );
XOR2_X1 U810 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U811 ( .A1(n1143), .A2(G478), .ZN(n1142) );
NOR3_X1 U812 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(G60) );
NOR3_X1 U813 ( .A1(n1147), .A2(G953), .A3(G952), .ZN(n1146) );
AND2_X1 U814 ( .A1(n1147), .A2(n1134), .ZN(n1145) );
INV_X1 U815 ( .A(KEYINPUT31), .ZN(n1147) );
NOR2_X1 U816 ( .A1(n1148), .A2(n1149), .ZN(n1144) );
XOR2_X1 U817 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U818 ( .A1(n1143), .A2(G475), .ZN(n1151) );
NAND2_X1 U819 ( .A1(n1152), .A2(n1153), .ZN(n1150) );
NOR2_X1 U820 ( .A1(n1152), .A2(n1153), .ZN(n1148) );
INV_X1 U821 ( .A(KEYINPUT35), .ZN(n1153) );
XNOR2_X1 U822 ( .A(G104), .B(n1154), .ZN(G6) );
NOR2_X1 U823 ( .A1(n1155), .A2(n1156), .ZN(G57) );
XNOR2_X1 U824 ( .A(n1134), .B(KEYINPUT49), .ZN(n1156) );
NOR2_X1 U825 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
XOR2_X1 U826 ( .A(KEYINPUT12), .B(n1159), .Z(n1158) );
NOR2_X1 U827 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
AND2_X1 U828 ( .A1(n1161), .A2(n1160), .ZN(n1157) );
XOR2_X1 U829 ( .A(n1162), .B(n1163), .Z(n1160) );
XOR2_X1 U830 ( .A(n1164), .B(n1165), .Z(n1162) );
NAND3_X1 U831 ( .A1(n1166), .A2(n1167), .A3(G472), .ZN(n1164) );
OR2_X1 U832 ( .A1(n1143), .A2(KEYINPUT53), .ZN(n1167) );
NAND2_X1 U833 ( .A1(KEYINPUT53), .A2(n1168), .ZN(n1166) );
NAND2_X1 U834 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
INV_X1 U835 ( .A(n1034), .ZN(n1170) );
NOR2_X1 U836 ( .A1(n1134), .A2(n1171), .ZN(G54) );
XOR2_X1 U837 ( .A(n1172), .B(n1173), .Z(n1171) );
XNOR2_X1 U838 ( .A(n1174), .B(n1175), .ZN(n1173) );
XNOR2_X1 U839 ( .A(n1176), .B(n1177), .ZN(n1172) );
NAND2_X1 U840 ( .A1(KEYINPUT61), .A2(n1178), .ZN(n1177) );
NAND2_X1 U841 ( .A1(n1143), .A2(G469), .ZN(n1178) );
INV_X1 U842 ( .A(n1139), .ZN(n1143) );
NAND3_X1 U843 ( .A1(n1179), .A2(n1180), .A3(KEYINPUT23), .ZN(n1176) );
NAND2_X1 U844 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U845 ( .A(n1183), .B(KEYINPUT2), .Z(n1181) );
NAND2_X1 U846 ( .A1(G140), .A2(n1184), .ZN(n1179) );
XOR2_X1 U847 ( .A(n1183), .B(KEYINPUT32), .Z(n1184) );
XNOR2_X1 U848 ( .A(G110), .B(n1185), .ZN(n1183) );
NOR2_X1 U849 ( .A1(n1134), .A2(n1186), .ZN(G51) );
NOR2_X1 U850 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U851 ( .A(n1189), .B(KEYINPUT47), .Z(n1188) );
NAND2_X1 U852 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U853 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
XNOR2_X1 U854 ( .A(n1192), .B(n1193), .ZN(n1191) );
NAND4_X1 U855 ( .A1(KEYINPUT62), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
OR2_X1 U856 ( .A1(n1197), .A2(KEYINPUT54), .ZN(n1196) );
NAND3_X1 U857 ( .A1(n1197), .A2(n1198), .A3(KEYINPUT54), .ZN(n1195) );
NOR2_X1 U858 ( .A1(n1139), .A2(n1083), .ZN(n1190) );
NAND2_X1 U859 ( .A1(n1169), .A2(n1034), .ZN(n1139) );
NAND4_X1 U860 ( .A1(n1199), .A2(n1097), .A3(n1200), .A4(n1099), .ZN(n1034) );
NAND4_X1 U861 ( .A1(n1201), .A2(n1202), .A3(n1068), .A4(n1061), .ZN(n1099) );
XNOR2_X1 U862 ( .A(n1203), .B(KEYINPUT55), .ZN(n1201) );
XNOR2_X1 U863 ( .A(KEYINPUT59), .B(n1096), .ZN(n1200) );
AND4_X1 U864 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1097) );
AND3_X1 U865 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1207) );
NAND2_X1 U866 ( .A1(n1211), .A2(n1212), .ZN(n1208) );
INV_X1 U867 ( .A(n1131), .ZN(n1199) );
NAND4_X1 U868 ( .A1(n1154), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1131) );
AND3_X1 U869 ( .A1(n1029), .A2(n1216), .A3(n1217), .ZN(n1215) );
NAND3_X1 U870 ( .A1(n1067), .A2(n1052), .A3(n1218), .ZN(n1029) );
NAND2_X1 U871 ( .A1(n1219), .A2(n1220), .ZN(n1214) );
NAND4_X1 U872 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1220) );
OR3_X1 U873 ( .A1(n1225), .A2(n1048), .A3(KEYINPUT36), .ZN(n1224) );
NAND2_X1 U874 ( .A1(KEYINPUT36), .A2(n1211), .ZN(n1223) );
NAND3_X1 U875 ( .A1(n1052), .A2(n1076), .A3(n1226), .ZN(n1222) );
NAND2_X1 U876 ( .A1(n1227), .A2(n1203), .ZN(n1221) );
NAND3_X1 U877 ( .A1(n1218), .A2(n1052), .A3(n1068), .ZN(n1154) );
XNOR2_X1 U878 ( .A(G902), .B(KEYINPUT8), .ZN(n1169) );
NOR2_X1 U879 ( .A1(n1098), .A2(G952), .ZN(n1134) );
XOR2_X1 U880 ( .A(G146), .B(n1228), .Z(G48) );
NOR2_X1 U881 ( .A1(n1225), .A2(n1229), .ZN(n1228) );
XNOR2_X1 U882 ( .A(G143), .B(n1210), .ZN(G45) );
NAND3_X1 U883 ( .A1(n1048), .A2(n1202), .A3(n1230), .ZN(n1210) );
AND3_X1 U884 ( .A1(n1226), .A2(n1076), .A3(n1061), .ZN(n1230) );
XNOR2_X1 U885 ( .A(G140), .B(n1209), .ZN(G42) );
NAND2_X1 U886 ( .A1(n1212), .A2(n1231), .ZN(n1209) );
XNOR2_X1 U887 ( .A(G137), .B(n1206), .ZN(G39) );
NAND3_X1 U888 ( .A1(n1227), .A2(n1203), .A3(n1212), .ZN(n1206) );
XNOR2_X1 U889 ( .A(G134), .B(n1096), .ZN(G36) );
NAND3_X1 U890 ( .A1(n1048), .A2(n1067), .A3(n1212), .ZN(n1096) );
AND2_X1 U891 ( .A1(n1202), .A2(n1066), .ZN(n1212) );
XNOR2_X1 U892 ( .A(G131), .B(n1232), .ZN(G33) );
NAND3_X1 U893 ( .A1(n1211), .A2(n1202), .A3(n1233), .ZN(n1232) );
XNOR2_X1 U894 ( .A(KEYINPUT14), .B(n1066), .ZN(n1233) );
NAND2_X1 U895 ( .A1(n1234), .A2(n1235), .ZN(n1066) );
OR3_X1 U896 ( .A1(n1236), .A2(n1085), .A3(KEYINPUT50), .ZN(n1235) );
INV_X1 U897 ( .A(n1064), .ZN(n1236) );
NAND2_X1 U898 ( .A1(KEYINPUT50), .A2(n1061), .ZN(n1234) );
INV_X1 U899 ( .A(n1237), .ZN(n1211) );
XNOR2_X1 U900 ( .A(n1204), .B(n1238), .ZN(G30) );
NOR2_X1 U901 ( .A1(KEYINPUT42), .A2(n1239), .ZN(n1238) );
INV_X1 U902 ( .A(G128), .ZN(n1239) );
OR2_X1 U903 ( .A1(n1229), .A2(n1240), .ZN(n1204) );
NAND3_X1 U904 ( .A1(n1203), .A2(n1061), .A3(n1202), .ZN(n1229) );
AND2_X1 U905 ( .A1(n1054), .A2(n1241), .ZN(n1202) );
XNOR2_X1 U906 ( .A(G101), .B(n1213), .ZN(G3) );
NAND3_X1 U907 ( .A1(n1227), .A2(n1218), .A3(n1048), .ZN(n1213) );
XNOR2_X1 U908 ( .A(n1242), .B(n1243), .ZN(G27) );
NAND2_X1 U909 ( .A1(KEYINPUT18), .A2(n1205), .ZN(n1242) );
NAND3_X1 U910 ( .A1(n1244), .A2(n1231), .A3(n1245), .ZN(n1205) );
AND3_X1 U911 ( .A1(n1061), .A2(n1241), .A3(n1053), .ZN(n1245) );
NAND2_X1 U912 ( .A1(n1246), .A2(n1036), .ZN(n1241) );
NAND2_X1 U913 ( .A1(n1247), .A2(n1102), .ZN(n1246) );
INV_X1 U914 ( .A(G900), .ZN(n1102) );
NOR3_X1 U915 ( .A1(n1051), .A2(n1050), .A3(n1225), .ZN(n1231) );
XNOR2_X1 U916 ( .A(G122), .B(n1248), .ZN(G24) );
NAND4_X1 U917 ( .A1(n1249), .A2(n1219), .A3(n1226), .A4(n1076), .ZN(n1248) );
XNOR2_X1 U918 ( .A(n1052), .B(KEYINPUT56), .ZN(n1249) );
NOR2_X1 U919 ( .A1(n1250), .A2(n1051), .ZN(n1052) );
XNOR2_X1 U920 ( .A(G119), .B(n1251), .ZN(G21) );
NAND4_X1 U921 ( .A1(n1252), .A2(n1253), .A3(n1227), .A4(n1203), .ZN(n1251) );
NOR2_X1 U922 ( .A1(n1254), .A2(n1050), .ZN(n1203) );
XNOR2_X1 U923 ( .A(n1061), .B(KEYINPUT27), .ZN(n1252) );
XNOR2_X1 U924 ( .A(G116), .B(n1217), .ZN(G18) );
NAND3_X1 U925 ( .A1(n1219), .A2(n1067), .A3(n1048), .ZN(n1217) );
INV_X1 U926 ( .A(n1240), .ZN(n1067) );
NAND2_X1 U927 ( .A1(n1255), .A2(n1076), .ZN(n1240) );
INV_X1 U928 ( .A(n1256), .ZN(n1219) );
XOR2_X1 U929 ( .A(G113), .B(n1257), .Z(G15) );
NOR3_X1 U930 ( .A1(n1237), .A2(KEYINPUT41), .A3(n1256), .ZN(n1257) );
NAND2_X1 U931 ( .A1(n1253), .A2(n1061), .ZN(n1256) );
AND3_X1 U932 ( .A1(n1053), .A2(n1258), .A3(n1244), .ZN(n1253) );
NAND2_X1 U933 ( .A1(n1048), .A2(n1068), .ZN(n1237) );
INV_X1 U934 ( .A(n1225), .ZN(n1068) );
NAND2_X1 U935 ( .A1(n1259), .A2(n1226), .ZN(n1225) );
XOR2_X1 U936 ( .A(n1255), .B(KEYINPUT57), .Z(n1226) );
NOR2_X1 U937 ( .A1(n1250), .A2(n1254), .ZN(n1048) );
XNOR2_X1 U938 ( .A(n1216), .B(n1260), .ZN(G12) );
NOR2_X1 U939 ( .A1(KEYINPUT25), .A2(n1261), .ZN(n1260) );
NAND4_X1 U940 ( .A1(n1227), .A2(n1218), .A3(n1254), .A4(n1250), .ZN(n1216) );
INV_X1 U941 ( .A(n1050), .ZN(n1250) );
NOR2_X1 U942 ( .A1(n1262), .A2(n1084), .ZN(n1050) );
NOR3_X1 U943 ( .A1(n1086), .A2(G902), .A3(n1263), .ZN(n1084) );
INV_X1 U944 ( .A(n1136), .ZN(n1263) );
AND2_X1 U945 ( .A1(n1264), .A2(n1087), .ZN(n1262) );
NAND2_X1 U946 ( .A1(n1136), .A2(n1265), .ZN(n1087) );
XNOR2_X1 U947 ( .A(n1266), .B(n1267), .ZN(n1136) );
NOR2_X1 U948 ( .A1(KEYINPUT44), .A2(n1268), .ZN(n1267) );
XOR2_X1 U949 ( .A(n1269), .B(n1270), .Z(n1268) );
XNOR2_X1 U950 ( .A(n1271), .B(n1272), .ZN(n1270) );
INV_X1 U951 ( .A(n1273), .ZN(n1271) );
XNOR2_X1 U952 ( .A(G119), .B(n1274), .ZN(n1269) );
XNOR2_X1 U953 ( .A(KEYINPUT51), .B(n1243), .ZN(n1274) );
INV_X1 U954 ( .A(G125), .ZN(n1243) );
NAND2_X1 U955 ( .A1(n1275), .A2(n1276), .ZN(n1266) );
NAND2_X1 U956 ( .A1(n1277), .A2(G137), .ZN(n1276) );
XOR2_X1 U957 ( .A(KEYINPUT34), .B(n1278), .Z(n1275) );
NOR2_X1 U958 ( .A1(n1277), .A2(G137), .ZN(n1278) );
AND2_X1 U959 ( .A1(n1279), .A2(G221), .ZN(n1277) );
XNOR2_X1 U960 ( .A(n1086), .B(KEYINPUT15), .ZN(n1264) );
INV_X1 U961 ( .A(n1138), .ZN(n1086) );
NAND2_X1 U962 ( .A1(G217), .A2(n1280), .ZN(n1138) );
INV_X1 U963 ( .A(n1051), .ZN(n1254) );
XNOR2_X1 U964 ( .A(n1078), .B(G472), .ZN(n1051) );
NAND2_X1 U965 ( .A1(n1281), .A2(n1265), .ZN(n1078) );
XOR2_X1 U966 ( .A(n1282), .B(n1283), .Z(n1281) );
XNOR2_X1 U967 ( .A(n1284), .B(n1161), .ZN(n1283) );
XNOR2_X1 U968 ( .A(n1285), .B(G101), .ZN(n1161) );
NAND2_X1 U969 ( .A1(n1286), .A2(G210), .ZN(n1285) );
NAND2_X1 U970 ( .A1(n1287), .A2(n1288), .ZN(n1284) );
NAND2_X1 U971 ( .A1(n1289), .A2(n1165), .ZN(n1288) );
XOR2_X1 U972 ( .A(KEYINPUT38), .B(n1290), .Z(n1287) );
NOR2_X1 U973 ( .A1(n1289), .A2(n1165), .ZN(n1290) );
XNOR2_X1 U974 ( .A(n1291), .B(n1292), .ZN(n1165) );
INV_X1 U975 ( .A(n1174), .ZN(n1291) );
XNOR2_X1 U976 ( .A(n1163), .B(KEYINPUT43), .ZN(n1289) );
XOR2_X1 U977 ( .A(n1293), .B(n1294), .Z(n1163) );
XOR2_X1 U978 ( .A(KEYINPUT30), .B(n1295), .Z(n1294) );
XOR2_X1 U979 ( .A(KEYINPUT48), .B(KEYINPUT40), .Z(n1282) );
AND3_X1 U980 ( .A1(n1061), .A2(n1258), .A3(n1054), .ZN(n1218) );
NOR2_X1 U981 ( .A1(n1244), .A2(n1047), .ZN(n1054) );
INV_X1 U982 ( .A(n1053), .ZN(n1047) );
NAND2_X1 U983 ( .A1(G221), .A2(n1280), .ZN(n1053) );
NAND2_X1 U984 ( .A1(G234), .A2(n1265), .ZN(n1280) );
INV_X1 U985 ( .A(n1044), .ZN(n1244) );
XOR2_X1 U986 ( .A(n1088), .B(n1090), .Z(n1044) );
INV_X1 U987 ( .A(G469), .ZN(n1090) );
NAND3_X1 U988 ( .A1(n1296), .A2(n1265), .A3(n1297), .ZN(n1088) );
NAND3_X1 U989 ( .A1(n1174), .A2(n1298), .A3(n1299), .ZN(n1297) );
XOR2_X1 U990 ( .A(n1300), .B(n1301), .Z(n1299) );
NAND2_X1 U991 ( .A1(KEYINPUT16), .A2(n1302), .ZN(n1300) );
NAND2_X1 U992 ( .A1(n1303), .A2(n1304), .ZN(n1296) );
NAND2_X1 U993 ( .A1(n1174), .A2(n1298), .ZN(n1304) );
INV_X1 U994 ( .A(KEYINPUT52), .ZN(n1298) );
XOR2_X1 U995 ( .A(n1305), .B(n1110), .Z(n1174) );
XNOR2_X1 U996 ( .A(G134), .B(G137), .ZN(n1110) );
XNOR2_X1 U997 ( .A(G131), .B(KEYINPUT7), .ZN(n1305) );
XNOR2_X1 U998 ( .A(n1301), .B(n1306), .ZN(n1303) );
NOR2_X1 U999 ( .A1(n1302), .A2(n1307), .ZN(n1306) );
INV_X1 U1000 ( .A(KEYINPUT16), .ZN(n1307) );
NAND2_X1 U1001 ( .A1(n1308), .A2(n1309), .ZN(n1302) );
NAND2_X1 U1002 ( .A1(n1175), .A2(n1310), .ZN(n1309) );
XOR2_X1 U1003 ( .A(n1311), .B(n1104), .Z(n1175) );
OR3_X1 U1004 ( .A1(n1311), .A2(n1104), .A3(n1310), .ZN(n1308) );
INV_X1 U1005 ( .A(KEYINPUT58), .ZN(n1310) );
XOR2_X1 U1006 ( .A(n1273), .B(n1312), .Z(n1104) );
XOR2_X1 U1007 ( .A(n1313), .B(n1314), .Z(n1311) );
XOR2_X1 U1008 ( .A(G104), .B(G101), .Z(n1314) );
NAND2_X1 U1009 ( .A1(KEYINPUT46), .A2(n1315), .ZN(n1313) );
XOR2_X1 U1010 ( .A(n1185), .B(n1272), .Z(n1301) );
XNOR2_X1 U1011 ( .A(n1261), .B(G140), .ZN(n1272) );
AND2_X1 U1012 ( .A1(G227), .A2(n1098), .ZN(n1185) );
NAND2_X1 U1013 ( .A1(n1036), .A2(n1316), .ZN(n1258) );
NAND2_X1 U1014 ( .A1(n1247), .A2(n1317), .ZN(n1316) );
XOR2_X1 U1015 ( .A(KEYINPUT19), .B(G898), .Z(n1317) );
AND3_X1 U1016 ( .A1(G902), .A2(n1318), .A3(G953), .ZN(n1247) );
NAND3_X1 U1017 ( .A1(n1318), .A2(n1098), .A3(G952), .ZN(n1036) );
NAND2_X1 U1018 ( .A1(G237), .A2(G234), .ZN(n1318) );
NOR2_X1 U1019 ( .A1(n1064), .A2(n1085), .ZN(n1061) );
INV_X1 U1020 ( .A(n1063), .ZN(n1085) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1319), .ZN(n1063) );
XOR2_X1 U1022 ( .A(n1320), .B(n1083), .Z(n1064) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1319), .ZN(n1083) );
NAND2_X1 U1024 ( .A1(n1321), .A2(n1265), .ZN(n1319) );
INV_X1 U1025 ( .A(G237), .ZN(n1321) );
NAND2_X1 U1026 ( .A1(KEYINPUT33), .A2(n1082), .ZN(n1320) );
NAND3_X1 U1027 ( .A1(n1322), .A2(n1265), .A3(n1323), .ZN(n1082) );
XOR2_X1 U1028 ( .A(n1324), .B(KEYINPUT9), .Z(n1323) );
OR2_X1 U1029 ( .A1(n1325), .A2(n1193), .ZN(n1324) );
NAND2_X1 U1030 ( .A1(n1193), .A2(n1325), .ZN(n1322) );
NAND2_X1 U1031 ( .A1(n1194), .A2(n1326), .ZN(n1325) );
NAND2_X1 U1032 ( .A1(n1197), .A2(n1198), .ZN(n1326) );
OR2_X1 U1033 ( .A1(n1198), .A2(n1197), .ZN(n1194) );
XNOR2_X1 U1034 ( .A(G125), .B(n1292), .ZN(n1197) );
XNOR2_X1 U1035 ( .A(n1327), .B(n1273), .ZN(n1292) );
XOR2_X1 U1036 ( .A(G128), .B(G146), .Z(n1273) );
XNOR2_X1 U1037 ( .A(KEYINPUT4), .B(n1328), .ZN(n1327) );
NOR2_X1 U1038 ( .A1(KEYINPUT17), .A2(n1312), .ZN(n1328) );
NAND2_X1 U1039 ( .A1(G224), .A2(n1098), .ZN(n1198) );
XNOR2_X1 U1040 ( .A(n1329), .B(n1130), .ZN(n1193) );
XNOR2_X1 U1041 ( .A(n1261), .B(G122), .ZN(n1130) );
INV_X1 U1042 ( .A(G110), .ZN(n1261) );
XNOR2_X1 U1043 ( .A(n1128), .B(n1129), .ZN(n1329) );
XNOR2_X1 U1044 ( .A(n1330), .B(G101), .ZN(n1129) );
NAND2_X1 U1045 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NAND2_X1 U1046 ( .A1(G104), .A2(n1315), .ZN(n1332) );
XOR2_X1 U1047 ( .A(KEYINPUT39), .B(n1333), .Z(n1331) );
NOR2_X1 U1048 ( .A1(G104), .A2(n1315), .ZN(n1333) );
AND2_X1 U1049 ( .A1(n1334), .A2(n1335), .ZN(n1128) );
OR2_X1 U1050 ( .A1(n1293), .A2(n1295), .ZN(n1335) );
XOR2_X1 U1051 ( .A(n1336), .B(KEYINPUT29), .Z(n1334) );
NAND2_X1 U1052 ( .A1(n1295), .A2(n1293), .ZN(n1336) );
XNOR2_X1 U1053 ( .A(G116), .B(n1337), .ZN(n1295) );
INV_X1 U1054 ( .A(G119), .ZN(n1337) );
INV_X1 U1055 ( .A(n1039), .ZN(n1227) );
NAND2_X1 U1056 ( .A1(n1259), .A2(n1255), .ZN(n1039) );
XOR2_X1 U1057 ( .A(n1079), .B(G475), .Z(n1255) );
NAND2_X1 U1058 ( .A1(n1152), .A2(n1265), .ZN(n1079) );
XOR2_X1 U1059 ( .A(n1338), .B(n1339), .Z(n1152) );
XOR2_X1 U1060 ( .A(n1340), .B(n1341), .Z(n1339) );
XNOR2_X1 U1061 ( .A(n1106), .B(n1293), .ZN(n1341) );
XOR2_X1 U1062 ( .A(G113), .B(KEYINPUT45), .Z(n1293) );
XNOR2_X1 U1063 ( .A(G125), .B(n1182), .ZN(n1106) );
INV_X1 U1064 ( .A(G140), .ZN(n1182) );
XOR2_X1 U1065 ( .A(n1342), .B(n1343), .Z(n1340) );
NOR2_X1 U1066 ( .A1(KEYINPUT1), .A2(n1312), .ZN(n1343) );
NAND2_X1 U1067 ( .A1(n1286), .A2(G214), .ZN(n1342) );
NOR2_X1 U1068 ( .A1(G953), .A2(G237), .ZN(n1286) );
XOR2_X1 U1069 ( .A(n1344), .B(n1345), .Z(n1338) );
XOR2_X1 U1070 ( .A(G122), .B(G104), .Z(n1345) );
XNOR2_X1 U1071 ( .A(G146), .B(G131), .ZN(n1344) );
XNOR2_X1 U1072 ( .A(n1076), .B(KEYINPUT5), .ZN(n1259) );
XOR2_X1 U1073 ( .A(G478), .B(n1346), .Z(n1076) );
AND2_X1 U1074 ( .A1(n1141), .A2(n1265), .ZN(n1346) );
INV_X1 U1075 ( .A(G902), .ZN(n1265) );
NAND2_X1 U1076 ( .A1(n1347), .A2(n1348), .ZN(n1141) );
NAND2_X1 U1077 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1078 ( .A1(G217), .A2(n1279), .ZN(n1350) );
INV_X1 U1079 ( .A(n1351), .ZN(n1279) );
XOR2_X1 U1080 ( .A(KEYINPUT63), .B(n1352), .Z(n1347) );
NOR3_X1 U1081 ( .A1(n1353), .A2(n1351), .A3(n1354), .ZN(n1352) );
INV_X1 U1082 ( .A(G217), .ZN(n1354) );
NAND2_X1 U1083 ( .A1(G234), .A2(n1098), .ZN(n1351) );
INV_X1 U1084 ( .A(G953), .ZN(n1098) );
XNOR2_X1 U1085 ( .A(KEYINPUT11), .B(n1349), .ZN(n1353) );
XOR2_X1 U1086 ( .A(n1355), .B(n1356), .Z(n1349) );
XNOR2_X1 U1087 ( .A(n1357), .B(n1312), .ZN(n1356) );
XOR2_X1 U1088 ( .A(G143), .B(KEYINPUT24), .Z(n1312) );
NAND2_X1 U1089 ( .A1(KEYINPUT3), .A2(n1358), .ZN(n1357) );
XOR2_X1 U1090 ( .A(n1359), .B(n1360), .Z(n1358) );
XNOR2_X1 U1091 ( .A(G122), .B(n1315), .ZN(n1360) );
INV_X1 U1092 ( .A(G107), .ZN(n1315) );
NOR2_X1 U1093 ( .A1(G116), .A2(KEYINPUT20), .ZN(n1359) );
XNOR2_X1 U1094 ( .A(G128), .B(G134), .ZN(n1355) );
endmodule


