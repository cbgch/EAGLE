//Key = 1101100010000011111100010101010111001011010101011011000110001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361;

XOR2_X1 U748 ( .A(G107), .B(n1032), .Z(G9) );
NOR2_X1 U749 ( .A1(n1033), .A2(n1034), .ZN(G75) );
NOR3_X1 U750 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NAND3_X1 U751 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1035) );
NAND4_X1 U752 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1040) );
NAND2_X1 U753 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND3_X1 U754 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND2_X1 U755 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
OR3_X1 U756 ( .A1(n1052), .A2(n1053), .A3(n1050), .ZN(n1047) );
AND2_X1 U757 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U758 ( .A1(n1056), .A2(n1057), .ZN(n1045) );
NAND4_X1 U759 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1038) );
NAND2_X1 U760 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND3_X1 U761 ( .A1(n1063), .A2(n1064), .A3(n1042), .ZN(n1061) );
INV_X1 U762 ( .A(KEYINPUT0), .ZN(n1064) );
NAND3_X1 U763 ( .A1(n1065), .A2(n1066), .A3(n1041), .ZN(n1059) );
INV_X1 U764 ( .A(n1062), .ZN(n1041) );
NAND2_X1 U765 ( .A1(n1042), .A2(n1067), .ZN(n1066) );
NAND2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U767 ( .A1(KEYINPUT0), .A2(n1063), .ZN(n1069) );
NAND2_X1 U768 ( .A1(n1043), .A2(n1070), .ZN(n1065) );
NAND2_X1 U769 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U770 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XNOR2_X1 U771 ( .A(n1075), .B(KEYINPUT60), .ZN(n1073) );
INV_X1 U772 ( .A(n1076), .ZN(n1071) );
NOR3_X1 U773 ( .A1(n1037), .A2(G952), .A3(n1077), .ZN(n1033) );
INV_X1 U774 ( .A(n1039), .ZN(n1077) );
NAND4_X1 U775 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1039) );
NOR4_X1 U776 ( .A1(n1082), .A2(n1083), .A3(n1050), .A4(n1084), .ZN(n1081) );
XOR2_X1 U777 ( .A(n1085), .B(n1086), .Z(n1083) );
XOR2_X1 U778 ( .A(n1087), .B(KEYINPUT50), .Z(n1086) );
NAND2_X1 U779 ( .A1(KEYINPUT36), .A2(n1088), .ZN(n1085) );
NAND3_X1 U780 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1082) );
XNOR2_X1 U781 ( .A(n1092), .B(G472), .ZN(n1091) );
OR3_X1 U782 ( .A1(n1093), .A2(n1094), .A3(KEYINPUT7), .ZN(n1090) );
NAND2_X1 U783 ( .A1(KEYINPUT7), .A2(n1094), .ZN(n1089) );
NOR3_X1 U784 ( .A1(n1054), .A2(n1075), .A3(n1095), .ZN(n1080) );
XOR2_X1 U785 ( .A(KEYINPUT8), .B(n1096), .Z(n1078) );
NOR2_X1 U786 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XNOR2_X1 U787 ( .A(G469), .B(KEYINPUT37), .ZN(n1098) );
INV_X1 U788 ( .A(n1099), .ZN(n1097) );
NAND2_X1 U789 ( .A1(n1100), .A2(n1101), .ZN(G72) );
NAND4_X1 U790 ( .A1(G953), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1101) );
NAND2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1100) );
NAND2_X1 U792 ( .A1(n1107), .A2(n1103), .ZN(n1106) );
NAND4_X1 U793 ( .A1(n1108), .A2(n1109), .A3(n1110), .A4(n1111), .ZN(n1103) );
NAND2_X1 U794 ( .A1(G953), .A2(n1112), .ZN(n1111) );
NAND2_X1 U795 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
XNOR2_X1 U796 ( .A(n1115), .B(n1104), .ZN(n1107) );
INV_X1 U797 ( .A(KEYINPUT11), .ZN(n1104) );
NAND3_X1 U798 ( .A1(n1113), .A2(n1114), .A3(n1116), .ZN(n1115) );
NAND2_X1 U799 ( .A1(n1108), .A2(n1109), .ZN(n1116) );
NAND2_X1 U800 ( .A1(n1117), .A2(n1118), .ZN(n1109) );
XNOR2_X1 U801 ( .A(n1119), .B(n1120), .ZN(n1117) );
XOR2_X1 U802 ( .A(n1121), .B(KEYINPUT49), .Z(n1108) );
NAND2_X1 U803 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XOR2_X1 U804 ( .A(n1119), .B(n1120), .Z(n1123) );
NAND2_X1 U805 ( .A1(n1124), .A2(n1125), .ZN(n1119) );
NAND2_X1 U806 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U807 ( .A(KEYINPUT4), .B(n1128), .Z(n1124) );
NOR2_X1 U808 ( .A1(n1126), .A2(n1127), .ZN(n1128) );
XNOR2_X1 U809 ( .A(KEYINPUT52), .B(n1118), .ZN(n1122) );
NAND2_X1 U810 ( .A1(n1129), .A2(n1130), .ZN(n1118) );
NAND2_X1 U811 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U812 ( .A1(KEYINPUT45), .A2(n1133), .ZN(n1131) );
NAND2_X1 U813 ( .A1(KEYINPUT45), .A2(n1134), .ZN(n1129) );
NAND2_X1 U814 ( .A1(n1135), .A2(n1136), .ZN(n1113) );
XOR2_X1 U815 ( .A(KEYINPUT57), .B(n1137), .Z(n1136) );
NAND2_X1 U816 ( .A1(G953), .A2(n1102), .ZN(n1105) );
NAND2_X1 U817 ( .A1(G900), .A2(G227), .ZN(n1102) );
XOR2_X1 U818 ( .A(n1138), .B(n1139), .Z(G69) );
NOR2_X1 U819 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U820 ( .A(n1142), .B(KEYINPUT29), .Z(n1141) );
NAND3_X1 U821 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1142) );
NAND2_X1 U822 ( .A1(G953), .A2(n1146), .ZN(n1144) );
NAND2_X1 U823 ( .A1(n1147), .A2(n1114), .ZN(n1143) );
NAND2_X1 U824 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NOR3_X1 U825 ( .A1(n1145), .A2(G953), .A3(n1150), .ZN(n1140) );
AND2_X1 U826 ( .A1(n1149), .A2(n1148), .ZN(n1150) );
XNOR2_X1 U827 ( .A(KEYINPUT17), .B(n1151), .ZN(n1145) );
NAND2_X1 U828 ( .A1(G953), .A2(n1152), .ZN(n1138) );
NAND2_X1 U829 ( .A1(G898), .A2(G224), .ZN(n1152) );
NOR2_X1 U830 ( .A1(n1153), .A2(n1154), .ZN(G66) );
XOR2_X1 U831 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND3_X1 U832 ( .A1(n1157), .A2(G217), .A3(KEYINPUT48), .ZN(n1155) );
NOR2_X1 U833 ( .A1(n1153), .A2(n1158), .ZN(G63) );
XOR2_X1 U834 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND3_X1 U835 ( .A1(G478), .A2(n1036), .A3(n1161), .ZN(n1159) );
XNOR2_X1 U836 ( .A(G902), .B(KEYINPUT39), .ZN(n1161) );
NOR2_X1 U837 ( .A1(n1153), .A2(n1162), .ZN(G60) );
NOR3_X1 U838 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1162) );
NOR3_X1 U839 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1165) );
NOR3_X1 U840 ( .A1(n1169), .A2(n1093), .A3(n1170), .ZN(n1167) );
NOR2_X1 U841 ( .A1(KEYINPUT33), .A2(n1171), .ZN(n1164) );
NOR3_X1 U842 ( .A1(n1170), .A2(n1172), .A3(n1093), .ZN(n1163) );
NOR2_X1 U843 ( .A1(n1173), .A2(n1166), .ZN(n1172) );
INV_X1 U844 ( .A(KEYINPUT33), .ZN(n1166) );
NOR2_X1 U845 ( .A1(n1171), .A2(n1169), .ZN(n1173) );
INV_X1 U846 ( .A(KEYINPUT55), .ZN(n1169) );
INV_X1 U847 ( .A(n1168), .ZN(n1171) );
XNOR2_X1 U848 ( .A(G104), .B(n1174), .ZN(G6) );
NOR2_X1 U849 ( .A1(n1153), .A2(n1175), .ZN(G57) );
XOR2_X1 U850 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U851 ( .A(n1178), .B(n1179), .Z(n1177) );
AND2_X1 U852 ( .A1(G472), .A2(n1157), .ZN(n1178) );
INV_X1 U853 ( .A(n1170), .ZN(n1157) );
XOR2_X1 U854 ( .A(n1180), .B(n1181), .Z(n1176) );
XNOR2_X1 U855 ( .A(n1182), .B(n1183), .ZN(n1181) );
NAND2_X1 U856 ( .A1(n1184), .A2(KEYINPUT16), .ZN(n1183) );
XNOR2_X1 U857 ( .A(G101), .B(KEYINPUT12), .ZN(n1184) );
NAND3_X1 U858 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1180) );
NAND2_X1 U859 ( .A1(KEYINPUT42), .A2(n1188), .ZN(n1187) );
NAND3_X1 U860 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1186) );
INV_X1 U861 ( .A(KEYINPUT42), .ZN(n1190) );
OR2_X1 U862 ( .A1(n1191), .A2(n1189), .ZN(n1185) );
NOR2_X1 U863 ( .A1(KEYINPUT30), .A2(n1188), .ZN(n1189) );
NOR2_X1 U864 ( .A1(n1153), .A2(n1192), .ZN(G54) );
XOR2_X1 U865 ( .A(n1193), .B(n1194), .Z(n1192) );
XNOR2_X1 U866 ( .A(n1195), .B(n1120), .ZN(n1194) );
XNOR2_X1 U867 ( .A(n1196), .B(n1191), .ZN(n1193) );
XOR2_X1 U868 ( .A(n1197), .B(n1198), .Z(n1196) );
NOR2_X1 U869 ( .A1(n1199), .A2(n1170), .ZN(n1198) );
NAND2_X1 U870 ( .A1(n1200), .A2(n1201), .ZN(n1197) );
NAND2_X1 U871 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NAND2_X1 U872 ( .A1(G227), .A2(n1114), .ZN(n1203) );
XNOR2_X1 U873 ( .A(n1204), .B(KEYINPUT2), .ZN(n1200) );
NOR2_X1 U874 ( .A1(n1153), .A2(n1205), .ZN(G51) );
XOR2_X1 U875 ( .A(n1206), .B(n1207), .Z(n1205) );
XNOR2_X1 U876 ( .A(n1208), .B(n1151), .ZN(n1207) );
NOR2_X1 U877 ( .A1(n1209), .A2(n1170), .ZN(n1208) );
NAND2_X1 U878 ( .A1(G902), .A2(n1036), .ZN(n1170) );
NAND4_X1 U879 ( .A1(n1210), .A2(n1137), .A3(n1148), .A4(n1135), .ZN(n1036) );
AND3_X1 U880 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1135) );
NAND3_X1 U881 ( .A1(n1057), .A2(n1214), .A3(n1215), .ZN(n1213) );
NAND2_X1 U882 ( .A1(n1068), .A2(n1216), .ZN(n1214) );
AND4_X1 U883 ( .A1(n1217), .A2(n1218), .A3(n1174), .A4(n1219), .ZN(n1148) );
NOR4_X1 U884 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1032), .ZN(n1219) );
AND3_X1 U885 ( .A1(n1063), .A2(n1058), .A3(n1223), .ZN(n1032) );
NAND3_X1 U886 ( .A1(n1223), .A2(n1058), .A3(n1224), .ZN(n1174) );
NAND2_X1 U887 ( .A1(n1225), .A2(n1226), .ZN(n1217) );
AND4_X1 U888 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1137) );
NAND3_X1 U889 ( .A1(n1231), .A2(n1057), .A3(n1043), .ZN(n1227) );
XOR2_X1 U890 ( .A(n1149), .B(KEYINPUT21), .Z(n1210) );
XNOR2_X1 U891 ( .A(G210), .B(KEYINPUT59), .ZN(n1209) );
NOR2_X1 U892 ( .A1(n1114), .A2(G952), .ZN(n1153) );
XNOR2_X1 U893 ( .A(G146), .B(n1228), .ZN(G48) );
NAND3_X1 U894 ( .A1(n1224), .A2(n1052), .A3(n1231), .ZN(n1228) );
XNOR2_X1 U895 ( .A(n1232), .B(n1229), .ZN(G45) );
NAND2_X1 U896 ( .A1(n1233), .A2(n1215), .ZN(n1229) );
NAND2_X1 U897 ( .A1(KEYINPUT43), .A2(n1234), .ZN(n1232) );
XNOR2_X1 U898 ( .A(G140), .B(n1230), .ZN(G42) );
NAND3_X1 U899 ( .A1(n1235), .A2(n1076), .A3(n1057), .ZN(n1230) );
XOR2_X1 U900 ( .A(G137), .B(n1236), .Z(G39) );
NOR3_X1 U901 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1236) );
INV_X1 U902 ( .A(n1043), .ZN(n1239) );
XNOR2_X1 U903 ( .A(KEYINPUT41), .B(n1051), .ZN(n1237) );
NAND2_X1 U904 ( .A1(n1240), .A2(n1241), .ZN(G36) );
NAND2_X1 U905 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U906 ( .A(KEYINPUT51), .B(n1244), .Z(n1240) );
NOR2_X1 U907 ( .A1(n1242), .A2(n1243), .ZN(n1244) );
INV_X1 U908 ( .A(G134), .ZN(n1243) );
AND2_X1 U909 ( .A1(n1057), .A2(n1245), .ZN(n1242) );
XOR2_X1 U910 ( .A(KEYINPUT9), .B(n1246), .Z(n1245) );
NOR2_X1 U911 ( .A1(n1216), .A2(n1247), .ZN(n1246) );
INV_X1 U912 ( .A(n1063), .ZN(n1216) );
XOR2_X1 U913 ( .A(n1248), .B(n1249), .Z(G33) );
NAND2_X1 U914 ( .A1(KEYINPUT18), .A2(G131), .ZN(n1249) );
NAND3_X1 U915 ( .A1(n1215), .A2(n1057), .A3(n1250), .ZN(n1248) );
XNOR2_X1 U916 ( .A(n1224), .B(KEYINPUT25), .ZN(n1250) );
INV_X1 U917 ( .A(n1051), .ZN(n1057) );
NAND2_X1 U918 ( .A1(n1055), .A2(n1251), .ZN(n1051) );
INV_X1 U919 ( .A(n1247), .ZN(n1215) );
NAND3_X1 U920 ( .A1(n1076), .A2(n1252), .A3(n1056), .ZN(n1247) );
XOR2_X1 U921 ( .A(n1211), .B(n1253), .Z(G30) );
NAND2_X1 U922 ( .A1(KEYINPUT61), .A2(G128), .ZN(n1253) );
NAND3_X1 U923 ( .A1(n1063), .A2(n1052), .A3(n1231), .ZN(n1211) );
INV_X1 U924 ( .A(n1238), .ZN(n1231) );
NAND4_X1 U925 ( .A1(n1254), .A2(n1076), .A3(n1050), .A4(n1252), .ZN(n1238) );
XNOR2_X1 U926 ( .A(G101), .B(n1218), .ZN(G3) );
NAND3_X1 U927 ( .A1(n1056), .A2(n1223), .A3(n1043), .ZN(n1218) );
XNOR2_X1 U928 ( .A(G125), .B(n1212), .ZN(G27) );
NAND3_X1 U929 ( .A1(n1235), .A2(n1052), .A3(n1042), .ZN(n1212) );
AND4_X1 U930 ( .A1(n1224), .A2(n1050), .A3(n1049), .A4(n1252), .ZN(n1235) );
NAND2_X1 U931 ( .A1(n1062), .A2(n1255), .ZN(n1252) );
NAND4_X1 U932 ( .A1(G953), .A2(G902), .A3(n1256), .A4(n1112), .ZN(n1255) );
INV_X1 U933 ( .A(G900), .ZN(n1112) );
XNOR2_X1 U934 ( .A(G122), .B(n1149), .ZN(G24) );
NAND4_X1 U935 ( .A1(n1042), .A2(n1233), .A3(n1058), .A4(n1257), .ZN(n1149) );
NOR2_X1 U936 ( .A1(n1050), .A2(n1254), .ZN(n1058) );
AND3_X1 U937 ( .A1(n1052), .A2(n1258), .A3(n1259), .ZN(n1233) );
XNOR2_X1 U938 ( .A(n1084), .B(KEYINPUT23), .ZN(n1259) );
XNOR2_X1 U939 ( .A(G119), .B(n1260), .ZN(G21) );
NAND2_X1 U940 ( .A1(KEYINPUT3), .A2(n1222), .ZN(n1260) );
AND4_X1 U941 ( .A1(n1261), .A2(n1043), .A3(n1254), .A4(n1050), .ZN(n1222) );
INV_X1 U942 ( .A(n1049), .ZN(n1254) );
XNOR2_X1 U943 ( .A(G116), .B(n1262), .ZN(G18) );
NAND2_X1 U944 ( .A1(KEYINPUT1), .A2(n1221), .ZN(n1262) );
AND3_X1 U945 ( .A1(n1056), .A2(n1063), .A3(n1261), .ZN(n1221) );
AND3_X1 U946 ( .A1(n1052), .A2(n1257), .A3(n1042), .ZN(n1261) );
XOR2_X1 U947 ( .A(n1226), .B(KEYINPUT62), .Z(n1052) );
NOR2_X1 U948 ( .A1(n1258), .A2(n1263), .ZN(n1063) );
XNOR2_X1 U949 ( .A(G113), .B(n1264), .ZN(G15) );
NAND3_X1 U950 ( .A1(n1225), .A2(n1265), .A3(KEYINPUT14), .ZN(n1264) );
XOR2_X1 U951 ( .A(KEYINPUT54), .B(n1226), .Z(n1265) );
AND4_X1 U952 ( .A1(n1042), .A2(n1056), .A3(n1224), .A4(n1257), .ZN(n1225) );
INV_X1 U953 ( .A(n1068), .ZN(n1224) );
NAND2_X1 U954 ( .A1(n1263), .A2(n1258), .ZN(n1068) );
INV_X1 U955 ( .A(n1084), .ZN(n1263) );
NOR2_X1 U956 ( .A1(n1049), .A2(n1050), .ZN(n1056) );
NOR2_X1 U957 ( .A1(n1266), .A2(n1267), .ZN(n1042) );
INV_X1 U958 ( .A(n1074), .ZN(n1266) );
XOR2_X1 U959 ( .A(G110), .B(n1220), .Z(G12) );
AND4_X1 U960 ( .A1(n1043), .A2(n1223), .A3(n1050), .A4(n1049), .ZN(n1220) );
XOR2_X1 U961 ( .A(G472), .B(n1268), .Z(n1049) );
NOR2_X1 U962 ( .A1(n1092), .A2(KEYINPUT63), .ZN(n1268) );
AND2_X1 U963 ( .A1(n1269), .A2(n1270), .ZN(n1092) );
XOR2_X1 U964 ( .A(n1179), .B(n1271), .Z(n1269) );
XNOR2_X1 U965 ( .A(n1272), .B(n1273), .ZN(n1271) );
NOR2_X1 U966 ( .A1(KEYINPUT58), .A2(n1274), .ZN(n1273) );
XNOR2_X1 U967 ( .A(n1188), .B(n1191), .ZN(n1274) );
INV_X1 U968 ( .A(n1275), .ZN(n1191) );
NAND2_X1 U969 ( .A1(KEYINPUT19), .A2(n1276), .ZN(n1272) );
XOR2_X1 U970 ( .A(G101), .B(n1182), .Z(n1276) );
AND3_X1 U971 ( .A1(n1277), .A2(n1114), .A3(G210), .ZN(n1182) );
XNOR2_X1 U972 ( .A(n1278), .B(n1279), .ZN(n1179) );
NOR2_X1 U973 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
AND3_X1 U974 ( .A1(KEYINPUT10), .A2(n1282), .A3(G116), .ZN(n1281) );
NOR2_X1 U975 ( .A1(KEYINPUT10), .A2(n1283), .ZN(n1280) );
XNOR2_X1 U976 ( .A(n1284), .B(n1285), .ZN(n1050) );
NOR2_X1 U977 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XNOR2_X1 U978 ( .A(G217), .B(KEYINPUT26), .ZN(n1287) );
INV_X1 U979 ( .A(n1288), .ZN(n1286) );
NAND2_X1 U980 ( .A1(n1156), .A2(n1270), .ZN(n1284) );
XNOR2_X1 U981 ( .A(n1289), .B(n1290), .ZN(n1156) );
XOR2_X1 U982 ( .A(n1291), .B(n1292), .Z(n1290) );
XNOR2_X1 U983 ( .A(G110), .B(G119), .ZN(n1292) );
NAND2_X1 U984 ( .A1(KEYINPUT56), .A2(n1293), .ZN(n1291) );
XNOR2_X1 U985 ( .A(G137), .B(n1294), .ZN(n1293) );
NAND2_X1 U986 ( .A1(n1295), .A2(G221), .ZN(n1294) );
XOR2_X1 U987 ( .A(n1296), .B(n1297), .Z(n1289) );
NOR2_X1 U988 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NOR2_X1 U989 ( .A1(n1133), .A2(n1300), .ZN(n1298) );
NAND2_X1 U990 ( .A1(KEYINPUT32), .A2(G128), .ZN(n1296) );
AND3_X1 U991 ( .A1(n1226), .A2(n1257), .A3(n1076), .ZN(n1223) );
NOR2_X1 U992 ( .A1(n1267), .A2(n1074), .ZN(n1076) );
NOR2_X1 U993 ( .A1(n1301), .A2(n1095), .ZN(n1074) );
NOR2_X1 U994 ( .A1(n1099), .A2(G469), .ZN(n1095) );
AND2_X1 U995 ( .A1(n1302), .A2(n1099), .ZN(n1301) );
NAND2_X1 U996 ( .A1(n1303), .A2(n1270), .ZN(n1099) );
XOR2_X1 U997 ( .A(n1304), .B(n1305), .Z(n1303) );
XOR2_X1 U998 ( .A(n1306), .B(n1307), .Z(n1305) );
NOR2_X1 U999 ( .A1(KEYINPUT44), .A2(n1275), .ZN(n1307) );
XNOR2_X1 U1000 ( .A(n1126), .B(n1308), .ZN(n1275) );
XOR2_X1 U1001 ( .A(KEYINPUT5), .B(n1127), .Z(n1308) );
XOR2_X1 U1002 ( .A(G131), .B(KEYINPUT15), .Z(n1127) );
XNOR2_X1 U1003 ( .A(G137), .B(G134), .ZN(n1126) );
NOR2_X1 U1004 ( .A1(n1204), .A2(n1309), .ZN(n1306) );
NOR2_X1 U1005 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NOR2_X1 U1006 ( .A1(G953), .A2(n1312), .ZN(n1310) );
NOR3_X1 U1007 ( .A1(n1202), .A2(G953), .A3(n1312), .ZN(n1204) );
INV_X1 U1008 ( .A(G227), .ZN(n1312) );
INV_X1 U1009 ( .A(n1311), .ZN(n1202) );
XOR2_X1 U1010 ( .A(G110), .B(n1132), .Z(n1311) );
XNOR2_X1 U1011 ( .A(n1195), .B(n1313), .ZN(n1304) );
NOR2_X1 U1012 ( .A1(KEYINPUT53), .A2(n1120), .ZN(n1313) );
XNOR2_X1 U1013 ( .A(n1314), .B(n1315), .ZN(n1120) );
NOR2_X1 U1014 ( .A1(KEYINPUT24), .A2(n1316), .ZN(n1315) );
XOR2_X1 U1015 ( .A(G107), .B(n1317), .Z(n1195) );
XNOR2_X1 U1016 ( .A(KEYINPUT20), .B(n1199), .ZN(n1302) );
INV_X1 U1017 ( .A(G469), .ZN(n1199) );
XOR2_X1 U1018 ( .A(n1075), .B(KEYINPUT22), .Z(n1267) );
AND2_X1 U1019 ( .A1(G221), .A2(n1288), .ZN(n1075) );
NAND2_X1 U1020 ( .A1(G234), .A2(n1270), .ZN(n1288) );
NAND2_X1 U1021 ( .A1(n1062), .A2(n1318), .ZN(n1257) );
NAND4_X1 U1022 ( .A1(G953), .A2(G902), .A3(n1256), .A4(n1146), .ZN(n1318) );
INV_X1 U1023 ( .A(G898), .ZN(n1146) );
NAND3_X1 U1024 ( .A1(n1319), .A2(n1256), .A3(G952), .ZN(n1062) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1256) );
INV_X1 U1026 ( .A(n1037), .ZN(n1319) );
XOR2_X1 U1027 ( .A(G953), .B(KEYINPUT40), .Z(n1037) );
NOR2_X1 U1028 ( .A1(n1055), .A2(n1054), .ZN(n1226) );
INV_X1 U1029 ( .A(n1251), .ZN(n1054) );
NAND2_X1 U1030 ( .A1(n1320), .A2(n1321), .ZN(n1251) );
XOR2_X1 U1031 ( .A(KEYINPUT35), .B(G214), .Z(n1320) );
XNOR2_X1 U1032 ( .A(n1088), .B(n1087), .ZN(n1055) );
NAND2_X1 U1033 ( .A1(G210), .A2(n1321), .ZN(n1087) );
NAND2_X1 U1034 ( .A1(n1270), .A2(n1277), .ZN(n1321) );
NAND2_X1 U1035 ( .A1(n1322), .A2(n1270), .ZN(n1088) );
XNOR2_X1 U1036 ( .A(n1323), .B(n1151), .ZN(n1322) );
XOR2_X1 U1037 ( .A(n1324), .B(n1325), .Z(n1151) );
XOR2_X1 U1038 ( .A(n1326), .B(n1327), .Z(n1325) );
XNOR2_X1 U1039 ( .A(n1328), .B(n1329), .ZN(n1327) );
NAND2_X1 U1040 ( .A1(KEYINPUT31), .A2(n1278), .ZN(n1329) );
INV_X1 U1041 ( .A(G113), .ZN(n1278) );
NAND2_X1 U1042 ( .A1(KEYINPUT27), .A2(G110), .ZN(n1328) );
XNOR2_X1 U1043 ( .A(KEYINPUT38), .B(KEYINPUT28), .ZN(n1326) );
XNOR2_X1 U1044 ( .A(n1317), .B(n1330), .ZN(n1324) );
XOR2_X1 U1045 ( .A(n1283), .B(n1331), .Z(n1330) );
XNOR2_X1 U1046 ( .A(G116), .B(n1282), .ZN(n1283) );
INV_X1 U1047 ( .A(G119), .ZN(n1282) );
XOR2_X1 U1048 ( .A(G104), .B(G101), .Z(n1317) );
NAND2_X1 U1049 ( .A1(KEYINPUT47), .A2(n1206), .ZN(n1323) );
XOR2_X1 U1050 ( .A(n1332), .B(n1188), .Z(n1206) );
XNOR2_X1 U1051 ( .A(n1316), .B(n1314), .ZN(n1188) );
XOR2_X1 U1052 ( .A(G143), .B(G146), .Z(n1314) );
INV_X1 U1053 ( .A(G128), .ZN(n1316) );
XNOR2_X1 U1054 ( .A(G125), .B(n1333), .ZN(n1332) );
AND2_X1 U1055 ( .A1(n1114), .A2(G224), .ZN(n1333) );
NOR2_X1 U1056 ( .A1(n1084), .A2(n1258), .ZN(n1043) );
NAND2_X1 U1057 ( .A1(n1079), .A2(n1334), .ZN(n1258) );
OR2_X1 U1058 ( .A1(n1093), .A2(n1094), .ZN(n1334) );
NAND2_X1 U1059 ( .A1(n1094), .A2(n1093), .ZN(n1079) );
INV_X1 U1060 ( .A(G475), .ZN(n1093) );
NOR2_X1 U1061 ( .A1(n1168), .A2(G902), .ZN(n1094) );
XNOR2_X1 U1062 ( .A(n1335), .B(n1336), .ZN(n1168) );
XOR2_X1 U1063 ( .A(n1337), .B(n1338), .Z(n1336) );
XOR2_X1 U1064 ( .A(n1339), .B(n1340), .Z(n1338) );
NOR2_X1 U1065 ( .A1(G143), .A2(KEYINPUT46), .ZN(n1340) );
NAND3_X1 U1066 ( .A1(n1277), .A2(n1114), .A3(G214), .ZN(n1339) );
INV_X1 U1067 ( .A(G237), .ZN(n1277) );
NAND3_X1 U1068 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1337) );
OR2_X1 U1069 ( .A1(n1300), .A2(n1133), .ZN(n1343) );
INV_X1 U1070 ( .A(G125), .ZN(n1133) );
NAND2_X1 U1071 ( .A1(KEYINPUT6), .A2(n1344), .ZN(n1342) );
NAND3_X1 U1072 ( .A1(n1345), .A2(n1346), .A3(n1300), .ZN(n1344) );
NAND2_X1 U1073 ( .A1(G146), .A2(n1132), .ZN(n1300) );
NAND2_X1 U1074 ( .A1(n1134), .A2(n1347), .ZN(n1346) );
NAND2_X1 U1075 ( .A1(G125), .A2(G146), .ZN(n1345) );
NAND2_X1 U1076 ( .A1(n1299), .A2(n1348), .ZN(n1341) );
INV_X1 U1077 ( .A(KEYINPUT6), .ZN(n1348) );
NAND2_X1 U1078 ( .A1(n1349), .A2(n1350), .ZN(n1299) );
NAND2_X1 U1079 ( .A1(n1134), .A2(G146), .ZN(n1350) );
NOR2_X1 U1080 ( .A1(n1132), .A2(G125), .ZN(n1134) );
INV_X1 U1081 ( .A(G140), .ZN(n1132) );
NAND2_X1 U1082 ( .A1(n1351), .A2(n1347), .ZN(n1349) );
INV_X1 U1083 ( .A(G146), .ZN(n1347) );
XNOR2_X1 U1084 ( .A(G140), .B(G125), .ZN(n1351) );
XOR2_X1 U1085 ( .A(n1352), .B(n1353), .Z(n1335) );
XOR2_X1 U1086 ( .A(G131), .B(G122), .Z(n1353) );
XNOR2_X1 U1087 ( .A(G104), .B(G113), .ZN(n1352) );
XNOR2_X1 U1088 ( .A(n1354), .B(G478), .ZN(n1084) );
NAND2_X1 U1089 ( .A1(n1160), .A2(n1270), .ZN(n1354) );
INV_X1 U1090 ( .A(G902), .ZN(n1270) );
XNOR2_X1 U1091 ( .A(n1355), .B(n1356), .ZN(n1160) );
XOR2_X1 U1092 ( .A(n1357), .B(n1358), .Z(n1356) );
XNOR2_X1 U1093 ( .A(n1234), .B(G134), .ZN(n1358) );
INV_X1 U1094 ( .A(G143), .ZN(n1234) );
NOR2_X1 U1095 ( .A1(KEYINPUT34), .A2(G116), .ZN(n1357) );
XOR2_X1 U1096 ( .A(n1359), .B(n1331), .Z(n1355) );
XOR2_X1 U1097 ( .A(G107), .B(G122), .Z(n1331) );
XOR2_X1 U1098 ( .A(n1360), .B(n1361), .Z(n1359) );
NOR2_X1 U1099 ( .A1(G128), .A2(KEYINPUT13), .ZN(n1361) );
NAND2_X1 U1100 ( .A1(G217), .A2(n1295), .ZN(n1360) );
AND2_X1 U1101 ( .A1(G234), .A2(n1114), .ZN(n1295) );
INV_X1 U1102 ( .A(G953), .ZN(n1114) );
endmodule


