//Key = 0100001001001011111110100010001000110111111111111100101011000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377;

XNOR2_X1 U745 ( .A(n1047), .B(n1048), .ZN(G9) );
AND2_X1 U746 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U747 ( .A1(n1051), .A2(n1052), .ZN(G75) );
NOR4_X1 U748 ( .A1(n1053), .A2(n1054), .A3(G953), .A4(n1055), .ZN(n1052) );
NOR4_X1 U749 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1054) );
INV_X1 U750 ( .A(n1060), .ZN(n1057) );
NOR2_X1 U751 ( .A1(n1061), .A2(n1062), .ZN(n1056) );
NOR2_X1 U752 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NAND3_X1 U753 ( .A1(G952), .A2(n1065), .A3(n1066), .ZN(n1053) );
NAND3_X1 U754 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1065) );
NAND4_X1 U755 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1068) );
NAND3_X1 U756 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
NAND2_X1 U757 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NAND2_X1 U758 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
INV_X1 U759 ( .A(KEYINPUT10), .ZN(n1080) );
INV_X1 U760 ( .A(n1081), .ZN(n1077) );
NAND3_X1 U761 ( .A1(n1060), .A2(n1082), .A3(n1083), .ZN(n1072) );
NAND2_X1 U762 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NAND2_X1 U763 ( .A1(n1074), .A2(n1086), .ZN(n1085) );
NAND2_X1 U764 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
OR2_X1 U765 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
INV_X1 U766 ( .A(n1091), .ZN(n1087) );
NAND2_X1 U767 ( .A1(n1092), .A2(n1093), .ZN(n1084) );
NAND2_X1 U768 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U769 ( .A1(KEYINPUT49), .A2(n1096), .ZN(n1095) );
NAND2_X1 U770 ( .A1(KEYINPUT10), .A2(n1097), .ZN(n1071) );
NAND2_X1 U771 ( .A1(n1076), .A2(n1049), .ZN(n1097) );
INV_X1 U772 ( .A(n1098), .ZN(n1049) );
NAND2_X1 U773 ( .A1(n1099), .A2(n1100), .ZN(n1070) );
INV_X1 U774 ( .A(KEYINPUT49), .ZN(n1100) );
NAND3_X1 U775 ( .A1(n1096), .A2(n1060), .A3(n1076), .ZN(n1099) );
INV_X1 U776 ( .A(n1059), .ZN(n1076) );
NAND2_X1 U777 ( .A1(n1083), .A2(n1092), .ZN(n1059) );
INV_X1 U778 ( .A(n1101), .ZN(n1083) );
NOR3_X1 U779 ( .A1(n1102), .A2(G953), .A3(n1055), .ZN(n1051) );
AND4_X1 U780 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1055) );
NOR4_X1 U781 ( .A1(n1107), .A2(n1108), .A3(n1109), .A4(n1110), .ZN(n1106) );
INV_X1 U782 ( .A(n1111), .ZN(n1110) );
NOR2_X1 U783 ( .A1(n1112), .A2(n1113), .ZN(n1108) );
XNOR2_X1 U784 ( .A(KEYINPUT1), .B(n1114), .ZN(n1112) );
NAND3_X1 U785 ( .A1(n1089), .A2(n1115), .A3(n1116), .ZN(n1107) );
NOR3_X1 U786 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1105) );
XNOR2_X1 U787 ( .A(n1120), .B(n1121), .ZN(n1119) );
NAND2_X1 U788 ( .A1(KEYINPUT48), .A2(n1122), .ZN(n1120) );
INV_X1 U789 ( .A(G475), .ZN(n1122) );
XOR2_X1 U790 ( .A(n1123), .B(KEYINPUT14), .Z(n1118) );
NAND2_X1 U791 ( .A1(n1113), .A2(n1114), .ZN(n1123) );
XNOR2_X1 U792 ( .A(KEYINPUT0), .B(n1124), .ZN(n1113) );
XOR2_X1 U793 ( .A(n1125), .B(KEYINPUT17), .Z(n1117) );
XOR2_X1 U794 ( .A(KEYINPUT60), .B(G952), .Z(n1102) );
XOR2_X1 U795 ( .A(n1126), .B(n1127), .Z(G72) );
XOR2_X1 U796 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND2_X1 U797 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND3_X1 U798 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1128) );
XOR2_X1 U799 ( .A(KEYINPUT46), .B(n1135), .Z(n1134) );
NOR2_X1 U800 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
INV_X1 U801 ( .A(n1138), .ZN(n1133) );
NAND2_X1 U802 ( .A1(n1136), .A2(n1137), .ZN(n1132) );
XOR2_X1 U803 ( .A(n1139), .B(n1140), .Z(n1136) );
XNOR2_X1 U804 ( .A(G131), .B(n1141), .ZN(n1139) );
NOR2_X1 U805 ( .A1(n1142), .A2(n1130), .ZN(n1126) );
AND2_X1 U806 ( .A1(G227), .A2(G900), .ZN(n1142) );
XOR2_X1 U807 ( .A(n1143), .B(n1144), .Z(G69) );
XOR2_X1 U808 ( .A(n1145), .B(n1146), .Z(n1144) );
AND2_X1 U809 ( .A1(n1147), .A2(n1130), .ZN(n1146) );
NOR2_X1 U810 ( .A1(n1148), .A2(n1149), .ZN(n1145) );
XNOR2_X1 U811 ( .A(KEYINPUT53), .B(n1150), .ZN(n1149) );
NOR2_X1 U812 ( .A1(n1151), .A2(n1130), .ZN(n1143) );
AND2_X1 U813 ( .A1(G224), .A2(G898), .ZN(n1151) );
NOR2_X1 U814 ( .A1(n1152), .A2(n1153), .ZN(G66) );
XOR2_X1 U815 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR3_X1 U816 ( .A1(n1156), .A2(KEYINPUT36), .A3(n1157), .ZN(n1154) );
NOR2_X1 U817 ( .A1(n1152), .A2(n1158), .ZN(G63) );
XOR2_X1 U818 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND3_X1 U819 ( .A1(n1161), .A2(n1162), .A3(G478), .ZN(n1159) );
OR2_X1 U820 ( .A1(n1163), .A2(KEYINPUT21), .ZN(n1162) );
NAND2_X1 U821 ( .A1(KEYINPUT21), .A2(n1164), .ZN(n1161) );
OR2_X1 U822 ( .A1(G902), .A2(n1066), .ZN(n1164) );
NOR2_X1 U823 ( .A1(n1152), .A2(n1165), .ZN(G60) );
NOR2_X1 U824 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U825 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND2_X1 U826 ( .A1(G475), .A2(n1163), .ZN(n1169) );
NAND2_X1 U827 ( .A1(n1170), .A2(n1171), .ZN(n1168) );
NOR2_X1 U828 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
INV_X1 U829 ( .A(KEYINPUT8), .ZN(n1171) );
XNOR2_X1 U830 ( .A(G104), .B(n1172), .ZN(G6) );
NOR2_X1 U831 ( .A1(n1152), .A2(n1173), .ZN(G57) );
XOR2_X1 U832 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U833 ( .A(n1176), .B(KEYINPUT40), .Z(n1175) );
NAND2_X1 U834 ( .A1(n1163), .A2(G472), .ZN(n1176) );
NOR2_X1 U835 ( .A1(n1152), .A2(n1177), .ZN(G54) );
XOR2_X1 U836 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U837 ( .A(n1180), .B(n1181), .Z(n1179) );
XNOR2_X1 U838 ( .A(n1182), .B(n1183), .ZN(n1181) );
NOR2_X1 U839 ( .A1(KEYINPUT24), .A2(n1184), .ZN(n1183) );
XOR2_X1 U840 ( .A(n1185), .B(n1186), .Z(n1178) );
XOR2_X1 U841 ( .A(G140), .B(n1187), .Z(n1186) );
NOR2_X1 U842 ( .A1(G110), .A2(KEYINPUT28), .ZN(n1187) );
NAND2_X1 U843 ( .A1(n1163), .A2(G469), .ZN(n1185) );
NOR2_X1 U844 ( .A1(n1152), .A2(n1188), .ZN(G51) );
XOR2_X1 U845 ( .A(n1189), .B(n1190), .Z(n1188) );
OR2_X1 U846 ( .A1(n1156), .A2(n1114), .ZN(n1190) );
INV_X1 U847 ( .A(n1163), .ZN(n1156) );
NOR2_X1 U848 ( .A1(n1191), .A2(n1066), .ZN(n1163) );
NOR2_X1 U849 ( .A1(n1147), .A2(n1131), .ZN(n1066) );
NAND4_X1 U850 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1131) );
NOR3_X1 U851 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1195) );
NAND2_X1 U852 ( .A1(n1062), .A2(n1199), .ZN(n1194) );
NAND2_X1 U853 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XNOR2_X1 U854 ( .A(KEYINPUT18), .B(n1202), .ZN(n1200) );
NAND2_X1 U855 ( .A1(n1203), .A2(n1204), .ZN(n1192) );
NAND2_X1 U856 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NAND2_X1 U857 ( .A1(n1207), .A2(n1079), .ZN(n1206) );
XNOR2_X1 U858 ( .A(KEYINPUT34), .B(n1096), .ZN(n1207) );
NAND2_X1 U859 ( .A1(n1208), .A2(n1081), .ZN(n1205) );
NAND4_X1 U860 ( .A1(n1172), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1147) );
AND4_X1 U861 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1211) );
NOR2_X1 U862 ( .A1(n1216), .A2(n1217), .ZN(n1210) );
NOR2_X1 U863 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NOR3_X1 U864 ( .A1(n1098), .A2(n1220), .A3(n1221), .ZN(n1216) );
NOR2_X1 U865 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
INV_X1 U866 ( .A(KEYINPUT4), .ZN(n1223) );
NOR3_X1 U867 ( .A1(n1224), .A2(n1225), .A3(n1062), .ZN(n1222) );
NOR2_X1 U868 ( .A1(KEYINPUT4), .A2(n1050), .ZN(n1220) );
NAND2_X1 U869 ( .A1(n1079), .A2(n1074), .ZN(n1098) );
NAND3_X1 U870 ( .A1(n1050), .A2(n1074), .A3(n1081), .ZN(n1172) );
NAND3_X1 U871 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1189) );
NAND2_X1 U872 ( .A1(KEYINPUT50), .A2(n1229), .ZN(n1228) );
NAND3_X1 U873 ( .A1(n1230), .A2(n1231), .A3(n1150), .ZN(n1227) );
INV_X1 U874 ( .A(n1232), .ZN(n1150) );
NAND2_X1 U875 ( .A1(n1232), .A2(n1233), .ZN(n1226) );
NAND2_X1 U876 ( .A1(n1234), .A2(n1231), .ZN(n1233) );
INV_X1 U877 ( .A(KEYINPUT50), .ZN(n1231) );
XNOR2_X1 U878 ( .A(KEYINPUT7), .B(n1229), .ZN(n1234) );
INV_X1 U879 ( .A(n1230), .ZN(n1229) );
XNOR2_X1 U880 ( .A(n1235), .B(n1236), .ZN(n1230) );
NAND2_X1 U881 ( .A1(KEYINPUT12), .A2(n1237), .ZN(n1235) );
NOR2_X1 U882 ( .A1(n1130), .A2(G952), .ZN(n1152) );
XOR2_X1 U883 ( .A(G146), .B(n1196), .Z(G48) );
AND4_X1 U884 ( .A1(n1238), .A2(n1081), .A3(n1239), .A4(n1062), .ZN(n1196) );
AND2_X1 U885 ( .A1(n1240), .A2(n1091), .ZN(n1239) );
XNOR2_X1 U886 ( .A(G143), .B(n1193), .ZN(G45) );
NAND4_X1 U887 ( .A1(n1096), .A2(n1240), .A3(n1091), .A4(n1241), .ZN(n1193) );
NOR3_X1 U888 ( .A1(n1242), .A2(n1218), .A3(n1243), .ZN(n1241) );
XOR2_X1 U889 ( .A(G140), .B(n1244), .Z(G42) );
NOR3_X1 U890 ( .A1(n1245), .A2(n1246), .A3(n1094), .ZN(n1244) );
INV_X1 U891 ( .A(n1208), .ZN(n1094) );
XNOR2_X1 U892 ( .A(n1081), .B(KEYINPUT51), .ZN(n1246) );
XOR2_X1 U893 ( .A(G137), .B(n1198), .Z(G39) );
AND3_X1 U894 ( .A1(n1238), .A2(n1060), .A3(n1203), .ZN(n1198) );
XOR2_X1 U895 ( .A(G134), .B(n1247), .Z(G36) );
NOR2_X1 U896 ( .A1(n1248), .A2(n1245), .ZN(n1247) );
XNOR2_X1 U897 ( .A(n1249), .B(n1197), .ZN(G33) );
AND3_X1 U898 ( .A1(n1081), .A2(n1096), .A3(n1203), .ZN(n1197) );
INV_X1 U899 ( .A(n1245), .ZN(n1203) );
NAND4_X1 U900 ( .A1(n1069), .A2(n1067), .A3(n1091), .A4(n1240), .ZN(n1245) );
XOR2_X1 U901 ( .A(n1250), .B(KEYINPUT29), .Z(n1091) );
XNOR2_X1 U902 ( .A(n1063), .B(KEYINPUT63), .ZN(n1067) );
NAND2_X1 U903 ( .A1(n1251), .A2(n1252), .ZN(G30) );
OR2_X1 U904 ( .A1(G128), .A2(KEYINPUT57), .ZN(n1252) );
XOR2_X1 U905 ( .A(n1253), .B(n1254), .Z(n1251) );
NOR2_X1 U906 ( .A1(n1218), .A2(n1202), .ZN(n1254) );
NAND4_X1 U907 ( .A1(n1238), .A2(n1079), .A3(n1250), .A4(n1240), .ZN(n1202) );
INV_X1 U908 ( .A(n1224), .ZN(n1250) );
NAND2_X1 U909 ( .A1(KEYINPUT57), .A2(G128), .ZN(n1253) );
XNOR2_X1 U910 ( .A(G101), .B(n1212), .ZN(G3) );
NAND3_X1 U911 ( .A1(n1096), .A2(n1060), .A3(n1050), .ZN(n1212) );
XNOR2_X1 U912 ( .A(n1255), .B(n1256), .ZN(G27) );
NOR2_X1 U913 ( .A1(n1257), .A2(n1218), .ZN(n1256) );
XOR2_X1 U914 ( .A(n1201), .B(KEYINPUT55), .Z(n1257) );
NAND4_X1 U915 ( .A1(n1092), .A2(n1208), .A3(n1081), .A4(n1240), .ZN(n1201) );
NAND2_X1 U916 ( .A1(n1101), .A2(n1258), .ZN(n1240) );
NAND3_X1 U917 ( .A1(G902), .A2(n1259), .A3(n1138), .ZN(n1258) );
NOR2_X1 U918 ( .A1(n1260), .A2(G900), .ZN(n1138) );
XNOR2_X1 U919 ( .A(G122), .B(n1209), .ZN(G24) );
NAND4_X1 U920 ( .A1(n1261), .A2(n1074), .A3(n1262), .A4(n1263), .ZN(n1209) );
INV_X1 U921 ( .A(n1058), .ZN(n1074) );
NAND2_X1 U922 ( .A1(n1264), .A2(n1265), .ZN(n1058) );
XNOR2_X1 U923 ( .A(n1104), .B(n1266), .ZN(n1264) );
XNOR2_X1 U924 ( .A(G119), .B(n1267), .ZN(G21) );
NAND2_X1 U925 ( .A1(n1268), .A2(n1062), .ZN(n1267) );
XOR2_X1 U926 ( .A(n1219), .B(KEYINPUT19), .Z(n1268) );
NAND4_X1 U927 ( .A1(n1092), .A2(n1238), .A3(n1060), .A4(n1269), .ZN(n1219) );
NAND2_X1 U928 ( .A1(n1270), .A2(n1271), .ZN(G18) );
NAND2_X1 U929 ( .A1(G116), .A2(n1215), .ZN(n1271) );
XOR2_X1 U930 ( .A(KEYINPUT9), .B(n1272), .Z(n1270) );
NOR2_X1 U931 ( .A1(G116), .A2(n1215), .ZN(n1272) );
OR2_X1 U932 ( .A1(n1248), .A2(n1273), .ZN(n1215) );
NAND2_X1 U933 ( .A1(n1079), .A2(n1096), .ZN(n1248) );
AND2_X1 U934 ( .A1(n1262), .A2(n1274), .ZN(n1079) );
XNOR2_X1 U935 ( .A(KEYINPUT3), .B(n1263), .ZN(n1274) );
XNOR2_X1 U936 ( .A(G113), .B(n1214), .ZN(G15) );
NAND3_X1 U937 ( .A1(n1081), .A2(n1096), .A3(n1261), .ZN(n1214) );
INV_X1 U938 ( .A(n1273), .ZN(n1261) );
NAND3_X1 U939 ( .A1(n1062), .A2(n1269), .A3(n1092), .ZN(n1273) );
NOR2_X1 U940 ( .A1(n1090), .A2(n1275), .ZN(n1092) );
INV_X1 U941 ( .A(n1089), .ZN(n1275) );
NAND2_X1 U942 ( .A1(n1276), .A2(n1277), .ZN(n1096) );
NAND3_X1 U943 ( .A1(n1104), .A2(n1278), .A3(n1266), .ZN(n1277) );
INV_X1 U944 ( .A(KEYINPUT33), .ZN(n1266) );
NAND2_X1 U945 ( .A1(KEYINPUT33), .A2(n1238), .ZN(n1276) );
NOR2_X1 U946 ( .A1(n1104), .A2(n1265), .ZN(n1238) );
INV_X1 U947 ( .A(n1278), .ZN(n1265) );
NAND2_X1 U948 ( .A1(n1279), .A2(n1280), .ZN(G12) );
NAND2_X1 U949 ( .A1(G110), .A2(n1213), .ZN(n1280) );
XOR2_X1 U950 ( .A(KEYINPUT43), .B(n1281), .Z(n1279) );
NOR2_X1 U951 ( .A1(G110), .A2(n1213), .ZN(n1281) );
NAND3_X1 U952 ( .A1(n1050), .A2(n1060), .A3(n1208), .ZN(n1213) );
NOR2_X1 U953 ( .A1(n1278), .A2(n1104), .ZN(n1208) );
XNOR2_X1 U954 ( .A(n1282), .B(n1157), .ZN(n1104) );
NAND2_X1 U955 ( .A1(G217), .A2(n1283), .ZN(n1157) );
OR2_X1 U956 ( .A1(n1155), .A2(n1284), .ZN(n1282) );
INV_X1 U957 ( .A(n1285), .ZN(n1284) );
XNOR2_X1 U958 ( .A(n1286), .B(n1287), .ZN(n1155) );
XOR2_X1 U959 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U960 ( .A(G140), .B(G137), .Z(n1289) );
XOR2_X1 U961 ( .A(KEYINPUT5), .B(KEYINPUT27), .Z(n1288) );
XOR2_X1 U962 ( .A(n1290), .B(n1291), .Z(n1286) );
XOR2_X1 U963 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U964 ( .A(n1294), .B(n1295), .Z(n1290) );
AND3_X1 U965 ( .A1(G221), .A2(n1130), .A3(G234), .ZN(n1295) );
NAND2_X1 U966 ( .A1(KEYINPUT54), .A2(n1255), .ZN(n1294) );
NAND2_X1 U967 ( .A1(n1125), .A2(n1111), .ZN(n1278) );
NAND2_X1 U968 ( .A1(G472), .A2(n1296), .ZN(n1111) );
OR2_X1 U969 ( .A1(n1296), .A2(G472), .ZN(n1125) );
NAND2_X1 U970 ( .A1(n1297), .A2(n1285), .ZN(n1296) );
XOR2_X1 U971 ( .A(n1174), .B(n1298), .Z(n1297) );
XOR2_X1 U972 ( .A(KEYINPUT52), .B(KEYINPUT31), .Z(n1298) );
XOR2_X1 U973 ( .A(n1299), .B(n1300), .Z(n1174) );
XOR2_X1 U974 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U975 ( .A(n1303), .B(n1304), .Z(n1302) );
NAND2_X1 U976 ( .A1(KEYINPUT41), .A2(n1305), .ZN(n1304) );
NAND2_X1 U977 ( .A1(n1306), .A2(G210), .ZN(n1303) );
XOR2_X1 U978 ( .A(KEYINPUT58), .B(G119), .Z(n1301) );
XNOR2_X1 U979 ( .A(n1307), .B(n1308), .ZN(n1299) );
INV_X1 U980 ( .A(n1182), .ZN(n1308) );
XNOR2_X1 U981 ( .A(n1309), .B(n1310), .ZN(n1307) );
INV_X1 U982 ( .A(n1311), .ZN(n1310) );
NAND2_X1 U983 ( .A1(n1312), .A2(n1313), .ZN(n1060) );
OR3_X1 U984 ( .A1(n1263), .A2(n1262), .A3(KEYINPUT3), .ZN(n1313) );
INV_X1 U985 ( .A(n1243), .ZN(n1263) );
NAND2_X1 U986 ( .A1(KEYINPUT3), .A2(n1081), .ZN(n1312) );
NOR2_X1 U987 ( .A1(n1243), .A2(n1262), .ZN(n1081) );
INV_X1 U988 ( .A(n1242), .ZN(n1262) );
XNOR2_X1 U989 ( .A(n1103), .B(KEYINPUT47), .ZN(n1242) );
XOR2_X1 U990 ( .A(n1314), .B(G478), .Z(n1103) );
NAND2_X1 U991 ( .A1(n1160), .A2(n1285), .ZN(n1314) );
XNOR2_X1 U992 ( .A(n1315), .B(n1316), .ZN(n1160) );
NOR3_X1 U993 ( .A1(n1317), .A2(G953), .A3(n1318), .ZN(n1316) );
INV_X1 U994 ( .A(G217), .ZN(n1318) );
XOR2_X1 U995 ( .A(KEYINPUT6), .B(G234), .Z(n1317) );
NAND2_X1 U996 ( .A1(KEYINPUT42), .A2(n1319), .ZN(n1315) );
XOR2_X1 U997 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U998 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U999 ( .A(n1324), .B(n1325), .Z(n1322) );
NAND2_X1 U1000 ( .A1(KEYINPUT26), .A2(G128), .ZN(n1324) );
XNOR2_X1 U1001 ( .A(G134), .B(n1326), .ZN(n1320) );
XOR2_X1 U1002 ( .A(KEYINPUT45), .B(G143), .Z(n1326) );
XNOR2_X1 U1003 ( .A(n1121), .B(n1327), .ZN(n1243) );
NOR2_X1 U1004 ( .A1(G475), .A2(KEYINPUT23), .ZN(n1327) );
NAND2_X1 U1005 ( .A1(n1170), .A2(n1285), .ZN(n1121) );
XOR2_X1 U1006 ( .A(n1328), .B(n1329), .Z(n1170) );
XOR2_X1 U1007 ( .A(n1330), .B(n1331), .Z(n1329) );
NAND2_X1 U1008 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
NAND2_X1 U1009 ( .A1(G113), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1010 ( .A(KEYINPUT35), .B(n1335), .Z(n1332) );
NOR2_X1 U1011 ( .A1(G113), .A2(n1334), .ZN(n1335) );
INV_X1 U1012 ( .A(G122), .ZN(n1334) );
NAND3_X1 U1013 ( .A1(n1336), .A2(n1337), .A3(n1338), .ZN(n1330) );
NAND2_X1 U1014 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
INV_X1 U1015 ( .A(KEYINPUT37), .ZN(n1340) );
NAND3_X1 U1016 ( .A1(KEYINPUT37), .A2(n1341), .A3(n1342), .ZN(n1337) );
OR2_X1 U1017 ( .A1(n1342), .A2(n1341), .ZN(n1336) );
NOR2_X1 U1018 ( .A1(n1339), .A2(KEYINPUT11), .ZN(n1341) );
AND2_X1 U1019 ( .A1(n1343), .A2(n1344), .ZN(n1339) );
NAND2_X1 U1020 ( .A1(G146), .A2(n1137), .ZN(n1344) );
XOR2_X1 U1021 ( .A(KEYINPUT22), .B(n1345), .Z(n1343) );
NOR2_X1 U1022 ( .A1(G146), .A2(n1137), .ZN(n1345) );
XNOR2_X1 U1023 ( .A(n1255), .B(G140), .ZN(n1137) );
XNOR2_X1 U1024 ( .A(n1346), .B(n1347), .ZN(n1342) );
XNOR2_X1 U1025 ( .A(G143), .B(n1249), .ZN(n1347) );
NAND2_X1 U1026 ( .A1(n1306), .A2(G214), .ZN(n1346) );
NOR2_X1 U1027 ( .A1(G953), .A2(G237), .ZN(n1306) );
XNOR2_X1 U1028 ( .A(G104), .B(KEYINPUT30), .ZN(n1328) );
NOR3_X1 U1029 ( .A1(n1218), .A2(n1225), .A3(n1224), .ZN(n1050) );
NAND2_X1 U1030 ( .A1(n1089), .A2(n1090), .ZN(n1224) );
NAND2_X1 U1031 ( .A1(n1348), .A2(n1116), .ZN(n1090) );
OR2_X1 U1032 ( .A1(n1349), .A2(G469), .ZN(n1116) );
XOR2_X1 U1033 ( .A(n1115), .B(KEYINPUT2), .Z(n1348) );
NAND2_X1 U1034 ( .A1(G469), .A2(n1349), .ZN(n1115) );
NAND2_X1 U1035 ( .A1(n1350), .A2(n1285), .ZN(n1349) );
XOR2_X1 U1036 ( .A(n1351), .B(n1352), .Z(n1350) );
XNOR2_X1 U1037 ( .A(n1353), .B(n1354), .ZN(n1352) );
NOR2_X1 U1038 ( .A1(KEYINPUT59), .A2(n1355), .ZN(n1354) );
XNOR2_X1 U1039 ( .A(G110), .B(n1356), .ZN(n1355) );
XOR2_X1 U1040 ( .A(KEYINPUT25), .B(G140), .Z(n1356) );
NAND2_X1 U1041 ( .A1(KEYINPUT56), .A2(n1182), .ZN(n1353) );
XOR2_X1 U1042 ( .A(n1357), .B(n1249), .Z(n1182) );
INV_X1 U1043 ( .A(G131), .ZN(n1249) );
NAND2_X1 U1044 ( .A1(KEYINPUT61), .A2(n1141), .ZN(n1357) );
XOR2_X1 U1045 ( .A(G134), .B(G137), .Z(n1141) );
XNOR2_X1 U1046 ( .A(n1180), .B(n1184), .ZN(n1351) );
NAND2_X1 U1047 ( .A1(G227), .A2(n1130), .ZN(n1184) );
XNOR2_X1 U1048 ( .A(n1140), .B(n1358), .ZN(n1180) );
XNOR2_X1 U1049 ( .A(G101), .B(n1359), .ZN(n1358) );
NAND2_X1 U1050 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NAND2_X1 U1051 ( .A1(G107), .A2(n1362), .ZN(n1361) );
XNOR2_X1 U1052 ( .A(KEYINPUT38), .B(n1363), .ZN(n1362) );
XOR2_X1 U1053 ( .A(n1364), .B(KEYINPUT13), .Z(n1360) );
NAND2_X1 U1054 ( .A1(n1365), .A2(n1047), .ZN(n1364) );
XNOR2_X1 U1055 ( .A(G104), .B(KEYINPUT62), .ZN(n1365) );
XNOR2_X1 U1056 ( .A(n1366), .B(G128), .ZN(n1140) );
NAND2_X1 U1057 ( .A1(KEYINPUT44), .A2(n1367), .ZN(n1366) );
XOR2_X1 U1058 ( .A(G146), .B(G143), .Z(n1367) );
NAND2_X1 U1059 ( .A1(G221), .A2(n1283), .ZN(n1089) );
NAND2_X1 U1060 ( .A1(G234), .A2(n1191), .ZN(n1283) );
INV_X1 U1061 ( .A(n1269), .ZN(n1225) );
NAND2_X1 U1062 ( .A1(n1101), .A2(n1368), .ZN(n1269) );
NAND3_X1 U1063 ( .A1(G902), .A2(n1259), .A3(n1148), .ZN(n1368) );
NOR2_X1 U1064 ( .A1(n1260), .A2(G898), .ZN(n1148) );
XNOR2_X1 U1065 ( .A(G953), .B(KEYINPUT32), .ZN(n1260) );
NAND3_X1 U1066 ( .A1(n1259), .A2(n1130), .A3(G952), .ZN(n1101) );
NAND2_X1 U1067 ( .A1(G237), .A2(G234), .ZN(n1259) );
INV_X1 U1068 ( .A(n1062), .ZN(n1218) );
NOR2_X1 U1069 ( .A1(n1069), .A2(n1109), .ZN(n1062) );
INV_X1 U1070 ( .A(n1063), .ZN(n1109) );
NAND2_X1 U1071 ( .A1(G214), .A2(n1369), .ZN(n1063) );
INV_X1 U1072 ( .A(n1064), .ZN(n1069) );
XOR2_X1 U1073 ( .A(n1124), .B(n1114), .Z(n1064) );
NAND2_X1 U1074 ( .A1(G210), .A2(n1369), .ZN(n1114) );
NAND2_X1 U1075 ( .A1(n1370), .A2(n1191), .ZN(n1369) );
INV_X1 U1076 ( .A(G902), .ZN(n1191) );
INV_X1 U1077 ( .A(G237), .ZN(n1370) );
NAND2_X1 U1078 ( .A1(n1371), .A2(n1372), .ZN(n1124) );
XNOR2_X1 U1079 ( .A(n1232), .B(n1373), .ZN(n1372) );
XNOR2_X1 U1080 ( .A(n1236), .B(n1237), .ZN(n1373) );
AND2_X1 U1081 ( .A1(G224), .A2(n1130), .ZN(n1237) );
INV_X1 U1082 ( .A(G953), .ZN(n1130) );
XNOR2_X1 U1083 ( .A(n1311), .B(n1255), .ZN(n1236) );
INV_X1 U1084 ( .A(G125), .ZN(n1255) );
XOR2_X1 U1085 ( .A(G143), .B(n1292), .Z(n1311) );
XOR2_X1 U1086 ( .A(G128), .B(G146), .Z(n1292) );
XNOR2_X1 U1087 ( .A(n1374), .B(n1375), .ZN(n1232) );
XNOR2_X1 U1088 ( .A(n1363), .B(n1376), .ZN(n1375) );
XNOR2_X1 U1089 ( .A(KEYINPUT20), .B(n1305), .ZN(n1376) );
INV_X1 U1090 ( .A(G113), .ZN(n1305) );
INV_X1 U1091 ( .A(G104), .ZN(n1363) );
XOR2_X1 U1092 ( .A(n1377), .B(n1323), .Z(n1374) );
XNOR2_X1 U1093 ( .A(n1047), .B(G122), .ZN(n1323) );
INV_X1 U1094 ( .A(G107), .ZN(n1047) );
XOR2_X1 U1095 ( .A(n1309), .B(n1293), .Z(n1377) );
XOR2_X1 U1096 ( .A(G119), .B(G110), .Z(n1293) );
XNOR2_X1 U1097 ( .A(G101), .B(n1325), .ZN(n1309) );
XOR2_X1 U1098 ( .A(G116), .B(KEYINPUT39), .Z(n1325) );
XNOR2_X1 U1099 ( .A(n1285), .B(KEYINPUT16), .ZN(n1371) );
XOR2_X1 U1100 ( .A(G902), .B(KEYINPUT15), .Z(n1285) );
endmodule


