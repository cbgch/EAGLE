//Key = 1100010110011100110011001101011110111010011001110100000001011011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383;

XNOR2_X1 U753 ( .A(n1042), .B(n1043), .ZN(G9) );
NOR2_X1 U754 ( .A1(n1044), .A2(n1045), .ZN(G75) );
NOR3_X1 U755 ( .A1(n1046), .A2(G952), .A3(n1047), .ZN(n1045) );
INV_X1 U756 ( .A(n1048), .ZN(n1047) );
NOR4_X1 U757 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1046), .ZN(n1044) );
NAND4_X1 U758 ( .A1(n1052), .A2(n1053), .A3(n1048), .A4(n1054), .ZN(n1049) );
NAND2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND3_X1 U760 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
NAND2_X1 U761 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
OR2_X1 U762 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND3_X1 U763 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1058) );
NAND2_X1 U764 ( .A1(n1067), .A2(n1068), .ZN(n1057) );
INV_X1 U765 ( .A(KEYINPUT52), .ZN(n1068) );
NAND4_X1 U766 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1048) );
NOR4_X1 U767 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1072) );
XOR2_X1 U768 ( .A(KEYINPUT33), .B(n1077), .Z(n1076) );
AND2_X1 U769 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XNOR2_X1 U770 ( .A(G475), .B(n1080), .ZN(n1075) );
XNOR2_X1 U771 ( .A(n1081), .B(n1082), .ZN(n1074) );
NOR2_X1 U772 ( .A1(n1083), .A2(n1084), .ZN(n1071) );
NAND4_X1 U773 ( .A1(n1085), .A2(n1060), .A3(n1066), .A4(n1086), .ZN(n1053) );
NAND2_X1 U774 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U775 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U776 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U777 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U778 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U779 ( .A1(n1084), .A2(n1097), .ZN(n1096) );
NAND2_X1 U780 ( .A1(n1098), .A2(n1099), .ZN(n1091) );
NAND2_X1 U781 ( .A1(n1100), .A2(n1098), .ZN(n1087) );
NAND2_X1 U782 ( .A1(KEYINPUT52), .A2(n1101), .ZN(n1052) );
NAND2_X1 U783 ( .A1(n1055), .A2(n1067), .ZN(n1101) );
AND4_X1 U784 ( .A1(n1085), .A2(n1098), .A3(n1093), .A4(n1089), .ZN(n1055) );
NAND2_X1 U785 ( .A1(n1102), .A2(n1103), .ZN(G72) );
NAND3_X1 U786 ( .A1(G953), .A2(n1104), .A3(n1105), .ZN(n1103) );
XOR2_X1 U787 ( .A(KEYINPUT5), .B(n1106), .Z(n1102) );
NOR2_X1 U788 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U789 ( .A(n1105), .B(KEYINPUT60), .ZN(n1108) );
AND2_X1 U790 ( .A1(n1109), .A2(n1110), .ZN(n1105) );
NAND2_X1 U791 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U792 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NAND2_X1 U793 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U794 ( .A1(G900), .A2(G953), .ZN(n1113) );
OR3_X1 U795 ( .A1(n1115), .A2(G953), .A3(n1112), .ZN(n1109) );
XNOR2_X1 U796 ( .A(n1117), .B(n1118), .ZN(n1112) );
XNOR2_X1 U797 ( .A(n1119), .B(KEYINPUT44), .ZN(n1118) );
NAND2_X1 U798 ( .A1(n1120), .A2(KEYINPUT35), .ZN(n1119) );
XOR2_X1 U799 ( .A(n1121), .B(n1122), .Z(n1120) );
XNOR2_X1 U800 ( .A(G131), .B(KEYINPUT58), .ZN(n1121) );
NAND2_X1 U801 ( .A1(n1123), .A2(n1124), .ZN(n1117) );
NAND2_X1 U802 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
OR2_X1 U803 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
INV_X1 U804 ( .A(n1129), .ZN(n1125) );
NAND2_X1 U805 ( .A1(n1130), .A2(n1129), .ZN(n1123) );
XNOR2_X1 U806 ( .A(n1131), .B(G125), .ZN(n1130) );
INV_X1 U807 ( .A(n1051), .ZN(n1115) );
AND2_X1 U808 ( .A1(n1104), .A2(G953), .ZN(n1107) );
NAND2_X1 U809 ( .A1(G900), .A2(G227), .ZN(n1104) );
XOR2_X1 U810 ( .A(n1132), .B(n1133), .Z(G69) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U812 ( .A1(n1136), .A2(n1116), .ZN(n1135) );
NOR2_X1 U813 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND3_X1 U814 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1134) );
XOR2_X1 U815 ( .A(n1142), .B(KEYINPUT43), .Z(n1141) );
NAND2_X1 U816 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
OR2_X1 U817 ( .A1(n1144), .A2(n1143), .ZN(n1140) );
NAND2_X1 U818 ( .A1(G953), .A2(n1138), .ZN(n1139) );
INV_X1 U819 ( .A(G898), .ZN(n1138) );
NAND2_X1 U820 ( .A1(n1116), .A2(n1050), .ZN(n1132) );
NOR2_X1 U821 ( .A1(n1145), .A2(n1146), .ZN(G66) );
XOR2_X1 U822 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U823 ( .A(n1149), .B(KEYINPUT40), .Z(n1147) );
NAND2_X1 U824 ( .A1(n1150), .A2(n1082), .ZN(n1149) );
INV_X1 U825 ( .A(n1151), .ZN(n1082) );
NOR2_X1 U826 ( .A1(n1145), .A2(n1152), .ZN(G63) );
NOR3_X1 U827 ( .A1(n1079), .A2(n1153), .A3(n1154), .ZN(n1152) );
AND3_X1 U828 ( .A1(n1155), .A2(G478), .A3(n1150), .ZN(n1154) );
NOR2_X1 U829 ( .A1(n1156), .A2(n1155), .ZN(n1153) );
NOR2_X1 U830 ( .A1(n1157), .A2(n1078), .ZN(n1156) );
NOR2_X1 U831 ( .A1(n1051), .A2(n1050), .ZN(n1157) );
NOR2_X1 U832 ( .A1(n1145), .A2(n1158), .ZN(G60) );
XOR2_X1 U833 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND2_X1 U834 ( .A1(n1150), .A2(G475), .ZN(n1159) );
XOR2_X1 U835 ( .A(G104), .B(n1161), .Z(G6) );
NOR2_X1 U836 ( .A1(n1145), .A2(n1162), .ZN(G57) );
XOR2_X1 U837 ( .A(n1163), .B(KEYINPUT63), .Z(n1162) );
NAND3_X1 U838 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1163) );
NAND2_X1 U839 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND2_X1 U840 ( .A1(n1169), .A2(n1170), .ZN(n1165) );
INV_X1 U841 ( .A(KEYINPUT27), .ZN(n1170) );
NAND2_X1 U842 ( .A1(n1171), .A2(n1172), .ZN(n1169) );
XNOR2_X1 U843 ( .A(n1173), .B(n1167), .ZN(n1171) );
NAND2_X1 U844 ( .A1(KEYINPUT27), .A2(n1174), .ZN(n1164) );
NAND2_X1 U845 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND2_X1 U846 ( .A1(n1167), .A2(n1173), .ZN(n1176) );
OR3_X1 U847 ( .A1(n1168), .A2(n1167), .A3(n1173), .ZN(n1175) );
INV_X1 U848 ( .A(KEYINPUT0), .ZN(n1173) );
XNOR2_X1 U849 ( .A(n1177), .B(n1178), .ZN(n1167) );
NOR2_X1 U850 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NOR2_X1 U851 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U852 ( .A(n1183), .B(KEYINPUT41), .Z(n1182) );
NOR2_X1 U853 ( .A1(n1184), .A2(n1183), .ZN(n1179) );
INV_X1 U854 ( .A(n1181), .ZN(n1184) );
NAND2_X1 U855 ( .A1(n1150), .A2(G472), .ZN(n1177) );
INV_X1 U856 ( .A(n1172), .ZN(n1168) );
NOR2_X1 U857 ( .A1(n1185), .A2(n1186), .ZN(n1172) );
NOR2_X1 U858 ( .A1(G101), .A2(n1187), .ZN(n1185) );
NOR2_X1 U859 ( .A1(n1188), .A2(n1189), .ZN(G54) );
XOR2_X1 U860 ( .A(n1190), .B(n1191), .Z(n1189) );
XNOR2_X1 U861 ( .A(n1192), .B(n1193), .ZN(n1191) );
NOR2_X1 U862 ( .A1(KEYINPUT3), .A2(n1194), .ZN(n1193) );
NOR2_X1 U863 ( .A1(KEYINPUT18), .A2(n1195), .ZN(n1192) );
XNOR2_X1 U864 ( .A(n1196), .B(n1197), .ZN(n1190) );
NAND2_X1 U865 ( .A1(n1150), .A2(G469), .ZN(n1196) );
XNOR2_X1 U866 ( .A(n1145), .B(KEYINPUT7), .ZN(n1188) );
NOR2_X1 U867 ( .A1(n1145), .A2(n1198), .ZN(G51) );
XOR2_X1 U868 ( .A(n1199), .B(n1200), .Z(n1198) );
XOR2_X1 U869 ( .A(n1201), .B(n1202), .Z(n1199) );
NAND2_X1 U870 ( .A1(n1150), .A2(n1203), .ZN(n1201) );
AND2_X1 U871 ( .A1(G902), .A2(n1204), .ZN(n1150) );
OR2_X1 U872 ( .A1(n1050), .A2(n1051), .ZN(n1204) );
NAND4_X1 U873 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1051) );
NOR4_X1 U874 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1208) );
NOR2_X1 U875 ( .A1(n1213), .A2(n1214), .ZN(n1207) );
INV_X1 U876 ( .A(n1215), .ZN(n1213) );
NAND3_X1 U877 ( .A1(n1060), .A2(n1216), .A3(n1217), .ZN(n1206) );
NAND2_X1 U878 ( .A1(n1218), .A2(n1098), .ZN(n1205) );
XOR2_X1 U879 ( .A(n1219), .B(KEYINPUT16), .Z(n1218) );
NAND4_X1 U880 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1050) );
NOR4_X1 U881 ( .A1(n1224), .A2(n1043), .A3(n1225), .A4(n1226), .ZN(n1223) );
AND3_X1 U882 ( .A1(n1093), .A2(n1227), .A3(n1063), .ZN(n1043) );
INV_X1 U883 ( .A(n1228), .ZN(n1224) );
NOR2_X1 U884 ( .A1(n1229), .A2(n1161), .ZN(n1222) );
AND3_X1 U885 ( .A1(n1093), .A2(n1227), .A3(n1062), .ZN(n1161) );
INV_X1 U886 ( .A(n1230), .ZN(n1229) );
NOR2_X1 U887 ( .A1(n1116), .A2(G952), .ZN(n1145) );
NAND2_X1 U888 ( .A1(n1231), .A2(n1232), .ZN(G48) );
NAND2_X1 U889 ( .A1(n1211), .A2(n1233), .ZN(n1232) );
XOR2_X1 U890 ( .A(KEYINPUT11), .B(n1234), .Z(n1231) );
NOR2_X1 U891 ( .A1(n1211), .A2(n1233), .ZN(n1234) );
AND3_X1 U892 ( .A1(n1062), .A2(n1216), .A3(n1235), .ZN(n1211) );
XNOR2_X1 U893 ( .A(n1210), .B(n1236), .ZN(G45) );
XNOR2_X1 U894 ( .A(G143), .B(KEYINPUT55), .ZN(n1236) );
AND4_X1 U895 ( .A1(n1237), .A2(n1216), .A3(n1238), .A4(n1239), .ZN(n1210) );
XOR2_X1 U896 ( .A(n1214), .B(n1240), .Z(G42) );
XNOR2_X1 U897 ( .A(KEYINPUT2), .B(n1131), .ZN(n1240) );
AND3_X1 U898 ( .A1(n1098), .A2(n1241), .A3(n1217), .ZN(n1214) );
INV_X1 U899 ( .A(n1242), .ZN(n1217) );
XNOR2_X1 U900 ( .A(G137), .B(n1243), .ZN(G39) );
NAND2_X1 U901 ( .A1(n1098), .A2(n1244), .ZN(n1243) );
XNOR2_X1 U902 ( .A(KEYINPUT37), .B(n1219), .ZN(n1244) );
NAND2_X1 U903 ( .A1(n1235), .A2(n1066), .ZN(n1219) );
XNOR2_X1 U904 ( .A(n1245), .B(n1209), .ZN(G36) );
AND3_X1 U905 ( .A1(n1098), .A2(n1063), .A3(n1237), .ZN(n1209) );
XNOR2_X1 U906 ( .A(n1246), .B(n1247), .ZN(G33) );
NOR2_X1 U907 ( .A1(KEYINPUT53), .A2(n1215), .ZN(n1247) );
NAND3_X1 U908 ( .A1(n1062), .A2(n1098), .A3(n1237), .ZN(n1215) );
AND3_X1 U909 ( .A1(n1241), .A2(n1248), .A3(n1100), .ZN(n1237) );
NOR2_X1 U910 ( .A1(n1249), .A2(n1084), .ZN(n1098) );
XOR2_X1 U911 ( .A(n1212), .B(n1250), .Z(G30) );
NOR2_X1 U912 ( .A1(KEYINPUT14), .A2(n1251), .ZN(n1250) );
AND3_X1 U913 ( .A1(n1063), .A2(n1216), .A3(n1235), .ZN(n1212) );
AND4_X1 U914 ( .A1(n1252), .A2(n1099), .A3(n1241), .A4(n1248), .ZN(n1235) );
XNOR2_X1 U915 ( .A(G101), .B(n1228), .ZN(G3) );
NAND3_X1 U916 ( .A1(n1067), .A2(n1253), .A3(n1100), .ZN(n1228) );
AND2_X1 U917 ( .A1(n1066), .A2(n1241), .ZN(n1067) );
XNOR2_X1 U918 ( .A(n1254), .B(n1255), .ZN(G27) );
NOR3_X1 U919 ( .A1(n1256), .A2(n1073), .A3(n1242), .ZN(n1255) );
NAND4_X1 U920 ( .A1(n1099), .A2(n1062), .A3(n1089), .A4(n1248), .ZN(n1242) );
NAND2_X1 U921 ( .A1(n1257), .A2(n1258), .ZN(n1248) );
OR4_X1 U922 ( .A1(n1259), .A2(n1116), .A3(n1260), .A4(G900), .ZN(n1258) );
XNOR2_X1 U923 ( .A(KEYINPUT46), .B(n1261), .ZN(n1257) );
XNOR2_X1 U924 ( .A(KEYINPUT8), .B(n1095), .ZN(n1256) );
INV_X1 U925 ( .A(n1216), .ZN(n1095) );
XNOR2_X1 U926 ( .A(G122), .B(n1230), .ZN(G24) );
NAND3_X1 U927 ( .A1(n1093), .A2(n1262), .A3(n1263), .ZN(n1230) );
NOR3_X1 U928 ( .A1(n1252), .A2(n1264), .A3(n1265), .ZN(n1263) );
NAND2_X1 U929 ( .A1(n1266), .A2(n1267), .ZN(G21) );
NAND2_X1 U930 ( .A1(G119), .A2(n1220), .ZN(n1267) );
XOR2_X1 U931 ( .A(n1268), .B(KEYINPUT50), .Z(n1266) );
OR2_X1 U932 ( .A1(n1220), .A2(G119), .ZN(n1268) );
NAND4_X1 U933 ( .A1(n1252), .A2(n1262), .A3(n1099), .A4(n1066), .ZN(n1220) );
XNOR2_X1 U934 ( .A(G116), .B(n1221), .ZN(G18) );
NAND3_X1 U935 ( .A1(n1100), .A2(n1063), .A3(n1262), .ZN(n1221) );
NOR2_X1 U936 ( .A1(n1239), .A2(n1265), .ZN(n1063) );
INV_X1 U937 ( .A(n1238), .ZN(n1265) );
XOR2_X1 U938 ( .A(G113), .B(n1226), .Z(G15) );
AND3_X1 U939 ( .A1(n1262), .A2(n1100), .A3(n1062), .ZN(n1226) );
NOR2_X1 U940 ( .A1(n1238), .A2(n1264), .ZN(n1062) );
INV_X1 U941 ( .A(n1239), .ZN(n1264) );
AND2_X1 U942 ( .A1(n1252), .A2(n1093), .ZN(n1100) );
XOR2_X1 U943 ( .A(n1099), .B(KEYINPUT12), .Z(n1093) );
INV_X1 U944 ( .A(n1089), .ZN(n1252) );
AND2_X1 U945 ( .A1(n1060), .A2(n1253), .ZN(n1262) );
INV_X1 U946 ( .A(n1073), .ZN(n1060) );
NAND2_X1 U947 ( .A1(n1064), .A2(n1269), .ZN(n1073) );
XNOR2_X1 U948 ( .A(n1270), .B(n1225), .ZN(G12) );
AND3_X1 U949 ( .A1(n1099), .A2(n1227), .A3(n1066), .ZN(n1225) );
NOR2_X1 U950 ( .A1(n1238), .A2(n1239), .ZN(n1066) );
XOR2_X1 U951 ( .A(G475), .B(n1271), .Z(n1239) );
NOR2_X1 U952 ( .A1(KEYINPUT48), .A2(n1080), .ZN(n1271) );
NAND2_X1 U953 ( .A1(n1160), .A2(n1259), .ZN(n1080) );
XNOR2_X1 U954 ( .A(n1272), .B(n1273), .ZN(n1160) );
XOR2_X1 U955 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U956 ( .A(n1276), .B(G113), .ZN(n1275) );
XNOR2_X1 U957 ( .A(KEYINPUT19), .B(n1246), .ZN(n1274) );
XOR2_X1 U958 ( .A(n1277), .B(n1278), .Z(n1272) );
XNOR2_X1 U959 ( .A(G104), .B(n1279), .ZN(n1278) );
NAND4_X1 U960 ( .A1(KEYINPUT21), .A2(G214), .A3(n1280), .A4(n1116), .ZN(n1279) );
XOR2_X1 U961 ( .A(n1281), .B(n1282), .Z(n1277) );
NOR3_X1 U962 ( .A1(n1127), .A2(n1283), .A3(n1284), .ZN(n1282) );
AND2_X1 U963 ( .A1(KEYINPUT62), .A2(n1128), .ZN(n1284) );
NOR2_X1 U964 ( .A1(KEYINPUT62), .A2(n1131), .ZN(n1283) );
NAND2_X1 U965 ( .A1(n1285), .A2(n1286), .ZN(n1238) );
NAND2_X1 U966 ( .A1(KEYINPUT29), .A2(n1287), .ZN(n1286) );
NAND2_X1 U967 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U968 ( .A1(n1079), .A2(n1078), .ZN(n1289) );
INV_X1 U969 ( .A(n1083), .ZN(n1288) );
NOR2_X1 U970 ( .A1(n1078), .A2(n1079), .ZN(n1083) );
INV_X1 U971 ( .A(G478), .ZN(n1078) );
NAND2_X1 U972 ( .A1(n1290), .A2(n1291), .ZN(n1285) );
INV_X1 U973 ( .A(KEYINPUT29), .ZN(n1291) );
XNOR2_X1 U974 ( .A(n1079), .B(G478), .ZN(n1290) );
NOR2_X1 U975 ( .A1(n1155), .A2(G902), .ZN(n1079) );
XNOR2_X1 U976 ( .A(n1292), .B(n1293), .ZN(n1155) );
XOR2_X1 U977 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U978 ( .A(n1296), .B(n1297), .Z(n1295) );
NAND2_X1 U979 ( .A1(KEYINPUT32), .A2(n1276), .ZN(n1297) );
NAND2_X1 U980 ( .A1(G217), .A2(n1298), .ZN(n1296) );
XOR2_X1 U981 ( .A(n1299), .B(n1300), .Z(n1292) );
XNOR2_X1 U982 ( .A(n1245), .B(G107), .ZN(n1300) );
NAND3_X1 U983 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1299) );
NAND2_X1 U984 ( .A1(KEYINPUT56), .A2(n1304), .ZN(n1303) );
NAND3_X1 U985 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1302) );
INV_X1 U986 ( .A(KEYINPUT56), .ZN(n1306) );
OR2_X1 U987 ( .A1(n1307), .A2(n1305), .ZN(n1301) );
NOR2_X1 U988 ( .A1(KEYINPUT26), .A2(n1304), .ZN(n1305) );
XNOR2_X1 U989 ( .A(n1251), .B(KEYINPUT47), .ZN(n1304) );
AND3_X1 U990 ( .A1(n1253), .A2(n1089), .A3(n1241), .ZN(n1227) );
NOR2_X1 U991 ( .A1(n1064), .A2(n1065), .ZN(n1241) );
INV_X1 U992 ( .A(n1269), .ZN(n1065) );
NAND2_X1 U993 ( .A1(G221), .A2(n1308), .ZN(n1269) );
XOR2_X1 U994 ( .A(KEYINPUT31), .B(n1309), .Z(n1308) );
NOR2_X1 U995 ( .A1(G902), .A2(n1310), .ZN(n1309) );
XOR2_X1 U996 ( .A(n1311), .B(G469), .Z(n1064) );
NAND3_X1 U997 ( .A1(n1312), .A2(n1313), .A3(n1259), .ZN(n1311) );
NAND2_X1 U998 ( .A1(KEYINPUT57), .A2(n1314), .ZN(n1313) );
XOR2_X1 U999 ( .A(n1194), .B(n1315), .Z(n1314) );
NAND3_X1 U1000 ( .A1(n1315), .A2(n1194), .A3(n1316), .ZN(n1312) );
INV_X1 U1001 ( .A(KEYINPUT57), .ZN(n1316) );
XOR2_X1 U1002 ( .A(n1317), .B(n1318), .Z(n1194) );
XNOR2_X1 U1003 ( .A(G101), .B(n1319), .ZN(n1318) );
NAND2_X1 U1004 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NAND2_X1 U1005 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NAND2_X1 U1006 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
NAND2_X1 U1007 ( .A1(G107), .A2(n1326), .ZN(n1325) );
INV_X1 U1008 ( .A(KEYINPUT39), .ZN(n1324) );
NAND2_X1 U1009 ( .A1(n1327), .A2(n1042), .ZN(n1320) );
INV_X1 U1010 ( .A(G107), .ZN(n1042) );
NAND2_X1 U1011 ( .A1(n1326), .A2(n1328), .ZN(n1327) );
OR2_X1 U1012 ( .A1(n1322), .A2(KEYINPUT39), .ZN(n1328) );
XOR2_X1 U1013 ( .A(G104), .B(KEYINPUT6), .Z(n1322) );
INV_X1 U1014 ( .A(KEYINPUT15), .ZN(n1326) );
XNOR2_X1 U1015 ( .A(n1181), .B(n1129), .ZN(n1317) );
XNOR2_X1 U1016 ( .A(n1329), .B(n1330), .ZN(n1129) );
XNOR2_X1 U1017 ( .A(KEYINPUT45), .B(n1251), .ZN(n1330) );
NAND2_X1 U1018 ( .A1(KEYINPUT17), .A2(n1281), .ZN(n1329) );
AND2_X1 U1019 ( .A1(n1331), .A2(n1332), .ZN(n1315) );
NAND2_X1 U1020 ( .A1(n1333), .A2(n1197), .ZN(n1332) );
XOR2_X1 U1021 ( .A(n1195), .B(KEYINPUT25), .Z(n1333) );
NAND2_X1 U1022 ( .A1(n1334), .A2(n1335), .ZN(n1331) );
XOR2_X1 U1023 ( .A(n1195), .B(KEYINPUT61), .Z(n1335) );
XNOR2_X1 U1024 ( .A(G110), .B(G140), .ZN(n1195) );
INV_X1 U1025 ( .A(n1197), .ZN(n1334) );
NAND2_X1 U1026 ( .A1(n1336), .A2(n1116), .ZN(n1197) );
XOR2_X1 U1027 ( .A(KEYINPUT23), .B(G227), .Z(n1336) );
XNOR2_X1 U1028 ( .A(n1070), .B(KEYINPUT20), .ZN(n1089) );
XOR2_X1 U1029 ( .A(n1337), .B(G472), .Z(n1070) );
NAND2_X1 U1030 ( .A1(n1338), .A2(n1259), .ZN(n1337) );
XNOR2_X1 U1031 ( .A(n1181), .B(n1339), .ZN(n1338) );
XOR2_X1 U1032 ( .A(n1183), .B(n1340), .Z(n1339) );
NOR2_X1 U1033 ( .A1(n1186), .A2(n1341), .ZN(n1340) );
XOR2_X1 U1034 ( .A(KEYINPUT51), .B(n1342), .Z(n1341) );
NOR2_X1 U1035 ( .A1(n1187), .A2(n1343), .ZN(n1342) );
XNOR2_X1 U1036 ( .A(G101), .B(KEYINPUT30), .ZN(n1343) );
INV_X1 U1037 ( .A(n1344), .ZN(n1187) );
NOR2_X1 U1038 ( .A1(n1344), .A2(n1345), .ZN(n1186) );
NAND3_X1 U1039 ( .A1(n1280), .A2(n1116), .A3(G210), .ZN(n1344) );
XOR2_X1 U1040 ( .A(n1346), .B(n1347), .Z(n1183) );
XOR2_X1 U1041 ( .A(n1348), .B(KEYINPUT42), .Z(n1346) );
XNOR2_X1 U1042 ( .A(n1349), .B(n1350), .ZN(n1181) );
NOR2_X1 U1043 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
NOR3_X1 U1044 ( .A1(KEYINPUT13), .A2(G137), .A3(n1245), .ZN(n1352) );
NOR2_X1 U1045 ( .A1(n1122), .A2(n1353), .ZN(n1351) );
INV_X1 U1046 ( .A(KEYINPUT13), .ZN(n1353) );
XNOR2_X1 U1047 ( .A(n1245), .B(G137), .ZN(n1122) );
INV_X1 U1048 ( .A(G134), .ZN(n1245) );
NAND2_X1 U1049 ( .A1(KEYINPUT34), .A2(n1246), .ZN(n1349) );
INV_X1 U1050 ( .A(G131), .ZN(n1246) );
AND2_X1 U1051 ( .A1(n1216), .A2(n1354), .ZN(n1253) );
NAND2_X1 U1052 ( .A1(n1355), .A2(n1261), .ZN(n1354) );
INV_X1 U1053 ( .A(n1085), .ZN(n1261) );
NOR3_X1 U1054 ( .A1(n1046), .A2(n1260), .A3(n1356), .ZN(n1085) );
INV_X1 U1055 ( .A(G952), .ZN(n1356) );
XOR2_X1 U1056 ( .A(G953), .B(KEYINPUT54), .Z(n1046) );
OR4_X1 U1057 ( .A1(n1259), .A2(n1116), .A3(n1260), .A4(G898), .ZN(n1355) );
NOR2_X1 U1058 ( .A1(n1280), .A2(n1310), .ZN(n1260) );
INV_X1 U1059 ( .A(G237), .ZN(n1280) );
INV_X1 U1060 ( .A(G953), .ZN(n1116) );
NOR2_X1 U1061 ( .A1(n1097), .A2(n1084), .ZN(n1216) );
AND2_X1 U1062 ( .A1(G214), .A2(n1357), .ZN(n1084) );
INV_X1 U1063 ( .A(n1249), .ZN(n1097) );
XNOR2_X1 U1064 ( .A(n1069), .B(KEYINPUT22), .ZN(n1249) );
XOR2_X1 U1065 ( .A(n1358), .B(n1203), .Z(n1069) );
AND2_X1 U1066 ( .A1(G210), .A2(n1357), .ZN(n1203) );
NAND2_X1 U1067 ( .A1(n1359), .A2(n1259), .ZN(n1357) );
XNOR2_X1 U1068 ( .A(G237), .B(KEYINPUT28), .ZN(n1359) );
NAND2_X1 U1069 ( .A1(n1360), .A2(n1259), .ZN(n1358) );
XNOR2_X1 U1070 ( .A(n1361), .B(n1202), .ZN(n1360) );
XOR2_X1 U1071 ( .A(n1362), .B(n1143), .Z(n1202) );
XNOR2_X1 U1072 ( .A(n1270), .B(n1276), .ZN(n1143) );
INV_X1 U1073 ( .A(G122), .ZN(n1276) );
XNOR2_X1 U1074 ( .A(n1144), .B(n1363), .ZN(n1362) );
NOR2_X1 U1075 ( .A1(G953), .A2(n1137), .ZN(n1363) );
INV_X1 U1076 ( .A(G224), .ZN(n1137) );
XOR2_X1 U1077 ( .A(n1347), .B(n1364), .Z(n1144) );
NOR2_X1 U1078 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
XOR2_X1 U1079 ( .A(n1367), .B(KEYINPUT38), .Z(n1366) );
NAND2_X1 U1080 ( .A1(n1368), .A2(n1345), .ZN(n1367) );
NOR2_X1 U1081 ( .A1(n1368), .A2(n1345), .ZN(n1365) );
INV_X1 U1082 ( .A(G101), .ZN(n1345) );
XNOR2_X1 U1083 ( .A(G104), .B(G107), .ZN(n1368) );
XNOR2_X1 U1084 ( .A(n1369), .B(n1370), .ZN(n1347) );
XOR2_X1 U1085 ( .A(KEYINPUT4), .B(G119), .Z(n1370) );
XNOR2_X1 U1086 ( .A(G113), .B(n1294), .ZN(n1369) );
XOR2_X1 U1087 ( .A(G116), .B(KEYINPUT10), .Z(n1294) );
NAND2_X1 U1088 ( .A1(KEYINPUT24), .A2(n1200), .ZN(n1361) );
XNOR2_X1 U1089 ( .A(n1348), .B(G125), .ZN(n1200) );
XNOR2_X1 U1090 ( .A(n1281), .B(n1251), .ZN(n1348) );
INV_X1 U1091 ( .A(G128), .ZN(n1251) );
XNOR2_X1 U1092 ( .A(G146), .B(n1307), .ZN(n1281) );
XOR2_X1 U1093 ( .A(G143), .B(KEYINPUT9), .Z(n1307) );
XNOR2_X1 U1094 ( .A(n1371), .B(n1081), .ZN(n1099) );
NAND2_X1 U1095 ( .A1(n1148), .A2(n1259), .ZN(n1081) );
XNOR2_X1 U1096 ( .A(n1372), .B(n1373), .ZN(n1148) );
XOR2_X1 U1097 ( .A(n1374), .B(n1375), .Z(n1373) );
XNOR2_X1 U1098 ( .A(n1376), .B(n1270), .ZN(n1375) );
NAND4_X1 U1099 ( .A1(n1377), .A2(n1378), .A3(n1379), .A4(n1380), .ZN(n1376) );
OR2_X1 U1100 ( .A1(n1131), .A2(KEYINPUT36), .ZN(n1380) );
NAND2_X1 U1101 ( .A1(KEYINPUT36), .A2(n1128), .ZN(n1379) );
NOR2_X1 U1102 ( .A1(G125), .A2(G140), .ZN(n1128) );
INV_X1 U1103 ( .A(n1127), .ZN(n1378) );
NOR2_X1 U1104 ( .A1(n1131), .A2(n1254), .ZN(n1127) );
INV_X1 U1105 ( .A(G125), .ZN(n1254) );
INV_X1 U1106 ( .A(G140), .ZN(n1131) );
XNOR2_X1 U1107 ( .A(KEYINPUT59), .B(KEYINPUT1), .ZN(n1377) );
NAND2_X1 U1108 ( .A1(G221), .A2(n1298), .ZN(n1374) );
NOR2_X1 U1109 ( .A1(n1310), .A2(G953), .ZN(n1298) );
INV_X1 U1110 ( .A(G234), .ZN(n1310) );
XOR2_X1 U1111 ( .A(n1381), .B(n1382), .Z(n1372) );
XNOR2_X1 U1112 ( .A(n1233), .B(G137), .ZN(n1382) );
INV_X1 U1113 ( .A(G146), .ZN(n1233) );
XNOR2_X1 U1114 ( .A(G119), .B(G128), .ZN(n1381) );
NAND2_X1 U1115 ( .A1(KEYINPUT49), .A2(n1151), .ZN(n1371) );
NAND2_X1 U1116 ( .A1(G217), .A2(n1383), .ZN(n1151) );
NAND2_X1 U1117 ( .A1(G234), .A2(n1259), .ZN(n1383) );
INV_X1 U1118 ( .A(G902), .ZN(n1259) );
INV_X1 U1119 ( .A(G110), .ZN(n1270) );
endmodule


