//Key = 1110011111010101010010110101010101001000001100000100110110100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278;

NAND2_X1 U707 ( .A1(n971), .A2(n972), .ZN(G9) );
NAND2_X1 U708 ( .A1(n973), .A2(n974), .ZN(n972) );
XOR2_X1 U709 ( .A(KEYINPUT5), .B(n975), .Z(n971) );
NOR2_X1 U710 ( .A1(n973), .A2(n974), .ZN(n975) );
NOR2_X1 U711 ( .A1(n976), .A2(n977), .ZN(G75) );
NOR3_X1 U712 ( .A1(n978), .A2(n979), .A3(n980), .ZN(n977) );
NOR2_X1 U713 ( .A1(n981), .A2(n982), .ZN(n979) );
NOR3_X1 U714 ( .A1(n983), .A2(n984), .A3(n985), .ZN(n981) );
NOR2_X1 U715 ( .A1(n986), .A2(n987), .ZN(n985) );
INV_X1 U716 ( .A(n988), .ZN(n987) );
NOR2_X1 U717 ( .A1(n989), .A2(n990), .ZN(n986) );
XNOR2_X1 U718 ( .A(n991), .B(KEYINPUT31), .ZN(n990) );
NOR3_X1 U719 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n984) );
NOR2_X1 U720 ( .A1(n995), .A2(n996), .ZN(n993) );
NOR2_X1 U721 ( .A1(n997), .A2(n998), .ZN(n996) );
NOR2_X1 U722 ( .A1(n999), .A2(n1000), .ZN(n997) );
NOR2_X1 U723 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NOR2_X1 U724 ( .A1(n1003), .A2(n1004), .ZN(n995) );
NOR2_X1 U725 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
NOR2_X1 U726 ( .A1(KEYINPUT26), .A2(n1007), .ZN(n1006) );
NOR2_X1 U727 ( .A1(n1008), .A2(n1009), .ZN(n1005) );
NOR2_X1 U728 ( .A1(n1010), .A2(n1011), .ZN(n983) );
INV_X1 U729 ( .A(KEYINPUT26), .ZN(n1011) );
NOR4_X1 U730 ( .A1(n1007), .A2(n1004), .A3(n994), .A4(n992), .ZN(n1010) );
NAND3_X1 U731 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n978) );
NAND2_X1 U732 ( .A1(n988), .A2(n1015), .ZN(n1014) );
NAND2_X1 U733 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND4_X1 U734 ( .A1(n1018), .A2(n1019), .A3(G214), .A4(n1020), .ZN(n1017) );
XNOR2_X1 U735 ( .A(n1021), .B(KEYINPUT7), .ZN(n1018) );
NAND2_X1 U736 ( .A1(n1021), .A2(n1022), .ZN(n1016) );
NOR3_X1 U737 ( .A1(n998), .A2(n1004), .A3(n992), .ZN(n988) );
NOR3_X1 U738 ( .A1(n1023), .A2(G953), .A3(G952), .ZN(n976) );
INV_X1 U739 ( .A(n1012), .ZN(n1023) );
NAND4_X1 U740 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1012) );
NOR3_X1 U741 ( .A1(n1028), .A2(n1029), .A3(n1004), .ZN(n1027) );
XOR2_X1 U742 ( .A(n1030), .B(n1031), .Z(n1026) );
NOR2_X1 U743 ( .A1(KEYINPUT30), .A2(n1032), .ZN(n1031) );
NAND2_X1 U744 ( .A1(n1033), .A2(n1034), .ZN(G72) );
NAND2_X1 U745 ( .A1(n1035), .A2(n1013), .ZN(n1034) );
XOR2_X1 U746 ( .A(n1036), .B(n1037), .Z(n1035) );
NAND2_X1 U747 ( .A1(KEYINPUT33), .A2(n1038), .ZN(n1037) );
NAND2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
INV_X1 U749 ( .A(n1041), .ZN(n1040) );
NAND2_X1 U750 ( .A1(n1042), .A2(G953), .ZN(n1033) );
XOR2_X1 U751 ( .A(n1036), .B(n1043), .Z(n1042) );
AND2_X1 U752 ( .A1(G227), .A2(G900), .ZN(n1043) );
NAND2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(n1036) );
NAND2_X1 U754 ( .A1(G953), .A2(n1046), .ZN(n1045) );
XOR2_X1 U755 ( .A(n1047), .B(n1048), .Z(n1044) );
XOR2_X1 U756 ( .A(n1049), .B(n1050), .Z(n1048) );
NAND2_X1 U757 ( .A1(KEYINPUT17), .A2(G125), .ZN(n1050) );
NAND2_X1 U758 ( .A1(KEYINPUT9), .A2(n1051), .ZN(n1049) );
XNOR2_X1 U759 ( .A(n1052), .B(G134), .ZN(n1051) );
XOR2_X1 U760 ( .A(n1053), .B(n1054), .Z(n1047) );
XOR2_X1 U761 ( .A(n1055), .B(n1056), .Z(G69) );
XOR2_X1 U762 ( .A(n1057), .B(n1058), .Z(n1056) );
NOR2_X1 U763 ( .A1(n1059), .A2(G953), .ZN(n1058) );
NOR2_X1 U764 ( .A1(n1060), .A2(n1061), .ZN(n1057) );
XOR2_X1 U765 ( .A(n1062), .B(n1063), .Z(n1061) );
NAND2_X1 U766 ( .A1(KEYINPUT11), .A2(n1064), .ZN(n1062) );
NOR2_X1 U767 ( .A1(G898), .A2(n1013), .ZN(n1060) );
NOR2_X1 U768 ( .A1(n1065), .A2(n1013), .ZN(n1055) );
NOR2_X1 U769 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U770 ( .A1(n1068), .A2(n1069), .ZN(G66) );
XNOR2_X1 U771 ( .A(n1070), .B(n1071), .ZN(n1069) );
NOR2_X1 U772 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U773 ( .A1(n1068), .A2(n1074), .ZN(G63) );
XOR2_X1 U774 ( .A(n1075), .B(n1076), .Z(n1074) );
AND2_X1 U775 ( .A1(G478), .A2(n1077), .ZN(n1075) );
NOR2_X1 U776 ( .A1(n1068), .A2(n1078), .ZN(G60) );
XNOR2_X1 U777 ( .A(n1079), .B(n1080), .ZN(n1078) );
NOR2_X1 U778 ( .A1(n1032), .A2(n1073), .ZN(n1080) );
XOR2_X1 U779 ( .A(n1081), .B(n1082), .Z(G6) );
XNOR2_X1 U780 ( .A(G104), .B(KEYINPUT51), .ZN(n1082) );
NAND3_X1 U781 ( .A1(n1083), .A2(n1084), .A3(n991), .ZN(n1081) );
XNOR2_X1 U782 ( .A(KEYINPUT50), .B(n1004), .ZN(n1084) );
NOR2_X1 U783 ( .A1(n1068), .A2(n1085), .ZN(G57) );
XOR2_X1 U784 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND2_X1 U785 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NAND2_X1 U786 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U787 ( .A(n1092), .B(KEYINPUT38), .Z(n1088) );
OR2_X1 U788 ( .A1(n1091), .A2(n1090), .ZN(n1092) );
XNOR2_X1 U789 ( .A(n1093), .B(n1094), .ZN(n1090) );
NOR2_X1 U790 ( .A1(KEYINPUT14), .A2(n1095), .ZN(n1094) );
XOR2_X1 U791 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U792 ( .A1(n1077), .A2(G472), .ZN(n1091) );
NOR2_X1 U793 ( .A1(n1068), .A2(n1098), .ZN(G54) );
XOR2_X1 U794 ( .A(n1099), .B(n1100), .Z(n1098) );
XOR2_X1 U795 ( .A(n1101), .B(n1102), .Z(n1100) );
NAND3_X1 U796 ( .A1(n1077), .A2(G469), .A3(KEYINPUT42), .ZN(n1101) );
XOR2_X1 U797 ( .A(n1103), .B(n1104), .Z(n1099) );
NOR2_X1 U798 ( .A1(KEYINPUT59), .A2(n1105), .ZN(n1104) );
XOR2_X1 U799 ( .A(n1106), .B(KEYINPUT55), .Z(n1103) );
NAND2_X1 U800 ( .A1(n1107), .A2(KEYINPUT1), .ZN(n1106) );
XOR2_X1 U801 ( .A(n1053), .B(n1108), .Z(n1107) );
XNOR2_X1 U802 ( .A(n1096), .B(n1109), .ZN(n1108) );
NOR2_X1 U803 ( .A1(n1068), .A2(n1110), .ZN(G51) );
XOR2_X1 U804 ( .A(n1111), .B(n1112), .Z(n1110) );
XNOR2_X1 U805 ( .A(n1113), .B(n1114), .ZN(n1112) );
XOR2_X1 U806 ( .A(n1115), .B(KEYINPUT19), .Z(n1111) );
NAND2_X1 U807 ( .A1(n1077), .A2(G210), .ZN(n1115) );
INV_X1 U808 ( .A(n1073), .ZN(n1077) );
NAND2_X1 U809 ( .A1(G902), .A2(n980), .ZN(n1073) );
NAND3_X1 U810 ( .A1(n1059), .A2(n1039), .A3(n1116), .ZN(n980) );
XNOR2_X1 U811 ( .A(n1041), .B(KEYINPUT41), .ZN(n1116) );
AND4_X1 U812 ( .A1(n1117), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1039) );
NOR3_X1 U813 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1120) );
NOR3_X1 U814 ( .A1(n1124), .A2(n982), .A3(n994), .ZN(n1123) );
NOR2_X1 U815 ( .A1(n1125), .A2(n1126), .ZN(n1121) );
NOR2_X1 U816 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
XOR2_X1 U817 ( .A(KEYINPUT3), .B(n1129), .Z(n1128) );
NOR2_X1 U818 ( .A1(n998), .A2(n1130), .ZN(n1127) );
AND4_X1 U819 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1059) );
AND4_X1 U820 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1134) );
OR3_X1 U821 ( .A1(n1139), .A2(n1004), .A3(n1140), .ZN(n1138) );
INV_X1 U822 ( .A(n1141), .ZN(n1135) );
NOR2_X1 U823 ( .A1(n973), .A2(n1142), .ZN(n1133) );
NOR3_X1 U824 ( .A1(n1143), .A2(n1004), .A3(n1140), .ZN(n973) );
NAND2_X1 U825 ( .A1(n1144), .A2(n1145), .ZN(n1131) );
INV_X1 U826 ( .A(n1146), .ZN(n1145) );
XNOR2_X1 U827 ( .A(n1147), .B(KEYINPUT20), .ZN(n1144) );
NOR2_X1 U828 ( .A1(n1013), .A2(G952), .ZN(n1068) );
XNOR2_X1 U829 ( .A(n1148), .B(n1041), .ZN(G48) );
NOR3_X1 U830 ( .A1(n1139), .A2(n1126), .A3(n1124), .ZN(n1041) );
INV_X1 U831 ( .A(n1022), .ZN(n1126) );
XOR2_X1 U832 ( .A(G143), .B(n1122), .Z(G45) );
AND4_X1 U833 ( .A1(n1149), .A2(n1022), .A3(n1028), .A4(n1150), .ZN(n1122) );
NAND2_X1 U834 ( .A1(n1151), .A2(n1152), .ZN(G42) );
NAND2_X1 U835 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U836 ( .A(n1118), .B(KEYINPUT27), .Z(n1153) );
NAND2_X1 U837 ( .A1(G140), .A2(n1155), .ZN(n1151) );
XOR2_X1 U838 ( .A(n1118), .B(KEYINPUT34), .Z(n1155) );
OR3_X1 U839 ( .A1(n982), .A2(n1007), .A3(n1130), .ZN(n1118) );
INV_X1 U840 ( .A(n1156), .ZN(n1007) );
XNOR2_X1 U841 ( .A(G137), .B(n1157), .ZN(G39) );
NAND3_X1 U842 ( .A1(n1025), .A2(n1158), .A3(KEYINPUT43), .ZN(n1157) );
XOR2_X1 U843 ( .A(KEYINPUT32), .B(n1159), .Z(n1158) );
NOR2_X1 U844 ( .A1(n994), .A2(n1124), .ZN(n1159) );
XNOR2_X1 U845 ( .A(G134), .B(n1119), .ZN(G36) );
NAND3_X1 U846 ( .A1(n1025), .A2(n989), .A3(n1149), .ZN(n1119) );
XNOR2_X1 U847 ( .A(G131), .B(n1117), .ZN(G33) );
NAND3_X1 U848 ( .A1(n991), .A2(n1025), .A3(n1149), .ZN(n1117) );
AND3_X1 U849 ( .A1(n1156), .A2(n1160), .A3(n1000), .ZN(n1149) );
INV_X1 U850 ( .A(n982), .ZN(n1025) );
NAND2_X1 U851 ( .A1(n1019), .A2(n1161), .ZN(n982) );
NAND2_X1 U852 ( .A1(G214), .A2(n1020), .ZN(n1161) );
XNOR2_X1 U853 ( .A(G128), .B(n1162), .ZN(G30) );
NAND3_X1 U854 ( .A1(n1129), .A2(n1022), .A3(KEYINPUT58), .ZN(n1162) );
NOR2_X1 U855 ( .A1(n1124), .A2(n1143), .ZN(n1129) );
INV_X1 U856 ( .A(n989), .ZN(n1143) );
NAND4_X1 U857 ( .A1(n1156), .A2(n1163), .A3(n1002), .A4(n1160), .ZN(n1124) );
XNOR2_X1 U858 ( .A(G101), .B(n1137), .ZN(G3) );
NAND3_X1 U859 ( .A1(n1021), .A2(n1083), .A3(n1000), .ZN(n1137) );
INV_X1 U860 ( .A(n1140), .ZN(n1083) );
XOR2_X1 U861 ( .A(G125), .B(n1164), .Z(G27) );
NOR3_X1 U862 ( .A1(n1130), .A2(n1165), .A3(n998), .ZN(n1164) );
XNOR2_X1 U863 ( .A(n1022), .B(KEYINPUT47), .ZN(n1165) );
NAND4_X1 U864 ( .A1(n1166), .A2(n991), .A3(n1163), .A4(n1160), .ZN(n1130) );
NAND2_X1 U865 ( .A1(n992), .A2(n1167), .ZN(n1160) );
NAND4_X1 U866 ( .A1(G953), .A2(G902), .A3(n1168), .A4(n1046), .ZN(n1167) );
INV_X1 U867 ( .A(G900), .ZN(n1046) );
XNOR2_X1 U868 ( .A(G122), .B(n1132), .ZN(G24) );
NAND4_X1 U869 ( .A1(n1028), .A2(n1150), .A3(n1169), .A4(n1170), .ZN(n1132) );
NOR2_X1 U870 ( .A1(n1004), .A2(n998), .ZN(n1170) );
NAND2_X1 U871 ( .A1(n1166), .A2(n1001), .ZN(n1004) );
XOR2_X1 U872 ( .A(G119), .B(n1142), .Z(G21) );
AND4_X1 U873 ( .A1(n1163), .A2(n1002), .A3(n1169), .A4(n1171), .ZN(n1142) );
NOR2_X1 U874 ( .A1(n994), .A2(n998), .ZN(n1171) );
XOR2_X1 U875 ( .A(G116), .B(n1172), .Z(G18) );
NOR2_X1 U876 ( .A1(n998), .A2(n1146), .ZN(n1172) );
NAND3_X1 U877 ( .A1(n989), .A2(n1169), .A3(n1000), .ZN(n1146) );
NOR2_X1 U878 ( .A1(n1150), .A2(n1173), .ZN(n989) );
INV_X1 U879 ( .A(n1028), .ZN(n1173) );
INV_X1 U880 ( .A(n1147), .ZN(n998) );
XNOR2_X1 U881 ( .A(G113), .B(n1136), .ZN(G15) );
NAND4_X1 U882 ( .A1(n1000), .A2(n991), .A3(n1147), .A4(n1169), .ZN(n1136) );
NOR2_X1 U883 ( .A1(n1008), .A2(n1029), .ZN(n1147) );
XOR2_X1 U884 ( .A(n1174), .B(KEYINPUT35), .Z(n1008) );
INV_X1 U885 ( .A(n1139), .ZN(n991) );
NAND2_X1 U886 ( .A1(n1175), .A2(n1150), .ZN(n1139) );
XOR2_X1 U887 ( .A(n1176), .B(KEYINPUT0), .Z(n1175) );
NOR2_X1 U888 ( .A1(n1163), .A2(n1166), .ZN(n1000) );
INV_X1 U889 ( .A(n1002), .ZN(n1166) );
NAND2_X1 U890 ( .A1(n1177), .A2(n1178), .ZN(G12) );
NAND2_X1 U891 ( .A1(n1141), .A2(n1179), .ZN(n1178) );
XOR2_X1 U892 ( .A(n1180), .B(KEYINPUT46), .Z(n1177) );
OR2_X1 U893 ( .A1(n1179), .A2(n1141), .ZN(n1180) );
NOR4_X1 U894 ( .A1(n994), .A2(n1140), .A3(n1002), .A4(n1001), .ZN(n1141) );
INV_X1 U895 ( .A(n1163), .ZN(n1001) );
XOR2_X1 U896 ( .A(n1181), .B(n1072), .Z(n1163) );
NAND2_X1 U897 ( .A1(G217), .A2(n1182), .ZN(n1072) );
NAND2_X1 U898 ( .A1(n1070), .A2(n1183), .ZN(n1181) );
XNOR2_X1 U899 ( .A(n1184), .B(n1185), .ZN(n1070) );
XOR2_X1 U900 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U901 ( .A(n1188), .B(n1189), .Z(n1187) );
NOR3_X1 U902 ( .A1(KEYINPUT39), .A2(n1190), .A3(n1191), .ZN(n1189) );
NOR2_X1 U903 ( .A1(n1148), .A2(n1192), .ZN(n1191) );
XOR2_X1 U904 ( .A(n1193), .B(KEYINPUT13), .Z(n1192) );
NOR2_X1 U905 ( .A1(G146), .A2(n1194), .ZN(n1190) );
XOR2_X1 U906 ( .A(n1193), .B(KEYINPUT63), .Z(n1194) );
XOR2_X1 U907 ( .A(n1195), .B(G125), .Z(n1193) );
NAND2_X1 U908 ( .A1(KEYINPUT49), .A2(n1154), .ZN(n1195) );
INV_X1 U909 ( .A(G140), .ZN(n1154) );
NOR2_X1 U910 ( .A1(n1196), .A2(n1197), .ZN(n1188) );
XOR2_X1 U911 ( .A(KEYINPUT16), .B(n1198), .Z(n1197) );
AND2_X1 U912 ( .A1(n1199), .A2(n1052), .ZN(n1198) );
NOR2_X1 U913 ( .A1(n1052), .A2(n1199), .ZN(n1196) );
NAND3_X1 U914 ( .A1(G234), .A2(n1013), .A3(G221), .ZN(n1199) );
INV_X1 U915 ( .A(G137), .ZN(n1052) );
XOR2_X1 U916 ( .A(G119), .B(G110), .Z(n1186) );
XOR2_X1 U917 ( .A(n1200), .B(n1201), .Z(n1184) );
XNOR2_X1 U918 ( .A(KEYINPUT56), .B(n1202), .ZN(n1201) );
XNOR2_X1 U919 ( .A(KEYINPUT8), .B(KEYINPUT61), .ZN(n1200) );
XNOR2_X1 U920 ( .A(n1203), .B(G472), .ZN(n1002) );
NAND2_X1 U921 ( .A1(n1204), .A2(n1183), .ZN(n1203) );
XOR2_X1 U922 ( .A(n1205), .B(n1206), .Z(n1204) );
XNOR2_X1 U923 ( .A(n1087), .B(n1093), .ZN(n1206) );
XOR2_X1 U924 ( .A(n1207), .B(n1208), .Z(n1093) );
INV_X1 U925 ( .A(n1209), .ZN(n1208) );
XNOR2_X1 U926 ( .A(G119), .B(G113), .ZN(n1207) );
XNOR2_X1 U927 ( .A(n1210), .B(G101), .ZN(n1087) );
NAND2_X1 U928 ( .A1(n1211), .A2(G210), .ZN(n1210) );
XNOR2_X1 U929 ( .A(n1212), .B(n1096), .ZN(n1205) );
NAND2_X1 U930 ( .A1(KEYINPUT53), .A2(n1097), .ZN(n1212) );
NAND2_X1 U931 ( .A1(n1156), .A2(n1169), .ZN(n1140) );
AND2_X1 U932 ( .A1(n1022), .A2(n1213), .ZN(n1169) );
NAND2_X1 U933 ( .A1(n1214), .A2(n992), .ZN(n1213) );
NAND3_X1 U934 ( .A1(n1168), .A2(n1013), .A3(G952), .ZN(n992) );
NAND4_X1 U935 ( .A1(G953), .A2(G902), .A3(n1168), .A4(n1067), .ZN(n1214) );
INV_X1 U936 ( .A(G898), .ZN(n1067) );
NAND2_X1 U937 ( .A1(G237), .A2(G234), .ZN(n1168) );
NOR2_X1 U938 ( .A1(n1019), .A2(n1215), .ZN(n1022) );
AND2_X1 U939 ( .A1(G214), .A2(n1020), .ZN(n1215) );
XOR2_X1 U940 ( .A(n1216), .B(n1217), .Z(n1019) );
NOR2_X1 U941 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XNOR2_X1 U942 ( .A(KEYINPUT44), .B(n1020), .ZN(n1219) );
NAND2_X1 U943 ( .A1(n1220), .A2(n1183), .ZN(n1020) );
XOR2_X1 U944 ( .A(KEYINPUT25), .B(G237), .Z(n1220) );
INV_X1 U945 ( .A(G210), .ZN(n1218) );
NAND4_X1 U946 ( .A1(n1221), .A2(n1183), .A3(n1222), .A4(n1223), .ZN(n1216) );
NAND3_X1 U947 ( .A1(KEYINPUT2), .A2(n1114), .A3(n1224), .ZN(n1223) );
INV_X1 U948 ( .A(n1225), .ZN(n1114) );
OR2_X1 U949 ( .A1(n1224), .A2(KEYINPUT2), .ZN(n1222) );
NAND2_X1 U950 ( .A1(n1225), .A2(n1226), .ZN(n1221) );
NAND2_X1 U951 ( .A1(KEYINPUT2), .A2(n1227), .ZN(n1226) );
XOR2_X1 U952 ( .A(KEYINPUT10), .B(n1224), .Z(n1227) );
XOR2_X1 U953 ( .A(n1113), .B(KEYINPUT22), .Z(n1224) );
XNOR2_X1 U954 ( .A(n1097), .B(n1228), .ZN(n1113) );
XOR2_X1 U955 ( .A(G125), .B(n1229), .Z(n1228) );
NOR2_X1 U956 ( .A1(G953), .A2(n1066), .ZN(n1229) );
INV_X1 U957 ( .A(G224), .ZN(n1066) );
XOR2_X1 U958 ( .A(n1230), .B(KEYINPUT62), .Z(n1097) );
XNOR2_X1 U959 ( .A(n1063), .B(n1064), .ZN(n1225) );
XNOR2_X1 U960 ( .A(G110), .B(G122), .ZN(n1064) );
XOR2_X1 U961 ( .A(n1109), .B(n1231), .Z(n1063) );
NOR2_X1 U962 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
XOR2_X1 U963 ( .A(KEYINPUT40), .B(n1234), .Z(n1233) );
NOR2_X1 U964 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
AND2_X1 U965 ( .A1(n1236), .A2(n1235), .ZN(n1232) );
XOR2_X1 U966 ( .A(n1209), .B(n1237), .Z(n1235) );
NOR2_X1 U967 ( .A1(G119), .A2(KEYINPUT12), .ZN(n1237) );
NOR2_X1 U968 ( .A1(n1024), .A2(n1029), .ZN(n1156) );
INV_X1 U969 ( .A(n1009), .ZN(n1029) );
NAND2_X1 U970 ( .A1(G221), .A2(n1182), .ZN(n1009) );
NAND2_X1 U971 ( .A1(G234), .A2(n1183), .ZN(n1182) );
INV_X1 U972 ( .A(n1174), .ZN(n1024) );
XNOR2_X1 U973 ( .A(n1238), .B(G469), .ZN(n1174) );
NAND2_X1 U974 ( .A1(n1239), .A2(n1183), .ZN(n1238) );
XOR2_X1 U975 ( .A(n1102), .B(n1240), .Z(n1239) );
XOR2_X1 U976 ( .A(n1105), .B(n1241), .Z(n1240) );
NOR3_X1 U977 ( .A1(n1242), .A2(KEYINPUT48), .A3(n1243), .ZN(n1241) );
AND2_X1 U978 ( .A1(n1244), .A2(n1096), .ZN(n1243) );
XOR2_X1 U979 ( .A(KEYINPUT21), .B(n1245), .Z(n1242) );
NOR2_X1 U980 ( .A1(n1096), .A2(n1244), .ZN(n1245) );
XOR2_X1 U981 ( .A(n1246), .B(n1247), .Z(n1244) );
INV_X1 U982 ( .A(n1109), .ZN(n1247) );
XOR2_X1 U983 ( .A(G101), .B(n1248), .Z(n1109) );
XNOR2_X1 U984 ( .A(n974), .B(G104), .ZN(n1248) );
NAND2_X1 U985 ( .A1(KEYINPUT52), .A2(n1053), .ZN(n1246) );
XOR2_X1 U986 ( .A(n1230), .B(KEYINPUT36), .Z(n1053) );
XNOR2_X1 U987 ( .A(G128), .B(n1249), .ZN(n1230) );
XOR2_X1 U988 ( .A(n1250), .B(n1251), .Z(n1096) );
NOR2_X1 U989 ( .A1(G134), .A2(KEYINPUT28), .ZN(n1251) );
XNOR2_X1 U990 ( .A(G137), .B(n1252), .ZN(n1250) );
NOR2_X1 U991 ( .A1(KEYINPUT60), .A2(n1253), .ZN(n1252) );
NAND2_X1 U992 ( .A1(G227), .A2(n1013), .ZN(n1105) );
XNOR2_X1 U993 ( .A(G110), .B(G140), .ZN(n1102) );
INV_X1 U994 ( .A(n1021), .ZN(n994) );
NOR2_X1 U995 ( .A1(n1150), .A2(n1176), .ZN(n1021) );
XNOR2_X1 U996 ( .A(n1028), .B(KEYINPUT6), .ZN(n1176) );
XOR2_X1 U997 ( .A(G478), .B(n1254), .Z(n1028) );
NOR2_X1 U998 ( .A1(G902), .A2(n1076), .ZN(n1254) );
XNOR2_X1 U999 ( .A(n1255), .B(n1256), .ZN(n1076) );
XOR2_X1 U1000 ( .A(n1257), .B(n1258), .Z(n1256) );
XNOR2_X1 U1001 ( .A(n1259), .B(n974), .ZN(n1258) );
INV_X1 U1002 ( .A(G107), .ZN(n974) );
NAND3_X1 U1003 ( .A1(G234), .A2(n1013), .A3(G217), .ZN(n1259) );
INV_X1 U1004 ( .A(G953), .ZN(n1013) );
NAND3_X1 U1005 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1257) );
NAND2_X1 U1006 ( .A1(n1209), .A2(n1263), .ZN(n1262) );
OR3_X1 U1007 ( .A1(n1263), .A2(n1209), .A3(KEYINPUT54), .ZN(n1261) );
XOR2_X1 U1008 ( .A(G116), .B(KEYINPUT45), .Z(n1209) );
NAND2_X1 U1009 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
XNOR2_X1 U1010 ( .A(KEYINPUT4), .B(KEYINPUT37), .ZN(n1264) );
NAND2_X1 U1011 ( .A1(KEYINPUT54), .A2(G122), .ZN(n1260) );
XOR2_X1 U1012 ( .A(n1266), .B(n1267), .Z(n1255) );
XNOR2_X1 U1013 ( .A(G134), .B(n1202), .ZN(n1267) );
INV_X1 U1014 ( .A(G128), .ZN(n1202) );
XNOR2_X1 U1015 ( .A(G143), .B(KEYINPUT15), .ZN(n1266) );
XOR2_X1 U1016 ( .A(n1030), .B(n1032), .Z(n1150) );
INV_X1 U1017 ( .A(G475), .ZN(n1032) );
NAND2_X1 U1018 ( .A1(n1079), .A2(n1183), .ZN(n1030) );
INV_X1 U1019 ( .A(G902), .ZN(n1183) );
XNOR2_X1 U1020 ( .A(n1268), .B(n1269), .ZN(n1079) );
XNOR2_X1 U1021 ( .A(n1054), .B(n1270), .ZN(n1269) );
XOR2_X1 U1022 ( .A(n1271), .B(n1249), .Z(n1270) );
XNOR2_X1 U1023 ( .A(G143), .B(n1148), .ZN(n1249) );
INV_X1 U1024 ( .A(G146), .ZN(n1148) );
NAND2_X1 U1025 ( .A1(n1211), .A2(G214), .ZN(n1271) );
NOR2_X1 U1026 ( .A1(G953), .A2(G237), .ZN(n1211) );
XOR2_X1 U1027 ( .A(G140), .B(n1253), .Z(n1054) );
XOR2_X1 U1028 ( .A(G131), .B(KEYINPUT29), .Z(n1253) );
XOR2_X1 U1029 ( .A(n1272), .B(n1273), .Z(n1268) );
NOR2_X1 U1030 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XOR2_X1 U1031 ( .A(KEYINPUT24), .B(n1276), .Z(n1275) );
NOR2_X1 U1032 ( .A1(G122), .A2(n1236), .ZN(n1276) );
INV_X1 U1033 ( .A(G113), .ZN(n1236) );
NOR2_X1 U1034 ( .A1(G113), .A2(n1265), .ZN(n1274) );
INV_X1 U1035 ( .A(G122), .ZN(n1265) );
XNOR2_X1 U1036 ( .A(G104), .B(n1277), .ZN(n1272) );
NOR2_X1 U1037 ( .A1(KEYINPUT18), .A2(n1278), .ZN(n1277) );
XNOR2_X1 U1038 ( .A(G125), .B(KEYINPUT57), .ZN(n1278) );
XOR2_X1 U1039 ( .A(G110), .B(KEYINPUT23), .Z(n1179) );
endmodule


