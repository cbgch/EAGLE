//Key = 1001000001001010111011001001101110011101100101110000001010110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
n1456;

XOR2_X1 U797 ( .A(n1106), .B(n1107), .Z(G9) );
NAND3_X1 U798 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(G75) );
NAND2_X1 U799 ( .A1(G952), .A2(n1111), .ZN(n1110) );
NAND3_X1 U800 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
NAND2_X1 U801 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NAND2_X1 U802 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND4_X1 U803 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1118) );
NAND2_X1 U804 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND3_X1 U805 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1117) );
NAND2_X1 U806 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NAND2_X1 U807 ( .A1(n1120), .A2(n1130), .ZN(n1129) );
NAND2_X1 U808 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND3_X1 U809 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
INV_X1 U810 ( .A(KEYINPUT63), .ZN(n1134) );
NAND2_X1 U811 ( .A1(n1121), .A2(n1136), .ZN(n1131) );
NAND2_X1 U812 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U813 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NAND2_X1 U814 ( .A1(n1119), .A2(n1133), .ZN(n1128) );
NAND3_X1 U815 ( .A1(n1141), .A2(n1142), .A3(n1119), .ZN(n1133) );
NAND2_X1 U816 ( .A1(n1121), .A2(n1143), .ZN(n1142) );
OR2_X1 U817 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND2_X1 U818 ( .A1(n1120), .A2(n1146), .ZN(n1141) );
NAND2_X1 U819 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND3_X1 U820 ( .A1(G221), .A2(n1149), .A3(n1150), .ZN(n1148) );
NAND2_X1 U821 ( .A1(KEYINPUT63), .A2(n1135), .ZN(n1147) );
XNOR2_X1 U822 ( .A(KEYINPUT45), .B(n1151), .ZN(n1115) );
NAND4_X1 U823 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1108) );
NOR4_X1 U824 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
NOR3_X1 U825 ( .A1(KEYINPUT61), .A2(n1160), .A3(n1161), .ZN(n1158) );
NOR2_X1 U826 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
INV_X1 U827 ( .A(KEYINPUT14), .ZN(n1163) );
NOR2_X1 U828 ( .A1(G472), .A2(n1164), .ZN(n1162) );
NOR2_X1 U829 ( .A1(KEYINPUT14), .A2(G472), .ZN(n1160) );
NAND3_X1 U830 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1156) );
XOR2_X1 U831 ( .A(n1168), .B(KEYINPUT8), .Z(n1167) );
OR2_X1 U832 ( .A1(n1169), .A2(KEYINPUT40), .ZN(n1166) );
NAND2_X1 U833 ( .A1(n1170), .A2(KEYINPUT40), .ZN(n1165) );
NOR3_X1 U834 ( .A1(n1139), .A2(n1171), .A3(n1172), .ZN(n1154) );
NAND2_X1 U835 ( .A1(n1173), .A2(n1174), .ZN(n1153) );
NAND2_X1 U836 ( .A1(n1175), .A2(n1164), .ZN(n1152) );
NAND2_X1 U837 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NAND2_X1 U838 ( .A1(KEYINPUT61), .A2(KEYINPUT14), .ZN(n1177) );
INV_X1 U839 ( .A(G472), .ZN(n1176) );
NAND3_X1 U840 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(G72) );
XOR2_X1 U841 ( .A(n1181), .B(KEYINPUT1), .Z(n1180) );
NAND3_X1 U842 ( .A1(n1182), .A2(n1183), .A3(G953), .ZN(n1181) );
NAND2_X1 U843 ( .A1(G900), .A2(G227), .ZN(n1182) );
NAND2_X1 U844 ( .A1(n1184), .A2(n1109), .ZN(n1179) );
XOR2_X1 U845 ( .A(n1112), .B(n1183), .Z(n1184) );
NAND3_X1 U846 ( .A1(n1185), .A2(G227), .A3(G953), .ZN(n1178) );
INV_X1 U847 ( .A(n1183), .ZN(n1185) );
NAND3_X1 U848 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1183) );
XOR2_X1 U849 ( .A(KEYINPUT32), .B(n1189), .Z(n1188) );
NOR2_X1 U850 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND2_X1 U851 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
NAND2_X1 U852 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
OR2_X1 U853 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
XOR2_X1 U854 ( .A(n1196), .B(KEYINPUT23), .Z(n1192) );
NAND2_X1 U855 ( .A1(n1194), .A2(n1195), .ZN(n1196) );
XNOR2_X1 U856 ( .A(n1197), .B(n1198), .ZN(n1194) );
NAND2_X1 U857 ( .A1(G953), .A2(n1199), .ZN(n1186) );
XOR2_X1 U858 ( .A(n1200), .B(n1201), .Z(G69) );
NOR2_X1 U859 ( .A1(n1202), .A2(n1109), .ZN(n1201) );
AND2_X1 U860 ( .A1(G224), .A2(G898), .ZN(n1202) );
NAND2_X1 U861 ( .A1(n1203), .A2(n1204), .ZN(n1200) );
NAND2_X1 U862 ( .A1(n1205), .A2(n1109), .ZN(n1204) );
XOR2_X1 U863 ( .A(n1114), .B(n1206), .Z(n1205) );
OR3_X1 U864 ( .A1(n1207), .A2(n1206), .A3(n1109), .ZN(n1203) );
XNOR2_X1 U865 ( .A(n1208), .B(n1209), .ZN(n1206) );
NOR2_X1 U866 ( .A1(n1210), .A2(n1211), .ZN(G66) );
XOR2_X1 U867 ( .A(n1212), .B(n1213), .Z(n1211) );
NOR2_X1 U868 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NOR2_X1 U869 ( .A1(n1210), .A2(n1216), .ZN(G63) );
XOR2_X1 U870 ( .A(n1217), .B(n1218), .Z(n1216) );
XNOR2_X1 U871 ( .A(n1219), .B(KEYINPUT59), .ZN(n1218) );
NAND2_X1 U872 ( .A1(KEYINPUT54), .A2(n1220), .ZN(n1219) );
NAND2_X1 U873 ( .A1(n1221), .A2(G478), .ZN(n1220) );
NOR2_X1 U874 ( .A1(n1222), .A2(n1223), .ZN(G60) );
XOR2_X1 U875 ( .A(n1224), .B(n1225), .Z(n1223) );
NAND3_X1 U876 ( .A1(n1221), .A2(G475), .A3(KEYINPUT43), .ZN(n1224) );
NOR2_X1 U877 ( .A1(n1226), .A2(n1227), .ZN(n1222) );
XOR2_X1 U878 ( .A(KEYINPUT39), .B(G953), .Z(n1227) );
XOR2_X1 U879 ( .A(KEYINPUT49), .B(G952), .Z(n1226) );
NAND2_X1 U880 ( .A1(n1228), .A2(n1229), .ZN(G6) );
NAND2_X1 U881 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U882 ( .A(KEYINPUT0), .B(n1232), .Z(n1228) );
NOR2_X1 U883 ( .A1(n1230), .A2(n1231), .ZN(n1232) );
NOR2_X1 U884 ( .A1(n1210), .A2(n1233), .ZN(G57) );
XOR2_X1 U885 ( .A(n1234), .B(n1235), .Z(n1233) );
NAND2_X1 U886 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U887 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND3_X1 U888 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1239) );
NAND2_X1 U889 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
INV_X1 U890 ( .A(n1245), .ZN(n1238) );
NAND3_X1 U891 ( .A1(n1246), .A2(n1241), .A3(n1245), .ZN(n1236) );
NAND2_X1 U892 ( .A1(n1221), .A2(G472), .ZN(n1245) );
NAND2_X1 U893 ( .A1(KEYINPUT29), .A2(n1247), .ZN(n1241) );
XOR2_X1 U894 ( .A(n1248), .B(n1249), .Z(n1247) );
NAND2_X1 U895 ( .A1(n1250), .A2(n1244), .ZN(n1246) );
INV_X1 U896 ( .A(KEYINPUT29), .ZN(n1244) );
NAND2_X1 U897 ( .A1(n1251), .A2(n1252), .ZN(n1234) );
NOR2_X1 U898 ( .A1(n1210), .A2(n1253), .ZN(G54) );
XOR2_X1 U899 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U900 ( .A(n1256), .B(n1257), .Z(n1255) );
NAND2_X1 U901 ( .A1(KEYINPUT36), .A2(n1258), .ZN(n1256) );
XOR2_X1 U902 ( .A(n1259), .B(n1260), .Z(n1254) );
XOR2_X1 U903 ( .A(KEYINPUT7), .B(n1261), .Z(n1260) );
AND2_X1 U904 ( .A1(G469), .A2(n1221), .ZN(n1261) );
INV_X1 U905 ( .A(n1215), .ZN(n1221) );
NAND3_X1 U906 ( .A1(n1262), .A2(n1263), .A3(KEYINPUT30), .ZN(n1259) );
OR3_X1 U907 ( .A1(n1209), .A2(n1195), .A3(KEYINPUT27), .ZN(n1263) );
NAND2_X1 U908 ( .A1(n1264), .A2(KEYINPUT27), .ZN(n1262) );
NOR2_X1 U909 ( .A1(n1210), .A2(n1265), .ZN(G51) );
XOR2_X1 U910 ( .A(n1266), .B(n1267), .Z(n1265) );
NOR2_X1 U911 ( .A1(n1268), .A2(KEYINPUT60), .ZN(n1267) );
NOR2_X1 U912 ( .A1(n1269), .A2(n1215), .ZN(n1268) );
NAND2_X1 U913 ( .A1(G902), .A2(n1270), .ZN(n1215) );
NAND2_X1 U914 ( .A1(n1114), .A2(n1112), .ZN(n1270) );
AND4_X1 U915 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1112) );
NOR2_X1 U916 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NOR2_X1 U917 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NOR2_X1 U918 ( .A1(n1279), .A2(n1280), .ZN(n1277) );
XNOR2_X1 U919 ( .A(KEYINPUT10), .B(n1281), .ZN(n1280) );
NOR3_X1 U920 ( .A1(n1137), .A2(n1282), .A3(n1283), .ZN(n1275) );
NOR2_X1 U921 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NOR2_X1 U922 ( .A1(n1286), .A2(n1287), .ZN(n1284) );
NOR2_X1 U923 ( .A1(n1288), .A2(n1289), .ZN(n1286) );
NOR3_X1 U924 ( .A1(n1290), .A2(n1127), .A3(n1125), .ZN(n1289) );
AND2_X1 U925 ( .A1(n1291), .A2(n1292), .ZN(n1114) );
AND4_X1 U926 ( .A1(n1293), .A2(n1294), .A3(n1295), .A4(n1107), .ZN(n1292) );
NAND3_X1 U927 ( .A1(n1145), .A2(n1296), .A3(n1135), .ZN(n1107) );
NOR4_X1 U928 ( .A1(n1297), .A2(n1230), .A3(n1298), .A4(n1299), .ZN(n1291) );
NOR2_X1 U929 ( .A1(n1137), .A2(n1300), .ZN(n1299) );
AND3_X1 U930 ( .A1(n1135), .A2(n1296), .A3(n1144), .ZN(n1230) );
INV_X1 U931 ( .A(n1301), .ZN(n1297) );
NAND3_X1 U932 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1266) );
NAND2_X1 U933 ( .A1(KEYINPUT38), .A2(n1305), .ZN(n1304) );
OR3_X1 U934 ( .A1(n1305), .A2(KEYINPUT38), .A3(n1306), .ZN(n1303) );
NAND2_X1 U935 ( .A1(n1306), .A2(n1307), .ZN(n1302) );
NAND2_X1 U936 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
INV_X1 U937 ( .A(KEYINPUT38), .ZN(n1309) );
XNOR2_X1 U938 ( .A(KEYINPUT19), .B(n1305), .ZN(n1308) );
XNOR2_X1 U939 ( .A(G125), .B(n1310), .ZN(n1305) );
AND2_X1 U940 ( .A1(n1311), .A2(G953), .ZN(n1210) );
XNOR2_X1 U941 ( .A(KEYINPUT49), .B(G952), .ZN(n1311) );
XNOR2_X1 U942 ( .A(G146), .B(n1312), .ZN(G48) );
NAND3_X1 U943 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1312) );
NOR3_X1 U944 ( .A1(n1290), .A2(KEYINPUT5), .A3(n1287), .ZN(n1315) );
XOR2_X1 U945 ( .A(n1316), .B(KEYINPUT33), .Z(n1313) );
XOR2_X1 U946 ( .A(n1317), .B(n1318), .Z(G45) );
NAND3_X1 U947 ( .A1(n1319), .A2(n1320), .A3(n1288), .ZN(n1318) );
NOR3_X1 U948 ( .A1(n1124), .A2(n1168), .A3(n1321), .ZN(n1288) );
XOR2_X1 U949 ( .A(n1137), .B(KEYINPUT47), .Z(n1319) );
XOR2_X1 U950 ( .A(G140), .B(n1322), .Z(G42) );
NOR2_X1 U951 ( .A1(n1278), .A2(n1281), .ZN(n1322) );
NAND3_X1 U952 ( .A1(n1323), .A2(n1144), .A3(n1320), .ZN(n1281) );
XOR2_X1 U953 ( .A(n1197), .B(n1273), .Z(G39) );
NAND3_X1 U954 ( .A1(n1119), .A2(n1320), .A3(n1324), .ZN(n1273) );
AND3_X1 U955 ( .A1(n1120), .A2(n1325), .A3(n1326), .ZN(n1324) );
XNOR2_X1 U956 ( .A(G134), .B(n1271), .ZN(G36) );
NAND4_X1 U957 ( .A1(n1119), .A2(n1320), .A3(n1327), .A4(n1145), .ZN(n1271) );
XNOR2_X1 U958 ( .A(G131), .B(n1328), .ZN(G33) );
NAND2_X1 U959 ( .A1(n1329), .A2(n1119), .ZN(n1328) );
INV_X1 U960 ( .A(n1278), .ZN(n1119) );
NAND2_X1 U961 ( .A1(n1140), .A2(n1330), .ZN(n1278) );
XNOR2_X1 U962 ( .A(n1279), .B(KEYINPUT46), .ZN(n1329) );
AND3_X1 U963 ( .A1(n1144), .A2(n1327), .A3(n1320), .ZN(n1279) );
XNOR2_X1 U964 ( .A(G128), .B(n1272), .ZN(G30) );
NAND3_X1 U965 ( .A1(n1314), .A2(n1145), .A3(n1320), .ZN(n1272) );
NOR2_X1 U966 ( .A1(n1287), .A2(n1282), .ZN(n1320) );
INV_X1 U967 ( .A(n1316), .ZN(n1282) );
INV_X1 U968 ( .A(n1135), .ZN(n1287) );
XOR2_X1 U969 ( .A(G101), .B(n1298), .Z(G3) );
AND2_X1 U970 ( .A1(n1331), .A2(n1327), .ZN(n1298) );
XNOR2_X1 U971 ( .A(G125), .B(n1332), .ZN(G27) );
NAND4_X1 U972 ( .A1(KEYINPUT20), .A2(n1285), .A3(n1333), .A4(n1316), .ZN(n1332) );
NAND2_X1 U973 ( .A1(n1334), .A2(n1335), .ZN(n1316) );
XOR2_X1 U974 ( .A(n1336), .B(KEYINPUT15), .Z(n1334) );
NAND4_X1 U975 ( .A1(G953), .A2(G902), .A3(n1151), .A4(n1199), .ZN(n1336) );
INV_X1 U976 ( .A(G900), .ZN(n1199) );
NOR3_X1 U977 ( .A1(n1290), .A2(n1157), .A3(n1123), .ZN(n1285) );
XOR2_X1 U978 ( .A(n1337), .B(n1301), .Z(G24) );
NAND4_X1 U979 ( .A1(n1121), .A2(n1296), .A3(n1159), .A4(n1338), .ZN(n1301) );
NOR4_X1 U980 ( .A1(n1137), .A2(n1325), .A3(n1326), .A4(n1339), .ZN(n1296) );
XOR2_X1 U981 ( .A(n1294), .B(n1340), .Z(G21) );
NAND2_X1 U982 ( .A1(n1341), .A2(G119), .ZN(n1340) );
XNOR2_X1 U983 ( .A(KEYINPUT17), .B(KEYINPUT12), .ZN(n1341) );
NAND4_X1 U984 ( .A1(n1120), .A2(n1314), .A3(n1121), .A4(n1342), .ZN(n1294) );
NOR3_X1 U985 ( .A1(n1125), .A2(n1127), .A3(n1137), .ZN(n1314) );
XNOR2_X1 U986 ( .A(G116), .B(n1343), .ZN(G18) );
NAND2_X1 U987 ( .A1(n1344), .A2(n1333), .ZN(n1343) );
XOR2_X1 U988 ( .A(n1300), .B(KEYINPUT31), .Z(n1344) );
NAND4_X1 U989 ( .A1(n1327), .A2(n1121), .A3(n1145), .A4(n1342), .ZN(n1300) );
NOR2_X1 U990 ( .A1(n1338), .A2(n1321), .ZN(n1145) );
XOR2_X1 U991 ( .A(n1345), .B(n1293), .Z(G15) );
NAND4_X1 U992 ( .A1(n1144), .A2(n1327), .A3(n1346), .A4(n1121), .ZN(n1293) );
INV_X1 U993 ( .A(n1157), .ZN(n1121) );
NAND2_X1 U994 ( .A1(n1150), .A2(n1347), .ZN(n1157) );
NAND2_X1 U995 ( .A1(G221), .A2(n1149), .ZN(n1347) );
NOR2_X1 U996 ( .A1(n1339), .A2(n1137), .ZN(n1346) );
INV_X1 U997 ( .A(n1333), .ZN(n1137) );
INV_X1 U998 ( .A(n1342), .ZN(n1339) );
INV_X1 U999 ( .A(n1124), .ZN(n1327) );
NAND2_X1 U1000 ( .A1(n1127), .A2(n1326), .ZN(n1124) );
INV_X1 U1001 ( .A(n1125), .ZN(n1326) );
INV_X1 U1002 ( .A(n1290), .ZN(n1144) );
NAND2_X1 U1003 ( .A1(n1321), .A2(n1338), .ZN(n1290) );
XOR2_X1 U1004 ( .A(n1348), .B(G110), .Z(G12) );
NAND2_X1 U1005 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND3_X1 U1006 ( .A1(n1331), .A2(n1123), .A3(n1351), .ZN(n1350) );
OR2_X1 U1007 ( .A1(n1295), .A2(n1351), .ZN(n1349) );
INV_X1 U1008 ( .A(KEYINPUT37), .ZN(n1351) );
NAND2_X1 U1009 ( .A1(n1323), .A2(n1331), .ZN(n1295) );
AND4_X1 U1010 ( .A1(n1120), .A2(n1135), .A3(n1333), .A4(n1342), .ZN(n1331) );
NAND2_X1 U1011 ( .A1(n1335), .A2(n1352), .ZN(n1342) );
NAND4_X1 U1012 ( .A1(G953), .A2(G902), .A3(n1151), .A4(n1207), .ZN(n1352) );
INV_X1 U1013 ( .A(G898), .ZN(n1207) );
NAND3_X1 U1014 ( .A1(n1151), .A2(n1109), .A3(G952), .ZN(n1335) );
NAND2_X1 U1015 ( .A1(G237), .A2(G234), .ZN(n1151) );
NOR2_X1 U1016 ( .A1(n1140), .A2(n1139), .ZN(n1333) );
INV_X1 U1017 ( .A(n1330), .ZN(n1139) );
NAND2_X1 U1018 ( .A1(G214), .A2(n1353), .ZN(n1330) );
NOR2_X1 U1019 ( .A1(n1171), .A2(n1170), .ZN(n1140) );
AND2_X1 U1020 ( .A1(n1169), .A2(n1354), .ZN(n1170) );
NOR2_X1 U1021 ( .A1(n1354), .A2(n1169), .ZN(n1171) );
INV_X1 U1022 ( .A(n1269), .ZN(n1169) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1353), .ZN(n1269) );
NAND2_X1 U1024 ( .A1(n1355), .A2(n1356), .ZN(n1353) );
NAND2_X1 U1025 ( .A1(n1357), .A2(n1358), .ZN(n1354) );
XOR2_X1 U1026 ( .A(n1310), .B(n1359), .Z(n1357) );
XNOR2_X1 U1027 ( .A(n1360), .B(n1361), .ZN(n1359) );
NOR2_X1 U1028 ( .A1(KEYINPUT55), .A2(n1306), .ZN(n1361) );
XOR2_X1 U1029 ( .A(n1208), .B(n1362), .Z(n1306) );
NOR2_X1 U1030 ( .A1(KEYINPUT4), .A2(n1209), .ZN(n1362) );
XOR2_X1 U1031 ( .A(n1363), .B(n1364), .Z(n1208) );
NOR2_X1 U1032 ( .A1(KEYINPUT57), .A2(n1337), .ZN(n1364) );
XOR2_X1 U1033 ( .A(n1365), .B(G110), .Z(n1363) );
NAND2_X1 U1034 ( .A1(n1366), .A2(n1367), .ZN(n1365) );
NAND2_X1 U1035 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
XOR2_X1 U1036 ( .A(G119), .B(n1370), .Z(n1369) );
XOR2_X1 U1037 ( .A(KEYINPUT48), .B(n1345), .Z(n1368) );
INV_X1 U1038 ( .A(G113), .ZN(n1345) );
XOR2_X1 U1039 ( .A(n1371), .B(KEYINPUT6), .Z(n1366) );
NAND2_X1 U1040 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
XOR2_X1 U1041 ( .A(KEYINPUT48), .B(G113), .Z(n1373) );
XNOR2_X1 U1042 ( .A(G119), .B(n1370), .ZN(n1372) );
NAND2_X1 U1043 ( .A1(n1374), .A2(KEYINPUT18), .ZN(n1360) );
XNOR2_X1 U1044 ( .A(G125), .B(KEYINPUT26), .ZN(n1374) );
XNOR2_X1 U1045 ( .A(n1375), .B(n1195), .ZN(n1310) );
NAND2_X1 U1046 ( .A1(G224), .A2(n1109), .ZN(n1375) );
NOR2_X1 U1047 ( .A1(n1150), .A2(n1376), .ZN(n1135) );
AND2_X1 U1048 ( .A1(G221), .A2(n1149), .ZN(n1376) );
XOR2_X1 U1049 ( .A(n1377), .B(G469), .Z(n1150) );
NAND2_X1 U1050 ( .A1(n1378), .A2(n1358), .ZN(n1377) );
XOR2_X1 U1051 ( .A(n1379), .B(n1380), .Z(n1378) );
XNOR2_X1 U1052 ( .A(n1264), .B(n1257), .ZN(n1380) );
XNOR2_X1 U1053 ( .A(n1381), .B(n1382), .ZN(n1257) );
XOR2_X1 U1054 ( .A(G110), .B(n1383), .Z(n1382) );
AND2_X1 U1055 ( .A1(n1109), .A2(G227), .ZN(n1383) );
XOR2_X1 U1056 ( .A(n1209), .B(n1195), .Z(n1264) );
XOR2_X1 U1057 ( .A(G101), .B(n1384), .Z(n1209) );
XOR2_X1 U1058 ( .A(G107), .B(G104), .Z(n1384) );
XOR2_X1 U1059 ( .A(n1258), .B(KEYINPUT21), .Z(n1379) );
NOR2_X1 U1060 ( .A1(n1159), .A2(n1338), .ZN(n1120) );
INV_X1 U1061 ( .A(n1168), .ZN(n1338) );
XOR2_X1 U1062 ( .A(n1385), .B(G475), .Z(n1168) );
NAND2_X1 U1063 ( .A1(n1225), .A2(n1358), .ZN(n1385) );
XOR2_X1 U1064 ( .A(n1386), .B(n1387), .Z(n1225) );
XOR2_X1 U1065 ( .A(n1388), .B(n1389), .Z(n1387) );
XOR2_X1 U1066 ( .A(G146), .B(G131), .Z(n1389) );
NOR3_X1 U1067 ( .A1(KEYINPUT44), .A2(n1390), .A3(n1391), .ZN(n1388) );
NOR4_X1 U1068 ( .A1(n1317), .A2(n1392), .A3(G953), .A4(n1393), .ZN(n1391) );
INV_X1 U1069 ( .A(G143), .ZN(n1317) );
NOR2_X1 U1070 ( .A1(G143), .A2(n1394), .ZN(n1390) );
NOR3_X1 U1071 ( .A1(n1392), .A2(G953), .A3(n1393), .ZN(n1394) );
XOR2_X1 U1072 ( .A(G237), .B(KEYINPUT53), .Z(n1393) );
INV_X1 U1073 ( .A(G214), .ZN(n1392) );
XOR2_X1 U1074 ( .A(n1395), .B(n1190), .Z(n1386) );
XOR2_X1 U1075 ( .A(G140), .B(G125), .Z(n1190) );
NAND2_X1 U1076 ( .A1(KEYINPUT58), .A2(n1396), .ZN(n1395) );
XOR2_X1 U1077 ( .A(n1231), .B(n1397), .Z(n1396) );
NAND2_X1 U1078 ( .A1(n1398), .A2(n1399), .ZN(n1397) );
NAND2_X1 U1079 ( .A1(G113), .A2(n1337), .ZN(n1399) );
XOR2_X1 U1080 ( .A(KEYINPUT24), .B(n1400), .Z(n1398) );
NOR2_X1 U1081 ( .A1(G113), .A2(n1337), .ZN(n1400) );
INV_X1 U1082 ( .A(G104), .ZN(n1231) );
INV_X1 U1083 ( .A(n1321), .ZN(n1159) );
XOR2_X1 U1084 ( .A(n1401), .B(G478), .Z(n1321) );
OR2_X1 U1085 ( .A1(n1217), .A2(G902), .ZN(n1401) );
XNOR2_X1 U1086 ( .A(n1402), .B(n1403), .ZN(n1217) );
XNOR2_X1 U1087 ( .A(n1404), .B(n1405), .ZN(n1403) );
NAND2_X1 U1088 ( .A1(G217), .A2(n1406), .ZN(n1404) );
INV_X1 U1089 ( .A(n1407), .ZN(n1406) );
XOR2_X1 U1090 ( .A(n1408), .B(G134), .Z(n1402) );
NAND2_X1 U1091 ( .A1(n1409), .A2(n1410), .ZN(n1408) );
NAND2_X1 U1092 ( .A1(n1411), .A2(n1412), .ZN(n1410) );
NAND2_X1 U1093 ( .A1(KEYINPUT3), .A2(n1413), .ZN(n1412) );
NAND2_X1 U1094 ( .A1(n1106), .A2(n1414), .ZN(n1413) );
INV_X1 U1095 ( .A(G107), .ZN(n1106) );
NAND2_X1 U1096 ( .A1(G107), .A2(n1415), .ZN(n1409) );
NAND2_X1 U1097 ( .A1(n1414), .A2(n1416), .ZN(n1415) );
NAND2_X1 U1098 ( .A1(KEYINPUT3), .A2(n1417), .ZN(n1416) );
INV_X1 U1099 ( .A(n1411), .ZN(n1417) );
XOR2_X1 U1100 ( .A(n1337), .B(n1370), .Z(n1411) );
INV_X1 U1101 ( .A(G122), .ZN(n1337) );
INV_X1 U1102 ( .A(KEYINPUT2), .ZN(n1414) );
INV_X1 U1103 ( .A(n1123), .ZN(n1323) );
NAND2_X1 U1104 ( .A1(n1125), .A2(n1325), .ZN(n1123) );
INV_X1 U1105 ( .A(n1127), .ZN(n1325) );
NOR2_X1 U1106 ( .A1(n1418), .A2(n1172), .ZN(n1127) );
NOR3_X1 U1107 ( .A1(n1173), .A2(G902), .A3(n1212), .ZN(n1172) );
INV_X1 U1108 ( .A(n1214), .ZN(n1173) );
AND2_X1 U1109 ( .A1(n1419), .A2(n1174), .ZN(n1418) );
NAND2_X1 U1110 ( .A1(n1420), .A2(n1358), .ZN(n1174) );
INV_X1 U1111 ( .A(n1212), .ZN(n1420) );
XOR2_X1 U1112 ( .A(n1421), .B(n1422), .Z(n1212) );
XOR2_X1 U1113 ( .A(n1423), .B(n1424), .Z(n1422) );
XNOR2_X1 U1114 ( .A(n1425), .B(n1426), .ZN(n1424) );
NOR2_X1 U1115 ( .A1(KEYINPUT25), .A2(n1427), .ZN(n1426) );
INV_X1 U1116 ( .A(G110), .ZN(n1427) );
NOR3_X1 U1117 ( .A1(n1407), .A2(KEYINPUT41), .A3(n1428), .ZN(n1425) );
INV_X1 U1118 ( .A(G221), .ZN(n1428) );
NAND2_X1 U1119 ( .A1(G234), .A2(n1109), .ZN(n1407) );
XOR2_X1 U1120 ( .A(n1429), .B(n1430), .Z(n1423) );
NOR2_X1 U1121 ( .A1(KEYINPUT52), .A2(n1431), .ZN(n1430) );
XNOR2_X1 U1122 ( .A(G146), .B(KEYINPUT16), .ZN(n1431) );
NAND2_X1 U1123 ( .A1(n1432), .A2(n1433), .ZN(n1429) );
OR2_X1 U1124 ( .A1(n1434), .A2(G125), .ZN(n1433) );
XOR2_X1 U1125 ( .A(n1435), .B(KEYINPUT42), .Z(n1432) );
NAND2_X1 U1126 ( .A1(G125), .A2(n1434), .ZN(n1435) );
XNOR2_X1 U1127 ( .A(n1258), .B(KEYINPUT56), .ZN(n1434) );
INV_X1 U1128 ( .A(G140), .ZN(n1258) );
XOR2_X1 U1129 ( .A(n1436), .B(n1437), .Z(n1421) );
XOR2_X1 U1130 ( .A(KEYINPUT51), .B(G137), .Z(n1437) );
XNOR2_X1 U1131 ( .A(G128), .B(G119), .ZN(n1436) );
XOR2_X1 U1132 ( .A(n1214), .B(KEYINPUT35), .Z(n1419) );
NAND2_X1 U1133 ( .A1(G217), .A2(n1149), .ZN(n1214) );
NAND2_X1 U1134 ( .A1(G234), .A2(n1355), .ZN(n1149) );
XOR2_X1 U1135 ( .A(n1358), .B(KEYINPUT13), .Z(n1355) );
XOR2_X1 U1136 ( .A(n1164), .B(G472), .Z(n1125) );
NAND2_X1 U1137 ( .A1(n1438), .A2(n1358), .ZN(n1164) );
INV_X1 U1138 ( .A(G902), .ZN(n1358) );
XOR2_X1 U1139 ( .A(n1439), .B(n1440), .Z(n1438) );
NOR2_X1 U1140 ( .A1(KEYINPUT34), .A2(n1441), .ZN(n1440) );
XOR2_X1 U1141 ( .A(n1250), .B(KEYINPUT62), .Z(n1441) );
NAND2_X1 U1142 ( .A1(n1442), .A2(n1240), .ZN(n1250) );
NAND3_X1 U1143 ( .A1(n1443), .A2(n1195), .A3(n1381), .ZN(n1240) );
INV_X1 U1144 ( .A(n1243), .ZN(n1442) );
NAND2_X1 U1145 ( .A1(n1444), .A2(n1445), .ZN(n1243) );
NAND3_X1 U1146 ( .A1(n1249), .A2(n1446), .A3(n1248), .ZN(n1445) );
INV_X1 U1147 ( .A(n1447), .ZN(n1248) );
NAND2_X1 U1148 ( .A1(n1381), .A2(n1195), .ZN(n1446) );
NAND2_X1 U1149 ( .A1(n1447), .A2(n1443), .ZN(n1444) );
INV_X1 U1150 ( .A(n1249), .ZN(n1443) );
XOR2_X1 U1151 ( .A(n1448), .B(n1449), .Z(n1249) );
XOR2_X1 U1152 ( .A(G119), .B(G113), .Z(n1449) );
NAND2_X1 U1153 ( .A1(n1450), .A2(n1370), .ZN(n1448) );
XOR2_X1 U1154 ( .A(G116), .B(KEYINPUT28), .Z(n1370) );
XOR2_X1 U1155 ( .A(KEYINPUT9), .B(KEYINPUT22), .Z(n1450) );
NOR2_X1 U1156 ( .A1(n1195), .A2(n1381), .ZN(n1447) );
AND2_X1 U1157 ( .A1(n1451), .A2(n1452), .ZN(n1381) );
NAND2_X1 U1158 ( .A1(n1198), .A2(G137), .ZN(n1452) );
NAND2_X1 U1159 ( .A1(n1453), .A2(n1197), .ZN(n1451) );
INV_X1 U1160 ( .A(G137), .ZN(n1197) );
XNOR2_X1 U1161 ( .A(n1198), .B(KEYINPUT50), .ZN(n1453) );
XOR2_X1 U1162 ( .A(G131), .B(G134), .Z(n1198) );
XOR2_X1 U1163 ( .A(G146), .B(n1405), .Z(n1195) );
XOR2_X1 U1164 ( .A(G128), .B(G143), .Z(n1405) );
NOR2_X1 U1165 ( .A1(n1454), .A2(n1455), .ZN(n1439) );
XNOR2_X1 U1166 ( .A(KEYINPUT11), .B(n1251), .ZN(n1455) );
OR2_X1 U1167 ( .A1(G101), .A2(n1456), .ZN(n1251) );
AND3_X1 U1168 ( .A1(n1356), .A2(n1109), .A3(G210), .ZN(n1456) );
INV_X1 U1169 ( .A(n1252), .ZN(n1454) );
NAND4_X1 U1170 ( .A1(G210), .A2(G101), .A3(n1356), .A4(n1109), .ZN(n1252) );
INV_X1 U1171 ( .A(G953), .ZN(n1109) );
INV_X1 U1172 ( .A(G237), .ZN(n1356) );
endmodule


