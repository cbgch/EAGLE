//Key = 0011001000100101110000000111110111001001000001111101010000001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379;

XNOR2_X1 U755 ( .A(G107), .B(n1051), .ZN(G9) );
NOR2_X1 U756 ( .A1(n1052), .A2(n1053), .ZN(G75) );
NOR3_X1 U757 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NOR3_X1 U758 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1055) );
NOR2_X1 U759 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR3_X1 U760 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
XNOR2_X1 U761 ( .A(KEYINPUT45), .B(n1065), .ZN(n1062) );
NOR4_X1 U762 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1065), .ZN(n1060) );
NOR2_X1 U763 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR2_X1 U764 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NAND3_X1 U765 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1054) );
NAND4_X1 U766 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1075) );
NOR3_X1 U767 ( .A1(n1065), .A2(n1063), .A3(n1068), .ZN(n1079) );
INV_X1 U768 ( .A(n1080), .ZN(n1063) );
NAND2_X1 U769 ( .A1(n1057), .A2(n1081), .ZN(n1078) );
OR3_X1 U770 ( .A1(n1082), .A2(n1066), .A3(n1059), .ZN(n1081) );
NAND3_X1 U771 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1077) );
XNOR2_X1 U772 ( .A(KEYINPUT2), .B(n1086), .ZN(n1085) );
OR2_X1 U773 ( .A1(n1087), .A2(n1088), .ZN(n1084) );
NAND3_X1 U774 ( .A1(n1089), .A2(n1090), .A3(n1087), .ZN(n1083) );
NAND2_X1 U775 ( .A1(n1082), .A2(n1091), .ZN(n1090) );
NOR2_X1 U776 ( .A1(n1092), .A2(n1093), .ZN(n1082) );
NAND2_X1 U777 ( .A1(n1066), .A2(n1059), .ZN(n1076) );
NOR3_X1 U778 ( .A1(n1094), .A2(G953), .A3(G952), .ZN(n1052) );
INV_X1 U779 ( .A(n1073), .ZN(n1094) );
NAND4_X1 U780 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1073) );
NOR4_X1 U781 ( .A1(n1099), .A2(n1066), .A3(n1100), .A4(n1101), .ZN(n1098) );
NAND3_X1 U782 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1099) );
NAND2_X1 U783 ( .A1(G469), .A2(n1105), .ZN(n1104) );
NOR3_X1 U784 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1097) );
XNOR2_X1 U785 ( .A(n1109), .B(n1110), .ZN(n1108) );
NAND2_X1 U786 ( .A1(KEYINPUT3), .A2(n1111), .ZN(n1109) );
AND2_X1 U787 ( .A1(n1112), .A2(n1113), .ZN(n1107) );
XOR2_X1 U788 ( .A(n1114), .B(KEYINPUT47), .Z(n1106) );
OR2_X1 U789 ( .A1(n1105), .A2(G469), .ZN(n1114) );
XOR2_X1 U790 ( .A(n1115), .B(n1116), .Z(G72) );
NOR2_X1 U791 ( .A1(n1117), .A2(n1074), .ZN(n1116) );
AND2_X1 U792 ( .A1(G227), .A2(G900), .ZN(n1117) );
NAND2_X1 U793 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
NAND3_X1 U794 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
INV_X1 U795 ( .A(n1123), .ZN(n1121) );
OR2_X1 U796 ( .A1(n1122), .A2(n1120), .ZN(n1118) );
XNOR2_X1 U797 ( .A(n1124), .B(n1125), .ZN(n1120) );
XNOR2_X1 U798 ( .A(KEYINPUT36), .B(n1126), .ZN(n1124) );
NOR2_X1 U799 ( .A1(KEYINPUT19), .A2(n1127), .ZN(n1126) );
XOR2_X1 U800 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND2_X1 U801 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
OR2_X1 U802 ( .A1(n1132), .A2(G134), .ZN(n1131) );
NAND2_X1 U803 ( .A1(n1133), .A2(G134), .ZN(n1130) );
XOR2_X1 U804 ( .A(KEYINPUT4), .B(n1132), .Z(n1133) );
NAND2_X1 U805 ( .A1(n1074), .A2(n1134), .ZN(n1122) );
NAND2_X1 U806 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U807 ( .A(KEYINPUT11), .B(n1137), .Z(n1136) );
XOR2_X1 U808 ( .A(n1138), .B(n1139), .Z(G69) );
NOR2_X1 U809 ( .A1(n1140), .A2(n1074), .ZN(n1139) );
AND2_X1 U810 ( .A1(G224), .A2(G898), .ZN(n1140) );
NAND2_X1 U811 ( .A1(n1141), .A2(n1142), .ZN(n1138) );
NAND3_X1 U812 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1142) );
INV_X1 U813 ( .A(n1146), .ZN(n1144) );
OR2_X1 U814 ( .A1(n1143), .A2(n1145), .ZN(n1141) );
NAND2_X1 U815 ( .A1(n1074), .A2(n1147), .ZN(n1145) );
NAND2_X1 U816 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U817 ( .A(n1150), .B(n1151), .Z(n1143) );
XNOR2_X1 U818 ( .A(G122), .B(n1152), .ZN(n1151) );
NAND2_X1 U819 ( .A1(n1153), .A2(n1154), .ZN(n1150) );
NAND2_X1 U820 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U821 ( .A(n1157), .B(KEYINPUT38), .Z(n1153) );
OR2_X1 U822 ( .A1(n1156), .A2(n1155), .ZN(n1157) );
XOR2_X1 U823 ( .A(n1158), .B(KEYINPUT51), .Z(n1155) );
XNOR2_X1 U824 ( .A(n1159), .B(n1160), .ZN(n1156) );
XNOR2_X1 U825 ( .A(G101), .B(G107), .ZN(n1159) );
NOR2_X1 U826 ( .A1(n1161), .A2(n1162), .ZN(G66) );
XOR2_X1 U827 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U828 ( .A(KEYINPUT32), .B(n1165), .Z(n1164) );
NOR2_X1 U829 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NOR2_X1 U830 ( .A1(n1161), .A2(n1168), .ZN(G63) );
XNOR2_X1 U831 ( .A(n1169), .B(n1170), .ZN(n1168) );
NOR2_X1 U832 ( .A1(n1171), .A2(n1167), .ZN(n1170) );
NOR2_X1 U833 ( .A1(n1161), .A2(n1172), .ZN(G60) );
XNOR2_X1 U834 ( .A(n1173), .B(n1174), .ZN(n1172) );
NOR2_X1 U835 ( .A1(n1111), .A2(n1167), .ZN(n1174) );
XNOR2_X1 U836 ( .A(G104), .B(n1175), .ZN(G6) );
NAND3_X1 U837 ( .A1(n1176), .A2(n1080), .A3(n1177), .ZN(n1175) );
XNOR2_X1 U838 ( .A(n1092), .B(KEYINPUT15), .ZN(n1177) );
NOR2_X1 U839 ( .A1(n1161), .A2(n1178), .ZN(G57) );
XOR2_X1 U840 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U841 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U842 ( .A(KEYINPUT25), .B(n1183), .Z(n1179) );
NOR2_X1 U843 ( .A1(n1184), .A2(n1167), .ZN(n1183) );
NOR3_X1 U844 ( .A1(n1161), .A2(n1185), .A3(n1186), .ZN(G54) );
NOR4_X1 U845 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1167), .ZN(n1186) );
INV_X1 U846 ( .A(KEYINPUT33), .ZN(n1188) );
NOR2_X1 U847 ( .A1(n1190), .A2(n1191), .ZN(n1185) );
NOR3_X1 U848 ( .A1(n1167), .A2(n1192), .A3(n1189), .ZN(n1191) );
NOR2_X1 U849 ( .A1(KEYINPUT33), .A2(n1193), .ZN(n1192) );
INV_X1 U850 ( .A(n1187), .ZN(n1190) );
NAND2_X1 U851 ( .A1(KEYINPUT29), .A2(n1193), .ZN(n1187) );
XOR2_X1 U852 ( .A(n1194), .B(n1195), .Z(n1193) );
XNOR2_X1 U853 ( .A(n1196), .B(n1197), .ZN(n1195) );
NOR3_X1 U854 ( .A1(n1198), .A2(KEYINPUT54), .A3(G953), .ZN(n1197) );
NOR2_X1 U855 ( .A1(n1161), .A2(n1199), .ZN(G51) );
XOR2_X1 U856 ( .A(n1200), .B(n1201), .Z(n1199) );
NOR2_X1 U857 ( .A1(n1202), .A2(n1167), .ZN(n1201) );
NAND2_X1 U858 ( .A1(G902), .A2(n1056), .ZN(n1167) );
NAND4_X1 U859 ( .A1(n1203), .A2(n1137), .A3(n1135), .A4(n1148), .ZN(n1056) );
AND4_X1 U860 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1148) );
AND4_X1 U861 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1135) );
NAND3_X1 U862 ( .A1(n1212), .A2(n1072), .A3(n1213), .ZN(n1208) );
XNOR2_X1 U863 ( .A(KEYINPUT35), .B(n1086), .ZN(n1212) );
AND4_X1 U864 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1137) );
XNOR2_X1 U865 ( .A(n1149), .B(KEYINPUT53), .ZN(n1203) );
AND3_X1 U866 ( .A1(n1218), .A2(n1051), .A3(n1219), .ZN(n1149) );
NAND2_X1 U867 ( .A1(n1176), .A2(n1220), .ZN(n1219) );
NAND2_X1 U868 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NAND2_X1 U869 ( .A1(n1092), .A2(n1080), .ZN(n1222) );
OR2_X1 U870 ( .A1(n1057), .A2(n1223), .ZN(n1221) );
NAND3_X1 U871 ( .A1(n1080), .A2(n1093), .A3(n1176), .ZN(n1051) );
NOR2_X1 U872 ( .A1(n1224), .A2(n1225), .ZN(n1200) );
XOR2_X1 U873 ( .A(KEYINPUT50), .B(n1226), .Z(n1225) );
NOR2_X1 U874 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
XOR2_X1 U875 ( .A(KEYINPUT20), .B(n1229), .Z(n1228) );
AND2_X1 U876 ( .A1(n1227), .A2(n1229), .ZN(n1224) );
XOR2_X1 U877 ( .A(n1230), .B(n1231), .Z(n1229) );
XNOR2_X1 U878 ( .A(n1232), .B(n1233), .ZN(n1231) );
NOR2_X1 U879 ( .A1(n1074), .A2(G952), .ZN(n1161) );
XNOR2_X1 U880 ( .A(G146), .B(n1234), .ZN(G48) );
NAND3_X1 U881 ( .A1(n1235), .A2(n1072), .A3(n1213), .ZN(n1234) );
XNOR2_X1 U882 ( .A(G143), .B(n1211), .ZN(G45) );
NAND4_X1 U883 ( .A1(n1236), .A2(n1237), .A3(n1070), .A4(n1238), .ZN(n1211) );
NOR3_X1 U884 ( .A1(n1086), .A2(n1239), .A3(n1096), .ZN(n1238) );
INV_X1 U885 ( .A(n1240), .ZN(n1096) );
XOR2_X1 U886 ( .A(G140), .B(n1241), .Z(G42) );
NOR2_X1 U887 ( .A1(KEYINPUT40), .A2(n1209), .ZN(n1241) );
NAND4_X1 U888 ( .A1(n1242), .A2(n1092), .A3(n1095), .A4(n1243), .ZN(n1209) );
XNOR2_X1 U889 ( .A(G137), .B(n1210), .ZN(G39) );
NAND3_X1 U890 ( .A1(n1242), .A2(n1072), .A3(n1244), .ZN(n1210) );
XNOR2_X1 U891 ( .A(G134), .B(n1214), .ZN(G36) );
NAND3_X1 U892 ( .A1(n1242), .A2(n1093), .A3(n1070), .ZN(n1214) );
XNOR2_X1 U893 ( .A(G131), .B(n1215), .ZN(G33) );
NAND3_X1 U894 ( .A1(n1242), .A2(n1092), .A3(n1070), .ZN(n1215) );
NOR4_X1 U895 ( .A1(n1068), .A2(n1086), .A3(n1239), .A4(n1066), .ZN(n1242) );
INV_X1 U896 ( .A(n1245), .ZN(n1068) );
XNOR2_X1 U897 ( .A(G128), .B(n1216), .ZN(G30) );
NAND4_X1 U898 ( .A1(n1246), .A2(n1093), .A3(n1235), .A4(n1072), .ZN(n1216) );
XNOR2_X1 U899 ( .A(n1247), .B(n1248), .ZN(G3) );
NOR4_X1 U900 ( .A1(KEYINPUT42), .A2(n1249), .A3(n1223), .A4(n1057), .ZN(n1248) );
XNOR2_X1 U901 ( .A(G125), .B(n1217), .ZN(G27) );
NAND3_X1 U902 ( .A1(n1095), .A2(n1213), .A3(n1250), .ZN(n1217) );
AND2_X1 U903 ( .A1(n1092), .A2(n1246), .ZN(n1213) );
NOR3_X1 U904 ( .A1(n1239), .A2(n1071), .A3(n1064), .ZN(n1246) );
AND2_X1 U905 ( .A1(n1065), .A2(n1251), .ZN(n1239) );
NAND3_X1 U906 ( .A1(G902), .A2(n1252), .A3(n1123), .ZN(n1251) );
NOR2_X1 U907 ( .A1(n1074), .A2(G900), .ZN(n1123) );
XOR2_X1 U908 ( .A(G122), .B(n1253), .Z(G24) );
NOR2_X1 U909 ( .A1(KEYINPUT30), .A2(n1204), .ZN(n1253) );
NAND4_X1 U910 ( .A1(n1254), .A2(n1080), .A3(n1237), .A4(n1240), .ZN(n1204) );
NOR2_X1 U911 ( .A1(n1243), .A2(n1072), .ZN(n1080) );
XNOR2_X1 U912 ( .A(n1255), .B(n1205), .ZN(G21) );
NAND3_X1 U913 ( .A1(n1244), .A2(n1072), .A3(n1254), .ZN(n1205) );
NAND2_X1 U914 ( .A1(KEYINPUT27), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U915 ( .A(G116), .B(n1257), .ZN(G18) );
NAND2_X1 U916 ( .A1(KEYINPUT17), .A2(n1258), .ZN(n1257) );
INV_X1 U917 ( .A(n1206), .ZN(n1258) );
NAND3_X1 U918 ( .A1(n1070), .A2(n1093), .A3(n1254), .ZN(n1206) );
AND3_X1 U919 ( .A1(n1236), .A2(n1259), .A3(n1250), .ZN(n1254) );
INV_X1 U920 ( .A(n1059), .ZN(n1250) );
INV_X1 U921 ( .A(n1064), .ZN(n1236) );
XOR2_X1 U922 ( .A(n1260), .B(KEYINPUT49), .Z(n1064) );
AND2_X1 U923 ( .A1(n1261), .A2(n1240), .ZN(n1093) );
XNOR2_X1 U924 ( .A(KEYINPUT52), .B(n1237), .ZN(n1261) );
NAND2_X1 U925 ( .A1(n1262), .A2(n1263), .ZN(G15) );
NAND2_X1 U926 ( .A1(G113), .A2(n1207), .ZN(n1263) );
XOR2_X1 U927 ( .A(n1264), .B(KEYINPUT56), .Z(n1262) );
OR2_X1 U928 ( .A1(n1207), .A2(G113), .ZN(n1264) );
NAND4_X1 U929 ( .A1(n1260), .A2(n1259), .A3(n1092), .A4(n1265), .ZN(n1207) );
NOR2_X1 U930 ( .A1(n1059), .A2(n1223), .ZN(n1265) );
INV_X1 U931 ( .A(n1070), .ZN(n1223) );
NOR2_X1 U932 ( .A1(n1243), .A2(n1095), .ZN(n1070) );
NAND2_X1 U933 ( .A1(n1089), .A2(n1087), .ZN(n1059) );
XNOR2_X1 U934 ( .A(n1088), .B(KEYINPUT18), .ZN(n1089) );
AND2_X1 U935 ( .A1(n1266), .A2(n1237), .ZN(n1092) );
INV_X1 U936 ( .A(n1267), .ZN(n1237) );
XNOR2_X1 U937 ( .A(G110), .B(n1218), .ZN(G12) );
NAND3_X1 U938 ( .A1(n1095), .A2(n1176), .A3(n1244), .ZN(n1218) );
NOR2_X1 U939 ( .A1(n1057), .A2(n1071), .ZN(n1244) );
INV_X1 U940 ( .A(n1243), .ZN(n1071) );
NAND2_X1 U941 ( .A1(n1268), .A2(n1102), .ZN(n1243) );
NAND2_X1 U942 ( .A1(n1269), .A2(n1270), .ZN(n1102) );
XOR2_X1 U943 ( .A(n1103), .B(KEYINPUT14), .Z(n1268) );
OR2_X1 U944 ( .A1(n1270), .A2(n1269), .ZN(n1103) );
INV_X1 U945 ( .A(n1166), .ZN(n1269) );
NAND2_X1 U946 ( .A1(G217), .A2(n1271), .ZN(n1166) );
NAND2_X1 U947 ( .A1(n1163), .A2(n1272), .ZN(n1270) );
XOR2_X1 U948 ( .A(n1273), .B(n1274), .Z(n1163) );
NOR2_X1 U949 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NOR2_X1 U950 ( .A1(n1277), .A2(G137), .ZN(n1276) );
NOR3_X1 U951 ( .A1(n1278), .A2(G953), .A3(n1279), .ZN(n1277) );
NOR4_X1 U952 ( .A1(G953), .A2(n1279), .A3(n1278), .A4(n1280), .ZN(n1275) );
XOR2_X1 U953 ( .A(KEYINPUT48), .B(G137), .Z(n1280) );
INV_X1 U954 ( .A(G221), .ZN(n1278) );
INV_X1 U955 ( .A(G234), .ZN(n1279) );
NAND3_X1 U956 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1273) );
OR2_X1 U957 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NAND2_X1 U958 ( .A1(KEYINPUT63), .A2(n1286), .ZN(n1282) );
NAND2_X1 U959 ( .A1(n1285), .A2(n1287), .ZN(n1286) );
XNOR2_X1 U960 ( .A(KEYINPUT43), .B(n1288), .ZN(n1287) );
NAND2_X1 U961 ( .A1(n1289), .A2(n1290), .ZN(n1281) );
INV_X1 U962 ( .A(KEYINPUT63), .ZN(n1290) );
NAND2_X1 U963 ( .A1(n1291), .A2(n1292), .ZN(n1289) );
NAND2_X1 U964 ( .A1(KEYINPUT43), .A2(n1288), .ZN(n1292) );
INV_X1 U965 ( .A(n1284), .ZN(n1288) );
NAND3_X1 U966 ( .A1(n1285), .A2(n1293), .A3(n1284), .ZN(n1291) );
XNOR2_X1 U967 ( .A(n1294), .B(n1295), .ZN(n1284) );
XNOR2_X1 U968 ( .A(n1296), .B(G119), .ZN(n1295) );
NAND2_X1 U969 ( .A1(KEYINPUT46), .A2(n1152), .ZN(n1294) );
INV_X1 U970 ( .A(G110), .ZN(n1152) );
INV_X1 U971 ( .A(KEYINPUT43), .ZN(n1293) );
XNOR2_X1 U972 ( .A(n1297), .B(G146), .ZN(n1285) );
NAND2_X1 U973 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NAND2_X1 U974 ( .A1(G125), .A2(n1300), .ZN(n1299) );
NAND2_X1 U975 ( .A1(n1301), .A2(n1232), .ZN(n1298) );
XOR2_X1 U976 ( .A(n1300), .B(KEYINPUT16), .Z(n1301) );
XNOR2_X1 U977 ( .A(G140), .B(KEYINPUT39), .ZN(n1300) );
NAND2_X1 U978 ( .A1(n1266), .A2(n1267), .ZN(n1057) );
XNOR2_X1 U979 ( .A(n1110), .B(n1302), .ZN(n1267) );
XNOR2_X1 U980 ( .A(KEYINPUT26), .B(n1111), .ZN(n1302) );
INV_X1 U981 ( .A(G475), .ZN(n1111) );
NAND2_X1 U982 ( .A1(n1303), .A2(n1173), .ZN(n1110) );
XNOR2_X1 U983 ( .A(n1304), .B(n1305), .ZN(n1173) );
XOR2_X1 U984 ( .A(n1306), .B(n1307), .Z(n1305) );
XNOR2_X1 U985 ( .A(G131), .B(n1308), .ZN(n1307) );
NAND2_X1 U986 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
OR2_X1 U987 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U988 ( .A(n1313), .B(KEYINPUT12), .Z(n1309) );
NAND2_X1 U989 ( .A1(n1311), .A2(n1312), .ZN(n1313) );
XOR2_X1 U990 ( .A(G113), .B(n1314), .Z(n1311) );
NOR2_X1 U991 ( .A1(G122), .A2(KEYINPUT23), .ZN(n1314) );
AND2_X1 U992 ( .A1(G214), .A2(n1315), .ZN(n1306) );
XNOR2_X1 U993 ( .A(n1316), .B(n1125), .ZN(n1304) );
XOR2_X1 U994 ( .A(G140), .B(G125), .Z(n1125) );
XNOR2_X1 U995 ( .A(KEYINPUT28), .B(n1272), .ZN(n1303) );
XNOR2_X1 U996 ( .A(n1240), .B(KEYINPUT34), .ZN(n1266) );
XOR2_X1 U997 ( .A(n1317), .B(n1171), .Z(n1240) );
INV_X1 U998 ( .A(G478), .ZN(n1171) );
NAND2_X1 U999 ( .A1(n1169), .A2(n1272), .ZN(n1317) );
XNOR2_X1 U1000 ( .A(n1318), .B(n1319), .ZN(n1169) );
XNOR2_X1 U1001 ( .A(n1320), .B(n1321), .ZN(n1319) );
XOR2_X1 U1002 ( .A(n1322), .B(n1323), .Z(n1321) );
AND3_X1 U1003 ( .A1(G217), .A2(n1074), .A3(G234), .ZN(n1323) );
NOR2_X1 U1004 ( .A1(KEYINPUT0), .A2(n1324), .ZN(n1322) );
INV_X1 U1005 ( .A(G116), .ZN(n1324) );
INV_X1 U1006 ( .A(n1325), .ZN(n1320) );
XNOR2_X1 U1007 ( .A(G128), .B(n1326), .ZN(n1318) );
XNOR2_X1 U1008 ( .A(n1327), .B(G134), .ZN(n1326) );
INV_X1 U1009 ( .A(G143), .ZN(n1327) );
INV_X1 U1010 ( .A(n1249), .ZN(n1176) );
NAND3_X1 U1011 ( .A1(n1260), .A2(n1259), .A3(n1235), .ZN(n1249) );
INV_X1 U1012 ( .A(n1086), .ZN(n1235) );
NAND2_X1 U1013 ( .A1(n1328), .A2(n1088), .ZN(n1086) );
XNOR2_X1 U1014 ( .A(n1105), .B(n1329), .ZN(n1088) );
XNOR2_X1 U1015 ( .A(KEYINPUT58), .B(n1189), .ZN(n1329) );
INV_X1 U1016 ( .A(G469), .ZN(n1189) );
NAND3_X1 U1017 ( .A1(n1330), .A2(n1331), .A3(n1272), .ZN(n1105) );
NAND2_X1 U1018 ( .A1(n1332), .A2(G227), .ZN(n1331) );
NAND2_X1 U1019 ( .A1(n1333), .A2(n1198), .ZN(n1330) );
INV_X1 U1020 ( .A(G227), .ZN(n1198) );
XNOR2_X1 U1021 ( .A(KEYINPUT62), .B(n1332), .ZN(n1333) );
XOR2_X1 U1022 ( .A(n1194), .B(n1334), .Z(n1332) );
NOR2_X1 U1023 ( .A1(KEYINPUT5), .A2(n1196), .ZN(n1334) );
XOR2_X1 U1024 ( .A(n1335), .B(n1336), .Z(n1194) );
XNOR2_X1 U1025 ( .A(n1337), .B(n1128), .ZN(n1336) );
NAND2_X1 U1026 ( .A1(n1338), .A2(n1339), .ZN(n1128) );
NAND2_X1 U1027 ( .A1(n1340), .A2(n1296), .ZN(n1339) );
XOR2_X1 U1028 ( .A(n1341), .B(KEYINPUT6), .Z(n1340) );
NAND2_X1 U1029 ( .A1(G128), .A2(n1342), .ZN(n1338) );
XOR2_X1 U1030 ( .A(n1341), .B(KEYINPUT24), .Z(n1342) );
XNOR2_X1 U1031 ( .A(n1316), .B(KEYINPUT44), .ZN(n1341) );
XOR2_X1 U1032 ( .A(n1343), .B(G140), .Z(n1335) );
NAND2_X1 U1033 ( .A1(KEYINPUT60), .A2(n1344), .ZN(n1343) );
XNOR2_X1 U1034 ( .A(n1345), .B(n1346), .ZN(n1344) );
INV_X1 U1035 ( .A(G107), .ZN(n1345) );
XNOR2_X1 U1036 ( .A(n1101), .B(KEYINPUT61), .ZN(n1328) );
INV_X1 U1037 ( .A(n1087), .ZN(n1101) );
NAND2_X1 U1038 ( .A1(G221), .A2(n1271), .ZN(n1087) );
NAND2_X1 U1039 ( .A1(G234), .A2(n1272), .ZN(n1271) );
NAND2_X1 U1040 ( .A1(n1065), .A2(n1347), .ZN(n1259) );
NAND3_X1 U1041 ( .A1(n1146), .A2(n1252), .A3(G902), .ZN(n1347) );
NOR2_X1 U1042 ( .A1(n1074), .A2(G898), .ZN(n1146) );
NAND3_X1 U1043 ( .A1(n1252), .A2(n1074), .A3(G952), .ZN(n1065) );
NAND2_X1 U1044 ( .A1(G237), .A2(G234), .ZN(n1252) );
NOR2_X1 U1045 ( .A1(n1245), .A2(n1066), .ZN(n1260) );
INV_X1 U1046 ( .A(n1091), .ZN(n1066) );
NAND2_X1 U1047 ( .A1(G214), .A2(n1348), .ZN(n1091) );
NOR2_X1 U1048 ( .A1(n1349), .A2(n1100), .ZN(n1245) );
NOR2_X1 U1049 ( .A1(n1112), .A2(n1113), .ZN(n1100) );
AND2_X1 U1050 ( .A1(n1350), .A2(n1113), .ZN(n1349) );
INV_X1 U1051 ( .A(n1202), .ZN(n1113) );
NAND2_X1 U1052 ( .A1(G210), .A2(n1348), .ZN(n1202) );
NAND2_X1 U1053 ( .A1(n1351), .A2(n1272), .ZN(n1348) );
INV_X1 U1054 ( .A(G237), .ZN(n1351) );
XOR2_X1 U1055 ( .A(n1112), .B(KEYINPUT55), .Z(n1350) );
NAND2_X1 U1056 ( .A1(n1352), .A2(n1272), .ZN(n1112) );
INV_X1 U1057 ( .A(G902), .ZN(n1272) );
XNOR2_X1 U1058 ( .A(n1227), .B(n1353), .ZN(n1352) );
XOR2_X1 U1059 ( .A(n1233), .B(n1354), .Z(n1353) );
NOR2_X1 U1060 ( .A1(KEYINPUT21), .A2(n1355), .ZN(n1354) );
XNOR2_X1 U1061 ( .A(n1232), .B(n1356), .ZN(n1355) );
NOR2_X1 U1062 ( .A1(KEYINPUT9), .A2(n1230), .ZN(n1356) );
INV_X1 U1063 ( .A(G125), .ZN(n1232) );
AND2_X1 U1064 ( .A1(G224), .A2(n1074), .ZN(n1233) );
INV_X1 U1065 ( .A(G953), .ZN(n1074) );
XNOR2_X1 U1066 ( .A(n1357), .B(n1358), .ZN(n1227) );
XOR2_X1 U1067 ( .A(n1337), .B(n1158), .Z(n1358) );
XOR2_X1 U1068 ( .A(n1359), .B(n1360), .Z(n1158) );
NAND3_X1 U1069 ( .A1(n1361), .A2(n1362), .A3(n1363), .ZN(n1359) );
NAND2_X1 U1070 ( .A1(KEYINPUT8), .A2(G119), .ZN(n1363) );
OR3_X1 U1071 ( .A1(n1364), .A2(KEYINPUT8), .A3(n1365), .ZN(n1362) );
NAND2_X1 U1072 ( .A1(n1365), .A2(n1364), .ZN(n1361) );
NAND2_X1 U1073 ( .A1(n1366), .A2(n1256), .ZN(n1364) );
INV_X1 U1074 ( .A(G119), .ZN(n1256) );
XOR2_X1 U1075 ( .A(KEYINPUT41), .B(KEYINPUT31), .Z(n1366) );
XOR2_X1 U1076 ( .A(G101), .B(G110), .Z(n1337) );
XNOR2_X1 U1077 ( .A(n1325), .B(n1160), .ZN(n1357) );
NOR2_X1 U1078 ( .A1(KEYINPUT22), .A2(n1367), .ZN(n1160) );
XOR2_X1 U1079 ( .A(KEYINPUT7), .B(n1346), .Z(n1367) );
XNOR2_X1 U1080 ( .A(n1312), .B(KEYINPUT37), .ZN(n1346) );
INV_X1 U1081 ( .A(G104), .ZN(n1312) );
XOR2_X1 U1082 ( .A(G107), .B(G122), .Z(n1325) );
INV_X1 U1083 ( .A(n1072), .ZN(n1095) );
XOR2_X1 U1084 ( .A(n1368), .B(n1184), .Z(n1072) );
INV_X1 U1085 ( .A(G472), .ZN(n1184) );
NAND2_X1 U1086 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
XOR2_X1 U1087 ( .A(n1371), .B(n1182), .Z(n1370) );
XOR2_X1 U1088 ( .A(n1372), .B(n1373), .Z(n1182) );
XNOR2_X1 U1089 ( .A(n1360), .B(n1374), .ZN(n1373) );
NOR2_X1 U1090 ( .A1(KEYINPUT1), .A2(n1375), .ZN(n1374) );
XNOR2_X1 U1091 ( .A(G119), .B(n1365), .ZN(n1375) );
XOR2_X1 U1092 ( .A(G116), .B(KEYINPUT59), .Z(n1365) );
INV_X1 U1093 ( .A(G113), .ZN(n1360) );
XNOR2_X1 U1094 ( .A(n1230), .B(n1376), .ZN(n1372) );
INV_X1 U1095 ( .A(n1196), .ZN(n1376) );
XNOR2_X1 U1096 ( .A(G134), .B(n1132), .ZN(n1196) );
XOR2_X1 U1097 ( .A(G131), .B(G137), .Z(n1132) );
XNOR2_X1 U1098 ( .A(n1296), .B(n1316), .ZN(n1230) );
XOR2_X1 U1099 ( .A(G143), .B(G146), .Z(n1316) );
INV_X1 U1100 ( .A(G128), .ZN(n1296) );
NAND2_X1 U1101 ( .A1(n1377), .A2(n1378), .ZN(n1371) );
OR2_X1 U1102 ( .A1(KEYINPUT10), .A2(n1181), .ZN(n1378) );
NAND2_X1 U1103 ( .A1(KEYINPUT13), .A2(n1181), .ZN(n1377) );
XNOR2_X1 U1104 ( .A(n1379), .B(n1247), .ZN(n1181) );
INV_X1 U1105 ( .A(G101), .ZN(n1247) );
NAND2_X1 U1106 ( .A1(n1315), .A2(G210), .ZN(n1379) );
NOR2_X1 U1107 ( .A1(G953), .A2(G237), .ZN(n1315) );
XNOR2_X1 U1108 ( .A(G902), .B(KEYINPUT57), .ZN(n1369) );
endmodule


