//Key = 0101011100011110001000011010000011110101110001000000100110100111


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
n2339, n2340;

OR2_X1 U1308 ( .A1(n2340), .A2(n1908), .ZN(U280) );
INV_X2 U1309 ( .A(U280), .ZN(n1759) );
AND2_X2 U1310 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1783), .ZN(n1908) );
NAND2_X1 U1311 ( .A1(n1760), .A2(n1761), .ZN(U344) );
NAND2_X1 U1312 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1762), .ZN(n1761) );
NAND2_X1 U1313 ( .A1(n1763), .A2(DATA_IN_7_), .ZN(n1760) );
NAND2_X1 U1314 ( .A1(n1764), .A2(n1765), .ZN(U343) );
NAND2_X1 U1315 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1766), .ZN(n1765) );
XNOR2_X1 U1316 ( .A(KEYINPUT1), .B(n1762), .ZN(n1766) );
NAND2_X1 U1317 ( .A1(n1763), .A2(DATA_IN_6_), .ZN(n1764) );
NAND2_X1 U1318 ( .A1(n1767), .A2(n1768), .ZN(U342) );
NAND2_X1 U1319 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1762), .ZN(n1768) );
NAND2_X1 U1320 ( .A1(n1763), .A2(DATA_IN_5_), .ZN(n1767) );
NAND2_X1 U1321 ( .A1(n1769), .A2(n1770), .ZN(U341) );
NAND2_X1 U1322 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1762), .ZN(n1770) );
NAND2_X1 U1323 ( .A1(n1763), .A2(DATA_IN_4_), .ZN(n1769) );
NAND2_X1 U1324 ( .A1(n1771), .A2(n1772), .ZN(U340) );
NAND2_X1 U1325 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1762), .ZN(n1772) );
NAND2_X1 U1326 ( .A1(n1763), .A2(DATA_IN_3_), .ZN(n1771) );
NAND2_X1 U1327 ( .A1(n1773), .A2(n1774), .ZN(U339) );
NAND2_X1 U1328 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1762), .ZN(n1774) );
NAND2_X1 U1329 ( .A1(n1763), .A2(DATA_IN_2_), .ZN(n1773) );
NAND2_X1 U1330 ( .A1(n1775), .A2(n1776), .ZN(U338) );
NAND2_X1 U1331 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1762), .ZN(n1776) );
NAND2_X1 U1332 ( .A1(n1777), .A2(n1763), .ZN(n1775) );
XNOR2_X1 U1333 ( .A(DATA_IN_1_), .B(KEYINPUT23), .ZN(n1777) );
NAND2_X1 U1334 ( .A1(n1778), .A2(n1779), .ZN(U337) );
NAND2_X1 U1335 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1762), .ZN(n1779) );
NAND2_X1 U1336 ( .A1(n1763), .A2(DATA_IN_0_), .ZN(n1778) );
INV_X1 U1337 ( .A(n1762), .ZN(n1763) );
NAND2_X1 U1338 ( .A1(n1780), .A2(n1781), .ZN(n1762) );
NAND3_X1 U1339 ( .A1(n1782), .A2(n1783), .A3(n1784), .ZN(n1781) );
NAND2_X1 U1340 ( .A1(n1785), .A2(n1786), .ZN(U336) );
NAND2_X1 U1341 ( .A1(n1787), .A2(DATA_IN_7_), .ZN(n1786) );
NAND2_X1 U1342 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1788), .ZN(n1785) );
NAND2_X1 U1343 ( .A1(n1789), .A2(n1790), .ZN(U335) );
NAND2_X1 U1344 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1788), .ZN(n1790) );
XOR2_X1 U1345 ( .A(n1791), .B(KEYINPUT16), .Z(n1789) );
NAND2_X1 U1346 ( .A1(n1787), .A2(DATA_IN_6_), .ZN(n1791) );
NAND2_X1 U1347 ( .A1(n1792), .A2(n1793), .ZN(U334) );
NAND2_X1 U1348 ( .A1(n1787), .A2(DATA_IN_5_), .ZN(n1793) );
NAND2_X1 U1349 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1788), .ZN(n1792) );
NAND2_X1 U1350 ( .A1(n1794), .A2(n1795), .ZN(U333) );
NAND2_X1 U1351 ( .A1(n1787), .A2(DATA_IN_4_), .ZN(n1795) );
NAND2_X1 U1352 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1788), .ZN(n1794) );
NAND2_X1 U1353 ( .A1(n1796), .A2(n1797), .ZN(U332) );
NAND2_X1 U1354 ( .A1(n1787), .A2(DATA_IN_3_), .ZN(n1797) );
NAND2_X1 U1355 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1788), .ZN(n1796) );
NAND2_X1 U1356 ( .A1(n1798), .A2(n1799), .ZN(U331) );
NAND2_X1 U1357 ( .A1(n1787), .A2(DATA_IN_2_), .ZN(n1799) );
NAND2_X1 U1358 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1788), .ZN(n1798) );
NAND2_X1 U1359 ( .A1(n1800), .A2(n1801), .ZN(U330) );
NAND2_X1 U1360 ( .A1(n1787), .A2(DATA_IN_1_), .ZN(n1801) );
NAND2_X1 U1361 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1788), .ZN(n1800) );
NAND2_X1 U1362 ( .A1(n1802), .A2(n1803), .ZN(U329) );
NAND2_X1 U1363 ( .A1(n1787), .A2(DATA_IN_0_), .ZN(n1803) );
AND2_X1 U1364 ( .A1(n1804), .A2(n1780), .ZN(n1787) );
NAND2_X1 U1365 ( .A1(n1783), .A2(n1805), .ZN(n1804) );
NAND2_X1 U1366 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1788), .ZN(n1802) );
NAND2_X1 U1367 ( .A1(n1806), .A2(n1780), .ZN(n1788) );
XOR2_X1 U1368 ( .A(KEYINPUT14), .B(n1807), .Z(n1806) );
NOR2_X1 U1369 ( .A1(n1808), .A2(n1809), .ZN(n1807) );
XNOR2_X1 U1370 ( .A(n1783), .B(KEYINPUT48), .ZN(n1809) );
INV_X1 U1371 ( .A(n1805), .ZN(n1808) );
NAND3_X1 U1372 ( .A1(n1784), .A2(n1782), .A3(n1810), .ZN(n1805) );
NAND2_X1 U1373 ( .A1(n1811), .A2(n1812), .ZN(n1810) );
NAND3_X1 U1374 ( .A1(n1813), .A2(n1814), .A3(n1815), .ZN(n1812) );
NAND2_X1 U1375 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1816), .ZN(n1815) );
NAND3_X1 U1376 ( .A1(n1817), .A2(n1818), .A3(n1819), .ZN(n1814) );
XOR2_X1 U1377 ( .A(n1820), .B(KEYINPUT46), .Z(n1819) );
NAND3_X1 U1378 ( .A1(n1821), .A2(n1822), .A3(n1823), .ZN(n1820) );
NAND2_X1 U1379 ( .A1(DATA_IN_5_), .A2(n1824), .ZN(n1823) );
NAND3_X1 U1380 ( .A1(n1825), .A2(n1826), .A3(n1827), .ZN(n1822) );
NAND2_X1 U1381 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1828), .ZN(n1827) );
NAND3_X1 U1382 ( .A1(n1829), .A2(n1830), .A3(n1831), .ZN(n1826) );
NAND2_X1 U1383 ( .A1(n1832), .A2(DATA_IN_3_), .ZN(n1831) );
XNOR2_X1 U1384 ( .A(RMIN_REG_3__SCAN_IN), .B(KEYINPUT51), .ZN(n1832) );
NAND3_X1 U1385 ( .A1(n1833), .A2(n1834), .A3(n1835), .ZN(n1830) );
NAND2_X1 U1386 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1836), .ZN(n1835) );
NAND3_X1 U1387 ( .A1(n1837), .A2(n1838), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1834) );
NAND2_X1 U1388 ( .A1(DATA_IN_1_), .A2(n1839), .ZN(n1837) );
NAND2_X1 U1389 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1840), .ZN(n1833) );
NAND2_X1 U1390 ( .A1(n1841), .A2(DATA_IN_2_), .ZN(n1829) );
XNOR2_X1 U1391 ( .A(RMIN_REG_2__SCAN_IN), .B(KEYINPUT60), .ZN(n1841) );
NAND2_X1 U1392 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1842), .ZN(n1825) );
XNOR2_X1 U1393 ( .A(KEYINPUT63), .B(n1843), .ZN(n1842) );
NAND2_X1 U1394 ( .A1(DATA_IN_4_), .A2(n1844), .ZN(n1821) );
NAND2_X1 U1395 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1845), .ZN(n1818) );
NAND2_X1 U1396 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1846), .ZN(n1817) );
NAND2_X1 U1397 ( .A1(n1847), .A2(n1848), .ZN(n1813) );
XNOR2_X1 U1398 ( .A(DATA_IN_6_), .B(KEYINPUT58), .ZN(n1847) );
NAND2_X1 U1399 ( .A1(DATA_IN_7_), .A2(n1849), .ZN(n1811) );
NAND3_X1 U1400 ( .A1(n1850), .A2(n1851), .A3(n1852), .ZN(n1782) );
NAND2_X1 U1401 ( .A1(DATA_IN_7_), .A2(n1853), .ZN(n1852) );
NAND3_X1 U1402 ( .A1(n1854), .A2(n1855), .A3(n1856), .ZN(n1851) );
NAND2_X1 U1403 ( .A1(DATA_IN_6_), .A2(n1857), .ZN(n1856) );
NAND3_X1 U1404 ( .A1(n1858), .A2(n1859), .A3(n1860), .ZN(n1855) );
NAND2_X1 U1405 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1828), .ZN(n1860) );
INV_X1 U1406 ( .A(DATA_IN_4_), .ZN(n1828) );
NAND3_X1 U1407 ( .A1(n1861), .A2(n1862), .A3(n1863), .ZN(n1859) );
NAND2_X1 U1408 ( .A1(DATA_IN_4_), .A2(n1864), .ZN(n1863) );
NAND3_X1 U1409 ( .A1(n1865), .A2(n1866), .A3(n1867), .ZN(n1862) );
NAND2_X1 U1410 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1843), .ZN(n1867) );
NAND3_X1 U1411 ( .A1(n1868), .A2(n1869), .A3(n1870), .ZN(n1866) );
XOR2_X1 U1412 ( .A(KEYINPUT45), .B(n1871), .Z(n1870) );
NOR2_X1 U1413 ( .A1(n1836), .A2(n1872), .ZN(n1871) );
XNOR2_X1 U1414 ( .A(n1873), .B(KEYINPUT43), .ZN(n1872) );
NAND3_X1 U1415 ( .A1(n1874), .A2(n1875), .A3(DATA_IN_0_), .ZN(n1869) );
NAND2_X1 U1416 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1840), .ZN(n1874) );
NAND2_X1 U1417 ( .A1(n1876), .A2(DATA_IN_1_), .ZN(n1868) );
XNOR2_X1 U1418 ( .A(RMAX_REG_1__SCAN_IN), .B(KEYINPUT8), .ZN(n1876) );
NAND2_X1 U1419 ( .A1(n1877), .A2(RMAX_REG_2__SCAN_IN), .ZN(n1865) );
XNOR2_X1 U1420 ( .A(DATA_IN_2_), .B(KEYINPUT36), .ZN(n1877) );
NAND2_X1 U1421 ( .A1(DATA_IN_3_), .A2(n1878), .ZN(n1861) );
NAND2_X1 U1422 ( .A1(n1879), .A2(RMAX_REG_5__SCAN_IN), .ZN(n1858) );
XNOR2_X1 U1423 ( .A(DATA_IN_5_), .B(KEYINPUT10), .ZN(n1879) );
NAND2_X1 U1424 ( .A1(n1880), .A2(DATA_IN_5_), .ZN(n1854) );
XNOR2_X1 U1425 ( .A(RMAX_REG_5__SCAN_IN), .B(KEYINPUT9), .ZN(n1880) );
NAND2_X1 U1426 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1846), .ZN(n1850) );
NAND2_X1 U1427 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1816), .ZN(n1784) );
NAND2_X1 U1428 ( .A1(n1881), .A2(n1882), .ZN(U328) );
NAND2_X1 U1429 ( .A1(n1883), .A2(DATA_IN_7_), .ZN(n1882) );
NAND2_X1 U1430 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1884), .ZN(n1881) );
NAND2_X1 U1431 ( .A1(n1885), .A2(n1886), .ZN(U327) );
NAND2_X1 U1432 ( .A1(n1883), .A2(DATA_IN_6_), .ZN(n1886) );
NAND2_X1 U1433 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1884), .ZN(n1885) );
NAND2_X1 U1434 ( .A1(n1887), .A2(n1888), .ZN(U326) );
NAND2_X1 U1435 ( .A1(n1883), .A2(DATA_IN_5_), .ZN(n1888) );
NAND2_X1 U1436 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1884), .ZN(n1887) );
NAND2_X1 U1437 ( .A1(n1889), .A2(n1890), .ZN(U325) );
NAND2_X1 U1438 ( .A1(n1891), .A2(DATA_IN_4_), .ZN(n1890) );
XNOR2_X1 U1439 ( .A(n1883), .B(KEYINPUT24), .ZN(n1891) );
XOR2_X1 U1440 ( .A(KEYINPUT6), .B(n1892), .Z(n1889) );
AND2_X1 U1441 ( .A1(n1884), .A2(RLAST_REG_4__SCAN_IN), .ZN(n1892) );
NAND2_X1 U1442 ( .A1(n1893), .A2(n1894), .ZN(U324) );
NAND2_X1 U1443 ( .A1(n1883), .A2(DATA_IN_3_), .ZN(n1894) );
NAND2_X1 U1444 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1884), .ZN(n1893) );
NAND2_X1 U1445 ( .A1(n1895), .A2(n1896), .ZN(U323) );
NAND2_X1 U1446 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1897), .ZN(n1896) );
XNOR2_X1 U1447 ( .A(KEYINPUT11), .B(n1884), .ZN(n1897) );
NAND2_X1 U1448 ( .A1(n1883), .A2(DATA_IN_2_), .ZN(n1895) );
NAND2_X1 U1449 ( .A1(n1898), .A2(n1899), .ZN(U322) );
NAND2_X1 U1450 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1884), .ZN(n1899) );
XOR2_X1 U1451 ( .A(KEYINPUT40), .B(n1900), .Z(n1898) );
NOR2_X1 U1452 ( .A1(n1840), .A2(n1901), .ZN(n1900) );
NAND2_X1 U1453 ( .A1(n1902), .A2(n1903), .ZN(U321) );
NAND2_X1 U1454 ( .A1(n1883), .A2(DATA_IN_0_), .ZN(n1903) );
INV_X1 U1455 ( .A(n1901), .ZN(n1883) );
NAND2_X1 U1456 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1904), .ZN(n1901) );
NAND2_X1 U1457 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1884), .ZN(n1902) );
NAND2_X1 U1458 ( .A1(n1780), .A2(n1904), .ZN(n1884) );
NAND2_X1 U1459 ( .A1(n1905), .A2(n1783), .ZN(n1904) );
INV_X1 U1460 ( .A(U375), .ZN(n1780) );
NOR2_X1 U1461 ( .A1(STATO_REG_0__SCAN_IN), .A2(STATO_REG_1__SCAN_IN), .ZN(U375) );
NAND2_X1 U1462 ( .A1(n1906), .A2(n1907), .ZN(U320) );
NAND2_X1 U1463 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1759), .ZN(n1907) );
NAND2_X1 U1464 ( .A1(n1908), .A2(DATA_IN_7_), .ZN(n1906) );
NAND2_X1 U1465 ( .A1(n1909), .A2(n1910), .ZN(U319) );
NAND2_X1 U1466 ( .A1(n1911), .A2(n1908), .ZN(n1910) );
XNOR2_X1 U1467 ( .A(DATA_IN_6_), .B(KEYINPUT18), .ZN(n1911) );
NAND2_X1 U1468 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1759), .ZN(n1909) );
NAND2_X1 U1469 ( .A1(n1912), .A2(n1913), .ZN(U318) );
NAND2_X1 U1470 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1759), .ZN(n1913) );
NAND2_X1 U1471 ( .A1(n1908), .A2(DATA_IN_5_), .ZN(n1912) );
NAND2_X1 U1472 ( .A1(n1914), .A2(n1915), .ZN(U317) );
NAND2_X1 U1473 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1759), .ZN(n1915) );
NAND2_X1 U1474 ( .A1(n1908), .A2(DATA_IN_4_), .ZN(n1914) );
NAND2_X1 U1475 ( .A1(n1916), .A2(n1917), .ZN(U316) );
NAND2_X1 U1476 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1759), .ZN(n1917) );
NAND2_X1 U1477 ( .A1(n1908), .A2(DATA_IN_3_), .ZN(n1916) );
NAND2_X1 U1478 ( .A1(n1918), .A2(n1919), .ZN(U315) );
NAND2_X1 U1479 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1759), .ZN(n1919) );
NAND2_X1 U1480 ( .A1(n1908), .A2(DATA_IN_2_), .ZN(n1918) );
NAND2_X1 U1481 ( .A1(n1920), .A2(n1921), .ZN(U314) );
NAND2_X1 U1482 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1759), .ZN(n1921) );
NAND2_X1 U1483 ( .A1(n1908), .A2(DATA_IN_1_), .ZN(n1920) );
NAND2_X1 U1484 ( .A1(n1922), .A2(n1923), .ZN(U313) );
NAND2_X1 U1485 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1759), .ZN(n1923) );
NAND2_X1 U1486 ( .A1(n1908), .A2(DATA_IN_0_), .ZN(n1922) );
NAND2_X1 U1487 ( .A1(n1924), .A2(n1925), .ZN(U312) );
NAND2_X1 U1488 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1759), .ZN(n1925) );
NAND2_X1 U1489 ( .A1(n1908), .A2(REG1_REG_7__SCAN_IN), .ZN(n1924) );
NAND2_X1 U1490 ( .A1(n1926), .A2(n1927), .ZN(U311) );
NAND2_X1 U1491 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1759), .ZN(n1927) );
NAND2_X1 U1492 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1908), .ZN(n1926) );
NAND2_X1 U1493 ( .A1(n1928), .A2(n1929), .ZN(U310) );
NAND2_X1 U1494 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1759), .ZN(n1929) );
NAND2_X1 U1495 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1908), .ZN(n1928) );
NAND2_X1 U1496 ( .A1(n1930), .A2(n1931), .ZN(U309) );
NAND2_X1 U1497 ( .A1(n1932), .A2(n1908), .ZN(n1931) );
XNOR2_X1 U1498 ( .A(REG1_REG_4__SCAN_IN), .B(KEYINPUT61), .ZN(n1932) );
XOR2_X1 U1499 ( .A(n1933), .B(KEYINPUT53), .Z(n1930) );
NAND2_X1 U1500 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1759), .ZN(n1933) );
NAND2_X1 U1501 ( .A1(n1934), .A2(n1935), .ZN(U308) );
NAND2_X1 U1502 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1759), .ZN(n1935) );
NAND2_X1 U1503 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1908), .ZN(n1934) );
NAND2_X1 U1504 ( .A1(n1936), .A2(n1937), .ZN(U307) );
NAND2_X1 U1505 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1759), .ZN(n1937) );
NAND2_X1 U1506 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1908), .ZN(n1936) );
NAND2_X1 U1507 ( .A1(n1938), .A2(n1939), .ZN(U306) );
NAND2_X1 U1508 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1759), .ZN(n1939) );
NAND2_X1 U1509 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1908), .ZN(n1938) );
NAND2_X1 U1510 ( .A1(n1940), .A2(n1941), .ZN(U305) );
NAND2_X1 U1511 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1759), .ZN(n1941) );
NAND2_X1 U1512 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1908), .ZN(n1940) );
NAND2_X1 U1513 ( .A1(n1942), .A2(n1943), .ZN(U304) );
NAND2_X1 U1514 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1759), .ZN(n1943) );
NAND2_X1 U1515 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1908), .ZN(n1942) );
NAND2_X1 U1516 ( .A1(n1944), .A2(n1945), .ZN(U303) );
NAND2_X1 U1517 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1759), .ZN(n1945) );
NAND2_X1 U1518 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1908), .ZN(n1944) );
NAND2_X1 U1519 ( .A1(n1946), .A2(n1947), .ZN(U302) );
NAND2_X1 U1520 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1759), .ZN(n1947) );
NAND2_X1 U1521 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1908), .ZN(n1946) );
NAND2_X1 U1522 ( .A1(n1948), .A2(n1949), .ZN(U301) );
NAND2_X1 U1523 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1759), .ZN(n1949) );
NAND2_X1 U1524 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1908), .ZN(n1948) );
NAND2_X1 U1525 ( .A1(n1950), .A2(n1951), .ZN(U300) );
NAND2_X1 U1526 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1759), .ZN(n1951) );
NAND2_X1 U1527 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1908), .ZN(n1950) );
NAND2_X1 U1528 ( .A1(n1952), .A2(n1953), .ZN(U299) );
NAND2_X1 U1529 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1759), .ZN(n1953) );
NAND2_X1 U1530 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1908), .ZN(n1952) );
NAND2_X1 U1531 ( .A1(n1954), .A2(n1955), .ZN(U298) );
NAND2_X1 U1532 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1759), .ZN(n1955) );
NAND2_X1 U1533 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1908), .ZN(n1954) );
NAND2_X1 U1534 ( .A1(n1956), .A2(n1957), .ZN(U297) );
NAND2_X1 U1535 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1759), .ZN(n1957) );
NAND2_X1 U1536 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1908), .ZN(n1956) );
NAND2_X1 U1537 ( .A1(n1958), .A2(n1959), .ZN(U296) );
NAND2_X1 U1538 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1759), .ZN(n1959) );
NAND2_X1 U1539 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1908), .ZN(n1958) );
NAND2_X1 U1540 ( .A1(n1960), .A2(n1961), .ZN(U295) );
NAND2_X1 U1541 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1759), .ZN(n1961) );
NAND2_X1 U1542 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1908), .ZN(n1960) );
NAND2_X1 U1543 ( .A1(n1962), .A2(n1963), .ZN(U294) );
NAND2_X1 U1544 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1759), .ZN(n1963) );
NAND2_X1 U1545 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1908), .ZN(n1962) );
NAND2_X1 U1546 ( .A1(n1964), .A2(n1965), .ZN(U293) );
NAND2_X1 U1547 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1759), .ZN(n1965) );
NAND2_X1 U1548 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1908), .ZN(n1964) );
NAND2_X1 U1549 ( .A1(n1966), .A2(n1967), .ZN(U292) );
NAND2_X1 U1550 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1759), .ZN(n1967) );
NAND2_X1 U1551 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1908), .ZN(n1966) );
NAND2_X1 U1552 ( .A1(n1968), .A2(n1969), .ZN(U291) );
NAND2_X1 U1553 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1759), .ZN(n1969) );
NAND2_X1 U1554 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1908), .ZN(n1968) );
NAND2_X1 U1555 ( .A1(n1970), .A2(n1971), .ZN(U290) );
NAND2_X1 U1556 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1759), .ZN(n1971) );
NAND2_X1 U1557 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1908), .ZN(n1970) );
NAND2_X1 U1558 ( .A1(n1972), .A2(n1973), .ZN(U289) );
NAND2_X1 U1559 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1759), .ZN(n1973) );
NAND2_X1 U1560 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1908), .ZN(n1972) );
NAND4_X1 U1561 ( .A1(n1974), .A2(n1975), .A3(n1976), .A4(n1977), .ZN(U288));
NAND2_X1 U1562 ( .A1(n1978), .A2(REG4_REG_7__SCAN_IN), .ZN(n1977) );
NAND2_X1 U1563 ( .A1(n1979), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1976) );
NAND2_X1 U1564 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1759), .ZN(n1975) );
NAND4_X1 U1565 ( .A1(n1980), .A2(n1981), .A3(n1974), .A4(n1982), .ZN(U287));
NOR3_X1 U1566 ( .A1(n1983), .A2(n1984), .A3(n1985), .ZN(n1982) );
NOR3_X1 U1567 ( .A1(n1986), .A2(n1987), .A3(n1988), .ZN(n1985) );
NOR2_X1 U1568 ( .A1(n1989), .A2(n1990), .ZN(n1988) );
NOR2_X1 U1569 ( .A1(KEYINPUT27), .A2(n1991), .ZN(n1989) );
NOR2_X1 U1570 ( .A1(KEYINPUT27), .A2(n1992), .ZN(n1987) );
INV_X1 U1571 ( .A(n1990), .ZN(n1992) );
NOR3_X1 U1572 ( .A1(n1993), .A2(n1994), .A3(n1995), .ZN(n1984) );
XNOR2_X1 U1573 ( .A(n1996), .B(KEYINPUT55), .ZN(n1995) );
XOR2_X1 U1574 ( .A(n1997), .B(KEYINPUT38), .Z(n1994) );
NOR2_X1 U1575 ( .A1(n1998), .A2(n1999), .ZN(n1983) );
XNOR2_X1 U1576 ( .A(n1978), .B(KEYINPUT20), .ZN(n1998) );
AND2_X1 U1577 ( .A1(n2000), .A2(n2001), .ZN(n1974) );
NAND3_X1 U1578 ( .A1(n2002), .A2(n1997), .A3(n1996), .ZN(n2001) );
NAND3_X1 U1579 ( .A1(n1991), .A2(n1990), .A3(n2003), .ZN(n2000) );
NAND2_X1 U1580 ( .A1(n2004), .A2(n2005), .ZN(n1990) );
NAND2_X1 U1581 ( .A1(n1979), .A2(RLAST_REG_6__SCAN_IN), .ZN(n1981) );
NAND2_X1 U1582 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1759), .ZN(n1980) );
NAND4_X1 U1583 ( .A1(n2006), .A2(n2007), .A3(n2008), .A4(n2009), .ZN(U286));
NOR3_X1 U1584 ( .A1(n2010), .A2(n2011), .A3(n2012), .ZN(n2009) );
NOR2_X1 U1585 ( .A1(n2013), .A2(n2014), .ZN(n2012) );
NOR2_X1 U1586 ( .A1(n2015), .A2(n2016), .ZN(n2011) );
AND2_X1 U1587 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1979), .ZN(n2010) );
NAND2_X1 U1588 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n2017), .ZN(n2008) );
XNOR2_X1 U1589 ( .A(KEYINPUT57), .B(U280), .ZN(n2017) );
NAND3_X1 U1590 ( .A1(n2002), .A2(n1997), .A3(n2018), .ZN(n2007) );
XOR2_X1 U1591 ( .A(n2019), .B(KEYINPUT42), .Z(n2018) );
OR2_X1 U1592 ( .A1(n2020), .A2(n2021), .ZN(n2019) );
NAND2_X1 U1593 ( .A1(n2021), .A2(n2020), .ZN(n1997) );
NAND2_X1 U1594 ( .A1(n2022), .A2(n2023), .ZN(n2020) );
NAND2_X1 U1595 ( .A1(n2024), .A2(n2025), .ZN(n2023) );
NAND2_X1 U1596 ( .A1(n2026), .A2(n2027), .ZN(n2025) );
INV_X1 U1597 ( .A(n1996), .ZN(n2022) );
NOR3_X1 U1598 ( .A1(n2028), .A2(n2024), .A3(n2029), .ZN(n1996) );
INV_X1 U1599 ( .A(n1993), .ZN(n2002) );
NAND2_X1 U1600 ( .A1(n2030), .A2(n2003), .ZN(n2006) );
XOR2_X1 U1601 ( .A(n2005), .B(n2004), .Z(n2030) );
NAND2_X1 U1602 ( .A1(n2031), .A2(n2032), .ZN(n2005) );
NAND2_X1 U1603 ( .A1(n2024), .A2(n2033), .ZN(n2032) );
INV_X1 U1604 ( .A(n1991), .ZN(n2031) );
NOR2_X1 U1605 ( .A1(n2033), .A2(n2024), .ZN(n1991) );
INV_X1 U1606 ( .A(n2015), .ZN(n2024) );
NAND2_X1 U1607 ( .A1(n2034), .A2(n2035), .ZN(n2015) );
NAND4_X1 U1608 ( .A1(n2036), .A2(n2037), .A3(n2038), .A4(n2039), .ZN(n2035));
NAND2_X1 U1609 ( .A1(n2040), .A2(n2041), .ZN(n2037) );
XNOR2_X1 U1610 ( .A(KEYINPUT19), .B(n2042), .ZN(n2040) );
NAND2_X1 U1611 ( .A1(n2043), .A2(n2044), .ZN(n2036) );
NAND2_X1 U1612 ( .A1(n2045), .A2(n2046), .ZN(n2044) );
NAND3_X1 U1613 ( .A1(n2047), .A2(n2048), .A3(n2049), .ZN(n2034) );
NOR3_X1 U1614 ( .A1(n2050), .A2(n2051), .A3(n2052), .ZN(n2049) );
NOR3_X1 U1615 ( .A1(n2053), .A2(n2041), .A3(n2054), .ZN(n2052) );
INV_X1 U1616 ( .A(KEYINPUT56), .ZN(n2053) );
NOR2_X1 U1617 ( .A1(KEYINPUT56), .A2(n2055), .ZN(n2051) );
NOR2_X1 U1618 ( .A1(n2056), .A2(n2057), .ZN(n2050) );
NAND2_X1 U1619 ( .A1(n2058), .A2(n2059), .ZN(n2048) );
XOR2_X1 U1620 ( .A(n2038), .B(KEYINPUT59), .Z(n2058) );
NAND2_X1 U1621 ( .A1(n2056), .A2(n2057), .ZN(n2038) );
NAND2_X1 U1622 ( .A1(n2042), .A2(n2039), .ZN(n2047) );
NAND2_X1 U1623 ( .A1(n2055), .A2(n2054), .ZN(n2039) );
XOR2_X1 U1624 ( .A(n2042), .B(KEYINPUT50), .Z(n2054) );
INV_X1 U1625 ( .A(n2041), .ZN(n2055) );
NAND2_X1 U1626 ( .A1(n2060), .A2(n2061), .ZN(n2041) );
NAND2_X1 U1627 ( .A1(n2062), .A2(n2063), .ZN(n2061) );
NAND2_X1 U1628 ( .A1(REG4_REG_6__SCAN_IN), .A2(n2064), .ZN(n2062) );
NAND2_X1 U1629 ( .A1(n2065), .A2(n1848), .ZN(n2060) );
INV_X1 U1630 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1848) );
NAND2_X1 U1631 ( .A1(REG4_REG_6__SCAN_IN), .A2(n2066), .ZN(n2065) );
NAND2_X1 U1632 ( .A1(RESTART), .A2(n2064), .ZN(n2066) );
INV_X1 U1633 ( .A(KEYINPUT25), .ZN(n2064) );
NAND2_X1 U1634 ( .A1(n2067), .A2(n2068), .ZN(n2042) );
NAND2_X1 U1635 ( .A1(RESTART), .A2(n1857), .ZN(n2068) );
NAND2_X1 U1636 ( .A1(n1846), .A2(n2063), .ZN(n2067) );
INV_X1 U1637 ( .A(DATA_IN_6_), .ZN(n1846) );
NAND4_X1 U1638 ( .A1(n2069), .A2(n2070), .A3(n2071), .A4(n2072), .ZN(U285));
NOR3_X1 U1639 ( .A1(n2073), .A2(n2074), .A3(n2075), .ZN(n2072) );
NOR3_X1 U1640 ( .A1(n1993), .A2(n2021), .A3(n2076), .ZN(n2075) );
XOR2_X1 U1641 ( .A(n2077), .B(KEYINPUT13), .Z(n2076) );
NAND2_X1 U1642 ( .A1(n2078), .A2(n2079), .ZN(n2077) );
XOR2_X1 U1643 ( .A(n2080), .B(KEYINPUT47), .Z(n2078) );
NAND2_X1 U1644 ( .A1(n2081), .A2(n2082), .ZN(n2080) );
AND3_X1 U1645 ( .A1(n2081), .A2(n2082), .A3(n2083), .ZN(n2021) );
XOR2_X1 U1646 ( .A(n2079), .B(KEYINPUT34), .Z(n2083) );
XNOR2_X1 U1647 ( .A(n2026), .B(n2028), .ZN(n2079) );
INV_X1 U1648 ( .A(n2029), .ZN(n2026) );
NOR3_X1 U1649 ( .A1(n1986), .A2(n2004), .A3(n2084), .ZN(n2074) );
NOR3_X1 U1650 ( .A1(n2028), .A2(n2085), .A3(n2086), .ZN(n2084) );
INV_X1 U1651 ( .A(n2033), .ZN(n2086) );
AND2_X1 U1652 ( .A1(n2085), .A2(n2087), .ZN(n2004) );
NAND2_X1 U1653 ( .A1(n2033), .A2(n2088), .ZN(n2087) );
NAND2_X1 U1654 ( .A1(n2028), .A2(n2029), .ZN(n2088) );
NAND2_X1 U1655 ( .A1(n2027), .A2(n2089), .ZN(n2033) );
XNOR2_X1 U1656 ( .A(KEYINPUT21), .B(n2029), .ZN(n2089) );
NOR2_X1 U1657 ( .A1(n2027), .A2(n2016), .ZN(n2073) );
INV_X1 U1658 ( .A(n2028), .ZN(n2027) );
XOR2_X1 U1659 ( .A(n2057), .B(n2090), .Z(n2028) );
NOR2_X1 U1660 ( .A1(n2091), .A2(n2092), .ZN(n2090) );
NOR3_X1 U1661 ( .A1(n2059), .A2(KEYINPUT30), .A3(n2046), .ZN(n2092) );
NOR2_X1 U1662 ( .A1(n2043), .A2(n2056), .ZN(n2091) );
INV_X1 U1663 ( .A(n2046), .ZN(n2056) );
NAND2_X1 U1664 ( .A1(n2093), .A2(n2094), .ZN(n2046) );
OR2_X1 U1665 ( .A1(n2063), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2094) );
NAND2_X1 U1666 ( .A1(n1845), .A2(n2063), .ZN(n2093) );
INV_X1 U1667 ( .A(n2059), .ZN(n2043) );
NAND2_X1 U1668 ( .A1(n2095), .A2(n2096), .ZN(n2059) );
NAND2_X1 U1669 ( .A1(n2097), .A2(n2098), .ZN(n2096) );
OR2_X1 U1670 ( .A1(n2099), .A2(n2100), .ZN(n2097) );
NAND2_X1 U1671 ( .A1(n2099), .A2(n2100), .ZN(n2095) );
INV_X1 U1672 ( .A(n2045), .ZN(n2057) );
NAND2_X1 U1673 ( .A1(n2101), .A2(n2102), .ZN(n2045) );
NAND2_X1 U1674 ( .A1(RESTART), .A2(n1824), .ZN(n2102) );
NAND2_X1 U1675 ( .A1(n2013), .A2(n2063), .ZN(n2101) );
NAND2_X1 U1676 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1759), .ZN(n2071) );
NAND2_X1 U1677 ( .A1(n1978), .A2(REG4_REG_4__SCAN_IN), .ZN(n2070) );
NAND2_X1 U1678 ( .A1(n1979), .A2(RLAST_REG_4__SCAN_IN), .ZN(n2069) );
NAND4_X1 U1679 ( .A1(n2103), .A2(n2104), .A3(n2105), .A4(n2106), .ZN(U284));
NOR3_X1 U1680 ( .A1(n2107), .A2(n2108), .A3(n2109), .ZN(n2106) );
NOR2_X1 U1681 ( .A1(n2110), .A2(n1993), .ZN(n2109) );
XOR2_X1 U1682 ( .A(n2082), .B(n2111), .Z(n2110) );
NOR2_X1 U1683 ( .A1(n2081), .A2(KEYINPUT17), .ZN(n2111) );
NOR3_X1 U1684 ( .A1(n1986), .A2(n2085), .A3(n2112), .ZN(n2108) );
NOR2_X1 U1685 ( .A1(n2113), .A2(n2082), .ZN(n2112) );
AND2_X1 U1686 ( .A1(n2113), .A2(n2082), .ZN(n2085) );
NAND2_X1 U1687 ( .A1(n2029), .A2(n2114), .ZN(n2082) );
NAND2_X1 U1688 ( .A1(n2115), .A2(n2116), .ZN(n2114) );
NAND2_X1 U1689 ( .A1(n2117), .A2(n2118), .ZN(n2116) );
NAND3_X1 U1690 ( .A1(n2119), .A2(n2118), .A3(n2117), .ZN(n2029) );
NOR2_X1 U1691 ( .A1(n2119), .A2(n2016), .ZN(n2107) );
INV_X1 U1692 ( .A(n2115), .ZN(n2119) );
XOR2_X1 U1693 ( .A(n2120), .B(n2099), .Z(n2115) );
NAND2_X1 U1694 ( .A1(n2121), .A2(n2122), .ZN(n2099) );
NAND2_X1 U1695 ( .A1(RESTART), .A2(n1844), .ZN(n2122) );
OR2_X1 U1696 ( .A1(REG4_REG_4__SCAN_IN), .A2(RESTART), .ZN(n2121) );
XNOR2_X1 U1697 ( .A(n2098), .B(n2100), .ZN(n2120) );
NAND2_X1 U1698 ( .A1(n2123), .A2(n2124), .ZN(n2100) );
NAND2_X1 U1699 ( .A1(n2125), .A2(n2063), .ZN(n2124) );
NAND2_X1 U1700 ( .A1(DATA_IN_4_), .A2(n2126), .ZN(n2125) );
NAND2_X1 U1701 ( .A1(n2127), .A2(n1864), .ZN(n2123) );
NAND2_X1 U1702 ( .A1(DATA_IN_4_), .A2(n2128), .ZN(n2127) );
NAND2_X1 U1703 ( .A1(RESTART), .A2(n2126), .ZN(n2128) );
INV_X1 U1704 ( .A(KEYINPUT22), .ZN(n2126) );
NAND2_X1 U1705 ( .A1(n2129), .A2(n2130), .ZN(n2098) );
NAND2_X1 U1706 ( .A1(n2131), .A2(n2132), .ZN(n2130) );
OR2_X1 U1707 ( .A1(n2133), .A2(n2134), .ZN(n2132) );
NAND2_X1 U1708 ( .A1(n2134), .A2(n2133), .ZN(n2129) );
NAND2_X1 U1709 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1759), .ZN(n2105) );
NAND2_X1 U1710 ( .A1(n1978), .A2(REG4_REG_3__SCAN_IN), .ZN(n2104) );
NAND2_X1 U1711 ( .A1(n1979), .A2(RLAST_REG_3__SCAN_IN), .ZN(n2103) );
NAND4_X1 U1712 ( .A1(n2135), .A2(n2136), .A3(n2137), .A4(n2138), .ZN(U283));
NOR3_X1 U1713 ( .A1(n2139), .A2(n2140), .A3(n2141), .ZN(n2138) );
NOR3_X1 U1714 ( .A1(n1993), .A2(n2081), .A3(n2142), .ZN(n2141) );
NOR2_X1 U1715 ( .A1(n2143), .A2(n2144), .ZN(n2142) );
AND2_X1 U1716 ( .A1(n2145), .A2(n2146), .ZN(n2143) );
AND3_X1 U1717 ( .A1(n2146), .A2(n2145), .A3(n2144), .ZN(n2081) );
NOR3_X1 U1718 ( .A1(n1986), .A2(n2113), .A3(n2147), .ZN(n2140) );
NOR2_X1 U1719 ( .A1(n2148), .A2(n2144), .ZN(n2147) );
AND2_X1 U1720 ( .A1(n2148), .A2(n2144), .ZN(n2113) );
XNOR2_X1 U1721 ( .A(n2118), .B(n2117), .ZN(n2144) );
INV_X1 U1722 ( .A(n2149), .ZN(n2148) );
NOR2_X1 U1723 ( .A1(n2118), .A2(n2016), .ZN(n2139) );
XOR2_X1 U1724 ( .A(n2131), .B(n2150), .Z(n2118) );
XOR2_X1 U1725 ( .A(n2133), .B(n2151), .Z(n2150) );
NAND2_X1 U1726 ( .A1(KEYINPUT33), .A2(n2152), .ZN(n2151) );
INV_X1 U1727 ( .A(n2134), .ZN(n2152) );
NAND2_X1 U1728 ( .A1(n2153), .A2(n2154), .ZN(n2134) );
NAND2_X1 U1729 ( .A1(RESTART), .A2(n2155), .ZN(n2154) );
NAND2_X1 U1730 ( .A1(n2156), .A2(n2063), .ZN(n2153) );
NAND2_X1 U1731 ( .A1(n2157), .A2(n2158), .ZN(n2133) );
NAND2_X1 U1732 ( .A1(n2159), .A2(n2160), .ZN(n2158) );
NAND2_X1 U1733 ( .A1(n2161), .A2(n2162), .ZN(n2160) );
XNOR2_X1 U1734 ( .A(KEYINPUT41), .B(n2163), .ZN(n2159) );
NAND2_X1 U1735 ( .A1(n2164), .A2(n2165), .ZN(n2157) );
NAND2_X1 U1736 ( .A1(n2166), .A2(n2167), .ZN(n2131) );
NAND2_X1 U1737 ( .A1(RESTART), .A2(n1878), .ZN(n2167) );
NAND2_X1 U1738 ( .A1(n1843), .A2(n2063), .ZN(n2166) );
NAND2_X1 U1739 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1759), .ZN(n2137) );
NAND2_X1 U1740 ( .A1(n1978), .A2(REG4_REG_2__SCAN_IN), .ZN(n2136) );
NAND2_X1 U1741 ( .A1(n1979), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2135) );
NAND4_X1 U1742 ( .A1(n2168), .A2(n2169), .A3(n2170), .A4(n2171), .ZN(U282));
NOR3_X1 U1743 ( .A1(n2172), .A2(n2173), .A3(n2174), .ZN(n2171) );
NOR2_X1 U1744 ( .A1(n2175), .A2(n1993), .ZN(n2174) );
XNOR2_X1 U1745 ( .A(n2145), .B(n2146), .ZN(n2175) );
NAND2_X1 U1746 ( .A1(n2176), .A2(n2177), .ZN(n2146) );
NAND2_X1 U1747 ( .A1(n2178), .A2(n2179), .ZN(n2177) );
XNOR2_X1 U1748 ( .A(n2180), .B(KEYINPUT15), .ZN(n2178) );
NOR3_X1 U1749 ( .A1(n1986), .A2(n2181), .A3(n2182), .ZN(n2173) );
NOR2_X1 U1750 ( .A1(n2183), .A2(n2149), .ZN(n2182) );
NAND2_X1 U1751 ( .A1(n2184), .A2(n2185), .ZN(n2149) );
NOR2_X1 U1752 ( .A1(KEYINPUT31), .A2(KEYINPUT12), .ZN(n2183) );
NOR2_X1 U1753 ( .A1(n2186), .A2(n2185), .ZN(n2181) );
NOR2_X1 U1754 ( .A1(n2187), .A2(n2188), .ZN(n2186) );
XNOR2_X1 U1755 ( .A(KEYINPUT31), .B(n2184), .ZN(n2188) );
NAND2_X1 U1756 ( .A1(n2176), .A2(n2189), .ZN(n2184) );
NAND2_X1 U1757 ( .A1(n2190), .A2(n2179), .ZN(n2189) );
NOR2_X1 U1758 ( .A1(n2117), .A2(n2191), .ZN(n2176) );
AND2_X1 U1759 ( .A1(n2192), .A2(n2179), .ZN(n2191) );
NOR2_X1 U1760 ( .A1(n2193), .A2(n2179), .ZN(n2117) );
INV_X1 U1761 ( .A(KEYINPUT12), .ZN(n2187) );
NOR2_X1 U1762 ( .A1(n2194), .A2(n2016), .ZN(n2172) );
INV_X1 U1763 ( .A(n2179), .ZN(n2194) );
NAND3_X1 U1764 ( .A1(n2195), .A2(n2196), .A3(n2197), .ZN(n2179) );
OR2_X1 U1765 ( .A1(n2198), .A2(KEYINPUT5), .ZN(n2197) );
NAND2_X1 U1766 ( .A1(n2161), .A2(n2199), .ZN(n2196) );
NAND2_X1 U1767 ( .A1(n2200), .A2(n2201), .ZN(n2199) );
OR2_X1 U1768 ( .A1(n2198), .A2(KEYINPUT62), .ZN(n2201) );
XNOR2_X1 U1769 ( .A(n2202), .B(n2162), .ZN(n2200) );
NAND2_X1 U1770 ( .A1(KEYINPUT5), .A2(n2198), .ZN(n2202) );
INV_X1 U1771 ( .A(n2165), .ZN(n2161) );
NAND2_X1 U1772 ( .A1(n2203), .A2(n2165), .ZN(n2195) );
NAND2_X1 U1773 ( .A1(n2204), .A2(n2205), .ZN(n2165) );
NAND2_X1 U1774 ( .A1(n2206), .A2(n2063), .ZN(n2205) );
NAND2_X1 U1775 ( .A1(REG4_REG_2__SCAN_IN), .A2(n2207), .ZN(n2206) );
NAND2_X1 U1776 ( .A1(n2208), .A2(n2209), .ZN(n2204) );
NAND2_X1 U1777 ( .A1(REG4_REG_2__SCAN_IN), .A2(n2210), .ZN(n2208) );
NAND2_X1 U1778 ( .A1(RESTART), .A2(n2207), .ZN(n2210) );
INV_X1 U1779 ( .A(KEYINPUT2), .ZN(n2207) );
NAND2_X1 U1780 ( .A1(n2211), .A2(n2212), .ZN(n2203) );
NAND2_X1 U1781 ( .A1(n2162), .A2(n2213), .ZN(n2212) );
NAND2_X1 U1782 ( .A1(KEYINPUT5), .A2(n2214), .ZN(n2213) );
NAND2_X1 U1783 ( .A1(KEYINPUT62), .A2(n2163), .ZN(n2214) );
INV_X1 U1784 ( .A(n2164), .ZN(n2162) );
NAND3_X1 U1785 ( .A1(KEYINPUT5), .A2(n2198), .A3(n2164), .ZN(n2211) );
NAND2_X1 U1786 ( .A1(n2215), .A2(n2216), .ZN(n2164) );
NAND2_X1 U1787 ( .A1(RESTART), .A2(n1873), .ZN(n2216) );
NAND2_X1 U1788 ( .A1(n1836), .A2(n2063), .ZN(n2215) );
INV_X1 U1789 ( .A(DATA_IN_2_), .ZN(n1836) );
INV_X1 U1790 ( .A(n2163), .ZN(n2198) );
NAND2_X1 U1791 ( .A1(n2217), .A2(n2218), .ZN(n2163) );
NAND2_X1 U1792 ( .A1(n2219), .A2(n2220), .ZN(n2218) );
INV_X1 U1793 ( .A(n2221), .ZN(n2220) );
XNOR2_X1 U1794 ( .A(KEYINPUT44), .B(n2222), .ZN(n2219) );
NAND2_X1 U1795 ( .A1(n2223), .A2(n2224), .ZN(n2217) );
NAND2_X1 U1796 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1759), .ZN(n2170) );
NAND2_X1 U1797 ( .A1(n1978), .A2(REG4_REG_1__SCAN_IN), .ZN(n2169) );
INV_X1 U1798 ( .A(n2014), .ZN(n1978) );
NAND2_X1 U1799 ( .A1(n1979), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2168) );
NAND4_X1 U1800 ( .A1(n2225), .A2(n2226), .A3(n2227), .A4(n2228), .ZN(U281));
NOR3_X1 U1801 ( .A1(n2229), .A2(n2230), .A3(n2231), .ZN(n2228) );
NOR2_X1 U1802 ( .A1(n2232), .A2(n2014), .ZN(n2231) );
NAND2_X1 U1803 ( .A1(AVERAGE), .A2(n2233), .ZN(n2014) );
NOR2_X1 U1804 ( .A1(n1986), .A2(n2185), .ZN(n2230) );
NAND2_X1 U1805 ( .A1(n2193), .A2(n2234), .ZN(n2185) );
NAND2_X1 U1806 ( .A1(n2192), .A2(n2190), .ZN(n2234) );
INV_X1 U1807 ( .A(n2003), .ZN(n1986) );
NOR2_X1 U1808 ( .A1(n2235), .A2(n2236), .ZN(n2003) );
NOR2_X1 U1809 ( .A1(n1993), .A2(n2145), .ZN(n2229) );
NAND3_X1 U1810 ( .A1(n2237), .A2(n2238), .A3(n2193), .ZN(n2145) );
OR2_X1 U1811 ( .A1(n2190), .A2(n2192), .ZN(n2193) );
OR2_X1 U1812 ( .A1(n2190), .A2(KEYINPUT37), .ZN(n2238) );
NAND3_X1 U1813 ( .A1(n2192), .A2(n2190), .A3(KEYINPUT37), .ZN(n2237) );
NAND3_X1 U1814 ( .A1(n2239), .A2(n2240), .A3(n2241), .ZN(n2192) );
NAND2_X1 U1815 ( .A1(n2242), .A2(n2243), .ZN(n2241) );
NAND2_X1 U1816 ( .A1(n2244), .A2(n2245), .ZN(n2240) );
INV_X1 U1817 ( .A(KEYINPUT32), .ZN(n2245) );
NAND2_X1 U1818 ( .A1(n2246), .A2(n2247), .ZN(n2244) );
XNOR2_X1 U1819 ( .A(n2243), .B(n2248), .ZN(n2246) );
NAND2_X1 U1820 ( .A1(KEYINPUT32), .A2(n2249), .ZN(n2239) );
NAND2_X1 U1821 ( .A1(n2250), .A2(n2251), .ZN(n2249) );
NAND2_X1 U1822 ( .A1(n2243), .A2(n2248), .ZN(n2251) );
OR3_X1 U1823 ( .A1(n2242), .A2(n2243), .A3(n2248), .ZN(n2250) );
INV_X1 U1824 ( .A(KEYINPUT39), .ZN(n2248) );
INV_X1 U1825 ( .A(n2247), .ZN(n2242) );
NAND4_X1 U1826 ( .A1(n2233), .A2(n2252), .A3(n2253), .A4(n2254), .ZN(n1993));
NAND2_X1 U1827 ( .A1(n2255), .A2(n2256), .ZN(n2253) );
INV_X1 U1828 ( .A(REG4_REG_7__SCAN_IN), .ZN(n2256) );
NOR3_X1 U1829 ( .A1(n2236), .A2(RESTART), .A3(n1905), .ZN(n2233) );
INV_X1 U1830 ( .A(ENABLE), .ZN(n1905) );
XOR2_X1 U1831 ( .A(n2257), .B(KEYINPUT4), .Z(n2227) );
NAND2_X1 U1832 ( .A1(n1979), .A2(RLAST_REG_0__SCAN_IN), .ZN(n2257) );
NOR3_X1 U1833 ( .A1(ENABLE), .A2(RESTART), .A3(n2236), .ZN(n1979) );
NAND2_X1 U1834 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1759), .ZN(n2226) );
XOR2_X1 U1835 ( .A(KEYINPUT7), .B(n2258), .Z(n2225) );
NOR2_X1 U1836 ( .A1(n2180), .A2(n2016), .ZN(n2258) );
NAND3_X1 U1837 ( .A1(n2259), .A2(n2235), .A3(n2260), .ZN(n2016) );
INV_X1 U1838 ( .A(n2236), .ZN(n2260) );
NAND2_X1 U1839 ( .A1(STATO_REG_1__SCAN_IN), .A2(U280), .ZN(n2236) );
NAND3_X1 U1840 ( .A1(n2261), .A2(n2262), .A3(RESTART), .ZN(n2235) );
NAND2_X1 U1841 ( .A1(n2263), .A2(n1849), .ZN(n2262) );
INV_X1 U1842 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1849) );
OR2_X1 U1843 ( .A1(n2264), .A2(n1853), .ZN(n2263) );
NAND2_X1 U1844 ( .A1(n2264), .A2(n1853), .ZN(n2261) );
INV_X1 U1845 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1853) );
NAND2_X1 U1846 ( .A1(n2265), .A2(n2266), .ZN(n2264) );
NAND2_X1 U1847 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n2267), .ZN(n2266) );
NAND2_X1 U1848 ( .A1(n2268), .A2(n1857), .ZN(n2267) );
INV_X1 U1849 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1857) );
XOR2_X1 U1850 ( .A(KEYINPUT26), .B(n2269), .Z(n2268) );
NAND2_X1 U1851 ( .A1(n2269), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2265) );
AND2_X1 U1852 ( .A1(n2270), .A2(n2271), .ZN(n2269) );
NAND2_X1 U1853 ( .A1(n1824), .A2(n2272), .ZN(n2271) );
NAND2_X1 U1854 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n2273), .ZN(n2272) );
INV_X1 U1855 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1824) );
OR2_X1 U1856 ( .A1(n2273), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2270) );
NAND2_X1 U1857 ( .A1(n2274), .A2(n2275), .ZN(n2273) );
NAND2_X1 U1858 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2275) );
NAND3_X1 U1859 ( .A1(n2276), .A2(n2277), .A3(n2278), .ZN(n2274) );
NAND2_X1 U1860 ( .A1(n1864), .A2(n1844), .ZN(n2278) );
INV_X1 U1861 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1844) );
INV_X1 U1862 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1864) );
NAND3_X1 U1863 ( .A1(n2279), .A2(n2280), .A3(n2281), .ZN(n2277) );
NAND2_X1 U1864 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2281) );
NAND3_X1 U1865 ( .A1(n2282), .A2(n2283), .A3(n2284), .ZN(n2280) );
NAND2_X1 U1866 ( .A1(n1873), .A2(n2209), .ZN(n2284) );
INV_X1 U1867 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n2209) );
INV_X1 U1868 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1873) );
NAND2_X1 U1869 ( .A1(n2285), .A2(n2286), .ZN(n2283) );
NAND2_X1 U1870 ( .A1(RMIN_REG_1__SCAN_IN), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2286) );
NAND2_X1 U1871 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2285) );
NAND2_X1 U1872 ( .A1(n2287), .A2(n1839), .ZN(n2282) );
NAND2_X1 U1873 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2279) );
NAND2_X1 U1874 ( .A1(n1878), .A2(n2155), .ZN(n2276) );
INV_X1 U1875 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n2155) );
INV_X1 U1876 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1878) );
NAND2_X1 U1877 ( .A1(n2288), .A2(n2063), .ZN(n2259) );
XOR2_X1 U1878 ( .A(n2289), .B(KEYINPUT54), .Z(n2288) );
NAND4_X1 U1879 ( .A1(ENABLE), .A2(n2255), .A3(n2290), .A4(n2254), .ZN(n2289));
INV_X1 U1880 ( .A(AVERAGE), .ZN(n2254) );
NAND2_X1 U1881 ( .A1(REG4_REG_7__SCAN_IN), .A2(n2252), .ZN(n2290) );
NAND2_X1 U1882 ( .A1(n2291), .A2(n1816), .ZN(n2252) );
INV_X1 U1883 ( .A(DATA_IN_7_), .ZN(n1816) );
INV_X1 U1884 ( .A(n2292), .ZN(n2291) );
NAND2_X1 U1885 ( .A1(DATA_IN_7_), .A2(n2292), .ZN(n2255) );
NAND2_X1 U1886 ( .A1(n2293), .A2(n2294), .ZN(n2292) );
NAND2_X1 U1887 ( .A1(n2295), .A2(n1999), .ZN(n2294) );
INV_X1 U1888 ( .A(REG4_REG_6__SCAN_IN), .ZN(n1999) );
XOR2_X1 U1889 ( .A(n2296), .B(KEYINPUT49), .Z(n2295) );
NAND2_X1 U1890 ( .A1(n2297), .A2(DATA_IN_6_), .ZN(n2296) );
XOR2_X1 U1891 ( .A(n2298), .B(KEYINPUT0), .Z(n2297) );
OR2_X1 U1892 ( .A1(n2298), .A2(DATA_IN_6_), .ZN(n2293) );
NAND2_X1 U1893 ( .A1(n2299), .A2(n2300), .ZN(n2298) );
NAND2_X1 U1894 ( .A1(n2301), .A2(n2302), .ZN(n2300) );
NAND2_X1 U1895 ( .A1(n2013), .A2(n1845), .ZN(n2302) );
INV_X1 U1896 ( .A(DATA_IN_5_), .ZN(n1845) );
INV_X1 U1897 ( .A(REG4_REG_5__SCAN_IN), .ZN(n2013) );
NAND2_X1 U1898 ( .A1(n2303), .A2(n2304), .ZN(n2301) );
NAND2_X1 U1899 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2304) );
NAND3_X1 U1900 ( .A1(n2305), .A2(n2306), .A3(n2307), .ZN(n2303) );
XOR2_X1 U1901 ( .A(KEYINPUT35), .B(n2308), .Z(n2307) );
NOR2_X1 U1902 ( .A1(DATA_IN_4_), .A2(REG4_REG_4__SCAN_IN), .ZN(n2308) );
NAND3_X1 U1903 ( .A1(n2309), .A2(n2310), .A3(n2311), .ZN(n2306) );
NAND2_X1 U1904 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2311) );
NAND3_X1 U1905 ( .A1(n2312), .A2(n2313), .A3(n2314), .ZN(n2310) );
OR2_X1 U1906 ( .A1(DATA_IN_2_), .A2(REG4_REG_2__SCAN_IN), .ZN(n2314) );
NAND2_X1 U1907 ( .A1(n2315), .A2(n2316), .ZN(n2313) );
NAND2_X1 U1908 ( .A1(REG4_REG_1__SCAN_IN), .A2(DATA_IN_1_), .ZN(n2316) );
NAND2_X1 U1909 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2315) );
NAND2_X1 U1910 ( .A1(n1840), .A2(n2317), .ZN(n2312) );
NAND2_X1 U1911 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2309) );
NAND2_X1 U1912 ( .A1(n1843), .A2(n2156), .ZN(n2305) );
INV_X1 U1913 ( .A(REG4_REG_3__SCAN_IN), .ZN(n2156) );
INV_X1 U1914 ( .A(DATA_IN_3_), .ZN(n1843) );
NAND2_X1 U1915 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2299) );
INV_X1 U1916 ( .A(n2190), .ZN(n2180) );
NAND3_X1 U1917 ( .A1(n2318), .A2(n2319), .A3(n2320), .ZN(n2190) );
NAND2_X1 U1918 ( .A1(n2221), .A2(n2222), .ZN(n2320) );
NOR2_X1 U1919 ( .A1(n2223), .A2(n2224), .ZN(n2221) );
OR3_X1 U1920 ( .A1(n2222), .A2(n2321), .A3(n2223), .ZN(n2319) );
NAND2_X1 U1921 ( .A1(n2322), .A2(n2223), .ZN(n2318) );
NAND3_X1 U1922 ( .A1(n2323), .A2(n2324), .A3(n2325), .ZN(n2223) );
NAND2_X1 U1923 ( .A1(n2326), .A2(n2287), .ZN(n2325) );
INV_X1 U1924 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n2287) );
NAND2_X1 U1925 ( .A1(DATA_IN_1_), .A2(n2063), .ZN(n2326) );
OR2_X1 U1926 ( .A1(n2063), .A2(KEYINPUT52), .ZN(n2324) );
NAND3_X1 U1927 ( .A1(n1840), .A2(n2063), .A3(KEYINPUT52), .ZN(n2323) );
INV_X1 U1928 ( .A(DATA_IN_1_), .ZN(n1840) );
NAND2_X1 U1929 ( .A1(n2327), .A2(n2328), .ZN(n2322) );
NAND2_X1 U1930 ( .A1(n2222), .A2(n2224), .ZN(n2328) );
INV_X1 U1931 ( .A(n2321), .ZN(n2224) );
XOR2_X1 U1932 ( .A(KEYINPUT3), .B(n2329), .Z(n2327) );
NOR2_X1 U1933 ( .A1(n2330), .A2(n2222), .ZN(n2329) );
NAND3_X1 U1934 ( .A1(n2331), .A2(n2332), .A3(n2333), .ZN(n2222) );
NAND2_X1 U1935 ( .A1(KEYINPUT28), .A2(n2317), .ZN(n2333) );
INV_X1 U1936 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2317) );
NAND3_X1 U1937 ( .A1(REG4_REG_1__SCAN_IN), .A2(n2334), .A3(n2063), .ZN(n2332) );
NAND2_X1 U1938 ( .A1(RESTART), .A2(n2335), .ZN(n2331) );
NAND2_X1 U1939 ( .A1(n1839), .A2(n2334), .ZN(n2335) );
INV_X1 U1940 ( .A(KEYINPUT28), .ZN(n2334) );
INV_X1 U1941 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1839) );
XNOR2_X1 U1942 ( .A(n2321), .B(KEYINPUT29), .ZN(n2330) );
NOR2_X1 U1943 ( .A1(n2243), .A2(n2247), .ZN(n2321) );
NAND2_X1 U1944 ( .A1(n2336), .A2(n2337), .ZN(n2247) );
NAND2_X1 U1945 ( .A1(RESTART), .A2(n1875), .ZN(n2337) );
INV_X1 U1946 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1875) );
NAND2_X1 U1947 ( .A1(n1838), .A2(n2063), .ZN(n2336) );
INV_X1 U1948 ( .A(DATA_IN_0_), .ZN(n1838) );
NAND2_X1 U1949 ( .A1(n2338), .A2(n2339), .ZN(n2243) );
OR2_X1 U1950 ( .A1(n2063), .A2(RMIN_REG_0__SCAN_IN), .ZN(n2339) );
NAND2_X1 U1951 ( .A1(n2232), .A2(n2063), .ZN(n2338) );
INV_X1 U1952 ( .A(RESTART), .ZN(n2063) );
INV_X1 U1953 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2232) );
NOR2_X1 U1954 ( .A1(n1783), .A2(STATO_REG_1__SCAN_IN), .ZN(n2340) );
INV_X1 U1955 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1783) );
endmodule


