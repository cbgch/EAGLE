//Key = 1001000001000111101011101010001110011000111100100110000111110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304;

XOR2_X1 U714 ( .A(G107), .B(n978), .Z(G9) );
NAND4_X1 U715 ( .A1(n979), .A2(n980), .A3(n981), .A4(n982), .ZN(G75) );
NAND2_X1 U716 ( .A1(n983), .A2(n984), .ZN(n982) );
NAND2_X1 U717 ( .A1(n985), .A2(n986), .ZN(n984) );
NAND3_X1 U718 ( .A1(n987), .A2(n988), .A3(n989), .ZN(n986) );
NAND2_X1 U719 ( .A1(n990), .A2(n991), .ZN(n987) );
NAND3_X1 U720 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
NAND2_X1 U721 ( .A1(n995), .A2(n996), .ZN(n993) );
NAND2_X1 U722 ( .A1(n997), .A2(n998), .ZN(n990) );
NAND2_X1 U723 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND2_X1 U724 ( .A1(n994), .A2(n1001), .ZN(n1000) );
NAND2_X1 U725 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NAND2_X1 U726 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
INV_X1 U727 ( .A(n1006), .ZN(n1002) );
NAND2_X1 U728 ( .A1(n992), .A2(n1007), .ZN(n999) );
NAND2_X1 U729 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND2_X1 U730 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND4_X1 U731 ( .A1(n994), .A2(n997), .A3(n992), .A4(n1012), .ZN(n985) );
NAND2_X1 U732 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
XOR2_X1 U733 ( .A(KEYINPUT59), .B(n1015), .Z(n1013) );
NOR2_X1 U734 ( .A1(n1016), .A2(n988), .ZN(n1015) );
INV_X1 U735 ( .A(n1017), .ZN(n983) );
NOR2_X1 U736 ( .A1(G953), .A2(n1018), .ZN(n981) );
NOR4_X1 U737 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
XOR2_X1 U738 ( .A(n1023), .B(n1024), .Z(n1022) );
NOR2_X1 U739 ( .A1(n1025), .A2(KEYINPUT51), .ZN(n1024) );
NOR2_X1 U740 ( .A1(n1026), .A2(n1027), .ZN(n1021) );
XNOR2_X1 U741 ( .A(KEYINPUT41), .B(n1028), .ZN(n1027) );
NAND3_X1 U742 ( .A1(n1029), .A2(n1030), .A3(n988), .ZN(n1020) );
NAND4_X1 U743 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1019) );
XOR2_X1 U744 ( .A(KEYINPUT37), .B(n1035), .Z(n1034) );
NOR3_X1 U745 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
AND3_X1 U746 ( .A1(KEYINPUT30), .A2(n1039), .A3(G475), .ZN(n1038) );
NOR2_X1 U747 ( .A1(KEYINPUT30), .A2(G475), .ZN(n1037) );
XOR2_X1 U748 ( .A(n1040), .B(G478), .Z(n1031) );
XOR2_X1 U749 ( .A(n1041), .B(n1042), .Z(G72) );
XOR2_X1 U750 ( .A(n1043), .B(n1044), .Z(n1042) );
NOR2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
XOR2_X1 U752 ( .A(KEYINPUT57), .B(G953), .Z(n1046) );
NOR2_X1 U753 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND2_X1 U754 ( .A1(n1049), .A2(n1050), .ZN(n1043) );
NAND2_X1 U755 ( .A1(G953), .A2(n1048), .ZN(n1050) );
XOR2_X1 U756 ( .A(n1051), .B(n1052), .Z(n1049) );
XOR2_X1 U757 ( .A(n1053), .B(n1054), .Z(n1051) );
NAND3_X1 U758 ( .A1(n1055), .A2(n1056), .A3(KEYINPUT56), .ZN(n1041) );
XOR2_X1 U759 ( .A(n1057), .B(n1058), .Z(G69) );
XOR2_X1 U760 ( .A(n1059), .B(n1060), .Z(n1058) );
NOR2_X1 U761 ( .A1(n1061), .A2(n1056), .ZN(n1060) );
NOR2_X1 U762 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U763 ( .A1(n1064), .A2(n1065), .ZN(n1059) );
NAND2_X1 U764 ( .A1(G953), .A2(n1063), .ZN(n1065) );
XOR2_X1 U765 ( .A(n1066), .B(n1067), .Z(n1064) );
XNOR2_X1 U766 ( .A(n1068), .B(KEYINPUT61), .ZN(n1067) );
NAND2_X1 U767 ( .A1(n1069), .A2(KEYINPUT3), .ZN(n1068) );
XOR2_X1 U768 ( .A(n1070), .B(KEYINPUT11), .Z(n1069) );
NAND2_X1 U769 ( .A1(n1056), .A2(n1071), .ZN(n1057) );
NOR3_X1 U770 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(G66) );
AND2_X1 U771 ( .A1(KEYINPUT55), .A2(n1075), .ZN(n1074) );
NOR3_X1 U772 ( .A1(KEYINPUT55), .A2(G953), .A3(G952), .ZN(n1073) );
XOR2_X1 U773 ( .A(n1076), .B(n1077), .Z(n1072) );
NOR2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U775 ( .A1(KEYINPUT45), .A2(n1080), .ZN(n1076) );
NOR2_X1 U776 ( .A1(n1081), .A2(n1082), .ZN(G63) );
XOR2_X1 U777 ( .A(KEYINPUT63), .B(n1075), .Z(n1082) );
XNOR2_X1 U778 ( .A(n1083), .B(n1084), .ZN(n1081) );
NOR2_X1 U779 ( .A1(n1085), .A2(n1079), .ZN(n1084) );
NOR2_X1 U780 ( .A1(n1075), .A2(n1086), .ZN(G60) );
XNOR2_X1 U781 ( .A(n1087), .B(n1088), .ZN(n1086) );
AND2_X1 U782 ( .A1(G475), .A2(n1089), .ZN(n1088) );
XOR2_X1 U783 ( .A(G104), .B(n1090), .Z(G6) );
NOR2_X1 U784 ( .A1(n1091), .A2(n1092), .ZN(G57) );
XNOR2_X1 U785 ( .A(n1093), .B(n1094), .ZN(n1092) );
XOR2_X1 U786 ( .A(n1095), .B(KEYINPUT27), .Z(n1093) );
NAND3_X1 U787 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
OR2_X1 U788 ( .A1(n1099), .A2(KEYINPUT49), .ZN(n1098) );
NAND3_X1 U789 ( .A1(KEYINPUT49), .A2(n1099), .A3(n1100), .ZN(n1097) );
NAND2_X1 U790 ( .A1(n1101), .A2(n1102), .ZN(n1096) );
NAND2_X1 U791 ( .A1(n1103), .A2(KEYINPUT49), .ZN(n1102) );
XNOR2_X1 U792 ( .A(n1099), .B(KEYINPUT50), .ZN(n1103) );
AND2_X1 U793 ( .A1(n1089), .A2(G472), .ZN(n1099) );
NOR2_X1 U794 ( .A1(G952), .A2(n1104), .ZN(n1091) );
XOR2_X1 U795 ( .A(KEYINPUT35), .B(G953), .Z(n1104) );
NOR2_X1 U796 ( .A1(n1075), .A2(n1105), .ZN(G54) );
XOR2_X1 U797 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U798 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U799 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U800 ( .A1(KEYINPUT23), .A2(n1112), .ZN(n1111) );
NOR2_X1 U801 ( .A1(KEYINPUT60), .A2(n1113), .ZN(n1108) );
XNOR2_X1 U802 ( .A(n1054), .B(n1114), .ZN(n1106) );
AND2_X1 U803 ( .A1(G469), .A2(n1089), .ZN(n1114) );
NOR2_X1 U804 ( .A1(n1075), .A2(n1115), .ZN(G51) );
XOR2_X1 U805 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U806 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR3_X1 U807 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
NOR2_X1 U808 ( .A1(KEYINPUT29), .A2(n1123), .ZN(n1122) );
NOR2_X1 U809 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
AND3_X1 U810 ( .A1(KEYINPUT36), .A2(n1053), .A3(n1126), .ZN(n1125) );
NOR2_X1 U811 ( .A1(KEYINPUT36), .A2(n1053), .ZN(n1124) );
NOR2_X1 U812 ( .A1(n1127), .A2(n1128), .ZN(n1121) );
INV_X1 U813 ( .A(KEYINPUT29), .ZN(n1128) );
NOR2_X1 U814 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
XOR2_X1 U815 ( .A(KEYINPUT36), .B(n1053), .Z(n1130) );
NAND3_X1 U816 ( .A1(n1089), .A2(n1025), .A3(KEYINPUT32), .ZN(n1118) );
INV_X1 U817 ( .A(n1079), .ZN(n1089) );
NAND2_X1 U818 ( .A1(G902), .A2(n1131), .ZN(n1079) );
NAND2_X1 U819 ( .A1(n979), .A2(n980), .ZN(n1131) );
INV_X1 U820 ( .A(n1055), .ZN(n980) );
NAND4_X1 U821 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1055) );
NOR4_X1 U822 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1135) );
NAND2_X1 U823 ( .A1(n994), .A2(n1140), .ZN(n1134) );
NAND2_X1 U824 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NAND2_X1 U825 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U826 ( .A(KEYINPUT25), .B(n1145), .Z(n1144) );
OR2_X1 U827 ( .A1(n1146), .A2(n1147), .ZN(n1141) );
INV_X1 U828 ( .A(n1071), .ZN(n979) );
NAND2_X1 U829 ( .A1(n1148), .A2(n1149), .ZN(n1071) );
NOR4_X1 U830 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1090), .ZN(n1149) );
AND3_X1 U831 ( .A1(n1153), .A2(n992), .A3(n1145), .ZN(n1090) );
NOR4_X1 U832 ( .A1(n978), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1148) );
INV_X1 U833 ( .A(n1157), .ZN(n1154) );
AND3_X1 U834 ( .A1(n1153), .A2(n992), .A3(n1158), .ZN(n978) );
NOR2_X1 U835 ( .A1(n1056), .A2(G952), .ZN(n1075) );
XOR2_X1 U836 ( .A(G146), .B(n1139), .Z(G48) );
NOR3_X1 U837 ( .A1(n995), .A2(n1008), .A3(n1146), .ZN(n1139) );
XNOR2_X1 U838 ( .A(n1138), .B(n1159), .ZN(G45) );
XOR2_X1 U839 ( .A(KEYINPUT9), .B(G143), .Z(n1159) );
AND4_X1 U840 ( .A1(n1143), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1138) );
INV_X1 U841 ( .A(n1163), .ZN(n1143) );
NAND2_X1 U842 ( .A1(n1164), .A2(n1165), .ZN(G42) );
NAND2_X1 U843 ( .A1(G140), .A2(n1132), .ZN(n1165) );
XOR2_X1 U844 ( .A(n1166), .B(KEYINPUT4), .Z(n1164) );
OR2_X1 U845 ( .A1(n1132), .A2(G140), .ZN(n1166) );
NAND3_X1 U846 ( .A1(n994), .A2(n1167), .A3(n1168), .ZN(n1132) );
XOR2_X1 U847 ( .A(G137), .B(n1169), .Z(G39) );
NOR4_X1 U848 ( .A1(KEYINPUT62), .A2(n1147), .A3(n1146), .A4(n1170), .ZN(n1169) );
XOR2_X1 U849 ( .A(G134), .B(n1137), .Z(G36) );
NOR3_X1 U850 ( .A1(n1163), .A2(n996), .A3(n1170), .ZN(n1137) );
XOR2_X1 U851 ( .A(G131), .B(n1171), .Z(G33) );
NOR3_X1 U852 ( .A1(n1172), .A2(n995), .A3(n1163), .ZN(n1171) );
NAND3_X1 U853 ( .A1(n1167), .A2(n1173), .A3(n1006), .ZN(n1163) );
XOR2_X1 U854 ( .A(KEYINPUT20), .B(n994), .Z(n1172) );
INV_X1 U855 ( .A(n1170), .ZN(n994) );
NAND2_X1 U856 ( .A1(n1011), .A2(n1030), .ZN(n1170) );
XOR2_X1 U857 ( .A(G128), .B(n1136), .Z(G30) );
NOR3_X1 U858 ( .A1(n996), .A2(n1008), .A3(n1146), .ZN(n1136) );
NAND4_X1 U859 ( .A1(n1167), .A2(n1174), .A3(n1173), .A4(n1005), .ZN(n1146) );
INV_X1 U860 ( .A(n1160), .ZN(n1008) );
XOR2_X1 U861 ( .A(n1152), .B(n1175), .Z(G3) );
NOR2_X1 U862 ( .A1(KEYINPUT10), .A2(n1176), .ZN(n1175) );
AND3_X1 U863 ( .A1(n1153), .A2(n1006), .A3(n997), .ZN(n1152) );
XOR2_X1 U864 ( .A(n1053), .B(n1133), .Z(G27) );
NAND4_X1 U865 ( .A1(n989), .A2(n1168), .A3(n1160), .A4(n988), .ZN(n1133) );
AND4_X1 U866 ( .A1(n1004), .A2(n1145), .A3(n1173), .A4(n1005), .ZN(n1168) );
NAND2_X1 U867 ( .A1(n1017), .A2(n1177), .ZN(n1173) );
NAND4_X1 U868 ( .A1(G953), .A2(G902), .A3(n1178), .A4(n1048), .ZN(n1177) );
INV_X1 U869 ( .A(G900), .ZN(n1048) );
NAND2_X1 U870 ( .A1(n1179), .A2(n1180), .ZN(G24) );
OR2_X1 U871 ( .A1(n1181), .A2(G122), .ZN(n1180) );
NAND2_X1 U872 ( .A1(G122), .A2(n1182), .ZN(n1179) );
NAND2_X1 U873 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NAND2_X1 U874 ( .A1(n1151), .A2(n1185), .ZN(n1184) );
INV_X1 U875 ( .A(KEYINPUT14), .ZN(n1185) );
NAND2_X1 U876 ( .A1(KEYINPUT14), .A2(n1181), .ZN(n1183) );
NAND2_X1 U877 ( .A1(KEYINPUT58), .A2(n1151), .ZN(n1181) );
AND4_X1 U878 ( .A1(n1186), .A2(n992), .A3(n1161), .A4(n1162), .ZN(n1151) );
NAND2_X1 U879 ( .A1(n1187), .A2(n1188), .ZN(n992) );
OR3_X1 U880 ( .A1(n1005), .A2(n1174), .A3(KEYINPUT52), .ZN(n1188) );
NAND2_X1 U881 ( .A1(KEYINPUT52), .A2(n1006), .ZN(n1187) );
NAND3_X1 U882 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(G21) );
OR2_X1 U883 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NAND2_X1 U884 ( .A1(n1194), .A2(n1195), .ZN(n1190) );
INV_X1 U885 ( .A(KEYINPUT42), .ZN(n1195) );
NAND2_X1 U886 ( .A1(n1196), .A2(n1193), .ZN(n1194) );
XOR2_X1 U887 ( .A(n1197), .B(n1156), .Z(n1196) );
NAND2_X1 U888 ( .A1(KEYINPUT42), .A2(n1198), .ZN(n1189) );
NAND2_X1 U889 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND3_X1 U890 ( .A1(n1197), .A2(n1193), .A3(n1192), .ZN(n1200) );
XNOR2_X1 U891 ( .A(G119), .B(KEYINPUT13), .ZN(n1193) );
NAND2_X1 U892 ( .A1(n1201), .A2(n1156), .ZN(n1199) );
INV_X1 U893 ( .A(n1192), .ZN(n1156) );
NAND4_X1 U894 ( .A1(n1186), .A2(n997), .A3(n1174), .A4(n1005), .ZN(n1192) );
INV_X1 U895 ( .A(n1032), .ZN(n1174) );
INV_X1 U896 ( .A(n1197), .ZN(n1201) );
XNOR2_X1 U897 ( .A(KEYINPUT24), .B(KEYINPUT15), .ZN(n1197) );
XOR2_X1 U898 ( .A(n1155), .B(n1202), .Z(G18) );
XOR2_X1 U899 ( .A(KEYINPUT19), .B(G116), .Z(n1202) );
AND3_X1 U900 ( .A1(n1158), .A2(n1006), .A3(n1186), .ZN(n1155) );
INV_X1 U901 ( .A(n996), .ZN(n1158) );
NAND2_X1 U902 ( .A1(n1203), .A2(n1161), .ZN(n996) );
XNOR2_X1 U903 ( .A(n1204), .B(KEYINPUT47), .ZN(n1161) );
NAND2_X1 U904 ( .A1(n1205), .A2(n1206), .ZN(G15) );
NAND2_X1 U905 ( .A1(G113), .A2(n1157), .ZN(n1206) );
XOR2_X1 U906 ( .A(KEYINPUT31), .B(n1207), .Z(n1205) );
NOR2_X1 U907 ( .A1(G113), .A2(n1157), .ZN(n1207) );
NAND3_X1 U908 ( .A1(n1186), .A2(n1006), .A3(n1145), .ZN(n1157) );
INV_X1 U909 ( .A(n995), .ZN(n1145) );
NAND2_X1 U910 ( .A1(n1204), .A2(n1162), .ZN(n995) );
INV_X1 U911 ( .A(n1203), .ZN(n1162) );
NOR2_X1 U912 ( .A1(n1005), .A2(n1032), .ZN(n1006) );
AND3_X1 U913 ( .A1(n1208), .A2(n988), .A3(n989), .ZN(n1186) );
NAND2_X1 U914 ( .A1(n1209), .A2(n1210), .ZN(G12) );
NAND2_X1 U915 ( .A1(G110), .A2(n1211), .ZN(n1210) );
NAND2_X1 U916 ( .A1(n1150), .A2(n1212), .ZN(n1211) );
NAND2_X1 U917 ( .A1(KEYINPUT8), .A2(n1213), .ZN(n1212) );
NAND3_X1 U918 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1209) );
INV_X1 U919 ( .A(KEYINPUT8), .ZN(n1216) );
NAND2_X1 U920 ( .A1(n1217), .A2(n1213), .ZN(n1215) );
NAND2_X1 U921 ( .A1(n1150), .A2(n1218), .ZN(n1214) );
NAND2_X1 U922 ( .A1(n1219), .A2(n1213), .ZN(n1218) );
INV_X1 U923 ( .A(KEYINPUT48), .ZN(n1213) );
INV_X1 U924 ( .A(n1217), .ZN(n1150) );
NAND4_X1 U925 ( .A1(n1004), .A2(n997), .A3(n1153), .A4(n1005), .ZN(n1217) );
NAND2_X1 U926 ( .A1(n1029), .A2(n1220), .ZN(n1005) );
OR2_X1 U927 ( .A1(n1028), .A2(n1026), .ZN(n1220) );
NAND2_X1 U928 ( .A1(n1026), .A2(n1028), .ZN(n1029) );
NAND2_X1 U929 ( .A1(n1080), .A2(n1221), .ZN(n1028) );
XNOR2_X1 U930 ( .A(n1222), .B(n1223), .ZN(n1080) );
XOR2_X1 U931 ( .A(n1224), .B(n1225), .Z(n1223) );
XOR2_X1 U932 ( .A(G125), .B(G119), .Z(n1225) );
XOR2_X1 U933 ( .A(KEYINPUT40), .B(G128), .Z(n1224) );
XOR2_X1 U934 ( .A(n1226), .B(n1227), .Z(n1222) );
XOR2_X1 U935 ( .A(n1228), .B(n1229), .Z(n1227) );
NAND2_X1 U936 ( .A1(KEYINPUT46), .A2(G110), .ZN(n1229) );
NAND3_X1 U937 ( .A1(G234), .A2(n1056), .A3(G221), .ZN(n1228) );
XNOR2_X1 U938 ( .A(n1230), .B(n1231), .ZN(n1226) );
NOR2_X1 U939 ( .A1(G137), .A2(KEYINPUT54), .ZN(n1231) );
INV_X1 U940 ( .A(n1078), .ZN(n1026) );
NAND2_X1 U941 ( .A1(G217), .A2(n1232), .ZN(n1078) );
AND2_X1 U942 ( .A1(n1208), .A2(n1167), .ZN(n1153) );
INV_X1 U943 ( .A(n1014), .ZN(n1167) );
NAND2_X1 U944 ( .A1(n1016), .A2(n988), .ZN(n1014) );
NAND2_X1 U945 ( .A1(G221), .A2(n1232), .ZN(n988) );
NAND2_X1 U946 ( .A1(G234), .A2(n1233), .ZN(n1232) );
INV_X1 U947 ( .A(n989), .ZN(n1016) );
XOR2_X1 U948 ( .A(n1033), .B(KEYINPUT5), .Z(n989) );
XOR2_X1 U949 ( .A(n1234), .B(G469), .Z(n1033) );
NAND2_X1 U950 ( .A1(n1235), .A2(n1221), .ZN(n1234) );
XOR2_X1 U951 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U952 ( .A(n1238), .B(n1113), .Z(n1237) );
AND2_X1 U953 ( .A1(n1239), .A2(n1240), .ZN(n1113) );
NAND2_X1 U954 ( .A1(G101), .A2(n1241), .ZN(n1240) );
NAND2_X1 U955 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND3_X1 U956 ( .A1(n1242), .A2(n1243), .A3(n1176), .ZN(n1239) );
NAND2_X1 U957 ( .A1(G104), .A2(n1244), .ZN(n1243) );
XOR2_X1 U958 ( .A(n1245), .B(KEYINPUT33), .Z(n1242) );
OR2_X1 U959 ( .A1(n1244), .A2(G104), .ZN(n1245) );
INV_X1 U960 ( .A(G107), .ZN(n1244) );
XNOR2_X1 U961 ( .A(n1112), .B(n1246), .ZN(n1238) );
XNOR2_X1 U962 ( .A(n1219), .B(n1052), .ZN(n1112) );
INV_X1 U963 ( .A(G110), .ZN(n1219) );
XOR2_X1 U964 ( .A(n1247), .B(n1248), .Z(n1236) );
NOR2_X1 U965 ( .A1(KEYINPUT34), .A2(n1129), .ZN(n1248) );
INV_X1 U966 ( .A(n1126), .ZN(n1129) );
XNOR2_X1 U967 ( .A(n1110), .B(KEYINPUT28), .ZN(n1247) );
NOR2_X1 U968 ( .A1(n1047), .A2(G953), .ZN(n1110) );
INV_X1 U969 ( .A(G227), .ZN(n1047) );
AND2_X1 U970 ( .A1(n1160), .A2(n1249), .ZN(n1208) );
NAND2_X1 U971 ( .A1(n1017), .A2(n1250), .ZN(n1249) );
NAND4_X1 U972 ( .A1(G953), .A2(G902), .A3(n1178), .A4(n1063), .ZN(n1250) );
INV_X1 U973 ( .A(G898), .ZN(n1063) );
NAND3_X1 U974 ( .A1(n1178), .A2(n1056), .A3(G952), .ZN(n1017) );
NAND2_X1 U975 ( .A1(G237), .A2(G234), .ZN(n1178) );
NOR2_X1 U976 ( .A1(n1011), .A2(n1010), .ZN(n1160) );
INV_X1 U977 ( .A(n1030), .ZN(n1010) );
NAND2_X1 U978 ( .A1(G214), .A2(n1251), .ZN(n1030) );
XNOR2_X1 U979 ( .A(n1023), .B(n1252), .ZN(n1011) );
NOR2_X1 U980 ( .A1(KEYINPUT38), .A2(n1253), .ZN(n1252) );
XNOR2_X1 U981 ( .A(n1025), .B(KEYINPUT21), .ZN(n1253) );
AND2_X1 U982 ( .A1(G210), .A2(n1251), .ZN(n1025) );
NAND2_X1 U983 ( .A1(n1233), .A2(n1254), .ZN(n1251) );
INV_X1 U984 ( .A(G237), .ZN(n1254) );
XOR2_X1 U985 ( .A(G902), .B(KEYINPUT18), .Z(n1233) );
NAND4_X1 U986 ( .A1(n1255), .A2(n1221), .A3(n1256), .A4(n1257), .ZN(n1023) );
NAND3_X1 U987 ( .A1(n1126), .A2(n1116), .A3(G125), .ZN(n1257) );
NAND2_X1 U988 ( .A1(n1258), .A2(n1053), .ZN(n1256) );
XOR2_X1 U989 ( .A(n1116), .B(n1126), .Z(n1258) );
NAND2_X1 U990 ( .A1(n1120), .A2(n1259), .ZN(n1255) );
INV_X1 U991 ( .A(n1116), .ZN(n1259) );
XOR2_X1 U992 ( .A(n1260), .B(n1261), .Z(n1116) );
INV_X1 U993 ( .A(n1070), .ZN(n1261) );
XNOR2_X1 U994 ( .A(G113), .B(n1262), .ZN(n1070) );
NOR2_X1 U995 ( .A1(KEYINPUT39), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U996 ( .A(n1066), .B(n1264), .ZN(n1260) );
NOR2_X1 U997 ( .A1(G953), .A2(n1062), .ZN(n1264) );
INV_X1 U998 ( .A(G224), .ZN(n1062) );
XNOR2_X1 U999 ( .A(n1265), .B(n1266), .ZN(n1066) );
XOR2_X1 U1000 ( .A(G110), .B(n1267), .Z(n1266) );
XOR2_X1 U1001 ( .A(KEYINPUT43), .B(G122), .Z(n1267) );
XOR2_X1 U1002 ( .A(n1176), .B(n1268), .Z(n1265) );
XOR2_X1 U1003 ( .A(G107), .B(G104), .Z(n1268) );
NOR2_X1 U1004 ( .A1(n1126), .A2(n1053), .ZN(n1120) );
INV_X1 U1005 ( .A(n1147), .ZN(n997) );
NAND2_X1 U1006 ( .A1(n1203), .A2(n1204), .ZN(n1147) );
XOR2_X1 U1007 ( .A(n1040), .B(n1269), .Z(n1204) );
NOR2_X1 U1008 ( .A1(KEYINPUT7), .A2(n1085), .ZN(n1269) );
INV_X1 U1009 ( .A(G478), .ZN(n1085) );
NAND2_X1 U1010 ( .A1(n1083), .A2(n1221), .ZN(n1040) );
XNOR2_X1 U1011 ( .A(n1270), .B(n1271), .ZN(n1083) );
XOR2_X1 U1012 ( .A(n1272), .B(n1273), .Z(n1271) );
NAND3_X1 U1013 ( .A1(n1274), .A2(n1056), .A3(G217), .ZN(n1272) );
INV_X1 U1014 ( .A(G953), .ZN(n1056) );
XOR2_X1 U1015 ( .A(KEYINPUT17), .B(G234), .Z(n1274) );
XOR2_X1 U1016 ( .A(n1275), .B(n1276), .Z(n1270) );
NOR2_X1 U1017 ( .A1(KEYINPUT44), .A2(n1277), .ZN(n1276) );
XNOR2_X1 U1018 ( .A(G116), .B(G122), .ZN(n1277) );
XOR2_X1 U1019 ( .A(n1278), .B(G107), .Z(n1275) );
INV_X1 U1020 ( .A(G134), .ZN(n1278) );
NOR2_X1 U1021 ( .A1(n1036), .A2(n1279), .ZN(n1203) );
AND2_X1 U1022 ( .A1(G475), .A2(n1039), .ZN(n1279) );
NOR2_X1 U1023 ( .A1(n1039), .A2(G475), .ZN(n1036) );
NAND2_X1 U1024 ( .A1(n1221), .A2(n1087), .ZN(n1039) );
NAND3_X1 U1025 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1087) );
OR2_X1 U1026 ( .A1(n1283), .A2(KEYINPUT26), .ZN(n1282) );
NAND3_X1 U1027 ( .A1(KEYINPUT26), .A2(n1283), .A3(n1284), .ZN(n1281) );
INV_X1 U1028 ( .A(n1285), .ZN(n1284) );
NAND2_X1 U1029 ( .A1(n1285), .A2(n1286), .ZN(n1280) );
NAND2_X1 U1030 ( .A1(KEYINPUT26), .A2(n1287), .ZN(n1286) );
XNOR2_X1 U1031 ( .A(KEYINPUT16), .B(n1283), .ZN(n1287) );
XOR2_X1 U1032 ( .A(n1288), .B(n1289), .Z(n1283) );
XOR2_X1 U1033 ( .A(KEYINPUT6), .B(G104), .Z(n1289) );
NAND2_X1 U1034 ( .A1(KEYINPUT0), .A2(n1290), .ZN(n1288) );
XOR2_X1 U1035 ( .A(G122), .B(G113), .Z(n1290) );
XOR2_X1 U1036 ( .A(n1291), .B(n1292), .Z(n1285) );
XOR2_X1 U1037 ( .A(n1293), .B(n1230), .Z(n1292) );
XNOR2_X1 U1038 ( .A(n1294), .B(n1052), .ZN(n1230) );
XOR2_X1 U1039 ( .A(G140), .B(KEYINPUT1), .Z(n1052) );
XNOR2_X1 U1040 ( .A(G146), .B(KEYINPUT53), .ZN(n1294) );
NOR2_X1 U1041 ( .A1(KEYINPUT12), .A2(n1053), .ZN(n1293) );
INV_X1 U1042 ( .A(G125), .ZN(n1053) );
XOR2_X1 U1043 ( .A(n1295), .B(n1296), .Z(n1291) );
XOR2_X1 U1044 ( .A(G143), .B(G131), .Z(n1296) );
NAND3_X1 U1045 ( .A1(G214), .A2(n1297), .A3(KEYINPUT22), .ZN(n1295) );
XOR2_X1 U1046 ( .A(KEYINPUT52), .B(n1032), .Z(n1004) );
XOR2_X1 U1047 ( .A(n1298), .B(G472), .Z(n1032) );
NAND2_X1 U1048 ( .A1(n1299), .A2(n1221), .ZN(n1298) );
INV_X1 U1049 ( .A(G902), .ZN(n1221) );
XOR2_X1 U1050 ( .A(n1300), .B(n1100), .Z(n1299) );
INV_X1 U1051 ( .A(n1101), .ZN(n1100) );
XNOR2_X1 U1052 ( .A(n1263), .B(n1301), .ZN(n1101) );
XOR2_X1 U1053 ( .A(G113), .B(n1054), .Z(n1301) );
XOR2_X1 U1054 ( .A(n1246), .B(n1126), .Z(n1054) );
XOR2_X1 U1055 ( .A(G146), .B(n1302), .Z(n1126) );
INV_X1 U1056 ( .A(n1273), .ZN(n1302) );
XNOR2_X1 U1057 ( .A(G128), .B(G143), .ZN(n1273) );
XOR2_X1 U1058 ( .A(G131), .B(n1303), .Z(n1246) );
XOR2_X1 U1059 ( .A(G137), .B(G134), .Z(n1303) );
XOR2_X1 U1060 ( .A(G116), .B(G119), .Z(n1263) );
NOR2_X1 U1061 ( .A1(KEYINPUT2), .A2(n1094), .ZN(n1300) );
XNOR2_X1 U1062 ( .A(n1304), .B(n1176), .ZN(n1094) );
INV_X1 U1063 ( .A(G101), .ZN(n1176) );
NAND2_X1 U1064 ( .A1(G210), .A2(n1297), .ZN(n1304) );
NOR2_X1 U1065 ( .A1(G953), .A2(G237), .ZN(n1297) );
endmodule


