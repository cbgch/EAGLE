//Key = 0010100110111111010011010110110111100000001001111111111100010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358;

NAND3_X1 U742 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(G9) );
NAND2_X1 U743 ( .A1(G107), .A2(n1044), .ZN(n1043) );
OR3_X1 U744 ( .A1(n1044), .A2(G107), .A3(n1045), .ZN(n1042) );
INV_X1 U745 ( .A(KEYINPUT33), .ZN(n1044) );
NAND2_X1 U746 ( .A1(n1046), .A2(n1045), .ZN(n1041) );
NAND2_X1 U747 ( .A1(n1047), .A2(KEYINPUT33), .ZN(n1046) );
XNOR2_X1 U748 ( .A(G107), .B(KEYINPUT43), .ZN(n1047) );
NOR2_X1 U749 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR3_X1 U750 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
NOR4_X1 U751 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1051) );
NOR3_X1 U752 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1053) );
NOR2_X1 U753 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
INV_X1 U754 ( .A(n1062), .ZN(n1061) );
XNOR2_X1 U755 ( .A(n1063), .B(KEYINPUT1), .ZN(n1060) );
NOR2_X1 U756 ( .A1(n1064), .A2(n1065), .ZN(n1058) );
NOR2_X1 U757 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U758 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
AND2_X1 U759 ( .A1(n1070), .A2(n1063), .ZN(n1057) );
NAND3_X1 U760 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1050) );
NAND4_X1 U761 ( .A1(n1063), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1073) );
NAND2_X1 U762 ( .A1(n1077), .A2(n1056), .ZN(n1076) );
NAND3_X1 U763 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
INV_X1 U764 ( .A(KEYINPUT15), .ZN(n1079) );
NAND3_X1 U765 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1075) );
INV_X1 U766 ( .A(n1056), .ZN(n1083) );
NAND2_X1 U767 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
OR2_X1 U768 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U769 ( .A1(n1080), .A2(n1088), .ZN(n1081) );
NAND2_X1 U770 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND3_X1 U771 ( .A1(G221), .A2(n1091), .A3(n1092), .ZN(n1090) );
NAND2_X1 U772 ( .A1(KEYINPUT15), .A2(n1078), .ZN(n1089) );
NOR3_X1 U773 ( .A1(n1093), .A2(G953), .A3(G952), .ZN(n1048) );
INV_X1 U774 ( .A(n1071), .ZN(n1093) );
NAND4_X1 U775 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1071) );
NOR4_X1 U776 ( .A1(n1098), .A2(n1099), .A3(n1054), .A4(n1100), .ZN(n1097) );
XNOR2_X1 U777 ( .A(n1101), .B(n1102), .ZN(n1099) );
INV_X1 U778 ( .A(n1103), .ZN(n1098) );
NOR3_X1 U779 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1096) );
NOR3_X1 U780 ( .A1(n1107), .A2(KEYINPUT38), .A3(n1108), .ZN(n1106) );
AND2_X1 U781 ( .A1(n1107), .A2(KEYINPUT38), .ZN(n1105) );
XOR2_X1 U782 ( .A(n1109), .B(n1110), .Z(n1104) );
XOR2_X1 U783 ( .A(n1111), .B(n1112), .Z(n1095) );
XOR2_X1 U784 ( .A(KEYINPUT42), .B(KEYINPUT10), .Z(n1112) );
XNOR2_X1 U785 ( .A(n1113), .B(n1114), .ZN(n1111) );
XNOR2_X1 U786 ( .A(n1115), .B(KEYINPUT0), .ZN(n1094) );
XOR2_X1 U787 ( .A(n1116), .B(n1117), .Z(G72) );
XOR2_X1 U788 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND2_X1 U789 ( .A1(G953), .A2(n1120), .ZN(n1119) );
NAND2_X1 U790 ( .A1(G900), .A2(G227), .ZN(n1120) );
NAND2_X1 U791 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
NAND2_X1 U792 ( .A1(G953), .A2(n1123), .ZN(n1122) );
XOR2_X1 U793 ( .A(n1124), .B(n1125), .Z(n1121) );
XNOR2_X1 U794 ( .A(n1126), .B(n1127), .ZN(n1125) );
XNOR2_X1 U795 ( .A(n1128), .B(n1129), .ZN(n1126) );
NAND3_X1 U796 ( .A1(n1130), .A2(n1131), .A3(KEYINPUT52), .ZN(n1129) );
OR3_X1 U797 ( .A1(n1132), .A2(G134), .A3(KEYINPUT2), .ZN(n1131) );
NAND2_X1 U798 ( .A1(n1133), .A2(KEYINPUT2), .ZN(n1130) );
XNOR2_X1 U799 ( .A(G134), .B(n1134), .ZN(n1133) );
NAND2_X1 U800 ( .A1(KEYINPUT49), .A2(n1132), .ZN(n1134) );
NAND2_X1 U801 ( .A1(n1135), .A2(KEYINPUT12), .ZN(n1128) );
XNOR2_X1 U802 ( .A(n1136), .B(KEYINPUT35), .ZN(n1135) );
XOR2_X1 U803 ( .A(n1137), .B(G131), .Z(n1124) );
XNOR2_X1 U804 ( .A(KEYINPUT30), .B(KEYINPUT16), .ZN(n1137) );
NOR2_X1 U805 ( .A1(n1138), .A2(G953), .ZN(n1116) );
AND2_X1 U806 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U807 ( .A(n1141), .B(n1142), .Z(G69) );
XOR2_X1 U808 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U809 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XNOR2_X1 U810 ( .A(KEYINPUT41), .B(n1072), .ZN(n1146) );
NAND2_X1 U811 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
INV_X1 U812 ( .A(n1149), .ZN(n1148) );
XOR2_X1 U813 ( .A(n1150), .B(n1151), .Z(n1147) );
NOR2_X1 U814 ( .A1(KEYINPUT36), .A2(n1152), .ZN(n1151) );
NAND2_X1 U815 ( .A1(G953), .A2(n1153), .ZN(n1141) );
NAND2_X1 U816 ( .A1(G898), .A2(G224), .ZN(n1153) );
NOR2_X1 U817 ( .A1(n1154), .A2(n1155), .ZN(G66) );
XOR2_X1 U818 ( .A(n1156), .B(KEYINPUT48), .Z(n1155) );
NAND2_X1 U819 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
OR3_X1 U820 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1158) );
XOR2_X1 U821 ( .A(n1162), .B(KEYINPUT40), .Z(n1157) );
NAND2_X1 U822 ( .A1(n1163), .A2(n1161), .ZN(n1162) );
XOR2_X1 U823 ( .A(KEYINPUT29), .B(n1164), .Z(n1163) );
NOR2_X1 U824 ( .A1(n1160), .A2(n1159), .ZN(n1164) );
NOR2_X1 U825 ( .A1(n1154), .A2(n1165), .ZN(G63) );
XOR2_X1 U826 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U827 ( .A(KEYINPUT58), .B(n1168), .Z(n1167) );
NOR2_X1 U828 ( .A1(n1114), .A2(n1159), .ZN(n1168) );
NOR2_X1 U829 ( .A1(n1154), .A2(n1169), .ZN(G60) );
XOR2_X1 U830 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U831 ( .A1(n1107), .A2(n1159), .ZN(n1170) );
XNOR2_X1 U832 ( .A(G104), .B(n1172), .ZN(G6) );
NOR2_X1 U833 ( .A1(n1154), .A2(n1173), .ZN(G57) );
XOR2_X1 U834 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U835 ( .A(n1176), .B(n1177), .ZN(n1175) );
XNOR2_X1 U836 ( .A(n1178), .B(n1179), .ZN(n1177) );
NOR2_X1 U837 ( .A1(KEYINPUT56), .A2(n1180), .ZN(n1179) );
NOR2_X1 U838 ( .A1(KEYINPUT19), .A2(n1181), .ZN(n1178) );
XOR2_X1 U839 ( .A(n1182), .B(n1183), .Z(n1174) );
NOR3_X1 U840 ( .A1(n1159), .A2(KEYINPUT18), .A3(n1184), .ZN(n1183) );
XOR2_X1 U841 ( .A(n1185), .B(n1186), .Z(n1182) );
NOR2_X1 U842 ( .A1(KEYINPUT39), .A2(n1187), .ZN(n1186) );
NOR2_X1 U843 ( .A1(n1154), .A2(n1188), .ZN(G54) );
XOR2_X1 U844 ( .A(n1189), .B(n1190), .Z(n1188) );
XNOR2_X1 U845 ( .A(n1176), .B(n1191), .ZN(n1190) );
NAND2_X1 U846 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
OR2_X1 U847 ( .A1(n1194), .A2(KEYINPUT61), .ZN(n1193) );
NAND3_X1 U848 ( .A1(n1195), .A2(n1196), .A3(KEYINPUT61), .ZN(n1192) );
XOR2_X1 U849 ( .A(n1197), .B(n1198), .Z(n1189) );
NOR2_X1 U850 ( .A1(n1199), .A2(n1159), .ZN(n1198) );
INV_X1 U851 ( .A(G469), .ZN(n1199) );
NAND3_X1 U852 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1197) );
NAND2_X1 U853 ( .A1(G140), .A2(n1203), .ZN(n1201) );
XNOR2_X1 U854 ( .A(G110), .B(n1204), .ZN(n1203) );
NAND3_X1 U855 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1200) );
NOR2_X1 U856 ( .A1(n1154), .A2(n1207), .ZN(G51) );
XOR2_X1 U857 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U858 ( .A(n1210), .B(n1211), .Z(n1209) );
NOR2_X1 U859 ( .A1(n1110), .A2(n1159), .ZN(n1211) );
NAND2_X1 U860 ( .A1(G902), .A2(n1052), .ZN(n1159) );
NAND3_X1 U861 ( .A1(n1140), .A2(n1212), .A3(n1145), .ZN(n1052) );
AND4_X1 U862 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1145) );
AND4_X1 U863 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1172), .ZN(n1216) );
NAND4_X1 U864 ( .A1(n1086), .A2(n1220), .A3(n1074), .A4(n1221), .ZN(n1172) );
NOR2_X1 U865 ( .A1(n1222), .A2(n1223), .ZN(n1215) );
INV_X1 U866 ( .A(n1045), .ZN(n1222) );
NAND4_X1 U867 ( .A1(n1087), .A2(n1220), .A3(n1074), .A4(n1221), .ZN(n1045) );
NAND2_X1 U868 ( .A1(n1224), .A2(n1225), .ZN(n1213) );
XOR2_X1 U869 ( .A(n1221), .B(KEYINPUT22), .Z(n1224) );
XNOR2_X1 U870 ( .A(KEYINPUT8), .B(n1139), .ZN(n1212) );
AND4_X1 U871 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1140) );
AND4_X1 U872 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1229) );
NAND2_X1 U873 ( .A1(n1234), .A2(n1067), .ZN(n1228) );
NAND2_X1 U874 ( .A1(n1063), .A2(n1235), .ZN(n1226) );
XNOR2_X1 U875 ( .A(KEYINPUT63), .B(n1236), .ZN(n1235) );
NOR2_X1 U876 ( .A1(n1237), .A2(n1238), .ZN(n1210) );
XOR2_X1 U877 ( .A(n1239), .B(KEYINPUT31), .Z(n1238) );
NAND2_X1 U878 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NOR2_X1 U879 ( .A1(n1242), .A2(n1241), .ZN(n1237) );
XNOR2_X1 U880 ( .A(n1240), .B(KEYINPUT17), .ZN(n1242) );
NOR2_X1 U881 ( .A1(n1072), .A2(G952), .ZN(n1154) );
XNOR2_X1 U882 ( .A(n1243), .B(n1244), .ZN(G48) );
NAND2_X1 U883 ( .A1(KEYINPUT53), .A2(n1230), .ZN(n1243) );
NAND4_X1 U884 ( .A1(n1245), .A2(n1246), .A3(n1220), .A4(n1100), .ZN(n1230) );
XNOR2_X1 U885 ( .A(n1227), .B(n1247), .ZN(G45) );
NOR2_X1 U886 ( .A1(KEYINPUT37), .A2(n1248), .ZN(n1247) );
NAND3_X1 U887 ( .A1(n1070), .A2(n1220), .A3(n1249), .ZN(n1227) );
NOR3_X1 U888 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1249) );
XNOR2_X1 U889 ( .A(G140), .B(n1233), .ZN(G42) );
NAND3_X1 U890 ( .A1(n1062), .A2(n1086), .A3(n1253), .ZN(n1233) );
XOR2_X1 U891 ( .A(n1232), .B(n1254), .Z(G39) );
NAND2_X1 U892 ( .A1(KEYINPUT47), .A2(G137), .ZN(n1254) );
NAND2_X1 U893 ( .A1(n1253), .A2(n1255), .ZN(n1232) );
XNOR2_X1 U894 ( .A(G134), .B(n1139), .ZN(G36) );
NAND3_X1 U895 ( .A1(n1070), .A2(n1087), .A3(n1253), .ZN(n1139) );
AND3_X1 U896 ( .A1(n1078), .A2(n1256), .A3(n1063), .ZN(n1253) );
XOR2_X1 U897 ( .A(G131), .B(n1257), .Z(G33) );
NOR2_X1 U898 ( .A1(n1258), .A2(n1236), .ZN(n1257) );
NAND3_X1 U899 ( .A1(n1070), .A2(n1078), .A3(n1246), .ZN(n1236) );
XNOR2_X1 U900 ( .A(n1063), .B(KEYINPUT9), .ZN(n1258) );
NOR2_X1 U901 ( .A1(n1068), .A2(n1115), .ZN(n1063) );
INV_X1 U902 ( .A(n1069), .ZN(n1115) );
XNOR2_X1 U903 ( .A(G128), .B(n1231), .ZN(G30) );
NAND4_X1 U904 ( .A1(n1245), .A2(n1087), .A3(n1259), .A4(n1220), .ZN(n1231) );
NOR2_X1 U905 ( .A1(n1252), .A2(n1260), .ZN(n1259) );
INV_X1 U906 ( .A(n1256), .ZN(n1252) );
XNOR2_X1 U907 ( .A(G101), .B(n1219), .ZN(G3) );
NAND4_X1 U908 ( .A1(n1080), .A2(n1070), .A3(n1220), .A4(n1221), .ZN(n1219) );
NAND2_X1 U909 ( .A1(n1261), .A2(n1262), .ZN(G27) );
NAND2_X1 U910 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
XOR2_X1 U911 ( .A(KEYINPUT23), .B(n1265), .Z(n1261) );
NOR2_X1 U912 ( .A1(n1263), .A2(n1264), .ZN(n1265) );
INV_X1 U913 ( .A(G125), .ZN(n1264) );
AND2_X1 U914 ( .A1(n1266), .A2(n1067), .ZN(n1263) );
XNOR2_X1 U915 ( .A(n1234), .B(KEYINPUT25), .ZN(n1266) );
AND3_X1 U916 ( .A1(n1062), .A2(n1084), .A3(n1246), .ZN(n1234) );
AND2_X1 U917 ( .A1(n1086), .A2(n1256), .ZN(n1246) );
NAND2_X1 U918 ( .A1(n1056), .A2(n1267), .ZN(n1256) );
NAND4_X1 U919 ( .A1(G953), .A2(G902), .A3(n1268), .A4(n1123), .ZN(n1267) );
INV_X1 U920 ( .A(G900), .ZN(n1123) );
XNOR2_X1 U921 ( .A(G122), .B(n1214), .ZN(G24) );
NAND4_X1 U922 ( .A1(n1269), .A2(n1074), .A3(n1270), .A4(n1271), .ZN(n1214) );
INV_X1 U923 ( .A(n1065), .ZN(n1074) );
NAND2_X1 U924 ( .A1(n1272), .A2(n1273), .ZN(n1065) );
XNOR2_X1 U925 ( .A(n1274), .B(n1223), .ZN(G21) );
AND2_X1 U926 ( .A1(n1255), .A2(n1269), .ZN(n1223) );
NOR3_X1 U927 ( .A1(n1272), .A2(n1260), .A3(n1055), .ZN(n1255) );
INV_X1 U928 ( .A(n1080), .ZN(n1055) );
XNOR2_X1 U929 ( .A(G116), .B(n1218), .ZN(G18) );
NAND3_X1 U930 ( .A1(n1070), .A2(n1087), .A3(n1269), .ZN(n1218) );
NOR2_X1 U931 ( .A1(n1271), .A2(n1250), .ZN(n1087) );
INV_X1 U932 ( .A(n1270), .ZN(n1250) );
XOR2_X1 U933 ( .A(n1217), .B(n1275), .Z(G15) );
XOR2_X1 U934 ( .A(KEYINPUT32), .B(G113), .Z(n1275) );
NAND3_X1 U935 ( .A1(n1269), .A2(n1070), .A3(n1086), .ZN(n1217) );
NOR2_X1 U936 ( .A1(n1270), .A2(n1251), .ZN(n1086) );
INV_X1 U937 ( .A(n1271), .ZN(n1251) );
AND2_X1 U938 ( .A1(n1245), .A2(n1273), .ZN(n1070) );
XNOR2_X1 U939 ( .A(n1260), .B(KEYINPUT14), .ZN(n1273) );
AND3_X1 U940 ( .A1(n1067), .A2(n1221), .A3(n1084), .ZN(n1269) );
INV_X1 U941 ( .A(n1054), .ZN(n1084) );
NAND2_X1 U942 ( .A1(n1092), .A2(n1276), .ZN(n1054) );
NAND2_X1 U943 ( .A1(G221), .A2(n1091), .ZN(n1276) );
XNOR2_X1 U944 ( .A(n1205), .B(n1277), .ZN(G12) );
AND2_X1 U945 ( .A1(n1221), .A2(n1225), .ZN(n1277) );
AND3_X1 U946 ( .A1(n1080), .A2(n1220), .A3(n1062), .ZN(n1225) );
NOR2_X1 U947 ( .A1(n1245), .A2(n1260), .ZN(n1062) );
INV_X1 U948 ( .A(n1100), .ZN(n1260) );
XNOR2_X1 U949 ( .A(n1160), .B(n1278), .ZN(n1100) );
AND2_X1 U950 ( .A1(n1161), .A2(n1279), .ZN(n1278) );
NAND2_X1 U951 ( .A1(n1280), .A2(n1281), .ZN(n1161) );
NAND2_X1 U952 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
XOR2_X1 U953 ( .A(KEYINPUT50), .B(n1284), .Z(n1280) );
NOR2_X1 U954 ( .A1(n1283), .A2(n1282), .ZN(n1284) );
XOR2_X1 U955 ( .A(n1285), .B(n1286), .Z(n1282) );
NAND2_X1 U956 ( .A1(KEYINPUT54), .A2(n1132), .ZN(n1286) );
NAND3_X1 U957 ( .A1(G234), .A2(n1072), .A3(G221), .ZN(n1285) );
XNOR2_X1 U958 ( .A(n1287), .B(n1288), .ZN(n1283) );
XNOR2_X1 U959 ( .A(n1289), .B(n1290), .ZN(n1288) );
INV_X1 U960 ( .A(n1136), .ZN(n1289) );
XNOR2_X1 U961 ( .A(G119), .B(G110), .ZN(n1287) );
NAND2_X1 U962 ( .A1(G217), .A2(n1091), .ZN(n1160) );
INV_X1 U963 ( .A(n1272), .ZN(n1245) );
XNOR2_X1 U964 ( .A(n1101), .B(n1291), .ZN(n1272) );
NOR2_X1 U965 ( .A1(KEYINPUT6), .A2(n1102), .ZN(n1291) );
XOR2_X1 U966 ( .A(n1184), .B(KEYINPUT11), .Z(n1102) );
INV_X1 U967 ( .A(G472), .ZN(n1184) );
NAND2_X1 U968 ( .A1(n1292), .A2(n1279), .ZN(n1101) );
XOR2_X1 U969 ( .A(n1293), .B(n1294), .Z(n1292) );
XNOR2_X1 U970 ( .A(n1176), .B(n1180), .ZN(n1294) );
NAND2_X1 U971 ( .A1(n1295), .A2(n1296), .ZN(n1180) );
NAND2_X1 U972 ( .A1(n1297), .A2(n1274), .ZN(n1296) );
INV_X1 U973 ( .A(G119), .ZN(n1274) );
XOR2_X1 U974 ( .A(KEYINPUT21), .B(n1298), .Z(n1297) );
NAND2_X1 U975 ( .A1(n1298), .A2(G119), .ZN(n1295) );
XNOR2_X1 U976 ( .A(n1181), .B(n1299), .ZN(n1293) );
XNOR2_X1 U977 ( .A(n1185), .B(n1300), .ZN(n1299) );
NAND2_X1 U978 ( .A1(G210), .A2(n1301), .ZN(n1185) );
XNOR2_X1 U979 ( .A(n1302), .B(KEYINPUT27), .ZN(n1181) );
AND2_X1 U980 ( .A1(n1078), .A2(n1067), .ZN(n1220) );
AND2_X1 U981 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U982 ( .A1(G214), .A2(n1303), .ZN(n1069) );
XNOR2_X1 U983 ( .A(n1304), .B(n1109), .ZN(n1068) );
NAND3_X1 U984 ( .A1(n1305), .A2(n1279), .A3(n1306), .ZN(n1109) );
XOR2_X1 U985 ( .A(KEYINPUT7), .B(n1307), .Z(n1306) );
NOR2_X1 U986 ( .A1(n1308), .A2(n1208), .ZN(n1307) );
NAND2_X1 U987 ( .A1(n1308), .A2(n1208), .ZN(n1305) );
XNOR2_X1 U988 ( .A(n1150), .B(n1309), .ZN(n1208) );
XOR2_X1 U989 ( .A(KEYINPUT46), .B(n1152), .Z(n1309) );
XNOR2_X1 U990 ( .A(G122), .B(n1205), .ZN(n1152) );
XOR2_X1 U991 ( .A(n1310), .B(n1311), .Z(n1150) );
XNOR2_X1 U992 ( .A(G119), .B(n1298), .ZN(n1310) );
XOR2_X1 U993 ( .A(G113), .B(G116), .Z(n1298) );
XNOR2_X1 U994 ( .A(n1240), .B(n1312), .ZN(n1308) );
XNOR2_X1 U995 ( .A(n1241), .B(KEYINPUT13), .ZN(n1312) );
NAND2_X1 U996 ( .A1(G224), .A2(n1072), .ZN(n1241) );
XNOR2_X1 U997 ( .A(G125), .B(n1302), .ZN(n1240) );
XNOR2_X1 U998 ( .A(G146), .B(n1313), .ZN(n1302) );
NAND2_X1 U999 ( .A1(KEYINPUT26), .A2(n1110), .ZN(n1304) );
NAND2_X1 U1000 ( .A1(G210), .A2(n1303), .ZN(n1110) );
NAND2_X1 U1001 ( .A1(n1314), .A2(n1279), .ZN(n1303) );
INV_X1 U1002 ( .A(G902), .ZN(n1279) );
INV_X1 U1003 ( .A(G237), .ZN(n1314) );
NOR2_X1 U1004 ( .A1(n1092), .A2(n1315), .ZN(n1078) );
AND2_X1 U1005 ( .A1(G221), .A2(n1091), .ZN(n1315) );
NAND2_X1 U1006 ( .A1(n1316), .A2(G234), .ZN(n1091) );
XNOR2_X1 U1007 ( .A(G902), .B(KEYINPUT44), .ZN(n1316) );
XNOR2_X1 U1008 ( .A(G469), .B(n1317), .ZN(n1092) );
NOR2_X1 U1009 ( .A1(n1318), .A2(G902), .ZN(n1317) );
NOR2_X1 U1010 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
XOR2_X1 U1011 ( .A(n1321), .B(KEYINPUT59), .Z(n1320) );
NAND2_X1 U1012 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NOR2_X1 U1013 ( .A1(n1322), .A2(n1323), .ZN(n1319) );
NAND3_X1 U1014 ( .A1(n1324), .A2(n1325), .A3(n1202), .ZN(n1323) );
NAND3_X1 U1015 ( .A1(n1326), .A2(n1206), .A3(G110), .ZN(n1202) );
NAND2_X1 U1016 ( .A1(n1327), .A2(n1326), .ZN(n1325) );
XNOR2_X1 U1017 ( .A(KEYINPUT3), .B(n1328), .ZN(n1327) );
NAND3_X1 U1018 ( .A1(n1329), .A2(n1330), .A3(n1204), .ZN(n1324) );
INV_X1 U1019 ( .A(n1326), .ZN(n1204) );
NAND2_X1 U1020 ( .A1(G227), .A2(n1072), .ZN(n1326) );
NAND2_X1 U1021 ( .A1(G110), .A2(n1206), .ZN(n1330) );
XOR2_X1 U1022 ( .A(n1328), .B(KEYINPUT3), .Z(n1329) );
NAND2_X1 U1023 ( .A1(n1331), .A2(n1205), .ZN(n1328) );
XNOR2_X1 U1024 ( .A(G140), .B(KEYINPUT20), .ZN(n1331) );
XNOR2_X1 U1025 ( .A(n1332), .B(n1194), .ZN(n1322) );
XNOR2_X1 U1026 ( .A(n1196), .B(n1195), .ZN(n1194) );
XOR2_X1 U1027 ( .A(n1311), .B(KEYINPUT62), .Z(n1195) );
XOR2_X1 U1028 ( .A(n1333), .B(n1187), .Z(n1311) );
INV_X1 U1029 ( .A(n1300), .ZN(n1187) );
XOR2_X1 U1030 ( .A(G101), .B(KEYINPUT55), .Z(n1300) );
XNOR2_X1 U1031 ( .A(G104), .B(G107), .ZN(n1333) );
XOR2_X1 U1032 ( .A(n1127), .B(KEYINPUT60), .Z(n1196) );
NAND2_X1 U1033 ( .A1(n1334), .A2(n1335), .ZN(n1127) );
OR2_X1 U1034 ( .A1(n1290), .A2(G143), .ZN(n1335) );
NAND2_X1 U1035 ( .A1(n1336), .A2(G143), .ZN(n1334) );
XOR2_X1 U1036 ( .A(KEYINPUT24), .B(n1290), .Z(n1336) );
XNOR2_X1 U1037 ( .A(G128), .B(n1244), .ZN(n1290) );
INV_X1 U1038 ( .A(n1176), .ZN(n1332) );
XNOR2_X1 U1039 ( .A(n1337), .B(G131), .ZN(n1176) );
NAND2_X1 U1040 ( .A1(KEYINPUT45), .A2(n1338), .ZN(n1337) );
XNOR2_X1 U1041 ( .A(n1132), .B(G134), .ZN(n1338) );
INV_X1 U1042 ( .A(G137), .ZN(n1132) );
NOR2_X1 U1043 ( .A1(n1270), .A2(n1271), .ZN(n1080) );
NAND2_X1 U1044 ( .A1(n1339), .A2(n1103), .ZN(n1271) );
NAND2_X1 U1045 ( .A1(n1108), .A2(n1107), .ZN(n1103) );
OR2_X1 U1046 ( .A1(n1107), .A2(n1108), .ZN(n1339) );
NOR2_X1 U1047 ( .A1(n1171), .A2(G902), .ZN(n1108) );
XNOR2_X1 U1048 ( .A(n1340), .B(G113), .ZN(n1171) );
XOR2_X1 U1049 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1050 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1051 ( .A(G122), .B(G104), .Z(n1344) );
XOR2_X1 U1052 ( .A(KEYINPUT5), .B(G131), .Z(n1343) );
XOR2_X1 U1053 ( .A(n1345), .B(n1346), .Z(n1341) );
XNOR2_X1 U1054 ( .A(n1347), .B(n1136), .ZN(n1346) );
XNOR2_X1 U1055 ( .A(G125), .B(n1206), .ZN(n1136) );
INV_X1 U1056 ( .A(G140), .ZN(n1206) );
NAND2_X1 U1057 ( .A1(G214), .A2(n1301), .ZN(n1347) );
NOR2_X1 U1058 ( .A1(G953), .A2(G237), .ZN(n1301) );
XNOR2_X1 U1059 ( .A(n1348), .B(n1349), .ZN(n1345) );
NAND2_X1 U1060 ( .A1(KEYINPUT51), .A2(n1244), .ZN(n1349) );
INV_X1 U1061 ( .A(G146), .ZN(n1244) );
NAND2_X1 U1062 ( .A1(n1350), .A2(KEYINPUT28), .ZN(n1348) );
XNOR2_X1 U1063 ( .A(G143), .B(KEYINPUT34), .ZN(n1350) );
INV_X1 U1064 ( .A(G475), .ZN(n1107) );
XNOR2_X1 U1065 ( .A(n1113), .B(n1351), .ZN(n1270) );
NOR2_X1 U1066 ( .A1(KEYINPUT57), .A2(n1114), .ZN(n1351) );
INV_X1 U1067 ( .A(G478), .ZN(n1114) );
OR2_X1 U1068 ( .A1(n1166), .A2(G902), .ZN(n1113) );
XNOR2_X1 U1069 ( .A(n1352), .B(n1353), .ZN(n1166) );
XOR2_X1 U1070 ( .A(n1354), .B(n1355), .Z(n1353) );
NAND3_X1 U1071 ( .A1(G217), .A2(n1072), .A3(G234), .ZN(n1355) );
NAND2_X1 U1072 ( .A1(n1356), .A2(KEYINPUT4), .ZN(n1354) );
XNOR2_X1 U1073 ( .A(G134), .B(n1313), .ZN(n1356) );
XNOR2_X1 U1074 ( .A(G128), .B(n1248), .ZN(n1313) );
INV_X1 U1075 ( .A(G143), .ZN(n1248) );
XNOR2_X1 U1076 ( .A(G107), .B(n1357), .ZN(n1352) );
XOR2_X1 U1077 ( .A(G122), .B(G116), .Z(n1357) );
NAND2_X1 U1078 ( .A1(n1056), .A2(n1358), .ZN(n1221) );
NAND3_X1 U1079 ( .A1(G902), .A2(n1268), .A3(n1149), .ZN(n1358) );
NOR2_X1 U1080 ( .A1(n1072), .A2(G898), .ZN(n1149) );
NAND3_X1 U1081 ( .A1(n1268), .A2(n1072), .A3(G952), .ZN(n1056) );
INV_X1 U1082 ( .A(G953), .ZN(n1072) );
NAND2_X1 U1083 ( .A1(G237), .A2(G234), .ZN(n1268) );
INV_X1 U1084 ( .A(G110), .ZN(n1205) );
endmodule


