//Key = 1111101010100001100010100011011001001111101011100101000100001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339;

XOR2_X1 U725 ( .A(G107), .B(n1019), .Z(G9) );
NOR2_X1 U726 ( .A1(n1020), .A2(n1021), .ZN(G75) );
NOR4_X1 U727 ( .A1(G953), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1021) );
NOR2_X1 U728 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U729 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR3_X1 U730 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NOR2_X1 U731 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
AND2_X1 U732 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR2_X1 U733 ( .A1(n1036), .A2(n1037), .ZN(n1032) );
NOR3_X1 U734 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1036) );
AND4_X1 U735 ( .A1(KEYINPUT45), .A2(n1041), .A3(n1042), .A4(G214), .ZN(n1040) );
INV_X1 U736 ( .A(n1043), .ZN(n1041) );
NOR2_X1 U737 ( .A1(KEYINPUT45), .A2(n1044), .ZN(n1039) );
NOR3_X1 U738 ( .A1(n1044), .A2(n1045), .A3(n1037), .ZN(n1027) );
NOR2_X1 U739 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U740 ( .A1(n1048), .A2(n1029), .ZN(n1047) );
NOR2_X1 U741 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U742 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
XOR2_X1 U743 ( .A(n1053), .B(KEYINPUT56), .Z(n1051) );
NOR2_X1 U744 ( .A1(n1054), .A2(n1031), .ZN(n1046) );
NOR2_X1 U745 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
INV_X1 U746 ( .A(n1035), .ZN(n1044) );
NOR3_X1 U747 ( .A1(n1022), .A2(G953), .A3(G952), .ZN(n1020) );
AND4_X1 U748 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1022) );
NOR4_X1 U749 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1060) );
NOR2_X1 U750 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
XNOR2_X1 U751 ( .A(G469), .B(KEYINPUT19), .ZN(n1066) );
INV_X1 U752 ( .A(n1067), .ZN(n1065) );
INV_X1 U753 ( .A(n1052), .ZN(n1063) );
INV_X1 U754 ( .A(n1068), .ZN(n1061) );
NOR3_X1 U755 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1059) );
NOR2_X1 U756 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
INV_X1 U757 ( .A(KEYINPUT28), .ZN(n1073) );
NOR2_X1 U758 ( .A1(G214), .A2(n1074), .ZN(n1072) );
NOR2_X1 U759 ( .A1(KEYINPUT28), .A2(n1035), .ZN(n1070) );
XOR2_X1 U760 ( .A(KEYINPUT54), .B(n1075), .Z(n1069) );
NOR2_X1 U761 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U762 ( .A(n1078), .B(KEYINPUT31), .Z(n1077) );
XOR2_X1 U763 ( .A(n1079), .B(n1080), .Z(G72) );
XOR2_X1 U764 ( .A(n1081), .B(n1082), .Z(n1080) );
NOR2_X1 U765 ( .A1(G953), .A2(n1083), .ZN(n1082) );
NAND2_X1 U766 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
INV_X1 U767 ( .A(n1086), .ZN(n1085) );
XOR2_X1 U768 ( .A(n1087), .B(n1088), .Z(n1084) );
XNOR2_X1 U769 ( .A(n1089), .B(n1090), .ZN(n1088) );
NAND2_X1 U770 ( .A1(n1091), .A2(KEYINPUT63), .ZN(n1089) );
XNOR2_X1 U771 ( .A(G137), .B(KEYINPUT17), .ZN(n1091) );
XOR2_X1 U772 ( .A(n1092), .B(n1093), .Z(n1087) );
XNOR2_X1 U773 ( .A(KEYINPUT60), .B(n1094), .ZN(n1093) );
NOR2_X1 U774 ( .A1(KEYINPUT18), .A2(n1095), .ZN(n1094) );
XOR2_X1 U775 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U776 ( .A1(G125), .A2(KEYINPUT11), .ZN(n1097) );
INV_X1 U777 ( .A(G140), .ZN(n1096) );
NAND2_X1 U778 ( .A1(G953), .A2(n1098), .ZN(n1079) );
NAND2_X1 U779 ( .A1(G900), .A2(G227), .ZN(n1098) );
NAND3_X1 U780 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(G69) );
NAND3_X1 U781 ( .A1(n1102), .A2(n1103), .A3(KEYINPUT4), .ZN(n1101) );
NAND2_X1 U782 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NAND2_X1 U783 ( .A1(G953), .A2(n1106), .ZN(n1105) );
NAND3_X1 U784 ( .A1(n1107), .A2(n1108), .A3(G953), .ZN(n1100) );
NAND2_X1 U785 ( .A1(KEYINPUT4), .A2(n1106), .ZN(n1108) );
XOR2_X1 U786 ( .A(KEYINPUT16), .B(G224), .Z(n1106) );
INV_X1 U787 ( .A(n1103), .ZN(n1107) );
NAND2_X1 U788 ( .A1(n1109), .A2(n1110), .ZN(n1099) );
XOR2_X1 U789 ( .A(n1103), .B(n1111), .Z(n1109) );
NAND2_X1 U790 ( .A1(n1112), .A2(n1104), .ZN(n1103) );
INV_X1 U791 ( .A(n1113), .ZN(n1104) );
XOR2_X1 U792 ( .A(n1114), .B(n1115), .Z(n1112) );
XNOR2_X1 U793 ( .A(n1116), .B(n1117), .ZN(n1114) );
NOR2_X1 U794 ( .A1(KEYINPUT48), .A2(n1118), .ZN(n1117) );
NOR2_X1 U795 ( .A1(n1119), .A2(n1120), .ZN(G66) );
XOR2_X1 U796 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U797 ( .A(KEYINPUT1), .B(n1123), .Z(n1122) );
NOR2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NOR2_X1 U799 ( .A1(n1119), .A2(n1126), .ZN(G63) );
XOR2_X1 U800 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U801 ( .A(KEYINPUT7), .B(n1129), .Z(n1128) );
NOR2_X1 U802 ( .A1(n1078), .A2(n1125), .ZN(n1129) );
NOR2_X1 U803 ( .A1(n1130), .A2(n1131), .ZN(G60) );
XNOR2_X1 U804 ( .A(n1132), .B(n1133), .ZN(n1131) );
AND2_X1 U805 ( .A1(G475), .A2(n1134), .ZN(n1133) );
XNOR2_X1 U806 ( .A(n1119), .B(KEYINPUT27), .ZN(n1130) );
XNOR2_X1 U807 ( .A(G104), .B(n1135), .ZN(G6) );
NOR2_X1 U808 ( .A1(n1119), .A2(n1136), .ZN(G57) );
XOR2_X1 U809 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U810 ( .A(n1139), .B(G101), .Z(n1138) );
NAND2_X1 U811 ( .A1(KEYINPUT29), .A2(n1140), .ZN(n1137) );
NAND2_X1 U812 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NAND2_X1 U813 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XNOR2_X1 U814 ( .A(KEYINPUT26), .B(n1145), .ZN(n1143) );
XOR2_X1 U815 ( .A(KEYINPUT36), .B(n1146), .Z(n1141) );
NOR2_X1 U816 ( .A1(n1147), .A2(n1145), .ZN(n1146) );
NAND2_X1 U817 ( .A1(n1134), .A2(G472), .ZN(n1145) );
XNOR2_X1 U818 ( .A(n1144), .B(KEYINPUT42), .ZN(n1147) );
XNOR2_X1 U819 ( .A(n1148), .B(n1149), .ZN(n1144) );
NOR2_X1 U820 ( .A1(KEYINPUT21), .A2(n1150), .ZN(n1149) );
XOR2_X1 U821 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U822 ( .A(KEYINPUT23), .B(n1153), .Z(n1152) );
NOR2_X1 U823 ( .A1(n1119), .A2(n1154), .ZN(G54) );
NOR2_X1 U824 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U825 ( .A(KEYINPUT58), .B(n1157), .Z(n1156) );
NOR2_X1 U826 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XNOR2_X1 U827 ( .A(KEYINPUT50), .B(n1160), .ZN(n1159) );
NOR2_X1 U828 ( .A1(n1161), .A2(n1160), .ZN(n1155) );
NAND2_X1 U829 ( .A1(n1134), .A2(G469), .ZN(n1160) );
INV_X1 U830 ( .A(n1158), .ZN(n1161) );
XOR2_X1 U831 ( .A(n1162), .B(n1163), .Z(n1158) );
NAND2_X1 U832 ( .A1(KEYINPUT51), .A2(n1164), .ZN(n1162) );
XOR2_X1 U833 ( .A(G140), .B(n1165), .Z(n1164) );
NOR2_X1 U834 ( .A1(G110), .A2(KEYINPUT41), .ZN(n1165) );
NOR3_X1 U835 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(G51) );
AND3_X1 U836 ( .A1(KEYINPUT47), .A2(G953), .A3(G952), .ZN(n1168) );
NOR2_X1 U837 ( .A1(KEYINPUT47), .A2(n1169), .ZN(n1167) );
INV_X1 U838 ( .A(n1119), .ZN(n1169) );
NOR2_X1 U839 ( .A1(n1110), .A2(G952), .ZN(n1119) );
XOR2_X1 U840 ( .A(n1170), .B(n1171), .Z(n1166) );
XNOR2_X1 U841 ( .A(n1172), .B(n1173), .ZN(n1171) );
AND2_X1 U842 ( .A1(G210), .A2(n1134), .ZN(n1173) );
INV_X1 U843 ( .A(n1125), .ZN(n1134) );
NAND2_X1 U844 ( .A1(G902), .A2(n1024), .ZN(n1125) );
NAND2_X1 U845 ( .A1(n1111), .A2(n1083), .ZN(n1024) );
AND4_X1 U846 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1083) );
AND4_X1 U847 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1177) );
NAND2_X1 U848 ( .A1(n1182), .A2(n1034), .ZN(n1176) );
NAND2_X1 U849 ( .A1(n1183), .A2(n1184), .ZN(n1034) );
NAND2_X1 U850 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
INV_X1 U851 ( .A(n1187), .ZN(n1182) );
NAND3_X1 U852 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1174) );
NAND2_X1 U853 ( .A1(KEYINPUT22), .A2(n1191), .ZN(n1189) );
NAND2_X1 U854 ( .A1(n1192), .A2(n1193), .ZN(n1188) );
INV_X1 U855 ( .A(KEYINPUT22), .ZN(n1193) );
NAND2_X1 U856 ( .A1(n1194), .A2(n1056), .ZN(n1192) );
AND4_X1 U857 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1111) );
NOR4_X1 U858 ( .A1(n1019), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1198) );
AND3_X1 U859 ( .A1(n1058), .A2(n1202), .A3(n1055), .ZN(n1019) );
AND2_X1 U860 ( .A1(n1203), .A2(n1135), .ZN(n1197) );
NAND3_X1 U861 ( .A1(n1058), .A2(n1202), .A3(n1056), .ZN(n1135) );
NAND4_X1 U862 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1196) );
NAND2_X1 U863 ( .A1(n1208), .A2(n1031), .ZN(n1207) );
NAND2_X1 U864 ( .A1(n1185), .A2(n1209), .ZN(n1206) );
NAND2_X1 U865 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
OR2_X1 U866 ( .A1(n1211), .A2(n1212), .ZN(n1195) );
INV_X1 U867 ( .A(KEYINPUT33), .ZN(n1211) );
XNOR2_X1 U868 ( .A(KEYINPUT43), .B(n1213), .ZN(n1170) );
NOR2_X1 U869 ( .A1(KEYINPUT5), .A2(n1214), .ZN(n1213) );
XOR2_X1 U870 ( .A(n1215), .B(n1216), .Z(G48) );
XOR2_X1 U871 ( .A(n1217), .B(KEYINPUT32), .Z(n1216) );
NAND3_X1 U872 ( .A1(n1190), .A2(n1218), .A3(KEYINPUT37), .ZN(n1215) );
XOR2_X1 U873 ( .A(n1219), .B(n1175), .Z(G45) );
NAND3_X1 U874 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1175) );
NOR3_X1 U875 ( .A1(n1223), .A2(n1224), .A3(n1057), .ZN(n1222) );
XOR2_X1 U876 ( .A(n1225), .B(n1226), .Z(G42) );
XOR2_X1 U877 ( .A(KEYINPUT20), .B(G140), .Z(n1226) );
NAND3_X1 U878 ( .A1(n1035), .A2(n1227), .A3(n1228), .ZN(n1225) );
XOR2_X1 U879 ( .A(n1210), .B(KEYINPUT8), .Z(n1228) );
NAND3_X1 U880 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(G39) );
NAND2_X1 U881 ( .A1(G137), .A2(n1232), .ZN(n1231) );
NAND2_X1 U882 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
INV_X1 U883 ( .A(KEYINPUT57), .ZN(n1234) );
XNOR2_X1 U884 ( .A(KEYINPUT59), .B(n1181), .ZN(n1233) );
OR3_X1 U885 ( .A1(n1181), .A2(G137), .A3(KEYINPUT57), .ZN(n1230) );
NAND2_X1 U886 ( .A1(KEYINPUT57), .A2(n1181), .ZN(n1229) );
NAND4_X1 U887 ( .A1(n1035), .A2(n1220), .A3(n1204), .A4(n1208), .ZN(n1181) );
XNOR2_X1 U888 ( .A(G134), .B(n1180), .ZN(G36) );
NAND4_X1 U889 ( .A1(n1035), .A2(n1220), .A3(n1221), .A4(n1055), .ZN(n1180) );
NOR2_X1 U890 ( .A1(n1210), .A2(n1194), .ZN(n1220) );
INV_X1 U891 ( .A(n1235), .ZN(n1194) );
XOR2_X1 U892 ( .A(G131), .B(n1236), .Z(G33) );
NOR2_X1 U893 ( .A1(n1237), .A2(n1187), .ZN(n1236) );
NAND3_X1 U894 ( .A1(n1218), .A2(n1050), .A3(n1035), .ZN(n1187) );
NOR2_X1 U895 ( .A1(n1043), .A2(n1238), .ZN(n1035) );
AND2_X1 U896 ( .A1(G214), .A2(n1042), .ZN(n1238) );
XOR2_X1 U897 ( .A(n1183), .B(KEYINPUT9), .Z(n1237) );
INV_X1 U898 ( .A(n1221), .ZN(n1183) );
XNOR2_X1 U899 ( .A(G128), .B(n1179), .ZN(G30) );
NAND3_X1 U900 ( .A1(n1055), .A2(n1235), .A3(n1190), .ZN(n1179) );
AND4_X1 U901 ( .A1(n1050), .A2(n1038), .A3(n1208), .A4(n1186), .ZN(n1190) );
XNOR2_X1 U902 ( .A(G101), .B(n1203), .ZN(G3) );
NAND3_X1 U903 ( .A1(n1221), .A2(n1202), .A3(n1239), .ZN(n1203) );
XOR2_X1 U904 ( .A(n1240), .B(n1178), .Z(G27) );
NAND3_X1 U905 ( .A1(n1241), .A2(n1038), .A3(n1227), .ZN(n1178) );
AND3_X1 U906 ( .A1(n1185), .A2(n1186), .A3(n1218), .ZN(n1227) );
INV_X1 U907 ( .A(n1191), .ZN(n1218) );
NAND2_X1 U908 ( .A1(n1056), .A2(n1235), .ZN(n1191) );
NAND2_X1 U909 ( .A1(n1026), .A2(n1242), .ZN(n1235) );
NAND3_X1 U910 ( .A1(G902), .A2(n1243), .A3(n1086), .ZN(n1242) );
NOR2_X1 U911 ( .A1(n1110), .A2(G900), .ZN(n1086) );
XOR2_X1 U912 ( .A(G122), .B(n1201), .Z(G24) );
NOR4_X1 U913 ( .A1(n1244), .A2(n1037), .A3(n1057), .A4(n1224), .ZN(n1201) );
INV_X1 U914 ( .A(n1058), .ZN(n1037) );
NOR2_X1 U915 ( .A1(n1186), .A2(n1208), .ZN(n1058) );
XNOR2_X1 U916 ( .A(G119), .B(n1245), .ZN(G21) );
NAND4_X1 U917 ( .A1(n1204), .A2(n1205), .A3(n1246), .A4(n1208), .ZN(n1245) );
INV_X1 U918 ( .A(n1185), .ZN(n1208) );
XOR2_X1 U919 ( .A(KEYINPUT25), .B(n1241), .Z(n1246) );
XOR2_X1 U920 ( .A(G116), .B(n1200), .Z(G18) );
AND3_X1 U921 ( .A1(n1247), .A2(n1055), .A3(n1221), .ZN(n1200) );
AND2_X1 U922 ( .A1(n1248), .A2(n1249), .ZN(n1055) );
XOR2_X1 U923 ( .A(n1250), .B(KEYINPUT14), .Z(n1248) );
XOR2_X1 U924 ( .A(n1251), .B(n1199), .Z(G15) );
AND3_X1 U925 ( .A1(n1221), .A2(n1247), .A3(n1056), .ZN(n1199) );
NOR2_X1 U926 ( .A1(n1249), .A2(n1057), .ZN(n1056) );
INV_X1 U927 ( .A(n1244), .ZN(n1247) );
NAND2_X1 U928 ( .A1(n1241), .A2(n1205), .ZN(n1244) );
INV_X1 U929 ( .A(n1031), .ZN(n1241) );
NAND2_X1 U930 ( .A1(n1252), .A2(n1052), .ZN(n1031) );
NOR2_X1 U931 ( .A1(n1186), .A2(n1185), .ZN(n1221) );
XNOR2_X1 U932 ( .A(G113), .B(KEYINPUT10), .ZN(n1251) );
XOR2_X1 U933 ( .A(n1253), .B(n1212), .Z(G12) );
NAND3_X1 U934 ( .A1(n1185), .A2(n1202), .A3(n1204), .ZN(n1212) );
AND2_X1 U935 ( .A1(n1239), .A2(n1186), .ZN(n1204) );
XOR2_X1 U936 ( .A(n1254), .B(n1124), .Z(n1186) );
NAND2_X1 U937 ( .A1(G217), .A2(n1255), .ZN(n1124) );
NAND2_X1 U938 ( .A1(n1121), .A2(n1256), .ZN(n1254) );
XOR2_X1 U939 ( .A(n1257), .B(KEYINPUT3), .Z(n1121) );
XOR2_X1 U940 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U941 ( .A(n1260), .B(n1261), .Z(n1259) );
XOR2_X1 U942 ( .A(G137), .B(G128), .Z(n1261) );
XOR2_X1 U943 ( .A(KEYINPUT35), .B(G146), .Z(n1260) );
XOR2_X1 U944 ( .A(n1262), .B(n1263), .Z(n1258) );
XOR2_X1 U945 ( .A(G119), .B(n1264), .Z(n1263) );
AND3_X1 U946 ( .A1(G221), .A2(n1110), .A3(G234), .ZN(n1264) );
XNOR2_X1 U947 ( .A(n1265), .B(n1266), .ZN(n1262) );
NAND2_X1 U948 ( .A1(KEYINPUT39), .A2(n1253), .ZN(n1266) );
NAND2_X1 U949 ( .A1(KEYINPUT40), .A2(n1267), .ZN(n1265) );
INV_X1 U950 ( .A(n1029), .ZN(n1239) );
NAND2_X1 U951 ( .A1(n1224), .A2(n1250), .ZN(n1029) );
XOR2_X1 U952 ( .A(n1057), .B(KEYINPUT12), .Z(n1250) );
XOR2_X1 U953 ( .A(n1268), .B(G475), .Z(n1057) );
NAND2_X1 U954 ( .A1(n1256), .A2(n1132), .ZN(n1268) );
NAND2_X1 U955 ( .A1(n1269), .A2(n1270), .ZN(n1132) );
NAND2_X1 U956 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XOR2_X1 U957 ( .A(n1273), .B(KEYINPUT34), .Z(n1269) );
OR2_X1 U958 ( .A1(n1272), .A2(n1271), .ZN(n1273) );
XOR2_X1 U959 ( .A(n1274), .B(G104), .Z(n1271) );
NAND2_X1 U960 ( .A1(n1275), .A2(KEYINPUT2), .ZN(n1274) );
XNOR2_X1 U961 ( .A(G113), .B(n1276), .ZN(n1275) );
XOR2_X1 U962 ( .A(KEYINPUT61), .B(G122), .Z(n1276) );
XNOR2_X1 U963 ( .A(n1277), .B(n1278), .ZN(n1272) );
XOR2_X1 U964 ( .A(n1279), .B(n1280), .Z(n1278) );
NAND2_X1 U965 ( .A1(G214), .A2(n1281), .ZN(n1280) );
NAND2_X1 U966 ( .A1(n1282), .A2(n1283), .ZN(n1279) );
NAND2_X1 U967 ( .A1(n1267), .A2(n1217), .ZN(n1283) );
XOR2_X1 U968 ( .A(KEYINPUT38), .B(n1284), .Z(n1282) );
NOR2_X1 U969 ( .A1(n1267), .A2(n1217), .ZN(n1284) );
INV_X1 U970 ( .A(G146), .ZN(n1217) );
XOR2_X1 U971 ( .A(n1240), .B(G140), .Z(n1267) );
INV_X1 U972 ( .A(G125), .ZN(n1240) );
XOR2_X1 U973 ( .A(G131), .B(n1219), .Z(n1277) );
INV_X1 U974 ( .A(G143), .ZN(n1219) );
INV_X1 U975 ( .A(n1249), .ZN(n1224) );
NAND2_X1 U976 ( .A1(n1285), .A2(n1068), .ZN(n1249) );
NAND2_X1 U977 ( .A1(n1076), .A2(n1078), .ZN(n1068) );
OR2_X1 U978 ( .A1(n1078), .A2(n1076), .ZN(n1285) );
NOR2_X1 U979 ( .A1(n1127), .A2(G902), .ZN(n1076) );
XNOR2_X1 U980 ( .A(n1286), .B(n1287), .ZN(n1127) );
NOR2_X1 U981 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
XOR2_X1 U982 ( .A(n1290), .B(KEYINPUT55), .Z(n1289) );
NAND2_X1 U983 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
NOR2_X1 U984 ( .A1(n1291), .A2(n1292), .ZN(n1288) );
XOR2_X1 U985 ( .A(G128), .B(n1293), .Z(n1292) );
XOR2_X1 U986 ( .A(G143), .B(G134), .Z(n1293) );
XOR2_X1 U987 ( .A(n1294), .B(n1295), .Z(n1291) );
XOR2_X1 U988 ( .A(G122), .B(G116), .Z(n1295) );
NAND3_X1 U989 ( .A1(G217), .A2(n1110), .A3(G234), .ZN(n1286) );
INV_X1 U990 ( .A(G478), .ZN(n1078) );
AND2_X1 U991 ( .A1(n1050), .A2(n1205), .ZN(n1202) );
AND2_X1 U992 ( .A1(n1038), .A2(n1296), .ZN(n1205) );
NAND2_X1 U993 ( .A1(n1026), .A2(n1297), .ZN(n1296) );
NAND3_X1 U994 ( .A1(n1113), .A2(n1243), .A3(G902), .ZN(n1297) );
NOR2_X1 U995 ( .A1(G898), .A2(n1110), .ZN(n1113) );
NAND3_X1 U996 ( .A1(n1243), .A2(n1110), .A3(G952), .ZN(n1026) );
NAND2_X1 U997 ( .A1(G237), .A2(G234), .ZN(n1243) );
INV_X1 U998 ( .A(n1223), .ZN(n1038) );
NAND2_X1 U999 ( .A1(n1298), .A2(n1043), .ZN(n1223) );
NAND2_X1 U1000 ( .A1(n1299), .A2(n1074), .ZN(n1043) );
NAND3_X1 U1001 ( .A1(n1042), .A2(n1300), .A3(G210), .ZN(n1074) );
NAND2_X1 U1002 ( .A1(n1301), .A2(n1302), .ZN(n1299) );
NAND2_X1 U1003 ( .A1(G210), .A2(n1042), .ZN(n1302) );
INV_X1 U1004 ( .A(n1300), .ZN(n1301) );
NAND3_X1 U1005 ( .A1(n1303), .A2(n1256), .A3(n1304), .ZN(n1300) );
XOR2_X1 U1006 ( .A(KEYINPUT0), .B(n1305), .Z(n1304) );
NOR2_X1 U1007 ( .A1(n1214), .A2(n1172), .ZN(n1305) );
NAND2_X1 U1008 ( .A1(n1214), .A2(n1172), .ZN(n1303) );
XNOR2_X1 U1009 ( .A(n1306), .B(n1307), .ZN(n1172) );
XOR2_X1 U1010 ( .A(KEYINPUT6), .B(G125), .Z(n1307) );
XOR2_X1 U1011 ( .A(n1308), .B(n1309), .Z(n1306) );
AND2_X1 U1012 ( .A1(n1110), .A2(G224), .ZN(n1309) );
XNOR2_X1 U1013 ( .A(n1310), .B(n1116), .ZN(n1214) );
XNOR2_X1 U1014 ( .A(n1311), .B(G101), .ZN(n1116) );
NAND2_X1 U1015 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NAND2_X1 U1016 ( .A1(G104), .A2(n1294), .ZN(n1313) );
XOR2_X1 U1017 ( .A(KEYINPUT30), .B(n1314), .Z(n1312) );
NOR2_X1 U1018 ( .A1(G104), .A2(n1294), .ZN(n1314) );
INV_X1 U1019 ( .A(G107), .ZN(n1294) );
XOR2_X1 U1020 ( .A(n1315), .B(n1118), .Z(n1310) );
INV_X1 U1021 ( .A(n1148), .ZN(n1118) );
NAND2_X1 U1022 ( .A1(KEYINPUT49), .A2(n1115), .ZN(n1315) );
XOR2_X1 U1023 ( .A(G122), .B(n1316), .Z(n1115) );
NOR2_X1 U1024 ( .A1(KEYINPUT13), .A2(n1253), .ZN(n1316) );
NAND2_X1 U1025 ( .A1(G214), .A2(n1042), .ZN(n1298) );
NAND2_X1 U1026 ( .A1(n1317), .A2(n1256), .ZN(n1042) );
XOR2_X1 U1027 ( .A(KEYINPUT46), .B(G237), .Z(n1317) );
INV_X1 U1028 ( .A(n1210), .ZN(n1050) );
NAND2_X1 U1029 ( .A1(n1052), .A2(n1053), .ZN(n1210) );
INV_X1 U1030 ( .A(n1252), .ZN(n1053) );
NOR2_X1 U1031 ( .A1(n1318), .A2(n1062), .ZN(n1252) );
NOR2_X1 U1032 ( .A1(n1067), .A2(G469), .ZN(n1062) );
AND2_X1 U1033 ( .A1(G469), .A2(n1067), .ZN(n1318) );
NAND2_X1 U1034 ( .A1(n1319), .A2(n1256), .ZN(n1067) );
XOR2_X1 U1035 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1036 ( .A(KEYINPUT24), .B(G140), .Z(n1321) );
XOR2_X1 U1037 ( .A(n1163), .B(n1253), .Z(n1320) );
XNOR2_X1 U1038 ( .A(n1322), .B(n1323), .ZN(n1163) );
XOR2_X1 U1039 ( .A(G104), .B(n1324), .Z(n1323) );
XOR2_X1 U1040 ( .A(KEYINPUT62), .B(G107), .Z(n1324) );
XOR2_X1 U1041 ( .A(n1325), .B(n1326), .Z(n1322) );
XOR2_X1 U1042 ( .A(n1092), .B(n1327), .Z(n1325) );
AND2_X1 U1043 ( .A1(n1110), .A2(G227), .ZN(n1327) );
INV_X1 U1044 ( .A(G953), .ZN(n1110) );
NAND2_X1 U1045 ( .A1(n1328), .A2(n1329), .ZN(n1092) );
NAND2_X1 U1046 ( .A1(G128), .A2(n1330), .ZN(n1329) );
XOR2_X1 U1047 ( .A(KEYINPUT44), .B(n1331), .Z(n1328) );
NOR2_X1 U1048 ( .A1(G128), .A2(n1330), .ZN(n1331) );
NAND2_X1 U1049 ( .A1(G221), .A2(n1255), .ZN(n1052) );
NAND2_X1 U1050 ( .A1(G234), .A2(n1256), .ZN(n1255) );
XOR2_X1 U1051 ( .A(n1332), .B(G472), .Z(n1185) );
NAND2_X1 U1052 ( .A1(n1333), .A2(n1256), .ZN(n1332) );
INV_X1 U1053 ( .A(G902), .ZN(n1256) );
XOR2_X1 U1054 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1055 ( .A(n1139), .B(n1336), .Z(n1335) );
XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n1336) );
NAND2_X1 U1057 ( .A1(G210), .A2(n1281), .ZN(n1139) );
NOR2_X1 U1058 ( .A1(G953), .A2(G237), .ZN(n1281) );
XOR2_X1 U1059 ( .A(n1337), .B(n1338), .Z(n1334) );
INV_X1 U1060 ( .A(n1151), .ZN(n1338) );
XOR2_X1 U1061 ( .A(n1308), .B(KEYINPUT15), .Z(n1151) );
XNOR2_X1 U1062 ( .A(G128), .B(n1330), .ZN(n1308) );
XOR2_X1 U1063 ( .A(G143), .B(G146), .Z(n1330) );
XOR2_X1 U1064 ( .A(n1326), .B(n1148), .Z(n1337) );
XNOR2_X1 U1065 ( .A(G113), .B(n1339), .ZN(n1148) );
XOR2_X1 U1066 ( .A(G119), .B(G116), .Z(n1339) );
XOR2_X1 U1067 ( .A(n1153), .B(G101), .Z(n1326) );
XOR2_X1 U1068 ( .A(G137), .B(n1090), .Z(n1153) );
XOR2_X1 U1069 ( .A(G131), .B(G134), .Z(n1090) );
INV_X1 U1070 ( .A(G110), .ZN(n1253) );
endmodule


