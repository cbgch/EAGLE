//Key = 0111111010010111000110100010110110011100100010101101010101101101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460;

XNOR2_X1 U810 ( .A(n1123), .B(n1124), .ZN(G9) );
NOR2_X1 U811 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR2_X1 U812 ( .A1(n1127), .A2(n1128), .ZN(G75) );
NOR3_X1 U813 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1128) );
NAND3_X1 U814 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1129) );
NAND3_X1 U815 ( .A1(n1135), .A2(n1136), .A3(KEYINPUT13), .ZN(n1134) );
NAND2_X1 U816 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
NAND3_X1 U817 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1138) );
NAND3_X1 U818 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1140) );
NAND2_X1 U819 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U820 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
XNOR2_X1 U821 ( .A(n1145), .B(KEYINPUT4), .ZN(n1147) );
NAND2_X1 U822 ( .A1(n1149), .A2(n1150), .ZN(n1142) );
NAND2_X1 U823 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NAND2_X1 U824 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND3_X1 U825 ( .A1(n1149), .A2(n1155), .A3(n1145), .ZN(n1137) );
NAND3_X1 U826 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1155) );
NAND2_X1 U827 ( .A1(n1141), .A2(n1159), .ZN(n1158) );
NAND2_X1 U828 ( .A1(n1126), .A2(n1160), .ZN(n1159) );
NAND2_X1 U829 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U830 ( .A1(n1163), .A2(n1164), .ZN(n1156) );
XNOR2_X1 U831 ( .A(n1139), .B(KEYINPUT28), .ZN(n1163) );
AND3_X1 U832 ( .A1(n1132), .A2(n1133), .A3(n1165), .ZN(n1127) );
NAND4_X1 U833 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1132) );
NOR3_X1 U834 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1169) );
XNOR2_X1 U835 ( .A(n1173), .B(KEYINPUT2), .ZN(n1171) );
NAND3_X1 U836 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1170) );
NAND2_X1 U837 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
INV_X1 U838 ( .A(KEYINPUT12), .ZN(n1178) );
NAND2_X1 U839 ( .A1(KEYINPUT12), .A2(n1179), .ZN(n1174) );
NOR3_X1 U840 ( .A1(n1153), .A2(n1162), .A3(n1180), .ZN(n1168) );
XNOR2_X1 U841 ( .A(n1181), .B(n1182), .ZN(n1167) );
NOR2_X1 U842 ( .A1(G469), .A2(KEYINPUT45), .ZN(n1182) );
XNOR2_X1 U843 ( .A(KEYINPUT49), .B(n1183), .ZN(n1166) );
XOR2_X1 U844 ( .A(n1184), .B(n1185), .Z(G72) );
XOR2_X1 U845 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U846 ( .A1(n1188), .A2(n1133), .ZN(n1187) );
AND2_X1 U847 ( .A1(G227), .A2(G900), .ZN(n1188) );
NAND2_X1 U848 ( .A1(n1189), .A2(n1190), .ZN(n1186) );
NAND2_X1 U849 ( .A1(G953), .A2(n1191), .ZN(n1190) );
XOR2_X1 U850 ( .A(n1192), .B(n1193), .Z(n1189) );
XOR2_X1 U851 ( .A(n1194), .B(n1195), .Z(n1193) );
XNOR2_X1 U852 ( .A(n1196), .B(n1197), .ZN(n1195) );
NOR2_X1 U853 ( .A1(G125), .A2(KEYINPUT7), .ZN(n1197) );
NOR2_X1 U854 ( .A1(KEYINPUT62), .A2(n1198), .ZN(n1196) );
XOR2_X1 U855 ( .A(n1199), .B(n1200), .Z(n1192) );
XNOR2_X1 U856 ( .A(KEYINPUT8), .B(n1201), .ZN(n1200) );
NOR2_X1 U857 ( .A1(KEYINPUT18), .A2(n1202), .ZN(n1199) );
NAND2_X1 U858 ( .A1(n1133), .A2(n1131), .ZN(n1184) );
NAND2_X1 U859 ( .A1(n1203), .A2(n1204), .ZN(G69) );
NAND2_X1 U860 ( .A1(n1205), .A2(n1133), .ZN(n1204) );
XNOR2_X1 U861 ( .A(n1130), .B(n1206), .ZN(n1205) );
NAND2_X1 U862 ( .A1(n1207), .A2(G953), .ZN(n1203) );
NAND2_X1 U863 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U864 ( .A1(n1206), .A2(n1210), .ZN(n1209) );
NAND2_X1 U865 ( .A1(G224), .A2(n1211), .ZN(n1208) );
NAND2_X1 U866 ( .A1(G898), .A2(n1206), .ZN(n1211) );
NAND4_X1 U867 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1206) );
NAND3_X1 U868 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
NAND3_X1 U869 ( .A1(KEYINPUT5), .A2(n1219), .A3(n1220), .ZN(n1214) );
NAND2_X1 U870 ( .A1(G953), .A2(n1221), .ZN(n1213) );
NAND3_X1 U871 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1212) );
INV_X1 U872 ( .A(n1217), .ZN(n1224) );
NAND2_X1 U873 ( .A1(n1220), .A2(KEYINPUT5), .ZN(n1223) );
NAND2_X1 U874 ( .A1(n1218), .A2(n1216), .ZN(n1222) );
NAND2_X1 U875 ( .A1(KEYINPUT5), .A2(n1225), .ZN(n1216) );
INV_X1 U876 ( .A(n1220), .ZN(n1218) );
NOR3_X1 U877 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(G66) );
AND2_X1 U878 ( .A1(KEYINPUT51), .A2(n1229), .ZN(n1228) );
NOR3_X1 U879 ( .A1(KEYINPUT51), .A2(n1133), .A3(n1165), .ZN(n1227) );
INV_X1 U880 ( .A(G952), .ZN(n1165) );
XOR2_X1 U881 ( .A(n1230), .B(n1231), .Z(n1226) );
NAND3_X1 U882 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1230) );
NAND2_X1 U883 ( .A1(KEYINPUT48), .A2(n1235), .ZN(n1233) );
NAND2_X1 U884 ( .A1(n1236), .A2(n1237), .ZN(n1232) );
INV_X1 U885 ( .A(KEYINPUT48), .ZN(n1237) );
NAND3_X1 U886 ( .A1(n1238), .A2(G902), .A3(n1239), .ZN(n1236) );
NOR3_X1 U887 ( .A1(n1240), .A2(n1229), .A3(n1241), .ZN(G63) );
NOR4_X1 U888 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1235), .ZN(n1241) );
NOR2_X1 U889 ( .A1(KEYINPUT29), .A2(n1245), .ZN(n1243) );
NOR2_X1 U890 ( .A1(n1246), .A2(n1247), .ZN(n1242) );
INV_X1 U891 ( .A(KEYINPUT29), .ZN(n1247) );
NOR2_X1 U892 ( .A1(n1248), .A2(n1246), .ZN(n1240) );
NOR2_X1 U893 ( .A1(KEYINPUT52), .A2(n1245), .ZN(n1246) );
NOR2_X1 U894 ( .A1(n1244), .A2(n1235), .ZN(n1248) );
INV_X1 U895 ( .A(G478), .ZN(n1244) );
NOR2_X1 U896 ( .A1(n1229), .A2(n1249), .ZN(G60) );
XNOR2_X1 U897 ( .A(n1250), .B(n1251), .ZN(n1249) );
NOR2_X1 U898 ( .A1(n1252), .A2(n1235), .ZN(n1251) );
XNOR2_X1 U899 ( .A(G104), .B(n1253), .ZN(G6) );
NAND2_X1 U900 ( .A1(KEYINPUT44), .A2(n1254), .ZN(n1253) );
NOR2_X1 U901 ( .A1(n1229), .A2(n1255), .ZN(G57) );
XOR2_X1 U902 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U903 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U904 ( .A(n1260), .B(n1261), .Z(n1256) );
NOR2_X1 U905 ( .A1(n1262), .A2(n1235), .ZN(n1261) );
NAND2_X1 U906 ( .A1(KEYINPUT36), .A2(n1263), .ZN(n1260) );
NOR2_X1 U907 ( .A1(n1229), .A2(n1264), .ZN(G54) );
NOR2_X1 U908 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
XOR2_X1 U909 ( .A(n1267), .B(KEYINPUT63), .Z(n1266) );
NAND2_X1 U910 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NOR2_X1 U911 ( .A1(n1268), .A2(n1269), .ZN(n1265) );
XNOR2_X1 U912 ( .A(n1270), .B(n1271), .ZN(n1269) );
XNOR2_X1 U913 ( .A(n1201), .B(G110), .ZN(n1271) );
XNOR2_X1 U914 ( .A(n1272), .B(n1273), .ZN(n1270) );
NAND2_X1 U915 ( .A1(KEYINPUT46), .A2(n1274), .ZN(n1272) );
NOR2_X1 U916 ( .A1(n1235), .A2(n1275), .ZN(n1268) );
INV_X1 U917 ( .A(G469), .ZN(n1275) );
NOR2_X1 U918 ( .A1(n1229), .A2(n1276), .ZN(G51) );
NOR2_X1 U919 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
XOR2_X1 U920 ( .A(KEYINPUT16), .B(n1279), .Z(n1278) );
NOR3_X1 U921 ( .A1(n1235), .A2(n1280), .A3(n1281), .ZN(n1279) );
XNOR2_X1 U922 ( .A(n1282), .B(KEYINPUT39), .ZN(n1280) );
NOR2_X1 U923 ( .A1(n1283), .A2(n1282), .ZN(n1277) );
XOR2_X1 U924 ( .A(n1284), .B(n1285), .Z(n1282) );
NOR2_X1 U925 ( .A1(KEYINPUT0), .A2(n1286), .ZN(n1285) );
NOR2_X1 U926 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XOR2_X1 U927 ( .A(n1289), .B(KEYINPUT57), .Z(n1288) );
NAND2_X1 U928 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NOR2_X1 U929 ( .A1(n1290), .A2(n1291), .ZN(n1287) );
NOR2_X1 U930 ( .A1(n1281), .A2(n1235), .ZN(n1283) );
NAND2_X1 U931 ( .A1(G902), .A2(n1292), .ZN(n1235) );
NAND2_X1 U932 ( .A1(n1239), .A2(n1238), .ZN(n1292) );
INV_X1 U933 ( .A(n1130), .ZN(n1238) );
NAND4_X1 U934 ( .A1(n1293), .A2(n1294), .A3(n1295), .A4(n1296), .ZN(n1130) );
NOR4_X1 U935 ( .A1(n1297), .A2(n1298), .A3(n1299), .A4(n1254), .ZN(n1296) );
AND3_X1 U936 ( .A1(n1300), .A2(n1149), .A3(n1301), .ZN(n1254) );
NOR2_X1 U937 ( .A1(n1302), .A2(n1303), .ZN(n1295) );
NOR2_X1 U938 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NOR2_X1 U939 ( .A1(n1306), .A2(n1307), .ZN(n1304) );
NOR2_X1 U940 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
XNOR2_X1 U941 ( .A(KEYINPUT19), .B(n1310), .ZN(n1309) );
AND3_X1 U942 ( .A1(KEYINPUT31), .A2(n1146), .A3(n1300), .ZN(n1306) );
INV_X1 U943 ( .A(n1311), .ZN(n1302) );
NAND2_X1 U944 ( .A1(n1312), .A2(n1313), .ZN(n1294) );
XOR2_X1 U945 ( .A(n1125), .B(KEYINPUT58), .Z(n1312) );
NAND4_X1 U946 ( .A1(n1149), .A2(n1164), .A3(n1314), .A4(n1315), .ZN(n1125) );
NAND4_X1 U947 ( .A1(n1145), .A2(n1300), .A3(n1316), .A4(n1126), .ZN(n1293) );
AND3_X1 U948 ( .A1(n1146), .A2(n1317), .A3(n1315), .ZN(n1316) );
INV_X1 U949 ( .A(KEYINPUT31), .ZN(n1317) );
XOR2_X1 U950 ( .A(n1131), .B(KEYINPUT14), .Z(n1239) );
NAND4_X1 U951 ( .A1(n1318), .A2(n1319), .A3(n1320), .A4(n1321), .ZN(n1131) );
NOR4_X1 U952 ( .A1(n1322), .A2(n1323), .A3(n1324), .A4(n1325), .ZN(n1321) );
NOR2_X1 U953 ( .A1(n1326), .A2(n1327), .ZN(n1320) );
NOR2_X1 U954 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NOR2_X1 U955 ( .A1(n1330), .A2(n1331), .ZN(n1326) );
XOR2_X1 U956 ( .A(n1332), .B(KEYINPUT21), .Z(n1330) );
NAND4_X1 U957 ( .A1(n1164), .A2(n1333), .A3(n1146), .A4(n1334), .ZN(n1332) );
XNOR2_X1 U958 ( .A(KEYINPUT30), .B(n1151), .ZN(n1333) );
INV_X1 U959 ( .A(n1335), .ZN(n1151) );
NAND3_X1 U960 ( .A1(n1336), .A2(n1313), .A3(n1337), .ZN(n1318) );
NOR2_X1 U961 ( .A1(n1133), .A2(G952), .ZN(n1229) );
XOR2_X1 U962 ( .A(G146), .B(n1338), .Z(G48) );
NOR3_X1 U963 ( .A1(n1329), .A2(KEYINPUT23), .A3(n1328), .ZN(n1338) );
NAND3_X1 U964 ( .A1(n1313), .A2(n1335), .A3(n1300), .ZN(n1329) );
XNOR2_X1 U965 ( .A(n1339), .B(n1340), .ZN(G45) );
NOR3_X1 U966 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1340) );
XNOR2_X1 U967 ( .A(n1337), .B(KEYINPUT59), .ZN(n1342) );
XNOR2_X1 U968 ( .A(KEYINPUT3), .B(n1126), .ZN(n1341) );
INV_X1 U969 ( .A(n1313), .ZN(n1126) );
NAND2_X1 U970 ( .A1(n1344), .A2(n1345), .ZN(G42) );
NAND2_X1 U971 ( .A1(n1346), .A2(n1201), .ZN(n1345) );
XOR2_X1 U972 ( .A(KEYINPUT33), .B(n1324), .Z(n1346) );
NAND2_X1 U973 ( .A1(n1347), .A2(G140), .ZN(n1344) );
XOR2_X1 U974 ( .A(KEYINPUT32), .B(n1324), .Z(n1347) );
AND4_X1 U975 ( .A1(n1348), .A2(n1148), .A3(n1335), .A4(n1334), .ZN(n1324) );
INV_X1 U976 ( .A(n1157), .ZN(n1348) );
XNOR2_X1 U977 ( .A(G137), .B(n1319), .ZN(G39) );
NAND4_X1 U978 ( .A1(n1141), .A2(n1349), .A3(n1139), .A4(n1335), .ZN(n1319) );
XOR2_X1 U979 ( .A(G134), .B(n1350), .Z(G36) );
AND3_X1 U980 ( .A1(n1336), .A2(n1164), .A3(n1139), .ZN(n1350) );
INV_X1 U981 ( .A(n1343), .ZN(n1336) );
XNOR2_X1 U982 ( .A(n1198), .B(n1323), .ZN(G33) );
NOR2_X1 U983 ( .A1(n1157), .A2(n1343), .ZN(n1323) );
NAND3_X1 U984 ( .A1(n1146), .A2(n1334), .A3(n1335), .ZN(n1343) );
NAND2_X1 U985 ( .A1(n1139), .A2(n1300), .ZN(n1157) );
INV_X1 U986 ( .A(n1331), .ZN(n1139) );
NAND2_X1 U987 ( .A1(n1161), .A2(n1351), .ZN(n1331) );
XOR2_X1 U988 ( .A(KEYINPUT60), .B(n1162), .Z(n1351) );
XOR2_X1 U989 ( .A(G128), .B(n1325), .Z(G30) );
AND4_X1 U990 ( .A1(n1349), .A2(n1313), .A3(n1314), .A4(n1164), .ZN(n1325) );
INV_X1 U991 ( .A(n1328), .ZN(n1349) );
NAND3_X1 U992 ( .A1(n1172), .A2(n1334), .A3(n1173), .ZN(n1328) );
XNOR2_X1 U993 ( .A(n1299), .B(n1352), .ZN(G3) );
NAND2_X1 U994 ( .A1(KEYINPUT11), .A2(G101), .ZN(n1352) );
AND3_X1 U995 ( .A1(n1141), .A2(n1146), .A3(n1301), .ZN(n1299) );
XOR2_X1 U996 ( .A(G125), .B(n1322), .Z(G27) );
AND4_X1 U997 ( .A1(n1148), .A2(n1145), .A3(n1353), .A4(n1300), .ZN(n1322) );
AND2_X1 U998 ( .A1(n1334), .A2(n1313), .ZN(n1353) );
NAND2_X1 U999 ( .A1(n1354), .A2(n1355), .ZN(n1334) );
NAND2_X1 U1000 ( .A1(n1356), .A2(n1191), .ZN(n1355) );
INV_X1 U1001 ( .A(G900), .ZN(n1191) );
XOR2_X1 U1002 ( .A(n1357), .B(n1358), .Z(G24) );
NOR3_X1 U1003 ( .A1(n1305), .A2(n1308), .A3(n1310), .ZN(n1358) );
INV_X1 U1004 ( .A(n1337), .ZN(n1310) );
NOR2_X1 U1005 ( .A1(n1183), .A2(n1176), .ZN(n1337) );
INV_X1 U1006 ( .A(n1149), .ZN(n1308) );
NOR2_X1 U1007 ( .A1(KEYINPUT10), .A2(n1359), .ZN(n1357) );
INV_X1 U1008 ( .A(G122), .ZN(n1359) );
XNOR2_X1 U1009 ( .A(G119), .B(n1311), .ZN(G21) );
NAND4_X1 U1010 ( .A1(n1360), .A2(n1141), .A3(n1173), .A4(n1172), .ZN(n1311) );
XOR2_X1 U1011 ( .A(G116), .B(n1298), .Z(G18) );
AND3_X1 U1012 ( .A1(n1164), .A2(n1146), .A3(n1360), .ZN(n1298) );
NOR2_X1 U1013 ( .A1(n1361), .A2(n1176), .ZN(n1164) );
XNOR2_X1 U1014 ( .A(G113), .B(n1362), .ZN(G15) );
NAND4_X1 U1015 ( .A1(KEYINPUT1), .A2(n1360), .A3(n1300), .A4(n1146), .ZN(n1362) );
NAND2_X1 U1016 ( .A1(n1363), .A2(n1364), .ZN(n1146) );
NAND3_X1 U1017 ( .A1(n1173), .A2(n1365), .A3(n1366), .ZN(n1364) );
INV_X1 U1018 ( .A(KEYINPUT50), .ZN(n1366) );
NAND2_X1 U1019 ( .A1(KEYINPUT50), .A2(n1149), .ZN(n1363) );
NOR2_X1 U1020 ( .A1(n1172), .A2(n1173), .ZN(n1149) );
AND2_X1 U1021 ( .A1(n1176), .A2(n1361), .ZN(n1300) );
INV_X1 U1022 ( .A(n1305), .ZN(n1360) );
NAND3_X1 U1023 ( .A1(n1313), .A2(n1315), .A3(n1145), .ZN(n1305) );
NOR2_X1 U1024 ( .A1(n1367), .A2(n1153), .ZN(n1145) );
INV_X1 U1025 ( .A(n1154), .ZN(n1367) );
XNOR2_X1 U1026 ( .A(n1368), .B(n1297), .ZN(G12) );
AND3_X1 U1027 ( .A1(n1141), .A2(n1148), .A3(n1301), .ZN(n1297) );
AND3_X1 U1028 ( .A1(n1314), .A2(n1315), .A3(n1313), .ZN(n1301) );
NOR2_X1 U1029 ( .A1(n1161), .A2(n1162), .ZN(n1313) );
AND2_X1 U1030 ( .A1(G214), .A2(n1369), .ZN(n1162) );
NOR2_X1 U1031 ( .A1(n1180), .A2(n1177), .ZN(n1161) );
NOR2_X1 U1032 ( .A1(n1281), .A2(n1179), .ZN(n1177) );
AND2_X1 U1033 ( .A1(n1179), .A2(n1281), .ZN(n1180) );
NAND2_X1 U1034 ( .A1(G210), .A2(n1369), .ZN(n1281) );
OR2_X1 U1035 ( .A1(G902), .A2(G237), .ZN(n1369) );
AND2_X1 U1036 ( .A1(n1370), .A2(n1371), .ZN(n1179) );
XNOR2_X1 U1037 ( .A(n1372), .B(n1373), .ZN(n1370) );
INV_X1 U1038 ( .A(n1284), .ZN(n1373) );
XOR2_X1 U1039 ( .A(n1220), .B(n1219), .Z(n1284) );
XNOR2_X1 U1040 ( .A(n1217), .B(n1225), .ZN(n1219) );
XNOR2_X1 U1041 ( .A(n1374), .B(n1375), .ZN(n1225) );
NAND2_X1 U1042 ( .A1(n1376), .A2(n1377), .ZN(n1217) );
NAND2_X1 U1043 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
XOR2_X1 U1044 ( .A(KEYINPUT53), .B(n1380), .Z(n1376) );
NOR2_X1 U1045 ( .A1(n1378), .A2(n1379), .ZN(n1380) );
XNOR2_X1 U1046 ( .A(G104), .B(n1381), .ZN(n1378) );
NOR2_X1 U1047 ( .A1(KEYINPUT34), .A2(n1123), .ZN(n1381) );
INV_X1 U1048 ( .A(G107), .ZN(n1123) );
XOR2_X1 U1049 ( .A(G110), .B(n1382), .Z(n1220) );
NOR2_X1 U1050 ( .A1(n1383), .A2(n1384), .ZN(n1372) );
NOR3_X1 U1051 ( .A1(n1385), .A2(KEYINPUT43), .A3(n1210), .ZN(n1384) );
INV_X1 U1052 ( .A(n1291), .ZN(n1385) );
NOR2_X1 U1053 ( .A1(n1386), .A2(n1291), .ZN(n1383) );
XOR2_X1 U1054 ( .A(G125), .B(n1387), .Z(n1291) );
NOR2_X1 U1055 ( .A1(KEYINPUT43), .A2(n1388), .ZN(n1386) );
INV_X1 U1056 ( .A(n1290), .ZN(n1388) );
NOR2_X1 U1057 ( .A1(n1210), .A2(G953), .ZN(n1290) );
INV_X1 U1058 ( .A(G224), .ZN(n1210) );
NAND2_X1 U1059 ( .A1(n1354), .A2(n1389), .ZN(n1315) );
NAND2_X1 U1060 ( .A1(n1356), .A2(n1221), .ZN(n1389) );
INV_X1 U1061 ( .A(G898), .ZN(n1221) );
AND3_X1 U1062 ( .A1(G902), .A2(n1136), .A3(G953), .ZN(n1356) );
NAND3_X1 U1063 ( .A1(n1136), .A2(n1133), .A3(G952), .ZN(n1354) );
NAND2_X1 U1064 ( .A1(G237), .A2(G234), .ZN(n1136) );
XNOR2_X1 U1065 ( .A(n1335), .B(KEYINPUT6), .ZN(n1314) );
NOR2_X1 U1066 ( .A1(n1154), .A2(n1153), .ZN(n1335) );
AND2_X1 U1067 ( .A1(G221), .A2(n1390), .ZN(n1153) );
XOR2_X1 U1068 ( .A(n1181), .B(G469), .Z(n1154) );
NAND2_X1 U1069 ( .A1(n1391), .A2(n1371), .ZN(n1181) );
XOR2_X1 U1070 ( .A(n1392), .B(n1393), .Z(n1391) );
XNOR2_X1 U1071 ( .A(G140), .B(n1394), .ZN(n1393) );
NAND2_X1 U1072 ( .A1(KEYINPUT55), .A2(n1368), .ZN(n1394) );
XOR2_X1 U1073 ( .A(n1274), .B(n1395), .Z(n1392) );
NOR2_X1 U1074 ( .A1(KEYINPUT24), .A2(n1273), .ZN(n1395) );
NAND2_X1 U1075 ( .A1(G227), .A2(n1133), .ZN(n1273) );
XOR2_X1 U1076 ( .A(n1396), .B(n1397), .Z(n1274) );
XOR2_X1 U1077 ( .A(n1398), .B(n1399), .Z(n1397) );
XNOR2_X1 U1078 ( .A(G104), .B(n1379), .ZN(n1399) );
NOR2_X1 U1079 ( .A1(G107), .A2(KEYINPUT56), .ZN(n1398) );
XOR2_X1 U1080 ( .A(n1194), .B(n1400), .Z(n1396) );
XOR2_X1 U1081 ( .A(n1401), .B(n1402), .Z(n1194) );
XOR2_X1 U1082 ( .A(n1403), .B(G134), .Z(n1401) );
NAND2_X1 U1083 ( .A1(KEYINPUT37), .A2(n1339), .ZN(n1403) );
NOR2_X1 U1084 ( .A1(n1173), .A2(n1365), .ZN(n1148) );
INV_X1 U1085 ( .A(n1172), .ZN(n1365) );
XNOR2_X1 U1086 ( .A(n1404), .B(n1234), .ZN(n1172) );
AND2_X1 U1087 ( .A1(G217), .A2(n1390), .ZN(n1234) );
NAND2_X1 U1088 ( .A1(G234), .A2(n1371), .ZN(n1390) );
NAND2_X1 U1089 ( .A1(n1231), .A2(n1371), .ZN(n1404) );
XOR2_X1 U1090 ( .A(n1405), .B(n1406), .Z(n1231) );
XOR2_X1 U1091 ( .A(n1407), .B(n1408), .Z(n1406) );
NAND3_X1 U1092 ( .A1(n1409), .A2(n1410), .A3(n1411), .ZN(n1408) );
NAND2_X1 U1093 ( .A1(G110), .A2(n1412), .ZN(n1411) );
NAND2_X1 U1094 ( .A1(n1413), .A2(n1414), .ZN(n1410) );
INV_X1 U1095 ( .A(KEYINPUT26), .ZN(n1414) );
NAND2_X1 U1096 ( .A1(n1415), .A2(n1416), .ZN(n1413) );
INV_X1 U1097 ( .A(n1412), .ZN(n1416) );
XNOR2_X1 U1098 ( .A(KEYINPUT47), .B(G110), .ZN(n1415) );
NAND2_X1 U1099 ( .A1(KEYINPUT26), .A2(n1417), .ZN(n1409) );
NAND2_X1 U1100 ( .A1(n1418), .A2(n1419), .ZN(n1417) );
OR3_X1 U1101 ( .A1(n1412), .A2(G110), .A3(KEYINPUT47), .ZN(n1419) );
XOR2_X1 U1102 ( .A(G119), .B(G128), .Z(n1412) );
NAND2_X1 U1103 ( .A1(KEYINPUT47), .A2(G110), .ZN(n1418) );
NAND2_X1 U1104 ( .A1(KEYINPUT40), .A2(n1420), .ZN(n1407) );
XOR2_X1 U1105 ( .A(n1421), .B(n1422), .Z(n1420) );
NOR2_X1 U1106 ( .A1(G146), .A2(KEYINPUT27), .ZN(n1421) );
XNOR2_X1 U1107 ( .A(n1423), .B(n1202), .ZN(n1405) );
INV_X1 U1108 ( .A(G137), .ZN(n1202) );
NAND2_X1 U1109 ( .A1(G221), .A2(n1424), .ZN(n1423) );
XOR2_X1 U1110 ( .A(n1425), .B(n1262), .Z(n1173) );
INV_X1 U1111 ( .A(G472), .ZN(n1262) );
NAND2_X1 U1112 ( .A1(n1426), .A2(n1371), .ZN(n1425) );
XOR2_X1 U1113 ( .A(n1427), .B(n1428), .Z(n1426) );
XNOR2_X1 U1114 ( .A(n1259), .B(n1258), .ZN(n1428) );
XNOR2_X1 U1115 ( .A(n1429), .B(n1379), .ZN(n1258) );
INV_X1 U1116 ( .A(G101), .ZN(n1379) );
NAND2_X1 U1117 ( .A1(n1430), .A2(G210), .ZN(n1429) );
XNOR2_X1 U1118 ( .A(n1431), .B(n1387), .ZN(n1259) );
XOR2_X1 U1119 ( .A(n1402), .B(n1432), .Z(n1387) );
NOR2_X1 U1120 ( .A1(G143), .A2(KEYINPUT25), .ZN(n1432) );
XOR2_X1 U1121 ( .A(G128), .B(G146), .Z(n1402) );
NAND2_X1 U1122 ( .A1(n1433), .A2(n1434), .ZN(n1431) );
NAND2_X1 U1123 ( .A1(n1375), .A2(G119), .ZN(n1434) );
NAND2_X1 U1124 ( .A1(n1435), .A2(n1374), .ZN(n1433) );
INV_X1 U1125 ( .A(G119), .ZN(n1374) );
XNOR2_X1 U1126 ( .A(n1375), .B(KEYINPUT41), .ZN(n1435) );
XOR2_X1 U1127 ( .A(G113), .B(G116), .Z(n1375) );
XNOR2_X1 U1128 ( .A(n1263), .B(KEYINPUT9), .ZN(n1427) );
XOR2_X1 U1129 ( .A(G134), .B(n1400), .Z(n1263) );
XNOR2_X1 U1130 ( .A(n1198), .B(G137), .ZN(n1400) );
INV_X1 U1131 ( .A(G131), .ZN(n1198) );
AND2_X1 U1132 ( .A1(n1176), .A2(n1183), .ZN(n1141) );
INV_X1 U1133 ( .A(n1361), .ZN(n1183) );
XNOR2_X1 U1134 ( .A(n1436), .B(n1437), .ZN(n1361) );
XNOR2_X1 U1135 ( .A(KEYINPUT38), .B(n1252), .ZN(n1437) );
INV_X1 U1136 ( .A(G475), .ZN(n1252) );
NAND2_X1 U1137 ( .A1(n1250), .A2(n1371), .ZN(n1436) );
INV_X1 U1138 ( .A(G902), .ZN(n1371) );
XNOR2_X1 U1139 ( .A(n1438), .B(n1439), .ZN(n1250) );
XOR2_X1 U1140 ( .A(G113), .B(G104), .Z(n1439) );
XNOR2_X1 U1141 ( .A(n1382), .B(n1440), .ZN(n1438) );
NOR2_X1 U1142 ( .A1(KEYINPUT54), .A2(n1441), .ZN(n1440) );
XOR2_X1 U1143 ( .A(n1442), .B(n1443), .Z(n1441) );
XOR2_X1 U1144 ( .A(n1444), .B(n1445), .Z(n1443) );
NAND2_X1 U1145 ( .A1(n1430), .A2(G214), .ZN(n1445) );
NOR2_X1 U1146 ( .A1(G953), .A2(G237), .ZN(n1430) );
NAND2_X1 U1147 ( .A1(KEYINPUT61), .A2(n1446), .ZN(n1444) );
XOR2_X1 U1148 ( .A(G146), .B(n1422), .Z(n1446) );
XNOR2_X1 U1149 ( .A(G125), .B(n1201), .ZN(n1422) );
INV_X1 U1150 ( .A(G140), .ZN(n1201) );
XNOR2_X1 U1151 ( .A(n1339), .B(G131), .ZN(n1442) );
XNOR2_X1 U1152 ( .A(G478), .B(n1447), .ZN(n1176) );
NOR2_X1 U1153 ( .A1(G902), .A2(n1245), .ZN(n1447) );
XNOR2_X1 U1154 ( .A(n1448), .B(n1449), .ZN(n1245) );
AND2_X1 U1155 ( .A1(G217), .A2(n1424), .ZN(n1449) );
AND2_X1 U1156 ( .A1(G234), .A2(n1133), .ZN(n1424) );
INV_X1 U1157 ( .A(G953), .ZN(n1133) );
NAND2_X1 U1158 ( .A1(n1450), .A2(KEYINPUT20), .ZN(n1448) );
XOR2_X1 U1159 ( .A(n1451), .B(n1452), .Z(n1450) );
XOR2_X1 U1160 ( .A(G134), .B(n1453), .Z(n1452) );
NOR2_X1 U1161 ( .A1(KEYINPUT17), .A2(n1454), .ZN(n1453) );
XNOR2_X1 U1162 ( .A(n1339), .B(n1455), .ZN(n1454) );
NOR2_X1 U1163 ( .A1(G128), .A2(KEYINPUT42), .ZN(n1455) );
INV_X1 U1164 ( .A(G143), .ZN(n1339) );
NAND2_X1 U1165 ( .A1(n1456), .A2(n1457), .ZN(n1451) );
NAND2_X1 U1166 ( .A1(G107), .A2(n1458), .ZN(n1457) );
XOR2_X1 U1167 ( .A(KEYINPUT35), .B(n1459), .Z(n1456) );
NOR2_X1 U1168 ( .A1(G107), .A2(n1458), .ZN(n1459) );
XNOR2_X1 U1169 ( .A(n1460), .B(n1382), .ZN(n1458) );
XOR2_X1 U1170 ( .A(G122), .B(KEYINPUT15), .Z(n1382) );
XNOR2_X1 U1171 ( .A(G116), .B(KEYINPUT22), .ZN(n1460) );
INV_X1 U1172 ( .A(G110), .ZN(n1368) );
endmodule


