//Key = 0101011000101001110111011110001011011010101001110101110000110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341;

XOR2_X1 U721 ( .A(n1020), .B(n1021), .Z(G9) );
NAND4_X1 U722 ( .A1(KEYINPUT20), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1021) );
NAND3_X1 U723 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(G75) );
NAND2_X1 U724 ( .A1(G952), .A2(n1028), .ZN(n1027) );
NAND4_X1 U725 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1028) );
NAND4_X1 U726 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1032) );
NOR2_X1 U727 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U728 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NAND4_X1 U729 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1035) );
NAND2_X1 U730 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U731 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U732 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U733 ( .A1(n1024), .A2(n1051), .ZN(n1043) );
NAND2_X1 U734 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U735 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XOR2_X1 U736 ( .A(KEYINPUT61), .B(n1056), .Z(n1052) );
NAND2_X1 U737 ( .A1(n1057), .A2(n1058), .ZN(n1034) );
NAND2_X1 U738 ( .A1(n1059), .A2(n1042), .ZN(n1058) );
NAND2_X1 U739 ( .A1(n1045), .A2(n1024), .ZN(n1057) );
NAND2_X1 U740 ( .A1(n1060), .A2(n1061), .ZN(n1033) );
NAND2_X1 U741 ( .A1(n1042), .A2(n1062), .ZN(n1060) );
XOR2_X1 U742 ( .A(n1063), .B(KEYINPUT43), .Z(n1029) );
INV_X1 U743 ( .A(n1064), .ZN(n1026) );
NAND4_X1 U744 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1025) );
NOR4_X1 U745 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1068) );
XNOR2_X1 U746 ( .A(KEYINPUT44), .B(n1073), .ZN(n1072) );
XOR2_X1 U747 ( .A(KEYINPUT12), .B(n1074), .Z(n1070) );
NOR2_X1 U748 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U749 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U750 ( .A(KEYINPUT18), .B(G478), .Z(n1078) );
AND2_X1 U751 ( .A1(G478), .A2(n1077), .ZN(n1075) );
XNOR2_X1 U752 ( .A(n1079), .B(KEYINPUT32), .ZN(n1077) );
NOR3_X1 U753 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1067) );
INV_X1 U754 ( .A(n1083), .ZN(n1080) );
NAND2_X1 U755 ( .A1(n1084), .A2(n1085), .ZN(n1066) );
XNOR2_X1 U756 ( .A(n1086), .B(n1087), .ZN(n1065) );
XOR2_X1 U757 ( .A(n1088), .B(KEYINPUT21), .Z(n1087) );
NAND2_X1 U758 ( .A1(n1089), .A2(n1090), .ZN(G72) );
NAND2_X1 U759 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U760 ( .A1(G953), .A2(n1093), .ZN(n1091) );
NAND3_X1 U761 ( .A1(G953), .A2(n1094), .A3(n1095), .ZN(n1089) );
INV_X1 U762 ( .A(n1092), .ZN(n1095) );
NAND2_X1 U763 ( .A1(n1096), .A2(n1097), .ZN(n1092) );
NAND4_X1 U764 ( .A1(n1098), .A2(KEYINPUT51), .A3(n1031), .A4(n1099), .ZN(n1097) );
NAND2_X1 U765 ( .A1(G953), .A2(n1100), .ZN(n1099) );
NAND4_X1 U766 ( .A1(n1101), .A2(n1063), .A3(n1102), .A4(n1103), .ZN(n1096) );
NAND3_X1 U767 ( .A1(KEYINPUT51), .A2(n1098), .A3(n1104), .ZN(n1103) );
OR2_X1 U768 ( .A1(n1098), .A2(n1104), .ZN(n1102) );
INV_X1 U769 ( .A(KEYINPUT27), .ZN(n1104) );
XOR2_X1 U770 ( .A(n1105), .B(n1106), .Z(n1098) );
XNOR2_X1 U771 ( .A(n1107), .B(n1108), .ZN(n1106) );
XOR2_X1 U772 ( .A(KEYINPUT60), .B(KEYINPUT22), .Z(n1108) );
XNOR2_X1 U773 ( .A(n1109), .B(n1110), .ZN(n1105) );
NAND2_X1 U774 ( .A1(G900), .A2(G227), .ZN(n1094) );
XOR2_X1 U775 ( .A(n1111), .B(n1112), .Z(G69) );
NOR2_X1 U776 ( .A1(n1113), .A2(n1063), .ZN(n1112) );
NOR2_X1 U777 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U778 ( .A1(n1116), .A2(n1117), .ZN(n1111) );
NAND2_X1 U779 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XOR2_X1 U780 ( .A(n1120), .B(n1121), .Z(n1116) );
NOR2_X1 U781 ( .A1(n1030), .A2(G953), .ZN(n1121) );
OR2_X1 U782 ( .A1(n1119), .A2(n1118), .ZN(n1120) );
NAND2_X1 U783 ( .A1(n1122), .A2(n1123), .ZN(n1118) );
NAND2_X1 U784 ( .A1(G953), .A2(n1115), .ZN(n1123) );
XOR2_X1 U785 ( .A(n1124), .B(n1125), .Z(n1122) );
INV_X1 U786 ( .A(KEYINPUT5), .ZN(n1119) );
NOR2_X1 U787 ( .A1(n1064), .A2(n1126), .ZN(G66) );
XNOR2_X1 U788 ( .A(n1127), .B(n1128), .ZN(n1126) );
NOR2_X1 U789 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U790 ( .A1(n1064), .A2(n1131), .ZN(G63) );
NOR3_X1 U791 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
NOR3_X1 U792 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1134) );
NOR3_X1 U793 ( .A1(n1130), .A2(KEYINPUT29), .A3(n1138), .ZN(n1136) );
NOR2_X1 U794 ( .A1(KEYINPUT40), .A2(n1139), .ZN(n1133) );
NOR3_X1 U795 ( .A1(n1130), .A2(n1140), .A3(n1138), .ZN(n1132) );
NOR2_X1 U796 ( .A1(n1141), .A2(n1135), .ZN(n1140) );
INV_X1 U797 ( .A(KEYINPUT40), .ZN(n1135) );
NOR2_X1 U798 ( .A1(KEYINPUT29), .A2(n1139), .ZN(n1141) );
NOR2_X1 U799 ( .A1(n1064), .A2(n1142), .ZN(G60) );
XNOR2_X1 U800 ( .A(n1143), .B(n1144), .ZN(n1142) );
NOR2_X1 U801 ( .A1(n1088), .A2(n1130), .ZN(n1144) );
XOR2_X1 U802 ( .A(n1145), .B(n1146), .Z(G6) );
NOR2_X1 U803 ( .A1(n1064), .A2(n1147), .ZN(G57) );
NOR2_X1 U804 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U805 ( .A(n1150), .B(KEYINPUT36), .Z(n1149) );
NAND2_X1 U806 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U807 ( .A1(n1152), .A2(n1151), .ZN(n1148) );
XOR2_X1 U808 ( .A(n1153), .B(n1154), .Z(n1151) );
XOR2_X1 U809 ( .A(n1155), .B(n1109), .Z(n1154) );
NOR2_X1 U810 ( .A1(KEYINPUT9), .A2(n1156), .ZN(n1155) );
XOR2_X1 U811 ( .A(n1157), .B(n1158), .Z(n1153) );
NOR2_X1 U812 ( .A1(n1159), .A2(n1130), .ZN(n1158) );
INV_X1 U813 ( .A(G472), .ZN(n1159) );
NAND2_X1 U814 ( .A1(KEYINPUT26), .A2(n1160), .ZN(n1157) );
NOR2_X1 U815 ( .A1(n1161), .A2(n1162), .ZN(G54) );
XOR2_X1 U816 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U817 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND2_X1 U818 ( .A1(n1167), .A2(KEYINPUT58), .ZN(n1165) );
XOR2_X1 U819 ( .A(n1168), .B(KEYINPUT55), .Z(n1167) );
XOR2_X1 U820 ( .A(n1169), .B(n1170), .Z(n1163) );
NOR2_X1 U821 ( .A1(n1171), .A2(n1130), .ZN(n1170) );
XOR2_X1 U822 ( .A(n1172), .B(KEYINPUT28), .Z(n1169) );
NAND2_X1 U823 ( .A1(n1173), .A2(KEYINPUT25), .ZN(n1172) );
XOR2_X1 U824 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U825 ( .A(KEYINPUT19), .B(KEYINPUT11), .Z(n1175) );
NOR2_X1 U826 ( .A1(n1063), .A2(n1176), .ZN(n1161) );
XOR2_X1 U827 ( .A(KEYINPUT50), .B(G952), .Z(n1176) );
NOR2_X1 U828 ( .A1(n1064), .A2(n1177), .ZN(G51) );
XOR2_X1 U829 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U830 ( .A(n1180), .B(n1181), .Z(n1179) );
NAND2_X1 U831 ( .A1(KEYINPUT24), .A2(n1182), .ZN(n1180) );
XOR2_X1 U832 ( .A(n1183), .B(n1184), .Z(n1178) );
NOR2_X1 U833 ( .A1(n1185), .A2(n1130), .ZN(n1184) );
NAND2_X1 U834 ( .A1(G902), .A2(n1186), .ZN(n1130) );
NAND2_X1 U835 ( .A1(n1030), .A2(n1031), .ZN(n1186) );
INV_X1 U836 ( .A(n1101), .ZN(n1031) );
NAND4_X1 U837 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1101) );
AND3_X1 U838 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1190) );
NAND2_X1 U839 ( .A1(n1194), .A2(n1062), .ZN(n1189) );
INV_X1 U840 ( .A(n1041), .ZN(n1062) );
NOR2_X1 U841 ( .A1(n1195), .A2(n1023), .ZN(n1041) );
NAND2_X1 U842 ( .A1(n1196), .A2(n1197), .ZN(n1194) );
NAND3_X1 U843 ( .A1(n1198), .A2(n1047), .A3(n1199), .ZN(n1188) );
OR2_X1 U844 ( .A1(n1200), .A2(n1199), .ZN(n1187) );
INV_X1 U845 ( .A(KEYINPUT23), .ZN(n1199) );
AND2_X1 U846 ( .A1(n1201), .A2(n1202), .ZN(n1030) );
NOR4_X1 U847 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
INV_X1 U848 ( .A(n1207), .ZN(n1206) );
AND4_X1 U849 ( .A1(n1208), .A2(n1209), .A3(n1146), .A4(n1210), .ZN(n1201) );
NAND3_X1 U850 ( .A1(n1022), .A2(n1024), .A3(n1023), .ZN(n1210) );
NAND3_X1 U851 ( .A1(n1022), .A2(n1024), .A3(n1195), .ZN(n1146) );
XNOR2_X1 U852 ( .A(n1211), .B(KEYINPUT62), .ZN(n1183) );
NOR2_X1 U853 ( .A1(n1063), .A2(G952), .ZN(n1064) );
XOR2_X1 U854 ( .A(n1212), .B(n1213), .Z(G48) );
NAND2_X1 U855 ( .A1(KEYINPUT49), .A2(G146), .ZN(n1213) );
NAND2_X1 U856 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
XOR2_X1 U857 ( .A(KEYINPUT39), .B(n1195), .Z(n1215) );
XNOR2_X1 U858 ( .A(G143), .B(n1200), .ZN(G45) );
NAND2_X1 U859 ( .A1(n1198), .A2(n1216), .ZN(n1200) );
AND4_X1 U860 ( .A1(n1217), .A2(n1218), .A3(n1056), .A4(n1219), .ZN(n1198) );
XOR2_X1 U861 ( .A(n1220), .B(n1221), .Z(G42) );
NAND2_X1 U862 ( .A1(KEYINPUT59), .A2(n1222), .ZN(n1221) );
INV_X1 U863 ( .A(n1191), .ZN(n1222) );
NAND3_X1 U864 ( .A1(n1049), .A2(n1050), .A3(n1223), .ZN(n1191) );
XNOR2_X1 U865 ( .A(G137), .B(n1193), .ZN(G39) );
NAND4_X1 U866 ( .A1(n1218), .A2(n1224), .A3(n1225), .A4(n1045), .ZN(n1193) );
XOR2_X1 U867 ( .A(G134), .B(n1226), .Z(G36) );
NOR2_X1 U868 ( .A1(n1197), .A2(n1227), .ZN(n1226) );
XOR2_X1 U869 ( .A(KEYINPUT52), .B(n1023), .Z(n1227) );
NAND3_X1 U870 ( .A1(n1216), .A2(n1045), .A3(n1218), .ZN(n1197) );
XNOR2_X1 U871 ( .A(G131), .B(n1228), .ZN(G33) );
NAND2_X1 U872 ( .A1(n1223), .A2(n1216), .ZN(n1228) );
AND3_X1 U873 ( .A1(n1195), .A2(n1045), .A3(n1218), .ZN(n1223) );
INV_X1 U874 ( .A(n1071), .ZN(n1045) );
NAND2_X1 U875 ( .A1(n1055), .A2(n1229), .ZN(n1071) );
NAND2_X1 U876 ( .A1(n1230), .A2(n1231), .ZN(G30) );
NAND2_X1 U877 ( .A1(G128), .A2(n1232), .ZN(n1231) );
XOR2_X1 U878 ( .A(KEYINPUT46), .B(n1233), .Z(n1230) );
NOR2_X1 U879 ( .A1(G128), .A2(n1232), .ZN(n1233) );
NAND2_X1 U880 ( .A1(n1214), .A2(n1023), .ZN(n1232) );
INV_X1 U881 ( .A(n1196), .ZN(n1214) );
NAND4_X1 U882 ( .A1(n1225), .A2(n1218), .A3(n1056), .A4(n1050), .ZN(n1196) );
NOR3_X1 U883 ( .A1(n1234), .A2(n1039), .A3(n1082), .ZN(n1218) );
INV_X1 U884 ( .A(n1235), .ZN(n1039) );
XOR2_X1 U885 ( .A(G101), .B(n1205), .Z(G3) );
NOR3_X1 U886 ( .A1(n1047), .A2(n1236), .A3(n1061), .ZN(n1205) );
XOR2_X1 U887 ( .A(G125), .B(n1237), .Z(G27) );
NOR2_X1 U888 ( .A1(KEYINPUT37), .A2(n1192), .ZN(n1237) );
NAND4_X1 U889 ( .A1(n1042), .A2(n1056), .A3(n1195), .A4(n1238), .ZN(n1192) );
NOR3_X1 U890 ( .A1(n1225), .A2(n1239), .A3(n1234), .ZN(n1238) );
AND2_X1 U891 ( .A1(n1240), .A2(n1241), .ZN(n1234) );
NAND2_X1 U892 ( .A1(n1242), .A2(n1100), .ZN(n1240) );
INV_X1 U893 ( .A(G900), .ZN(n1100) );
XOR2_X1 U894 ( .A(n1243), .B(n1209), .Z(G24) );
NAND3_X1 U895 ( .A1(n1042), .A2(n1024), .A3(n1244), .ZN(n1209) );
AND3_X1 U896 ( .A1(n1217), .A2(n1219), .A3(n1245), .ZN(n1244) );
NOR2_X1 U897 ( .A1(n1050), .A2(n1225), .ZN(n1024) );
INV_X1 U898 ( .A(n1239), .ZN(n1050) );
XOR2_X1 U899 ( .A(n1246), .B(n1208), .Z(G21) );
NAND4_X1 U900 ( .A1(n1224), .A2(n1042), .A3(n1225), .A4(n1245), .ZN(n1208) );
XOR2_X1 U901 ( .A(G116), .B(n1204), .Z(G18) );
AND2_X1 U902 ( .A1(n1247), .A2(n1023), .ZN(n1204) );
NOR2_X1 U903 ( .A1(n1219), .A2(n1248), .ZN(n1023) );
XOR2_X1 U904 ( .A(G113), .B(n1203), .Z(G15) );
AND2_X1 U905 ( .A1(n1247), .A2(n1195), .ZN(n1203) );
AND2_X1 U906 ( .A1(n1248), .A2(n1219), .ZN(n1195) );
INV_X1 U907 ( .A(n1217), .ZN(n1248) );
AND3_X1 U908 ( .A1(n1042), .A2(n1245), .A3(n1216), .ZN(n1247) );
INV_X1 U909 ( .A(n1047), .ZN(n1216) );
NAND2_X1 U910 ( .A1(n1225), .A2(n1239), .ZN(n1047) );
NOR2_X1 U911 ( .A1(n1235), .A2(n1082), .ZN(n1042) );
INV_X1 U912 ( .A(n1040), .ZN(n1082) );
NAND3_X1 U913 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(G12) );
OR2_X1 U914 ( .A1(n1207), .A2(KEYINPUT16), .ZN(n1251) );
NAND3_X1 U915 ( .A1(KEYINPUT16), .A2(n1207), .A3(G110), .ZN(n1250) );
NAND2_X1 U916 ( .A1(n1252), .A2(n1253), .ZN(n1249) );
NAND2_X1 U917 ( .A1(n1254), .A2(KEYINPUT16), .ZN(n1252) );
XOR2_X1 U918 ( .A(n1207), .B(KEYINPUT7), .Z(n1254) );
NAND3_X1 U919 ( .A1(n1022), .A2(n1049), .A3(n1224), .ZN(n1207) );
NOR2_X1 U920 ( .A1(n1061), .A2(n1239), .ZN(n1224) );
NOR2_X1 U921 ( .A1(n1255), .A2(n1081), .ZN(n1239) );
NOR2_X1 U922 ( .A1(n1085), .A2(n1084), .ZN(n1081) );
AND2_X1 U923 ( .A1(n1084), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U924 ( .A(KEYINPUT17), .B(n1085), .ZN(n1256) );
NAND2_X1 U925 ( .A1(n1257), .A2(n1258), .ZN(n1085) );
XOR2_X1 U926 ( .A(n1127), .B(KEYINPUT13), .Z(n1257) );
NAND2_X1 U927 ( .A1(n1259), .A2(n1260), .ZN(n1127) );
NAND2_X1 U928 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U929 ( .A(KEYINPUT42), .B(n1263), .Z(n1259) );
NOR2_X1 U930 ( .A1(n1261), .A2(n1262), .ZN(n1263) );
XOR2_X1 U931 ( .A(n1264), .B(n1265), .Z(n1262) );
XOR2_X1 U932 ( .A(G146), .B(n1266), .Z(n1265) );
NOR2_X1 U933 ( .A1(KEYINPUT34), .A2(n1267), .ZN(n1266) );
XOR2_X1 U934 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U935 ( .A(n1253), .B(G128), .Z(n1269) );
NAND2_X1 U936 ( .A1(KEYINPUT10), .A2(n1246), .ZN(n1268) );
XOR2_X1 U937 ( .A(n1270), .B(G137), .Z(n1261) );
NAND2_X1 U938 ( .A1(n1271), .A2(G221), .ZN(n1270) );
INV_X1 U939 ( .A(n1129), .ZN(n1084) );
NAND2_X1 U940 ( .A1(G217), .A2(n1272), .ZN(n1129) );
INV_X1 U941 ( .A(n1059), .ZN(n1061) );
NOR2_X1 U942 ( .A1(n1219), .A2(n1217), .ZN(n1059) );
XOR2_X1 U943 ( .A(n1079), .B(n1273), .Z(n1217) );
NOR2_X1 U944 ( .A1(KEYINPUT4), .A2(n1274), .ZN(n1273) );
XOR2_X1 U945 ( .A(n1138), .B(KEYINPUT6), .Z(n1274) );
INV_X1 U946 ( .A(G478), .ZN(n1138) );
NAND2_X1 U947 ( .A1(n1258), .A2(n1139), .ZN(n1079) );
INV_X1 U948 ( .A(n1137), .ZN(n1139) );
XOR2_X1 U949 ( .A(n1275), .B(n1276), .Z(n1137) );
XOR2_X1 U950 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U951 ( .A(G134), .B(G122), .Z(n1278) );
XOR2_X1 U952 ( .A(KEYINPUT53), .B(G143), .Z(n1277) );
XOR2_X1 U953 ( .A(n1279), .B(n1280), .Z(n1275) );
XOR2_X1 U954 ( .A(G116), .B(G107), .Z(n1280) );
XOR2_X1 U955 ( .A(n1281), .B(n1282), .Z(n1279) );
NOR2_X1 U956 ( .A1(KEYINPUT63), .A2(G128), .ZN(n1282) );
NAND2_X1 U957 ( .A1(G217), .A2(n1271), .ZN(n1281) );
NOR2_X1 U958 ( .A1(n1283), .A2(n1284), .ZN(n1271) );
INV_X1 U959 ( .A(G234), .ZN(n1283) );
NAND2_X1 U960 ( .A1(n1285), .A2(n1286), .ZN(n1219) );
NAND2_X1 U961 ( .A1(n1086), .A2(n1088), .ZN(n1286) );
XOR2_X1 U962 ( .A(KEYINPUT30), .B(n1287), .Z(n1285) );
NOR2_X1 U963 ( .A1(n1086), .A2(n1088), .ZN(n1287) );
INV_X1 U964 ( .A(G475), .ZN(n1088) );
AND2_X1 U965 ( .A1(n1258), .A2(n1143), .ZN(n1086) );
XNOR2_X1 U966 ( .A(n1288), .B(n1289), .ZN(n1143) );
XOR2_X1 U967 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U968 ( .A(G113), .B(G104), .Z(n1291) );
NOR2_X1 U969 ( .A1(KEYINPUT56), .A2(n1243), .ZN(n1290) );
INV_X1 U970 ( .A(G122), .ZN(n1243) );
XOR2_X1 U971 ( .A(n1292), .B(n1110), .Z(n1288) );
XOR2_X1 U972 ( .A(G131), .B(n1264), .Z(n1110) );
XOR2_X1 U973 ( .A(G125), .B(G140), .Z(n1264) );
XOR2_X1 U974 ( .A(n1293), .B(n1294), .Z(n1292) );
NAND2_X1 U975 ( .A1(n1295), .A2(G214), .ZN(n1293) );
INV_X1 U976 ( .A(n1225), .ZN(n1049) );
XNOR2_X1 U977 ( .A(n1069), .B(KEYINPUT47), .ZN(n1225) );
XNOR2_X1 U978 ( .A(n1296), .B(G472), .ZN(n1069) );
NAND2_X1 U979 ( .A1(n1297), .A2(n1258), .ZN(n1296) );
XOR2_X1 U980 ( .A(n1298), .B(n1299), .Z(n1297) );
XOR2_X1 U981 ( .A(n1109), .B(n1152), .Z(n1299) );
AND2_X1 U982 ( .A1(n1300), .A2(n1301), .ZN(n1152) );
NAND2_X1 U983 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NAND2_X1 U984 ( .A1(n1295), .A2(G210), .ZN(n1303) );
NAND3_X1 U985 ( .A1(n1295), .A2(G210), .A3(n1304), .ZN(n1300) );
NOR2_X1 U986 ( .A1(n1284), .A2(G237), .ZN(n1295) );
XOR2_X1 U987 ( .A(n1305), .B(n1156), .Z(n1298) );
XNOR2_X1 U988 ( .A(n1306), .B(G113), .ZN(n1156) );
NAND3_X1 U989 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1306) );
NAND2_X1 U990 ( .A1(G116), .A2(n1310), .ZN(n1309) );
INV_X1 U991 ( .A(KEYINPUT35), .ZN(n1310) );
NAND3_X1 U992 ( .A1(KEYINPUT35), .A2(n1311), .A3(n1246), .ZN(n1308) );
OR2_X1 U993 ( .A1(n1246), .A2(n1311), .ZN(n1307) );
NOR2_X1 U994 ( .A1(G116), .A2(KEYINPUT0), .ZN(n1311) );
INV_X1 U995 ( .A(G119), .ZN(n1246) );
NOR2_X1 U996 ( .A1(KEYINPUT57), .A2(n1160), .ZN(n1305) );
INV_X1 U997 ( .A(n1236), .ZN(n1022) );
NAND3_X1 U998 ( .A1(n1040), .A2(n1235), .A3(n1245), .ZN(n1236) );
AND2_X1 U999 ( .A1(n1056), .A2(n1312), .ZN(n1245) );
NAND2_X1 U1000 ( .A1(n1313), .A2(n1241), .ZN(n1312) );
NAND2_X1 U1001 ( .A1(n1314), .A2(n1315), .ZN(n1241) );
INV_X1 U1002 ( .A(n1038), .ZN(n1315) );
NAND2_X1 U1003 ( .A1(n1063), .A2(n1316), .ZN(n1038) );
XNOR2_X1 U1004 ( .A(G952), .B(KEYINPUT38), .ZN(n1314) );
NAND2_X1 U1005 ( .A1(n1242), .A2(n1115), .ZN(n1313) );
INV_X1 U1006 ( .A(G898), .ZN(n1115) );
AND3_X1 U1007 ( .A1(G902), .A2(n1316), .A3(G953), .ZN(n1242) );
NAND2_X1 U1008 ( .A1(G237), .A2(G234), .ZN(n1316) );
NOR2_X1 U1009 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
INV_X1 U1010 ( .A(n1229), .ZN(n1054) );
NAND2_X1 U1011 ( .A1(G214), .A2(n1317), .ZN(n1229) );
XNOR2_X1 U1012 ( .A(n1318), .B(n1185), .ZN(n1055) );
NAND2_X1 U1013 ( .A1(G210), .A2(n1317), .ZN(n1185) );
NAND2_X1 U1014 ( .A1(n1319), .A2(n1320), .ZN(n1317) );
INV_X1 U1015 ( .A(G237), .ZN(n1319) );
NAND2_X1 U1016 ( .A1(n1258), .A2(n1321), .ZN(n1318) );
XOR2_X1 U1017 ( .A(n1182), .B(n1322), .Z(n1321) );
XNOR2_X1 U1018 ( .A(n1181), .B(n1211), .ZN(n1322) );
NOR2_X1 U1019 ( .A1(n1114), .A2(n1284), .ZN(n1211) );
INV_X1 U1020 ( .A(G224), .ZN(n1114) );
XNOR2_X1 U1021 ( .A(n1124), .B(n1323), .ZN(n1181) );
XNOR2_X1 U1022 ( .A(n1324), .B(KEYINPUT41), .ZN(n1323) );
NAND2_X1 U1023 ( .A1(KEYINPUT15), .A2(n1125), .ZN(n1324) );
XOR2_X1 U1024 ( .A(n1253), .B(n1325), .Z(n1125) );
XOR2_X1 U1025 ( .A(KEYINPUT3), .B(G122), .Z(n1325) );
INV_X1 U1026 ( .A(G110), .ZN(n1253) );
XOR2_X1 U1027 ( .A(n1326), .B(n1327), .Z(n1124) );
XNOR2_X1 U1028 ( .A(n1328), .B(n1329), .ZN(n1327) );
NAND2_X1 U1029 ( .A1(KEYINPUT1), .A2(G119), .ZN(n1328) );
XOR2_X1 U1030 ( .A(n1330), .B(n1331), .Z(n1326) );
XOR2_X1 U1031 ( .A(G116), .B(G113), .Z(n1331) );
NAND2_X1 U1032 ( .A1(KEYINPUT45), .A2(n1304), .ZN(n1330) );
XNOR2_X1 U1033 ( .A(G125), .B(n1109), .ZN(n1182) );
NAND2_X1 U1034 ( .A1(n1083), .A2(n1073), .ZN(n1235) );
NAND2_X1 U1035 ( .A1(G469), .A2(n1332), .ZN(n1073) );
NAND2_X1 U1036 ( .A1(n1258), .A2(n1333), .ZN(n1332) );
NAND3_X1 U1037 ( .A1(n1333), .A2(n1171), .A3(n1258), .ZN(n1083) );
XOR2_X1 U1038 ( .A(n1320), .B(KEYINPUT31), .Z(n1258) );
INV_X1 U1039 ( .A(G469), .ZN(n1171) );
XNOR2_X1 U1040 ( .A(n1168), .B(n1334), .ZN(n1333) );
XOR2_X1 U1041 ( .A(n1166), .B(n1335), .Z(n1334) );
INV_X1 U1042 ( .A(n1174), .ZN(n1335) );
XOR2_X1 U1043 ( .A(n1336), .B(n1337), .Z(n1174) );
NOR2_X1 U1044 ( .A1(n1284), .A2(n1093), .ZN(n1337) );
INV_X1 U1045 ( .A(G227), .ZN(n1093) );
XNOR2_X1 U1046 ( .A(n1063), .B(KEYINPUT2), .ZN(n1284) );
INV_X1 U1047 ( .A(G953), .ZN(n1063) );
XOR2_X1 U1048 ( .A(n1220), .B(G110), .Z(n1336) );
INV_X1 U1049 ( .A(G140), .ZN(n1220) );
XOR2_X1 U1050 ( .A(n1304), .B(n1338), .Z(n1166) );
XNOR2_X1 U1051 ( .A(n1339), .B(n1160), .ZN(n1338) );
XNOR2_X1 U1052 ( .A(G131), .B(n1340), .ZN(n1160) );
NOR2_X1 U1053 ( .A1(KEYINPUT14), .A2(n1107), .ZN(n1340) );
XNOR2_X1 U1054 ( .A(G134), .B(n1341), .ZN(n1107) );
XOR2_X1 U1055 ( .A(KEYINPUT8), .B(G137), .Z(n1341) );
NOR2_X1 U1056 ( .A1(KEYINPUT54), .A2(n1329), .ZN(n1339) );
XOR2_X1 U1057 ( .A(n1145), .B(n1020), .Z(n1329) );
INV_X1 U1058 ( .A(G107), .ZN(n1020) );
INV_X1 U1059 ( .A(G104), .ZN(n1145) );
INV_X1 U1060 ( .A(n1302), .ZN(n1304) );
XNOR2_X1 U1061 ( .A(G101), .B(KEYINPUT48), .ZN(n1302) );
XNOR2_X1 U1062 ( .A(n1109), .B(KEYINPUT33), .ZN(n1168) );
XOR2_X1 U1063 ( .A(G128), .B(n1294), .Z(n1109) );
XOR2_X1 U1064 ( .A(G143), .B(G146), .Z(n1294) );
NAND2_X1 U1065 ( .A1(G221), .A2(n1272), .ZN(n1040) );
NAND2_X1 U1066 ( .A1(G234), .A2(n1320), .ZN(n1272) );
INV_X1 U1067 ( .A(G902), .ZN(n1320) );
endmodule


