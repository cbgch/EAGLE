//Key = 0100101111000000101100110010111101000001110000100110100011010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263;

XOR2_X1 U697 ( .A(n958), .B(n959), .Z(G9) );
NOR2_X1 U698 ( .A1(n960), .A2(n961), .ZN(G75) );
NOR2_X1 U699 ( .A1(n962), .A2(n963), .ZN(n961) );
NAND4_X1 U700 ( .A1(n964), .A2(n965), .A3(G952), .A4(n966), .ZN(n963) );
XOR2_X1 U701 ( .A(KEYINPUT56), .B(n967), .Z(n966) );
AND4_X1 U702 ( .A1(n968), .A2(n969), .A3(n970), .A4(n971), .ZN(n967) );
NAND4_X1 U703 ( .A1(n972), .A2(n973), .A3(n974), .A4(n975), .ZN(n962) );
NAND2_X1 U704 ( .A1(n976), .A2(n968), .ZN(n972) );
NAND2_X1 U705 ( .A1(n977), .A2(n978), .ZN(n976) );
NAND3_X1 U706 ( .A1(n979), .A2(n980), .A3(n969), .ZN(n978) );
NAND2_X1 U707 ( .A1(n981), .A2(n982), .ZN(n980) );
NAND2_X1 U708 ( .A1(n983), .A2(n984), .ZN(n982) );
NAND2_X1 U709 ( .A1(n985), .A2(n986), .ZN(n984) );
NAND2_X1 U710 ( .A1(n987), .A2(n988), .ZN(n986) );
NAND2_X1 U711 ( .A1(n970), .A2(n989), .ZN(n981) );
NAND3_X1 U712 ( .A1(n983), .A2(n990), .A3(n970), .ZN(n977) );
NAND2_X1 U713 ( .A1(n991), .A2(n992), .ZN(n990) );
NAND2_X1 U714 ( .A1(n969), .A2(n993), .ZN(n992) );
OR2_X1 U715 ( .A1(n994), .A2(n995), .ZN(n993) );
NAND2_X1 U716 ( .A1(n979), .A2(n996), .ZN(n991) );
NAND2_X1 U717 ( .A1(n997), .A2(n998), .ZN(n996) );
NAND2_X1 U718 ( .A1(n999), .A2(n1000), .ZN(n998) );
NOR3_X1 U719 ( .A1(n1001), .A2(G953), .A3(n1002), .ZN(n960) );
INV_X1 U720 ( .A(n974), .ZN(n1002) );
NAND4_X1 U721 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n974) );
NOR4_X1 U722 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1006) );
XOR2_X1 U723 ( .A(n1011), .B(n1012), .Z(n1007) );
NOR2_X1 U724 ( .A1(KEYINPUT38), .A2(n1013), .ZN(n1012) );
XOR2_X1 U725 ( .A(KEYINPUT32), .B(G478), .Z(n1013) );
NOR3_X1 U726 ( .A1(n999), .A2(n1014), .A3(n987), .ZN(n1005) );
NAND2_X1 U727 ( .A1(G472), .A2(n1015), .ZN(n1004) );
XOR2_X1 U728 ( .A(n1016), .B(KEYINPUT37), .Z(n1003) );
NAND2_X1 U729 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND2_X1 U730 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
XOR2_X1 U731 ( .A(n1021), .B(KEYINPUT20), .Z(n1019) );
NAND2_X1 U732 ( .A1(n1022), .A2(n1023), .ZN(n1017) );
XOR2_X1 U733 ( .A(n1021), .B(KEYINPUT4), .Z(n1022) );
XNOR2_X1 U734 ( .A(G952), .B(KEYINPUT31), .ZN(n1001) );
XOR2_X1 U735 ( .A(n1024), .B(n1025), .Z(G72) );
XOR2_X1 U736 ( .A(n1026), .B(n1027), .Z(n1025) );
NOR2_X1 U737 ( .A1(G953), .A2(n1028), .ZN(n1027) );
XOR2_X1 U738 ( .A(KEYINPUT47), .B(n964), .Z(n1028) );
NOR2_X1 U739 ( .A1(n1029), .A2(n1030), .ZN(n1026) );
XNOR2_X1 U740 ( .A(n1031), .B(n1032), .ZN(n1030) );
XOR2_X1 U741 ( .A(n1033), .B(KEYINPUT11), .Z(n1032) );
NOR2_X1 U742 ( .A1(G900), .A2(n975), .ZN(n1029) );
NOR3_X1 U743 ( .A1(n975), .A2(KEYINPUT12), .A3(n1034), .ZN(n1024) );
AND2_X1 U744 ( .A1(G227), .A2(G900), .ZN(n1034) );
XOR2_X1 U745 ( .A(n1035), .B(n1036), .Z(G69) );
NOR2_X1 U746 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U747 ( .A1(G898), .A2(n975), .ZN(n1037) );
NAND2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1035) );
NAND2_X1 U749 ( .A1(n1041), .A2(n975), .ZN(n1040) );
NAND2_X1 U750 ( .A1(n1042), .A2(n965), .ZN(n1041) );
XOR2_X1 U751 ( .A(n973), .B(KEYINPUT54), .Z(n1042) );
NAND2_X1 U752 ( .A1(G953), .A2(n1043), .ZN(n1039) );
NAND2_X1 U753 ( .A1(G898), .A2(n1044), .ZN(n1043) );
XOR2_X1 U754 ( .A(KEYINPUT25), .B(G224), .Z(n1044) );
NOR2_X1 U755 ( .A1(n1045), .A2(n1046), .ZN(G66) );
NOR2_X1 U756 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
XOR2_X1 U757 ( .A(KEYINPUT5), .B(n1049), .Z(n1048) );
NOR2_X1 U758 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
XNOR2_X1 U759 ( .A(KEYINPUT10), .B(n1052), .ZN(n1051) );
NOR2_X1 U760 ( .A1(n1053), .A2(n1052), .ZN(n1047) );
NAND2_X1 U761 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U762 ( .A1(n1045), .A2(n1056), .ZN(G63) );
XOR2_X1 U763 ( .A(n1057), .B(n1058), .Z(n1056) );
AND2_X1 U764 ( .A1(G478), .A2(n1054), .ZN(n1058) );
NAND2_X1 U765 ( .A1(KEYINPUT59), .A2(n1059), .ZN(n1057) );
NOR2_X1 U766 ( .A1(n1045), .A2(n1060), .ZN(G60) );
XOR2_X1 U767 ( .A(n1061), .B(n1062), .Z(n1060) );
NAND3_X1 U768 ( .A1(n1054), .A2(G475), .A3(KEYINPUT18), .ZN(n1061) );
XOR2_X1 U769 ( .A(G104), .B(n1063), .Z(G6) );
AND2_X1 U770 ( .A1(n1064), .A2(n971), .ZN(n1063) );
NOR2_X1 U771 ( .A1(n1045), .A2(n1065), .ZN(G57) );
NOR2_X1 U772 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
XOR2_X1 U773 ( .A(KEYINPUT43), .B(n1068), .Z(n1067) );
NOR2_X1 U774 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XOR2_X1 U775 ( .A(n1071), .B(n1072), .Z(n1070) );
NOR2_X1 U776 ( .A1(n1073), .A2(n1074), .ZN(n1066) );
XNOR2_X1 U777 ( .A(n1072), .B(n1071), .ZN(n1073) );
XOR2_X1 U778 ( .A(n1075), .B(n1076), .Z(n1072) );
NOR2_X1 U779 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR2_X1 U780 ( .A1(n1045), .A2(n1079), .ZN(G54) );
XOR2_X1 U781 ( .A(n1080), .B(n1081), .Z(n1079) );
XNOR2_X1 U782 ( .A(n1082), .B(n1083), .ZN(n1081) );
NOR3_X1 U783 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1082) );
NOR2_X1 U784 ( .A1(G110), .A2(n1087), .ZN(n1086) );
NOR2_X1 U785 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U786 ( .A(KEYINPUT53), .B(G140), .Z(n1089) );
NOR3_X1 U787 ( .A1(n1090), .A2(G140), .A3(n1088), .ZN(n1085) );
INV_X1 U788 ( .A(KEYINPUT16), .ZN(n1088) );
NOR2_X1 U789 ( .A1(KEYINPUT16), .A2(n1091), .ZN(n1084) );
XOR2_X1 U790 ( .A(n1092), .B(n1093), .Z(n1080) );
AND2_X1 U791 ( .A1(G469), .A2(n1054), .ZN(n1093) );
INV_X1 U792 ( .A(n1078), .ZN(n1054) );
NOR2_X1 U793 ( .A1(n1045), .A2(n1094), .ZN(G51) );
XOR2_X1 U794 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U795 ( .A1(n1020), .A2(n1078), .ZN(n1096) );
NAND2_X1 U796 ( .A1(G902), .A2(n1097), .ZN(n1078) );
NAND3_X1 U797 ( .A1(n965), .A2(n973), .A3(n964), .ZN(n1097) );
AND4_X1 U798 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n964) );
NOR4_X1 U799 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1101) );
INV_X1 U800 ( .A(n1106), .ZN(n1102) );
AND2_X1 U801 ( .A1(n1107), .A2(n1108), .ZN(n1100) );
NAND4_X1 U802 ( .A1(n971), .A2(n1109), .A3(n1110), .A4(n1111), .ZN(n973) );
XOR2_X1 U803 ( .A(KEYINPUT61), .B(n1112), .Z(n1111) );
AND2_X1 U804 ( .A1(n1113), .A2(n979), .ZN(n971) );
AND4_X1 U805 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n965) );
AND3_X1 U806 ( .A1(n959), .A2(n1118), .A3(n1119), .ZN(n1117) );
NAND3_X1 U807 ( .A1(n1064), .A2(n989), .A3(n979), .ZN(n959) );
NAND2_X1 U808 ( .A1(n1120), .A2(n1121), .ZN(n1116) );
NAND2_X1 U809 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND3_X1 U810 ( .A1(n1124), .A2(n1009), .A3(n979), .ZN(n1123) );
NAND2_X1 U811 ( .A1(n994), .A2(n989), .ZN(n1122) );
NOR2_X1 U812 ( .A1(n1125), .A2(n1126), .ZN(n1095) );
XOR2_X1 U813 ( .A(n1127), .B(KEYINPUT1), .Z(n1126) );
NAND2_X1 U814 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR2_X1 U815 ( .A1(n1130), .A2(n1128), .ZN(n1125) );
XOR2_X1 U816 ( .A(KEYINPUT58), .B(n1131), .Z(n1128) );
XOR2_X1 U817 ( .A(KEYINPUT27), .B(n1129), .Z(n1130) );
XNOR2_X1 U818 ( .A(n1132), .B(n1133), .ZN(n1129) );
XOR2_X1 U819 ( .A(n1134), .B(n1135), .Z(n1132) );
NOR2_X1 U820 ( .A1(n975), .A2(G952), .ZN(n1045) );
XOR2_X1 U821 ( .A(n1136), .B(G146), .Z(G48) );
NAND2_X1 U822 ( .A1(KEYINPUT7), .A2(n1098), .ZN(n1136) );
NAND3_X1 U823 ( .A1(n1137), .A2(n1112), .A3(n1113), .ZN(n1098) );
XOR2_X1 U824 ( .A(G143), .B(n1105), .Z(G45) );
AND3_X1 U825 ( .A1(n994), .A2(n1138), .A3(n1139), .ZN(n1105) );
NOR3_X1 U826 ( .A1(n997), .A2(n1140), .A3(n1141), .ZN(n1139) );
XOR2_X1 U827 ( .A(G140), .B(n1104), .Z(G42) );
AND2_X1 U828 ( .A1(n1142), .A2(n995), .ZN(n1104) );
XNOR2_X1 U829 ( .A(G137), .B(n1099), .ZN(G39) );
NAND3_X1 U830 ( .A1(n969), .A2(n1137), .A3(n983), .ZN(n1099) );
XOR2_X1 U831 ( .A(n1108), .B(n1143), .Z(G36) );
XNOR2_X1 U832 ( .A(G134), .B(KEYINPUT2), .ZN(n1143) );
NAND4_X1 U833 ( .A1(n994), .A2(n969), .A3(n1138), .A4(n989), .ZN(n1108) );
XOR2_X1 U834 ( .A(G131), .B(n1103), .Z(G33) );
AND2_X1 U835 ( .A1(n1142), .A2(n994), .ZN(n1103) );
AND3_X1 U836 ( .A1(n969), .A2(n1138), .A3(n1113), .ZN(n1142) );
NOR2_X1 U837 ( .A1(n1144), .A2(n999), .ZN(n969) );
INV_X1 U838 ( .A(n1000), .ZN(n1144) );
XOR2_X1 U839 ( .A(n1145), .B(n1107), .Z(G30) );
NAND3_X1 U840 ( .A1(n989), .A2(n1112), .A3(n1137), .ZN(n1107) );
AND3_X1 U841 ( .A1(n1146), .A2(n1008), .A3(n1138), .ZN(n1137) );
NOR2_X1 U842 ( .A1(n1147), .A2(n985), .ZN(n1138) );
XOR2_X1 U843 ( .A(n1119), .B(n1148), .Z(G3) );
XOR2_X1 U844 ( .A(KEYINPUT9), .B(G101), .Z(n1148) );
NAND3_X1 U845 ( .A1(n994), .A2(n1064), .A3(n983), .ZN(n1119) );
XOR2_X1 U846 ( .A(n1134), .B(n1106), .Z(G27) );
NAND3_X1 U847 ( .A1(n970), .A2(n995), .A3(n1149), .ZN(n1106) );
NOR3_X1 U848 ( .A1(n1150), .A2(n997), .A3(n1147), .ZN(n1149) );
NAND2_X1 U849 ( .A1(n1151), .A2(n968), .ZN(n1147) );
NAND2_X1 U850 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
OR3_X1 U851 ( .A1(n1154), .A2(G900), .A3(n975), .ZN(n1153) );
INV_X1 U852 ( .A(n1155), .ZN(n970) );
XOR2_X1 U853 ( .A(n1156), .B(n1157), .Z(G24) );
NAND4_X1 U854 ( .A1(n1120), .A2(n1158), .A3(n1124), .A4(n1009), .ZN(n1157) );
XOR2_X1 U855 ( .A(KEYINPUT45), .B(n979), .Z(n1158) );
NOR2_X1 U856 ( .A1(n1159), .A2(n1008), .ZN(n979) );
XOR2_X1 U857 ( .A(n1114), .B(n1160), .Z(G21) );
XNOR2_X1 U858 ( .A(G119), .B(KEYINPUT60), .ZN(n1160) );
NAND4_X1 U859 ( .A1(n1120), .A2(n983), .A3(n1146), .A4(n1008), .ZN(n1114) );
XNOR2_X1 U860 ( .A(G116), .B(n1161), .ZN(G18) );
NAND3_X1 U861 ( .A1(n1162), .A2(n994), .A3(n1163), .ZN(n1161) );
AND3_X1 U862 ( .A1(n989), .A2(n1112), .A3(n1110), .ZN(n1163) );
INV_X1 U863 ( .A(n1164), .ZN(n1110) );
NOR2_X1 U864 ( .A1(n1009), .A2(n1141), .ZN(n989) );
XOR2_X1 U865 ( .A(n1155), .B(KEYINPUT29), .Z(n1162) );
XOR2_X1 U866 ( .A(n1165), .B(n1115), .Z(G15) );
NAND3_X1 U867 ( .A1(n1113), .A2(n994), .A3(n1120), .ZN(n1115) );
NOR3_X1 U868 ( .A1(n1164), .A2(n997), .A3(n1155), .ZN(n1120) );
NAND2_X1 U869 ( .A1(n988), .A2(n1166), .ZN(n1155) );
AND2_X1 U870 ( .A1(n1146), .A2(n1167), .ZN(n994) );
XOR2_X1 U871 ( .A(n1159), .B(KEYINPUT48), .Z(n1146) );
INV_X1 U872 ( .A(n1150), .ZN(n1113) );
NAND2_X1 U873 ( .A1(n1141), .A2(n1009), .ZN(n1150) );
XNOR2_X1 U874 ( .A(n1168), .B(n1118), .ZN(G12) );
NAND3_X1 U875 ( .A1(n983), .A2(n1064), .A3(n995), .ZN(n1118) );
NOR2_X1 U876 ( .A1(n1159), .A2(n1167), .ZN(n995) );
INV_X1 U877 ( .A(n1008), .ZN(n1167) );
XNOR2_X1 U878 ( .A(n1169), .B(n1055), .ZN(n1008) );
AND2_X1 U879 ( .A1(G217), .A2(n1170), .ZN(n1055) );
NAND2_X1 U880 ( .A1(n1053), .A2(n1154), .ZN(n1169) );
INV_X1 U881 ( .A(n1050), .ZN(n1053) );
XOR2_X1 U882 ( .A(n1171), .B(n1172), .Z(n1050) );
NOR2_X1 U883 ( .A1(G137), .A2(KEYINPUT17), .ZN(n1172) );
XOR2_X1 U884 ( .A(n1173), .B(n1174), .Z(n1171) );
NOR2_X1 U885 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
INV_X1 U886 ( .A(G221), .ZN(n1176) );
NAND2_X1 U887 ( .A1(n1177), .A2(n1178), .ZN(n1173) );
OR2_X1 U888 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XOR2_X1 U889 ( .A(n1181), .B(KEYINPUT3), .Z(n1177) );
NAND2_X1 U890 ( .A1(n1180), .A2(n1179), .ZN(n1181) );
XNOR2_X1 U891 ( .A(n1182), .B(n1183), .ZN(n1179) );
XOR2_X1 U892 ( .A(KEYINPUT8), .B(KEYINPUT36), .Z(n1183) );
XOR2_X1 U893 ( .A(n1184), .B(n1031), .Z(n1182) );
XOR2_X1 U894 ( .A(n1134), .B(n1091), .Z(n1031) );
XNOR2_X1 U895 ( .A(n1090), .B(n1185), .ZN(n1180) );
XOR2_X1 U896 ( .A(G128), .B(G119), .Z(n1185) );
NAND3_X1 U897 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1159) );
INV_X1 U898 ( .A(n1014), .ZN(n1188) );
NOR2_X1 U899 ( .A1(n1015), .A2(G472), .ZN(n1014) );
NAND2_X1 U900 ( .A1(KEYINPUT14), .A2(n1077), .ZN(n1187) );
INV_X1 U901 ( .A(G472), .ZN(n1077) );
NAND3_X1 U902 ( .A1(n1015), .A2(n1189), .A3(G472), .ZN(n1186) );
INV_X1 U903 ( .A(KEYINPUT14), .ZN(n1189) );
NAND2_X1 U904 ( .A1(n1190), .A2(n1154), .ZN(n1015) );
XOR2_X1 U905 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U906 ( .A(n1071), .B(n1074), .Z(n1192) );
INV_X1 U907 ( .A(n1069), .ZN(n1074) );
XOR2_X1 U908 ( .A(n1193), .B(G101), .Z(n1069) );
NAND2_X1 U909 ( .A1(G210), .A2(n1194), .ZN(n1193) );
XNOR2_X1 U910 ( .A(n1195), .B(KEYINPUT42), .ZN(n1191) );
NAND2_X1 U911 ( .A1(KEYINPUT19), .A2(n1075), .ZN(n1195) );
XNOR2_X1 U912 ( .A(n1165), .B(n1196), .ZN(n1075) );
NOR2_X1 U913 ( .A1(KEYINPUT62), .A2(n1197), .ZN(n1196) );
NOR3_X1 U914 ( .A1(n1164), .A2(n997), .A3(n985), .ZN(n1064) );
INV_X1 U915 ( .A(n1109), .ZN(n985) );
NOR2_X1 U916 ( .A1(n1198), .A2(n988), .ZN(n1109) );
XOR2_X1 U917 ( .A(n1010), .B(KEYINPUT40), .Z(n988) );
XNOR2_X1 U918 ( .A(n1199), .B(G469), .ZN(n1010) );
NAND2_X1 U919 ( .A1(n1200), .A2(n1154), .ZN(n1199) );
XOR2_X1 U920 ( .A(n1201), .B(n1202), .Z(n1200) );
XNOR2_X1 U921 ( .A(n1203), .B(n1092), .ZN(n1202) );
NAND2_X1 U922 ( .A1(G227), .A2(n975), .ZN(n1092) );
NAND2_X1 U923 ( .A1(KEYINPUT22), .A2(n1083), .ZN(n1203) );
XOR2_X1 U924 ( .A(n1204), .B(n1205), .Z(n1083) );
XOR2_X1 U925 ( .A(G107), .B(G104), .Z(n1205) );
XOR2_X1 U926 ( .A(n1206), .B(n1071), .Z(n1204) );
XNOR2_X1 U927 ( .A(n1033), .B(KEYINPUT24), .ZN(n1071) );
XOR2_X1 U928 ( .A(n1207), .B(n1208), .Z(n1033) );
XOR2_X1 U929 ( .A(G137), .B(G131), .Z(n1208) );
XNOR2_X1 U930 ( .A(n1133), .B(n1209), .ZN(n1207) );
XOR2_X1 U931 ( .A(n1090), .B(G140), .Z(n1201) );
XOR2_X1 U932 ( .A(n987), .B(KEYINPUT63), .Z(n1198) );
INV_X1 U933 ( .A(n1166), .ZN(n987) );
NAND2_X1 U934 ( .A1(G221), .A2(n1170), .ZN(n1166) );
NAND2_X1 U935 ( .A1(G234), .A2(n1210), .ZN(n1170) );
XOR2_X1 U936 ( .A(KEYINPUT35), .B(n1211), .Z(n1210) );
INV_X1 U937 ( .A(n1112), .ZN(n997) );
NOR2_X1 U938 ( .A1(n1000), .A2(n999), .ZN(n1112) );
AND2_X1 U939 ( .A1(G214), .A2(n1212), .ZN(n999) );
XOR2_X1 U940 ( .A(n1213), .B(n1023), .Z(n1000) );
INV_X1 U941 ( .A(n1020), .ZN(n1023) );
NAND2_X1 U942 ( .A1(G210), .A2(n1212), .ZN(n1020) );
NAND2_X1 U943 ( .A1(n1211), .A2(n1214), .ZN(n1212) );
INV_X1 U944 ( .A(G237), .ZN(n1214) );
XOR2_X1 U945 ( .A(G902), .B(KEYINPUT49), .Z(n1211) );
XOR2_X1 U946 ( .A(n1021), .B(KEYINPUT15), .Z(n1213) );
NAND2_X1 U947 ( .A1(n1215), .A2(n1154), .ZN(n1021) );
XOR2_X1 U948 ( .A(n1216), .B(KEYINPUT26), .Z(n1215) );
NAND3_X1 U949 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1216) );
OR2_X1 U950 ( .A1(n1131), .A2(KEYINPUT33), .ZN(n1219) );
NAND2_X1 U951 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
NAND2_X1 U952 ( .A1(KEYINPUT33), .A2(n1222), .ZN(n1221) );
XOR2_X1 U953 ( .A(KEYINPUT51), .B(n1131), .Z(n1222) );
NAND3_X1 U954 ( .A1(KEYINPUT33), .A2(n1131), .A3(n1223), .ZN(n1217) );
INV_X1 U955 ( .A(n1220), .ZN(n1223) );
XOR2_X1 U956 ( .A(n1224), .B(n1225), .Z(n1220) );
NOR2_X1 U957 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
NOR2_X1 U958 ( .A1(n1134), .A2(n1228), .ZN(n1227) );
XNOR2_X1 U959 ( .A(n1133), .B(KEYINPUT50), .ZN(n1228) );
INV_X1 U960 ( .A(G125), .ZN(n1134) );
NOR2_X1 U961 ( .A1(G125), .A2(n1229), .ZN(n1226) );
XOR2_X1 U962 ( .A(KEYINPUT46), .B(n1133), .Z(n1229) );
XNOR2_X1 U963 ( .A(n1184), .B(n1230), .ZN(n1133) );
INV_X1 U964 ( .A(G146), .ZN(n1184) );
NAND2_X1 U965 ( .A1(KEYINPUT6), .A2(n1135), .ZN(n1224) );
AND2_X1 U966 ( .A1(G224), .A2(n975), .ZN(n1135) );
INV_X1 U967 ( .A(n1038), .ZN(n1131) );
XOR2_X1 U968 ( .A(n1231), .B(n1232), .Z(n1038) );
XOR2_X1 U969 ( .A(n1233), .B(n1234), .Z(n1232) );
XNOR2_X1 U970 ( .A(n1235), .B(n1236), .ZN(n1234) );
NOR2_X1 U971 ( .A1(KEYINPUT21), .A2(n1165), .ZN(n1236) );
NAND2_X1 U972 ( .A1(KEYINPUT28), .A2(n958), .ZN(n1235) );
INV_X1 U973 ( .A(G107), .ZN(n958) );
XOR2_X1 U974 ( .A(G110), .B(G104), .Z(n1233) );
XOR2_X1 U975 ( .A(n1237), .B(n1238), .Z(n1231) );
INV_X1 U976 ( .A(n1206), .ZN(n1238) );
XNOR2_X1 U977 ( .A(G101), .B(KEYINPUT23), .ZN(n1206) );
XNOR2_X1 U978 ( .A(n1239), .B(n1197), .ZN(n1237) );
XNOR2_X1 U979 ( .A(G116), .B(G119), .ZN(n1197) );
NAND2_X1 U980 ( .A1(KEYINPUT57), .A2(n1156), .ZN(n1239) );
INV_X1 U981 ( .A(G122), .ZN(n1156) );
NAND2_X1 U982 ( .A1(n968), .A2(n1240), .ZN(n1164) );
NAND2_X1 U983 ( .A1(n1241), .A2(n1152), .ZN(n1240) );
NAND2_X1 U984 ( .A1(n1242), .A2(n975), .ZN(n1152) );
XOR2_X1 U985 ( .A(KEYINPUT34), .B(G952), .Z(n1242) );
NAND3_X1 U986 ( .A1(n1243), .A2(n1244), .A3(G902), .ZN(n1241) );
INV_X1 U987 ( .A(G898), .ZN(n1244) );
XOR2_X1 U988 ( .A(KEYINPUT44), .B(G953), .Z(n1243) );
NAND2_X1 U989 ( .A1(G237), .A2(G234), .ZN(n968) );
NOR2_X1 U990 ( .A1(n1124), .A2(n1009), .ZN(n983) );
INV_X1 U991 ( .A(n1140), .ZN(n1009) );
XOR2_X1 U992 ( .A(n1245), .B(G475), .Z(n1140) );
NAND2_X1 U993 ( .A1(n1062), .A2(n1154), .ZN(n1245) );
XNOR2_X1 U994 ( .A(n1246), .B(n1247), .ZN(n1062) );
XNOR2_X1 U995 ( .A(G104), .B(n1248), .ZN(n1247) );
NAND2_X1 U996 ( .A1(n1249), .A2(KEYINPUT41), .ZN(n1248) );
XOR2_X1 U997 ( .A(n1250), .B(n1251), .Z(n1249) );
XOR2_X1 U998 ( .A(G131), .B(n1252), .Z(n1251) );
XOR2_X1 U999 ( .A(G146), .B(G143), .Z(n1252) );
XOR2_X1 U1000 ( .A(n1253), .B(n1254), .Z(n1250) );
NOR2_X1 U1001 ( .A1(KEYINPUT13), .A2(n1091), .ZN(n1254) );
INV_X1 U1002 ( .A(G140), .ZN(n1091) );
XOR2_X1 U1003 ( .A(n1255), .B(G125), .Z(n1253) );
NAND3_X1 U1004 ( .A1(G214), .A2(n1194), .A3(KEYINPUT30), .ZN(n1255) );
NOR2_X1 U1005 ( .A1(G953), .A2(G237), .ZN(n1194) );
XOR2_X1 U1006 ( .A(n1165), .B(n1256), .Z(n1246) );
XOR2_X1 U1007 ( .A(KEYINPUT39), .B(G122), .Z(n1256) );
INV_X1 U1008 ( .A(G113), .ZN(n1165) );
INV_X1 U1009 ( .A(n1141), .ZN(n1124) );
XOR2_X1 U1010 ( .A(n1011), .B(G478), .Z(n1141) );
NAND2_X1 U1011 ( .A1(n1059), .A2(n1154), .ZN(n1011) );
INV_X1 U1012 ( .A(G902), .ZN(n1154) );
XOR2_X1 U1013 ( .A(n1257), .B(n1258), .Z(n1059) );
XOR2_X1 U1014 ( .A(G107), .B(n1259), .Z(n1258) );
XOR2_X1 U1015 ( .A(G122), .B(G116), .Z(n1259) );
XNOR2_X1 U1016 ( .A(n1230), .B(n1260), .ZN(n1257) );
XOR2_X1 U1017 ( .A(n1261), .B(n1209), .Z(n1260) );
XOR2_X1 U1018 ( .A(G134), .B(KEYINPUT55), .Z(n1209) );
NOR2_X1 U1019 ( .A1(n1262), .A2(KEYINPUT0), .ZN(n1261) );
NOR2_X1 U1020 ( .A1(n1263), .A2(n1175), .ZN(n1262) );
NAND2_X1 U1021 ( .A1(G234), .A2(n975), .ZN(n1175) );
INV_X1 U1022 ( .A(G953), .ZN(n975) );
INV_X1 U1023 ( .A(G217), .ZN(n1263) );
XNOR2_X1 U1024 ( .A(n1145), .B(G143), .ZN(n1230) );
INV_X1 U1025 ( .A(G128), .ZN(n1145) );
NAND2_X1 U1026 ( .A1(KEYINPUT52), .A2(n1090), .ZN(n1168) );
INV_X1 U1027 ( .A(G110), .ZN(n1090) );
endmodule


