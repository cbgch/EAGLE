//Key = 1111110000001101000000011000001011111100100110001110001100011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346;

XNOR2_X1 U751 ( .A(G107), .B(n1030), .ZN(G9) );
NAND4_X1 U752 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
NOR2_X1 U753 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U754 ( .A1(KEYINPUT43), .A2(n1037), .ZN(n1032) );
NAND2_X1 U755 ( .A1(n1038), .A2(n1039), .ZN(n1031) );
INV_X1 U756 ( .A(KEYINPUT43), .ZN(n1039) );
NAND2_X1 U757 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U758 ( .A1(n1042), .A2(n1043), .ZN(G75) );
NOR4_X1 U759 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
NOR3_X1 U760 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
XOR2_X1 U761 ( .A(KEYINPUT40), .B(n1051), .Z(n1050) );
NAND3_X1 U762 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1048) );
XNOR2_X1 U763 ( .A(KEYINPUT22), .B(n1055), .ZN(n1053) );
NOR4_X1 U764 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1045) );
NOR2_X1 U765 ( .A1(n1040), .A2(n1060), .ZN(n1058) );
NAND3_X1 U766 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1056) );
OR2_X1 U767 ( .A1(n1033), .A2(n1064), .ZN(n1063) );
NAND3_X1 U768 ( .A1(n1065), .A2(n1036), .A3(n1066), .ZN(n1062) );
NAND2_X1 U769 ( .A1(n1064), .A2(n1067), .ZN(n1066) );
NAND4_X1 U770 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1067) );
NAND2_X1 U771 ( .A1(n1072), .A2(n1055), .ZN(n1061) );
NAND3_X1 U772 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1044) );
NAND3_X1 U773 ( .A1(n1054), .A2(n1052), .A3(n1076), .ZN(n1074) );
INV_X1 U774 ( .A(n1072), .ZN(n1052) );
NAND2_X1 U775 ( .A1(n1064), .A2(n1033), .ZN(n1072) );
INV_X1 U776 ( .A(n1057), .ZN(n1054) );
NOR3_X1 U777 ( .A1(n1077), .A2(G952), .A3(n1046), .ZN(n1042) );
AND4_X1 U778 ( .A1(n1078), .A2(n1064), .A3(n1079), .A4(n1080), .ZN(n1046) );
NOR4_X1 U779 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1080) );
NOR2_X1 U780 ( .A1(n1085), .A2(n1086), .ZN(n1079) );
XOR2_X1 U781 ( .A(n1087), .B(n1088), .Z(n1085) );
XOR2_X1 U782 ( .A(KEYINPUT50), .B(G469), .Z(n1088) );
XOR2_X1 U783 ( .A(n1089), .B(KEYINPUT26), .Z(n1078) );
INV_X1 U784 ( .A(n1073), .ZN(n1077) );
XOR2_X1 U785 ( .A(n1090), .B(n1091), .Z(G72) );
XOR2_X1 U786 ( .A(n1092), .B(n1093), .Z(n1091) );
NOR2_X1 U787 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
XNOR2_X1 U788 ( .A(KEYINPUT41), .B(n1096), .ZN(n1095) );
INV_X1 U789 ( .A(n1097), .ZN(n1094) );
NAND2_X1 U790 ( .A1(n1098), .A2(n1099), .ZN(n1092) );
NAND2_X1 U791 ( .A1(G953), .A2(n1100), .ZN(n1099) );
XOR2_X1 U792 ( .A(n1101), .B(n1102), .Z(n1098) );
XOR2_X1 U793 ( .A(n1103), .B(n1104), .Z(n1102) );
XNOR2_X1 U794 ( .A(n1105), .B(G131), .ZN(n1104) );
XOR2_X1 U795 ( .A(KEYINPUT27), .B(KEYINPUT10), .Z(n1103) );
XOR2_X1 U796 ( .A(n1106), .B(n1107), .Z(n1101) );
XOR2_X1 U797 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U798 ( .A1(KEYINPUT34), .A2(n1110), .ZN(n1108) );
XNOR2_X1 U799 ( .A(G125), .B(n1111), .ZN(n1110) );
NAND2_X1 U800 ( .A1(KEYINPUT2), .A2(n1112), .ZN(n1111) );
NAND2_X1 U801 ( .A1(G953), .A2(n1113), .ZN(n1090) );
NAND2_X1 U802 ( .A1(G900), .A2(G227), .ZN(n1113) );
NAND2_X1 U803 ( .A1(n1114), .A2(n1115), .ZN(G69) );
NAND2_X1 U804 ( .A1(n1116), .A2(n1096), .ZN(n1115) );
XNOR2_X1 U805 ( .A(n1117), .B(n1118), .ZN(n1116) );
NAND2_X1 U806 ( .A1(n1119), .A2(G953), .ZN(n1114) );
NAND2_X1 U807 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U808 ( .A1(n1118), .A2(n1122), .ZN(n1121) );
INV_X1 U809 ( .A(G224), .ZN(n1122) );
NAND2_X1 U810 ( .A1(G224), .A2(n1123), .ZN(n1120) );
NAND2_X1 U811 ( .A1(G898), .A2(n1118), .ZN(n1123) );
NAND2_X1 U812 ( .A1(n1124), .A2(n1125), .ZN(n1118) );
NAND2_X1 U813 ( .A1(G953), .A2(n1126), .ZN(n1125) );
XOR2_X1 U814 ( .A(n1127), .B(n1128), .Z(n1124) );
XNOR2_X1 U815 ( .A(KEYINPUT33), .B(n1129), .ZN(n1127) );
NOR2_X1 U816 ( .A1(KEYINPUT38), .A2(n1130), .ZN(n1129) );
NOR2_X1 U817 ( .A1(n1131), .A2(n1132), .ZN(G66) );
NOR2_X1 U818 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U819 ( .A(n1135), .B(n1136), .Z(n1134) );
NAND2_X1 U820 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U821 ( .A1(KEYINPUT48), .A2(n1139), .ZN(n1135) );
NOR2_X1 U822 ( .A1(KEYINPUT48), .A2(n1139), .ZN(n1133) );
XNOR2_X1 U823 ( .A(n1140), .B(KEYINPUT59), .ZN(n1139) );
NOR2_X1 U824 ( .A1(n1131), .A2(n1141), .ZN(G63) );
XOR2_X1 U825 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND2_X1 U826 ( .A1(n1137), .A2(G478), .ZN(n1142) );
NOR2_X1 U827 ( .A1(n1131), .A2(n1144), .ZN(G60) );
XOR2_X1 U828 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND2_X1 U829 ( .A1(n1137), .A2(G475), .ZN(n1145) );
XOR2_X1 U830 ( .A(n1147), .B(G104), .Z(G6) );
NAND2_X1 U831 ( .A1(KEYINPUT55), .A2(n1148), .ZN(n1147) );
NAND4_X1 U832 ( .A1(n1149), .A2(n1150), .A3(n1033), .A4(n1151), .ZN(n1148) );
NOR2_X1 U833 ( .A1(n1131), .A2(n1152), .ZN(G57) );
XOR2_X1 U834 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U835 ( .A1(n1155), .A2(KEYINPUT44), .ZN(n1153) );
XNOR2_X1 U836 ( .A(n1156), .B(n1157), .ZN(n1155) );
XOR2_X1 U837 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND2_X1 U838 ( .A1(n1137), .A2(G472), .ZN(n1158) );
NOR2_X1 U839 ( .A1(n1131), .A2(n1160), .ZN(G54) );
XOR2_X1 U840 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U841 ( .A(n1163), .B(n1106), .ZN(n1162) );
XNOR2_X1 U842 ( .A(n1164), .B(n1165), .ZN(n1161) );
XOR2_X1 U843 ( .A(n1166), .B(n1167), .Z(n1165) );
NAND2_X1 U844 ( .A1(n1137), .A2(G469), .ZN(n1167) );
NAND2_X1 U845 ( .A1(n1168), .A2(KEYINPUT49), .ZN(n1166) );
XOR2_X1 U846 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U847 ( .A1(KEYINPUT8), .A2(n1171), .ZN(n1170) );
XOR2_X1 U848 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U849 ( .A1(KEYINPUT47), .A2(G110), .ZN(n1173) );
XNOR2_X1 U850 ( .A(G140), .B(KEYINPUT4), .ZN(n1172) );
NOR2_X1 U851 ( .A1(n1131), .A2(n1174), .ZN(G51) );
XOR2_X1 U852 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U853 ( .A(n1177), .B(n1178), .Z(n1176) );
NAND2_X1 U854 ( .A1(n1137), .A2(n1179), .ZN(n1177) );
NOR2_X1 U855 ( .A1(n1180), .A2(n1075), .ZN(n1137) );
NOR2_X1 U856 ( .A1(n1097), .A2(n1117), .ZN(n1075) );
NAND4_X1 U857 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1117) );
AND4_X1 U858 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1184) );
NAND2_X1 U859 ( .A1(n1189), .A2(n1190), .ZN(n1183) );
XOR2_X1 U860 ( .A(n1191), .B(KEYINPUT1), .Z(n1189) );
NAND4_X1 U861 ( .A1(n1150), .A2(n1033), .A3(n1192), .A4(n1193), .ZN(n1181) );
NAND2_X1 U862 ( .A1(n1035), .A2(n1194), .ZN(n1193) );
NAND2_X1 U863 ( .A1(KEYINPUT31), .A2(n1149), .ZN(n1194) );
INV_X1 U864 ( .A(n1151), .ZN(n1035) );
NAND3_X1 U865 ( .A1(n1195), .A2(n1036), .A3(n1151), .ZN(n1192) );
OR2_X1 U866 ( .A1(n1065), .A2(KEYINPUT31), .ZN(n1195) );
NAND4_X1 U867 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1097) );
NOR4_X1 U868 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
NOR2_X1 U869 ( .A1(n1204), .A2(n1205), .ZN(n1198) );
NOR4_X1 U870 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1205) );
XNOR2_X1 U871 ( .A(n1064), .B(KEYINPUT63), .ZN(n1208) );
INV_X1 U872 ( .A(n1210), .ZN(n1204) );
NAND4_X1 U873 ( .A1(n1076), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1197) );
OR2_X1 U874 ( .A1(n1214), .A2(KEYINPUT18), .ZN(n1213) );
NAND2_X1 U875 ( .A1(KEYINPUT18), .A2(n1215), .ZN(n1212) );
NAND2_X1 U876 ( .A1(n1149), .A2(n1068), .ZN(n1215) );
NAND3_X1 U877 ( .A1(n1216), .A2(n1217), .A3(n1214), .ZN(n1196) );
NAND2_X1 U878 ( .A1(KEYINPUT30), .A2(n1209), .ZN(n1217) );
NAND2_X1 U879 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
INV_X1 U880 ( .A(KEYINPUT30), .ZN(n1219) );
NAND3_X1 U881 ( .A1(n1040), .A2(n1220), .A3(n1221), .ZN(n1218) );
XOR2_X1 U882 ( .A(KEYINPUT54), .B(n1222), .Z(n1175) );
NOR3_X1 U883 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1222) );
AND2_X1 U884 ( .A1(n1226), .A2(KEYINPUT17), .ZN(n1225) );
NOR3_X1 U885 ( .A1(KEYINPUT17), .A2(G125), .A3(n1227), .ZN(n1224) );
INV_X1 U886 ( .A(n1228), .ZN(n1227) );
NOR2_X1 U887 ( .A1(n1228), .A2(n1229), .ZN(n1223) );
NOR2_X1 U888 ( .A1(KEYINPUT58), .A2(n1226), .ZN(n1228) );
XNOR2_X1 U889 ( .A(n1230), .B(KEYINPUT62), .ZN(n1226) );
NOR2_X1 U890 ( .A1(n1231), .A2(G952), .ZN(n1131) );
XNOR2_X1 U891 ( .A(n1096), .B(KEYINPUT35), .ZN(n1231) );
INV_X1 U892 ( .A(G953), .ZN(n1096) );
XOR2_X1 U893 ( .A(G146), .B(n1203), .Z(G48) );
AND2_X1 U894 ( .A1(n1149), .A2(n1232), .ZN(n1203) );
XNOR2_X1 U895 ( .A(G143), .B(n1210), .ZN(G45) );
NAND3_X1 U896 ( .A1(n1150), .A2(n1233), .A3(n1234), .ZN(n1210) );
NOR3_X1 U897 ( .A1(n1235), .A2(n1221), .A3(n1236), .ZN(n1234) );
XNOR2_X1 U898 ( .A(G140), .B(n1237), .ZN(G42) );
NAND2_X1 U899 ( .A1(n1214), .A2(n1238), .ZN(n1237) );
XNOR2_X1 U900 ( .A(n1105), .B(n1239), .ZN(G39) );
AND2_X1 U901 ( .A1(n1238), .A2(n1240), .ZN(n1239) );
XNOR2_X1 U902 ( .A(G134), .B(n1241), .ZN(G36) );
NOR2_X1 U903 ( .A1(n1202), .A2(KEYINPUT51), .ZN(n1241) );
NOR3_X1 U904 ( .A1(n1036), .A2(n1069), .A3(n1209), .ZN(n1202) );
INV_X1 U905 ( .A(n1242), .ZN(n1036) );
XNOR2_X1 U906 ( .A(n1201), .B(n1243), .ZN(G33) );
NAND2_X1 U907 ( .A1(KEYINPUT36), .A2(G131), .ZN(n1243) );
NOR3_X1 U908 ( .A1(n1065), .A2(n1069), .A3(n1209), .ZN(n1201) );
INV_X1 U909 ( .A(n1238), .ZN(n1209) );
NOR3_X1 U910 ( .A1(n1059), .A2(n1221), .A3(n1071), .ZN(n1238) );
INV_X1 U911 ( .A(n1040), .ZN(n1071) );
INV_X1 U912 ( .A(n1220), .ZN(n1059) );
NAND2_X1 U913 ( .A1(n1244), .A2(n1245), .ZN(n1220) );
OR2_X1 U914 ( .A1(n1041), .A2(KEYINPUT40), .ZN(n1245) );
NAND3_X1 U915 ( .A1(n1051), .A2(n1049), .A3(KEYINPUT40), .ZN(n1244) );
INV_X1 U916 ( .A(n1233), .ZN(n1069) );
XOR2_X1 U917 ( .A(G128), .B(n1200), .Z(G30) );
AND2_X1 U918 ( .A1(n1232), .A2(n1242), .ZN(n1200) );
NOR4_X1 U919 ( .A1(n1037), .A2(n1207), .A3(n1206), .A4(n1221), .ZN(n1232) );
INV_X1 U920 ( .A(n1211), .ZN(n1221) );
XOR2_X1 U921 ( .A(G101), .B(n1246), .Z(G3) );
NOR2_X1 U922 ( .A1(n1041), .A2(n1191), .ZN(n1246) );
NAND4_X1 U923 ( .A1(n1064), .A2(n1040), .A3(n1233), .A4(n1151), .ZN(n1191) );
XNOR2_X1 U924 ( .A(G125), .B(n1247), .ZN(G27) );
NAND3_X1 U925 ( .A1(n1076), .A2(n1211), .A3(n1214), .ZN(n1247) );
NOR2_X1 U926 ( .A1(n1065), .A2(n1068), .ZN(n1214) );
INV_X1 U927 ( .A(n1248), .ZN(n1068) );
INV_X1 U928 ( .A(n1149), .ZN(n1065) );
NAND2_X1 U929 ( .A1(n1057), .A2(n1249), .ZN(n1211) );
NAND4_X1 U930 ( .A1(G902), .A2(G953), .A3(n1250), .A4(n1100), .ZN(n1249) );
INV_X1 U931 ( .A(G900), .ZN(n1100) );
XOR2_X1 U932 ( .A(n1182), .B(n1251), .Z(G24) );
XNOR2_X1 U933 ( .A(G122), .B(KEYINPUT56), .ZN(n1251) );
NAND4_X1 U934 ( .A1(n1252), .A2(n1033), .A3(n1253), .A4(n1254), .ZN(n1182) );
XNOR2_X1 U935 ( .A(G119), .B(n1188), .ZN(G21) );
NAND2_X1 U936 ( .A1(n1240), .A2(n1252), .ZN(n1188) );
NOR3_X1 U937 ( .A1(n1207), .A2(n1206), .A3(n1255), .ZN(n1240) );
INV_X1 U938 ( .A(n1064), .ZN(n1255) );
XNOR2_X1 U939 ( .A(n1256), .B(KEYINPUT39), .ZN(n1207) );
XNOR2_X1 U940 ( .A(G116), .B(n1187), .ZN(G18) );
NAND3_X1 U941 ( .A1(n1242), .A2(n1233), .A3(n1252), .ZN(n1187) );
NOR2_X1 U942 ( .A1(n1254), .A2(n1235), .ZN(n1242) );
INV_X1 U943 ( .A(n1253), .ZN(n1235) );
XNOR2_X1 U944 ( .A(G113), .B(n1186), .ZN(G15) );
NAND3_X1 U945 ( .A1(n1149), .A2(n1233), .A3(n1252), .ZN(n1186) );
AND2_X1 U946 ( .A1(n1076), .A2(n1151), .ZN(n1252) );
NOR2_X1 U947 ( .A1(n1055), .A2(n1041), .ZN(n1076) );
INV_X1 U948 ( .A(n1190), .ZN(n1041) );
NAND2_X1 U949 ( .A1(n1060), .A2(n1070), .ZN(n1055) );
NAND2_X1 U950 ( .A1(n1257), .A2(n1258), .ZN(n1233) );
OR3_X1 U951 ( .A1(n1259), .A2(n1086), .A3(KEYINPUT39), .ZN(n1258) );
INV_X1 U952 ( .A(n1256), .ZN(n1259) );
NAND2_X1 U953 ( .A1(KEYINPUT39), .A2(n1033), .ZN(n1257) );
NOR2_X1 U954 ( .A1(n1253), .A2(n1236), .ZN(n1149) );
INV_X1 U955 ( .A(n1254), .ZN(n1236) );
XNOR2_X1 U956 ( .A(G110), .B(n1185), .ZN(G12) );
NAND4_X1 U957 ( .A1(n1150), .A2(n1064), .A3(n1248), .A4(n1151), .ZN(n1185) );
NAND2_X1 U958 ( .A1(n1057), .A2(n1260), .ZN(n1151) );
NAND4_X1 U959 ( .A1(G902), .A2(G953), .A3(n1250), .A4(n1126), .ZN(n1260) );
INV_X1 U960 ( .A(G898), .ZN(n1126) );
NAND3_X1 U961 ( .A1(n1073), .A2(n1250), .A3(G952), .ZN(n1057) );
NAND2_X1 U962 ( .A1(G237), .A2(G234), .ZN(n1250) );
XOR2_X1 U963 ( .A(G953), .B(KEYINPUT13), .Z(n1073) );
NAND2_X1 U964 ( .A1(n1261), .A2(n1262), .ZN(n1248) );
OR3_X1 U965 ( .A1(n1206), .A2(n1256), .A3(KEYINPUT29), .ZN(n1262) );
INV_X1 U966 ( .A(n1086), .ZN(n1206) );
NAND2_X1 U967 ( .A1(KEYINPUT29), .A2(n1033), .ZN(n1261) );
NOR2_X1 U968 ( .A1(n1086), .A2(n1256), .ZN(n1033) );
XNOR2_X1 U969 ( .A(n1089), .B(KEYINPUT20), .ZN(n1256) );
XOR2_X1 U970 ( .A(n1263), .B(G472), .Z(n1089) );
NAND2_X1 U971 ( .A1(n1264), .A2(n1180), .ZN(n1263) );
XOR2_X1 U972 ( .A(n1154), .B(n1265), .Z(n1264) );
XOR2_X1 U973 ( .A(n1266), .B(KEYINPUT9), .Z(n1265) );
NAND2_X1 U974 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
OR2_X1 U975 ( .A1(n1156), .A2(n1269), .ZN(n1268) );
XOR2_X1 U976 ( .A(n1270), .B(KEYINPUT11), .Z(n1267) );
NAND2_X1 U977 ( .A1(n1269), .A2(n1156), .ZN(n1270) );
XNOR2_X1 U978 ( .A(n1271), .B(n1272), .ZN(n1156) );
NAND2_X1 U979 ( .A1(KEYINPUT24), .A2(G116), .ZN(n1271) );
XNOR2_X1 U980 ( .A(n1159), .B(KEYINPUT7), .ZN(n1269) );
XNOR2_X1 U981 ( .A(n1273), .B(n1274), .ZN(n1159) );
XNOR2_X1 U982 ( .A(n1230), .B(KEYINPUT46), .ZN(n1273) );
XOR2_X1 U983 ( .A(n1275), .B(G101), .Z(n1154) );
NAND2_X1 U984 ( .A1(G210), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U985 ( .A(n1277), .B(n1138), .ZN(n1086) );
AND2_X1 U986 ( .A1(G217), .A2(n1278), .ZN(n1138) );
NAND2_X1 U987 ( .A1(n1140), .A2(n1180), .ZN(n1277) );
XNOR2_X1 U988 ( .A(n1279), .B(n1280), .ZN(n1140) );
XOR2_X1 U989 ( .A(G110), .B(n1281), .Z(n1280) );
XOR2_X1 U990 ( .A(G128), .B(G119), .Z(n1281) );
XOR2_X1 U991 ( .A(n1282), .B(n1283), .Z(n1279) );
NOR2_X1 U992 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U993 ( .A(KEYINPUT42), .B(n1286), .Z(n1285) );
NOR2_X1 U994 ( .A1(n1287), .A2(n1105), .ZN(n1286) );
AND2_X1 U995 ( .A1(n1105), .A2(n1287), .ZN(n1284) );
NAND3_X1 U996 ( .A1(n1288), .A2(n1289), .A3(G221), .ZN(n1287) );
INV_X1 U997 ( .A(G137), .ZN(n1105) );
NAND2_X1 U998 ( .A1(KEYINPUT37), .A2(n1290), .ZN(n1282) );
NOR2_X1 U999 ( .A1(n1253), .A2(n1254), .ZN(n1064) );
XNOR2_X1 U1000 ( .A(n1291), .B(G475), .ZN(n1254) );
NAND2_X1 U1001 ( .A1(n1146), .A2(n1180), .ZN(n1291) );
XOR2_X1 U1002 ( .A(n1292), .B(n1293), .Z(n1146) );
XOR2_X1 U1003 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U1004 ( .A(n1296), .B(n1297), .ZN(n1295) );
NAND2_X1 U1005 ( .A1(KEYINPUT5), .A2(n1298), .ZN(n1297) );
INV_X1 U1006 ( .A(n1290), .ZN(n1298) );
XOR2_X1 U1007 ( .A(G125), .B(n1299), .Z(n1290) );
XNOR2_X1 U1008 ( .A(G146), .B(n1112), .ZN(n1299) );
NAND2_X1 U1009 ( .A1(KEYINPUT0), .A2(G104), .ZN(n1296) );
NAND2_X1 U1010 ( .A1(G214), .A2(n1276), .ZN(n1294) );
AND2_X1 U1011 ( .A1(n1289), .A2(n1300), .ZN(n1276) );
XOR2_X1 U1012 ( .A(n1301), .B(n1302), .Z(n1292) );
XNOR2_X1 U1013 ( .A(n1303), .B(G131), .ZN(n1302) );
XNOR2_X1 U1014 ( .A(G113), .B(G122), .ZN(n1301) );
XNOR2_X1 U1015 ( .A(n1304), .B(G478), .ZN(n1253) );
NAND2_X1 U1016 ( .A1(n1143), .A2(n1180), .ZN(n1304) );
XNOR2_X1 U1017 ( .A(n1305), .B(n1306), .ZN(n1143) );
XOR2_X1 U1018 ( .A(G107), .B(n1307), .Z(n1306) );
NOR2_X1 U1019 ( .A1(KEYINPUT61), .A2(n1308), .ZN(n1307) );
XNOR2_X1 U1020 ( .A(G116), .B(G122), .ZN(n1308) );
XOR2_X1 U1021 ( .A(n1309), .B(n1310), .Z(n1305) );
NOR2_X1 U1022 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U1023 ( .A(n1313), .B(KEYINPUT60), .Z(n1312) );
NAND2_X1 U1024 ( .A1(G134), .A2(n1314), .ZN(n1313) );
NOR2_X1 U1025 ( .A1(G134), .A2(n1314), .ZN(n1311) );
XNOR2_X1 U1026 ( .A(n1303), .B(G128), .ZN(n1314) );
INV_X1 U1027 ( .A(G143), .ZN(n1303) );
NAND3_X1 U1028 ( .A1(n1288), .A2(G217), .A3(n1289), .ZN(n1309) );
XNOR2_X1 U1029 ( .A(G234), .B(KEYINPUT23), .ZN(n1288) );
INV_X1 U1030 ( .A(n1037), .ZN(n1150) );
NAND2_X1 U1031 ( .A1(n1190), .A2(n1040), .ZN(n1037) );
NOR2_X1 U1032 ( .A1(n1060), .A2(n1084), .ZN(n1040) );
INV_X1 U1033 ( .A(n1070), .ZN(n1084) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1278), .ZN(n1070) );
NAND2_X1 U1035 ( .A1(G234), .A2(n1180), .ZN(n1278) );
XNOR2_X1 U1036 ( .A(n1315), .B(G469), .ZN(n1060) );
NAND2_X1 U1037 ( .A1(KEYINPUT15), .A2(n1087), .ZN(n1315) );
NAND2_X1 U1038 ( .A1(n1316), .A2(n1180), .ZN(n1087) );
XOR2_X1 U1039 ( .A(n1317), .B(n1318), .Z(n1316) );
XNOR2_X1 U1040 ( .A(n1319), .B(n1274), .ZN(n1318) );
INV_X1 U1041 ( .A(n1164), .ZN(n1274) );
XOR2_X1 U1042 ( .A(G131), .B(n1320), .Z(n1164) );
NOR2_X1 U1043 ( .A1(KEYINPUT14), .A2(n1321), .ZN(n1320) );
XNOR2_X1 U1044 ( .A(G137), .B(n1322), .ZN(n1321) );
NOR2_X1 U1045 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
AND2_X1 U1046 ( .A1(KEYINPUT6), .A2(n1109), .ZN(n1324) );
NOR2_X1 U1047 ( .A1(KEYINPUT53), .A2(n1109), .ZN(n1323) );
XNOR2_X1 U1048 ( .A(G134), .B(KEYINPUT12), .ZN(n1109) );
NOR3_X1 U1049 ( .A1(n1325), .A2(KEYINPUT16), .A3(n1326), .ZN(n1319) );
AND2_X1 U1050 ( .A1(n1163), .A2(n1106), .ZN(n1326) );
XOR2_X1 U1051 ( .A(KEYINPUT52), .B(n1327), .Z(n1325) );
NOR2_X1 U1052 ( .A1(n1106), .A2(n1163), .ZN(n1327) );
XOR2_X1 U1053 ( .A(n1328), .B(n1329), .Z(n1163) );
NOR2_X1 U1054 ( .A1(G104), .A2(KEYINPUT19), .ZN(n1329) );
XOR2_X1 U1055 ( .A(G128), .B(n1330), .Z(n1106) );
XNOR2_X1 U1056 ( .A(n1169), .B(n1331), .ZN(n1317) );
XNOR2_X1 U1057 ( .A(n1112), .B(G110), .ZN(n1331) );
INV_X1 U1058 ( .A(G140), .ZN(n1112) );
NAND2_X1 U1059 ( .A1(G227), .A2(n1289), .ZN(n1169) );
NOR2_X1 U1060 ( .A1(n1082), .A2(n1051), .ZN(n1190) );
NOR2_X1 U1061 ( .A1(n1332), .A2(n1083), .ZN(n1051) );
NOR2_X1 U1062 ( .A1(n1333), .A2(n1179), .ZN(n1083) );
XOR2_X1 U1063 ( .A(n1081), .B(KEYINPUT28), .Z(n1332) );
AND2_X1 U1064 ( .A1(n1179), .A2(n1333), .ZN(n1081) );
NAND2_X1 U1065 ( .A1(n1334), .A2(n1180), .ZN(n1333) );
XOR2_X1 U1066 ( .A(n1335), .B(n1336), .Z(n1334) );
XNOR2_X1 U1067 ( .A(KEYINPUT3), .B(n1229), .ZN(n1336) );
INV_X1 U1068 ( .A(G125), .ZN(n1229) );
XNOR2_X1 U1069 ( .A(n1178), .B(n1337), .ZN(n1335) );
INV_X1 U1070 ( .A(n1230), .ZN(n1337) );
XOR2_X1 U1071 ( .A(G128), .B(n1338), .Z(n1230) );
NOR2_X1 U1072 ( .A1(KEYINPUT57), .A2(n1330), .ZN(n1338) );
XNOR2_X1 U1073 ( .A(G146), .B(G143), .ZN(n1330) );
XNOR2_X1 U1074 ( .A(n1128), .B(n1339), .ZN(n1178) );
XNOR2_X1 U1075 ( .A(n1340), .B(n1130), .ZN(n1339) );
XNOR2_X1 U1076 ( .A(n1341), .B(n1342), .ZN(n1130) );
XOR2_X1 U1077 ( .A(G122), .B(G110), .Z(n1342) );
XNOR2_X1 U1078 ( .A(KEYINPUT45), .B(KEYINPUT32), .ZN(n1341) );
NAND2_X1 U1079 ( .A1(G224), .A2(n1289), .ZN(n1340) );
XNOR2_X1 U1080 ( .A(G953), .B(KEYINPUT25), .ZN(n1289) );
XNOR2_X1 U1081 ( .A(n1343), .B(n1344), .ZN(n1128) );
XOR2_X1 U1082 ( .A(n1272), .B(n1328), .Z(n1344) );
XOR2_X1 U1083 ( .A(G101), .B(G107), .Z(n1328) );
XOR2_X1 U1084 ( .A(G113), .B(G119), .Z(n1272) );
XNOR2_X1 U1085 ( .A(G104), .B(n1345), .ZN(n1343) );
NOR2_X1 U1086 ( .A1(G116), .A2(KEYINPUT21), .ZN(n1345) );
AND2_X1 U1087 ( .A1(G210), .A2(n1346), .ZN(n1179) );
INV_X1 U1088 ( .A(n1049), .ZN(n1082) );
NAND2_X1 U1089 ( .A1(G214), .A2(n1346), .ZN(n1049) );
NAND2_X1 U1090 ( .A1(n1300), .A2(n1180), .ZN(n1346) );
INV_X1 U1091 ( .A(G902), .ZN(n1180) );
INV_X1 U1092 ( .A(G237), .ZN(n1300) );
endmodule


