//Key = 0011111010110011100000110000110010101100111100100001000100100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326;

XNOR2_X1 U729 ( .A(G107), .B(n1010), .ZN(G9) );
NAND2_X1 U730 ( .A1(KEYINPUT23), .A2(n1011), .ZN(n1010) );
INV_X1 U731 ( .A(n1012), .ZN(n1011) );
NOR2_X1 U732 ( .A1(n1013), .A2(n1014), .ZN(G75) );
NOR4_X1 U733 ( .A1(n1015), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(n1014) );
NOR2_X1 U734 ( .A1(n1019), .A2(n1020), .ZN(n1016) );
NOR2_X1 U735 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR4_X1 U736 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1022) );
NOR3_X1 U737 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1023) );
AND2_X1 U738 ( .A1(n1030), .A2(KEYINPUT53), .ZN(n1027) );
NOR2_X1 U739 ( .A1(n1031), .A2(n1032), .ZN(n1021) );
INV_X1 U740 ( .A(n1033), .ZN(n1032) );
NOR2_X1 U741 ( .A1(n1034), .A2(n1035), .ZN(n1031) );
NOR2_X1 U742 ( .A1(n1036), .A2(n1025), .ZN(n1035) );
INV_X1 U743 ( .A(n1037), .ZN(n1025) );
NOR2_X1 U744 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U745 ( .A1(n1040), .A2(n1024), .ZN(n1039) );
NOR2_X1 U746 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR3_X1 U747 ( .A1(n1043), .A2(KEYINPUT53), .A3(n1044), .ZN(n1041) );
NOR2_X1 U748 ( .A1(n1045), .A2(n1026), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U750 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR3_X1 U751 ( .A1(n1026), .A2(n1050), .A3(n1024), .ZN(n1034) );
NOR2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U753 ( .A1(n1017), .A2(G952), .A3(n1015), .ZN(n1013) );
AND4_X1 U754 ( .A1(n1037), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1015) );
NOR3_X1 U755 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
XOR2_X1 U756 ( .A(n1059), .B(n1060), .Z(n1054) );
INV_X1 U757 ( .A(n1061), .ZN(n1017) );
XOR2_X1 U758 ( .A(n1062), .B(n1063), .Z(G72) );
NOR2_X1 U759 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
AND2_X1 U760 ( .A1(G227), .A2(G900), .ZN(n1064) );
NAND2_X1 U761 ( .A1(n1066), .A2(n1067), .ZN(n1062) );
NAND3_X1 U762 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
NAND2_X1 U763 ( .A1(G953), .A2(n1071), .ZN(n1069) );
OR2_X1 U764 ( .A1(n1068), .A2(n1070), .ZN(n1066) );
NAND2_X1 U765 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NAND4_X1 U766 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1073) );
NOR2_X1 U767 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
INV_X1 U768 ( .A(n1080), .ZN(n1078) );
XOR2_X1 U769 ( .A(n1081), .B(n1082), .Z(n1068) );
XNOR2_X1 U770 ( .A(n1083), .B(n1084), .ZN(n1082) );
NOR2_X1 U771 ( .A1(KEYINPUT47), .A2(n1085), .ZN(n1084) );
XNOR2_X1 U772 ( .A(n1086), .B(n1087), .ZN(n1085) );
NAND2_X1 U773 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U774 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U775 ( .A(KEYINPUT29), .B(n1092), .Z(n1090) );
NAND2_X1 U776 ( .A1(n1092), .A2(G137), .ZN(n1088) );
NAND2_X1 U777 ( .A1(KEYINPUT10), .A2(n1093), .ZN(n1081) );
XOR2_X1 U778 ( .A(n1094), .B(n1095), .Z(G69) );
NOR2_X1 U779 ( .A1(n1096), .A2(n1065), .ZN(n1095) );
XNOR2_X1 U780 ( .A(n1072), .B(KEYINPUT4), .ZN(n1065) );
NOR2_X1 U781 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND3_X1 U782 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1094) );
NAND2_X1 U783 ( .A1(KEYINPUT56), .A2(n1102), .ZN(n1101) );
OR3_X1 U784 ( .A1(n1102), .A2(KEYINPUT56), .A3(n1103), .ZN(n1100) );
OR2_X1 U785 ( .A1(G953), .A2(n1104), .ZN(n1102) );
NAND2_X1 U786 ( .A1(n1103), .A2(n1105), .ZN(n1099) );
NAND2_X1 U787 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U788 ( .A1(G898), .A2(G953), .ZN(n1107) );
NAND2_X1 U789 ( .A1(n1104), .A2(n1072), .ZN(n1106) );
XNOR2_X1 U790 ( .A(n1108), .B(n1109), .ZN(n1103) );
XNOR2_X1 U791 ( .A(n1110), .B(n1111), .ZN(n1108) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(G66) );
XOR2_X1 U793 ( .A(KEYINPUT38), .B(n1114), .Z(n1113) );
XOR2_X1 U794 ( .A(n1115), .B(n1116), .Z(n1112) );
NAND3_X1 U795 ( .A1(n1117), .A2(n1118), .A3(KEYINPUT32), .ZN(n1115) );
NOR3_X1 U796 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(G63) );
AND2_X1 U797 ( .A1(KEYINPUT61), .A2(n1114), .ZN(n1121) );
NOR3_X1 U798 ( .A1(KEYINPUT61), .A2(G953), .A3(G952), .ZN(n1120) );
NOR2_X1 U799 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
XOR2_X1 U800 ( .A(n1124), .B(n1125), .Z(n1123) );
AND2_X1 U801 ( .A1(G478), .A2(n1117), .ZN(n1125) );
AND2_X1 U802 ( .A1(n1126), .A2(KEYINPUT43), .ZN(n1124) );
NOR2_X1 U803 ( .A1(KEYINPUT43), .A2(n1126), .ZN(n1122) );
NOR2_X1 U804 ( .A1(n1114), .A2(n1127), .ZN(G60) );
XOR2_X1 U805 ( .A(n1128), .B(n1129), .Z(n1127) );
AND2_X1 U806 ( .A1(G475), .A2(n1117), .ZN(n1128) );
XOR2_X1 U807 ( .A(G104), .B(n1130), .Z(G6) );
NOR2_X1 U808 ( .A1(n1131), .A2(n1132), .ZN(G57) );
XOR2_X1 U809 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U810 ( .A(KEYINPUT11), .B(n1135), .Z(n1134) );
AND2_X1 U811 ( .A1(G472), .A2(n1117), .ZN(n1135) );
NOR2_X1 U812 ( .A1(G952), .A2(n1136), .ZN(n1131) );
XNOR2_X1 U813 ( .A(G953), .B(KEYINPUT44), .ZN(n1136) );
NOR2_X1 U814 ( .A1(n1114), .A2(n1137), .ZN(G54) );
XOR2_X1 U815 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U816 ( .A(n1110), .B(n1140), .Z(n1139) );
XOR2_X1 U817 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U818 ( .A1(KEYINPUT2), .A2(n1086), .ZN(n1141) );
XOR2_X1 U819 ( .A(n1143), .B(n1144), .Z(n1138) );
XNOR2_X1 U820 ( .A(n1093), .B(G110), .ZN(n1144) );
XOR2_X1 U821 ( .A(n1145), .B(n1146), .Z(n1143) );
AND2_X1 U822 ( .A1(G469), .A2(n1117), .ZN(n1146) );
INV_X1 U823 ( .A(n1147), .ZN(n1117) );
NOR2_X1 U824 ( .A1(n1114), .A2(n1148), .ZN(G51) );
XOR2_X1 U825 ( .A(n1149), .B(n1150), .Z(n1148) );
XNOR2_X1 U826 ( .A(n1151), .B(n1152), .ZN(n1150) );
XNOR2_X1 U827 ( .A(KEYINPUT12), .B(n1153), .ZN(n1152) );
NOR2_X1 U828 ( .A1(KEYINPUT33), .A2(n1154), .ZN(n1153) );
XOR2_X1 U829 ( .A(KEYINPUT27), .B(n1155), .Z(n1154) );
XOR2_X1 U830 ( .A(n1156), .B(n1157), .Z(n1149) );
XOR2_X1 U831 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U832 ( .A1(n1060), .A2(n1147), .ZN(n1158) );
NAND2_X1 U833 ( .A1(n1160), .A2(n1018), .ZN(n1147) );
NAND4_X1 U834 ( .A1(n1104), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1018) );
AND3_X1 U835 ( .A1(n1080), .A2(n1075), .A3(n1074), .ZN(n1163) );
NAND2_X1 U836 ( .A1(n1164), .A2(n1165), .ZN(n1080) );
XNOR2_X1 U837 ( .A(KEYINPUT7), .B(n1166), .ZN(n1165) );
XOR2_X1 U838 ( .A(n1079), .B(KEYINPUT5), .Z(n1162) );
NAND3_X1 U839 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1079) );
NAND2_X1 U840 ( .A1(n1051), .A2(n1170), .ZN(n1169) );
NAND2_X1 U841 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND3_X1 U842 ( .A1(n1173), .A2(n1056), .A3(n1174), .ZN(n1172) );
NOR3_X1 U843 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1174) );
NOR2_X1 U844 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
INV_X1 U845 ( .A(KEYINPUT20), .ZN(n1179) );
NOR2_X1 U846 ( .A1(n1180), .A2(n1181), .ZN(n1178) );
NOR2_X1 U847 ( .A1(KEYINPUT20), .A2(n1182), .ZN(n1176) );
NAND3_X1 U848 ( .A1(n1182), .A2(n1029), .A3(n1164), .ZN(n1171) );
XNOR2_X1 U849 ( .A(KEYINPUT40), .B(n1076), .ZN(n1161) );
AND4_X1 U850 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1104) );
AND4_X1 U851 ( .A1(n1187), .A2(n1012), .A3(n1188), .A4(n1189), .ZN(n1186) );
NAND3_X1 U852 ( .A1(n1190), .A2(n1033), .A3(n1051), .ZN(n1012) );
NOR2_X1 U853 ( .A1(n1130), .A2(n1191), .ZN(n1185) );
NOR2_X1 U854 ( .A1(n1175), .A2(n1192), .ZN(n1191) );
AND4_X1 U855 ( .A1(n1193), .A2(n1033), .A3(n1047), .A4(n1194), .ZN(n1130) );
XNOR2_X1 U856 ( .A(G902), .B(KEYINPUT58), .ZN(n1160) );
NOR2_X1 U857 ( .A1(n1072), .A2(G952), .ZN(n1114) );
XNOR2_X1 U858 ( .A(G146), .B(n1076), .ZN(G48) );
NAND2_X1 U859 ( .A1(n1195), .A2(n1193), .ZN(n1076) );
XNOR2_X1 U860 ( .A(G143), .B(n1074), .ZN(G45) );
NAND4_X1 U861 ( .A1(n1182), .A2(n1196), .A3(n1029), .A4(n1042), .ZN(n1074) );
XNOR2_X1 U862 ( .A(n1093), .B(n1197), .ZN(G42) );
NOR2_X1 U863 ( .A1(n1026), .A2(n1166), .ZN(n1197) );
NAND3_X1 U864 ( .A1(n1052), .A2(n1028), .A3(n1182), .ZN(n1166) );
XNOR2_X1 U865 ( .A(n1075), .B(n1198), .ZN(G39) );
NOR2_X1 U866 ( .A1(KEYINPUT52), .A2(n1091), .ZN(n1198) );
INV_X1 U867 ( .A(G137), .ZN(n1091) );
NAND3_X1 U868 ( .A1(n1195), .A2(n1037), .A3(n1164), .ZN(n1075) );
XOR2_X1 U869 ( .A(n1199), .B(n1200), .Z(G36) );
NOR3_X1 U870 ( .A1(n1201), .A2(n1026), .A3(n1202), .ZN(n1200) );
XNOR2_X1 U871 ( .A(KEYINPUT16), .B(n1180), .ZN(n1202) );
INV_X1 U872 ( .A(n1164), .ZN(n1026) );
NAND3_X1 U873 ( .A1(n1051), .A2(n1181), .A3(n1029), .ZN(n1201) );
XNOR2_X1 U874 ( .A(G134), .B(KEYINPUT42), .ZN(n1199) );
XOR2_X1 U875 ( .A(n1167), .B(n1203), .Z(G33) );
NAND2_X1 U876 ( .A1(KEYINPUT37), .A2(G131), .ZN(n1203) );
NAND4_X1 U877 ( .A1(n1164), .A2(n1182), .A3(n1052), .A4(n1029), .ZN(n1167) );
NOR2_X1 U878 ( .A1(n1044), .A2(n1057), .ZN(n1164) );
INV_X1 U879 ( .A(n1043), .ZN(n1057) );
XNOR2_X1 U880 ( .A(G128), .B(n1204), .ZN(G30) );
NAND3_X1 U881 ( .A1(n1195), .A2(n1051), .A3(n1205), .ZN(n1204) );
XNOR2_X1 U882 ( .A(n1042), .B(KEYINPUT3), .ZN(n1205) );
AND3_X1 U883 ( .A1(n1173), .A2(n1056), .A3(n1182), .ZN(n1195) );
AND2_X1 U884 ( .A1(n1047), .A2(n1181), .ZN(n1182) );
XNOR2_X1 U885 ( .A(G101), .B(n1206), .ZN(G3) );
NAND2_X1 U886 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
INV_X1 U887 ( .A(n1192), .ZN(n1208) );
NAND4_X1 U888 ( .A1(n1029), .A2(n1037), .A3(n1047), .A4(n1194), .ZN(n1192) );
XNOR2_X1 U889 ( .A(n1042), .B(KEYINPUT36), .ZN(n1207) );
XNOR2_X1 U890 ( .A(G125), .B(n1168), .ZN(G27) );
NAND4_X1 U891 ( .A1(n1193), .A2(n1028), .A3(n1053), .A4(n1181), .ZN(n1168) );
NAND2_X1 U892 ( .A1(n1209), .A2(n1210), .ZN(n1181) );
NAND2_X1 U893 ( .A1(n1211), .A2(n1071), .ZN(n1210) );
INV_X1 U894 ( .A(G900), .ZN(n1071) );
AND2_X1 U895 ( .A1(n1052), .A2(n1042), .ZN(n1193) );
XNOR2_X1 U896 ( .A(G122), .B(n1212), .ZN(G24) );
NOR2_X1 U897 ( .A1(n1213), .A2(KEYINPUT25), .ZN(n1212) );
INV_X1 U898 ( .A(n1183), .ZN(n1213) );
NAND3_X1 U899 ( .A1(n1214), .A2(n1033), .A3(n1196), .ZN(n1183) );
AND2_X1 U900 ( .A1(n1215), .A2(n1216), .ZN(n1196) );
XNOR2_X1 U901 ( .A(n1217), .B(KEYINPUT15), .ZN(n1215) );
NOR2_X1 U902 ( .A1(n1056), .A2(n1173), .ZN(n1033) );
XNOR2_X1 U903 ( .A(G119), .B(n1184), .ZN(G21) );
NAND4_X1 U904 ( .A1(n1214), .A2(n1037), .A3(n1173), .A4(n1056), .ZN(n1184) );
XNOR2_X1 U905 ( .A(G116), .B(n1189), .ZN(G18) );
NAND3_X1 U906 ( .A1(n1029), .A2(n1051), .A3(n1214), .ZN(n1189) );
AND2_X1 U907 ( .A1(n1218), .A2(n1216), .ZN(n1051) );
XNOR2_X1 U908 ( .A(G113), .B(n1188), .ZN(G15) );
NAND3_X1 U909 ( .A1(n1214), .A2(n1029), .A3(n1052), .ZN(n1188) );
NOR2_X1 U910 ( .A1(n1216), .A2(n1218), .ZN(n1052) );
INV_X1 U911 ( .A(n1217), .ZN(n1218) );
NOR2_X1 U912 ( .A1(n1173), .A2(n1030), .ZN(n1029) );
AND3_X1 U913 ( .A1(n1042), .A2(n1194), .A3(n1053), .ZN(n1214) );
INV_X1 U914 ( .A(n1024), .ZN(n1053) );
NAND2_X1 U915 ( .A1(n1219), .A2(n1049), .ZN(n1024) );
INV_X1 U916 ( .A(n1048), .ZN(n1219) );
XNOR2_X1 U917 ( .A(n1220), .B(n1221), .ZN(G12) );
NOR2_X1 U918 ( .A1(n1187), .A2(n1222), .ZN(n1221) );
XOR2_X1 U919 ( .A(KEYINPUT54), .B(KEYINPUT49), .Z(n1222) );
NAND3_X1 U920 ( .A1(n1037), .A2(n1190), .A3(n1028), .ZN(n1187) );
AND2_X1 U921 ( .A1(n1030), .A2(n1173), .ZN(n1028) );
XOR2_X1 U922 ( .A(n1058), .B(KEYINPUT57), .Z(n1173) );
XNOR2_X1 U923 ( .A(n1223), .B(n1118), .ZN(n1058) );
AND2_X1 U924 ( .A1(G217), .A2(n1224), .ZN(n1118) );
NAND2_X1 U925 ( .A1(n1116), .A2(n1225), .ZN(n1223) );
XOR2_X1 U926 ( .A(n1226), .B(n1227), .Z(n1116) );
NOR2_X1 U927 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
INV_X1 U928 ( .A(G221), .ZN(n1229) );
XNOR2_X1 U929 ( .A(G137), .B(n1230), .ZN(n1226) );
NOR2_X1 U930 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XOR2_X1 U931 ( .A(KEYINPUT26), .B(n1233), .Z(n1232) );
NOR2_X1 U932 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
AND2_X1 U933 ( .A1(n1235), .A2(n1234), .ZN(n1231) );
XOR2_X1 U934 ( .A(n1236), .B(n1237), .Z(n1234) );
XOR2_X1 U935 ( .A(KEYINPUT45), .B(G146), .Z(n1237) );
XNOR2_X1 U936 ( .A(G125), .B(G140), .ZN(n1236) );
NAND3_X1 U937 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1235) );
NAND2_X1 U938 ( .A1(KEYINPUT48), .A2(n1241), .ZN(n1240) );
OR3_X1 U939 ( .A1(n1242), .A2(KEYINPUT48), .A3(G110), .ZN(n1239) );
NAND2_X1 U940 ( .A1(G110), .A2(n1242), .ZN(n1238) );
NAND2_X1 U941 ( .A1(KEYINPUT22), .A2(n1243), .ZN(n1242) );
INV_X1 U942 ( .A(n1241), .ZN(n1243) );
XOR2_X1 U943 ( .A(G119), .B(n1244), .Z(n1241) );
INV_X1 U944 ( .A(n1056), .ZN(n1030) );
XNOR2_X1 U945 ( .A(n1245), .B(G472), .ZN(n1056) );
NAND2_X1 U946 ( .A1(n1133), .A2(n1225), .ZN(n1245) );
XOR2_X1 U947 ( .A(n1246), .B(n1247), .Z(n1133) );
XOR2_X1 U948 ( .A(n1111), .B(n1248), .Z(n1247) );
XNOR2_X1 U949 ( .A(G101), .B(n1249), .ZN(n1248) );
NAND2_X1 U950 ( .A1(G210), .A2(n1250), .ZN(n1249) );
XOR2_X1 U951 ( .A(n1142), .B(n1155), .Z(n1246) );
AND3_X1 U952 ( .A1(n1047), .A2(n1194), .A3(n1042), .ZN(n1190) );
INV_X1 U953 ( .A(n1175), .ZN(n1042) );
NAND2_X1 U954 ( .A1(n1044), .A2(n1043), .ZN(n1175) );
NAND2_X1 U955 ( .A1(G214), .A2(n1251), .ZN(n1043) );
XNOR2_X1 U956 ( .A(n1252), .B(n1060), .ZN(n1044) );
NAND2_X1 U957 ( .A1(G210), .A2(n1251), .ZN(n1060) );
NAND2_X1 U958 ( .A1(n1253), .A2(n1225), .ZN(n1251) );
XNOR2_X1 U959 ( .A(KEYINPUT17), .B(n1254), .ZN(n1252) );
NOR2_X1 U960 ( .A1(n1059), .A2(KEYINPUT0), .ZN(n1254) );
AND3_X1 U961 ( .A1(n1255), .A2(n1225), .A3(n1256), .ZN(n1059) );
XOR2_X1 U962 ( .A(KEYINPUT8), .B(n1257), .Z(n1256) );
NOR2_X1 U963 ( .A1(n1156), .A2(n1258), .ZN(n1257) );
NAND2_X1 U964 ( .A1(n1156), .A2(n1258), .ZN(n1255) );
XOR2_X1 U965 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U966 ( .A(KEYINPUT39), .B(n1261), .Z(n1260) );
NOR2_X1 U967 ( .A1(n1151), .A2(KEYINPUT31), .ZN(n1261) );
NOR2_X1 U968 ( .A1(n1097), .A2(G953), .ZN(n1151) );
INV_X1 U969 ( .A(G224), .ZN(n1097) );
XNOR2_X1 U970 ( .A(n1155), .B(n1159), .ZN(n1259) );
XNOR2_X1 U971 ( .A(n1083), .B(KEYINPUT35), .ZN(n1159) );
INV_X1 U972 ( .A(G125), .ZN(n1083) );
XOR2_X1 U973 ( .A(G146), .B(n1262), .Z(n1155) );
XOR2_X1 U974 ( .A(n1263), .B(n1264), .Z(n1156) );
NOR2_X1 U975 ( .A1(KEYINPUT30), .A2(n1109), .ZN(n1264) );
XNOR2_X1 U976 ( .A(G122), .B(n1220), .ZN(n1109) );
NAND2_X1 U977 ( .A1(n1265), .A2(n1266), .ZN(n1263) );
NAND2_X1 U978 ( .A1(n1267), .A2(n1110), .ZN(n1266) );
XOR2_X1 U979 ( .A(KEYINPUT62), .B(n1268), .Z(n1265) );
NOR2_X1 U980 ( .A1(n1110), .A2(n1267), .ZN(n1268) );
XOR2_X1 U981 ( .A(KEYINPUT28), .B(n1111), .Z(n1267) );
XNOR2_X1 U982 ( .A(n1269), .B(n1270), .ZN(n1111) );
XNOR2_X1 U983 ( .A(G113), .B(G119), .ZN(n1269) );
NAND2_X1 U984 ( .A1(n1209), .A2(n1271), .ZN(n1194) );
NAND2_X1 U985 ( .A1(n1211), .A2(n1098), .ZN(n1271) );
INV_X1 U986 ( .A(G898), .ZN(n1098) );
NOR3_X1 U987 ( .A1(n1225), .A2(n1020), .A3(n1072), .ZN(n1211) );
INV_X1 U988 ( .A(n1272), .ZN(n1020) );
NAND3_X1 U989 ( .A1(n1061), .A2(n1272), .A3(G952), .ZN(n1209) );
NAND2_X1 U990 ( .A1(G234), .A2(n1273), .ZN(n1272) );
XNOR2_X1 U991 ( .A(KEYINPUT19), .B(n1253), .ZN(n1273) );
INV_X1 U992 ( .A(G237), .ZN(n1253) );
XOR2_X1 U993 ( .A(G953), .B(KEYINPUT41), .Z(n1061) );
INV_X1 U994 ( .A(n1180), .ZN(n1047) );
NAND2_X1 U995 ( .A1(n1048), .A2(n1049), .ZN(n1180) );
NAND2_X1 U996 ( .A1(G221), .A2(n1224), .ZN(n1049) );
NAND2_X1 U997 ( .A1(G234), .A2(n1225), .ZN(n1224) );
XNOR2_X1 U998 ( .A(n1274), .B(G469), .ZN(n1048) );
NAND2_X1 U999 ( .A1(n1275), .A2(n1225), .ZN(n1274) );
INV_X1 U1000 ( .A(G902), .ZN(n1225) );
XOR2_X1 U1001 ( .A(n1276), .B(n1277), .Z(n1275) );
NOR2_X1 U1002 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
XNOR2_X1 U1003 ( .A(KEYINPUT50), .B(KEYINPUT34), .ZN(n1279) );
NOR3_X1 U1004 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1278) );
NOR2_X1 U1005 ( .A1(KEYINPUT21), .A2(n1283), .ZN(n1282) );
NOR2_X1 U1006 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NOR3_X1 U1007 ( .A1(n1220), .A2(KEYINPUT18), .A3(G140), .ZN(n1285) );
AND2_X1 U1008 ( .A1(n1220), .A2(KEYINPUT18), .ZN(n1284) );
NOR2_X1 U1009 ( .A1(n1286), .A2(n1287), .ZN(n1281) );
INV_X1 U1010 ( .A(KEYINPUT21), .ZN(n1287) );
NOR2_X1 U1011 ( .A1(G140), .A2(n1288), .ZN(n1286) );
XNOR2_X1 U1012 ( .A(KEYINPUT18), .B(G110), .ZN(n1288) );
NOR2_X1 U1013 ( .A1(G110), .A2(n1093), .ZN(n1280) );
XNOR2_X1 U1014 ( .A(n1289), .B(n1145), .ZN(n1276) );
NAND2_X1 U1015 ( .A1(G227), .A2(n1072), .ZN(n1145) );
NAND3_X1 U1016 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1289) );
NAND2_X1 U1017 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
INV_X1 U1018 ( .A(KEYINPUT46), .ZN(n1294) );
NAND3_X1 U1019 ( .A1(KEYINPUT46), .A2(n1295), .A3(n1142), .ZN(n1291) );
OR2_X1 U1020 ( .A1(n1142), .A2(n1295), .ZN(n1290) );
NOR2_X1 U1021 ( .A1(KEYINPUT24), .A2(n1293), .ZN(n1295) );
XNOR2_X1 U1022 ( .A(n1086), .B(n1110), .ZN(n1293) );
XOR2_X1 U1023 ( .A(G101), .B(n1296), .Z(n1110) );
XNOR2_X1 U1024 ( .A(n1297), .B(G104), .ZN(n1296) );
AND2_X1 U1025 ( .A1(n1298), .A2(n1299), .ZN(n1086) );
NAND2_X1 U1026 ( .A1(n1300), .A2(n1244), .ZN(n1299) );
INV_X1 U1027 ( .A(G128), .ZN(n1244) );
XNOR2_X1 U1028 ( .A(n1301), .B(n1302), .ZN(n1300) );
NAND2_X1 U1029 ( .A1(G128), .A2(n1303), .ZN(n1298) );
XNOR2_X1 U1030 ( .A(G143), .B(n1302), .ZN(n1303) );
NOR2_X1 U1031 ( .A1(G146), .A2(KEYINPUT63), .ZN(n1302) );
XNOR2_X1 U1032 ( .A(G137), .B(n1092), .ZN(n1142) );
XOR2_X1 U1033 ( .A(G131), .B(G134), .Z(n1092) );
NOR2_X1 U1034 ( .A1(n1217), .A2(n1216), .ZN(n1037) );
XOR2_X1 U1035 ( .A(n1304), .B(n1305), .Z(n1216) );
XOR2_X1 U1036 ( .A(KEYINPUT55), .B(G478), .Z(n1305) );
NAND2_X1 U1037 ( .A1(n1306), .A2(n1126), .ZN(n1304) );
XOR2_X1 U1038 ( .A(n1307), .B(n1308), .Z(n1126) );
XNOR2_X1 U1039 ( .A(n1262), .B(n1309), .ZN(n1308) );
XNOR2_X1 U1040 ( .A(n1270), .B(n1310), .ZN(n1309) );
NOR3_X1 U1041 ( .A1(n1311), .A2(KEYINPUT60), .A3(n1228), .ZN(n1310) );
NAND2_X1 U1042 ( .A1(G234), .A2(n1072), .ZN(n1228) );
INV_X1 U1043 ( .A(G953), .ZN(n1072) );
INV_X1 U1044 ( .A(G217), .ZN(n1311) );
XOR2_X1 U1045 ( .A(G116), .B(KEYINPUT14), .Z(n1270) );
XOR2_X1 U1046 ( .A(G128), .B(G143), .Z(n1262) );
XOR2_X1 U1047 ( .A(n1312), .B(n1313), .Z(n1307) );
XOR2_X1 U1048 ( .A(G122), .B(n1314), .Z(n1313) );
NOR2_X1 U1049 ( .A1(KEYINPUT1), .A2(n1297), .ZN(n1314) );
INV_X1 U1050 ( .A(G107), .ZN(n1297) );
XNOR2_X1 U1051 ( .A(G134), .B(KEYINPUT9), .ZN(n1312) );
XNOR2_X1 U1052 ( .A(G902), .B(KEYINPUT59), .ZN(n1306) );
XNOR2_X1 U1053 ( .A(n1315), .B(G475), .ZN(n1217) );
OR2_X1 U1054 ( .A1(n1129), .A2(G902), .ZN(n1315) );
XNOR2_X1 U1055 ( .A(n1316), .B(n1317), .ZN(n1129) );
XOR2_X1 U1056 ( .A(G122), .B(G113), .Z(n1317) );
XOR2_X1 U1057 ( .A(n1318), .B(G104), .Z(n1316) );
NAND2_X1 U1058 ( .A1(n1319), .A2(KEYINPUT51), .ZN(n1318) );
XOR2_X1 U1059 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1060 ( .A(G131), .B(n1322), .Z(n1321) );
XNOR2_X1 U1061 ( .A(G146), .B(n1301), .ZN(n1322) );
INV_X1 U1062 ( .A(G143), .ZN(n1301) );
XOR2_X1 U1063 ( .A(n1323), .B(n1324), .Z(n1320) );
NOR2_X1 U1064 ( .A1(KEYINPUT13), .A2(n1325), .ZN(n1324) );
XNOR2_X1 U1065 ( .A(G125), .B(n1326), .ZN(n1325) );
NAND2_X1 U1066 ( .A1(KEYINPUT6), .A2(n1093), .ZN(n1326) );
INV_X1 U1067 ( .A(G140), .ZN(n1093) );
NAND2_X1 U1068 ( .A1(G214), .A2(n1250), .ZN(n1323) );
NOR2_X1 U1069 ( .A1(G953), .A2(G237), .ZN(n1250) );
INV_X1 U1070 ( .A(G110), .ZN(n1220) );
endmodule


