//Key = 0110000101111011110111011000110111011110110100000101011000100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309;

XOR2_X1 U723 ( .A(n1004), .B(n1005), .Z(G9) );
XNOR2_X1 U724 ( .A(G107), .B(KEYINPUT44), .ZN(n1005) );
NAND3_X1 U725 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(G75) );
NAND2_X1 U726 ( .A1(G952), .A2(n1009), .ZN(n1008) );
NAND4_X1 U727 ( .A1(n1010), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1009) );
NAND4_X1 U728 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1013) );
NOR3_X1 U729 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1017) );
AND3_X1 U730 ( .A1(KEYINPUT55), .A2(n1021), .A3(n1022), .ZN(n1020) );
NOR2_X1 U731 ( .A1(KEYINPUT55), .A2(n1023), .ZN(n1019) );
XNOR2_X1 U732 ( .A(n1024), .B(n1025), .ZN(n1023) );
NAND4_X1 U733 ( .A1(n1021), .A2(n1026), .A3(n1027), .A4(n1015), .ZN(n1012) );
NAND2_X1 U734 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND3_X1 U735 ( .A1(n1014), .A2(n1030), .A3(n1031), .ZN(n1029) );
NAND2_X1 U736 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NAND2_X1 U737 ( .A1(n1016), .A2(n1034), .ZN(n1028) );
NAND2_X1 U738 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U739 ( .A1(n1031), .A2(n1037), .ZN(n1036) );
NAND2_X1 U740 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U741 ( .A1(n1014), .A2(n1040), .ZN(n1035) );
NAND2_X1 U742 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U743 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND3_X1 U744 ( .A1(n1045), .A2(n1021), .A3(n1046), .ZN(n1006) );
NOR3_X1 U745 ( .A1(n1047), .A2(n1043), .A3(n1022), .ZN(n1046) );
INV_X1 U746 ( .A(n1024), .ZN(n1022) );
XOR2_X1 U747 ( .A(n1048), .B(KEYINPUT43), .Z(n1045) );
NAND4_X1 U748 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
XNOR2_X1 U749 ( .A(G472), .B(n1053), .ZN(n1052) );
NAND2_X1 U750 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT16), .Z(n1054) );
XOR2_X1 U752 ( .A(n1056), .B(n1057), .Z(n1051) );
XNOR2_X1 U753 ( .A(G478), .B(KEYINPUT0), .ZN(n1056) );
XOR2_X1 U754 ( .A(n1058), .B(n1059), .Z(n1050) );
XOR2_X1 U755 ( .A(KEYINPUT9), .B(KEYINPUT49), .Z(n1059) );
XOR2_X1 U756 ( .A(n1060), .B(n1061), .Z(n1049) );
XOR2_X1 U757 ( .A(n1062), .B(n1063), .Z(G72) );
XOR2_X1 U758 ( .A(n1064), .B(n1065), .Z(n1063) );
NAND2_X1 U759 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
INV_X1 U760 ( .A(n1068), .ZN(n1067) );
XOR2_X1 U761 ( .A(n1069), .B(n1070), .Z(n1066) );
XOR2_X1 U762 ( .A(n1071), .B(n1072), .Z(n1070) );
XOR2_X1 U763 ( .A(n1073), .B(n1074), .Z(n1069) );
XNOR2_X1 U764 ( .A(G134), .B(KEYINPUT35), .ZN(n1073) );
NAND2_X1 U765 ( .A1(G953), .A2(n1075), .ZN(n1064) );
NAND2_X1 U766 ( .A1(G900), .A2(G227), .ZN(n1075) );
NAND2_X1 U767 ( .A1(n1076), .A2(n1077), .ZN(n1062) );
NAND2_X1 U768 ( .A1(KEYINPUT28), .A2(n1078), .ZN(n1077) );
OR2_X1 U769 ( .A1(KEYINPUT61), .A2(n1078), .ZN(n1076) );
NOR2_X1 U770 ( .A1(G953), .A2(n1011), .ZN(n1078) );
NAND2_X1 U771 ( .A1(n1079), .A2(n1080), .ZN(G69) );
NAND2_X1 U772 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U773 ( .A1(G953), .A2(n1083), .ZN(n1082) );
NAND3_X1 U774 ( .A1(G953), .A2(n1084), .A3(n1085), .ZN(n1079) );
XNOR2_X1 U775 ( .A(n1081), .B(KEYINPUT34), .ZN(n1085) );
XNOR2_X1 U776 ( .A(n1086), .B(n1087), .ZN(n1081) );
NOR2_X1 U777 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U778 ( .A(KEYINPUT53), .B(n1090), .Z(n1089) );
NOR2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR2_X1 U780 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1091) );
XNOR2_X1 U782 ( .A(KEYINPUT39), .B(n1093), .ZN(n1096) );
NAND2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1093) );
NAND3_X1 U784 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
INV_X1 U785 ( .A(KEYINPUT38), .ZN(n1101) );
NAND2_X1 U786 ( .A1(n1102), .A2(KEYINPUT38), .ZN(n1097) );
NOR2_X1 U787 ( .A1(G898), .A2(n1007), .ZN(n1088) );
NAND2_X1 U788 ( .A1(n1007), .A2(n1103), .ZN(n1086) );
NAND2_X1 U789 ( .A1(G898), .A2(G224), .ZN(n1084) );
NOR2_X1 U790 ( .A1(n1104), .A2(n1105), .ZN(G66) );
XOR2_X1 U791 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR3_X1 U792 ( .A1(n1108), .A2(KEYINPUT42), .A3(n1061), .ZN(n1106) );
NOR2_X1 U793 ( .A1(n1104), .A2(n1109), .ZN(G63) );
NOR3_X1 U794 ( .A1(n1057), .A2(n1110), .A3(n1111), .ZN(n1109) );
AND3_X1 U795 ( .A1(n1112), .A2(G478), .A3(n1113), .ZN(n1111) );
NOR2_X1 U796 ( .A1(n1114), .A2(n1112), .ZN(n1110) );
NOR2_X1 U797 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
INV_X1 U798 ( .A(G478), .ZN(n1116) );
NOR2_X1 U799 ( .A1(n1117), .A2(n1103), .ZN(n1115) );
NOR2_X1 U800 ( .A1(n1104), .A2(n1118), .ZN(G60) );
XOR2_X1 U801 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U802 ( .A1(n1113), .A2(G475), .ZN(n1119) );
XOR2_X1 U803 ( .A(n1121), .B(n1122), .Z(G6) );
XOR2_X1 U804 ( .A(KEYINPUT51), .B(G104), .Z(n1122) );
NAND3_X1 U805 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1121) );
XNOR2_X1 U806 ( .A(KEYINPUT3), .B(n1126), .ZN(n1124) );
NOR2_X1 U807 ( .A1(n1104), .A2(n1127), .ZN(G57) );
XOR2_X1 U808 ( .A(n1128), .B(n1129), .Z(n1127) );
XNOR2_X1 U809 ( .A(n1130), .B(n1131), .ZN(n1129) );
XOR2_X1 U810 ( .A(n1132), .B(n1133), .Z(n1128) );
NOR2_X1 U811 ( .A1(KEYINPUT5), .A2(n1134), .ZN(n1133) );
XOR2_X1 U812 ( .A(n1135), .B(KEYINPUT13), .Z(n1132) );
NAND2_X1 U813 ( .A1(n1113), .A2(G472), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1104), .A2(n1136), .ZN(G54) );
XOR2_X1 U815 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U816 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U817 ( .A1(KEYINPUT1), .A2(n1141), .ZN(n1139) );
XOR2_X1 U818 ( .A(n1142), .B(n1143), .Z(n1137) );
XNOR2_X1 U819 ( .A(n1144), .B(n1145), .ZN(n1143) );
NOR2_X1 U820 ( .A1(KEYINPUT48), .A2(n1146), .ZN(n1145) );
XNOR2_X1 U821 ( .A(n1147), .B(n1148), .ZN(n1146) );
NAND2_X1 U822 ( .A1(KEYINPUT19), .A2(n1149), .ZN(n1147) );
NAND2_X1 U823 ( .A1(n1113), .A2(G469), .ZN(n1142) );
NOR2_X1 U824 ( .A1(n1104), .A2(n1150), .ZN(G51) );
XOR2_X1 U825 ( .A(n1151), .B(n1152), .Z(n1150) );
XNOR2_X1 U826 ( .A(n1153), .B(n1154), .ZN(n1152) );
NAND2_X1 U827 ( .A1(n1113), .A2(n1155), .ZN(n1153) );
INV_X1 U828 ( .A(n1108), .ZN(n1113) );
NAND2_X1 U829 ( .A1(G902), .A2(n1156), .ZN(n1108) );
NAND2_X1 U830 ( .A1(n1010), .A2(n1011), .ZN(n1156) );
INV_X1 U831 ( .A(n1117), .ZN(n1011) );
NAND2_X1 U832 ( .A1(n1157), .A2(n1158), .ZN(n1117) );
NOR4_X1 U833 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1158) );
NOR4_X1 U834 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1157) );
NOR3_X1 U835 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1166) );
INV_X1 U836 ( .A(n1103), .ZN(n1010) );
NAND4_X1 U837 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1103) );
AND4_X1 U838 ( .A1(n1004), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1173) );
NAND3_X1 U839 ( .A1(n1177), .A2(n1123), .A3(n1178), .ZN(n1004) );
OR2_X1 U840 ( .A1(n1179), .A2(KEYINPUT18), .ZN(n1172) );
NAND2_X1 U841 ( .A1(n1180), .A2(n1181), .ZN(n1170) );
NAND2_X1 U842 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND4_X1 U843 ( .A1(KEYINPUT18), .A2(n1184), .A3(n1177), .A4(n1018), .ZN(n1183) );
NAND2_X1 U844 ( .A1(n1178), .A2(n1185), .ZN(n1182) );
NAND2_X1 U845 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NAND2_X1 U846 ( .A1(n1125), .A2(n1016), .ZN(n1187) );
NAND2_X1 U847 ( .A1(n1188), .A2(n1184), .ZN(n1186) );
XOR2_X1 U848 ( .A(KEYINPUT31), .B(n1168), .Z(n1188) );
INV_X1 U849 ( .A(n1014), .ZN(n1168) );
NOR2_X1 U850 ( .A1(n1007), .A2(G952), .ZN(n1104) );
XNOR2_X1 U851 ( .A(G146), .B(n1189), .ZN(G48) );
NAND2_X1 U852 ( .A1(KEYINPUT12), .A2(n1165), .ZN(n1189) );
NOR4_X1 U853 ( .A1(n1190), .A2(n1169), .A3(n1039), .A4(n1041), .ZN(n1165) );
INV_X1 U854 ( .A(n1191), .ZN(n1041) );
XNOR2_X1 U855 ( .A(n1164), .B(n1192), .ZN(G45) );
XNOR2_X1 U856 ( .A(G143), .B(KEYINPUT47), .ZN(n1192) );
AND4_X1 U857 ( .A1(n1191), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1164) );
NOR2_X1 U858 ( .A1(n1032), .A2(n1190), .ZN(n1195) );
XNOR2_X1 U859 ( .A(G140), .B(n1196), .ZN(G42) );
NAND2_X1 U860 ( .A1(KEYINPUT10), .A2(n1163), .ZN(n1196) );
NOR3_X1 U861 ( .A1(n1039), .A2(n1033), .A3(n1167), .ZN(n1163) );
XOR2_X1 U862 ( .A(G137), .B(n1197), .Z(G39) );
NOR3_X1 U863 ( .A1(n1198), .A2(n1169), .A3(n1167), .ZN(n1197) );
XOR2_X1 U864 ( .A(n1014), .B(KEYINPUT7), .Z(n1198) );
XNOR2_X1 U865 ( .A(n1199), .B(n1200), .ZN(G36) );
NOR2_X1 U866 ( .A1(KEYINPUT50), .A2(n1201), .ZN(n1200) );
INV_X1 U867 ( .A(n1162), .ZN(n1201) );
NOR3_X1 U868 ( .A1(n1032), .A2(n1038), .A3(n1167), .ZN(n1162) );
XOR2_X1 U869 ( .A(G131), .B(n1161), .Z(G33) );
NOR3_X1 U870 ( .A1(n1039), .A2(n1032), .A3(n1167), .ZN(n1161) );
NAND4_X1 U871 ( .A1(n1021), .A2(n1026), .A3(n1191), .A4(n1202), .ZN(n1167) );
XOR2_X1 U872 ( .A(n1178), .B(KEYINPUT26), .Z(n1191) );
XNOR2_X1 U873 ( .A(n1024), .B(KEYINPUT20), .ZN(n1026) );
INV_X1 U874 ( .A(n1025), .ZN(n1021) );
XOR2_X1 U875 ( .A(G128), .B(n1160), .Z(G30) );
NOR4_X1 U876 ( .A1(n1190), .A2(n1169), .A3(n1126), .A4(n1038), .ZN(n1160) );
INV_X1 U877 ( .A(n1177), .ZN(n1038) );
INV_X1 U878 ( .A(n1178), .ZN(n1126) );
XNOR2_X1 U879 ( .A(G101), .B(n1203), .ZN(G3) );
NAND2_X1 U880 ( .A1(n1184), .A2(n1204), .ZN(n1203) );
XNOR2_X1 U881 ( .A(G125), .B(n1205), .ZN(G27) );
NAND2_X1 U882 ( .A1(KEYINPUT11), .A2(n1159), .ZN(n1205) );
NOR4_X1 U883 ( .A1(n1190), .A2(n1039), .A3(n1018), .A4(n1033), .ZN(n1159) );
INV_X1 U884 ( .A(n1206), .ZN(n1033) );
NAND3_X1 U885 ( .A1(n1202), .A2(n1024), .A3(n1025), .ZN(n1190) );
NAND2_X1 U886 ( .A1(n1207), .A2(n1208), .ZN(n1202) );
NAND3_X1 U887 ( .A1(n1209), .A2(n1007), .A3(G952), .ZN(n1208) );
NAND3_X1 U888 ( .A1(G902), .A2(n1015), .A3(n1068), .ZN(n1207) );
NOR2_X1 U889 ( .A1(n1007), .A2(G900), .ZN(n1068) );
XNOR2_X1 U890 ( .A(G122), .B(n1171), .ZN(G24) );
NAND4_X1 U891 ( .A1(n1031), .A2(n1123), .A3(n1194), .A4(n1193), .ZN(n1171) );
AND2_X1 U892 ( .A1(n1180), .A2(n1016), .ZN(n1123) );
NOR2_X1 U893 ( .A1(n1210), .A2(n1211), .ZN(n1016) );
XNOR2_X1 U894 ( .A(G119), .B(n1176), .ZN(G21) );
NAND3_X1 U895 ( .A1(n1212), .A2(n1014), .A3(n1213), .ZN(n1176) );
INV_X1 U896 ( .A(n1169), .ZN(n1213) );
NAND2_X1 U897 ( .A1(n1211), .A2(n1210), .ZN(n1169) );
XNOR2_X1 U898 ( .A(G116), .B(n1179), .ZN(G18) );
NAND3_X1 U899 ( .A1(n1212), .A2(n1177), .A3(n1184), .ZN(n1179) );
XNOR2_X1 U900 ( .A(G113), .B(n1175), .ZN(G15) );
NAND3_X1 U901 ( .A1(n1184), .A2(n1212), .A3(n1125), .ZN(n1175) );
INV_X1 U902 ( .A(n1039), .ZN(n1125) );
NAND2_X1 U903 ( .A1(n1193), .A2(n1214), .ZN(n1039) );
AND2_X1 U904 ( .A1(n1031), .A2(n1180), .ZN(n1212) );
INV_X1 U905 ( .A(n1018), .ZN(n1031) );
NAND2_X1 U906 ( .A1(n1044), .A2(n1215), .ZN(n1018) );
INV_X1 U907 ( .A(n1032), .ZN(n1184) );
NAND2_X1 U908 ( .A1(n1216), .A2(n1211), .ZN(n1032) );
XOR2_X1 U909 ( .A(KEYINPUT32), .B(n1210), .Z(n1216) );
XNOR2_X1 U910 ( .A(G110), .B(n1174), .ZN(G12) );
NAND2_X1 U911 ( .A1(n1206), .A2(n1204), .ZN(n1174) );
AND3_X1 U912 ( .A1(n1180), .A2(n1014), .A3(n1178), .ZN(n1204) );
NOR2_X1 U913 ( .A1(n1044), .A2(n1043), .ZN(n1178) );
INV_X1 U914 ( .A(n1215), .ZN(n1043) );
NAND2_X1 U915 ( .A1(G221), .A2(n1217), .ZN(n1215) );
XOR2_X1 U916 ( .A(n1047), .B(KEYINPUT24), .Z(n1044) );
XOR2_X1 U917 ( .A(n1218), .B(n1219), .Z(n1047) );
XOR2_X1 U918 ( .A(KEYINPUT21), .B(G469), .Z(n1219) );
NAND2_X1 U919 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
XOR2_X1 U920 ( .A(n1222), .B(n1223), .Z(n1220) );
XNOR2_X1 U921 ( .A(n1149), .B(n1148), .ZN(n1223) );
XNOR2_X1 U922 ( .A(n1224), .B(n1225), .ZN(n1149) );
XOR2_X1 U923 ( .A(G104), .B(G101), .Z(n1225) );
XOR2_X1 U924 ( .A(n1226), .B(n1074), .Z(n1224) );
NAND2_X1 U925 ( .A1(KEYINPUT54), .A2(n1227), .ZN(n1226) );
XOR2_X1 U926 ( .A(n1228), .B(n1229), .Z(n1222) );
XNOR2_X1 U927 ( .A(n1144), .B(n1141), .ZN(n1229) );
AND2_X1 U928 ( .A1(G227), .A2(n1007), .ZN(n1141) );
INV_X1 U929 ( .A(G110), .ZN(n1144) );
NAND2_X1 U930 ( .A1(KEYINPUT14), .A2(n1140), .ZN(n1228) );
XNOR2_X1 U931 ( .A(G140), .B(KEYINPUT63), .ZN(n1140) );
NAND2_X1 U932 ( .A1(n1230), .A2(n1231), .ZN(n1014) );
OR3_X1 U933 ( .A1(n1194), .A2(n1193), .A3(KEYINPUT30), .ZN(n1231) );
INV_X1 U934 ( .A(n1214), .ZN(n1194) );
NAND2_X1 U935 ( .A1(KEYINPUT30), .A2(n1177), .ZN(n1230) );
NOR2_X1 U936 ( .A1(n1214), .A2(n1193), .ZN(n1177) );
XNOR2_X1 U937 ( .A(n1058), .B(KEYINPUT22), .ZN(n1193) );
XOR2_X1 U938 ( .A(n1232), .B(G475), .Z(n1058) );
NAND2_X1 U939 ( .A1(n1120), .A2(n1221), .ZN(n1232) );
XNOR2_X1 U940 ( .A(n1233), .B(n1234), .ZN(n1120) );
XOR2_X1 U941 ( .A(n1235), .B(n1236), .Z(n1234) );
XNOR2_X1 U942 ( .A(n1237), .B(n1238), .ZN(n1236) );
NOR2_X1 U943 ( .A1(KEYINPUT56), .A2(n1239), .ZN(n1238) );
XNOR2_X1 U944 ( .A(n1240), .B(n1241), .ZN(n1239) );
NAND2_X1 U945 ( .A1(G214), .A2(n1242), .ZN(n1240) );
XNOR2_X1 U946 ( .A(G104), .B(G113), .ZN(n1235) );
XOR2_X1 U947 ( .A(n1243), .B(n1244), .Z(n1233) );
XOR2_X1 U948 ( .A(KEYINPUT6), .B(G146), .Z(n1244) );
XNOR2_X1 U949 ( .A(G131), .B(G122), .ZN(n1243) );
XNOR2_X1 U950 ( .A(n1245), .B(n1057), .ZN(n1214) );
NOR2_X1 U951 ( .A1(n1112), .A2(G902), .ZN(n1057) );
XOR2_X1 U952 ( .A(n1246), .B(n1247), .Z(n1112) );
NOR2_X1 U953 ( .A1(KEYINPUT59), .A2(n1248), .ZN(n1247) );
XOR2_X1 U954 ( .A(n1249), .B(n1250), .Z(n1248) );
XNOR2_X1 U955 ( .A(n1251), .B(n1252), .ZN(n1250) );
XNOR2_X1 U956 ( .A(n1253), .B(n1254), .ZN(n1251) );
NAND2_X1 U957 ( .A1(KEYINPUT40), .A2(n1227), .ZN(n1253) );
INV_X1 U958 ( .A(G107), .ZN(n1227) );
XNOR2_X1 U959 ( .A(G122), .B(n1255), .ZN(n1249) );
XNOR2_X1 U960 ( .A(n1199), .B(G128), .ZN(n1255) );
INV_X1 U961 ( .A(G134), .ZN(n1199) );
NAND2_X1 U962 ( .A1(G217), .A2(n1256), .ZN(n1246) );
NAND2_X1 U963 ( .A1(n1257), .A2(KEYINPUT33), .ZN(n1245) );
XNOR2_X1 U964 ( .A(G478), .B(KEYINPUT52), .ZN(n1257) );
AND4_X1 U965 ( .A1(n1025), .A2(n1024), .A3(n1258), .A4(n1259), .ZN(n1180) );
NAND2_X1 U966 ( .A1(n1260), .A2(n1007), .ZN(n1259) );
NAND2_X1 U967 ( .A1(G952), .A2(n1209), .ZN(n1260) );
XOR2_X1 U968 ( .A(n1015), .B(KEYINPUT46), .Z(n1209) );
NAND2_X1 U969 ( .A1(G953), .A2(n1261), .ZN(n1258) );
NAND3_X1 U970 ( .A1(n1015), .A2(n1262), .A3(G902), .ZN(n1261) );
INV_X1 U971 ( .A(G898), .ZN(n1262) );
NAND2_X1 U972 ( .A1(G237), .A2(G234), .ZN(n1015) );
NAND2_X1 U973 ( .A1(G214), .A2(n1263), .ZN(n1024) );
XNOR2_X1 U974 ( .A(n1264), .B(n1155), .ZN(n1025) );
AND2_X1 U975 ( .A1(G210), .A2(n1263), .ZN(n1155) );
NAND2_X1 U976 ( .A1(n1265), .A2(n1221), .ZN(n1263) );
INV_X1 U977 ( .A(G237), .ZN(n1265) );
NAND2_X1 U978 ( .A1(n1266), .A2(n1221), .ZN(n1264) );
XOR2_X1 U979 ( .A(n1267), .B(n1154), .Z(n1266) );
XNOR2_X1 U980 ( .A(n1102), .B(n1094), .ZN(n1154) );
INV_X1 U981 ( .A(n1095), .ZN(n1094) );
XNOR2_X1 U982 ( .A(n1268), .B(n1269), .ZN(n1095) );
NOR2_X1 U983 ( .A1(KEYINPUT60), .A2(n1270), .ZN(n1269) );
INV_X1 U984 ( .A(G122), .ZN(n1270) );
XNOR2_X1 U985 ( .A(G110), .B(KEYINPUT25), .ZN(n1268) );
XOR2_X1 U986 ( .A(n1100), .B(n1099), .Z(n1102) );
AND3_X1 U987 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1099) );
NAND3_X1 U988 ( .A1(G116), .A2(n1274), .A3(G119), .ZN(n1273) );
AND2_X1 U989 ( .A1(n1275), .A2(n1276), .ZN(n1100) );
NAND2_X1 U990 ( .A1(n1277), .A2(G101), .ZN(n1276) );
XOR2_X1 U991 ( .A(KEYINPUT23), .B(n1278), .Z(n1275) );
NOR2_X1 U992 ( .A1(G101), .A2(n1277), .ZN(n1278) );
AND2_X1 U993 ( .A1(n1279), .A2(n1280), .ZN(n1277) );
OR2_X1 U994 ( .A1(G104), .A2(G107), .ZN(n1280) );
NAND2_X1 U995 ( .A1(G107), .A2(n1281), .ZN(n1279) );
XNOR2_X1 U996 ( .A(G104), .B(KEYINPUT17), .ZN(n1281) );
NAND2_X1 U997 ( .A1(KEYINPUT41), .A2(n1151), .ZN(n1267) );
XOR2_X1 U998 ( .A(n1282), .B(n1283), .Z(n1151) );
XOR2_X1 U999 ( .A(G125), .B(n1284), .Z(n1283) );
NOR2_X1 U1000 ( .A1(G953), .A2(n1083), .ZN(n1284) );
INV_X1 U1001 ( .A(G224), .ZN(n1083) );
NOR2_X1 U1002 ( .A1(n1211), .A2(n1285), .ZN(n1206) );
INV_X1 U1003 ( .A(n1210), .ZN(n1285) );
XOR2_X1 U1004 ( .A(n1286), .B(n1061), .Z(n1210) );
NAND2_X1 U1005 ( .A1(G217), .A2(n1217), .ZN(n1061) );
NAND2_X1 U1006 ( .A1(G234), .A2(n1221), .ZN(n1217) );
NAND2_X1 U1007 ( .A1(KEYINPUT37), .A2(n1060), .ZN(n1286) );
NOR2_X1 U1008 ( .A1(n1107), .A2(G902), .ZN(n1060) );
XNOR2_X1 U1009 ( .A(n1287), .B(n1288), .ZN(n1107) );
XOR2_X1 U1010 ( .A(n1237), .B(n1289), .Z(n1288) );
XOR2_X1 U1011 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U1012 ( .A(n1072), .B(KEYINPUT36), .Z(n1237) );
XOR2_X1 U1013 ( .A(G125), .B(G140), .Z(n1072) );
XOR2_X1 U1014 ( .A(n1292), .B(n1293), .Z(n1287) );
XNOR2_X1 U1015 ( .A(n1294), .B(n1295), .ZN(n1293) );
NOR2_X1 U1016 ( .A1(G110), .A2(KEYINPUT27), .ZN(n1295) );
NAND2_X1 U1017 ( .A1(n1256), .A2(G221), .ZN(n1292) );
AND2_X1 U1018 ( .A1(G234), .A2(n1007), .ZN(n1256) );
INV_X1 U1019 ( .A(G953), .ZN(n1007) );
XNOR2_X1 U1020 ( .A(n1055), .B(G472), .ZN(n1211) );
NAND3_X1 U1021 ( .A1(n1296), .A2(n1297), .A3(n1221), .ZN(n1055) );
INV_X1 U1022 ( .A(G902), .ZN(n1221) );
NAND3_X1 U1023 ( .A1(n1298), .A2(n1131), .A3(n1299), .ZN(n1297) );
INV_X1 U1024 ( .A(KEYINPUT29), .ZN(n1299) );
NAND2_X1 U1025 ( .A1(n1300), .A2(KEYINPUT29), .ZN(n1296) );
XOR2_X1 U1026 ( .A(n1131), .B(n1298), .Z(n1300) );
XOR2_X1 U1027 ( .A(n1301), .B(n1134), .Z(n1298) );
NAND4_X1 U1028 ( .A1(n1302), .A2(n1272), .A3(n1303), .A4(n1304), .ZN(n1134) );
NAND3_X1 U1029 ( .A1(KEYINPUT8), .A2(G113), .A3(n1254), .ZN(n1304) );
NAND3_X1 U1030 ( .A1(n1305), .A2(n1274), .A3(G116), .ZN(n1303) );
INV_X1 U1031 ( .A(G113), .ZN(n1274) );
OR2_X1 U1032 ( .A1(KEYINPUT8), .A2(G119), .ZN(n1305) );
NAND3_X1 U1033 ( .A1(G113), .A2(n1254), .A3(G119), .ZN(n1272) );
INV_X1 U1034 ( .A(G116), .ZN(n1254) );
OR2_X1 U1035 ( .A1(n1271), .A2(KEYINPUT8), .ZN(n1302) );
NAND2_X1 U1036 ( .A1(n1306), .A2(n1294), .ZN(n1271) );
INV_X1 U1037 ( .A(G119), .ZN(n1294) );
XNOR2_X1 U1038 ( .A(G113), .B(G116), .ZN(n1306) );
NAND2_X1 U1039 ( .A1(KEYINPUT58), .A2(n1130), .ZN(n1301) );
XOR2_X1 U1040 ( .A(n1148), .B(n1282), .Z(n1130) );
XNOR2_X1 U1041 ( .A(n1307), .B(n1074), .ZN(n1282) );
XNOR2_X1 U1042 ( .A(n1252), .B(n1290), .ZN(n1074) );
XOR2_X1 U1043 ( .A(G128), .B(G146), .Z(n1290) );
INV_X1 U1044 ( .A(n1241), .ZN(n1252) );
XOR2_X1 U1045 ( .A(G143), .B(KEYINPUT4), .Z(n1241) );
XNOR2_X1 U1046 ( .A(KEYINPUT62), .B(KEYINPUT2), .ZN(n1307) );
XOR2_X1 U1047 ( .A(n1071), .B(n1308), .Z(n1148) );
NOR2_X1 U1048 ( .A1(G134), .A2(KEYINPUT45), .ZN(n1308) );
XOR2_X1 U1049 ( .A(G131), .B(n1291), .Z(n1071) );
XOR2_X1 U1050 ( .A(G137), .B(KEYINPUT15), .Z(n1291) );
XNOR2_X1 U1051 ( .A(n1309), .B(G101), .ZN(n1131) );
NAND2_X1 U1052 ( .A1(G210), .A2(n1242), .ZN(n1309) );
NOR2_X1 U1053 ( .A1(G953), .A2(G237), .ZN(n1242) );
endmodule


