//Key = 1100001111100100101001001111001001000101011111110101100100011011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401;

XOR2_X1 U770 ( .A(n1061), .B(n1062), .Z(G9) );
XNOR2_X1 U771 ( .A(G107), .B(KEYINPUT35), .ZN(n1062) );
NOR2_X1 U772 ( .A1(n1063), .A2(n1064), .ZN(G75) );
XOR2_X1 U773 ( .A(n1065), .B(KEYINPUT45), .Z(n1064) );
NAND3_X1 U774 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
NOR4_X1 U775 ( .A1(n1069), .A2(n1070), .A3(n1066), .A4(n1071), .ZN(n1063) );
INV_X1 U776 ( .A(G952), .ZN(n1066) );
NAND3_X1 U777 ( .A1(n1072), .A2(n1068), .A3(n1073), .ZN(n1069) );
XOR2_X1 U778 ( .A(KEYINPUT59), .B(G953), .Z(n1073) );
NAND4_X1 U779 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1068) );
NOR4_X1 U780 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1077) );
XOR2_X1 U781 ( .A(n1082), .B(n1083), .Z(n1081) );
XOR2_X1 U782 ( .A(n1084), .B(KEYINPUT51), .Z(n1082) );
XNOR2_X1 U783 ( .A(n1085), .B(n1086), .ZN(n1080) );
NAND2_X1 U784 ( .A1(KEYINPUT7), .A2(n1087), .ZN(n1085) );
NOR3_X1 U785 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1076) );
NOR3_X1 U786 ( .A1(n1091), .A2(KEYINPUT17), .A3(n1092), .ZN(n1090) );
AND2_X1 U787 ( .A1(n1091), .A2(KEYINPUT17), .ZN(n1089) );
XOR2_X1 U788 ( .A(G475), .B(n1093), .Z(n1088) );
XOR2_X1 U789 ( .A(n1094), .B(n1095), .Z(n1074) );
NOR2_X1 U790 ( .A1(KEYINPUT23), .A2(n1096), .ZN(n1095) );
NAND2_X1 U791 ( .A1(n1097), .A2(n1098), .ZN(n1072) );
NAND2_X1 U792 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND3_X1 U793 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1100) );
NAND2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NAND2_X1 U795 ( .A1(n1075), .A2(n1106), .ZN(n1105) );
OR2_X1 U796 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U797 ( .A1(n1109), .A2(n1110), .ZN(n1104) );
NAND2_X1 U798 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U799 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND3_X1 U800 ( .A1(n1109), .A2(n1115), .A3(n1075), .ZN(n1099) );
NAND3_X1 U801 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
NAND2_X1 U802 ( .A1(n1101), .A2(n1119), .ZN(n1118) );
NAND3_X1 U803 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1117) );
XNOR2_X1 U804 ( .A(n1101), .B(KEYINPUT42), .ZN(n1122) );
XNOR2_X1 U805 ( .A(n1078), .B(KEYINPUT47), .ZN(n1120) );
NAND2_X1 U806 ( .A1(n1103), .A2(n1123), .ZN(n1116) );
NAND2_X1 U807 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND2_X1 U808 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
INV_X1 U809 ( .A(n1128), .ZN(n1097) );
XOR2_X1 U810 ( .A(n1129), .B(n1130), .Z(G72) );
XOR2_X1 U811 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U812 ( .A1(n1133), .A2(n1067), .ZN(n1132) );
NOR2_X1 U813 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NOR2_X1 U814 ( .A1(n1136), .A2(n1137), .ZN(n1131) );
XOR2_X1 U815 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U816 ( .A(n1140), .B(n1141), .Z(n1138) );
NOR2_X1 U817 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XOR2_X1 U818 ( .A(n1144), .B(KEYINPUT60), .Z(n1143) );
NAND2_X1 U819 ( .A1(G131), .A2(n1145), .ZN(n1144) );
NAND2_X1 U820 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NOR3_X1 U821 ( .A1(n1148), .A2(G131), .A3(n1149), .ZN(n1142) );
INV_X1 U822 ( .A(n1147), .ZN(n1148) );
NAND2_X1 U823 ( .A1(n1150), .A2(n1151), .ZN(n1147) );
XOR2_X1 U824 ( .A(n1152), .B(KEYINPUT46), .Z(n1150) );
NAND2_X1 U825 ( .A1(n1153), .A2(n1154), .ZN(n1140) );
NOR2_X1 U826 ( .A1(G900), .A2(n1067), .ZN(n1136) );
AND2_X1 U827 ( .A1(n1070), .A2(n1067), .ZN(n1129) );
NAND2_X1 U828 ( .A1(n1155), .A2(n1156), .ZN(G69) );
NAND2_X1 U829 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND2_X1 U830 ( .A1(G953), .A2(n1159), .ZN(n1158) );
NAND3_X1 U831 ( .A1(n1160), .A2(n1161), .A3(G953), .ZN(n1155) );
NAND2_X1 U832 ( .A1(G898), .A2(G224), .ZN(n1161) );
XOR2_X1 U833 ( .A(KEYINPUT10), .B(n1157), .Z(n1160) );
XNOR2_X1 U834 ( .A(n1162), .B(n1163), .ZN(n1157) );
NOR4_X1 U835 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1163) );
NOR2_X1 U836 ( .A1(KEYINPUT40), .A2(n1168), .ZN(n1167) );
NOR2_X1 U837 ( .A1(G898), .A2(n1067), .ZN(n1166) );
NOR2_X1 U838 ( .A1(n1169), .A2(n1170), .ZN(n1165) );
INV_X1 U839 ( .A(n1171), .ZN(n1170) );
NOR2_X1 U840 ( .A1(n1172), .A2(n1173), .ZN(n1169) );
XOR2_X1 U841 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U842 ( .A1(n1176), .A2(n1177), .ZN(n1172) );
NOR3_X1 U843 ( .A1(n1171), .A2(n1174), .A3(n1175), .ZN(n1164) );
INV_X1 U844 ( .A(KEYINPUT40), .ZN(n1174) );
NAND2_X1 U845 ( .A1(n1067), .A2(n1071), .ZN(n1162) );
NOR2_X1 U846 ( .A1(n1178), .A2(n1179), .ZN(G66) );
XOR2_X1 U847 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U848 ( .A1(n1182), .A2(KEYINPUT20), .ZN(n1181) );
NOR2_X1 U849 ( .A1(n1091), .A2(n1183), .ZN(n1182) );
NOR2_X1 U850 ( .A1(n1178), .A2(n1184), .ZN(G63) );
NOR3_X1 U851 ( .A1(n1083), .A2(n1185), .A3(n1186), .ZN(n1184) );
NOR3_X1 U852 ( .A1(n1187), .A2(n1084), .A3(n1183), .ZN(n1186) );
INV_X1 U853 ( .A(n1188), .ZN(n1187) );
NOR2_X1 U854 ( .A1(n1189), .A2(n1188), .ZN(n1185) );
NOR2_X1 U855 ( .A1(n1190), .A2(n1084), .ZN(n1189) );
NOR2_X1 U856 ( .A1(n1071), .A2(n1070), .ZN(n1190) );
NOR2_X1 U857 ( .A1(n1178), .A2(n1191), .ZN(G60) );
XNOR2_X1 U858 ( .A(n1192), .B(n1193), .ZN(n1191) );
NOR2_X1 U859 ( .A1(n1194), .A2(n1183), .ZN(n1193) );
INV_X1 U860 ( .A(G475), .ZN(n1194) );
XOR2_X1 U861 ( .A(n1195), .B(n1196), .Z(G6) );
NOR2_X1 U862 ( .A1(n1178), .A2(n1197), .ZN(G57) );
XOR2_X1 U863 ( .A(n1198), .B(n1199), .Z(n1197) );
NAND2_X1 U864 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
NAND2_X1 U865 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XOR2_X1 U866 ( .A(KEYINPUT8), .B(n1204), .Z(n1200) );
NOR2_X1 U867 ( .A1(n1203), .A2(n1205), .ZN(n1204) );
XOR2_X1 U868 ( .A(KEYINPUT2), .B(n1202), .Z(n1205) );
NOR2_X1 U869 ( .A1(n1183), .A2(n1087), .ZN(n1202) );
NOR2_X1 U870 ( .A1(n1178), .A2(n1206), .ZN(G54) );
XOR2_X1 U871 ( .A(n1207), .B(n1208), .Z(n1206) );
XOR2_X1 U872 ( .A(n1209), .B(n1210), .Z(n1208) );
XNOR2_X1 U873 ( .A(n1211), .B(n1212), .ZN(n1210) );
NOR2_X1 U874 ( .A1(KEYINPUT38), .A2(n1213), .ZN(n1212) );
NAND2_X1 U875 ( .A1(KEYINPUT9), .A2(n1214), .ZN(n1211) );
XOR2_X1 U876 ( .A(n1215), .B(n1216), .Z(n1207) );
XOR2_X1 U877 ( .A(G140), .B(G110), .Z(n1216) );
XOR2_X1 U878 ( .A(n1217), .B(n1218), .Z(n1215) );
NOR2_X1 U879 ( .A1(n1219), .A2(n1183), .ZN(n1218) );
INV_X1 U880 ( .A(G469), .ZN(n1219) );
NOR3_X1 U881 ( .A1(n1178), .A2(n1220), .A3(n1221), .ZN(G51) );
NOR2_X1 U882 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
XOR2_X1 U883 ( .A(KEYINPUT48), .B(n1224), .Z(n1223) );
NOR2_X1 U884 ( .A1(n1225), .A2(n1226), .ZN(n1220) );
XNOR2_X1 U885 ( .A(n1224), .B(KEYINPUT34), .ZN(n1226) );
XNOR2_X1 U886 ( .A(n1227), .B(n1228), .ZN(n1224) );
NOR3_X1 U887 ( .A1(n1183), .A2(KEYINPUT29), .A3(n1094), .ZN(n1228) );
NAND2_X1 U888 ( .A1(G902), .A2(n1229), .ZN(n1183) );
OR2_X1 U889 ( .A1(n1070), .A2(n1071), .ZN(n1229) );
NAND4_X1 U890 ( .A1(n1196), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1071) );
AND4_X1 U891 ( .A1(n1061), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1232) );
NAND3_X1 U892 ( .A1(n1108), .A2(n1101), .A3(n1236), .ZN(n1061) );
NAND2_X1 U893 ( .A1(n1109), .A2(n1237), .ZN(n1231) );
NAND2_X1 U894 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND3_X1 U895 ( .A1(n1240), .A2(n1127), .A3(n1241), .ZN(n1239) );
NAND2_X1 U896 ( .A1(n1242), .A2(n1236), .ZN(n1238) );
NAND3_X1 U897 ( .A1(n1236), .A2(n1101), .A3(n1107), .ZN(n1196) );
NAND4_X1 U898 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1070) );
NOR4_X1 U899 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1246) );
AND2_X1 U900 ( .A1(n1251), .A2(n1252), .ZN(n1245) );
NAND2_X1 U901 ( .A1(n1253), .A2(n1254), .ZN(n1227) );
NAND2_X1 U902 ( .A1(n1255), .A2(n1213), .ZN(n1254) );
XOR2_X1 U903 ( .A(n1256), .B(KEYINPUT5), .Z(n1255) );
NAND2_X1 U904 ( .A1(n1257), .A2(n1139), .ZN(n1253) );
XOR2_X1 U905 ( .A(n1256), .B(KEYINPUT33), .Z(n1257) );
INV_X1 U906 ( .A(n1222), .ZN(n1225) );
NOR2_X1 U907 ( .A1(n1067), .A2(G952), .ZN(n1178) );
XNOR2_X1 U908 ( .A(G146), .B(n1243), .ZN(G48) );
NAND2_X1 U909 ( .A1(n1258), .A2(n1107), .ZN(n1243) );
XOR2_X1 U910 ( .A(n1244), .B(n1259), .Z(G45) );
XNOR2_X1 U911 ( .A(G143), .B(KEYINPUT36), .ZN(n1259) );
NAND4_X1 U912 ( .A1(n1260), .A2(n1119), .A3(n1261), .A4(n1262), .ZN(n1244) );
XOR2_X1 U913 ( .A(n1263), .B(n1252), .Z(G42) );
NAND4_X1 U914 ( .A1(n1264), .A2(n1103), .A3(n1126), .A4(n1107), .ZN(n1252) );
XOR2_X1 U915 ( .A(n1151), .B(n1265), .Z(G39) );
NAND2_X1 U916 ( .A1(KEYINPUT27), .A2(n1250), .ZN(n1265) );
AND4_X1 U917 ( .A1(n1264), .A2(n1103), .A3(n1109), .A4(n1240), .ZN(n1250) );
XOR2_X1 U918 ( .A(G134), .B(n1249), .Z(G36) );
AND3_X1 U919 ( .A1(n1260), .A2(n1108), .A3(n1103), .ZN(n1249) );
XOR2_X1 U920 ( .A(G131), .B(n1248), .Z(G33) );
AND3_X1 U921 ( .A1(n1260), .A2(n1107), .A3(n1103), .ZN(n1248) );
NOR2_X1 U922 ( .A1(n1266), .A2(n1078), .ZN(n1103) );
INV_X1 U923 ( .A(n1121), .ZN(n1266) );
NOR3_X1 U924 ( .A1(n1111), .A2(n1267), .A3(n1124), .ZN(n1260) );
XOR2_X1 U925 ( .A(n1268), .B(n1251), .Z(G30) );
NAND2_X1 U926 ( .A1(n1258), .A2(n1108), .ZN(n1251) );
AND3_X1 U927 ( .A1(n1119), .A2(n1240), .A3(n1264), .ZN(n1258) );
NOR3_X1 U928 ( .A1(n1269), .A2(n1267), .A3(n1111), .ZN(n1264) );
XOR2_X1 U929 ( .A(n1270), .B(n1271), .Z(G3) );
NAND3_X1 U930 ( .A1(n1242), .A2(n1236), .A3(n1272), .ZN(n1271) );
XNOR2_X1 U931 ( .A(KEYINPUT37), .B(n1109), .ZN(n1272) );
XNOR2_X1 U932 ( .A(n1247), .B(n1273), .ZN(G27) );
NAND2_X1 U933 ( .A1(KEYINPUT44), .A2(G125), .ZN(n1273) );
AND4_X1 U934 ( .A1(n1126), .A2(n1075), .A3(n1107), .A4(n1274), .ZN(n1247) );
NOR3_X1 U935 ( .A1(n1275), .A2(n1267), .A3(n1269), .ZN(n1274) );
AND2_X1 U936 ( .A1(n1276), .A2(n1128), .ZN(n1267) );
NAND4_X1 U937 ( .A1(G953), .A2(G902), .A3(n1277), .A4(n1135), .ZN(n1276) );
INV_X1 U938 ( .A(G900), .ZN(n1135) );
XOR2_X1 U939 ( .A(n1278), .B(n1230), .Z(G24) );
NAND4_X1 U940 ( .A1(n1241), .A2(n1101), .A3(n1261), .A4(n1262), .ZN(n1230) );
NOR2_X1 U941 ( .A1(n1127), .A2(n1240), .ZN(n1101) );
XNOR2_X1 U942 ( .A(G119), .B(n1279), .ZN(G21) );
NAND4_X1 U943 ( .A1(n1280), .A2(n1109), .A3(n1075), .A4(n1281), .ZN(n1279) );
NOR3_X1 U944 ( .A1(n1126), .A2(n1282), .A3(n1269), .ZN(n1281) );
XOR2_X1 U945 ( .A(KEYINPUT57), .B(n1119), .Z(n1280) );
XNOR2_X1 U946 ( .A(G116), .B(n1235), .ZN(G18) );
NAND3_X1 U947 ( .A1(n1242), .A2(n1108), .A3(n1241), .ZN(n1235) );
NOR2_X1 U948 ( .A1(n1261), .A2(n1283), .ZN(n1108) );
XOR2_X1 U949 ( .A(n1234), .B(n1284), .Z(G15) );
XOR2_X1 U950 ( .A(n1285), .B(KEYINPUT22), .Z(n1284) );
NAND3_X1 U951 ( .A1(n1242), .A2(n1107), .A3(n1241), .ZN(n1234) );
AND3_X1 U952 ( .A1(n1119), .A2(n1286), .A3(n1075), .ZN(n1241) );
NOR2_X1 U953 ( .A1(n1287), .A2(n1113), .ZN(n1075) );
INV_X1 U954 ( .A(n1114), .ZN(n1287) );
INV_X1 U955 ( .A(n1124), .ZN(n1242) );
NAND2_X1 U956 ( .A1(n1269), .A2(n1240), .ZN(n1124) );
INV_X1 U957 ( .A(n1126), .ZN(n1240) );
XOR2_X1 U958 ( .A(n1233), .B(n1288), .Z(G12) );
NAND2_X1 U959 ( .A1(KEYINPUT63), .A2(G110), .ZN(n1288) );
NAND4_X1 U960 ( .A1(n1126), .A2(n1236), .A3(n1109), .A4(n1127), .ZN(n1233) );
INV_X1 U961 ( .A(n1269), .ZN(n1127) );
NOR2_X1 U962 ( .A1(n1079), .A2(n1289), .ZN(n1269) );
NOR2_X1 U963 ( .A1(n1091), .A2(n1092), .ZN(n1289) );
AND2_X1 U964 ( .A1(n1092), .A2(n1091), .ZN(n1079) );
NAND2_X1 U965 ( .A1(G217), .A2(n1290), .ZN(n1091) );
AND2_X1 U966 ( .A1(n1180), .A2(n1291), .ZN(n1092) );
XOR2_X1 U967 ( .A(n1292), .B(n1293), .Z(n1180) );
XOR2_X1 U968 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U969 ( .A(n1296), .B(n1297), .Z(n1295) );
NAND3_X1 U970 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1297) );
NAND2_X1 U971 ( .A1(KEYINPUT61), .A2(G119), .ZN(n1300) );
NAND3_X1 U972 ( .A1(n1301), .A2(n1302), .A3(n1268), .ZN(n1299) );
INV_X1 U973 ( .A(KEYINPUT61), .ZN(n1302) );
OR2_X1 U974 ( .A1(n1268), .A2(n1301), .ZN(n1298) );
NOR2_X1 U975 ( .A1(G119), .A2(KEYINPUT11), .ZN(n1301) );
NAND2_X1 U976 ( .A1(KEYINPUT26), .A2(n1303), .ZN(n1296) );
XOR2_X1 U977 ( .A(KEYINPUT1), .B(G110), .Z(n1303) );
AND2_X1 U978 ( .A1(G221), .A2(n1304), .ZN(n1294) );
XOR2_X1 U979 ( .A(n1305), .B(n1306), .Z(n1292) );
XOR2_X1 U980 ( .A(KEYINPUT31), .B(G146), .Z(n1306) );
XOR2_X1 U981 ( .A(n1151), .B(n1307), .Z(n1305) );
NOR2_X1 U982 ( .A1(KEYINPUT32), .A2(n1308), .ZN(n1307) );
NOR3_X1 U983 ( .A1(n1309), .A2(n1310), .A3(n1311), .ZN(n1308) );
NOR2_X1 U984 ( .A1(n1312), .A2(n1154), .ZN(n1311) );
INV_X1 U985 ( .A(KEYINPUT52), .ZN(n1312) );
NOR2_X1 U986 ( .A1(KEYINPUT52), .A2(n1313), .ZN(n1310) );
INV_X1 U987 ( .A(n1153), .ZN(n1309) );
NAND2_X1 U988 ( .A1(n1314), .A2(n1315), .ZN(n1109) );
NAND2_X1 U989 ( .A1(n1107), .A2(n1316), .ZN(n1315) );
AND2_X1 U990 ( .A1(n1283), .A2(n1261), .ZN(n1107) );
INV_X1 U991 ( .A(n1262), .ZN(n1283) );
OR3_X1 U992 ( .A1(n1262), .A2(n1261), .A3(n1316), .ZN(n1314) );
INV_X1 U993 ( .A(KEYINPUT18), .ZN(n1316) );
XNOR2_X1 U994 ( .A(n1317), .B(G475), .ZN(n1261) );
NAND2_X1 U995 ( .A1(KEYINPUT21), .A2(n1093), .ZN(n1317) );
AND2_X1 U996 ( .A1(n1291), .A2(n1192), .ZN(n1093) );
NAND3_X1 U997 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1192) );
NAND2_X1 U998 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
OR3_X1 U999 ( .A1(n1322), .A2(n1321), .A3(n1323), .ZN(n1319) );
INV_X1 U1000 ( .A(KEYINPUT41), .ZN(n1322) );
NAND2_X1 U1001 ( .A1(n1323), .A2(n1324), .ZN(n1318) );
NAND2_X1 U1002 ( .A1(n1325), .A2(KEYINPUT41), .ZN(n1324) );
XOR2_X1 U1003 ( .A(n1321), .B(KEYINPUT6), .Z(n1325) );
XOR2_X1 U1004 ( .A(n1326), .B(n1327), .Z(n1321) );
XNOR2_X1 U1005 ( .A(n1328), .B(n1329), .ZN(n1327) );
NAND2_X1 U1006 ( .A1(n1330), .A2(n1154), .ZN(n1328) );
NAND2_X1 U1007 ( .A1(G140), .A2(n1313), .ZN(n1154) );
XOR2_X1 U1008 ( .A(n1153), .B(KEYINPUT54), .Z(n1330) );
NAND2_X1 U1009 ( .A1(G125), .A2(n1263), .ZN(n1153) );
INV_X1 U1010 ( .A(G140), .ZN(n1263) );
XOR2_X1 U1011 ( .A(n1331), .B(n1332), .Z(n1326) );
XOR2_X1 U1012 ( .A(KEYINPUT39), .B(G131), .Z(n1332) );
NAND2_X1 U1013 ( .A1(n1333), .A2(G214), .ZN(n1331) );
XNOR2_X1 U1014 ( .A(n1334), .B(G104), .ZN(n1323) );
NAND3_X1 U1015 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1334) );
NAND2_X1 U1016 ( .A1(KEYINPUT56), .A2(n1338), .ZN(n1337) );
NAND3_X1 U1017 ( .A1(n1339), .A2(n1340), .A3(n1285), .ZN(n1336) );
INV_X1 U1018 ( .A(KEYINPUT56), .ZN(n1340) );
OR2_X1 U1019 ( .A1(n1285), .A2(n1339), .ZN(n1335) );
NOR2_X1 U1020 ( .A1(KEYINPUT19), .A2(n1338), .ZN(n1339) );
XOR2_X1 U1021 ( .A(n1278), .B(KEYINPUT30), .Z(n1338) );
INV_X1 U1022 ( .A(G113), .ZN(n1285) );
NAND2_X1 U1023 ( .A1(n1341), .A2(n1342), .ZN(n1262) );
OR2_X1 U1024 ( .A1(n1343), .A2(n1083), .ZN(n1342) );
XOR2_X1 U1025 ( .A(n1344), .B(KEYINPUT12), .Z(n1341) );
NAND2_X1 U1026 ( .A1(n1083), .A2(n1343), .ZN(n1344) );
XNOR2_X1 U1027 ( .A(n1084), .B(KEYINPUT0), .ZN(n1343) );
INV_X1 U1028 ( .A(G478), .ZN(n1084) );
NOR2_X1 U1029 ( .A1(n1188), .A2(G902), .ZN(n1083) );
XOR2_X1 U1030 ( .A(n1345), .B(n1346), .Z(n1188) );
NOR2_X1 U1031 ( .A1(KEYINPUT14), .A2(n1347), .ZN(n1346) );
XOR2_X1 U1032 ( .A(n1348), .B(n1349), .Z(n1347) );
XOR2_X1 U1033 ( .A(G107), .B(n1350), .Z(n1349) );
XOR2_X1 U1034 ( .A(G122), .B(G116), .Z(n1350) );
XOR2_X1 U1035 ( .A(n1351), .B(n1352), .Z(n1348) );
XOR2_X1 U1036 ( .A(G134), .B(G128), .Z(n1352) );
XNOR2_X1 U1037 ( .A(G143), .B(KEYINPUT28), .ZN(n1351) );
NAND2_X1 U1038 ( .A1(G217), .A2(n1304), .ZN(n1345) );
AND2_X1 U1039 ( .A1(G234), .A2(n1067), .ZN(n1304) );
NOR3_X1 U1040 ( .A1(n1111), .A2(n1282), .A3(n1275), .ZN(n1236) );
INV_X1 U1041 ( .A(n1119), .ZN(n1275) );
NOR2_X1 U1042 ( .A1(n1121), .A2(n1078), .ZN(n1119) );
AND2_X1 U1043 ( .A1(G214), .A2(n1353), .ZN(n1078) );
XNOR2_X1 U1044 ( .A(KEYINPUT49), .B(n1354), .ZN(n1353) );
XNOR2_X1 U1045 ( .A(n1096), .B(n1094), .ZN(n1121) );
NAND2_X1 U1046 ( .A1(G210), .A2(n1354), .ZN(n1094) );
OR2_X1 U1047 ( .A1(G902), .A2(G237), .ZN(n1354) );
NAND2_X1 U1048 ( .A1(n1355), .A2(n1291), .ZN(n1096) );
XOR2_X1 U1049 ( .A(n1256), .B(n1356), .Z(n1355) );
XOR2_X1 U1050 ( .A(n1222), .B(n1213), .Z(n1356) );
NAND2_X1 U1051 ( .A1(n1168), .A2(n1357), .ZN(n1222) );
NAND2_X1 U1052 ( .A1(n1171), .A2(n1358), .ZN(n1357) );
OR2_X1 U1053 ( .A1(n1358), .A2(n1171), .ZN(n1168) );
XNOR2_X1 U1054 ( .A(n1278), .B(G110), .ZN(n1171) );
INV_X1 U1055 ( .A(G122), .ZN(n1278) );
NAND2_X1 U1056 ( .A1(n1175), .A2(n1359), .ZN(n1358) );
OR2_X1 U1057 ( .A1(n1177), .A2(n1176), .ZN(n1359) );
NAND2_X1 U1058 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XNOR2_X1 U1059 ( .A(n1360), .B(n1361), .ZN(n1177) );
XOR2_X1 U1060 ( .A(G107), .B(G101), .Z(n1361) );
NAND2_X1 U1061 ( .A1(KEYINPUT25), .A2(n1195), .ZN(n1360) );
INV_X1 U1062 ( .A(G104), .ZN(n1195) );
XOR2_X1 U1063 ( .A(n1362), .B(n1363), .Z(n1176) );
XOR2_X1 U1064 ( .A(G116), .B(G113), .Z(n1363) );
NAND2_X1 U1065 ( .A1(KEYINPUT16), .A2(G119), .ZN(n1362) );
XOR2_X1 U1066 ( .A(n1313), .B(n1364), .Z(n1256) );
NOR2_X1 U1067 ( .A1(G953), .A2(n1159), .ZN(n1364) );
INV_X1 U1068 ( .A(G224), .ZN(n1159) );
INV_X1 U1069 ( .A(G125), .ZN(n1313) );
INV_X1 U1070 ( .A(n1286), .ZN(n1282) );
NAND2_X1 U1071 ( .A1(n1128), .A2(n1365), .ZN(n1286) );
NAND4_X1 U1072 ( .A1(G953), .A2(G902), .A3(n1277), .A4(n1366), .ZN(n1365) );
INV_X1 U1073 ( .A(G898), .ZN(n1366) );
NAND3_X1 U1074 ( .A1(n1277), .A2(n1067), .A3(G952), .ZN(n1128) );
INV_X1 U1075 ( .A(G953), .ZN(n1067) );
NAND2_X1 U1076 ( .A1(G237), .A2(G234), .ZN(n1277) );
OR2_X1 U1077 ( .A1(n1114), .A2(n1113), .ZN(n1111) );
AND2_X1 U1078 ( .A1(G221), .A2(n1290), .ZN(n1113) );
NAND2_X1 U1079 ( .A1(G234), .A2(n1291), .ZN(n1290) );
XOR2_X1 U1080 ( .A(n1367), .B(G469), .Z(n1114) );
NAND2_X1 U1081 ( .A1(n1368), .A2(n1291), .ZN(n1367) );
XOR2_X1 U1082 ( .A(n1369), .B(n1370), .Z(n1368) );
XOR2_X1 U1083 ( .A(n1217), .B(n1371), .Z(n1370) );
NAND3_X1 U1084 ( .A1(n1372), .A2(n1373), .A3(n1374), .ZN(n1217) );
NAND2_X1 U1085 ( .A1(n1375), .A2(G101), .ZN(n1374) );
NAND2_X1 U1086 ( .A1(n1376), .A2(n1377), .ZN(n1373) );
INV_X1 U1087 ( .A(KEYINPUT24), .ZN(n1377) );
NAND2_X1 U1088 ( .A1(n1378), .A2(n1270), .ZN(n1376) );
INV_X1 U1089 ( .A(G101), .ZN(n1270) );
XNOR2_X1 U1090 ( .A(KEYINPUT4), .B(n1375), .ZN(n1378) );
NAND2_X1 U1091 ( .A1(KEYINPUT24), .A2(n1379), .ZN(n1372) );
NAND2_X1 U1092 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
NAND2_X1 U1093 ( .A1(KEYINPUT4), .A2(n1375), .ZN(n1381) );
OR3_X1 U1094 ( .A1(G101), .A2(KEYINPUT4), .A3(n1375), .ZN(n1380) );
XOR2_X1 U1095 ( .A(n1382), .B(n1383), .Z(n1375) );
XOR2_X1 U1096 ( .A(G107), .B(G104), .Z(n1383) );
XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(KEYINPUT43), .ZN(n1382) );
XOR2_X1 U1098 ( .A(n1384), .B(n1214), .Z(n1369) );
NOR2_X1 U1099 ( .A1(n1134), .A2(G953), .ZN(n1214) );
INV_X1 U1100 ( .A(G227), .ZN(n1134) );
NAND3_X1 U1101 ( .A1(n1385), .A2(n1386), .A3(n1387), .ZN(n1384) );
NAND2_X1 U1102 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
INV_X1 U1103 ( .A(KEYINPUT55), .ZN(n1389) );
NAND3_X1 U1104 ( .A1(KEYINPUT55), .A2(n1390), .A3(n1391), .ZN(n1386) );
OR2_X1 U1105 ( .A1(n1391), .A2(n1390), .ZN(n1385) );
NOR2_X1 U1106 ( .A1(KEYINPUT50), .A2(n1388), .ZN(n1390) );
XOR2_X1 U1107 ( .A(G140), .B(KEYINPUT53), .Z(n1388) );
INV_X1 U1108 ( .A(G110), .ZN(n1391) );
XOR2_X1 U1109 ( .A(n1087), .B(n1392), .Z(n1126) );
NOR2_X1 U1110 ( .A1(KEYINPUT3), .A2(n1086), .ZN(n1392) );
NAND2_X1 U1111 ( .A1(n1393), .A2(n1394), .ZN(n1086) );
XOR2_X1 U1112 ( .A(n1199), .B(n1203), .Z(n1394) );
XNOR2_X1 U1113 ( .A(n1395), .B(n1396), .ZN(n1203) );
XOR2_X1 U1114 ( .A(G116), .B(n1397), .Z(n1396) );
XOR2_X1 U1115 ( .A(KEYINPUT62), .B(G119), .Z(n1397) );
XOR2_X1 U1116 ( .A(n1371), .B(G113), .Z(n1395) );
XOR2_X1 U1117 ( .A(n1209), .B(n1139), .Z(n1371) );
INV_X1 U1118 ( .A(n1213), .ZN(n1139) );
XOR2_X1 U1119 ( .A(n1268), .B(n1329), .Z(n1213) );
XOR2_X1 U1120 ( .A(G143), .B(G146), .Z(n1329) );
INV_X1 U1121 ( .A(G128), .ZN(n1268) );
XOR2_X1 U1122 ( .A(n1398), .B(G131), .Z(n1209) );
NAND2_X1 U1123 ( .A1(n1399), .A2(n1400), .ZN(n1398) );
NAND2_X1 U1124 ( .A1(G134), .A2(n1151), .ZN(n1400) );
INV_X1 U1125 ( .A(G137), .ZN(n1151) );
XOR2_X1 U1126 ( .A(KEYINPUT13), .B(n1149), .Z(n1399) );
INV_X1 U1127 ( .A(n1146), .ZN(n1149) );
NAND2_X1 U1128 ( .A1(G137), .A2(n1152), .ZN(n1146) );
INV_X1 U1129 ( .A(G134), .ZN(n1152) );
XNOR2_X1 U1130 ( .A(n1401), .B(G101), .ZN(n1199) );
NAND2_X1 U1131 ( .A1(n1333), .A2(G210), .ZN(n1401) );
NOR2_X1 U1132 ( .A1(G953), .A2(G237), .ZN(n1333) );
XOR2_X1 U1133 ( .A(n1291), .B(KEYINPUT15), .Z(n1393) );
INV_X1 U1134 ( .A(G902), .ZN(n1291) );
INV_X1 U1135 ( .A(G472), .ZN(n1087) );
endmodule


