//Key = 0111111010000111100100111110000100111001111010010001111100010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305;

XNOR2_X1 U725 ( .A(G107), .B(n1001), .ZN(G9) );
NOR2_X1 U726 ( .A1(n1002), .A2(n1003), .ZN(G75) );
NOR3_X1 U727 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1003) );
NAND3_X1 U728 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1004) );
NAND2_X1 U729 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND2_X1 U730 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND4_X1 U731 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1013) );
NAND2_X1 U732 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND2_X1 U733 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
INV_X1 U734 ( .A(n1022), .ZN(n1018) );
NAND2_X1 U735 ( .A1(n1023), .A2(n1024), .ZN(n1012) );
NAND2_X1 U736 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U737 ( .A1(n1015), .A2(n1027), .ZN(n1026) );
NAND2_X1 U738 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND3_X1 U739 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
INV_X1 U740 ( .A(KEYINPUT15), .ZN(n1031) );
NAND2_X1 U741 ( .A1(n1014), .A2(n1033), .ZN(n1028) );
NAND2_X1 U742 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U743 ( .A1(n1016), .A2(n1030), .ZN(n1025) );
NAND3_X1 U744 ( .A1(n1036), .A2(n1037), .A3(n1016), .ZN(n1030) );
NAND2_X1 U745 ( .A1(n1015), .A2(n1038), .ZN(n1037) );
NAND2_X1 U746 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U747 ( .A1(KEYINPUT15), .A2(n1032), .ZN(n1040) );
NAND2_X1 U748 ( .A1(n1014), .A2(n1041), .ZN(n1036) );
NAND2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
INV_X1 U751 ( .A(n1046), .ZN(n1010) );
NOR3_X1 U752 ( .A1(n1047), .A2(G953), .A3(G952), .ZN(n1002) );
INV_X1 U753 ( .A(n1007), .ZN(n1047) );
NAND4_X1 U754 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1007) );
NOR4_X1 U755 ( .A1(n1020), .A2(n1044), .A3(n1052), .A4(n1053), .ZN(n1051) );
XOR2_X1 U756 ( .A(n1054), .B(n1055), .Z(n1052) );
NOR2_X1 U757 ( .A1(G469), .A2(KEYINPUT62), .ZN(n1055) );
NOR3_X1 U758 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1050) );
NOR2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR2_X1 U760 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U761 ( .A1(KEYINPUT24), .A2(n1063), .ZN(n1062) );
NOR2_X1 U762 ( .A1(n1064), .A2(n1065), .ZN(n1061) );
INV_X1 U763 ( .A(KEYINPUT24), .ZN(n1065) );
NOR2_X1 U764 ( .A1(n1063), .A2(n1066), .ZN(n1064) );
NOR3_X1 U765 ( .A1(G475), .A2(n1063), .A3(n1066), .ZN(n1057) );
INV_X1 U766 ( .A(KEYINPUT3), .ZN(n1066) );
XOR2_X1 U767 ( .A(n1067), .B(KEYINPUT14), .Z(n1063) );
XNOR2_X1 U768 ( .A(G472), .B(n1068), .ZN(n1056) );
XNOR2_X1 U769 ( .A(n1069), .B(KEYINPUT60), .ZN(n1049) );
XOR2_X1 U770 ( .A(n1070), .B(n1071), .Z(n1048) );
XOR2_X1 U771 ( .A(n1072), .B(KEYINPUT9), .Z(n1070) );
XOR2_X1 U772 ( .A(n1073), .B(n1074), .Z(G72) );
XOR2_X1 U773 ( .A(n1075), .B(n1076), .Z(n1074) );
NAND2_X1 U774 ( .A1(n1008), .A2(n1005), .ZN(n1076) );
NAND2_X1 U775 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NAND2_X1 U776 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XNOR2_X1 U777 ( .A(G953), .B(KEYINPUT47), .ZN(n1079) );
XOR2_X1 U778 ( .A(n1081), .B(n1082), .Z(n1077) );
XOR2_X1 U779 ( .A(n1083), .B(n1084), .Z(n1082) );
XNOR2_X1 U780 ( .A(n1085), .B(n1086), .ZN(n1081) );
NOR2_X1 U781 ( .A1(n1087), .A2(n1008), .ZN(n1073) );
NOR2_X1 U782 ( .A1(n1088), .A2(n1080), .ZN(n1087) );
NAND2_X1 U783 ( .A1(n1089), .A2(n1090), .ZN(G69) );
NAND2_X1 U784 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U785 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
INV_X1 U786 ( .A(n1095), .ZN(n1093) );
NAND2_X1 U787 ( .A1(n1096), .A2(n1094), .ZN(n1089) );
NAND2_X1 U788 ( .A1(G953), .A2(n1097), .ZN(n1094) );
INV_X1 U789 ( .A(n1092), .ZN(n1096) );
NAND2_X1 U790 ( .A1(KEYINPUT36), .A2(n1098), .ZN(n1092) );
XOR2_X1 U791 ( .A(n1099), .B(n1100), .Z(n1098) );
AND2_X1 U792 ( .A1(n1006), .A2(n1008), .ZN(n1100) );
NOR2_X1 U793 ( .A1(n1095), .A2(n1101), .ZN(n1099) );
XOR2_X1 U794 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U795 ( .A(n1104), .B(KEYINPUT1), .Z(n1103) );
NAND2_X1 U796 ( .A1(KEYINPUT40), .A2(n1105), .ZN(n1104) );
INV_X1 U797 ( .A(n1106), .ZN(n1105) );
NOR2_X1 U798 ( .A1(n1107), .A2(n1108), .ZN(G66) );
XOR2_X1 U799 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND3_X1 U800 ( .A1(n1111), .A2(G217), .A3(n1112), .ZN(n1109) );
XOR2_X1 U801 ( .A(n1113), .B(KEYINPUT17), .Z(n1112) );
NOR2_X1 U802 ( .A1(n1107), .A2(n1114), .ZN(G63) );
XOR2_X1 U803 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U804 ( .A1(n1111), .A2(G478), .ZN(n1115) );
NOR2_X1 U805 ( .A1(n1107), .A2(n1117), .ZN(G60) );
NOR3_X1 U806 ( .A1(n1067), .A2(n1118), .A3(n1119), .ZN(n1117) );
AND3_X1 U807 ( .A1(n1120), .A2(G475), .A3(n1111), .ZN(n1119) );
NOR2_X1 U808 ( .A1(n1121), .A2(n1120), .ZN(n1118) );
NOR2_X1 U809 ( .A1(n1122), .A2(n1059), .ZN(n1121) );
NOR2_X1 U810 ( .A1(n1005), .A2(n1006), .ZN(n1122) );
XNOR2_X1 U811 ( .A(G104), .B(n1123), .ZN(G6) );
NOR2_X1 U812 ( .A1(n1107), .A2(n1124), .ZN(G57) );
XOR2_X1 U813 ( .A(n1125), .B(n1126), .Z(n1124) );
XNOR2_X1 U814 ( .A(n1106), .B(n1127), .ZN(n1126) );
NAND2_X1 U815 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U816 ( .A1(KEYINPUT4), .A2(n1130), .ZN(n1129) );
OR2_X1 U817 ( .A1(KEYINPUT2), .A2(n1130), .ZN(n1128) );
XNOR2_X1 U818 ( .A(n1131), .B(G101), .ZN(n1130) );
NAND2_X1 U819 ( .A1(KEYINPUT26), .A2(n1132), .ZN(n1131) );
XOR2_X1 U820 ( .A(n1133), .B(n1134), .Z(n1125) );
XNOR2_X1 U821 ( .A(KEYINPUT0), .B(n1135), .ZN(n1134) );
NOR2_X1 U822 ( .A1(KEYINPUT18), .A2(n1136), .ZN(n1135) );
XOR2_X1 U823 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U824 ( .A1(KEYINPUT34), .A2(n1139), .ZN(n1137) );
NAND2_X1 U825 ( .A1(n1111), .A2(G472), .ZN(n1133) );
NOR2_X1 U826 ( .A1(n1107), .A2(n1140), .ZN(G54) );
XNOR2_X1 U827 ( .A(n1141), .B(n1142), .ZN(n1140) );
XOR2_X1 U828 ( .A(n1143), .B(n1144), .Z(n1141) );
NAND2_X1 U829 ( .A1(n1145), .A2(n1111), .ZN(n1143) );
XNOR2_X1 U830 ( .A(G469), .B(KEYINPUT59), .ZN(n1145) );
NOR2_X1 U831 ( .A1(n1107), .A2(n1146), .ZN(G51) );
XOR2_X1 U832 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U833 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U834 ( .A(n1151), .B(KEYINPUT19), .Z(n1147) );
NAND2_X1 U835 ( .A1(n1111), .A2(n1071), .ZN(n1151) );
AND2_X1 U836 ( .A1(G902), .A2(n1152), .ZN(n1111) );
OR2_X1 U837 ( .A1(n1006), .A2(n1005), .ZN(n1152) );
NAND4_X1 U838 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1005) );
NOR4_X1 U839 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1156) );
NOR3_X1 U840 ( .A1(n1161), .A2(n1034), .A3(n1162), .ZN(n1158) );
XNOR2_X1 U841 ( .A(KEYINPUT49), .B(n1163), .ZN(n1161) );
NOR2_X1 U842 ( .A1(n1164), .A2(n1165), .ZN(n1157) );
XNOR2_X1 U843 ( .A(n1166), .B(KEYINPUT56), .ZN(n1164) );
NOR3_X1 U844 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1155) );
AND4_X1 U845 ( .A1(KEYINPUT29), .A2(n1170), .A3(n1171), .A4(n1022), .ZN(n1169) );
NAND2_X1 U846 ( .A1(n1053), .A2(n1172), .ZN(n1171) );
NOR2_X1 U847 ( .A1(KEYINPUT29), .A2(n1173), .ZN(n1168) );
INV_X1 U848 ( .A(n1174), .ZN(n1167) );
INV_X1 U849 ( .A(n1175), .ZN(n1153) );
NAND2_X1 U850 ( .A1(n1176), .A2(n1177), .ZN(n1006) );
AND4_X1 U851 ( .A1(n1178), .A2(n1001), .A3(n1179), .A4(n1180), .ZN(n1177) );
NAND3_X1 U852 ( .A1(n1032), .A2(n1016), .A3(n1181), .ZN(n1001) );
AND4_X1 U853 ( .A1(n1182), .A2(n1183), .A3(n1123), .A4(n1184), .ZN(n1176) );
OR2_X1 U854 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XNOR2_X1 U855 ( .A(n1187), .B(KEYINPUT30), .ZN(n1185) );
NAND3_X1 U856 ( .A1(n1181), .A2(n1016), .A3(n1188), .ZN(n1123) );
NOR2_X1 U857 ( .A1(n1008), .A2(G952), .ZN(n1107) );
XNOR2_X1 U858 ( .A(G146), .B(n1174), .ZN(G48) );
NAND4_X1 U859 ( .A1(n1189), .A2(n1188), .A3(n1022), .A4(n1190), .ZN(n1174) );
XNOR2_X1 U860 ( .A(G143), .B(n1173), .ZN(G45) );
NAND4_X1 U861 ( .A1(n1172), .A2(n1170), .A3(n1022), .A4(n1053), .ZN(n1173) );
XOR2_X1 U862 ( .A(n1191), .B(n1192), .Z(G42) );
XOR2_X1 U863 ( .A(KEYINPUT25), .B(G140), .Z(n1192) );
NOR2_X1 U864 ( .A1(n1175), .A2(KEYINPUT50), .ZN(n1191) );
NOR4_X1 U865 ( .A1(n1042), .A2(n1193), .A3(n1034), .A4(n1194), .ZN(n1175) );
NAND2_X1 U866 ( .A1(n1188), .A2(n1023), .ZN(n1194) );
XOR2_X1 U867 ( .A(n1154), .B(n1195), .Z(G39) );
XNOR2_X1 U868 ( .A(G137), .B(KEYINPUT45), .ZN(n1195) );
NAND4_X1 U869 ( .A1(n1189), .A2(n1023), .A3(n1014), .A4(n1190), .ZN(n1154) );
XNOR2_X1 U870 ( .A(G134), .B(n1196), .ZN(G36) );
NAND2_X1 U871 ( .A1(n1023), .A2(n1166), .ZN(n1196) );
AND2_X1 U872 ( .A1(n1170), .A2(n1032), .ZN(n1166) );
XOR2_X1 U873 ( .A(G131), .B(n1160), .Z(G33) );
AND3_X1 U874 ( .A1(n1170), .A2(n1188), .A3(n1023), .ZN(n1160) );
INV_X1 U875 ( .A(n1165), .ZN(n1023) );
NAND2_X1 U876 ( .A1(n1021), .A2(n1197), .ZN(n1165) );
NOR3_X1 U877 ( .A1(n1042), .A2(n1193), .A3(n1035), .ZN(n1170) );
INV_X1 U878 ( .A(n1190), .ZN(n1042) );
XOR2_X1 U879 ( .A(n1198), .B(KEYINPUT10), .Z(n1190) );
XOR2_X1 U880 ( .A(G128), .B(n1159), .Z(G30) );
AND4_X1 U881 ( .A1(n1189), .A2(n1032), .A3(n1022), .A4(n1198), .ZN(n1159) );
AND3_X1 U882 ( .A1(n1069), .A2(n1163), .A3(n1199), .ZN(n1189) );
XNOR2_X1 U883 ( .A(n1200), .B(n1201), .ZN(G3) );
NOR2_X1 U884 ( .A1(n1186), .A2(n1035), .ZN(n1201) );
XNOR2_X1 U885 ( .A(n1202), .B(n1203), .ZN(G27) );
NOR4_X1 U886 ( .A1(KEYINPUT7), .A2(n1193), .A3(n1034), .A4(n1162), .ZN(n1203) );
NAND3_X1 U887 ( .A1(n1015), .A2(n1022), .A3(n1188), .ZN(n1162) );
INV_X1 U888 ( .A(n1163), .ZN(n1193) );
NAND2_X1 U889 ( .A1(n1046), .A2(n1204), .ZN(n1163) );
NAND4_X1 U890 ( .A1(G902), .A2(G953), .A3(n1205), .A4(n1080), .ZN(n1204) );
INV_X1 U891 ( .A(G900), .ZN(n1080) );
XNOR2_X1 U892 ( .A(G122), .B(n1178), .ZN(G24) );
NAND4_X1 U893 ( .A1(n1172), .A2(n1206), .A3(n1016), .A4(n1053), .ZN(n1178) );
AND2_X1 U894 ( .A1(n1207), .A2(n1208), .ZN(n1016) );
XNOR2_X1 U895 ( .A(G119), .B(n1183), .ZN(G21) );
NAND4_X1 U896 ( .A1(n1199), .A2(n1014), .A3(n1206), .A4(n1069), .ZN(n1183) );
XNOR2_X1 U897 ( .A(G116), .B(n1182), .ZN(G18) );
NAND3_X1 U898 ( .A1(n1206), .A2(n1032), .A3(n1187), .ZN(n1182) );
NOR2_X1 U899 ( .A1(n1209), .A2(n1172), .ZN(n1032) );
XOR2_X1 U900 ( .A(n1180), .B(n1210), .Z(G15) );
NOR2_X1 U901 ( .A1(G113), .A2(KEYINPUT27), .ZN(n1210) );
NAND3_X1 U902 ( .A1(n1187), .A2(n1206), .A3(n1188), .ZN(n1180) );
INV_X1 U903 ( .A(n1039), .ZN(n1188) );
NAND2_X1 U904 ( .A1(n1172), .A2(n1209), .ZN(n1039) );
INV_X1 U905 ( .A(n1053), .ZN(n1209) );
AND3_X1 U906 ( .A1(n1022), .A2(n1211), .A3(n1015), .ZN(n1206) );
NOR2_X1 U907 ( .A1(n1212), .A2(n1044), .ZN(n1015) );
INV_X1 U908 ( .A(n1035), .ZN(n1187) );
NAND2_X1 U909 ( .A1(n1199), .A2(n1207), .ZN(n1035) );
XNOR2_X1 U910 ( .A(n1069), .B(KEYINPUT11), .ZN(n1207) );
INV_X1 U911 ( .A(n1208), .ZN(n1199) );
XNOR2_X1 U912 ( .A(G110), .B(n1179), .ZN(G12) );
OR2_X1 U913 ( .A1(n1034), .A2(n1186), .ZN(n1179) );
NAND2_X1 U914 ( .A1(n1014), .A2(n1181), .ZN(n1186) );
AND3_X1 U915 ( .A1(n1198), .A2(n1211), .A3(n1022), .ZN(n1181) );
NOR2_X1 U916 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
INV_X1 U917 ( .A(n1197), .ZN(n1020) );
NAND2_X1 U918 ( .A1(G214), .A2(n1213), .ZN(n1197) );
XNOR2_X1 U919 ( .A(n1072), .B(n1214), .ZN(n1021) );
NOR2_X1 U920 ( .A1(n1071), .A2(KEYINPUT12), .ZN(n1214) );
AND2_X1 U921 ( .A1(G210), .A2(n1213), .ZN(n1071) );
NAND2_X1 U922 ( .A1(n1215), .A2(n1216), .ZN(n1213) );
INV_X1 U923 ( .A(G237), .ZN(n1216) );
NAND2_X1 U924 ( .A1(n1217), .A2(n1218), .ZN(n1072) );
XOR2_X1 U925 ( .A(n1219), .B(n1149), .Z(n1217) );
XNOR2_X1 U926 ( .A(n1102), .B(n1220), .ZN(n1149) );
XOR2_X1 U927 ( .A(n1221), .B(n1222), .Z(n1220) );
NOR2_X1 U928 ( .A1(KEYINPUT33), .A2(n1106), .ZN(n1222) );
NOR2_X1 U929 ( .A1(G953), .A2(n1097), .ZN(n1221) );
INV_X1 U930 ( .A(G224), .ZN(n1097) );
XOR2_X1 U931 ( .A(n1223), .B(n1224), .Z(n1102) );
XNOR2_X1 U932 ( .A(n1225), .B(n1226), .ZN(n1224) );
XOR2_X1 U933 ( .A(KEYINPUT16), .B(G122), .Z(n1226) );
XOR2_X1 U934 ( .A(n1227), .B(n1228), .Z(n1223) );
XNOR2_X1 U935 ( .A(G101), .B(n1229), .ZN(n1228) );
NAND2_X1 U936 ( .A1(n1230), .A2(KEYINPUT53), .ZN(n1229) );
XNOR2_X1 U937 ( .A(G110), .B(KEYINPUT57), .ZN(n1230) );
NAND2_X1 U938 ( .A1(KEYINPUT51), .A2(G107), .ZN(n1227) );
NAND2_X1 U939 ( .A1(KEYINPUT5), .A2(n1150), .ZN(n1219) );
XNOR2_X1 U940 ( .A(G125), .B(n1138), .ZN(n1150) );
NAND2_X1 U941 ( .A1(n1046), .A2(n1231), .ZN(n1211) );
NAND3_X1 U942 ( .A1(n1095), .A2(n1205), .A3(G902), .ZN(n1231) );
NOR2_X1 U943 ( .A1(G898), .A2(n1008), .ZN(n1095) );
NAND3_X1 U944 ( .A1(n1205), .A2(n1008), .A3(G952), .ZN(n1046) );
NAND2_X1 U945 ( .A1(G237), .A2(G234), .ZN(n1205) );
NOR2_X1 U946 ( .A1(n1045), .A2(n1044), .ZN(n1198) );
AND2_X1 U947 ( .A1(G221), .A2(n1113), .ZN(n1044) );
INV_X1 U948 ( .A(n1212), .ZN(n1045) );
XNOR2_X1 U949 ( .A(n1054), .B(G469), .ZN(n1212) );
NAND2_X1 U950 ( .A1(n1232), .A2(n1218), .ZN(n1054) );
XOR2_X1 U951 ( .A(n1233), .B(n1144), .Z(n1232) );
XNOR2_X1 U952 ( .A(n1234), .B(n1235), .ZN(n1144) );
XOR2_X1 U953 ( .A(n1236), .B(n1139), .Z(n1235) );
NOR2_X1 U954 ( .A1(G953), .A2(n1088), .ZN(n1236) );
INV_X1 U955 ( .A(G227), .ZN(n1088) );
NAND2_X1 U956 ( .A1(KEYINPUT41), .A2(n1142), .ZN(n1233) );
XOR2_X1 U957 ( .A(n1237), .B(n1238), .Z(n1142) );
XNOR2_X1 U958 ( .A(n1239), .B(G104), .ZN(n1238) );
XNOR2_X1 U959 ( .A(n1085), .B(n1200), .ZN(n1237) );
INV_X1 U960 ( .A(G101), .ZN(n1200) );
XOR2_X1 U961 ( .A(n1240), .B(n1241), .Z(n1085) );
XOR2_X1 U962 ( .A(n1242), .B(n1243), .Z(n1241) );
NOR2_X1 U963 ( .A1(G146), .A2(KEYINPUT37), .ZN(n1242) );
XNOR2_X1 U964 ( .A(G143), .B(KEYINPUT20), .ZN(n1240) );
NOR2_X1 U965 ( .A1(n1053), .A2(n1172), .ZN(n1014) );
XOR2_X1 U966 ( .A(n1244), .B(n1067), .Z(n1172) );
NOR2_X1 U967 ( .A1(n1120), .A2(G902), .ZN(n1067) );
XOR2_X1 U968 ( .A(n1245), .B(n1246), .Z(n1120) );
XOR2_X1 U969 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U970 ( .A(G113), .B(n1249), .Z(n1248) );
NOR2_X1 U971 ( .A1(KEYINPUT46), .A2(n1250), .ZN(n1249) );
XOR2_X1 U972 ( .A(G131), .B(G122), .Z(n1247) );
XOR2_X1 U973 ( .A(n1251), .B(n1252), .Z(n1245) );
XOR2_X1 U974 ( .A(n1253), .B(n1254), .Z(n1252) );
NAND2_X1 U975 ( .A1(n1255), .A2(G214), .ZN(n1254) );
NAND3_X1 U976 ( .A1(n1256), .A2(n1257), .A3(KEYINPUT44), .ZN(n1253) );
NAND2_X1 U977 ( .A1(n1086), .A2(n1258), .ZN(n1257) );
NAND2_X1 U978 ( .A1(KEYINPUT8), .A2(n1259), .ZN(n1258) );
NAND2_X1 U979 ( .A1(G146), .A2(n1260), .ZN(n1259) );
NAND2_X1 U980 ( .A1(n1261), .A2(n1262), .ZN(n1256) );
NAND2_X1 U981 ( .A1(n1260), .A2(n1263), .ZN(n1261) );
NAND2_X1 U982 ( .A1(KEYINPUT8), .A2(n1264), .ZN(n1263) );
INV_X1 U983 ( .A(n1086), .ZN(n1264) );
XOR2_X1 U984 ( .A(G140), .B(n1202), .Z(n1086) );
INV_X1 U985 ( .A(KEYINPUT28), .ZN(n1260) );
NAND2_X1 U986 ( .A1(KEYINPUT22), .A2(n1225), .ZN(n1251) );
INV_X1 U987 ( .A(G104), .ZN(n1225) );
NAND2_X1 U988 ( .A1(KEYINPUT13), .A2(n1059), .ZN(n1244) );
INV_X1 U989 ( .A(G475), .ZN(n1059) );
XNOR2_X1 U990 ( .A(n1265), .B(G478), .ZN(n1053) );
NAND2_X1 U991 ( .A1(n1116), .A2(n1218), .ZN(n1265) );
XNOR2_X1 U992 ( .A(n1266), .B(n1267), .ZN(n1116) );
AND2_X1 U993 ( .A1(n1268), .A2(G217), .ZN(n1267) );
NAND2_X1 U994 ( .A1(KEYINPUT52), .A2(n1269), .ZN(n1266) );
XOR2_X1 U995 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U996 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U997 ( .A(G122), .B(G116), .Z(n1273) );
NAND2_X1 U998 ( .A1(KEYINPUT55), .A2(n1239), .ZN(n1272) );
INV_X1 U999 ( .A(G107), .ZN(n1239) );
XOR2_X1 U1000 ( .A(n1274), .B(n1275), .Z(n1270) );
XNOR2_X1 U1001 ( .A(KEYINPUT23), .B(n1250), .ZN(n1275) );
INV_X1 U1002 ( .A(G143), .ZN(n1250) );
XNOR2_X1 U1003 ( .A(G134), .B(G128), .ZN(n1274) );
NAND2_X1 U1004 ( .A1(n1069), .A2(n1208), .ZN(n1034) );
NAND3_X1 U1005 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1208) );
NAND2_X1 U1006 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
OR3_X1 U1007 ( .A1(n1280), .A2(n1279), .A3(KEYINPUT21), .ZN(n1277) );
INV_X1 U1008 ( .A(n1068), .ZN(n1279) );
NAND2_X1 U1009 ( .A1(n1281), .A2(n1218), .ZN(n1068) );
XOR2_X1 U1010 ( .A(n1282), .B(n1283), .Z(n1281) );
XOR2_X1 U1011 ( .A(n1132), .B(n1284), .Z(n1283) );
XNOR2_X1 U1012 ( .A(G101), .B(KEYINPUT32), .ZN(n1284) );
NAND2_X1 U1013 ( .A1(n1255), .A2(G210), .ZN(n1132) );
NOR2_X1 U1014 ( .A1(G953), .A2(G237), .ZN(n1255) );
XOR2_X1 U1015 ( .A(n1285), .B(n1139), .Z(n1282) );
XNOR2_X1 U1016 ( .A(n1286), .B(n1083), .ZN(n1139) );
XOR2_X1 U1017 ( .A(G131), .B(n1287), .Z(n1083) );
XNOR2_X1 U1018 ( .A(KEYINPUT39), .B(n1288), .ZN(n1286) );
NOR2_X1 U1019 ( .A1(KEYINPUT58), .A2(n1084), .ZN(n1288) );
XNOR2_X1 U1020 ( .A(n1289), .B(KEYINPUT48), .ZN(n1084) );
INV_X1 U1021 ( .A(G134), .ZN(n1289) );
XNOR2_X1 U1022 ( .A(n1138), .B(n1106), .ZN(n1285) );
XNOR2_X1 U1023 ( .A(n1290), .B(n1291), .ZN(n1106) );
XOR2_X1 U1024 ( .A(KEYINPUT43), .B(G119), .Z(n1291) );
XNOR2_X1 U1025 ( .A(G113), .B(G116), .ZN(n1290) );
XNOR2_X1 U1026 ( .A(n1292), .B(n1243), .ZN(n1138) );
XOR2_X1 U1027 ( .A(G128), .B(KEYINPUT6), .Z(n1243) );
NAND2_X1 U1028 ( .A1(KEYINPUT35), .A2(n1293), .ZN(n1292) );
XOR2_X1 U1029 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U1030 ( .A(G143), .B(KEYINPUT42), .ZN(n1295) );
NAND2_X1 U1031 ( .A1(KEYINPUT31), .A2(n1262), .ZN(n1294) );
NAND2_X1 U1032 ( .A1(n1296), .A2(n1297), .ZN(n1280) );
INV_X1 U1033 ( .A(G472), .ZN(n1297) );
XOR2_X1 U1034 ( .A(KEYINPUT63), .B(KEYINPUT61), .Z(n1296) );
NAND2_X1 U1035 ( .A1(KEYINPUT21), .A2(G472), .ZN(n1276) );
XNOR2_X1 U1036 ( .A(n1298), .B(n1299), .ZN(n1069) );
AND2_X1 U1037 ( .A1(n1113), .A2(G217), .ZN(n1299) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1215), .ZN(n1113) );
XNOR2_X1 U1039 ( .A(n1218), .B(KEYINPUT54), .ZN(n1215) );
NAND2_X1 U1040 ( .A1(n1110), .A2(n1218), .ZN(n1298) );
INV_X1 U1041 ( .A(G902), .ZN(n1218) );
XNOR2_X1 U1042 ( .A(n1300), .B(n1301), .ZN(n1110) );
XOR2_X1 U1043 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U1044 ( .A(n1202), .B(G119), .ZN(n1303) );
INV_X1 U1045 ( .A(G125), .ZN(n1202) );
XNOR2_X1 U1046 ( .A(n1262), .B(G128), .ZN(n1302) );
INV_X1 U1047 ( .A(G146), .ZN(n1262) );
XNOR2_X1 U1048 ( .A(n1304), .B(n1234), .ZN(n1300) );
XNOR2_X1 U1049 ( .A(G110), .B(G140), .ZN(n1234) );
XOR2_X1 U1050 ( .A(n1305), .B(n1287), .Z(n1304) );
XOR2_X1 U1051 ( .A(G137), .B(KEYINPUT38), .Z(n1287) );
NAND2_X1 U1052 ( .A1(n1268), .A2(G221), .ZN(n1305) );
AND2_X1 U1053 ( .A1(G234), .A2(n1008), .ZN(n1268) );
INV_X1 U1054 ( .A(G953), .ZN(n1008) );
endmodule


