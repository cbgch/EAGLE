//Key = 0110001111011100010101010001011001010110011011100001100101001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359;

XNOR2_X1 U736 ( .A(n1030), .B(n1031), .ZN(G9) );
NOR3_X1 U737 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NOR2_X1 U738 ( .A1(n1035), .A2(n1036), .ZN(G75) );
NOR4_X1 U739 ( .A1(n1037), .A2(n1038), .A3(G953), .A4(n1039), .ZN(n1036) );
NOR4_X1 U740 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1038) );
NOR2_X1 U741 ( .A1(n1044), .A2(n1045), .ZN(n1040) );
NOR2_X1 U742 ( .A1(n1046), .A2(n1032), .ZN(n1045) );
NOR2_X1 U743 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U744 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U745 ( .A1(n1051), .A2(n1052), .ZN(n1044) );
NOR2_X1 U746 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NAND2_X1 U747 ( .A1(n1055), .A2(n1056), .ZN(n1037) );
NAND4_X1 U748 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
NAND2_X1 U749 ( .A1(n1061), .A2(n1043), .ZN(n1060) );
OR3_X1 U750 ( .A1(n1033), .A2(KEYINPUT9), .A3(n1042), .ZN(n1061) );
NAND2_X1 U751 ( .A1(n1062), .A2(n1063), .ZN(n1059) );
INV_X1 U752 ( .A(n1043), .ZN(n1063) );
NAND2_X1 U753 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND2_X1 U754 ( .A1(n1066), .A2(n1042), .ZN(n1065) );
INV_X1 U755 ( .A(n1067), .ZN(n1042) );
NAND2_X1 U756 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NAND2_X1 U757 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND3_X1 U758 ( .A1(n1072), .A2(n1073), .A3(n1067), .ZN(n1064) );
NAND2_X1 U759 ( .A1(KEYINPUT9), .A2(n1074), .ZN(n1072) );
NOR3_X1 U760 ( .A1(n1039), .A2(G953), .A3(G952), .ZN(n1035) );
AND4_X1 U761 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1039) );
NOR4_X1 U762 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1082), .ZN(n1078) );
NOR2_X1 U763 ( .A1(KEYINPUT17), .A2(n1083), .ZN(n1082) );
XOR2_X1 U764 ( .A(n1049), .B(KEYINPUT34), .Z(n1081) );
NAND3_X1 U765 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1079) );
XOR2_X1 U766 ( .A(n1087), .B(G478), .Z(n1086) );
NAND3_X1 U767 ( .A1(KEYINPUT17), .A2(n1083), .A3(n1088), .ZN(n1085) );
NAND2_X1 U768 ( .A1(G469), .A2(n1089), .ZN(n1084) );
NAND2_X1 U769 ( .A1(KEYINPUT17), .A2(n1090), .ZN(n1089) );
XNOR2_X1 U770 ( .A(KEYINPUT20), .B(n1091), .ZN(n1090) );
NOR3_X1 U771 ( .A1(n1092), .A2(n1093), .A3(n1070), .ZN(n1077) );
XNOR2_X1 U772 ( .A(KEYINPUT21), .B(n1094), .ZN(n1075) );
XOR2_X1 U773 ( .A(n1095), .B(n1096), .Z(G72) );
XOR2_X1 U774 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U775 ( .A1(G953), .A2(n1099), .ZN(n1098) );
XOR2_X1 U776 ( .A(n1100), .B(KEYINPUT55), .Z(n1099) );
NAND2_X1 U777 ( .A1(n1101), .A2(n1102), .ZN(n1097) );
XOR2_X1 U778 ( .A(n1103), .B(n1104), .Z(n1101) );
XNOR2_X1 U779 ( .A(n1105), .B(n1106), .ZN(n1104) );
NOR3_X1 U780 ( .A1(KEYINPUT15), .A2(n1107), .A3(n1108), .ZN(n1106) );
NOR3_X1 U781 ( .A1(G131), .A2(n1109), .A3(n1110), .ZN(n1108) );
NOR2_X1 U782 ( .A1(n1111), .A2(n1112), .ZN(n1107) );
NOR2_X1 U783 ( .A1(n1109), .A2(n1110), .ZN(n1111) );
NAND2_X1 U784 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
OR2_X1 U785 ( .A1(n1115), .A2(KEYINPUT11), .ZN(n1114) );
NAND3_X1 U786 ( .A1(G134), .A2(n1115), .A3(KEYINPUT11), .ZN(n1113) );
NAND2_X1 U787 ( .A1(n1116), .A2(n1117), .ZN(n1095) );
NAND2_X1 U788 ( .A1(G900), .A2(G227), .ZN(n1117) );
XOR2_X1 U789 ( .A(n1118), .B(n1119), .Z(G69) );
XOR2_X1 U790 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U791 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U792 ( .A1(G898), .A2(n1124), .ZN(n1122) );
NAND2_X1 U793 ( .A1(n1125), .A2(n1126), .ZN(n1120) );
NAND2_X1 U794 ( .A1(n1116), .A2(n1127), .ZN(n1118) );
NAND2_X1 U795 ( .A1(G898), .A2(G224), .ZN(n1127) );
XNOR2_X1 U796 ( .A(G953), .B(KEYINPUT6), .ZN(n1116) );
NOR2_X1 U797 ( .A1(n1128), .A2(n1129), .ZN(G66) );
XOR2_X1 U798 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U799 ( .A1(n1132), .A2(n1133), .ZN(n1130) );
NOR2_X1 U800 ( .A1(n1128), .A2(n1134), .ZN(G63) );
XOR2_X1 U801 ( .A(n1135), .B(n1136), .Z(n1134) );
AND2_X1 U802 ( .A1(G478), .A2(n1132), .ZN(n1136) );
NAND2_X1 U803 ( .A1(KEYINPUT29), .A2(n1137), .ZN(n1135) );
NOR2_X1 U804 ( .A1(n1128), .A2(n1138), .ZN(G60) );
XOR2_X1 U805 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U806 ( .A1(n1132), .A2(G475), .ZN(n1139) );
XOR2_X1 U807 ( .A(n1141), .B(n1142), .Z(G6) );
NOR2_X1 U808 ( .A1(KEYINPUT18), .A2(n1143), .ZN(n1142) );
NOR2_X1 U809 ( .A1(n1128), .A2(n1144), .ZN(G57) );
XOR2_X1 U810 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U811 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U812 ( .A(n1149), .B(n1150), .Z(n1145) );
NAND2_X1 U813 ( .A1(n1132), .A2(G472), .ZN(n1149) );
NOR2_X1 U814 ( .A1(n1128), .A2(n1151), .ZN(G54) );
XOR2_X1 U815 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U816 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND3_X1 U817 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1154) );
INV_X1 U818 ( .A(n1159), .ZN(n1158) );
OR2_X1 U819 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NAND3_X1 U820 ( .A1(n1162), .A2(n1160), .A3(n1161), .ZN(n1156) );
NAND2_X1 U821 ( .A1(G140), .A2(n1163), .ZN(n1160) );
XOR2_X1 U822 ( .A(KEYINPUT8), .B(G110), .Z(n1163) );
XOR2_X1 U823 ( .A(n1164), .B(KEYINPUT57), .Z(n1152) );
NAND2_X1 U824 ( .A1(n1132), .A2(G469), .ZN(n1164) );
NOR2_X1 U825 ( .A1(n1128), .A2(n1165), .ZN(G51) );
XOR2_X1 U826 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U827 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U828 ( .A1(KEYINPUT14), .A2(n1170), .ZN(n1168) );
XOR2_X1 U829 ( .A(n1171), .B(KEYINPUT50), .Z(n1166) );
NAND2_X1 U830 ( .A1(n1132), .A2(G210), .ZN(n1171) );
NOR2_X1 U831 ( .A1(n1172), .A2(n1055), .ZN(n1132) );
NOR2_X1 U832 ( .A1(n1100), .A2(n1126), .ZN(n1055) );
NAND4_X1 U833 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1126) );
NOR4_X1 U834 ( .A1(n1177), .A2(n1141), .A3(n1178), .A4(n1179), .ZN(n1176) );
NOR3_X1 U835 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1179) );
XNOR2_X1 U836 ( .A(n1048), .B(KEYINPUT5), .ZN(n1182) );
XOR2_X1 U837 ( .A(n1183), .B(KEYINPUT12), .Z(n1181) );
NOR3_X1 U838 ( .A1(n1032), .A2(n1034), .A3(n1073), .ZN(n1141) );
OR2_X1 U839 ( .A1(n1184), .A2(n1185), .ZN(n1175) );
NAND3_X1 U840 ( .A1(n1074), .A2(n1186), .A3(n1187), .ZN(n1174) );
XNOR2_X1 U841 ( .A(KEYINPUT62), .B(n1032), .ZN(n1186) );
INV_X1 U842 ( .A(n1058), .ZN(n1032) );
NAND2_X1 U843 ( .A1(n1188), .A2(n1189), .ZN(n1173) );
NAND2_X1 U844 ( .A1(n1073), .A2(n1033), .ZN(n1189) );
INV_X1 U845 ( .A(n1190), .ZN(n1188) );
NAND4_X1 U846 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1100) );
NOR4_X1 U847 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1194) );
NAND3_X1 U848 ( .A1(n1199), .A2(n1200), .A3(n1054), .ZN(n1193) );
NAND2_X1 U849 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NAND3_X1 U850 ( .A1(n1203), .A2(n1204), .A3(n1067), .ZN(n1202) );
XNOR2_X1 U851 ( .A(KEYINPUT0), .B(n1185), .ZN(n1203) );
NAND3_X1 U852 ( .A1(n1205), .A2(n1074), .A3(n1206), .ZN(n1191) );
XNOR2_X1 U853 ( .A(n1207), .B(KEYINPUT44), .ZN(n1206) );
NOR2_X1 U854 ( .A1(n1125), .A2(G952), .ZN(n1128) );
NAND2_X1 U855 ( .A1(n1208), .A2(n1209), .ZN(G48) );
NAND2_X1 U856 ( .A1(G146), .A2(n1192), .ZN(n1209) );
XOR2_X1 U857 ( .A(KEYINPUT7), .B(n1210), .Z(n1208) );
NOR2_X1 U858 ( .A1(G146), .A2(n1192), .ZN(n1210) );
NAND3_X1 U859 ( .A1(n1207), .A2(n1199), .A3(n1205), .ZN(n1192) );
XNOR2_X1 U860 ( .A(n1211), .B(n1198), .ZN(G45) );
AND3_X1 U861 ( .A1(n1053), .A2(n1212), .A3(n1205), .ZN(n1198) );
XNOR2_X1 U862 ( .A(n1213), .B(n1214), .ZN(G42) );
NOR4_X1 U863 ( .A1(KEYINPUT22), .A2(n1201), .A3(n1073), .A4(n1215), .ZN(n1214) );
XNOR2_X1 U864 ( .A(n1197), .B(n1216), .ZN(G39) );
NAND2_X1 U865 ( .A1(KEYINPUT2), .A2(G137), .ZN(n1216) );
NOR3_X1 U866 ( .A1(n1217), .A2(n1201), .A3(n1041), .ZN(n1197) );
INV_X1 U867 ( .A(n1218), .ZN(n1201) );
XNOR2_X1 U868 ( .A(n1219), .B(n1196), .ZN(G36) );
AND3_X1 U869 ( .A1(n1218), .A2(n1074), .A3(n1053), .ZN(n1196) );
XNOR2_X1 U870 ( .A(n1112), .B(n1195), .ZN(G33) );
AND3_X1 U871 ( .A1(n1053), .A2(n1218), .A3(n1199), .ZN(n1195) );
NOR4_X1 U872 ( .A1(n1220), .A2(n1052), .A3(n1221), .A4(n1070), .ZN(n1218) );
INV_X1 U873 ( .A(n1057), .ZN(n1052) );
NOR2_X1 U874 ( .A1(n1049), .A2(n1222), .ZN(n1057) );
XNOR2_X1 U875 ( .A(KEYINPUT30), .B(n1092), .ZN(n1222) );
INV_X1 U876 ( .A(n1050), .ZN(n1092) );
XNOR2_X1 U877 ( .A(n1223), .B(n1224), .ZN(G30) );
AND3_X1 U878 ( .A1(n1205), .A2(n1074), .A3(n1207), .ZN(n1224) );
NOR4_X1 U879 ( .A1(n1220), .A2(n1185), .A3(n1221), .A4(n1070), .ZN(n1205) );
NAND2_X1 U880 ( .A1(n1225), .A2(n1226), .ZN(G3) );
NAND2_X1 U881 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
XNOR2_X1 U882 ( .A(KEYINPUT59), .B(n1229), .ZN(n1227) );
NAND2_X1 U883 ( .A1(G101), .A2(n1230), .ZN(n1225) );
XNOR2_X1 U884 ( .A(n1178), .B(KEYINPUT43), .ZN(n1230) );
INV_X1 U885 ( .A(n1229), .ZN(n1178) );
NAND3_X1 U886 ( .A1(n1053), .A2(n1187), .A3(n1068), .ZN(n1229) );
INV_X1 U887 ( .A(n1034), .ZN(n1187) );
XNOR2_X1 U888 ( .A(G125), .B(n1231), .ZN(G27) );
NAND3_X1 U889 ( .A1(n1054), .A2(n1067), .A3(n1232), .ZN(n1231) );
NOR3_X1 U890 ( .A1(n1185), .A2(n1221), .A3(n1233), .ZN(n1232) );
XNOR2_X1 U891 ( .A(n1199), .B(KEYINPUT26), .ZN(n1233) );
INV_X1 U892 ( .A(n1204), .ZN(n1221) );
NAND2_X1 U893 ( .A1(n1234), .A2(n1043), .ZN(n1204) );
XOR2_X1 U894 ( .A(KEYINPUT61), .B(n1235), .Z(n1234) );
NOR3_X1 U895 ( .A1(n1102), .A2(n1236), .A3(n1172), .ZN(n1235) );
OR2_X1 U896 ( .A1(n1124), .A2(G900), .ZN(n1102) );
INV_X1 U897 ( .A(n1215), .ZN(n1054) );
NAND2_X1 U898 ( .A1(n1237), .A2(n1238), .ZN(G24) );
NAND2_X1 U899 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
XOR2_X1 U900 ( .A(n1241), .B(KEYINPUT36), .Z(n1237) );
OR2_X1 U901 ( .A1(n1240), .A2(n1239), .ZN(n1241) );
NOR3_X1 U902 ( .A1(n1185), .A2(n1242), .A3(n1180), .ZN(n1239) );
NAND3_X1 U903 ( .A1(n1058), .A2(n1212), .A3(n1067), .ZN(n1180) );
NAND2_X1 U904 ( .A1(n1243), .A2(n1244), .ZN(n1212) );
OR3_X1 U905 ( .A1(n1245), .A2(n1246), .A3(KEYINPUT24), .ZN(n1244) );
NAND2_X1 U906 ( .A1(KEYINPUT24), .A2(n1199), .ZN(n1243) );
NOR2_X1 U907 ( .A1(n1247), .A2(n1248), .ZN(n1058) );
INV_X1 U908 ( .A(n1183), .ZN(n1242) );
INV_X1 U909 ( .A(G122), .ZN(n1240) );
XNOR2_X1 U910 ( .A(G119), .B(n1249), .ZN(G21) );
NAND2_X1 U911 ( .A1(n1250), .A2(n1048), .ZN(n1249) );
XOR2_X1 U912 ( .A(n1184), .B(KEYINPUT35), .Z(n1250) );
NAND4_X1 U913 ( .A1(n1067), .A2(n1068), .A3(n1207), .A4(n1183), .ZN(n1184) );
INV_X1 U914 ( .A(n1217), .ZN(n1207) );
NAND2_X1 U915 ( .A1(n1248), .A2(n1247), .ZN(n1217) );
XOR2_X1 U916 ( .A(n1251), .B(n1252), .Z(G18) );
NOR2_X1 U917 ( .A1(n1253), .A2(n1190), .ZN(n1252) );
XNOR2_X1 U918 ( .A(n1074), .B(KEYINPUT54), .ZN(n1253) );
INV_X1 U919 ( .A(n1033), .ZN(n1074) );
NAND2_X1 U920 ( .A1(n1246), .A2(n1254), .ZN(n1033) );
XNOR2_X1 U921 ( .A(KEYINPUT24), .B(n1245), .ZN(n1254) );
INV_X1 U922 ( .A(n1255), .ZN(n1245) );
NAND2_X1 U923 ( .A1(KEYINPUT23), .A2(n1256), .ZN(n1251) );
INV_X1 U924 ( .A(G116), .ZN(n1256) );
XOR2_X1 U925 ( .A(G113), .B(n1257), .Z(G15) );
NOR3_X1 U926 ( .A1(n1258), .A2(n1073), .A3(n1190), .ZN(n1257) );
NAND4_X1 U927 ( .A1(n1067), .A2(n1053), .A3(n1048), .A4(n1183), .ZN(n1190) );
NOR2_X1 U928 ( .A1(n1247), .A2(n1094), .ZN(n1053) );
NOR2_X1 U929 ( .A1(n1071), .A2(n1070), .ZN(n1067) );
INV_X1 U930 ( .A(n1259), .ZN(n1070) );
INV_X1 U931 ( .A(n1199), .ZN(n1073) );
NOR2_X1 U932 ( .A1(n1255), .A2(n1246), .ZN(n1199) );
INV_X1 U933 ( .A(n1080), .ZN(n1246) );
XOR2_X1 U934 ( .A(KEYINPUT28), .B(KEYINPUT16), .Z(n1258) );
XOR2_X1 U935 ( .A(G110), .B(n1177), .Z(G12) );
NOR3_X1 U936 ( .A1(n1041), .A2(n1034), .A3(n1215), .ZN(n1177) );
NAND2_X1 U937 ( .A1(n1094), .A2(n1247), .ZN(n1215) );
NAND2_X1 U938 ( .A1(n1260), .A2(n1076), .ZN(n1247) );
NAND2_X1 U939 ( .A1(n1133), .A2(n1261), .ZN(n1076) );
XOR2_X1 U940 ( .A(KEYINPUT63), .B(n1093), .Z(n1260) );
NOR2_X1 U941 ( .A1(n1261), .A2(n1133), .ZN(n1093) );
AND2_X1 U942 ( .A1(G217), .A2(n1262), .ZN(n1133) );
NAND2_X1 U943 ( .A1(n1131), .A2(n1172), .ZN(n1261) );
XNOR2_X1 U944 ( .A(n1263), .B(n1264), .ZN(n1131) );
XOR2_X1 U945 ( .A(G110), .B(n1265), .Z(n1264) );
XNOR2_X1 U946 ( .A(n1223), .B(G119), .ZN(n1265) );
XOR2_X1 U947 ( .A(n1266), .B(n1267), .Z(n1263) );
XOR2_X1 U948 ( .A(n1268), .B(n1269), .Z(n1267) );
NAND3_X1 U949 ( .A1(G234), .A2(n1125), .A3(G221), .ZN(n1269) );
NAND2_X1 U950 ( .A1(KEYINPUT46), .A2(n1115), .ZN(n1268) );
NAND2_X1 U951 ( .A1(n1270), .A2(n1271), .ZN(n1266) );
NAND3_X1 U952 ( .A1(G146), .A2(n1272), .A3(n1273), .ZN(n1271) );
INV_X1 U953 ( .A(KEYINPUT45), .ZN(n1273) );
XNOR2_X1 U954 ( .A(n1213), .B(G125), .ZN(n1272) );
NAND2_X1 U955 ( .A1(n1105), .A2(KEYINPUT45), .ZN(n1270) );
INV_X1 U956 ( .A(n1248), .ZN(n1094) );
XNOR2_X1 U957 ( .A(n1274), .B(G472), .ZN(n1248) );
NAND2_X1 U958 ( .A1(n1275), .A2(n1172), .ZN(n1274) );
XNOR2_X1 U959 ( .A(n1276), .B(n1150), .ZN(n1275) );
XNOR2_X1 U960 ( .A(n1277), .B(n1278), .ZN(n1150) );
NAND2_X1 U961 ( .A1(G210), .A2(n1279), .ZN(n1277) );
NAND2_X1 U962 ( .A1(n1280), .A2(n1281), .ZN(n1276) );
OR2_X1 U963 ( .A1(n1148), .A2(n1147), .ZN(n1281) );
XOR2_X1 U964 ( .A(n1282), .B(KEYINPUT32), .Z(n1280) );
NAND2_X1 U965 ( .A1(n1147), .A2(n1148), .ZN(n1282) );
XNOR2_X1 U966 ( .A(n1283), .B(n1284), .ZN(n1148) );
XNOR2_X1 U967 ( .A(G113), .B(KEYINPUT40), .ZN(n1283) );
XNOR2_X1 U968 ( .A(n1285), .B(n1286), .ZN(n1147) );
XOR2_X1 U969 ( .A(n1287), .B(KEYINPUT52), .Z(n1285) );
NAND4_X1 U970 ( .A1(n1071), .A2(n1048), .A3(n1183), .A4(n1259), .ZN(n1034) );
NAND2_X1 U971 ( .A1(n1288), .A2(n1262), .ZN(n1259) );
NAND2_X1 U972 ( .A1(G234), .A2(n1172), .ZN(n1262) );
XOR2_X1 U973 ( .A(KEYINPUT58), .B(G221), .Z(n1288) );
NAND2_X1 U974 ( .A1(n1043), .A2(n1289), .ZN(n1183) );
OR4_X1 U975 ( .A1(n1124), .A2(n1172), .A3(n1236), .A4(G898), .ZN(n1289) );
INV_X1 U976 ( .A(n1290), .ZN(n1236) );
XOR2_X1 U977 ( .A(G953), .B(KEYINPUT37), .Z(n1124) );
NAND3_X1 U978 ( .A1(n1290), .A2(n1125), .A3(G952), .ZN(n1043) );
NAND2_X1 U979 ( .A1(G237), .A2(G234), .ZN(n1290) );
INV_X1 U980 ( .A(n1185), .ZN(n1048) );
NAND2_X1 U981 ( .A1(n1049), .A2(n1050), .ZN(n1185) );
NAND2_X1 U982 ( .A1(G214), .A2(n1291), .ZN(n1050) );
OR2_X1 U983 ( .A1(G237), .A2(G902), .ZN(n1291) );
NAND2_X1 U984 ( .A1(n1292), .A2(n1293), .ZN(n1049) );
NAND2_X1 U985 ( .A1(G210), .A2(n1294), .ZN(n1293) );
NAND2_X1 U986 ( .A1(n1172), .A2(n1295), .ZN(n1294) );
NAND2_X1 U987 ( .A1(G237), .A2(n1296), .ZN(n1295) );
NAND3_X1 U988 ( .A1(n1297), .A2(n1172), .A3(n1298), .ZN(n1292) );
INV_X1 U989 ( .A(n1296), .ZN(n1298) );
XOR2_X1 U990 ( .A(n1170), .B(n1169), .Z(n1296) );
XNOR2_X1 U991 ( .A(n1299), .B(n1286), .ZN(n1169) );
XNOR2_X1 U992 ( .A(n1300), .B(n1301), .ZN(n1286) );
NOR2_X1 U993 ( .A1(KEYINPUT31), .A2(G128), .ZN(n1301) );
XNOR2_X1 U994 ( .A(G143), .B(KEYINPUT38), .ZN(n1300) );
XOR2_X1 U995 ( .A(n1302), .B(n1303), .Z(n1299) );
NAND2_X1 U996 ( .A1(G224), .A2(n1125), .ZN(n1302) );
XNOR2_X1 U997 ( .A(n1123), .B(KEYINPUT39), .ZN(n1170) );
XOR2_X1 U998 ( .A(n1304), .B(n1305), .Z(n1123) );
XOR2_X1 U999 ( .A(G110), .B(n1306), .Z(n1305) );
XOR2_X1 U1000 ( .A(KEYINPUT4), .B(G113), .Z(n1306) );
XOR2_X1 U1001 ( .A(n1307), .B(n1308), .Z(n1304) );
XNOR2_X1 U1002 ( .A(n1309), .B(n1310), .ZN(n1308) );
NAND2_X1 U1003 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
OR2_X1 U1004 ( .A1(n1284), .A2(KEYINPUT56), .ZN(n1312) );
XOR2_X1 U1005 ( .A(G116), .B(G119), .Z(n1284) );
NAND3_X1 U1006 ( .A1(G116), .A2(n1313), .A3(KEYINPUT56), .ZN(n1311) );
INV_X1 U1007 ( .A(G119), .ZN(n1313) );
NAND2_X1 U1008 ( .A1(n1314), .A2(n1315), .ZN(n1307) );
NAND2_X1 U1009 ( .A1(n1316), .A2(G107), .ZN(n1315) );
NAND2_X1 U1010 ( .A1(n1317), .A2(n1030), .ZN(n1314) );
XNOR2_X1 U1011 ( .A(n1316), .B(KEYINPUT53), .ZN(n1317) );
NAND2_X1 U1012 ( .A1(G237), .A2(G210), .ZN(n1297) );
INV_X1 U1013 ( .A(n1220), .ZN(n1071) );
XOR2_X1 U1014 ( .A(n1083), .B(n1318), .Z(n1220) );
XNOR2_X1 U1015 ( .A(KEYINPUT41), .B(n1088), .ZN(n1318) );
INV_X1 U1016 ( .A(G469), .ZN(n1088) );
INV_X1 U1017 ( .A(n1091), .ZN(n1083) );
NAND2_X1 U1018 ( .A1(n1319), .A2(n1172), .ZN(n1091) );
XOR2_X1 U1019 ( .A(n1155), .B(n1320), .Z(n1319) );
XOR2_X1 U1020 ( .A(KEYINPUT25), .B(n1321), .Z(n1320) );
NOR3_X1 U1021 ( .A1(n1159), .A2(n1322), .A3(n1323), .ZN(n1321) );
NOR3_X1 U1022 ( .A1(G140), .A2(G110), .A3(n1324), .ZN(n1323) );
NOR2_X1 U1023 ( .A1(n1213), .A2(n1325), .ZN(n1322) );
XNOR2_X1 U1024 ( .A(G110), .B(n1324), .ZN(n1325) );
NOR2_X1 U1025 ( .A1(n1162), .A2(n1161), .ZN(n1159) );
INV_X1 U1026 ( .A(n1324), .ZN(n1161) );
NAND2_X1 U1027 ( .A1(G227), .A2(n1125), .ZN(n1324) );
NAND2_X1 U1028 ( .A1(G110), .A2(n1213), .ZN(n1162) );
INV_X1 U1029 ( .A(G140), .ZN(n1213) );
XOR2_X1 U1030 ( .A(n1326), .B(n1327), .Z(n1155) );
XNOR2_X1 U1031 ( .A(G107), .B(n1287), .ZN(n1327) );
XOR2_X1 U1032 ( .A(n1328), .B(n1329), .Z(n1287) );
NOR2_X1 U1033 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
XOR2_X1 U1034 ( .A(n1332), .B(KEYINPUT13), .Z(n1331) );
NAND2_X1 U1035 ( .A1(G131), .A2(n1333), .ZN(n1332) );
NAND2_X1 U1036 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
INV_X1 U1037 ( .A(n1109), .ZN(n1335) );
NAND2_X1 U1038 ( .A1(G134), .A2(n1115), .ZN(n1334) );
NOR3_X1 U1039 ( .A1(n1336), .A2(G131), .A3(n1109), .ZN(n1330) );
NOR2_X1 U1040 ( .A1(n1115), .A2(G134), .ZN(n1109) );
INV_X1 U1041 ( .A(G137), .ZN(n1115) );
NOR2_X1 U1042 ( .A1(G137), .A2(n1219), .ZN(n1336) );
INV_X1 U1043 ( .A(G134), .ZN(n1219) );
XNOR2_X1 U1044 ( .A(G146), .B(KEYINPUT51), .ZN(n1328) );
XNOR2_X1 U1045 ( .A(n1103), .B(n1337), .ZN(n1326) );
INV_X1 U1046 ( .A(n1316), .ZN(n1337) );
XOR2_X1 U1047 ( .A(G104), .B(n1278), .Z(n1316) );
XNOR2_X1 U1048 ( .A(n1228), .B(KEYINPUT47), .ZN(n1278) );
INV_X1 U1049 ( .A(G101), .ZN(n1228) );
XNOR2_X1 U1050 ( .A(n1338), .B(n1223), .ZN(n1103) );
INV_X1 U1051 ( .A(G128), .ZN(n1223) );
NAND2_X1 U1052 ( .A1(n1339), .A2(KEYINPUT42), .ZN(n1338) );
XNOR2_X1 U1053 ( .A(G143), .B(KEYINPUT10), .ZN(n1339) );
INV_X1 U1054 ( .A(n1068), .ZN(n1041) );
NOR2_X1 U1055 ( .A1(n1080), .A2(n1255), .ZN(n1068) );
XNOR2_X1 U1056 ( .A(n1340), .B(n1341), .ZN(n1255) );
NOR2_X1 U1057 ( .A1(G478), .A2(KEYINPUT49), .ZN(n1341) );
XOR2_X1 U1058 ( .A(n1087), .B(KEYINPUT60), .Z(n1340) );
NAND2_X1 U1059 ( .A1(n1137), .A2(n1172), .ZN(n1087) );
XNOR2_X1 U1060 ( .A(n1342), .B(n1343), .ZN(n1137) );
XOR2_X1 U1061 ( .A(n1344), .B(n1345), .Z(n1343) );
XNOR2_X1 U1062 ( .A(n1346), .B(n1030), .ZN(n1345) );
INV_X1 U1063 ( .A(G107), .ZN(n1030) );
NAND3_X1 U1064 ( .A1(G234), .A2(n1125), .A3(G217), .ZN(n1346) );
INV_X1 U1065 ( .A(G953), .ZN(n1125) );
NAND2_X1 U1066 ( .A1(n1347), .A2(KEYINPUT1), .ZN(n1344) );
XNOR2_X1 U1067 ( .A(G116), .B(n1309), .ZN(n1347) );
XOR2_X1 U1068 ( .A(n1348), .B(n1349), .Z(n1342) );
XNOR2_X1 U1069 ( .A(KEYINPUT3), .B(n1211), .ZN(n1349) );
XNOR2_X1 U1070 ( .A(G128), .B(G134), .ZN(n1348) );
XNOR2_X1 U1071 ( .A(n1350), .B(G475), .ZN(n1080) );
NAND2_X1 U1072 ( .A1(n1140), .A2(n1172), .ZN(n1350) );
INV_X1 U1073 ( .A(G902), .ZN(n1172) );
XNOR2_X1 U1074 ( .A(n1351), .B(n1352), .ZN(n1140) );
XOR2_X1 U1075 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1076 ( .A(n1355), .B(n1356), .Z(n1354) );
NOR2_X1 U1077 ( .A1(G113), .A2(KEYINPUT48), .ZN(n1356) );
NAND2_X1 U1078 ( .A1(KEYINPUT19), .A2(n1112), .ZN(n1355) );
INV_X1 U1079 ( .A(G131), .ZN(n1112) );
XNOR2_X1 U1080 ( .A(n1357), .B(n1211), .ZN(n1353) );
INV_X1 U1081 ( .A(G143), .ZN(n1211) );
NAND2_X1 U1082 ( .A1(G214), .A2(n1279), .ZN(n1357) );
NOR2_X1 U1083 ( .A1(G953), .A2(G237), .ZN(n1279) );
XNOR2_X1 U1084 ( .A(n1105), .B(n1358), .ZN(n1351) );
XNOR2_X1 U1085 ( .A(n1359), .B(n1309), .ZN(n1358) );
XOR2_X1 U1086 ( .A(G122), .B(KEYINPUT27), .Z(n1309) );
NAND2_X1 U1087 ( .A1(KEYINPUT33), .A2(n1143), .ZN(n1359) );
INV_X1 U1088 ( .A(G104), .ZN(n1143) );
XOR2_X1 U1089 ( .A(G140), .B(n1303), .Z(n1105) );
XOR2_X1 U1090 ( .A(G125), .B(G146), .Z(n1303) );
endmodule


