//Key = 1000101001100110111110100011110111101011011100000100110001101110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382;

NAND2_X1 U759 ( .A1(n1040), .A2(n1041), .ZN(G9) );
NAND2_X1 U760 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
XOR2_X1 U761 ( .A(KEYINPUT0), .B(n1044), .Z(n1040) );
NOR2_X1 U762 ( .A1(n1042), .A2(n1043), .ZN(n1044) );
INV_X1 U763 ( .A(G107), .ZN(n1043) );
NOR2_X1 U764 ( .A1(n1045), .A2(n1046), .ZN(G75) );
NOR3_X1 U765 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND3_X1 U766 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1047) );
NAND2_X1 U767 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U768 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND3_X1 U769 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
NAND3_X1 U770 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1058) );
NAND2_X1 U771 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U772 ( .A1(n1065), .A2(n1066), .ZN(n1060) );
NAND2_X1 U773 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U774 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND3_X1 U775 ( .A1(n1065), .A2(n1071), .A3(n1064), .ZN(n1055) );
NAND3_X1 U776 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
INV_X1 U777 ( .A(n1075), .ZN(n1074) );
NAND3_X1 U778 ( .A1(n1076), .A2(n1059), .A3(n1077), .ZN(n1073) );
NAND2_X1 U779 ( .A1(n1057), .A2(n1078), .ZN(n1072) );
INV_X1 U780 ( .A(n1079), .ZN(n1053) );
NOR3_X1 U781 ( .A1(n1080), .A2(G953), .A3(G952), .ZN(n1045) );
INV_X1 U782 ( .A(n1050), .ZN(n1080) );
NAND4_X1 U783 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1050) );
NOR3_X1 U784 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
XNOR2_X1 U785 ( .A(n1088), .B(KEYINPUT22), .ZN(n1086) );
NAND3_X1 U786 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1085) );
OR3_X1 U787 ( .A1(n1092), .A2(n1093), .A3(KEYINPUT6), .ZN(n1090) );
INV_X1 U788 ( .A(n1094), .ZN(n1092) );
NAND2_X1 U789 ( .A1(n1093), .A2(KEYINPUT6), .ZN(n1089) );
NOR3_X1 U790 ( .A1(n1095), .A2(n1069), .A3(n1077), .ZN(n1083) );
INV_X1 U791 ( .A(n1096), .ZN(n1077) );
AND2_X1 U792 ( .A1(n1097), .A2(G469), .ZN(n1095) );
NAND2_X1 U793 ( .A1(n1098), .A2(n1099), .ZN(n1082) );
INV_X1 U794 ( .A(n1100), .ZN(n1098) );
NAND2_X1 U795 ( .A1(n1101), .A2(n1102), .ZN(n1081) );
NAND4_X1 U796 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1101) );
NAND3_X1 U797 ( .A1(n1107), .A2(n1108), .A3(KEYINPUT6), .ZN(n1106) );
NAND2_X1 U798 ( .A1(n1109), .A2(n1110), .ZN(n1105) );
NAND2_X1 U799 ( .A1(n1111), .A2(n1100), .ZN(n1104) );
NAND2_X1 U800 ( .A1(n1112), .A2(n1113), .ZN(n1103) );
XOR2_X1 U801 ( .A(n1114), .B(n1115), .Z(G72) );
NOR2_X1 U802 ( .A1(n1116), .A2(n1051), .ZN(n1115) );
AND2_X1 U803 ( .A1(G227), .A2(G900), .ZN(n1116) );
NAND2_X1 U804 ( .A1(n1117), .A2(KEYINPUT39), .ZN(n1114) );
XOR2_X1 U805 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U806 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U807 ( .A(n1122), .B(n1123), .Z(n1121) );
XNOR2_X1 U808 ( .A(n1124), .B(n1125), .ZN(n1123) );
XOR2_X1 U809 ( .A(n1126), .B(n1127), .Z(n1122) );
XNOR2_X1 U810 ( .A(G134), .B(KEYINPUT15), .ZN(n1127) );
NAND2_X1 U811 ( .A1(KEYINPUT52), .A2(n1128), .ZN(n1126) );
NAND2_X1 U812 ( .A1(n1051), .A2(n1049), .ZN(n1118) );
NAND2_X1 U813 ( .A1(n1129), .A2(n1130), .ZN(G69) );
NAND2_X1 U814 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U815 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
OR2_X1 U816 ( .A1(n1051), .A2(G224), .ZN(n1134) );
INV_X1 U817 ( .A(n1135), .ZN(n1133) );
NAND2_X1 U818 ( .A1(n1136), .A2(n1137), .ZN(n1129) );
NAND2_X1 U819 ( .A1(G953), .A2(n1138), .ZN(n1137) );
NAND2_X1 U820 ( .A1(G898), .A2(G224), .ZN(n1138) );
INV_X1 U821 ( .A(n1132), .ZN(n1136) );
NAND2_X1 U822 ( .A1(KEYINPUT20), .A2(n1139), .ZN(n1132) );
XOR2_X1 U823 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U824 ( .A1(n1135), .A2(n1142), .ZN(n1141) );
XOR2_X1 U825 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U826 ( .A1(n1145), .A2(n1146), .ZN(n1140) );
XNOR2_X1 U827 ( .A(KEYINPUT44), .B(n1051), .ZN(n1146) );
NOR2_X1 U828 ( .A1(n1147), .A2(n1148), .ZN(G66) );
XNOR2_X1 U829 ( .A(n1149), .B(n1112), .ZN(n1148) );
NOR2_X1 U830 ( .A1(n1113), .A2(n1150), .ZN(n1149) );
NOR2_X1 U831 ( .A1(n1147), .A2(n1151), .ZN(G63) );
XNOR2_X1 U832 ( .A(n1107), .B(n1152), .ZN(n1151) );
NOR2_X1 U833 ( .A1(n1108), .A2(n1150), .ZN(n1152) );
NOR2_X1 U834 ( .A1(n1147), .A2(n1153), .ZN(G60) );
XNOR2_X1 U835 ( .A(n1154), .B(n1155), .ZN(n1153) );
NOR2_X1 U836 ( .A1(n1156), .A2(n1150), .ZN(n1155) );
XNOR2_X1 U837 ( .A(G475), .B(KEYINPUT50), .ZN(n1156) );
NAND2_X1 U838 ( .A1(n1157), .A2(n1158), .ZN(G6) );
NAND2_X1 U839 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U840 ( .A(KEYINPUT18), .B(n1161), .Z(n1157) );
NOR2_X1 U841 ( .A1(n1159), .A2(n1160), .ZN(n1161) );
NOR2_X1 U842 ( .A1(n1147), .A2(n1162), .ZN(G57) );
XOR2_X1 U843 ( .A(n1163), .B(n1164), .Z(n1162) );
XNOR2_X1 U844 ( .A(n1165), .B(n1166), .ZN(n1164) );
XOR2_X1 U845 ( .A(n1167), .B(n1168), .Z(n1163) );
XNOR2_X1 U846 ( .A(KEYINPUT49), .B(n1169), .ZN(n1168) );
NOR2_X1 U847 ( .A1(n1170), .A2(n1150), .ZN(n1167) );
NOR2_X1 U848 ( .A1(n1147), .A2(n1171), .ZN(G54) );
XOR2_X1 U849 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U850 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U851 ( .A1(n1110), .A2(n1150), .ZN(n1174) );
XOR2_X1 U852 ( .A(n1176), .B(n1177), .Z(n1172) );
XOR2_X1 U853 ( .A(KEYINPUT5), .B(n1178), .Z(n1177) );
NOR2_X1 U854 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XOR2_X1 U855 ( .A(n1181), .B(KEYINPUT62), .Z(n1180) );
NAND2_X1 U856 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NOR2_X1 U857 ( .A1(n1182), .A2(n1183), .ZN(n1179) );
XNOR2_X1 U858 ( .A(KEYINPUT43), .B(G110), .ZN(n1182) );
NAND2_X1 U859 ( .A1(KEYINPUT61), .A2(n1184), .ZN(n1176) );
NOR2_X1 U860 ( .A1(n1147), .A2(n1185), .ZN(G51) );
XOR2_X1 U861 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U862 ( .A(n1188), .B(n1189), .Z(n1187) );
NAND2_X1 U863 ( .A1(KEYINPUT27), .A2(n1190), .ZN(n1189) );
NAND3_X1 U864 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1188) );
NAND2_X1 U865 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NAND2_X1 U866 ( .A1(n1196), .A2(n1197), .ZN(n1192) );
INV_X1 U867 ( .A(KEYINPUT31), .ZN(n1197) );
NAND2_X1 U868 ( .A1(n1198), .A2(n1199), .ZN(n1196) );
XNOR2_X1 U869 ( .A(KEYINPUT14), .B(n1200), .ZN(n1198) );
NAND2_X1 U870 ( .A1(KEYINPUT31), .A2(n1201), .ZN(n1191) );
NAND2_X1 U871 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
OR2_X1 U872 ( .A1(n1200), .A2(KEYINPUT14), .ZN(n1203) );
NAND3_X1 U873 ( .A1(n1200), .A2(n1199), .A3(KEYINPUT14), .ZN(n1202) );
INV_X1 U874 ( .A(n1195), .ZN(n1200) );
NOR3_X1 U875 ( .A1(n1150), .A2(KEYINPUT40), .A3(n1100), .ZN(n1186) );
NAND2_X1 U876 ( .A1(G902), .A2(n1204), .ZN(n1150) );
NAND2_X1 U877 ( .A1(n1205), .A2(n1145), .ZN(n1204) );
INV_X1 U878 ( .A(n1048), .ZN(n1145) );
NAND4_X1 U879 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1048) );
NOR4_X1 U880 ( .A1(n1159), .A2(n1042), .A3(n1210), .A4(n1211), .ZN(n1209) );
INV_X1 U881 ( .A(n1212), .ZN(n1210) );
AND4_X1 U882 ( .A1(n1213), .A2(n1078), .A3(n1065), .A4(n1214), .ZN(n1042) );
AND4_X1 U883 ( .A1(n1215), .A2(n1213), .A3(n1065), .A4(n1214), .ZN(n1159) );
OR2_X1 U884 ( .A1(n1216), .A2(n1217), .ZN(n1208) );
NAND3_X1 U885 ( .A1(n1213), .A2(n1075), .A3(n1218), .ZN(n1206) );
NAND2_X1 U886 ( .A1(n1219), .A2(n1220), .ZN(n1075) );
NAND2_X1 U887 ( .A1(n1057), .A2(n1215), .ZN(n1220) );
NAND2_X1 U888 ( .A1(n1059), .A2(n1214), .ZN(n1219) );
XOR2_X1 U889 ( .A(n1049), .B(KEYINPUT13), .Z(n1205) );
NAND4_X1 U890 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1049) );
NOR3_X1 U891 ( .A1(n1225), .A2(n1226), .A3(n1227), .ZN(n1224) );
INV_X1 U892 ( .A(n1228), .ZN(n1227) );
NOR3_X1 U893 ( .A1(n1229), .A2(n1061), .A3(n1230), .ZN(n1225) );
NAND3_X1 U894 ( .A1(n1231), .A2(n1232), .A3(n1078), .ZN(n1229) );
OR2_X1 U895 ( .A1(n1233), .A2(n1234), .ZN(n1223) );
NAND2_X1 U896 ( .A1(n1235), .A2(n1215), .ZN(n1222) );
INV_X1 U897 ( .A(n1236), .ZN(n1235) );
NAND2_X1 U898 ( .A1(n1237), .A2(n1238), .ZN(n1221) );
NAND4_X1 U899 ( .A1(n1239), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1238) );
NAND4_X1 U900 ( .A1(n1243), .A2(n1218), .A3(n1244), .A4(n1087), .ZN(n1242) );
NAND3_X1 U901 ( .A1(n1078), .A2(n1230), .A3(n1245), .ZN(n1241) );
INV_X1 U902 ( .A(KEYINPUT56), .ZN(n1230) );
NAND3_X1 U903 ( .A1(n1064), .A2(n1246), .A3(n1059), .ZN(n1240) );
NAND2_X1 U904 ( .A1(n1215), .A2(n1247), .ZN(n1239) );
NAND2_X1 U905 ( .A1(n1061), .A2(n1248), .ZN(n1247) );
NAND3_X1 U906 ( .A1(n1249), .A2(n1233), .A3(n1063), .ZN(n1248) );
INV_X1 U907 ( .A(KEYINPUT58), .ZN(n1233) );
NOR2_X1 U908 ( .A1(n1051), .A2(G952), .ZN(n1147) );
XNOR2_X1 U909 ( .A(G146), .B(n1228), .ZN(G48) );
NAND4_X1 U910 ( .A1(n1215), .A2(n1246), .A3(n1237), .A4(n1244), .ZN(n1228) );
XNOR2_X1 U911 ( .A(G143), .B(n1250), .ZN(G45) );
NAND4_X1 U912 ( .A1(n1218), .A2(n1237), .A3(n1251), .A4(n1243), .ZN(n1250) );
NOR2_X1 U913 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
XNOR2_X1 U914 ( .A(n1244), .B(KEYINPUT48), .ZN(n1253) );
XOR2_X1 U915 ( .A(n1234), .B(n1254), .Z(G42) );
NAND2_X1 U916 ( .A1(KEYINPUT36), .A2(G140), .ZN(n1254) );
NAND4_X1 U917 ( .A1(n1063), .A2(n1064), .A3(n1215), .A4(n1237), .ZN(n1234) );
NAND3_X1 U918 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(G39) );
NAND2_X1 U919 ( .A1(G137), .A2(n1258), .ZN(n1257) );
NAND2_X1 U920 ( .A1(KEYINPUT47), .A2(n1259), .ZN(n1256) );
NAND2_X1 U921 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
INV_X1 U922 ( .A(n1258), .ZN(n1261) );
XNOR2_X1 U923 ( .A(KEYINPUT59), .B(G137), .ZN(n1260) );
NAND2_X1 U924 ( .A1(n1262), .A2(n1263), .ZN(n1255) );
INV_X1 U925 ( .A(KEYINPUT47), .ZN(n1263) );
NAND2_X1 U926 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
OR3_X1 U927 ( .A1(n1258), .A2(G137), .A3(KEYINPUT59), .ZN(n1265) );
NAND4_X1 U928 ( .A1(n1064), .A2(n1246), .A3(n1237), .A4(n1266), .ZN(n1258) );
XOR2_X1 U929 ( .A(KEYINPUT25), .B(n1059), .Z(n1266) );
NAND2_X1 U930 ( .A1(KEYINPUT59), .A2(G137), .ZN(n1264) );
XOR2_X1 U931 ( .A(n1267), .B(n1268), .Z(G36) );
XNOR2_X1 U932 ( .A(KEYINPUT45), .B(n1269), .ZN(n1268) );
NOR2_X1 U933 ( .A1(n1270), .A2(n1061), .ZN(n1267) );
XNOR2_X1 U934 ( .A(G131), .B(n1271), .ZN(G33) );
NAND4_X1 U935 ( .A1(n1245), .A2(n1215), .A3(n1272), .A4(n1231), .ZN(n1271) );
XNOR2_X1 U936 ( .A(KEYINPUT1), .B(n1232), .ZN(n1272) );
INV_X1 U937 ( .A(n1061), .ZN(n1245) );
NAND2_X1 U938 ( .A1(n1218), .A2(n1064), .ZN(n1061) );
INV_X1 U939 ( .A(n1249), .ZN(n1064) );
NAND2_X1 U940 ( .A1(n1070), .A2(n1273), .ZN(n1249) );
XNOR2_X1 U941 ( .A(n1274), .B(n1226), .ZN(G30) );
NOR3_X1 U942 ( .A1(n1270), .A2(n1067), .A3(n1275), .ZN(n1226) );
NAND2_X1 U943 ( .A1(n1237), .A2(n1078), .ZN(n1270) );
AND2_X1 U944 ( .A1(n1214), .A2(n1231), .ZN(n1237) );
XNOR2_X1 U945 ( .A(G101), .B(n1276), .ZN(G3) );
NAND4_X1 U946 ( .A1(n1059), .A2(n1218), .A3(n1277), .A4(n1214), .ZN(n1276) );
NOR2_X1 U947 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
XNOR2_X1 U948 ( .A(n1244), .B(KEYINPUT3), .ZN(n1279) );
XOR2_X1 U949 ( .A(G125), .B(n1280), .Z(G27) );
NOR2_X1 U950 ( .A1(n1281), .A2(n1236), .ZN(n1280) );
NAND4_X1 U951 ( .A1(n1063), .A2(n1057), .A3(n1244), .A4(n1231), .ZN(n1236) );
NAND2_X1 U952 ( .A1(n1282), .A2(n1283), .ZN(n1231) );
NAND2_X1 U953 ( .A1(n1120), .A2(n1284), .ZN(n1283) );
NOR2_X1 U954 ( .A1(n1051), .A2(G900), .ZN(n1120) );
XNOR2_X1 U955 ( .A(KEYINPUT60), .B(n1079), .ZN(n1282) );
XNOR2_X1 U956 ( .A(n1215), .B(KEYINPUT23), .ZN(n1281) );
NAND2_X1 U957 ( .A1(n1285), .A2(n1286), .ZN(G24) );
OR2_X1 U958 ( .A1(n1207), .A2(n1287), .ZN(n1286) );
XOR2_X1 U959 ( .A(n1288), .B(KEYINPUT35), .Z(n1285) );
NAND2_X1 U960 ( .A1(n1287), .A2(n1207), .ZN(n1288) );
NAND3_X1 U961 ( .A1(n1057), .A2(n1213), .A3(n1289), .ZN(n1207) );
AND3_X1 U962 ( .A1(n1065), .A2(n1087), .A3(n1243), .ZN(n1289) );
NOR2_X1 U963 ( .A1(n1290), .A2(n1291), .ZN(n1065) );
XOR2_X1 U964 ( .A(G122), .B(KEYINPUT63), .Z(n1287) );
XOR2_X1 U965 ( .A(G119), .B(n1292), .Z(G21) );
NOR2_X1 U966 ( .A1(n1293), .A2(n1216), .ZN(n1292) );
NAND3_X1 U967 ( .A1(n1246), .A2(n1213), .A3(n1059), .ZN(n1216) );
INV_X1 U968 ( .A(n1275), .ZN(n1246) );
NAND2_X1 U969 ( .A1(n1291), .A2(n1290), .ZN(n1275) );
XNOR2_X1 U970 ( .A(n1057), .B(KEYINPUT2), .ZN(n1293) );
XOR2_X1 U971 ( .A(G116), .B(n1211), .Z(G18) );
AND4_X1 U972 ( .A1(n1057), .A2(n1218), .A3(n1213), .A4(n1078), .ZN(n1211) );
AND2_X1 U973 ( .A1(n1252), .A2(n1243), .ZN(n1078) );
XOR2_X1 U974 ( .A(n1294), .B(KEYINPUT21), .Z(n1243) );
INV_X1 U975 ( .A(n1217), .ZN(n1057) );
XNOR2_X1 U976 ( .A(G113), .B(n1295), .ZN(G15) );
NAND4_X1 U977 ( .A1(n1215), .A2(n1244), .A3(n1218), .A4(n1296), .ZN(n1295) );
NOR2_X1 U978 ( .A1(n1217), .A2(n1297), .ZN(n1296) );
XOR2_X1 U979 ( .A(KEYINPUT12), .B(n1278), .Z(n1297) );
NAND2_X1 U980 ( .A1(n1076), .A2(n1096), .ZN(n1217) );
XOR2_X1 U981 ( .A(n1298), .B(KEYINPUT29), .Z(n1076) );
NOR2_X1 U982 ( .A1(n1290), .A2(n1091), .ZN(n1218) );
NOR2_X1 U983 ( .A1(n1294), .A2(n1252), .ZN(n1215) );
INV_X1 U984 ( .A(n1087), .ZN(n1252) );
XNOR2_X1 U985 ( .A(G110), .B(n1212), .ZN(G12) );
NAND4_X1 U986 ( .A1(n1059), .A2(n1063), .A3(n1213), .A4(n1214), .ZN(n1212) );
INV_X1 U987 ( .A(n1232), .ZN(n1214) );
NAND2_X1 U988 ( .A1(n1298), .A2(n1096), .ZN(n1232) );
NAND2_X1 U989 ( .A1(n1299), .A2(n1300), .ZN(n1096) );
XOR2_X1 U990 ( .A(KEYINPUT54), .B(G221), .Z(n1299) );
XNOR2_X1 U991 ( .A(n1301), .B(n1110), .ZN(n1298) );
INV_X1 U992 ( .A(G469), .ZN(n1110) );
NAND2_X1 U993 ( .A1(KEYINPUT9), .A2(n1097), .ZN(n1301) );
NAND2_X1 U994 ( .A1(n1109), .A2(n1102), .ZN(n1097) );
XOR2_X1 U995 ( .A(n1302), .B(n1303), .Z(n1109) );
XNOR2_X1 U996 ( .A(n1183), .B(G110), .ZN(n1303) );
XNOR2_X1 U997 ( .A(n1175), .B(n1184), .ZN(n1302) );
AND2_X1 U998 ( .A1(G227), .A2(n1051), .ZN(n1184) );
XNOR2_X1 U999 ( .A(n1304), .B(n1305), .ZN(n1175) );
XNOR2_X1 U1000 ( .A(n1160), .B(n1306), .ZN(n1305) );
NOR2_X1 U1001 ( .A1(G107), .A2(KEYINPUT7), .ZN(n1306) );
XNOR2_X1 U1002 ( .A(n1165), .B(n1128), .ZN(n1304) );
NAND2_X1 U1003 ( .A1(n1307), .A2(n1308), .ZN(n1128) );
OR2_X1 U1004 ( .A1(n1309), .A2(KEYINPUT11), .ZN(n1308) );
NAND3_X1 U1005 ( .A1(n1310), .A2(n1274), .A3(KEYINPUT11), .ZN(n1307) );
XNOR2_X1 U1006 ( .A(n1311), .B(G101), .ZN(n1165) );
NOR2_X1 U1007 ( .A1(n1067), .A2(n1278), .ZN(n1213) );
AND2_X1 U1008 ( .A1(n1079), .A2(n1312), .ZN(n1278) );
NAND2_X1 U1009 ( .A1(n1135), .A2(n1284), .ZN(n1312) );
AND2_X1 U1010 ( .A1(n1313), .A2(n1314), .ZN(n1284) );
XNOR2_X1 U1011 ( .A(G902), .B(KEYINPUT41), .ZN(n1313) );
NOR2_X1 U1012 ( .A1(n1051), .A2(G898), .ZN(n1135) );
NAND3_X1 U1013 ( .A1(n1314), .A2(n1051), .A3(G952), .ZN(n1079) );
NAND2_X1 U1014 ( .A1(G237), .A2(G234), .ZN(n1314) );
INV_X1 U1015 ( .A(n1244), .ZN(n1067) );
NOR2_X1 U1016 ( .A1(n1070), .A2(n1069), .ZN(n1244) );
INV_X1 U1017 ( .A(n1273), .ZN(n1069) );
NAND2_X1 U1018 ( .A1(G214), .A2(n1315), .ZN(n1273) );
XOR2_X1 U1019 ( .A(n1316), .B(n1100), .Z(n1070) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1315), .ZN(n1100) );
NAND2_X1 U1021 ( .A1(n1317), .A2(n1102), .ZN(n1315) );
INV_X1 U1022 ( .A(G237), .ZN(n1317) );
NAND2_X1 U1023 ( .A1(KEYINPUT28), .A2(n1099), .ZN(n1316) );
NAND2_X1 U1024 ( .A1(n1111), .A2(n1102), .ZN(n1099) );
XNOR2_X1 U1025 ( .A(n1318), .B(n1319), .ZN(n1111) );
XNOR2_X1 U1026 ( .A(n1195), .B(n1194), .ZN(n1319) );
INV_X1 U1027 ( .A(n1199), .ZN(n1194) );
XOR2_X1 U1028 ( .A(G125), .B(n1309), .Z(n1199) );
NAND2_X1 U1029 ( .A1(G224), .A2(n1051), .ZN(n1195) );
XOR2_X1 U1030 ( .A(n1190), .B(KEYINPUT32), .Z(n1318) );
NAND2_X1 U1031 ( .A1(n1320), .A2(n1321), .ZN(n1190) );
OR2_X1 U1032 ( .A1(n1322), .A2(n1143), .ZN(n1321) );
XOR2_X1 U1033 ( .A(n1323), .B(KEYINPUT55), .Z(n1320) );
NAND2_X1 U1034 ( .A1(n1143), .A2(n1322), .ZN(n1323) );
XNOR2_X1 U1035 ( .A(n1144), .B(KEYINPUT46), .ZN(n1322) );
XNOR2_X1 U1036 ( .A(G110), .B(n1324), .ZN(n1144) );
NOR2_X1 U1037 ( .A1(G122), .A2(KEYINPUT51), .ZN(n1324) );
XOR2_X1 U1038 ( .A(n1325), .B(n1326), .Z(n1143) );
XOR2_X1 U1039 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1040 ( .A(G107), .B(KEYINPUT16), .ZN(n1328) );
NAND2_X1 U1041 ( .A1(KEYINPUT4), .A2(n1329), .ZN(n1327) );
INV_X1 U1042 ( .A(G101), .ZN(n1329) );
XOR2_X1 U1043 ( .A(n1330), .B(n1331), .Z(n1325) );
NAND2_X1 U1044 ( .A1(KEYINPUT57), .A2(n1160), .ZN(n1330) );
AND2_X1 U1045 ( .A1(n1091), .A2(n1290), .ZN(n1063) );
NAND2_X1 U1046 ( .A1(n1332), .A2(n1333), .ZN(n1290) );
NAND3_X1 U1047 ( .A1(n1112), .A2(n1102), .A3(n1334), .ZN(n1333) );
XOR2_X1 U1048 ( .A(n1113), .B(KEYINPUT24), .Z(n1334) );
XOR2_X1 U1049 ( .A(KEYINPUT33), .B(n1088), .Z(n1332) );
NOR2_X1 U1050 ( .A1(n1113), .A2(n1335), .ZN(n1088) );
AND2_X1 U1051 ( .A1(n1112), .A2(n1102), .ZN(n1335) );
XOR2_X1 U1052 ( .A(n1336), .B(n1337), .Z(n1112) );
XOR2_X1 U1053 ( .A(n1338), .B(n1339), .Z(n1337) );
XNOR2_X1 U1054 ( .A(G119), .B(n1340), .ZN(n1339) );
INV_X1 U1055 ( .A(G110), .ZN(n1340) );
XNOR2_X1 U1056 ( .A(n1341), .B(G137), .ZN(n1338) );
INV_X1 U1057 ( .A(G146), .ZN(n1341) );
XNOR2_X1 U1058 ( .A(n1342), .B(n1343), .ZN(n1336) );
XOR2_X1 U1059 ( .A(n1344), .B(n1345), .Z(n1343) );
NAND2_X1 U1060 ( .A1(G221), .A2(n1346), .ZN(n1345) );
NAND2_X1 U1061 ( .A1(KEYINPUT34), .A2(n1347), .ZN(n1344) );
XNOR2_X1 U1062 ( .A(KEYINPUT42), .B(n1274), .ZN(n1347) );
INV_X1 U1063 ( .A(n1125), .ZN(n1342) );
NAND2_X1 U1064 ( .A1(G217), .A2(n1300), .ZN(n1113) );
NAND2_X1 U1065 ( .A1(G234), .A2(n1102), .ZN(n1300) );
INV_X1 U1066 ( .A(n1291), .ZN(n1091) );
XOR2_X1 U1067 ( .A(n1348), .B(n1170), .Z(n1291) );
INV_X1 U1068 ( .A(G472), .ZN(n1170) );
NAND2_X1 U1069 ( .A1(n1349), .A2(n1102), .ZN(n1348) );
XNOR2_X1 U1070 ( .A(n1350), .B(n1351), .ZN(n1349) );
XNOR2_X1 U1071 ( .A(n1352), .B(n1353), .ZN(n1351) );
INV_X1 U1072 ( .A(n1311), .ZN(n1353) );
XNOR2_X1 U1073 ( .A(n1354), .B(n1124), .ZN(n1311) );
XOR2_X1 U1074 ( .A(G131), .B(G137), .Z(n1124) );
NAND2_X1 U1075 ( .A1(KEYINPUT26), .A2(n1269), .ZN(n1354) );
NOR2_X1 U1076 ( .A1(n1355), .A2(n1356), .ZN(n1352) );
XOR2_X1 U1077 ( .A(KEYINPUT30), .B(n1357), .Z(n1356) );
AND2_X1 U1078 ( .A1(n1358), .A2(G101), .ZN(n1357) );
NOR2_X1 U1079 ( .A1(G101), .A2(n1358), .ZN(n1355) );
XNOR2_X1 U1080 ( .A(n1169), .B(KEYINPUT37), .ZN(n1358) );
NAND2_X1 U1081 ( .A1(n1359), .A2(G210), .ZN(n1169) );
INV_X1 U1082 ( .A(n1166), .ZN(n1350) );
XNOR2_X1 U1083 ( .A(n1360), .B(n1331), .ZN(n1166) );
XOR2_X1 U1084 ( .A(G113), .B(n1361), .Z(n1331) );
XOR2_X1 U1085 ( .A(G119), .B(G116), .Z(n1361) );
XOR2_X1 U1086 ( .A(n1309), .B(KEYINPUT53), .Z(n1360) );
XOR2_X1 U1087 ( .A(G128), .B(n1310), .Z(n1309) );
NOR2_X1 U1088 ( .A1(n1087), .A2(n1294), .ZN(n1059) );
NAND3_X1 U1089 ( .A1(n1362), .A2(n1363), .A3(n1094), .ZN(n1294) );
NAND2_X1 U1090 ( .A1(n1364), .A2(n1108), .ZN(n1094) );
OR2_X1 U1091 ( .A1(G478), .A2(KEYINPUT38), .ZN(n1363) );
NAND2_X1 U1092 ( .A1(n1093), .A2(KEYINPUT38), .ZN(n1362) );
NOR2_X1 U1093 ( .A1(n1108), .A2(n1364), .ZN(n1093) );
NOR2_X1 U1094 ( .A1(n1365), .A2(G902), .ZN(n1364) );
INV_X1 U1095 ( .A(n1107), .ZN(n1365) );
XNOR2_X1 U1096 ( .A(n1366), .B(n1367), .ZN(n1107) );
XOR2_X1 U1097 ( .A(n1368), .B(n1369), .Z(n1367) );
XNOR2_X1 U1098 ( .A(G107), .B(n1370), .ZN(n1369) );
NOR2_X1 U1099 ( .A1(KEYINPUT8), .A2(n1371), .ZN(n1370) );
XNOR2_X1 U1100 ( .A(G143), .B(n1372), .ZN(n1371) );
NOR2_X1 U1101 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
AND2_X1 U1102 ( .A1(KEYINPUT10), .A2(n1274), .ZN(n1374) );
NOR2_X1 U1103 ( .A1(KEYINPUT17), .A2(n1274), .ZN(n1373) );
INV_X1 U1104 ( .A(G128), .ZN(n1274) );
NAND3_X1 U1105 ( .A1(G217), .A2(n1346), .A3(KEYINPUT19), .ZN(n1368) );
AND2_X1 U1106 ( .A1(G234), .A2(n1051), .ZN(n1346) );
INV_X1 U1107 ( .A(G953), .ZN(n1051) );
XNOR2_X1 U1108 ( .A(G116), .B(n1375), .ZN(n1366) );
XNOR2_X1 U1109 ( .A(n1269), .B(G122), .ZN(n1375) );
INV_X1 U1110 ( .A(G134), .ZN(n1269) );
INV_X1 U1111 ( .A(G478), .ZN(n1108) );
XNOR2_X1 U1112 ( .A(n1376), .B(G475), .ZN(n1087) );
NAND2_X1 U1113 ( .A1(n1154), .A2(n1102), .ZN(n1376) );
INV_X1 U1114 ( .A(G902), .ZN(n1102) );
XNOR2_X1 U1115 ( .A(n1377), .B(n1378), .ZN(n1154) );
XOR2_X1 U1116 ( .A(n1379), .B(n1380), .Z(n1378) );
XNOR2_X1 U1117 ( .A(G113), .B(n1160), .ZN(n1380) );
INV_X1 U1118 ( .A(G104), .ZN(n1160) );
XOR2_X1 U1119 ( .A(G131), .B(G122), .Z(n1379) );
XNOR2_X1 U1120 ( .A(n1381), .B(n1125), .ZN(n1377) );
XOR2_X1 U1121 ( .A(G125), .B(n1183), .Z(n1125) );
INV_X1 U1122 ( .A(G140), .ZN(n1183) );
XNOR2_X1 U1123 ( .A(n1382), .B(n1310), .ZN(n1381) );
XNOR2_X1 U1124 ( .A(G143), .B(G146), .ZN(n1310) );
NAND2_X1 U1125 ( .A1(n1359), .A2(G214), .ZN(n1382) );
NOR2_X1 U1126 ( .A1(G953), .A2(G237), .ZN(n1359) );
endmodule


