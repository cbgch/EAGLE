//Key = 0001100100110011101001010011010101111101011100011011000010001010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;

XOR2_X1 U764 ( .A(G107), .B(n1045), .Z(G9) );
NOR2_X1 U765 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U766 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR4_X1 U767 ( .A1(G953), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1049) );
NOR2_X1 U768 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U769 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U770 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U771 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U772 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U773 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U774 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U775 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR2_X1 U776 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR2_X1 U777 ( .A1(n1071), .A2(n1072), .ZN(n1063) );
NOR2_X1 U778 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U779 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NOR3_X1 U780 ( .A1(n1072), .A2(n1077), .A3(n1066), .ZN(n1059) );
NOR2_X1 U781 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U782 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR4_X1 U783 ( .A1(n1082), .A2(n1066), .A3(n1072), .A4(n1062), .ZN(n1055) );
NOR2_X1 U784 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR3_X1 U785 ( .A1(n1050), .A2(G953), .A3(G952), .ZN(n1048) );
AND4_X1 U786 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1050) );
NOR3_X1 U787 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
XNOR2_X1 U788 ( .A(n1092), .B(n1093), .ZN(n1091) );
NOR2_X1 U789 ( .A1(G478), .A2(KEYINPUT8), .ZN(n1093) );
NOR2_X1 U790 ( .A1(n1094), .A2(n1095), .ZN(n1090) );
NAND3_X1 U791 ( .A1(n1080), .A2(n1070), .A3(n1096), .ZN(n1089) );
NOR3_X1 U792 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1087) );
NOR2_X1 U793 ( .A1(KEYINPUT61), .A2(n1100), .ZN(n1099) );
AND2_X1 U794 ( .A1(n1101), .A2(KEYINPUT61), .ZN(n1098) );
XOR2_X1 U795 ( .A(n1102), .B(n1103), .Z(n1097) );
NOR2_X1 U796 ( .A1(KEYINPUT53), .A2(n1104), .ZN(n1103) );
XOR2_X1 U797 ( .A(n1105), .B(n1106), .Z(G72) );
NOR3_X1 U798 ( .A1(KEYINPUT55), .A2(n1107), .A3(n1108), .ZN(n1106) );
NOR2_X1 U799 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U800 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U801 ( .A1(G900), .A2(n1113), .ZN(n1111) );
INV_X1 U802 ( .A(n1114), .ZN(n1109) );
NOR2_X1 U803 ( .A1(n1112), .A2(n1114), .ZN(n1107) );
XOR2_X1 U804 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U805 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U806 ( .A1(KEYINPUT0), .A2(n1119), .ZN(n1117) );
INV_X1 U807 ( .A(G137), .ZN(n1119) );
XOR2_X1 U808 ( .A(n1120), .B(n1121), .Z(n1115) );
XOR2_X1 U809 ( .A(G134), .B(n1122), .Z(n1121) );
NOR2_X1 U810 ( .A1(KEYINPUT58), .A2(n1123), .ZN(n1122) );
XOR2_X1 U811 ( .A(G140), .B(G125), .Z(n1123) );
NAND2_X1 U812 ( .A1(KEYINPUT26), .A2(n1124), .ZN(n1120) );
XOR2_X1 U813 ( .A(KEYINPUT34), .B(G131), .Z(n1124) );
NOR2_X1 U814 ( .A1(G953), .A2(n1125), .ZN(n1112) );
AND2_X1 U815 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XNOR2_X1 U816 ( .A(KEYINPUT62), .B(n1128), .ZN(n1127) );
NOR2_X1 U817 ( .A1(n1113), .A2(n1129), .ZN(n1105) );
XOR2_X1 U818 ( .A(KEYINPUT20), .B(n1130), .Z(n1129) );
AND2_X1 U819 ( .A1(G227), .A2(G900), .ZN(n1130) );
XOR2_X1 U820 ( .A(n1131), .B(n1132), .Z(G69) );
XOR2_X1 U821 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U822 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U823 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XNOR2_X1 U824 ( .A(KEYINPUT21), .B(n1139), .ZN(n1138) );
XOR2_X1 U825 ( .A(KEYINPUT36), .B(G953), .Z(n1135) );
NAND4_X1 U826 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1133) );
NAND2_X1 U827 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
INV_X1 U828 ( .A(KEYINPUT19), .ZN(n1145) );
NAND2_X1 U829 ( .A1(n1146), .A2(KEYINPUT19), .ZN(n1142) );
XNOR2_X1 U830 ( .A(n1147), .B(n1148), .ZN(n1146) );
NAND2_X1 U831 ( .A1(n1149), .A2(n1147), .ZN(n1141) );
NAND2_X1 U832 ( .A1(G953), .A2(n1150), .ZN(n1140) );
NOR2_X1 U833 ( .A1(n1151), .A2(n1113), .ZN(n1131) );
NOR2_X1 U834 ( .A1(n1152), .A2(n1150), .ZN(n1151) );
NOR2_X1 U835 ( .A1(n1153), .A2(n1154), .ZN(G66) );
XOR2_X1 U836 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U837 ( .A1(n1095), .A2(n1157), .ZN(n1156) );
NOR2_X1 U838 ( .A1(n1153), .A2(n1158), .ZN(G63) );
NOR3_X1 U839 ( .A1(n1092), .A2(n1159), .A3(n1160), .ZN(n1158) );
NOR3_X1 U840 ( .A1(n1161), .A2(n1162), .A3(n1157), .ZN(n1160) );
INV_X1 U841 ( .A(G478), .ZN(n1162) );
NOR2_X1 U842 ( .A1(n1163), .A2(n1164), .ZN(n1159) );
AND2_X1 U843 ( .A1(n1052), .A2(G478), .ZN(n1163) );
NOR2_X1 U844 ( .A1(n1165), .A2(n1166), .ZN(G60) );
XOR2_X1 U845 ( .A(n1167), .B(KEYINPUT12), .Z(n1166) );
NAND2_X1 U846 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U847 ( .A1(n1153), .A2(n1170), .ZN(n1169) );
INV_X1 U848 ( .A(KEYINPUT17), .ZN(n1170) );
NAND3_X1 U849 ( .A1(G953), .A2(G952), .A3(KEYINPUT17), .ZN(n1168) );
XNOR2_X1 U850 ( .A(n1171), .B(n1172), .ZN(n1165) );
NOR2_X1 U851 ( .A1(n1101), .A2(n1157), .ZN(n1172) );
INV_X1 U852 ( .A(G475), .ZN(n1101) );
XNOR2_X1 U853 ( .A(G104), .B(n1173), .ZN(G6) );
NOR2_X1 U854 ( .A1(n1153), .A2(n1174), .ZN(G57) );
XOR2_X1 U855 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U856 ( .A(n1177), .B(n1178), .ZN(n1176) );
XOR2_X1 U857 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U858 ( .A1(G101), .A2(KEYINPUT6), .ZN(n1180) );
XOR2_X1 U859 ( .A(n1181), .B(n1182), .Z(n1175) );
XOR2_X1 U860 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U861 ( .A1(n1185), .A2(n1157), .ZN(n1184) );
INV_X1 U862 ( .A(G472), .ZN(n1185) );
NAND2_X1 U863 ( .A1(KEYINPUT3), .A2(n1186), .ZN(n1181) );
NOR2_X1 U864 ( .A1(n1153), .A2(n1187), .ZN(G54) );
XOR2_X1 U865 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U866 ( .A(n1190), .B(n1191), .Z(n1189) );
NOR2_X1 U867 ( .A1(n1192), .A2(n1193), .ZN(n1190) );
XOR2_X1 U868 ( .A(n1194), .B(KEYINPUT7), .Z(n1193) );
NAND2_X1 U869 ( .A1(G110), .A2(n1195), .ZN(n1194) );
XOR2_X1 U870 ( .A(n1196), .B(n1197), .Z(n1188) );
NOR2_X1 U871 ( .A1(n1198), .A2(n1157), .ZN(n1197) );
INV_X1 U872 ( .A(G469), .ZN(n1198) );
NAND2_X1 U873 ( .A1(KEYINPUT56), .A2(n1199), .ZN(n1196) );
XOR2_X1 U874 ( .A(n1200), .B(n1201), .Z(n1199) );
NAND2_X1 U875 ( .A1(KEYINPUT31), .A2(n1118), .ZN(n1200) );
NOR2_X1 U876 ( .A1(n1153), .A2(n1202), .ZN(G51) );
NOR2_X1 U877 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
XOR2_X1 U878 ( .A(n1205), .B(n1206), .Z(n1204) );
NOR2_X1 U879 ( .A1(n1207), .A2(n1157), .ZN(n1206) );
NAND2_X1 U880 ( .A1(G902), .A2(n1052), .ZN(n1157) );
NAND4_X1 U881 ( .A1(n1137), .A2(n1126), .A3(n1139), .A4(n1128), .ZN(n1052) );
AND4_X1 U882 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1126) );
NOR4_X1 U883 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1211) );
OR2_X1 U884 ( .A1(n1216), .A2(n1072), .ZN(n1210) );
NAND3_X1 U885 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1209) );
XOR2_X1 U886 ( .A(n1058), .B(KEYINPUT4), .Z(n1219) );
INV_X1 U887 ( .A(n1220), .ZN(n1058) );
XOR2_X1 U888 ( .A(KEYINPUT44), .B(n1221), .Z(n1218) );
NAND2_X1 U889 ( .A1(n1222), .A2(n1079), .ZN(n1208) );
AND4_X1 U890 ( .A1(n1223), .A2(n1173), .A3(n1224), .A4(n1225), .ZN(n1137) );
NOR4_X1 U891 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1225) );
NOR4_X1 U892 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1229) );
XOR2_X1 U893 ( .A(n1047), .B(KEYINPUT57), .Z(n1233) );
XOR2_X1 U894 ( .A(n1234), .B(KEYINPUT43), .Z(n1232) );
NAND2_X1 U895 ( .A1(n1084), .A2(n1235), .ZN(n1230) );
NAND2_X1 U896 ( .A1(n1068), .A2(n1236), .ZN(n1224) );
XNOR2_X1 U897 ( .A(KEYINPUT1), .B(n1046), .ZN(n1236) );
NAND2_X1 U898 ( .A1(n1083), .A2(n1237), .ZN(n1046) );
NAND3_X1 U899 ( .A1(n1068), .A2(n1237), .A3(n1084), .ZN(n1173) );
AND3_X1 U900 ( .A1(n1238), .A2(n1234), .A3(n1079), .ZN(n1237) );
NAND3_X1 U901 ( .A1(n1074), .A2(n1079), .A3(n1239), .ZN(n1223) );
NOR2_X1 U902 ( .A1(KEYINPUT52), .A2(n1240), .ZN(n1205) );
XOR2_X1 U903 ( .A(n1241), .B(n1242), .Z(n1240) );
NOR2_X1 U904 ( .A1(n1243), .A2(n1244), .ZN(n1203) );
INV_X1 U905 ( .A(KEYINPUT52), .ZN(n1244) );
XOR2_X1 U906 ( .A(n1242), .B(n1245), .Z(n1243) );
XOR2_X1 U907 ( .A(n1246), .B(n1247), .Z(n1242) );
NAND2_X1 U908 ( .A1(KEYINPUT11), .A2(n1248), .ZN(n1246) );
NOR2_X1 U909 ( .A1(n1113), .A2(G952), .ZN(n1153) );
XOR2_X1 U910 ( .A(G146), .B(n1214), .Z(G48) );
AND3_X1 U911 ( .A1(n1084), .A2(n1068), .A3(n1217), .ZN(n1214) );
NAND2_X1 U912 ( .A1(n1249), .A2(n1250), .ZN(G45) );
NAND3_X1 U913 ( .A1(n1251), .A2(n1252), .A3(n1222), .ZN(n1250) );
INV_X1 U914 ( .A(G143), .ZN(n1252) );
XOR2_X1 U915 ( .A(n1253), .B(KEYINPUT5), .Z(n1249) );
NAND2_X1 U916 ( .A1(G143), .A2(n1254), .ZN(n1253) );
NAND2_X1 U917 ( .A1(n1222), .A2(n1251), .ZN(n1254) );
XOR2_X1 U918 ( .A(n1079), .B(KEYINPUT28), .Z(n1251) );
AND4_X1 U919 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1222) );
NOR2_X1 U920 ( .A1(n1047), .A2(n1231), .ZN(n1258) );
XOR2_X1 U921 ( .A(n1195), .B(n1259), .Z(G42) );
NAND2_X1 U922 ( .A1(n1260), .A2(n1221), .ZN(n1259) );
XOR2_X1 U923 ( .A(n1216), .B(KEYINPUT10), .Z(n1260) );
NAND3_X1 U924 ( .A1(n1261), .A2(n1255), .A3(n1084), .ZN(n1216) );
NAND2_X1 U925 ( .A1(n1262), .A2(n1263), .ZN(G39) );
NAND2_X1 U926 ( .A1(G137), .A2(n1264), .ZN(n1263) );
XOR2_X1 U927 ( .A(n1265), .B(KEYINPUT22), .Z(n1262) );
OR2_X1 U928 ( .A1(n1264), .A2(G137), .ZN(n1265) );
NAND3_X1 U929 ( .A1(n1220), .A2(n1221), .A3(n1217), .ZN(n1264) );
INV_X1 U930 ( .A(n1072), .ZN(n1221) );
NAND2_X1 U931 ( .A1(n1266), .A2(n1267), .ZN(G36) );
NAND2_X1 U932 ( .A1(G134), .A2(n1128), .ZN(n1267) );
XOR2_X1 U933 ( .A(n1268), .B(KEYINPUT40), .Z(n1266) );
OR2_X1 U934 ( .A1(n1128), .A2(G134), .ZN(n1268) );
NAND2_X1 U935 ( .A1(n1269), .A2(n1083), .ZN(n1128) );
XOR2_X1 U936 ( .A(G131), .B(n1215), .Z(G33) );
AND2_X1 U937 ( .A1(n1084), .A2(n1269), .ZN(n1215) );
NOR4_X1 U938 ( .A1(n1231), .A2(n1072), .A3(n1270), .A4(n1271), .ZN(n1269) );
NAND2_X1 U939 ( .A1(n1272), .A2(n1070), .ZN(n1072) );
INV_X1 U940 ( .A(n1069), .ZN(n1272) );
XOR2_X1 U941 ( .A(G128), .B(n1213), .Z(G30) );
AND3_X1 U942 ( .A1(n1068), .A2(n1083), .A3(n1217), .ZN(n1213) );
NOR4_X1 U943 ( .A1(n1270), .A2(n1086), .A3(n1271), .A4(n1075), .ZN(n1217) );
XOR2_X1 U944 ( .A(n1273), .B(n1274), .Z(G3) );
NAND4_X1 U945 ( .A1(KEYINPUT42), .A2(n1239), .A3(n1074), .A4(n1079), .ZN(n1274) );
INV_X1 U946 ( .A(n1270), .ZN(n1079) );
XOR2_X1 U947 ( .A(n1275), .B(n1212), .Z(G27) );
AND4_X1 U948 ( .A1(n1235), .A2(n1068), .A3(n1084), .A4(n1276), .ZN(n1212) );
NOR3_X1 U949 ( .A1(n1076), .A2(n1075), .A3(n1271), .ZN(n1276) );
INV_X1 U950 ( .A(n1255), .ZN(n1271) );
NAND2_X1 U951 ( .A1(n1054), .A2(n1277), .ZN(n1255) );
NAND4_X1 U952 ( .A1(G953), .A2(G902), .A3(n1278), .A4(n1279), .ZN(n1277) );
INV_X1 U953 ( .A(G900), .ZN(n1279) );
NAND2_X1 U954 ( .A1(KEYINPUT51), .A2(n1280), .ZN(n1275) );
INV_X1 U955 ( .A(G125), .ZN(n1280) );
XOR2_X1 U956 ( .A(n1281), .B(n1282), .Z(G24) );
NAND2_X1 U957 ( .A1(KEYINPUT14), .A2(n1228), .ZN(n1282) );
AND4_X1 U958 ( .A1(n1283), .A2(n1238), .A3(n1257), .A4(n1256), .ZN(n1228) );
INV_X1 U959 ( .A(n1066), .ZN(n1238) );
NAND2_X1 U960 ( .A1(n1075), .A2(n1086), .ZN(n1066) );
XNOR2_X1 U961 ( .A(G119), .B(n1284), .ZN(G21) );
NOR2_X1 U962 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NOR2_X1 U963 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
NAND4_X1 U964 ( .A1(n1239), .A2(n1076), .A3(n1289), .A4(n1062), .ZN(n1288) );
INV_X1 U965 ( .A(n1235), .ZN(n1062) );
INV_X1 U966 ( .A(KEYINPUT30), .ZN(n1287) );
NOR2_X1 U967 ( .A1(KEYINPUT30), .A2(n1139), .ZN(n1285) );
NAND4_X1 U968 ( .A1(n1239), .A2(n1235), .A3(n1076), .A4(n1289), .ZN(n1139) );
XOR2_X1 U969 ( .A(G116), .B(n1227), .Z(G18) );
AND3_X1 U970 ( .A1(n1074), .A2(n1083), .A3(n1283), .ZN(n1227) );
AND2_X1 U971 ( .A1(n1100), .A2(n1257), .ZN(n1083) );
XNOR2_X1 U972 ( .A(G113), .B(n1290), .ZN(G15) );
NAND3_X1 U973 ( .A1(n1283), .A2(n1074), .A3(n1084), .ZN(n1290) );
NOR2_X1 U974 ( .A1(n1257), .A2(n1100), .ZN(n1084) );
INV_X1 U975 ( .A(n1231), .ZN(n1074) );
NAND2_X1 U976 ( .A1(n1075), .A2(n1076), .ZN(n1231) );
AND3_X1 U977 ( .A1(n1068), .A2(n1234), .A3(n1235), .ZN(n1283) );
NOR2_X1 U978 ( .A1(n1081), .A2(n1291), .ZN(n1235) );
XOR2_X1 U979 ( .A(KEYINPUT37), .B(n1080), .Z(n1291) );
XNOR2_X1 U980 ( .A(n1226), .B(n1292), .ZN(G12) );
NAND2_X1 U981 ( .A1(KEYINPUT15), .A2(G110), .ZN(n1292) );
AND2_X1 U982 ( .A1(n1261), .A2(n1239), .ZN(n1226) );
AND3_X1 U983 ( .A1(n1068), .A2(n1234), .A3(n1220), .ZN(n1239) );
NOR2_X1 U984 ( .A1(n1257), .A2(n1256), .ZN(n1220) );
INV_X1 U985 ( .A(n1100), .ZN(n1256) );
XOR2_X1 U986 ( .A(n1293), .B(G475), .Z(n1100) );
NAND2_X1 U987 ( .A1(n1171), .A2(n1294), .ZN(n1293) );
XNOR2_X1 U988 ( .A(n1295), .B(n1296), .ZN(n1171) );
XOR2_X1 U989 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U990 ( .A(n1299), .B(n1300), .Z(n1298) );
AND3_X1 U991 ( .A1(G214), .A2(n1113), .A3(n1301), .ZN(n1300) );
NAND2_X1 U992 ( .A1(KEYINPUT23), .A2(G104), .ZN(n1299) );
XNOR2_X1 U993 ( .A(G113), .B(G131), .ZN(n1297) );
XOR2_X1 U994 ( .A(n1302), .B(n1303), .Z(n1295) );
XNOR2_X1 U995 ( .A(n1304), .B(n1305), .ZN(n1303) );
NOR2_X1 U996 ( .A1(KEYINPUT2), .A2(n1281), .ZN(n1305) );
NAND2_X1 U997 ( .A1(KEYINPUT27), .A2(G143), .ZN(n1304) );
XOR2_X1 U998 ( .A(n1092), .B(G478), .Z(n1257) );
NOR2_X1 U999 ( .A1(n1164), .A2(G902), .ZN(n1092) );
INV_X1 U1000 ( .A(n1161), .ZN(n1164) );
XOR2_X1 U1001 ( .A(n1306), .B(n1307), .Z(n1161) );
XOR2_X1 U1002 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U1003 ( .A(n1310), .B(n1311), .Z(n1309) );
NOR2_X1 U1004 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
INV_X1 U1005 ( .A(G217), .ZN(n1313) );
NAND2_X1 U1006 ( .A1(KEYINPUT18), .A2(n1281), .ZN(n1310) );
NAND2_X1 U1007 ( .A1(KEYINPUT47), .A2(n1314), .ZN(n1308) );
XNOR2_X1 U1008 ( .A(G107), .B(n1315), .ZN(n1306) );
XOR2_X1 U1009 ( .A(G134), .B(G116), .Z(n1315) );
NAND2_X1 U1010 ( .A1(n1316), .A2(n1054), .ZN(n1234) );
NAND3_X1 U1011 ( .A1(n1278), .A2(n1113), .A3(G952), .ZN(n1054) );
NAND4_X1 U1012 ( .A1(G953), .A2(G902), .A3(n1278), .A4(n1150), .ZN(n1316) );
INV_X1 U1013 ( .A(G898), .ZN(n1150) );
NAND2_X1 U1014 ( .A1(G234), .A2(G237), .ZN(n1278) );
INV_X1 U1015 ( .A(n1047), .ZN(n1068) );
NAND2_X1 U1016 ( .A1(n1069), .A2(n1070), .ZN(n1047) );
NAND2_X1 U1017 ( .A1(G214), .A2(n1317), .ZN(n1070) );
NAND2_X1 U1018 ( .A1(n1318), .A2(n1319), .ZN(n1069) );
NAND2_X1 U1019 ( .A1(n1102), .A2(n1104), .ZN(n1319) );
XOR2_X1 U1020 ( .A(KEYINPUT16), .B(n1320), .Z(n1318) );
NOR2_X1 U1021 ( .A1(n1102), .A2(n1104), .ZN(n1320) );
NAND2_X1 U1022 ( .A1(n1321), .A2(n1294), .ZN(n1104) );
XOR2_X1 U1023 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1024 ( .A(n1248), .B(n1324), .ZN(n1323) );
NAND2_X1 U1025 ( .A1(KEYINPUT48), .A2(n1245), .ZN(n1324) );
INV_X1 U1026 ( .A(n1241), .ZN(n1245) );
XNOR2_X1 U1027 ( .A(n1325), .B(n1314), .ZN(n1241) );
NOR2_X1 U1028 ( .A1(n1152), .A2(G953), .ZN(n1248) );
INV_X1 U1029 ( .A(G224), .ZN(n1152) );
XOR2_X1 U1030 ( .A(KEYINPUT60), .B(n1247), .Z(n1322) );
NOR2_X1 U1031 ( .A1(n1144), .A2(n1326), .ZN(n1247) );
AND2_X1 U1032 ( .A1(n1149), .A2(n1147), .ZN(n1326) );
NAND2_X1 U1033 ( .A1(n1327), .A2(n1328), .ZN(n1144) );
OR3_X1 U1034 ( .A1(n1147), .A2(n1149), .A3(n1329), .ZN(n1328) );
AND2_X1 U1035 ( .A1(n1330), .A2(n1148), .ZN(n1149) );
NAND2_X1 U1036 ( .A1(n1329), .A2(n1147), .ZN(n1327) );
XNOR2_X1 U1037 ( .A(n1281), .B(G110), .ZN(n1147) );
INV_X1 U1038 ( .A(G122), .ZN(n1281) );
NOR2_X1 U1039 ( .A1(n1148), .A2(n1330), .ZN(n1329) );
XNOR2_X1 U1040 ( .A(G113), .B(n1331), .ZN(n1330) );
NOR2_X1 U1041 ( .A1(KEYINPUT38), .A2(n1332), .ZN(n1331) );
XNOR2_X1 U1042 ( .A(KEYINPUT41), .B(n1333), .ZN(n1332) );
XOR2_X1 U1043 ( .A(n1334), .B(n1335), .Z(n1148) );
XOR2_X1 U1044 ( .A(n1273), .B(KEYINPUT63), .Z(n1334) );
INV_X1 U1045 ( .A(n1207), .ZN(n1102) );
NAND2_X1 U1046 ( .A1(G210), .A2(n1317), .ZN(n1207) );
NAND2_X1 U1047 ( .A1(n1336), .A2(n1337), .ZN(n1317) );
XOR2_X1 U1048 ( .A(n1301), .B(KEYINPUT13), .Z(n1336) );
NOR3_X1 U1049 ( .A1(n1076), .A2(n1075), .A3(n1270), .ZN(n1261) );
NAND2_X1 U1050 ( .A1(n1081), .A2(n1080), .ZN(n1270) );
NAND2_X1 U1051 ( .A1(G221), .A2(n1338), .ZN(n1080) );
XNOR2_X1 U1052 ( .A(n1085), .B(KEYINPUT24), .ZN(n1081) );
XOR2_X1 U1053 ( .A(n1339), .B(G469), .Z(n1085) );
NAND2_X1 U1054 ( .A1(n1340), .A2(n1294), .ZN(n1339) );
XOR2_X1 U1055 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1056 ( .A(n1343), .B(n1191), .Z(n1342) );
XOR2_X1 U1057 ( .A(n1344), .B(n1179), .Z(n1191) );
NAND2_X1 U1058 ( .A1(G227), .A2(n1113), .ZN(n1344) );
INV_X1 U1059 ( .A(n1201), .ZN(n1343) );
XOR2_X1 U1060 ( .A(n1345), .B(n1335), .Z(n1201) );
XOR2_X1 U1061 ( .A(G104), .B(G107), .Z(n1335) );
NAND2_X1 U1062 ( .A1(KEYINPUT35), .A2(n1273), .ZN(n1345) );
INV_X1 U1063 ( .A(G101), .ZN(n1273) );
XOR2_X1 U1064 ( .A(n1346), .B(n1118), .Z(n1341) );
XOR2_X1 U1065 ( .A(n1347), .B(n1348), .Z(n1118) );
NAND2_X1 U1066 ( .A1(KEYINPUT33), .A2(n1349), .ZN(n1347) );
XOR2_X1 U1067 ( .A(G143), .B(n1350), .Z(n1349) );
XOR2_X1 U1068 ( .A(KEYINPUT25), .B(G146), .Z(n1350) );
NOR3_X1 U1069 ( .A1(n1192), .A2(n1351), .A3(n1352), .ZN(n1346) );
NOR2_X1 U1070 ( .A1(KEYINPUT46), .A2(n1353), .ZN(n1352) );
NOR2_X1 U1071 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NOR2_X1 U1072 ( .A1(G110), .A2(n1356), .ZN(n1355) );
AND3_X1 U1073 ( .A1(n1356), .A2(n1195), .A3(G110), .ZN(n1354) );
NOR2_X1 U1074 ( .A1(n1357), .A2(n1358), .ZN(n1351) );
INV_X1 U1075 ( .A(KEYINPUT46), .ZN(n1358) );
NOR2_X1 U1076 ( .A1(G140), .A2(n1359), .ZN(n1357) );
XOR2_X1 U1077 ( .A(n1356), .B(G110), .Z(n1359) );
INV_X1 U1078 ( .A(KEYINPUT59), .ZN(n1356) );
NOR2_X1 U1079 ( .A1(n1195), .A2(G110), .ZN(n1192) );
INV_X1 U1080 ( .A(n1289), .ZN(n1075) );
NAND3_X1 U1081 ( .A1(n1360), .A2(n1361), .A3(n1096), .ZN(n1289) );
NAND2_X1 U1082 ( .A1(n1094), .A2(n1095), .ZN(n1096) );
NAND2_X1 U1083 ( .A1(n1095), .A2(n1362), .ZN(n1361) );
OR3_X1 U1084 ( .A1(n1095), .A2(n1094), .A3(n1362), .ZN(n1360) );
INV_X1 U1085 ( .A(KEYINPUT39), .ZN(n1362) );
NOR2_X1 U1086 ( .A1(n1155), .A2(G902), .ZN(n1094) );
XOR2_X1 U1087 ( .A(n1363), .B(n1364), .Z(n1155) );
XOR2_X1 U1088 ( .A(n1302), .B(n1365), .Z(n1364) );
XOR2_X1 U1089 ( .A(n1366), .B(n1367), .Z(n1365) );
NOR2_X1 U1090 ( .A1(n1312), .A2(n1368), .ZN(n1367) );
INV_X1 U1091 ( .A(G221), .ZN(n1368) );
NAND2_X1 U1092 ( .A1(n1369), .A2(n1113), .ZN(n1312) );
XNOR2_X1 U1093 ( .A(G234), .B(KEYINPUT29), .ZN(n1369) );
NAND2_X1 U1094 ( .A1(n1370), .A2(KEYINPUT50), .ZN(n1366) );
XOR2_X1 U1095 ( .A(n1348), .B(n1371), .Z(n1370) );
NOR2_X1 U1096 ( .A1(G119), .A2(KEYINPUT45), .ZN(n1371) );
INV_X1 U1097 ( .A(G128), .ZN(n1348) );
XOR2_X1 U1098 ( .A(n1195), .B(n1325), .Z(n1302) );
XOR2_X1 U1099 ( .A(G125), .B(G146), .Z(n1325) );
INV_X1 U1100 ( .A(G140), .ZN(n1195) );
XNOR2_X1 U1101 ( .A(G110), .B(n1372), .ZN(n1363) );
XOR2_X1 U1102 ( .A(KEYINPUT9), .B(G137), .Z(n1372) );
NAND2_X1 U1103 ( .A1(G217), .A2(n1338), .ZN(n1095) );
NAND2_X1 U1104 ( .A1(G234), .A2(n1337), .ZN(n1338) );
XOR2_X1 U1105 ( .A(n1294), .B(KEYINPUT32), .Z(n1337) );
INV_X1 U1106 ( .A(n1086), .ZN(n1076) );
XOR2_X1 U1107 ( .A(n1373), .B(G472), .Z(n1086) );
NAND2_X1 U1108 ( .A1(n1374), .A2(n1294), .ZN(n1373) );
INV_X1 U1109 ( .A(G902), .ZN(n1294) );
XOR2_X1 U1110 ( .A(n1375), .B(n1376), .Z(n1374) );
XNOR2_X1 U1111 ( .A(n1186), .B(n1177), .ZN(n1376) );
XOR2_X1 U1112 ( .A(G113), .B(n1377), .Z(n1177) );
NOR2_X1 U1113 ( .A1(KEYINPUT54), .A2(n1333), .ZN(n1377) );
XNOR2_X1 U1114 ( .A(G116), .B(G119), .ZN(n1333) );
XNOR2_X1 U1115 ( .A(G146), .B(n1314), .ZN(n1186) );
XOR2_X1 U1116 ( .A(G128), .B(G143), .Z(n1314) );
XOR2_X1 U1117 ( .A(n1378), .B(n1379), .Z(n1375) );
XOR2_X1 U1118 ( .A(G101), .B(n1183), .Z(n1379) );
AND3_X1 U1119 ( .A1(n1301), .A2(n1113), .A3(G210), .ZN(n1183) );
INV_X1 U1120 ( .A(G953), .ZN(n1113) );
INV_X1 U1121 ( .A(G237), .ZN(n1301) );
INV_X1 U1122 ( .A(n1179), .ZN(n1378) );
XNOR2_X1 U1123 ( .A(G131), .B(n1380), .ZN(n1179) );
NOR2_X1 U1124 ( .A1(KEYINPUT49), .A2(n1381), .ZN(n1380) );
XOR2_X1 U1125 ( .A(n1382), .B(G137), .Z(n1381) );
INV_X1 U1126 ( .A(G134), .ZN(n1382) );
endmodule


