//Key = 1010110100010000010100110011110101011101000110000101001110101110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354;

XNOR2_X1 U746 ( .A(G107), .B(n1030), .ZN(G9) );
NOR2_X1 U747 ( .A1(n1031), .A2(n1032), .ZN(G75) );
NOR4_X1 U748 ( .A1(G953), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1032) );
INV_X1 U749 ( .A(n1036), .ZN(n1035) );
NOR2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1034) );
NOR2_X1 U751 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR2_X1 U752 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR2_X1 U753 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR2_X1 U754 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U756 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U760 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(n1051) );
NOR2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR3_X1 U764 ( .A1(n1060), .A2(n1065), .A3(n1066), .ZN(n1047) );
XNOR2_X1 U765 ( .A(n1067), .B(KEYINPUT41), .ZN(n1066) );
NOR3_X1 U766 ( .A1(n1060), .A2(n1068), .A3(n1054), .ZN(n1043) );
INV_X1 U767 ( .A(n1067), .ZN(n1054) );
NOR3_X1 U768 ( .A1(n1046), .A2(n1065), .A3(n1049), .ZN(n1039) );
AND2_X1 U769 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
NAND3_X1 U770 ( .A1(n1071), .A2(n1072), .A3(n1067), .ZN(n1069) );
NAND2_X1 U771 ( .A1(n1073), .A2(n1060), .ZN(n1072) );
NAND2_X1 U772 ( .A1(KEYINPUT50), .A2(n1074), .ZN(n1073) );
NAND2_X1 U773 ( .A1(n1075), .A2(n1076), .ZN(n1071) );
NAND2_X1 U774 ( .A1(n1074), .A2(n1077), .ZN(n1075) );
NAND2_X1 U775 ( .A1(KEYINPUT50), .A2(n1078), .ZN(n1077) );
INV_X1 U776 ( .A(n1079), .ZN(n1046) );
NOR3_X1 U777 ( .A1(n1033), .A2(G953), .A3(G952), .ZN(n1031) );
AND4_X1 U778 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1033) );
NOR4_X1 U779 ( .A1(n1084), .A2(n1085), .A3(n1060), .A4(n1064), .ZN(n1083) );
XOR2_X1 U780 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND2_X1 U781 ( .A1(KEYINPUT56), .A2(n1088), .ZN(n1086) );
NOR3_X1 U782 ( .A1(n1049), .A2(n1089), .A3(n1090), .ZN(n1082) );
NAND2_X1 U783 ( .A1(G469), .A2(n1091), .ZN(n1081) );
NAND2_X1 U784 ( .A1(n1092), .A2(n1093), .ZN(n1080) );
XNOR2_X1 U785 ( .A(n1094), .B(KEYINPUT5), .ZN(n1092) );
XOR2_X1 U786 ( .A(n1095), .B(n1096), .Z(G72) );
NOR2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XNOR2_X1 U788 ( .A(G953), .B(KEYINPUT14), .ZN(n1098) );
AND2_X1 U789 ( .A1(G227), .A2(G900), .ZN(n1097) );
NAND2_X1 U790 ( .A1(n1099), .A2(n1100), .ZN(n1095) );
NAND2_X1 U791 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U792 ( .A(n1103), .B(n1104), .Z(n1101) );
NAND3_X1 U793 ( .A1(G900), .A2(n1104), .A3(G953), .ZN(n1099) );
XNOR2_X1 U794 ( .A(n1105), .B(n1106), .ZN(n1104) );
XNOR2_X1 U795 ( .A(G140), .B(n1107), .ZN(n1106) );
NAND3_X1 U796 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1107) );
OR2_X1 U797 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U798 ( .A1(KEYINPUT46), .A2(n1113), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1114), .A2(n1112), .ZN(n1113) );
XNOR2_X1 U800 ( .A(n1111), .B(KEYINPUT22), .ZN(n1114) );
NAND2_X1 U801 ( .A1(n1115), .A2(n1116), .ZN(n1108) );
INV_X1 U802 ( .A(KEYINPUT46), .ZN(n1116) );
NAND2_X1 U803 ( .A1(n1117), .A2(n1118), .ZN(n1115) );
OR2_X1 U804 ( .A1(n1111), .A2(KEYINPUT22), .ZN(n1118) );
NAND3_X1 U805 ( .A1(n1111), .A2(n1112), .A3(KEYINPUT22), .ZN(n1117) );
NAND2_X1 U806 ( .A1(KEYINPUT54), .A2(n1119), .ZN(n1105) );
XOR2_X1 U807 ( .A(n1120), .B(n1121), .Z(G69) );
AND2_X1 U808 ( .A1(n1122), .A2(n1102), .ZN(n1121) );
NAND2_X1 U809 ( .A1(n1123), .A2(n1124), .ZN(n1120) );
NAND2_X1 U810 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
INV_X1 U811 ( .A(n1127), .ZN(n1125) );
NAND2_X1 U812 ( .A1(n1128), .A2(n1127), .ZN(n1123) );
NAND2_X1 U813 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
XOR2_X1 U814 ( .A(n1131), .B(n1132), .Z(n1129) );
NOR2_X1 U815 ( .A1(KEYINPUT52), .A2(n1133), .ZN(n1131) );
XOR2_X1 U816 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U817 ( .A1(n1130), .A2(n1126), .ZN(n1128) );
NAND2_X1 U818 ( .A1(G953), .A2(n1136), .ZN(n1126) );
INV_X1 U819 ( .A(G224), .ZN(n1136) );
INV_X1 U820 ( .A(n1137), .ZN(n1130) );
NOR2_X1 U821 ( .A1(n1138), .A2(n1139), .ZN(G66) );
NOR3_X1 U822 ( .A1(n1094), .A2(n1140), .A3(n1141), .ZN(n1139) );
AND3_X1 U823 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1141) );
INV_X1 U824 ( .A(n1093), .ZN(n1143) );
NOR2_X1 U825 ( .A1(n1145), .A2(n1142), .ZN(n1140) );
NOR2_X1 U826 ( .A1(n1036), .A2(n1093), .ZN(n1145) );
NOR2_X1 U827 ( .A1(n1138), .A2(n1146), .ZN(G63) );
NOR3_X1 U828 ( .A1(n1087), .A2(n1147), .A3(n1148), .ZN(n1146) );
AND3_X1 U829 ( .A1(n1149), .A2(G478), .A3(n1144), .ZN(n1148) );
NOR2_X1 U830 ( .A1(n1150), .A2(n1149), .ZN(n1147) );
NOR2_X1 U831 ( .A1(n1036), .A2(n1088), .ZN(n1150) );
NOR2_X1 U832 ( .A1(n1138), .A2(n1151), .ZN(G60) );
XOR2_X1 U833 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U834 ( .A1(n1144), .A2(G475), .ZN(n1152) );
XNOR2_X1 U835 ( .A(G104), .B(n1154), .ZN(G6) );
NOR2_X1 U836 ( .A1(n1138), .A2(n1155), .ZN(G57) );
XOR2_X1 U837 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR2_X1 U838 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U839 ( .A(n1160), .B(n1161), .Z(n1159) );
NAND2_X1 U840 ( .A1(n1144), .A2(G472), .ZN(n1161) );
NAND2_X1 U841 ( .A1(n1162), .A2(n1163), .ZN(n1160) );
NOR2_X1 U842 ( .A1(n1162), .A2(n1163), .ZN(n1158) );
INV_X1 U843 ( .A(KEYINPUT21), .ZN(n1163) );
XOR2_X1 U844 ( .A(n1164), .B(n1165), .Z(n1162) );
NAND2_X1 U845 ( .A1(n1166), .A2(n1167), .ZN(n1164) );
NAND2_X1 U846 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XNOR2_X1 U847 ( .A(KEYINPUT60), .B(n1170), .ZN(n1168) );
XOR2_X1 U848 ( .A(KEYINPUT35), .B(n1171), .Z(n1166) );
NOR2_X1 U849 ( .A1(n1172), .A2(n1169), .ZN(n1171) );
XNOR2_X1 U850 ( .A(n1173), .B(KEYINPUT3), .ZN(n1172) );
NOR2_X1 U851 ( .A1(n1138), .A2(n1174), .ZN(G54) );
XOR2_X1 U852 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U853 ( .A(n1177), .B(n1178), .Z(n1176) );
XNOR2_X1 U854 ( .A(G110), .B(n1179), .ZN(n1178) );
XOR2_X1 U855 ( .A(KEYINPUT6), .B(G140), .Z(n1177) );
XOR2_X1 U856 ( .A(n1180), .B(n1181), .Z(n1175) );
XNOR2_X1 U857 ( .A(n1182), .B(n1183), .ZN(n1180) );
NAND2_X1 U858 ( .A1(KEYINPUT49), .A2(n1184), .ZN(n1183) );
INV_X1 U859 ( .A(n1111), .ZN(n1184) );
NAND2_X1 U860 ( .A1(KEYINPUT7), .A2(n1185), .ZN(n1182) );
NAND2_X1 U861 ( .A1(n1144), .A2(G469), .ZN(n1185) );
NOR2_X1 U862 ( .A1(n1138), .A2(n1186), .ZN(G51) );
XOR2_X1 U863 ( .A(n1187), .B(n1188), .Z(n1186) );
XNOR2_X1 U864 ( .A(n1189), .B(n1190), .ZN(n1188) );
NAND2_X1 U865 ( .A1(n1144), .A2(n1191), .ZN(n1189) );
NOR2_X1 U866 ( .A1(n1192), .A2(n1036), .ZN(n1144) );
NOR2_X1 U867 ( .A1(n1122), .A2(n1103), .ZN(n1036) );
NAND4_X1 U868 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1103) );
AND4_X1 U869 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1196) );
NAND2_X1 U870 ( .A1(n1056), .A2(n1201), .ZN(n1195) );
XOR2_X1 U871 ( .A(KEYINPUT48), .B(n1202), .Z(n1201) );
NAND3_X1 U872 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1193) );
NAND2_X1 U873 ( .A1(n1206), .A2(n1207), .ZN(n1204) );
NAND3_X1 U874 ( .A1(n1208), .A2(n1209), .A3(KEYINPUT63), .ZN(n1206) );
NAND3_X1 U875 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1203) );
OR3_X1 U876 ( .A1(n1213), .A2(KEYINPUT63), .A3(n1076), .ZN(n1211) );
NAND2_X1 U877 ( .A1(n1214), .A2(n1074), .ZN(n1210) );
XNOR2_X1 U878 ( .A(n1213), .B(KEYINPUT34), .ZN(n1214) );
NAND4_X1 U879 ( .A1(n1154), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1122) );
NOR4_X1 U880 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1217) );
AND2_X1 U881 ( .A1(n1030), .A2(n1222), .ZN(n1216) );
NAND2_X1 U882 ( .A1(n1223), .A2(n1074), .ZN(n1030) );
NAND2_X1 U883 ( .A1(n1208), .A2(n1223), .ZN(n1154) );
AND3_X1 U884 ( .A1(n1067), .A2(n1224), .A3(n1205), .ZN(n1223) );
XOR2_X1 U885 ( .A(n1225), .B(n1226), .Z(n1187) );
NOR2_X1 U886 ( .A1(KEYINPUT10), .A2(n1227), .ZN(n1226) );
NAND2_X1 U887 ( .A1(n1228), .A2(n1119), .ZN(n1225) );
XNOR2_X1 U888 ( .A(KEYINPUT42), .B(KEYINPUT20), .ZN(n1228) );
NOR2_X1 U889 ( .A1(n1102), .A2(G952), .ZN(n1138) );
XOR2_X1 U890 ( .A(n1229), .B(n1230), .Z(G48) );
NOR2_X1 U891 ( .A1(n1076), .A2(n1231), .ZN(n1230) );
NOR2_X1 U892 ( .A1(KEYINPUT18), .A2(n1232), .ZN(n1229) );
XNOR2_X1 U893 ( .A(G143), .B(n1233), .ZN(G45) );
NAND3_X1 U894 ( .A1(n1202), .A2(n1056), .A3(KEYINPUT62), .ZN(n1233) );
AND4_X1 U895 ( .A1(n1234), .A2(n1062), .A3(n1235), .A4(n1236), .ZN(n1202) );
NOR2_X1 U896 ( .A1(n1213), .A2(n1237), .ZN(n1235) );
XNOR2_X1 U897 ( .A(G140), .B(n1200), .ZN(G42) );
NAND2_X1 U898 ( .A1(n1238), .A2(n1239), .ZN(n1200) );
XNOR2_X1 U899 ( .A(G137), .B(n1199), .ZN(G39) );
NAND3_X1 U900 ( .A1(n1212), .A2(n1240), .A3(n1238), .ZN(n1199) );
XNOR2_X1 U901 ( .A(G134), .B(n1198), .ZN(G36) );
NAND3_X1 U902 ( .A1(n1062), .A2(n1074), .A3(n1238), .ZN(n1198) );
NAND2_X1 U903 ( .A1(n1241), .A2(n1242), .ZN(G33) );
NAND2_X1 U904 ( .A1(G131), .A2(n1194), .ZN(n1242) );
XOR2_X1 U905 ( .A(n1243), .B(KEYINPUT59), .Z(n1241) );
OR2_X1 U906 ( .A1(n1194), .A2(G131), .ZN(n1243) );
NAND3_X1 U907 ( .A1(n1062), .A2(n1208), .A3(n1238), .ZN(n1194) );
NOR3_X1 U908 ( .A1(n1068), .A2(n1213), .A3(n1060), .ZN(n1238) );
INV_X1 U909 ( .A(n1078), .ZN(n1060) );
NOR2_X1 U910 ( .A1(n1057), .A2(n1244), .ZN(n1078) );
INV_X1 U911 ( .A(n1058), .ZN(n1244) );
XNOR2_X1 U912 ( .A(G128), .B(n1245), .ZN(G30) );
NAND2_X1 U913 ( .A1(n1246), .A2(n1074), .ZN(n1245) );
INV_X1 U914 ( .A(n1231), .ZN(n1246) );
NAND3_X1 U915 ( .A1(n1205), .A2(n1209), .A3(n1212), .ZN(n1231) );
XOR2_X1 U916 ( .A(n1221), .B(n1247), .Z(G3) );
NOR2_X1 U917 ( .A1(KEYINPUT1), .A2(n1248), .ZN(n1247) );
NOR2_X1 U918 ( .A1(n1249), .A2(n1250), .ZN(n1221) );
XNOR2_X1 U919 ( .A(G125), .B(n1197), .ZN(G27) );
NAND3_X1 U920 ( .A1(n1239), .A2(n1079), .A3(n1251), .ZN(n1197) );
NOR3_X1 U921 ( .A1(n1252), .A2(n1049), .A3(n1213), .ZN(n1251) );
INV_X1 U922 ( .A(n1209), .ZN(n1213) );
NAND2_X1 U923 ( .A1(n1038), .A2(n1253), .ZN(n1209) );
NAND4_X1 U924 ( .A1(n1254), .A2(G953), .A3(G902), .A4(n1255), .ZN(n1253) );
INV_X1 U925 ( .A(G900), .ZN(n1255) );
XOR2_X1 U926 ( .A(n1256), .B(KEYINPUT13), .Z(n1254) );
NOR3_X1 U927 ( .A1(n1064), .A2(n1063), .A3(n1076), .ZN(n1239) );
XNOR2_X1 U928 ( .A(G122), .B(n1215), .ZN(G24) );
NAND4_X1 U929 ( .A1(n1234), .A2(n1257), .A3(n1067), .A4(n1258), .ZN(n1215) );
NOR2_X1 U930 ( .A1(n1259), .A2(n1064), .ZN(n1067) );
XOR2_X1 U931 ( .A(n1220), .B(n1260), .Z(G21) );
NOR2_X1 U932 ( .A1(KEYINPUT15), .A2(n1261), .ZN(n1260) );
AND3_X1 U933 ( .A1(n1257), .A2(n1240), .A3(n1212), .ZN(n1220) );
INV_X1 U934 ( .A(n1207), .ZN(n1212) );
NAND2_X1 U935 ( .A1(n1064), .A2(n1259), .ZN(n1207) );
INV_X1 U936 ( .A(n1063), .ZN(n1259) );
XOR2_X1 U937 ( .A(n1222), .B(n1262), .Z(G18) );
NOR2_X1 U938 ( .A1(G116), .A2(KEYINPUT38), .ZN(n1262) );
NAND3_X1 U939 ( .A1(n1062), .A2(n1074), .A3(n1257), .ZN(n1222) );
NAND2_X1 U940 ( .A1(n1263), .A2(n1264), .ZN(n1074) );
NAND3_X1 U941 ( .A1(n1265), .A2(n1258), .A3(n1266), .ZN(n1264) );
INV_X1 U942 ( .A(KEYINPUT9), .ZN(n1266) );
NAND2_X1 U943 ( .A1(KEYINPUT9), .A2(n1240), .ZN(n1263) );
XNOR2_X1 U944 ( .A(n1219), .B(n1267), .ZN(G15) );
NAND2_X1 U945 ( .A1(KEYINPUT27), .A2(G113), .ZN(n1267) );
AND3_X1 U946 ( .A1(n1062), .A2(n1208), .A3(n1257), .ZN(n1219) );
AND4_X1 U947 ( .A1(n1079), .A2(n1056), .A3(n1070), .A4(n1224), .ZN(n1257) );
INV_X1 U948 ( .A(n1252), .ZN(n1056) );
INV_X1 U949 ( .A(n1076), .ZN(n1208) );
NAND2_X1 U950 ( .A1(n1237), .A2(n1234), .ZN(n1076) );
INV_X1 U951 ( .A(n1249), .ZN(n1062) );
NAND2_X1 U952 ( .A1(n1268), .A2(n1064), .ZN(n1249) );
XNOR2_X1 U953 ( .A(n1063), .B(KEYINPUT19), .ZN(n1268) );
XOR2_X1 U954 ( .A(n1269), .B(n1218), .Z(G12) );
NOR3_X1 U955 ( .A1(n1064), .A2(n1063), .A3(n1250), .ZN(n1218) );
NAND3_X1 U956 ( .A1(n1205), .A2(n1224), .A3(n1240), .ZN(n1250) );
INV_X1 U957 ( .A(n1042), .ZN(n1240) );
NAND2_X1 U958 ( .A1(n1237), .A2(n1265), .ZN(n1042) );
XNOR2_X1 U959 ( .A(n1234), .B(KEYINPUT12), .ZN(n1265) );
XOR2_X1 U960 ( .A(n1084), .B(KEYINPUT8), .Z(n1234) );
XOR2_X1 U961 ( .A(n1270), .B(n1271), .Z(n1084) );
XOR2_X1 U962 ( .A(KEYINPUT36), .B(G475), .Z(n1271) );
NAND2_X1 U963 ( .A1(n1153), .A2(n1192), .ZN(n1270) );
XOR2_X1 U964 ( .A(n1272), .B(n1273), .Z(n1153) );
XOR2_X1 U965 ( .A(n1274), .B(n1275), .Z(n1273) );
NAND2_X1 U966 ( .A1(KEYINPUT58), .A2(n1276), .ZN(n1275) );
NAND2_X1 U967 ( .A1(n1277), .A2(n1278), .ZN(n1274) );
NAND2_X1 U968 ( .A1(n1279), .A2(G143), .ZN(n1278) );
XOR2_X1 U969 ( .A(KEYINPUT29), .B(n1280), .Z(n1277) );
NOR2_X1 U970 ( .A1(G143), .A2(n1281), .ZN(n1280) );
XNOR2_X1 U971 ( .A(n1279), .B(KEYINPUT37), .ZN(n1281) );
AND3_X1 U972 ( .A1(n1282), .A2(n1102), .A3(G214), .ZN(n1279) );
XNOR2_X1 U973 ( .A(G131), .B(n1283), .ZN(n1272) );
NOR2_X1 U974 ( .A1(KEYINPUT25), .A2(n1284), .ZN(n1283) );
XOR2_X1 U975 ( .A(n1285), .B(n1286), .Z(n1284) );
XOR2_X1 U976 ( .A(G113), .B(G104), .Z(n1286) );
NAND2_X1 U977 ( .A1(KEYINPUT2), .A2(G122), .ZN(n1285) );
INV_X1 U978 ( .A(n1258), .ZN(n1237) );
XOR2_X1 U979 ( .A(n1087), .B(n1287), .Z(n1258) );
XNOR2_X1 U980 ( .A(KEYINPUT30), .B(n1088), .ZN(n1287) );
INV_X1 U981 ( .A(G478), .ZN(n1088) );
NOR2_X1 U982 ( .A1(n1149), .A2(G902), .ZN(n1087) );
XOR2_X1 U983 ( .A(n1288), .B(n1289), .Z(n1149) );
XOR2_X1 U984 ( .A(n1290), .B(n1291), .Z(n1289) );
XNOR2_X1 U985 ( .A(n1292), .B(G116), .ZN(n1291) );
INV_X1 U986 ( .A(G128), .ZN(n1292) );
XOR2_X1 U987 ( .A(KEYINPUT44), .B(G134), .Z(n1290) );
XOR2_X1 U988 ( .A(n1293), .B(n1294), .Z(n1288) );
XOR2_X1 U989 ( .A(G107), .B(n1295), .Z(n1294) );
AND3_X1 U990 ( .A1(G217), .A2(n1102), .A3(G234), .ZN(n1295) );
XOR2_X1 U991 ( .A(n1296), .B(n1297), .Z(n1293) );
NOR2_X1 U992 ( .A1(KEYINPUT24), .A2(n1298), .ZN(n1297) );
NAND2_X1 U993 ( .A1(KEYINPUT0), .A2(n1299), .ZN(n1296) );
NAND2_X1 U994 ( .A1(n1038), .A2(n1300), .ZN(n1224) );
NAND3_X1 U995 ( .A1(G902), .A2(n1256), .A3(n1137), .ZN(n1300) );
NOR2_X1 U996 ( .A1(G898), .A2(n1102), .ZN(n1137) );
NAND3_X1 U997 ( .A1(n1256), .A2(n1102), .A3(G952), .ZN(n1038) );
NAND2_X1 U998 ( .A1(G237), .A2(G234), .ZN(n1256) );
NOR2_X1 U999 ( .A1(n1068), .A2(n1252), .ZN(n1205) );
NAND2_X1 U1000 ( .A1(n1057), .A2(n1058), .ZN(n1252) );
NAND2_X1 U1001 ( .A1(G214), .A2(n1301), .ZN(n1058) );
XNOR2_X1 U1002 ( .A(n1302), .B(n1191), .ZN(n1057) );
AND2_X1 U1003 ( .A1(G210), .A2(n1301), .ZN(n1191) );
NAND2_X1 U1004 ( .A1(n1303), .A2(n1192), .ZN(n1301) );
NAND2_X1 U1005 ( .A1(n1304), .A2(n1192), .ZN(n1302) );
XOR2_X1 U1006 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1007 ( .A(n1227), .B(n1190), .ZN(n1306) );
XOR2_X1 U1008 ( .A(n1307), .B(n1170), .Z(n1190) );
INV_X1 U1009 ( .A(n1173), .ZN(n1170) );
NAND2_X1 U1010 ( .A1(G224), .A2(n1102), .ZN(n1307) );
XNOR2_X1 U1011 ( .A(n1135), .B(n1308), .ZN(n1227) );
XNOR2_X1 U1012 ( .A(n1309), .B(n1132), .ZN(n1308) );
XOR2_X1 U1013 ( .A(n1310), .B(n1311), .Z(n1132) );
NAND2_X1 U1014 ( .A1(KEYINPUT61), .A2(n1298), .ZN(n1310) );
INV_X1 U1015 ( .A(G122), .ZN(n1298) );
NAND2_X1 U1016 ( .A1(KEYINPUT23), .A2(n1134), .ZN(n1309) );
NAND2_X1 U1017 ( .A1(n1312), .A2(n1313), .ZN(n1134) );
NAND2_X1 U1018 ( .A1(n1314), .A2(n1261), .ZN(n1313) );
INV_X1 U1019 ( .A(G119), .ZN(n1261) );
XOR2_X1 U1020 ( .A(KEYINPUT17), .B(n1315), .Z(n1314) );
NAND2_X1 U1021 ( .A1(n1315), .A2(G119), .ZN(n1312) );
XNOR2_X1 U1022 ( .A(KEYINPUT28), .B(n1119), .ZN(n1305) );
INV_X1 U1023 ( .A(n1236), .ZN(n1068) );
NOR2_X1 U1024 ( .A1(n1049), .A2(n1079), .ZN(n1236) );
NOR2_X1 U1025 ( .A1(n1316), .A2(n1090), .ZN(n1079) );
NOR2_X1 U1026 ( .A1(n1091), .A2(G469), .ZN(n1090) );
AND2_X1 U1027 ( .A1(G469), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1028 ( .A(KEYINPUT43), .B(n1091), .ZN(n1317) );
NAND2_X1 U1029 ( .A1(n1318), .A2(n1192), .ZN(n1091) );
XNOR2_X1 U1030 ( .A(n1111), .B(n1319), .ZN(n1318) );
XOR2_X1 U1031 ( .A(n1320), .B(n1181), .Z(n1319) );
XNOR2_X1 U1032 ( .A(n1169), .B(n1135), .ZN(n1181) );
XOR2_X1 U1033 ( .A(G101), .B(n1321), .Z(n1135) );
XOR2_X1 U1034 ( .A(G107), .B(G104), .Z(n1321) );
NAND3_X1 U1035 ( .A1(n1322), .A2(n1323), .A3(n1324), .ZN(n1320) );
NAND2_X1 U1036 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
OR3_X1 U1037 ( .A1(n1326), .A2(n1325), .A3(KEYINPUT57), .ZN(n1323) );
XOR2_X1 U1038 ( .A(G110), .B(n1327), .Z(n1325) );
NOR2_X1 U1039 ( .A1(G140), .A2(KEYINPUT16), .ZN(n1327) );
OR2_X1 U1040 ( .A1(KEYINPUT53), .A2(n1179), .ZN(n1326) );
NAND2_X1 U1041 ( .A1(KEYINPUT57), .A2(n1179), .ZN(n1322) );
NAND2_X1 U1042 ( .A1(G227), .A2(n1102), .ZN(n1179) );
XNOR2_X1 U1043 ( .A(n1328), .B(n1329), .ZN(n1111) );
NOR2_X1 U1044 ( .A1(KEYINPUT47), .A2(n1330), .ZN(n1329) );
XNOR2_X1 U1045 ( .A(G128), .B(KEYINPUT51), .ZN(n1328) );
INV_X1 U1046 ( .A(n1070), .ZN(n1049) );
NAND2_X1 U1047 ( .A1(G221), .A2(n1331), .ZN(n1070) );
NOR2_X1 U1048 ( .A1(n1332), .A2(n1089), .ZN(n1063) );
NOR2_X1 U1049 ( .A1(n1093), .A2(n1094), .ZN(n1089) );
AND2_X1 U1050 ( .A1(n1094), .A2(n1093), .ZN(n1332) );
NAND2_X1 U1051 ( .A1(G217), .A2(n1331), .ZN(n1093) );
NAND2_X1 U1052 ( .A1(G234), .A2(n1333), .ZN(n1331) );
XNOR2_X1 U1053 ( .A(KEYINPUT39), .B(n1192), .ZN(n1333) );
NOR2_X1 U1054 ( .A1(n1142), .A2(G902), .ZN(n1094) );
XNOR2_X1 U1055 ( .A(n1334), .B(n1335), .ZN(n1142) );
XOR2_X1 U1056 ( .A(n1336), .B(n1337), .Z(n1335) );
XNOR2_X1 U1057 ( .A(G110), .B(n1338), .ZN(n1337) );
AND3_X1 U1058 ( .A1(G221), .A2(n1102), .A3(G234), .ZN(n1338) );
NAND2_X1 U1059 ( .A1(KEYINPUT11), .A2(n1339), .ZN(n1336) );
XNOR2_X1 U1060 ( .A(G128), .B(n1340), .ZN(n1339) );
NAND2_X1 U1061 ( .A1(KEYINPUT26), .A2(G119), .ZN(n1340) );
XNOR2_X1 U1062 ( .A(n1341), .B(n1276), .ZN(n1334) );
XOR2_X1 U1063 ( .A(n1119), .B(n1342), .Z(n1276) );
XNOR2_X1 U1064 ( .A(n1232), .B(G140), .ZN(n1342) );
INV_X1 U1065 ( .A(G125), .ZN(n1119) );
NAND2_X1 U1066 ( .A1(KEYINPUT31), .A2(n1343), .ZN(n1341) );
XNOR2_X1 U1067 ( .A(n1344), .B(G472), .ZN(n1064) );
NAND2_X1 U1068 ( .A1(n1345), .A2(n1192), .ZN(n1344) );
INV_X1 U1069 ( .A(G902), .ZN(n1192) );
XOR2_X1 U1070 ( .A(n1346), .B(n1347), .Z(n1345) );
XNOR2_X1 U1071 ( .A(n1165), .B(n1156), .ZN(n1347) );
XNOR2_X1 U1072 ( .A(n1348), .B(n1248), .ZN(n1156) );
INV_X1 U1073 ( .A(G101), .ZN(n1248) );
NAND3_X1 U1074 ( .A1(n1282), .A2(n1102), .A3(G210), .ZN(n1348) );
INV_X1 U1075 ( .A(G953), .ZN(n1102) );
XNOR2_X1 U1076 ( .A(n1303), .B(KEYINPUT33), .ZN(n1282) );
INV_X1 U1077 ( .A(G237), .ZN(n1303) );
XOR2_X1 U1078 ( .A(G119), .B(n1315), .Z(n1165) );
XOR2_X1 U1079 ( .A(G113), .B(G116), .Z(n1315) );
XNOR2_X1 U1080 ( .A(KEYINPUT45), .B(n1349), .ZN(n1346) );
NOR2_X1 U1081 ( .A1(KEYINPUT40), .A2(n1350), .ZN(n1349) );
XNOR2_X1 U1082 ( .A(n1169), .B(n1173), .ZN(n1350) );
XOR2_X1 U1083 ( .A(n1351), .B(n1330), .Z(n1173) );
XNOR2_X1 U1084 ( .A(n1232), .B(n1299), .ZN(n1330) );
INV_X1 U1085 ( .A(G143), .ZN(n1299) );
INV_X1 U1086 ( .A(G146), .ZN(n1232) );
XNOR2_X1 U1087 ( .A(G128), .B(KEYINPUT4), .ZN(n1351) );
NAND2_X1 U1088 ( .A1(n1352), .A2(n1353), .ZN(n1169) );
OR2_X1 U1089 ( .A1(n1112), .A2(KEYINPUT32), .ZN(n1353) );
XNOR2_X1 U1090 ( .A(G131), .B(n1354), .ZN(n1112) );
NAND3_X1 U1091 ( .A1(G131), .A2(n1354), .A3(KEYINPUT32), .ZN(n1352) );
XNOR2_X1 U1092 ( .A(G134), .B(n1343), .ZN(n1354) );
INV_X1 U1093 ( .A(G137), .ZN(n1343) );
NAND2_X1 U1094 ( .A1(KEYINPUT55), .A2(n1311), .ZN(n1269) );
INV_X1 U1095 ( .A(G110), .ZN(n1311) );
endmodule


