//Key = 0011100101101011111010010001111011001001001000110000101001000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
n1424, n1425;

XNOR2_X1 U776 ( .A(G107), .B(n1084), .ZN(G9) );
NOR2_X1 U777 ( .A1(n1085), .A2(n1086), .ZN(G75) );
NOR4_X1 U778 ( .A1(n1087), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1086) );
NAND3_X1 U779 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1087) );
NAND2_X1 U780 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U781 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NAND4_X1 U782 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
NAND2_X1 U783 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
OR2_X1 U784 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U785 ( .A1(n1106), .A2(n1107), .ZN(n1096) );
NAND2_X1 U786 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U787 ( .A1(n1099), .A2(n1110), .ZN(n1109) );
NAND2_X1 U788 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND3_X1 U789 ( .A1(n1113), .A2(n1114), .A3(KEYINPUT49), .ZN(n1112) );
NAND2_X1 U790 ( .A1(n1100), .A2(n1114), .ZN(n1108) );
NAND3_X1 U791 ( .A1(n1115), .A2(n1116), .A3(n1100), .ZN(n1114) );
NAND2_X1 U792 ( .A1(n1099), .A2(n1117), .ZN(n1116) );
NAND2_X1 U793 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U794 ( .A1(n1113), .A2(n1120), .ZN(n1119) );
INV_X1 U795 ( .A(KEYINPUT49), .ZN(n1120) );
NAND2_X1 U796 ( .A1(n1098), .A2(n1121), .ZN(n1115) );
NAND2_X1 U797 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
INV_X1 U799 ( .A(n1126), .ZN(n1122) );
NOR3_X1 U800 ( .A1(n1127), .A2(G953), .A3(n1128), .ZN(n1085) );
INV_X1 U801 ( .A(n1091), .ZN(n1128) );
NAND4_X1 U802 ( .A1(n1129), .A2(n1104), .A3(n1130), .A4(n1131), .ZN(n1091) );
NOR4_X1 U803 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1131) );
XOR2_X1 U804 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U805 ( .A(n1138), .B(n1139), .Z(n1132) );
NOR3_X1 U806 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1130) );
INV_X1 U807 ( .A(n1143), .ZN(n1142) );
NAND2_X1 U808 ( .A1(n1144), .A2(n1145), .ZN(n1129) );
XOR2_X1 U809 ( .A(n1089), .B(KEYINPUT7), .Z(n1127) );
XOR2_X1 U810 ( .A(n1146), .B(n1147), .Z(G72) );
XOR2_X1 U811 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U812 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND2_X1 U813 ( .A1(G953), .A2(n1152), .ZN(n1151) );
XOR2_X1 U814 ( .A(n1153), .B(n1154), .Z(n1150) );
XOR2_X1 U815 ( .A(G125), .B(n1155), .Z(n1154) );
NOR2_X1 U816 ( .A1(KEYINPUT0), .A2(n1156), .ZN(n1155) );
XOR2_X1 U817 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U818 ( .A(G134), .B(G131), .Z(n1158) );
XOR2_X1 U819 ( .A(n1159), .B(n1160), .Z(n1157) );
NOR2_X1 U820 ( .A1(G137), .A2(KEYINPUT48), .ZN(n1160) );
NAND2_X1 U821 ( .A1(KEYINPUT12), .A2(n1161), .ZN(n1153) );
NAND3_X1 U822 ( .A1(n1090), .A2(n1092), .A3(n1162), .ZN(n1148) );
XNOR2_X1 U823 ( .A(KEYINPUT62), .B(KEYINPUT32), .ZN(n1162) );
NOR2_X1 U824 ( .A1(n1163), .A2(n1092), .ZN(n1146) );
AND2_X1 U825 ( .A1(G227), .A2(G900), .ZN(n1163) );
XOR2_X1 U826 ( .A(n1164), .B(n1165), .Z(G69) );
XOR2_X1 U827 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U828 ( .A1(n1168), .A2(n1092), .ZN(n1167) );
AND2_X1 U829 ( .A1(G224), .A2(G898), .ZN(n1168) );
NAND3_X1 U830 ( .A1(n1169), .A2(n1170), .A3(n1171), .ZN(n1166) );
XOR2_X1 U831 ( .A(n1172), .B(KEYINPUT53), .Z(n1171) );
NAND2_X1 U832 ( .A1(G953), .A2(n1173), .ZN(n1169) );
NAND2_X1 U833 ( .A1(n1092), .A2(n1088), .ZN(n1164) );
NOR2_X1 U834 ( .A1(n1174), .A2(n1175), .ZN(G66) );
XOR2_X1 U835 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U836 ( .A1(n1178), .A2(n1179), .ZN(n1176) );
NOR2_X1 U837 ( .A1(n1174), .A2(n1180), .ZN(G63) );
NOR3_X1 U838 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
NOR2_X1 U839 ( .A1(KEYINPUT15), .A2(n1184), .ZN(n1183) );
AND3_X1 U840 ( .A1(n1184), .A2(n1185), .A3(KEYINPUT15), .ZN(n1182) );
NOR2_X1 U841 ( .A1(n1185), .A2(n1186), .ZN(n1181) );
NOR2_X1 U842 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
INV_X1 U843 ( .A(KEYINPUT15), .ZN(n1188) );
XNOR2_X1 U844 ( .A(n1184), .B(KEYINPUT5), .ZN(n1187) );
XNOR2_X1 U845 ( .A(n1189), .B(KEYINPUT37), .ZN(n1184) );
NOR2_X1 U846 ( .A1(n1190), .A2(n1136), .ZN(n1185) );
NOR2_X1 U847 ( .A1(n1174), .A2(n1191), .ZN(G60) );
NOR3_X1 U848 ( .A1(n1138), .A2(n1192), .A3(n1193), .ZN(n1191) );
AND3_X1 U849 ( .A1(n1194), .A2(G475), .A3(n1178), .ZN(n1193) );
NOR2_X1 U850 ( .A1(n1195), .A2(n1194), .ZN(n1192) );
NOR2_X1 U851 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NOR2_X1 U852 ( .A1(n1090), .A2(n1088), .ZN(n1196) );
XOR2_X1 U853 ( .A(G104), .B(n1198), .Z(G6) );
NOR3_X1 U854 ( .A1(n1199), .A2(n1118), .A3(n1200), .ZN(n1198) );
XOR2_X1 U855 ( .A(KEYINPUT18), .B(n1201), .Z(n1200) );
NAND3_X1 U856 ( .A1(n1126), .A2(n1202), .A3(n1100), .ZN(n1199) );
NOR2_X1 U857 ( .A1(n1174), .A2(n1203), .ZN(G57) );
XOR2_X1 U858 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U859 ( .A(n1206), .B(n1207), .Z(n1205) );
NOR2_X1 U860 ( .A1(KEYINPUT56), .A2(n1208), .ZN(n1206) );
XOR2_X1 U861 ( .A(n1209), .B(n1210), .Z(n1204) );
XNOR2_X1 U862 ( .A(G101), .B(n1211), .ZN(n1210) );
NOR2_X1 U863 ( .A1(KEYINPUT50), .A2(n1212), .ZN(n1211) );
NAND2_X1 U864 ( .A1(n1178), .A2(G472), .ZN(n1209) );
NOR3_X1 U865 ( .A1(n1174), .A2(n1213), .A3(n1214), .ZN(G54) );
NOR2_X1 U866 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XOR2_X1 U867 ( .A(n1217), .B(KEYINPUT24), .Z(n1215) );
NOR2_X1 U868 ( .A1(n1218), .A2(n1219), .ZN(n1213) );
XOR2_X1 U869 ( .A(KEYINPUT59), .B(n1220), .Z(n1219) );
INV_X1 U870 ( .A(n1217), .ZN(n1220) );
XOR2_X1 U871 ( .A(n1221), .B(n1222), .Z(n1217) );
XOR2_X1 U872 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U873 ( .A(n1225), .B(KEYINPUT39), .Z(n1221) );
NAND2_X1 U874 ( .A1(n1178), .A2(G469), .ZN(n1225) );
INV_X1 U875 ( .A(n1216), .ZN(n1218) );
NAND3_X1 U876 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1216) );
NAND2_X1 U877 ( .A1(n1229), .A2(G140), .ZN(n1227) );
XOR2_X1 U878 ( .A(n1230), .B(n1231), .Z(n1229) );
NAND3_X1 U879 ( .A1(n1231), .A2(n1230), .A3(n1161), .ZN(n1226) );
NOR2_X1 U880 ( .A1(n1174), .A2(n1232), .ZN(G51) );
XOR2_X1 U881 ( .A(n1233), .B(n1234), .Z(n1232) );
XNOR2_X1 U882 ( .A(n1235), .B(n1236), .ZN(n1234) );
NAND2_X1 U883 ( .A1(n1178), .A2(n1144), .ZN(n1235) );
INV_X1 U884 ( .A(n1190), .ZN(n1178) );
NAND2_X1 U885 ( .A1(G902), .A2(n1237), .ZN(n1190) );
OR2_X1 U886 ( .A1(n1088), .A2(n1090), .ZN(n1237) );
NAND4_X1 U887 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1090) );
NOR4_X1 U888 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1241) );
NOR2_X1 U889 ( .A1(n1246), .A2(n1247), .ZN(n1240) );
NOR3_X1 U890 ( .A1(n1248), .A2(n1102), .A3(n1118), .ZN(n1247) );
NAND4_X1 U891 ( .A1(n1249), .A2(n1250), .A3(n1084), .A4(n1251), .ZN(n1088) );
NOR3_X1 U892 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1251) );
NOR3_X1 U893 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1252) );
NOR2_X1 U894 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
INV_X1 U895 ( .A(n1111), .ZN(n1259) );
NAND2_X1 U896 ( .A1(n1098), .A2(n1260), .ZN(n1111) );
OR2_X1 U897 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
AND2_X1 U898 ( .A1(n1100), .A2(n1263), .ZN(n1258) );
NAND4_X1 U899 ( .A1(n1100), .A2(n1113), .A3(n1264), .A4(n1202), .ZN(n1084) );
NAND2_X1 U900 ( .A1(n1265), .A2(n1266), .ZN(n1233) );
NAND2_X1 U901 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
INV_X1 U902 ( .A(n1269), .ZN(n1267) );
NAND2_X1 U903 ( .A1(n1270), .A2(n1269), .ZN(n1265) );
XOR2_X1 U904 ( .A(n1271), .B(G125), .Z(n1269) );
NAND2_X1 U905 ( .A1(KEYINPUT63), .A2(n1272), .ZN(n1271) );
XNOR2_X1 U906 ( .A(n1273), .B(n1268), .ZN(n1270) );
XNOR2_X1 U907 ( .A(KEYINPUT41), .B(KEYINPUT10), .ZN(n1273) );
AND2_X1 U908 ( .A1(n1274), .A2(G953), .ZN(n1174) );
XOR2_X1 U909 ( .A(n1089), .B(KEYINPUT6), .Z(n1274) );
INV_X1 U910 ( .A(G952), .ZN(n1089) );
XOR2_X1 U911 ( .A(n1275), .B(n1276), .Z(G48) );
XOR2_X1 U912 ( .A(KEYINPUT44), .B(G146), .Z(n1276) );
NOR3_X1 U913 ( .A1(n1248), .A2(n1277), .A3(n1118), .ZN(n1275) );
XOR2_X1 U914 ( .A(n1102), .B(KEYINPUT38), .Z(n1277) );
XOR2_X1 U915 ( .A(G143), .B(n1246), .Z(G45) );
AND4_X1 U916 ( .A1(n1278), .A2(n1262), .A3(n1279), .A4(n1264), .ZN(n1246) );
AND2_X1 U917 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U918 ( .A1(n1282), .A2(n1283), .ZN(G42) );
OR2_X1 U919 ( .A1(n1238), .A2(G140), .ZN(n1283) );
XOR2_X1 U920 ( .A(n1284), .B(KEYINPUT40), .Z(n1282) );
NAND2_X1 U921 ( .A1(G140), .A2(n1238), .ZN(n1284) );
NAND3_X1 U922 ( .A1(n1106), .A2(n1126), .A3(n1285), .ZN(n1238) );
XNOR2_X1 U923 ( .A(n1245), .B(n1286), .ZN(G39) );
NAND2_X1 U924 ( .A1(KEYINPUT2), .A2(G137), .ZN(n1286) );
AND3_X1 U925 ( .A1(n1287), .A2(n1098), .A3(n1106), .ZN(n1245) );
XOR2_X1 U926 ( .A(G134), .B(n1244), .Z(G36) );
AND2_X1 U927 ( .A1(n1288), .A2(n1113), .ZN(n1244) );
XOR2_X1 U928 ( .A(G131), .B(n1243), .Z(G33) );
AND2_X1 U929 ( .A1(n1288), .A2(n1263), .ZN(n1243) );
AND4_X1 U930 ( .A1(n1106), .A2(n1262), .A3(n1126), .A4(n1280), .ZN(n1288) );
NOR2_X1 U931 ( .A1(n1105), .A2(n1289), .ZN(n1106) );
INV_X1 U932 ( .A(n1104), .ZN(n1289) );
XOR2_X1 U933 ( .A(G128), .B(n1242), .Z(G30) );
AND3_X1 U934 ( .A1(n1113), .A2(n1201), .A3(n1287), .ZN(n1242) );
INV_X1 U935 ( .A(n1248), .ZN(n1287) );
NAND4_X1 U936 ( .A1(n1126), .A2(n1133), .A3(n1280), .A4(n1290), .ZN(n1248) );
XNOR2_X1 U937 ( .A(G101), .B(n1291), .ZN(G3) );
NAND4_X1 U938 ( .A1(n1262), .A2(n1098), .A3(n1292), .A4(n1264), .ZN(n1291) );
NOR2_X1 U939 ( .A1(KEYINPUT51), .A2(n1256), .ZN(n1292) );
NAND3_X1 U940 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(G27) );
OR2_X1 U941 ( .A1(n1239), .A2(G125), .ZN(n1295) );
NAND2_X1 U942 ( .A1(KEYINPUT8), .A2(n1296), .ZN(n1294) );
NAND2_X1 U943 ( .A1(G125), .A2(n1297), .ZN(n1296) );
XNOR2_X1 U944 ( .A(KEYINPUT61), .B(n1239), .ZN(n1297) );
NAND2_X1 U945 ( .A1(n1298), .A2(n1299), .ZN(n1293) );
INV_X1 U946 ( .A(KEYINPUT8), .ZN(n1299) );
NAND2_X1 U947 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
NAND3_X1 U948 ( .A1(KEYINPUT61), .A2(G125), .A3(n1239), .ZN(n1301) );
OR2_X1 U949 ( .A1(n1239), .A2(KEYINPUT61), .ZN(n1300) );
NAND3_X1 U950 ( .A1(n1099), .A2(n1201), .A3(n1285), .ZN(n1239) );
AND3_X1 U951 ( .A1(n1263), .A2(n1280), .A3(n1261), .ZN(n1285) );
NAND2_X1 U952 ( .A1(n1302), .A2(n1303), .ZN(n1280) );
NAND2_X1 U953 ( .A1(n1304), .A2(n1152), .ZN(n1303) );
INV_X1 U954 ( .A(G900), .ZN(n1152) );
INV_X1 U955 ( .A(n1134), .ZN(n1099) );
XNOR2_X1 U956 ( .A(G122), .B(n1249), .ZN(G24) );
NAND4_X1 U957 ( .A1(n1278), .A2(n1305), .A3(n1100), .A4(n1281), .ZN(n1249) );
NOR2_X1 U958 ( .A1(n1290), .A2(n1133), .ZN(n1100) );
XNOR2_X1 U959 ( .A(n1250), .B(n1306), .ZN(G21) );
NOR2_X1 U960 ( .A1(KEYINPUT25), .A2(n1307), .ZN(n1306) );
NAND4_X1 U961 ( .A1(n1305), .A2(n1098), .A3(n1133), .A4(n1290), .ZN(n1250) );
XOR2_X1 U962 ( .A(G116), .B(n1254), .Z(G18) );
AND3_X1 U963 ( .A1(n1305), .A2(n1113), .A3(n1262), .ZN(n1254) );
AND2_X1 U964 ( .A1(n1281), .A2(n1308), .ZN(n1113) );
INV_X1 U965 ( .A(n1309), .ZN(n1281) );
XOR2_X1 U966 ( .A(G113), .B(n1253), .Z(G15) );
AND3_X1 U967 ( .A1(n1263), .A2(n1305), .A3(n1262), .ZN(n1253) );
AND2_X1 U968 ( .A1(n1310), .A2(n1133), .ZN(n1262) );
NOR3_X1 U969 ( .A1(n1102), .A2(n1256), .A3(n1134), .ZN(n1305) );
NAND2_X1 U970 ( .A1(n1125), .A2(n1311), .ZN(n1134) );
INV_X1 U971 ( .A(n1202), .ZN(n1256) );
INV_X1 U972 ( .A(n1118), .ZN(n1263) );
NAND2_X1 U973 ( .A1(n1312), .A2(n1309), .ZN(n1118) );
XOR2_X1 U974 ( .A(n1278), .B(KEYINPUT13), .Z(n1312) );
XOR2_X1 U975 ( .A(n1313), .B(KEYINPUT30), .Z(n1278) );
XOR2_X1 U976 ( .A(n1230), .B(n1314), .Z(G12) );
NAND4_X1 U977 ( .A1(n1315), .A2(n1261), .A3(n1098), .A4(n1264), .ZN(n1314) );
INV_X1 U978 ( .A(n1255), .ZN(n1264) );
NAND2_X1 U979 ( .A1(n1126), .A2(n1201), .ZN(n1255) );
INV_X1 U980 ( .A(n1102), .ZN(n1201) );
NAND2_X1 U981 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NAND3_X1 U982 ( .A1(n1316), .A2(n1317), .A3(n1318), .ZN(n1105) );
INV_X1 U983 ( .A(n1141), .ZN(n1318) );
NOR2_X1 U984 ( .A1(n1145), .A2(n1144), .ZN(n1141) );
NAND3_X1 U985 ( .A1(n1144), .A2(n1145), .A3(n1319), .ZN(n1317) );
INV_X1 U986 ( .A(KEYINPUT55), .ZN(n1319) );
NAND2_X1 U987 ( .A1(n1320), .A2(n1321), .ZN(n1145) );
XOR2_X1 U988 ( .A(n1322), .B(n1323), .Z(n1320) );
XOR2_X1 U989 ( .A(n1268), .B(n1272), .Z(n1323) );
NAND2_X1 U990 ( .A1(G224), .A2(n1092), .ZN(n1268) );
XOR2_X1 U991 ( .A(n1236), .B(G125), .Z(n1322) );
NAND2_X1 U992 ( .A1(n1324), .A2(n1170), .ZN(n1236) );
NAND2_X1 U993 ( .A1(n1325), .A2(n1326), .ZN(n1170) );
INV_X1 U994 ( .A(n1327), .ZN(n1326) );
XOR2_X1 U995 ( .A(G122), .B(n1230), .Z(n1325) );
XOR2_X1 U996 ( .A(n1172), .B(KEYINPUT58), .Z(n1324) );
NAND2_X1 U997 ( .A1(n1327), .A2(n1328), .ZN(n1172) );
XOR2_X1 U998 ( .A(G122), .B(G110), .Z(n1328) );
XOR2_X1 U999 ( .A(n1329), .B(n1330), .Z(n1327) );
XOR2_X1 U1000 ( .A(n1331), .B(n1332), .Z(n1330) );
XOR2_X1 U1001 ( .A(G113), .B(n1307), .Z(n1329) );
INV_X1 U1002 ( .A(G119), .ZN(n1307) );
INV_X1 U1003 ( .A(n1333), .ZN(n1144) );
NAND2_X1 U1004 ( .A1(KEYINPUT55), .A2(n1333), .ZN(n1316) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1334), .ZN(n1333) );
NAND2_X1 U1006 ( .A1(G214), .A2(n1335), .ZN(n1104) );
XNOR2_X1 U1007 ( .A(KEYINPUT46), .B(n1334), .ZN(n1335) );
NAND2_X1 U1008 ( .A1(n1336), .A2(n1321), .ZN(n1334) );
XNOR2_X1 U1009 ( .A(G237), .B(KEYINPUT60), .ZN(n1336) );
NOR2_X1 U1010 ( .A1(n1125), .A2(n1124), .ZN(n1126) );
INV_X1 U1011 ( .A(n1311), .ZN(n1124) );
NAND2_X1 U1012 ( .A1(G221), .A2(n1337), .ZN(n1311) );
XOR2_X1 U1013 ( .A(n1338), .B(G469), .Z(n1125) );
NAND2_X1 U1014 ( .A1(n1339), .A2(n1321), .ZN(n1338) );
XOR2_X1 U1015 ( .A(n1223), .B(n1340), .Z(n1339) );
XOR2_X1 U1016 ( .A(n1341), .B(n1342), .Z(n1340) );
NOR3_X1 U1017 ( .A1(n1343), .A2(n1344), .A3(n1345), .ZN(n1342) );
NOR3_X1 U1018 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1345) );
INV_X1 U1019 ( .A(n1349), .ZN(n1347) );
NOR2_X1 U1020 ( .A1(n1231), .A2(n1349), .ZN(n1344) );
NAND2_X1 U1021 ( .A1(n1350), .A2(n1230), .ZN(n1349) );
XOR2_X1 U1022 ( .A(n1161), .B(KEYINPUT23), .Z(n1350) );
INV_X1 U1023 ( .A(G140), .ZN(n1161) );
INV_X1 U1024 ( .A(n1346), .ZN(n1231) );
INV_X1 U1025 ( .A(n1228), .ZN(n1343) );
NAND2_X1 U1026 ( .A1(n1348), .A2(n1346), .ZN(n1228) );
NAND2_X1 U1027 ( .A1(G227), .A2(n1092), .ZN(n1346) );
NOR2_X1 U1028 ( .A1(n1230), .A2(G140), .ZN(n1348) );
NAND2_X1 U1029 ( .A1(KEYINPUT54), .A2(n1224), .ZN(n1341) );
XNOR2_X1 U1030 ( .A(G107), .B(n1331), .ZN(n1224) );
XOR2_X1 U1031 ( .A(G104), .B(G101), .Z(n1331) );
XOR2_X1 U1032 ( .A(n1159), .B(n1351), .Z(n1223) );
NAND2_X1 U1033 ( .A1(n1352), .A2(n1353), .ZN(n1159) );
NAND2_X1 U1034 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
INV_X1 U1035 ( .A(G146), .ZN(n1355) );
XOR2_X1 U1036 ( .A(n1356), .B(n1357), .Z(n1354) );
XOR2_X1 U1037 ( .A(KEYINPUT36), .B(KEYINPUT35), .Z(n1357) );
NAND2_X1 U1038 ( .A1(n1356), .A2(G146), .ZN(n1352) );
AND2_X1 U1039 ( .A1(n1308), .A2(n1309), .ZN(n1098) );
NAND3_X1 U1040 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1309) );
OR2_X1 U1041 ( .A1(n1137), .A2(n1361), .ZN(n1360) );
NAND3_X1 U1042 ( .A1(n1361), .A2(n1137), .A3(KEYINPUT57), .ZN(n1359) );
NAND2_X1 U1043 ( .A1(n1189), .A2(n1321), .ZN(n1137) );
XOR2_X1 U1044 ( .A(n1362), .B(n1363), .Z(n1189) );
XNOR2_X1 U1045 ( .A(n1364), .B(n1332), .ZN(n1363) );
XOR2_X1 U1046 ( .A(G107), .B(G116), .Z(n1332) );
NAND2_X1 U1047 ( .A1(n1365), .A2(KEYINPUT20), .ZN(n1364) );
XNOR2_X1 U1048 ( .A(G134), .B(n1356), .ZN(n1365) );
XOR2_X1 U1049 ( .A(G128), .B(G143), .Z(n1356) );
XOR2_X1 U1050 ( .A(n1366), .B(G122), .Z(n1362) );
NAND2_X1 U1051 ( .A1(n1367), .A2(G217), .ZN(n1366) );
AND2_X1 U1052 ( .A1(KEYINPUT29), .A2(n1136), .ZN(n1361) );
OR2_X1 U1053 ( .A1(n1136), .A2(KEYINPUT57), .ZN(n1358) );
INV_X1 U1054 ( .A(G478), .ZN(n1136) );
XNOR2_X1 U1055 ( .A(n1313), .B(KEYINPUT47), .ZN(n1308) );
NAND3_X1 U1056 ( .A1(n1368), .A2(n1369), .A3(n1370), .ZN(n1313) );
NAND2_X1 U1057 ( .A1(n1139), .A2(n1371), .ZN(n1370) );
OR3_X1 U1058 ( .A1(n1371), .A2(n1139), .A3(KEYINPUT19), .ZN(n1369) );
XOR2_X1 U1059 ( .A(n1197), .B(KEYINPUT16), .Z(n1139) );
INV_X1 U1060 ( .A(G475), .ZN(n1197) );
NAND2_X1 U1061 ( .A1(KEYINPUT52), .A2(n1372), .ZN(n1371) );
INV_X1 U1062 ( .A(n1138), .ZN(n1372) );
NAND2_X1 U1063 ( .A1(n1138), .A2(KEYINPUT19), .ZN(n1368) );
NOR2_X1 U1064 ( .A1(n1194), .A2(G902), .ZN(n1138) );
XNOR2_X1 U1065 ( .A(n1373), .B(n1374), .ZN(n1194) );
NOR2_X1 U1066 ( .A1(n1375), .A2(n1376), .ZN(n1374) );
XOR2_X1 U1067 ( .A(KEYINPUT45), .B(n1377), .Z(n1376) );
AND2_X1 U1068 ( .A1(n1378), .A2(G122), .ZN(n1377) );
NOR2_X1 U1069 ( .A1(G122), .A2(n1378), .ZN(n1375) );
XOR2_X1 U1070 ( .A(G113), .B(KEYINPUT27), .Z(n1378) );
XNOR2_X1 U1071 ( .A(G104), .B(n1379), .ZN(n1373) );
NOR2_X1 U1072 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
XOR2_X1 U1073 ( .A(n1382), .B(KEYINPUT42), .Z(n1381) );
NAND2_X1 U1074 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
NOR2_X1 U1075 ( .A1(n1384), .A2(n1383), .ZN(n1380) );
XOR2_X1 U1076 ( .A(n1385), .B(n1386), .Z(n1383) );
XOR2_X1 U1077 ( .A(n1387), .B(G143), .Z(n1386) );
NAND2_X1 U1078 ( .A1(G214), .A2(n1388), .ZN(n1387) );
NAND2_X1 U1079 ( .A1(KEYINPUT4), .A2(G131), .ZN(n1385) );
INV_X1 U1080 ( .A(n1389), .ZN(n1384) );
NOR2_X1 U1081 ( .A1(n1133), .A2(n1310), .ZN(n1261) );
INV_X1 U1082 ( .A(n1290), .ZN(n1310) );
NAND2_X1 U1083 ( .A1(n1390), .A2(n1143), .ZN(n1290) );
NAND3_X1 U1084 ( .A1(n1391), .A2(n1321), .A3(n1177), .ZN(n1143) );
XOR2_X1 U1085 ( .A(KEYINPUT33), .B(n1140), .Z(n1390) );
AND2_X1 U1086 ( .A1(n1179), .A2(n1392), .ZN(n1140) );
NAND2_X1 U1087 ( .A1(n1177), .A2(n1321), .ZN(n1392) );
XOR2_X1 U1088 ( .A(n1393), .B(n1394), .Z(n1177) );
AND2_X1 U1089 ( .A1(n1367), .A2(G221), .ZN(n1394) );
AND2_X1 U1090 ( .A1(G234), .A2(n1092), .ZN(n1367) );
XOR2_X1 U1091 ( .A(n1395), .B(G137), .Z(n1393) );
NAND2_X1 U1092 ( .A1(n1396), .A2(n1397), .ZN(n1395) );
NAND2_X1 U1093 ( .A1(n1389), .A2(n1398), .ZN(n1397) );
XOR2_X1 U1094 ( .A(n1399), .B(KEYINPUT11), .Z(n1396) );
OR2_X1 U1095 ( .A1(n1398), .A2(n1389), .ZN(n1399) );
XNOR2_X1 U1096 ( .A(G125), .B(n1400), .ZN(n1389) );
XOR2_X1 U1097 ( .A(G146), .B(G140), .Z(n1400) );
XNOR2_X1 U1098 ( .A(n1230), .B(n1401), .ZN(n1398) );
XOR2_X1 U1099 ( .A(G128), .B(G119), .Z(n1401) );
INV_X1 U1100 ( .A(n1391), .ZN(n1179) );
NAND2_X1 U1101 ( .A1(G217), .A2(n1337), .ZN(n1391) );
NAND2_X1 U1102 ( .A1(G234), .A2(n1321), .ZN(n1337) );
XNOR2_X1 U1103 ( .A(n1402), .B(n1403), .ZN(n1133) );
XOR2_X1 U1104 ( .A(KEYINPUT22), .B(G472), .Z(n1403) );
NAND2_X1 U1105 ( .A1(n1404), .A2(n1321), .ZN(n1402) );
INV_X1 U1106 ( .A(G902), .ZN(n1321) );
XOR2_X1 U1107 ( .A(n1405), .B(n1406), .Z(n1404) );
XNOR2_X1 U1108 ( .A(n1407), .B(n1212), .ZN(n1406) );
XOR2_X1 U1109 ( .A(n1408), .B(n1409), .Z(n1212) );
XOR2_X1 U1110 ( .A(KEYINPUT9), .B(G119), .Z(n1409) );
XOR2_X1 U1111 ( .A(n1410), .B(G116), .Z(n1408) );
NAND2_X1 U1112 ( .A1(KEYINPUT14), .A2(G113), .ZN(n1410) );
NOR2_X1 U1113 ( .A1(KEYINPUT26), .A2(n1207), .ZN(n1407) );
XNOR2_X1 U1114 ( .A(n1272), .B(n1351), .ZN(n1207) );
AND2_X1 U1115 ( .A1(n1411), .A2(n1412), .ZN(n1351) );
NAND2_X1 U1116 ( .A1(G131), .A2(n1413), .ZN(n1412) );
XOR2_X1 U1117 ( .A(n1414), .B(KEYINPUT1), .Z(n1411) );
OR2_X1 U1118 ( .A1(n1413), .A2(G131), .ZN(n1414) );
NAND2_X1 U1119 ( .A1(n1415), .A2(n1416), .ZN(n1413) );
NAND2_X1 U1120 ( .A1(G134), .A2(n1417), .ZN(n1416) );
XOR2_X1 U1121 ( .A(KEYINPUT17), .B(n1418), .Z(n1415) );
NOR2_X1 U1122 ( .A1(G134), .A2(n1417), .ZN(n1418) );
INV_X1 U1123 ( .A(G137), .ZN(n1417) );
XOR2_X1 U1124 ( .A(n1419), .B(n1420), .Z(n1272) );
XOR2_X1 U1125 ( .A(G146), .B(G128), .Z(n1420) );
NAND2_X1 U1126 ( .A1(KEYINPUT28), .A2(G143), .ZN(n1419) );
XNOR2_X1 U1127 ( .A(KEYINPUT21), .B(n1421), .ZN(n1405) );
NOR2_X1 U1128 ( .A1(KEYINPUT43), .A2(n1422), .ZN(n1421) );
XOR2_X1 U1129 ( .A(n1208), .B(n1423), .Z(n1422) );
XNOR2_X1 U1130 ( .A(G101), .B(KEYINPUT31), .ZN(n1423) );
NAND2_X1 U1131 ( .A1(G210), .A2(n1388), .ZN(n1208) );
NOR2_X1 U1132 ( .A1(G953), .A2(G237), .ZN(n1388) );
XOR2_X1 U1133 ( .A(n1202), .B(KEYINPUT34), .Z(n1315) );
NAND2_X1 U1134 ( .A1(n1302), .A2(n1424), .ZN(n1202) );
NAND2_X1 U1135 ( .A1(n1304), .A2(n1173), .ZN(n1424) );
INV_X1 U1136 ( .A(G898), .ZN(n1173) );
AND3_X1 U1137 ( .A1(G902), .A2(n1095), .A3(G953), .ZN(n1304) );
NAND3_X1 U1138 ( .A1(n1425), .A2(n1092), .A3(G952), .ZN(n1302) );
INV_X1 U1139 ( .A(G953), .ZN(n1092) );
XNOR2_X1 U1140 ( .A(KEYINPUT3), .B(n1095), .ZN(n1425) );
NAND2_X1 U1141 ( .A1(G237), .A2(G234), .ZN(n1095) );
INV_X1 U1142 ( .A(G110), .ZN(n1230) );
endmodule


