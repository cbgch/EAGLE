//Key = 0010111110010010100101110101011101101100011001100101000010110001


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
n2171, n2172, n2173, n2174, n2175, n2176;

NOR4_X2 U1227 ( .A1(n1773), .A2(n2093), .A3(n2089), .A4(AVERAGE), .ZN(n1897));
XOR2_X2 U1228 ( .A(RESTART), .B(KEYINPUT37), .Z(n1924) );
INV_X2 U1229 ( .A(n1812), .ZN(n1776) );
INV_X2 U1230 ( .A(U280), .ZN(n1779) );
NAND2_X1 U1231 ( .A1(n1641), .A2(n1642), .ZN(U344) );
NAND2_X1 U1232 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1643), .ZN(n1642) );
NAND2_X1 U1233 ( .A1(n1644), .A2(DATA_IN_7_), .ZN(n1641) );
NAND2_X1 U1234 ( .A1(n1645), .A2(n1646), .ZN(U343) );
NAND2_X1 U1235 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1643), .ZN(n1646) );
NAND2_X1 U1236 ( .A1(n1644), .A2(DATA_IN_6_), .ZN(n1645) );
NAND2_X1 U1237 ( .A1(n1647), .A2(n1648), .ZN(U342) );
NAND2_X1 U1238 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1643), .ZN(n1648) );
NAND2_X1 U1239 ( .A1(n1644), .A2(DATA_IN_5_), .ZN(n1647) );
NAND2_X1 U1240 ( .A1(n1649), .A2(n1650), .ZN(U341) );
NAND2_X1 U1241 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1643), .ZN(n1650) );
NAND2_X1 U1242 ( .A1(n1644), .A2(DATA_IN_4_), .ZN(n1649) );
NAND2_X1 U1243 ( .A1(n1651), .A2(n1652), .ZN(U340) );
NAND2_X1 U1244 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1643), .ZN(n1652) );
NAND2_X1 U1245 ( .A1(n1644), .A2(DATA_IN_3_), .ZN(n1651) );
NAND2_X1 U1246 ( .A1(n1653), .A2(n1654), .ZN(U339) );
NAND2_X1 U1247 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1643), .ZN(n1654) );
NAND2_X1 U1248 ( .A1(n1644), .A2(DATA_IN_2_), .ZN(n1653) );
NAND2_X1 U1249 ( .A1(n1655), .A2(n1656), .ZN(U338) );
NAND2_X1 U1250 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1643), .ZN(n1656) );
NAND2_X1 U1251 ( .A1(n1644), .A2(DATA_IN_1_), .ZN(n1655) );
NAND2_X1 U1252 ( .A1(n1657), .A2(n1658), .ZN(U337) );
NAND2_X1 U1253 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1643), .ZN(n1658) );
NAND2_X1 U1254 ( .A1(n1644), .A2(DATA_IN_0_), .ZN(n1657) );
INV_X1 U1255 ( .A(n1643), .ZN(n1644) );
NAND2_X1 U1256 ( .A1(n1659), .A2(n1660), .ZN(n1643) );
NAND3_X1 U1257 ( .A1(n1661), .A2(n1662), .A3(n1663), .ZN(n1660) );
NAND2_X1 U1258 ( .A1(n1664), .A2(n1665), .ZN(U336) );
NAND2_X1 U1259 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1666), .ZN(n1665) );
XNOR2_X1 U1260 ( .A(KEYINPUT34), .B(n1667), .ZN(n1666) );
NAND2_X1 U1261 ( .A1(n1668), .A2(DATA_IN_7_), .ZN(n1664) );
NAND2_X1 U1262 ( .A1(n1669), .A2(n1670), .ZN(U335) );
NAND2_X1 U1263 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1667), .ZN(n1670) );
NAND2_X1 U1264 ( .A1(n1668), .A2(DATA_IN_6_), .ZN(n1669) );
NAND2_X1 U1265 ( .A1(n1671), .A2(n1672), .ZN(U334) );
NAND2_X1 U1266 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1667), .ZN(n1672) );
NAND2_X1 U1267 ( .A1(n1668), .A2(DATA_IN_5_), .ZN(n1671) );
NAND2_X1 U1268 ( .A1(n1673), .A2(n1674), .ZN(U333) );
NAND2_X1 U1269 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1667), .ZN(n1674) );
NAND2_X1 U1270 ( .A1(n1668), .A2(DATA_IN_4_), .ZN(n1673) );
NAND2_X1 U1271 ( .A1(n1675), .A2(n1676), .ZN(U332) );
NAND2_X1 U1272 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1667), .ZN(n1676) );
NAND2_X1 U1273 ( .A1(n1668), .A2(DATA_IN_3_), .ZN(n1675) );
NAND2_X1 U1274 ( .A1(n1677), .A2(n1678), .ZN(U331) );
NAND2_X1 U1275 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1667), .ZN(n1678) );
NAND2_X1 U1276 ( .A1(n1668), .A2(DATA_IN_2_), .ZN(n1677) );
NAND2_X1 U1277 ( .A1(n1679), .A2(n1680), .ZN(U330) );
NAND2_X1 U1278 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1667), .ZN(n1680) );
NAND2_X1 U1279 ( .A1(n1668), .A2(DATA_IN_1_), .ZN(n1679) );
NAND2_X1 U1280 ( .A1(n1681), .A2(n1682), .ZN(U329) );
NAND2_X1 U1281 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1667), .ZN(n1682) );
NAND2_X1 U1282 ( .A1(n1668), .A2(DATA_IN_0_), .ZN(n1681) );
INV_X1 U1283 ( .A(n1667), .ZN(n1668) );
NAND2_X1 U1284 ( .A1(n1659), .A2(n1683), .ZN(n1667) );
NAND2_X1 U1285 ( .A1(n1684), .A2(n1662), .ZN(n1683) );
NAND3_X1 U1286 ( .A1(n1663), .A2(n1661), .A3(n1685), .ZN(n1684) );
NAND2_X1 U1287 ( .A1(n1686), .A2(n1687), .ZN(n1685) );
NAND3_X1 U1288 ( .A1(n1688), .A2(n1689), .A3(n1690), .ZN(n1687) );
NAND2_X1 U1289 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1691), .ZN(n1690) );
NAND3_X1 U1290 ( .A1(n1692), .A2(n1693), .A3(n1694), .ZN(n1689) );
NAND2_X1 U1291 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1695), .ZN(n1694) );
NAND3_X1 U1292 ( .A1(n1696), .A2(n1697), .A3(n1698), .ZN(n1693) );
OR2_X1 U1293 ( .A1(n1699), .A2(RMIN_REG_4__SCAN_IN), .ZN(n1698) );
NAND3_X1 U1294 ( .A1(n1700), .A2(n1701), .A3(n1702), .ZN(n1697) );
XOR2_X1 U1295 ( .A(n1703), .B(KEYINPUT20), .Z(n1702) );
NAND2_X1 U1296 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1699), .ZN(n1703) );
NAND3_X1 U1297 ( .A1(n1704), .A2(n1705), .A3(n1706), .ZN(n1701) );
NAND2_X1 U1298 ( .A1(DATA_IN_3_), .A2(n1707), .ZN(n1706) );
NAND3_X1 U1299 ( .A1(n1708), .A2(n1709), .A3(n1710), .ZN(n1705) );
NAND2_X1 U1300 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1711), .ZN(n1710) );
NAND3_X1 U1301 ( .A1(n1712), .A2(n1713), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1709) );
NAND2_X1 U1302 ( .A1(n1714), .A2(DATA_IN_1_), .ZN(n1712) );
XNOR2_X1 U1303 ( .A(RMIN_REG_1__SCAN_IN), .B(KEYINPUT13), .ZN(n1714) );
NAND2_X1 U1304 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1715), .ZN(n1708) );
NAND2_X1 U1305 ( .A1(DATA_IN_2_), .A2(n1716), .ZN(n1704) );
NAND2_X1 U1306 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1717), .ZN(n1700) );
NAND2_X1 U1307 ( .A1(DATA_IN_5_), .A2(n1718), .ZN(n1696) );
XOR2_X1 U1308 ( .A(KEYINPUT16), .B(n1719), .Z(n1718) );
XOR2_X1 U1309 ( .A(RMIN_REG_5__SCAN_IN), .B(KEYINPUT39), .Z(n1719) );
NAND2_X1 U1310 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1720), .ZN(n1692) );
NAND2_X1 U1311 ( .A1(DATA_IN_6_), .A2(n1721), .ZN(n1688) );
NAND2_X1 U1312 ( .A1(DATA_IN_7_), .A2(n1722), .ZN(n1686) );
NAND3_X1 U1313 ( .A1(n1723), .A2(n1724), .A3(n1725), .ZN(n1661) );
NAND2_X1 U1314 ( .A1(n1726), .A2(n1727), .ZN(n1725) );
XNOR2_X1 U1315 ( .A(DATA_IN_7_), .B(KEYINPUT29), .ZN(n1726) );
NAND3_X1 U1316 ( .A1(n1728), .A2(n1729), .A3(n1730), .ZN(n1724) );
OR2_X1 U1317 ( .A1(n1720), .A2(RMAX_REG_5__SCAN_IN), .ZN(n1730) );
NAND3_X1 U1318 ( .A1(n1731), .A2(n1732), .A3(n1733), .ZN(n1729) );
NAND2_X1 U1319 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1720), .ZN(n1733) );
INV_X1 U1320 ( .A(DATA_IN_5_), .ZN(n1720) );
NAND3_X1 U1321 ( .A1(n1734), .A2(n1735), .A3(n1736), .ZN(n1732) );
OR2_X1 U1322 ( .A1(n1699), .A2(RMAX_REG_4__SCAN_IN), .ZN(n1736) );
NAND3_X1 U1323 ( .A1(n1737), .A2(n1738), .A3(n1739), .ZN(n1735) );
XOR2_X1 U1324 ( .A(n1740), .B(KEYINPUT26), .Z(n1739) );
NAND2_X1 U1325 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1711), .ZN(n1740) );
NAND3_X1 U1326 ( .A1(n1741), .A2(n1742), .A3(n1743), .ZN(n1738) );
NAND2_X1 U1327 ( .A1(DATA_IN_2_), .A2(n1744), .ZN(n1743) );
NAND3_X1 U1328 ( .A1(n1745), .A2(n1746), .A3(DATA_IN_0_), .ZN(n1742) );
NAND2_X1 U1329 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1715), .ZN(n1745) );
NAND2_X1 U1330 ( .A1(DATA_IN_1_), .A2(n1747), .ZN(n1741) );
XOR2_X1 U1331 ( .A(RMAX_REG_1__SCAN_IN), .B(KEYINPUT5), .Z(n1747) );
NAND2_X1 U1332 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1717), .ZN(n1737) );
INV_X1 U1333 ( .A(DATA_IN_3_), .ZN(n1717) );
NAND2_X1 U1334 ( .A1(DATA_IN_3_), .A2(n1748), .ZN(n1734) );
NAND2_X1 U1335 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1699), .ZN(n1731) );
NAND2_X1 U1336 ( .A1(n1749), .A2(DATA_IN_6_), .ZN(n1728) );
XNOR2_X1 U1337 ( .A(RMAX_REG_6__SCAN_IN), .B(KEYINPUT0), .ZN(n1749) );
NAND2_X1 U1338 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1750), .ZN(n1723) );
XNOR2_X1 U1339 ( .A(KEYINPUT14), .B(n1695), .ZN(n1750) );
NAND2_X1 U1340 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1691), .ZN(n1663) );
NAND2_X1 U1341 ( .A1(n1751), .A2(n1752), .ZN(U328) );
NAND2_X1 U1342 ( .A1(n1753), .A2(DATA_IN_7_), .ZN(n1752) );
XOR2_X1 U1343 ( .A(KEYINPUT51), .B(n1754), .Z(n1751) );
AND2_X1 U1344 ( .A1(n1755), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1754) );
NAND2_X1 U1345 ( .A1(n1756), .A2(n1757), .ZN(U327) );
NAND2_X1 U1346 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1755), .ZN(n1757) );
NAND2_X1 U1347 ( .A1(n1753), .A2(DATA_IN_6_), .ZN(n1756) );
NAND2_X1 U1348 ( .A1(n1758), .A2(n1759), .ZN(U326) );
NAND2_X1 U1349 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1755), .ZN(n1759) );
NAND2_X1 U1350 ( .A1(n1753), .A2(DATA_IN_5_), .ZN(n1758) );
NAND2_X1 U1351 ( .A1(n1760), .A2(n1761), .ZN(U325) );
NAND2_X1 U1352 ( .A1(n1762), .A2(n1755), .ZN(n1761) );
XNOR2_X1 U1353 ( .A(RLAST_REG_4__SCAN_IN), .B(KEYINPUT36), .ZN(n1762) );
NAND2_X1 U1354 ( .A1(n1753), .A2(DATA_IN_4_), .ZN(n1760) );
NAND2_X1 U1355 ( .A1(n1763), .A2(n1764), .ZN(U324) );
NAND2_X1 U1356 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1755), .ZN(n1764) );
NAND2_X1 U1357 ( .A1(n1753), .A2(DATA_IN_3_), .ZN(n1763) );
NAND2_X1 U1358 ( .A1(n1765), .A2(n1766), .ZN(U323) );
NAND2_X1 U1359 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1755), .ZN(n1766) );
NAND2_X1 U1360 ( .A1(n1753), .A2(DATA_IN_2_), .ZN(n1765) );
NAND2_X1 U1361 ( .A1(n1767), .A2(n1768), .ZN(U322) );
NAND2_X1 U1362 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1755), .ZN(n1768) );
NAND2_X1 U1363 ( .A1(n1753), .A2(DATA_IN_1_), .ZN(n1767) );
NAND2_X1 U1364 ( .A1(n1769), .A2(n1770), .ZN(U321) );
NAND2_X1 U1365 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1771), .ZN(n1770) );
XNOR2_X1 U1366 ( .A(KEYINPUT6), .B(n1755), .ZN(n1771) );
NAND2_X1 U1367 ( .A1(n1659), .A2(n1772), .ZN(n1755) );
INV_X1 U1368 ( .A(U375), .ZN(n1659) );
NOR2_X1 U1369 ( .A1(STATO_REG_0__SCAN_IN), .A2(STATO_REG_1__SCAN_IN), .ZN(U375) );
NAND2_X1 U1370 ( .A1(n1753), .A2(DATA_IN_0_), .ZN(n1769) );
AND2_X1 U1371 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1772), .ZN(n1753) );
NAND2_X1 U1372 ( .A1(n1662), .A2(n1773), .ZN(n1772) );
NAND2_X1 U1373 ( .A1(n1774), .A2(n1775), .ZN(U320) );
NAND2_X1 U1374 ( .A1(n1776), .A2(DATA_IN_7_), .ZN(n1775) );
XOR2_X1 U1375 ( .A(n1777), .B(KEYINPUT60), .Z(n1774) );
NAND2_X1 U1376 ( .A1(n1778), .A2(n1779), .ZN(n1777) );
XOR2_X1 U1377 ( .A(REG1_REG_7__SCAN_IN), .B(KEYINPUT50), .Z(n1778) );
NAND2_X1 U1378 ( .A1(n1780), .A2(n1781), .ZN(U319) );
NAND2_X1 U1379 ( .A1(n1776), .A2(n1782), .ZN(n1781) );
XNOR2_X1 U1380 ( .A(KEYINPUT43), .B(n1695), .ZN(n1782) );
NAND2_X1 U1381 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1779), .ZN(n1780) );
NAND2_X1 U1382 ( .A1(n1783), .A2(n1784), .ZN(U318) );
NAND2_X1 U1383 ( .A1(n1776), .A2(DATA_IN_5_), .ZN(n1784) );
NAND2_X1 U1384 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1779), .ZN(n1783) );
NAND2_X1 U1385 ( .A1(n1785), .A2(n1786), .ZN(U317) );
NAND2_X1 U1386 ( .A1(n1776), .A2(DATA_IN_4_), .ZN(n1786) );
NAND2_X1 U1387 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1779), .ZN(n1785) );
NAND2_X1 U1388 ( .A1(n1787), .A2(n1788), .ZN(U316) );
NAND2_X1 U1389 ( .A1(n1776), .A2(DATA_IN_3_), .ZN(n1788) );
NAND2_X1 U1390 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1779), .ZN(n1787) );
NAND2_X1 U1391 ( .A1(n1789), .A2(n1790), .ZN(U315) );
NAND2_X1 U1392 ( .A1(n1791), .A2(n1776), .ZN(n1790) );
XNOR2_X1 U1393 ( .A(DATA_IN_2_), .B(KEYINPUT25), .ZN(n1791) );
NAND2_X1 U1394 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1779), .ZN(n1789) );
NAND2_X1 U1395 ( .A1(n1792), .A2(n1793), .ZN(U314) );
NAND2_X1 U1396 ( .A1(n1776), .A2(DATA_IN_1_), .ZN(n1793) );
NAND2_X1 U1397 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1779), .ZN(n1792) );
NAND2_X1 U1398 ( .A1(n1794), .A2(n1795), .ZN(U313) );
NAND2_X1 U1399 ( .A1(n1776), .A2(DATA_IN_0_), .ZN(n1795) );
NAND2_X1 U1400 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1779), .ZN(n1794) );
NAND2_X1 U1401 ( .A1(n1796), .A2(n1797), .ZN(U312) );
NAND2_X1 U1402 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1776), .ZN(n1797) );
NAND2_X1 U1403 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1779), .ZN(n1796) );
NAND2_X1 U1404 ( .A1(n1798), .A2(n1799), .ZN(U311) );
NAND2_X1 U1405 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1776), .ZN(n1799) );
NAND2_X1 U1406 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1779), .ZN(n1798) );
NAND2_X1 U1407 ( .A1(n1800), .A2(n1801), .ZN(U310) );
NAND2_X1 U1408 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1779), .ZN(n1801) );
XOR2_X1 U1409 ( .A(n1802), .B(KEYINPUT12), .Z(n1800) );
NAND2_X1 U1410 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1776), .ZN(n1802) );
NAND2_X1 U1411 ( .A1(n1803), .A2(n1804), .ZN(U309) );
NAND2_X1 U1412 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1776), .ZN(n1804) );
NAND2_X1 U1413 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1779), .ZN(n1803) );
NAND2_X1 U1414 ( .A1(n1805), .A2(n1806), .ZN(U308) );
NAND2_X1 U1415 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1776), .ZN(n1806) );
NAND2_X1 U1416 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1779), .ZN(n1805) );
NAND2_X1 U1417 ( .A1(n1807), .A2(n1808), .ZN(U307) );
NAND2_X1 U1418 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1776), .ZN(n1808) );
NAND2_X1 U1419 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1779), .ZN(n1807) );
NAND2_X1 U1420 ( .A1(n1809), .A2(n1810), .ZN(U306) );
NAND2_X1 U1421 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1811), .ZN(n1810) );
XNOR2_X1 U1422 ( .A(KEYINPUT17), .B(n1812), .ZN(n1811) );
NAND2_X1 U1423 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1779), .ZN(n1809) );
NAND2_X1 U1424 ( .A1(n1813), .A2(n1814), .ZN(U305) );
NAND2_X1 U1425 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1776), .ZN(n1814) );
NAND2_X1 U1426 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1779), .ZN(n1813) );
NAND2_X1 U1427 ( .A1(n1815), .A2(n1816), .ZN(U304) );
NAND2_X1 U1428 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1776), .ZN(n1816) );
NAND2_X1 U1429 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1779), .ZN(n1815) );
NAND2_X1 U1430 ( .A1(n1817), .A2(n1818), .ZN(U303) );
NAND2_X1 U1431 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1776), .ZN(n1818) );
NAND2_X1 U1432 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1779), .ZN(n1817) );
NAND2_X1 U1433 ( .A1(n1819), .A2(n1820), .ZN(U302) );
NAND2_X1 U1434 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1776), .ZN(n1820) );
NAND2_X1 U1435 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1779), .ZN(n1819) );
NAND2_X1 U1436 ( .A1(n1821), .A2(n1822), .ZN(U301) );
NAND2_X1 U1437 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1776), .ZN(n1822) );
NAND2_X1 U1438 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1779), .ZN(n1821) );
NAND2_X1 U1439 ( .A1(n1823), .A2(n1824), .ZN(U300) );
NAND2_X1 U1440 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1776), .ZN(n1824) );
NAND2_X1 U1441 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1779), .ZN(n1823) );
NAND2_X1 U1442 ( .A1(n1825), .A2(n1826), .ZN(U299) );
NAND2_X1 U1443 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1776), .ZN(n1826) );
NAND2_X1 U1444 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1779), .ZN(n1825) );
NAND2_X1 U1445 ( .A1(n1827), .A2(n1828), .ZN(U298) );
NAND2_X1 U1446 ( .A1(n1829), .A2(REG2_REG_1__SCAN_IN), .ZN(n1828) );
XNOR2_X1 U1447 ( .A(n1776), .B(KEYINPUT41), .ZN(n1829) );
NAND2_X1 U1448 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1779), .ZN(n1827) );
NAND2_X1 U1449 ( .A1(n1830), .A2(n1831), .ZN(U297) );
NAND2_X1 U1450 ( .A1(n1832), .A2(REG2_REG_0__SCAN_IN), .ZN(n1831) );
XNOR2_X1 U1451 ( .A(n1776), .B(KEYINPUT63), .ZN(n1832) );
NAND2_X1 U1452 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1779), .ZN(n1830) );
NAND2_X1 U1453 ( .A1(n1833), .A2(n1834), .ZN(U296) );
NAND2_X1 U1454 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1776), .ZN(n1834) );
NAND2_X1 U1455 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1779), .ZN(n1833) );
NAND2_X1 U1456 ( .A1(n1835), .A2(n1836), .ZN(U295) );
NAND2_X1 U1457 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1776), .ZN(n1836) );
NAND2_X1 U1458 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1779), .ZN(n1835) );
NAND2_X1 U1459 ( .A1(n1837), .A2(n1838), .ZN(U294) );
NAND2_X1 U1460 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1776), .ZN(n1838) );
NAND2_X1 U1461 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1779), .ZN(n1837) );
NAND2_X1 U1462 ( .A1(n1839), .A2(n1840), .ZN(U293) );
NAND2_X1 U1463 ( .A1(n1841), .A2(n1779), .ZN(n1840) );
XOR2_X1 U1464 ( .A(REG4_REG_4__SCAN_IN), .B(KEYINPUT18), .Z(n1841) );
NAND2_X1 U1465 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1776), .ZN(n1839) );
NAND2_X1 U1466 ( .A1(n1842), .A2(n1843), .ZN(U292) );
NAND2_X1 U1467 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1844), .ZN(n1843) );
XNOR2_X1 U1468 ( .A(KEYINPUT47), .B(U280), .ZN(n1844) );
NAND2_X1 U1469 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1776), .ZN(n1842) );
NAND2_X1 U1470 ( .A1(n1845), .A2(n1846), .ZN(U291) );
NAND2_X1 U1471 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1776), .ZN(n1846) );
NAND2_X1 U1472 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1779), .ZN(n1845) );
NAND2_X1 U1473 ( .A1(n1847), .A2(n1848), .ZN(U290) );
NAND2_X1 U1474 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1776), .ZN(n1848) );
NAND2_X1 U1475 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1779), .ZN(n1847) );
NAND2_X1 U1476 ( .A1(n1849), .A2(n1850), .ZN(U289) );
NAND2_X1 U1477 ( .A1(n1851), .A2(n1776), .ZN(n1850) );
XNOR2_X1 U1478 ( .A(REG3_REG_0__SCAN_IN), .B(KEYINPUT58), .ZN(n1851) );
NAND2_X1 U1479 ( .A1(n1852), .A2(REG4_REG_0__SCAN_IN), .ZN(n1849) );
XNOR2_X1 U1480 ( .A(n1779), .B(KEYINPUT8), .ZN(n1852) );
NAND4_X1 U1481 ( .A1(n1853), .A2(n1854), .A3(n1855), .A4(n1856), .ZN(U288));
NAND2_X1 U1482 ( .A1(n1857), .A2(REG4_REG_7__SCAN_IN), .ZN(n1856) );
NAND2_X1 U1483 ( .A1(n1858), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1855) );
NAND2_X1 U1484 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1779), .ZN(n1854) );
INV_X1 U1485 ( .A(n1859), .ZN(n1853) );
NAND4_X1 U1486 ( .A1(n1860), .A2(n1861), .A3(n1862), .A4(n1863), .ZN(U287));
NOR4_X1 U1487 ( .A1(n1864), .A2(n1865), .A3(n1866), .A4(n1859), .ZN(n1863));
NAND2_X1 U1488 ( .A1(n1867), .A2(n1868), .ZN(n1859) );
NAND3_X1 U1489 ( .A1(n1869), .A2(n1870), .A3(n1871), .ZN(n1868) );
OR2_X1 U1490 ( .A1(n1872), .A2(n1873), .ZN(n1867) );
AND2_X1 U1491 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1779), .ZN(n1866) );
NOR2_X1 U1492 ( .A1(n1873), .A2(n1874), .ZN(n1865) );
INV_X1 U1493 ( .A(KEYINPUT28), .ZN(n1874) );
NOR4_X1 U1494 ( .A1(KEYINPUT28), .A2(n1875), .A3(n1876), .A4(n1877), .ZN(n1864) );
NAND2_X1 U1495 ( .A1(n1858), .A2(RLAST_REG_6__SCAN_IN), .ZN(n1862) );
OR3_X1 U1496 ( .A1(n1878), .A2(n1871), .A3(n1870), .ZN(n1861) );
NAND2_X1 U1497 ( .A1(n1879), .A2(n1880), .ZN(n1870) );
XNOR2_X1 U1498 ( .A(n1881), .B(KEYINPUT61), .ZN(n1879) );
NAND2_X1 U1499 ( .A1(n1882), .A2(REG4_REG_6__SCAN_IN), .ZN(n1860) );
XNOR2_X1 U1500 ( .A(n1857), .B(KEYINPUT45), .ZN(n1882) );
NAND4_X1 U1501 ( .A1(n1883), .A2(n1884), .A3(n1885), .A4(n1886), .ZN(U286));
NOR3_X1 U1502 ( .A1(n1887), .A2(n1888), .A3(n1889), .ZN(n1886) );
NOR2_X1 U1503 ( .A1(n1878), .A2(n1890), .ZN(n1889) );
XOR2_X1 U1504 ( .A(n1881), .B(n1891), .Z(n1890) );
NOR2_X1 U1505 ( .A1(KEYINPUT61), .A2(n1892), .ZN(n1891) );
NOR2_X1 U1506 ( .A1(n1893), .A2(n1871), .ZN(n1881) );
NOR2_X1 U1507 ( .A1(n1894), .A2(n1895), .ZN(n1871) );
AND2_X1 U1508 ( .A1(n1895), .A2(n1894), .ZN(n1893) );
NOR2_X1 U1509 ( .A1(n1896), .A2(n1873), .ZN(n1888) );
NAND2_X1 U1510 ( .A1(n1897), .A2(n1875), .ZN(n1873) );
NAND2_X1 U1511 ( .A1(n1898), .A2(n1899), .ZN(n1875) );
NAND2_X1 U1512 ( .A1(n1900), .A2(n1872), .ZN(n1899) );
INV_X1 U1513 ( .A(n1876), .ZN(n1872) );
NAND2_X1 U1514 ( .A1(n1895), .A2(n1901), .ZN(n1900) );
XOR2_X1 U1515 ( .A(KEYINPUT55), .B(n1902), .Z(n1898) );
NOR3_X1 U1516 ( .A1(n1903), .A2(n1902), .A3(n1876), .ZN(n1896) );
NOR2_X1 U1517 ( .A1(n1901), .A2(n1895), .ZN(n1876) );
INV_X1 U1518 ( .A(n1904), .ZN(n1895) );
NOR2_X1 U1519 ( .A1(n1905), .A2(n1904), .ZN(n1903) );
NOR2_X1 U1520 ( .A1(n1904), .A2(n1906), .ZN(n1887) );
NAND2_X1 U1521 ( .A1(n1907), .A2(n1908), .ZN(n1904) );
NAND3_X1 U1522 ( .A1(n1909), .A2(n1910), .A3(n1911), .ZN(n1908) );
NAND2_X1 U1523 ( .A1(n1912), .A2(n1913), .ZN(n1909) );
NAND3_X1 U1524 ( .A1(n1914), .A2(n1913), .A3(n1915), .ZN(n1907) );
XNOR2_X1 U1525 ( .A(KEYINPUT32), .B(n1911), .ZN(n1915) );
XOR2_X1 U1526 ( .A(n1916), .B(n1917), .Z(n1911) );
NOR2_X1 U1527 ( .A1(n1918), .A2(n1919), .ZN(n1917) );
AND2_X1 U1528 ( .A1(RMAX_REG_6__SCAN_IN), .A2(RESTART), .ZN(n1919) );
NOR2_X1 U1529 ( .A1(n1920), .A2(n1921), .ZN(n1918) );
XNOR2_X1 U1530 ( .A(DATA_IN_6_), .B(KEYINPUT9), .ZN(n1921) );
NAND2_X1 U1531 ( .A1(n1922), .A2(n1923), .ZN(n1916) );
NAND2_X1 U1532 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1924), .ZN(n1923) );
NAND2_X1 U1533 ( .A1(RESTART), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1922) );
NAND2_X1 U1534 ( .A1(n1925), .A2(n1926), .ZN(n1914) );
XNOR2_X1 U1535 ( .A(KEYINPUT19), .B(n1910), .ZN(n1925) );
NAND2_X1 U1536 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1779), .ZN(n1885) );
NAND2_X1 U1537 ( .A1(n1857), .A2(REG4_REG_5__SCAN_IN), .ZN(n1884) );
NAND2_X1 U1538 ( .A1(n1858), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1883) );
NAND4_X1 U1539 ( .A1(n1927), .A2(n1928), .A3(n1929), .A4(n1930), .ZN(U285));
NOR3_X1 U1540 ( .A1(n1931), .A2(n1932), .A3(n1933), .ZN(n1930) );
NOR3_X1 U1541 ( .A1(n1878), .A2(n1880), .A3(n1934), .ZN(n1933) );
NOR2_X1 U1542 ( .A1(n1935), .A2(n1936), .ZN(n1934) );
AND2_X1 U1543 ( .A1(n1937), .A2(n1938), .ZN(n1935) );
INV_X1 U1544 ( .A(n1892), .ZN(n1880) );
NAND3_X1 U1545 ( .A1(n1939), .A2(n1937), .A3(n1938), .ZN(n1892) );
NAND2_X1 U1546 ( .A1(n1940), .A2(n1894), .ZN(n1939) );
OR2_X1 U1547 ( .A1(n1941), .A2(n1936), .ZN(n1894) );
NAND2_X1 U1548 ( .A1(n1936), .A2(n1941), .ZN(n1940) );
NOR3_X1 U1549 ( .A1(n1877), .A2(n1902), .A3(n1942), .ZN(n1932) );
NOR2_X1 U1550 ( .A1(n1943), .A2(n1944), .ZN(n1942) );
AND2_X1 U1551 ( .A1(n1945), .A2(n1946), .ZN(n1943) );
AND3_X1 U1552 ( .A1(n1944), .A2(n1945), .A3(n1946), .ZN(n1902) );
NAND2_X1 U1553 ( .A1(n1901), .A2(n1947), .ZN(n1944) );
NAND2_X1 U1554 ( .A1(n1936), .A2(n1948), .ZN(n1947) );
INV_X1 U1555 ( .A(n1905), .ZN(n1901) );
NOR2_X1 U1556 ( .A1(n1948), .A2(n1936), .ZN(n1905) );
AND2_X1 U1557 ( .A1(n1936), .A2(n1949), .ZN(n1931) );
NAND2_X1 U1558 ( .A1(n1950), .A2(n1951), .ZN(n1936) );
NAND2_X1 U1559 ( .A1(n1912), .A2(n1952), .ZN(n1951) );
NAND2_X1 U1560 ( .A1(n1910), .A2(n1913), .ZN(n1952) );
INV_X1 U1561 ( .A(n1926), .ZN(n1912) );
NAND4_X1 U1562 ( .A1(n1953), .A2(n1954), .A3(n1910), .A4(n1926), .ZN(n1950));
NAND2_X1 U1563 ( .A1(n1955), .A2(n1956), .ZN(n1926) );
NAND2_X1 U1564 ( .A1(n1957), .A2(n1958), .ZN(n1956) );
NAND2_X1 U1565 ( .A1(n1959), .A2(n1960), .ZN(n1957) );
OR2_X1 U1566 ( .A1(n1960), .A2(n1959), .ZN(n1955) );
NAND2_X1 U1567 ( .A1(n1961), .A2(n1962), .ZN(n1910) );
NAND2_X1 U1568 ( .A1(n1963), .A2(n1964), .ZN(n1962) );
NAND2_X1 U1569 ( .A1(KEYINPUT52), .A2(n1961), .ZN(n1954) );
OR2_X1 U1570 ( .A1(n1913), .A2(KEYINPUT52), .ZN(n1953) );
NAND3_X1 U1571 ( .A1(n1963), .A2(n1964), .A3(n1965), .ZN(n1913) );
INV_X1 U1572 ( .A(n1961), .ZN(n1965) );
NAND2_X1 U1573 ( .A1(n1966), .A2(n1967), .ZN(n1961) );
NAND2_X1 U1574 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1924), .ZN(n1967) );
NAND2_X1 U1575 ( .A1(RESTART), .A2(RMIN_REG_5__SCAN_IN), .ZN(n1966) );
NAND2_X1 U1576 ( .A1(DATA_IN_5_), .A2(n1924), .ZN(n1964) );
NAND2_X1 U1577 ( .A1(RESTART), .A2(RMAX_REG_5__SCAN_IN), .ZN(n1963) );
NAND2_X1 U1578 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1779), .ZN(n1929) );
NAND2_X1 U1579 ( .A1(n1857), .A2(REG4_REG_4__SCAN_IN), .ZN(n1928) );
NAND2_X1 U1580 ( .A1(n1858), .A2(RLAST_REG_4__SCAN_IN), .ZN(n1927) );
NAND4_X1 U1581 ( .A1(n1968), .A2(n1969), .A3(n1970), .A4(n1971), .ZN(U284));
NOR3_X1 U1582 ( .A1(n1972), .A2(n1973), .A3(n1974), .ZN(n1971) );
NOR2_X1 U1583 ( .A1(n1975), .A2(n1906), .ZN(n1974) );
NOR2_X1 U1584 ( .A1(n1877), .A2(n1976), .ZN(n1973) );
XNOR2_X1 U1585 ( .A(n1945), .B(n1977), .ZN(n1976) );
NOR2_X1 U1586 ( .A1(KEYINPUT54), .A2(n1978), .ZN(n1977) );
INV_X1 U1587 ( .A(n1946), .ZN(n1978) );
NAND2_X1 U1588 ( .A1(n1948), .A2(n1979), .ZN(n1945) );
NAND2_X1 U1589 ( .A1(n1980), .A2(n1981), .ZN(n1948) );
XNOR2_X1 U1590 ( .A(KEYINPUT22), .B(n1975), .ZN(n1980) );
INV_X1 U1591 ( .A(n1897), .ZN(n1877) );
AND2_X1 U1592 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1858), .ZN(n1972) );
NAND2_X1 U1593 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1982), .ZN(n1970) );
XNOR2_X1 U1594 ( .A(KEYINPUT57), .B(n1983), .ZN(n1982) );
NAND2_X1 U1595 ( .A1(n1984), .A2(n1869), .ZN(n1969) );
XOR2_X1 U1596 ( .A(n1938), .B(n1937), .Z(n1984) );
NAND2_X1 U1597 ( .A1(n1941), .A2(n1979), .ZN(n1937) );
NAND2_X1 U1598 ( .A1(n1985), .A2(n1986), .ZN(n1979) );
NAND2_X1 U1599 ( .A1(n1981), .A2(n1975), .ZN(n1941) );
INV_X1 U1600 ( .A(n1985), .ZN(n1975) );
XOR2_X1 U1601 ( .A(n1987), .B(n1960), .Z(n1985) );
NAND2_X1 U1602 ( .A1(n1988), .A2(n1989), .ZN(n1960) );
NAND2_X1 U1603 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1924), .ZN(n1989) );
NAND2_X1 U1604 ( .A1(RESTART), .A2(RMIN_REG_4__SCAN_IN), .ZN(n1988) );
NAND2_X1 U1605 ( .A1(n1990), .A2(n1991), .ZN(n1987) );
OR2_X1 U1606 ( .A1(n1958), .A2(n1959), .ZN(n1991) );
NAND2_X1 U1607 ( .A1(n1992), .A2(n1958), .ZN(n1990) );
NAND2_X1 U1608 ( .A1(n1993), .A2(n1994), .ZN(n1958) );
NAND2_X1 U1609 ( .A1(n1995), .A2(n1996), .ZN(n1994) );
NAND2_X1 U1610 ( .A1(n1997), .A2(n1998), .ZN(n1996) );
OR2_X1 U1611 ( .A1(n1998), .A2(n1997), .ZN(n1993) );
NAND2_X1 U1612 ( .A1(KEYINPUT46), .A2(n1999), .ZN(n1992) );
INV_X1 U1613 ( .A(n1959), .ZN(n1999) );
NAND2_X1 U1614 ( .A1(n2000), .A2(n2001), .ZN(n1959) );
NAND2_X1 U1615 ( .A1(DATA_IN_4_), .A2(n1924), .ZN(n2001) );
NAND2_X1 U1616 ( .A1(RESTART), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2000) );
NAND2_X1 U1617 ( .A1(n2002), .A2(DATA_OUT_REG_3__SCAN_IN), .ZN(n1968) );
XNOR2_X1 U1618 ( .A(n1779), .B(KEYINPUT23), .ZN(n2002) );
NAND4_X1 U1619 ( .A1(n2003), .A2(n2004), .A3(n2005), .A4(n2006), .ZN(U283));
NOR3_X1 U1620 ( .A1(n2007), .A2(n2008), .A3(n2009), .ZN(n2006) );
NOR3_X1 U1621 ( .A1(n1878), .A2(n1938), .A3(n2010), .ZN(n2009) );
NOR2_X1 U1622 ( .A1(n2011), .A2(n2012), .ZN(n2010) );
NOR2_X1 U1623 ( .A1(n2013), .A2(n2014), .ZN(n2011) );
NOR3_X1 U1624 ( .A1(n2015), .A2(n2013), .A3(n2014), .ZN(n1938) );
NOR3_X1 U1625 ( .A1(n2016), .A2(n1946), .A3(n2017), .ZN(n2008) );
NOR2_X1 U1626 ( .A1(n2018), .A2(n2012), .ZN(n2017) );
NOR2_X1 U1627 ( .A1(n2013), .A2(n2019), .ZN(n2018) );
NOR3_X1 U1628 ( .A1(n2015), .A2(n2013), .A3(n2019), .ZN(n1946) );
INV_X1 U1629 ( .A(n2012), .ZN(n2015) );
NAND2_X1 U1630 ( .A1(n1986), .A2(n2020), .ZN(n2012) );
NAND2_X1 U1631 ( .A1(n2021), .A2(n2022), .ZN(n2020) );
INV_X1 U1632 ( .A(n1981), .ZN(n1986) );
NOR2_X1 U1633 ( .A1(n2022), .A2(n2021), .ZN(n1981) );
XNOR2_X1 U1634 ( .A(n1897), .B(KEYINPUT44), .ZN(n2016) );
NOR2_X1 U1635 ( .A1(n2023), .A2(n2024), .ZN(n2007) );
XNOR2_X1 U1636 ( .A(n1857), .B(KEYINPUT10), .ZN(n2023) );
NAND2_X1 U1637 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1779), .ZN(n2005) );
NAND2_X1 U1638 ( .A1(n1949), .A2(n2021), .ZN(n2004) );
XOR2_X1 U1639 ( .A(n2025), .B(n2026), .Z(n2021) );
XOR2_X1 U1640 ( .A(n1998), .B(n1997), .Z(n2026) );
NAND2_X1 U1641 ( .A1(n2027), .A2(n2028), .ZN(n1997) );
NAND2_X1 U1642 ( .A1(n2029), .A2(RESTART), .ZN(n2028) );
XNOR2_X1 U1643 ( .A(RMAX_REG_3__SCAN_IN), .B(KEYINPUT7), .ZN(n2029) );
NAND2_X1 U1644 ( .A1(DATA_IN_3_), .A2(n1924), .ZN(n2027) );
NAND2_X1 U1645 ( .A1(n2030), .A2(n2031), .ZN(n1998) );
NAND2_X1 U1646 ( .A1(n2032), .A2(REG4_REG_3__SCAN_IN), .ZN(n2031) );
XNOR2_X1 U1647 ( .A(n1924), .B(KEYINPUT4), .ZN(n2032) );
NAND2_X1 U1648 ( .A1(RESTART), .A2(RMIN_REG_3__SCAN_IN), .ZN(n2030) );
NAND2_X1 U1649 ( .A1(KEYINPUT33), .A2(n1995), .ZN(n2025) );
AND2_X1 U1650 ( .A1(n2033), .A2(n2034), .ZN(n1995) );
NAND2_X1 U1651 ( .A1(n2035), .A2(n2036), .ZN(n2034) );
XOR2_X1 U1652 ( .A(KEYINPUT2), .B(n2037), .Z(n2033) );
NOR2_X1 U1653 ( .A1(n2038), .A2(n2039), .ZN(n2037) );
INV_X1 U1654 ( .A(n2040), .ZN(n2039) );
NOR2_X1 U1655 ( .A1(n2035), .A2(n2036), .ZN(n2038) );
NAND2_X1 U1656 ( .A1(n1858), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2003) );
NAND4_X1 U1657 ( .A1(n2041), .A2(n2042), .A3(n2043), .A4(n2044), .ZN(U282));
NOR3_X1 U1658 ( .A1(n2045), .A2(n2046), .A3(n2047), .ZN(n2044) );
AND2_X1 U1659 ( .A1(n2048), .A2(n1949), .ZN(n2047) );
INV_X1 U1660 ( .A(n1906), .ZN(n1949) );
NOR2_X1 U1661 ( .A1(n2049), .A2(n2050), .ZN(n2046) );
XNOR2_X1 U1662 ( .A(n1897), .B(KEYINPUT53), .ZN(n2050) );
XNOR2_X1 U1663 ( .A(n2051), .B(n2019), .ZN(n2049) );
NAND2_X1 U1664 ( .A1(KEYINPUT27), .A2(n2052), .ZN(n2051) );
NOR2_X1 U1665 ( .A1(n2053), .A2(n1983), .ZN(n2045) );
XOR2_X1 U1666 ( .A(KEYINPUT21), .B(n2054), .Z(n2043) );
NOR2_X1 U1667 ( .A1(n2055), .A2(n1878), .ZN(n2054) );
XNOR2_X1 U1668 ( .A(n2013), .B(n2014), .ZN(n2055) );
INV_X1 U1669 ( .A(n2052), .ZN(n2013) );
NAND2_X1 U1670 ( .A1(n2056), .A2(n2022), .ZN(n2052) );
OR3_X1 U1671 ( .A1(n2057), .A2(n2058), .A3(n2048), .ZN(n2022) );
NAND2_X1 U1672 ( .A1(n2048), .A2(n2059), .ZN(n2056) );
NAND2_X1 U1673 ( .A1(n2060), .A2(n2061), .ZN(n2059) );
NAND3_X1 U1674 ( .A1(n2062), .A2(n2063), .A3(n2064), .ZN(n2048) );
OR2_X1 U1675 ( .A1(n2040), .A2(n2065), .ZN(n2064) );
NAND3_X1 U1676 ( .A1(n2065), .A2(n2040), .A3(KEYINPUT59), .ZN(n2063) );
NAND2_X1 U1677 ( .A1(n2066), .A2(n2067), .ZN(n2040) );
NAND2_X1 U1678 ( .A1(n2068), .A2(n2069), .ZN(n2067) );
NAND2_X1 U1679 ( .A1(n2070), .A2(n2071), .ZN(n2068) );
XOR2_X1 U1680 ( .A(n2072), .B(KEYINPUT15), .Z(n2066) );
OR2_X1 U1681 ( .A1(n2071), .A2(n2070), .ZN(n2072) );
XOR2_X1 U1682 ( .A(n2073), .B(n2036), .Z(n2065) );
NAND2_X1 U1683 ( .A1(KEYINPUT31), .A2(n2035), .ZN(n2073) );
OR3_X1 U1684 ( .A1(n2035), .A2(n2074), .A3(KEYINPUT59), .ZN(n2062) );
INV_X1 U1685 ( .A(n2036), .ZN(n2074) );
NAND2_X1 U1686 ( .A1(n2075), .A2(n2076), .ZN(n2036) );
NAND2_X1 U1687 ( .A1(DATA_IN_2_), .A2(n1924), .ZN(n2076) );
NAND2_X1 U1688 ( .A1(RESTART), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2075) );
NAND2_X1 U1689 ( .A1(n2077), .A2(n2078), .ZN(n2035) );
NAND2_X1 U1690 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1924), .ZN(n2078) );
NAND2_X1 U1691 ( .A1(RESTART), .A2(RMIN_REG_2__SCAN_IN), .ZN(n2077) );
NAND2_X1 U1692 ( .A1(n1858), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2042) );
NAND2_X1 U1693 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1779), .ZN(n2041) );
NAND4_X1 U1694 ( .A1(n2079), .A2(n2080), .A3(n2081), .A4(n2082), .ZN(U281));
NOR3_X1 U1695 ( .A1(n2083), .A2(n2084), .A3(n2085), .ZN(n2082) );
NOR2_X1 U1696 ( .A1(n2060), .A2(n1906), .ZN(n2085) );
NAND4_X1 U1697 ( .A1(STATO_REG_1__SCAN_IN), .A2(n2086), .A3(n2087), .A4(U280), .ZN(n1906) );
NAND2_X1 U1698 ( .A1(n1924), .A2(n2088), .ZN(n2087) );
NAND3_X1 U1699 ( .A1(n2089), .A2(n2090), .A3(ENABLE), .ZN(n2088) );
NAND2_X1 U1700 ( .A1(RESTART), .A2(n2091), .ZN(n2086) );
NOR2_X1 U1701 ( .A1(n2092), .A2(n1983), .ZN(n2084) );
INV_X1 U1702 ( .A(n1857), .ZN(n1983) );
NOR3_X1 U1703 ( .A1(n1773), .A2(n2093), .A3(n2090), .ZN(n1857) );
INV_X1 U1704 ( .A(AVERAGE), .ZN(n2090) );
AND2_X1 U1705 ( .A1(n2014), .A2(n1869), .ZN(n2083) );
INV_X1 U1706 ( .A(n1878), .ZN(n1869) );
NAND4_X1 U1707 ( .A1(RESTART), .A2(STATO_REG_1__SCAN_IN), .A3(n2091), .A4(
U280), .ZN(n1878) );
XNOR2_X1 U1708 ( .A(n2094), .B(KEYINPUT62), .ZN(n2091) );
NAND2_X1 U1709 ( .A1(n2095), .A2(n2096), .ZN(n2094) );
NAND2_X1 U1710 ( .A1(n1727), .A2(n1722), .ZN(n2096) );
INV_X1 U1711 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1722) );
NAND3_X1 U1712 ( .A1(n2097), .A2(n2098), .A3(n2099), .ZN(n2095) );
OR2_X1 U1713 ( .A1(n2100), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2099) );
NAND2_X1 U1714 ( .A1(n2101), .A2(n1721), .ZN(n2098) );
INV_X1 U1715 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1721) );
NAND2_X1 U1716 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n2100), .ZN(n2101) );
NAND2_X1 U1717 ( .A1(n2102), .A2(n2103), .ZN(n2100) );
NAND2_X1 U1718 ( .A1(RMIN_REG_5__SCAN_IN), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2103) );
XOR2_X1 U1719 ( .A(KEYINPUT42), .B(n2104), .Z(n2102) );
NOR3_X1 U1720 ( .A1(n2105), .A2(n2106), .A3(n2107), .ZN(n2104) );
NOR2_X1 U1721 ( .A1(RMAX_REG_5__SCAN_IN), .A2(RMIN_REG_5__SCAN_IN), .ZN(n2107) );
NOR2_X1 U1722 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n2108), .ZN(n2106) );
NOR2_X1 U1723 ( .A1(n2109), .A2(n2110), .ZN(n2108) );
XOR2_X1 U1724 ( .A(RMAX_REG_4__SCAN_IN), .B(KEYINPUT49), .Z(n2110) );
NOR2_X1 U1725 ( .A1(n2111), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2105) );
INV_X1 U1726 ( .A(n2109), .ZN(n2111) );
NAND2_X1 U1727 ( .A1(n2112), .A2(n2113), .ZN(n2109) );
NAND3_X1 U1728 ( .A1(n2114), .A2(n2115), .A3(n2116), .ZN(n2113) );
NAND2_X1 U1729 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2116) );
NAND3_X1 U1730 ( .A1(n2117), .A2(n2118), .A3(n2119), .ZN(n2115) );
NAND2_X1 U1731 ( .A1(n1744), .A2(n1716), .ZN(n2119) );
INV_X1 U1732 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1716) );
INV_X1 U1733 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1744) );
NAND2_X1 U1734 ( .A1(n2120), .A2(n2121), .ZN(n2118) );
NAND2_X1 U1735 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2121) );
XOR2_X1 U1736 ( .A(n2122), .B(KEYINPUT1), .Z(n2120) );
NAND2_X1 U1737 ( .A1(RMIN_REG_1__SCAN_IN), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2122) );
NAND2_X1 U1738 ( .A1(n2123), .A2(n2124), .ZN(n2117) );
INV_X1 U1739 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n2124) );
XNOR2_X1 U1740 ( .A(RMAX_REG_1__SCAN_IN), .B(KEYINPUT40), .ZN(n2123) );
NAND2_X1 U1741 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2114) );
NAND2_X1 U1742 ( .A1(n1748), .A2(n1707), .ZN(n2112) );
INV_X1 U1743 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1707) );
INV_X1 U1744 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1748) );
NAND2_X1 U1745 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n2125), .ZN(n2097) );
XNOR2_X1 U1746 ( .A(n1727), .B(KEYINPUT24), .ZN(n2125) );
INV_X1 U1747 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1727) );
XOR2_X1 U1748 ( .A(n2057), .B(n2058), .Z(n2014) );
XOR2_X1 U1749 ( .A(n2126), .B(KEYINPUT38), .Z(n2081) );
NAND2_X1 U1750 ( .A1(n1897), .A2(n2019), .ZN(n2126) );
NAND2_X1 U1751 ( .A1(n2127), .A2(n2128), .ZN(n2019) );
NAND2_X1 U1752 ( .A1(n2058), .A2(n2060), .ZN(n2128) );
INV_X1 U1753 ( .A(n2057), .ZN(n2060) );
INV_X1 U1754 ( .A(n2061), .ZN(n2058) );
XOR2_X1 U1755 ( .A(n2129), .B(KEYINPUT3), .Z(n2127) );
NAND2_X1 U1756 ( .A1(n2057), .A2(n2061), .ZN(n2129) );
NAND2_X1 U1757 ( .A1(n2071), .A2(n2130), .ZN(n2061) );
NAND2_X1 U1758 ( .A1(n2131), .A2(n2132), .ZN(n2130) );
NAND2_X1 U1759 ( .A1(n1924), .A2(n2133), .ZN(n2132) );
NAND2_X1 U1760 ( .A1(n1713), .A2(n2092), .ZN(n2133) );
NAND2_X1 U1761 ( .A1(RESTART), .A2(n2134), .ZN(n2131) );
NAND2_X1 U1762 ( .A1(n1746), .A2(n2135), .ZN(n2134) );
XNOR2_X1 U1763 ( .A(n2071), .B(n2136), .ZN(n2057) );
XNOR2_X1 U1764 ( .A(n2070), .B(n2069), .ZN(n2136) );
NAND2_X1 U1765 ( .A1(n2137), .A2(n2138), .ZN(n2069) );
NAND2_X1 U1766 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1924), .ZN(n2138) );
NAND2_X1 U1767 ( .A1(RESTART), .A2(RMIN_REG_1__SCAN_IN), .ZN(n2137) );
AND2_X1 U1768 ( .A1(n2139), .A2(n2140), .ZN(n2070) );
NAND2_X1 U1769 ( .A1(DATA_IN_1_), .A2(n1924), .ZN(n2140) );
NAND2_X1 U1770 ( .A1(RESTART), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2139) );
NAND4_X1 U1771 ( .A1(n2141), .A2(n2142), .A3(n2143), .A4(n2144), .ZN(n2071));
NAND2_X1 U1772 ( .A1(n1920), .A2(n2145), .ZN(n2144) );
NAND3_X1 U1773 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .A3(
RESTART), .ZN(n2145) );
INV_X1 U1774 ( .A(n1924), .ZN(n1920) );
OR2_X1 U1775 ( .A1(n2146), .A2(RESTART), .ZN(n2143) );
NAND2_X1 U1776 ( .A1(n1713), .A2(n1746), .ZN(n2142) );
INV_X1 U1777 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1746) );
NAND2_X1 U1778 ( .A1(n2092), .A2(n2135), .ZN(n2141) );
INV_X1 U1779 ( .A(RMIN_REG_0__SCAN_IN), .ZN(n2135) );
NAND2_X1 U1780 ( .A1(n2147), .A2(n2148), .ZN(n2089) );
NAND2_X1 U1781 ( .A1(n2149), .A2(n2150), .ZN(n2148) );
INV_X1 U1782 ( .A(REG4_REG_7__SCAN_IN), .ZN(n2150) );
OR2_X1 U1783 ( .A1(n2151), .A2(n1691), .ZN(n2149) );
NAND2_X1 U1784 ( .A1(n2151), .A2(n1691), .ZN(n2147) );
INV_X1 U1785 ( .A(DATA_IN_7_), .ZN(n1691) );
NAND2_X1 U1786 ( .A1(n2152), .A2(n2153), .ZN(n2151) );
NAND2_X1 U1787 ( .A1(REG4_REG_6__SCAN_IN), .A2(n2154), .ZN(n2153) );
NAND2_X1 U1788 ( .A1(n2155), .A2(n1695), .ZN(n2154) );
XOR2_X1 U1789 ( .A(n2156), .B(KEYINPUT35), .Z(n2155) );
OR2_X1 U1790 ( .A1(n2156), .A2(n1695), .ZN(n2152) );
INV_X1 U1791 ( .A(DATA_IN_6_), .ZN(n1695) );
NAND2_X1 U1792 ( .A1(n2157), .A2(n2158), .ZN(n2156) );
OR2_X1 U1793 ( .A1(DATA_IN_5_), .A2(REG4_REG_5__SCAN_IN), .ZN(n2158) );
NAND3_X1 U1794 ( .A1(n2159), .A2(n2160), .A3(n2161), .ZN(n2157) );
NAND2_X1 U1795 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2161) );
NAND3_X1 U1796 ( .A1(n2162), .A2(n2163), .A3(n2164), .ZN(n2160) );
OR2_X1 U1797 ( .A1(DATA_IN_4_), .A2(REG4_REG_4__SCAN_IN), .ZN(n2164) );
NAND3_X1 U1798 ( .A1(n2165), .A2(n2166), .A3(n2167), .ZN(n2163) );
NAND2_X1 U1799 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2167) );
NAND3_X1 U1800 ( .A1(n2168), .A2(n2169), .A3(n2170), .ZN(n2166) );
NAND2_X1 U1801 ( .A1(n1711), .A2(n2024), .ZN(n2170) );
INV_X1 U1802 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2024) );
INV_X1 U1803 ( .A(DATA_IN_2_), .ZN(n1711) );
NAND2_X1 U1804 ( .A1(n2171), .A2(n2172), .ZN(n2169) );
NAND2_X1 U1805 ( .A1(REG4_REG_1__SCAN_IN), .A2(DATA_IN_1_), .ZN(n2172) );
XOR2_X1 U1806 ( .A(KEYINPUT11), .B(n2146), .Z(n2171) );
NOR2_X1 U1807 ( .A1(n2092), .A2(n1713), .ZN(n2146) );
INV_X1 U1808 ( .A(DATA_IN_0_), .ZN(n1713) );
INV_X1 U1809 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2092) );
NAND2_X1 U1810 ( .A1(n1715), .A2(n2053), .ZN(n2168) );
INV_X1 U1811 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2053) );
INV_X1 U1812 ( .A(DATA_IN_1_), .ZN(n1715) );
NAND2_X1 U1813 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2165) );
OR2_X1 U1814 ( .A1(DATA_IN_3_), .A2(REG4_REG_3__SCAN_IN), .ZN(n2162) );
NAND2_X1 U1815 ( .A1(REG4_REG_4__SCAN_IN), .A2(n2173), .ZN(n2159) );
XNOR2_X1 U1816 ( .A(KEYINPUT48), .B(n1699), .ZN(n2173) );
INV_X1 U1817 ( .A(DATA_IN_4_), .ZN(n1699) );
INV_X1 U1818 ( .A(ENABLE), .ZN(n1773) );
NAND2_X1 U1819 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1779), .ZN(n2080) );
XOR2_X1 U1820 ( .A(KEYINPUT30), .B(n2174), .Z(n2079) );
AND2_X1 U1821 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1858), .ZN(n2174) );
NOR2_X1 U1822 ( .A1(n2093), .A2(ENABLE), .ZN(n1858) );
NAND3_X1 U1823 ( .A1(n1924), .A2(U280), .A3(STATO_REG_1__SCAN_IN), .ZN(n2093) );
NAND2_X1 U1824 ( .A1(n1812), .A2(n2175), .ZN(U280) );
NAND2_X1 U1825 ( .A1(STATO_REG_0__SCAN_IN), .A2(n2176), .ZN(n2175) );
XOR2_X1 U1826 ( .A(STATO_REG_1__SCAN_IN), .B(KEYINPUT56), .Z(n2176) );
NAND2_X1 U1827 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1662), .ZN(n1812) );
INV_X1 U1828 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1662) );
endmodule


