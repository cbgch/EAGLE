//Key = 0010010110000010010100101011000000101001010101110011000001111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322;

XOR2_X1 U724 ( .A(n1006), .B(n1007), .Z(G9) );
NAND4_X1 U725 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(G75) );
NAND4_X1 U726 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1010) );
NOR4_X1 U727 ( .A1(n1016), .A2(n1017), .A3(n1018), .A4(n1019), .ZN(n1015) );
XNOR2_X1 U728 ( .A(G472), .B(n1020), .ZN(n1018) );
NOR2_X1 U729 ( .A1(n1021), .A2(KEYINPUT52), .ZN(n1020) );
NOR2_X1 U730 ( .A1(n1022), .A2(n1023), .ZN(n1014) );
XNOR2_X1 U731 ( .A(n1024), .B(n1025), .ZN(n1023) );
NOR2_X1 U732 ( .A1(KEYINPUT61), .A2(n1026), .ZN(n1025) );
XOR2_X1 U733 ( .A(n1027), .B(G469), .Z(n1013) );
NAND2_X1 U734 ( .A1(KEYINPUT41), .A2(n1028), .ZN(n1027) );
XNOR2_X1 U735 ( .A(KEYINPUT54), .B(n1029), .ZN(n1028) );
XOR2_X1 U736 ( .A(n1030), .B(n1031), .Z(n1012) );
NAND2_X1 U737 ( .A1(n1032), .A2(n1033), .ZN(n1009) );
NAND2_X1 U738 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND4_X1 U739 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
NAND2_X1 U740 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND3_X1 U741 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1040) );
INV_X1 U742 ( .A(KEYINPUT45), .ZN(n1043) );
NAND4_X1 U743 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1038) );
NAND2_X1 U744 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NAND3_X1 U745 ( .A1(n1044), .A2(n1042), .A3(KEYINPUT45), .ZN(n1046) );
NAND2_X1 U746 ( .A1(n1051), .A2(n1052), .ZN(n1045) );
NAND2_X1 U747 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND3_X1 U748 ( .A1(n1051), .A2(n1055), .A3(n1049), .ZN(n1034) );
NAND2_X1 U749 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U750 ( .A1(n1048), .A2(n1058), .ZN(n1057) );
NAND2_X1 U751 ( .A1(n1037), .A2(n1059), .ZN(n1056) );
NAND2_X1 U752 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U753 ( .A1(n1036), .A2(n1062), .ZN(n1061) );
NAND2_X1 U754 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U755 ( .A1(n1017), .A2(n1065), .ZN(n1064) );
NAND2_X1 U756 ( .A1(n1048), .A2(n1016), .ZN(n1060) );
INV_X1 U757 ( .A(n1066), .ZN(n1032) );
NAND2_X1 U758 ( .A1(n1067), .A2(n1068), .ZN(G72) );
NAND2_X1 U759 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U760 ( .A1(G953), .A2(n1071), .ZN(n1070) );
NAND2_X1 U761 ( .A1(G900), .A2(G227), .ZN(n1071) );
INV_X1 U762 ( .A(n1072), .ZN(n1069) );
NAND2_X1 U763 ( .A1(n1072), .A2(n1073), .ZN(n1067) );
NAND2_X1 U764 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U765 ( .A1(G953), .A2(n1076), .ZN(n1075) );
INV_X1 U766 ( .A(n1077), .ZN(n1074) );
XOR2_X1 U767 ( .A(n1078), .B(n1079), .Z(n1072) );
NOR3_X1 U768 ( .A1(n1080), .A2(n1081), .A3(n1077), .ZN(n1079) );
AND2_X1 U769 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XOR2_X1 U770 ( .A(KEYINPUT18), .B(n1084), .Z(n1080) );
NOR2_X1 U771 ( .A1(n1083), .A2(n1082), .ZN(n1084) );
NAND2_X1 U772 ( .A1(n1085), .A2(n1086), .ZN(n1078) );
XOR2_X1 U773 ( .A(n1011), .B(KEYINPUT33), .Z(n1085) );
XOR2_X1 U774 ( .A(n1087), .B(n1088), .Z(G69) );
XOR2_X1 U775 ( .A(n1089), .B(n1090), .Z(n1088) );
NAND2_X1 U776 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U777 ( .A1(G898), .A2(G224), .ZN(n1092) );
XOR2_X1 U778 ( .A(n1011), .B(KEYINPUT7), .Z(n1091) );
NAND4_X1 U779 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1089) );
NAND3_X1 U780 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
INV_X1 U781 ( .A(n1100), .ZN(n1099) );
NAND2_X1 U782 ( .A1(n1101), .A2(n1100), .ZN(n1095) );
NAND2_X1 U783 ( .A1(n1102), .A2(n1098), .ZN(n1101) );
XNOR2_X1 U784 ( .A(KEYINPUT17), .B(n1097), .ZN(n1102) );
NAND2_X1 U785 ( .A1(G953), .A2(n1103), .ZN(n1094) );
OR2_X1 U786 ( .A1(n1098), .A2(n1097), .ZN(n1093) );
NAND2_X1 U787 ( .A1(n1104), .A2(n1105), .ZN(n1097) );
INV_X1 U788 ( .A(KEYINPUT42), .ZN(n1098) );
AND2_X1 U789 ( .A1(n1106), .A2(n1011), .ZN(n1087) );
NOR2_X1 U790 ( .A1(n1107), .A2(n1108), .ZN(G66) );
XNOR2_X1 U791 ( .A(n1109), .B(n1110), .ZN(n1108) );
AND2_X1 U792 ( .A1(G217), .A2(n1111), .ZN(n1110) );
NOR2_X1 U793 ( .A1(n1107), .A2(n1112), .ZN(G63) );
XOR2_X1 U794 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U795 ( .A1(n1031), .A2(n1115), .ZN(n1113) );
NOR2_X1 U796 ( .A1(n1107), .A2(n1116), .ZN(G60) );
XOR2_X1 U797 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U798 ( .A1(KEYINPUT16), .A2(n1119), .ZN(n1118) );
NAND2_X1 U799 ( .A1(n1111), .A2(G475), .ZN(n1117) );
XNOR2_X1 U800 ( .A(G104), .B(n1120), .ZN(G6) );
NOR3_X1 U801 ( .A1(n1107), .A2(n1121), .A3(n1122), .ZN(G57) );
NOR3_X1 U802 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1122) );
NOR2_X1 U803 ( .A1(KEYINPUT40), .A2(n1126), .ZN(n1124) );
INV_X1 U804 ( .A(KEYINPUT3), .ZN(n1126) );
NOR2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1121) );
INV_X1 U806 ( .A(n1123), .ZN(n1128) );
XOR2_X1 U807 ( .A(n1129), .B(n1130), .Z(n1123) );
AND2_X1 U808 ( .A1(G472), .A2(n1111), .ZN(n1130) );
NAND2_X1 U809 ( .A1(KEYINPUT59), .A2(n1131), .ZN(n1129) );
XOR2_X1 U810 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U812 ( .A1(KEYINPUT50), .A2(n1136), .ZN(n1134) );
NOR2_X1 U813 ( .A1(KEYINPUT3), .A2(n1137), .ZN(n1127) );
XOR2_X1 U814 ( .A(n1125), .B(KEYINPUT40), .Z(n1137) );
NAND2_X1 U815 ( .A1(n1138), .A2(n1139), .ZN(n1125) );
NAND2_X1 U816 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR2_X1 U817 ( .A1(n1107), .A2(n1142), .ZN(G54) );
XOR2_X1 U818 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U819 ( .A(n1136), .B(n1145), .Z(n1144) );
XOR2_X1 U820 ( .A(n1146), .B(n1132), .Z(n1145) );
NAND2_X1 U821 ( .A1(KEYINPUT27), .A2(n1147), .ZN(n1146) );
XOR2_X1 U822 ( .A(n1148), .B(n1149), .Z(n1143) );
XOR2_X1 U823 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U824 ( .A1(G110), .A2(KEYINPUT32), .ZN(n1151) );
AND2_X1 U825 ( .A1(G469), .A2(n1111), .ZN(n1150) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1148) );
NOR2_X1 U827 ( .A1(n1107), .A2(n1154), .ZN(G51) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U829 ( .A(n1157), .B(n1158), .Z(n1155) );
NOR2_X1 U830 ( .A1(n1159), .A2(n1115), .ZN(n1158) );
INV_X1 U831 ( .A(n1111), .ZN(n1115) );
NOR2_X1 U832 ( .A1(n1160), .A2(n1008), .ZN(n1111) );
NOR2_X1 U833 ( .A1(n1106), .A2(n1086), .ZN(n1008) );
NAND4_X1 U834 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1086) );
NOR4_X1 U835 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
NOR3_X1 U836 ( .A1(n1169), .A2(n1170), .A3(n1054), .ZN(n1168) );
NOR3_X1 U837 ( .A1(n1171), .A2(n1172), .A3(n1053), .ZN(n1167) );
AND2_X1 U838 ( .A1(n1173), .A2(n1174), .ZN(n1163) );
NAND4_X1 U839 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1106) );
AND4_X1 U840 ( .A1(n1007), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1178) );
NAND3_X1 U841 ( .A1(n1182), .A2(n1051), .A3(n1183), .ZN(n1007) );
AND2_X1 U842 ( .A1(n1184), .A2(n1120), .ZN(n1177) );
NAND3_X1 U843 ( .A1(n1182), .A2(n1051), .A3(n1185), .ZN(n1120) );
NAND2_X1 U844 ( .A1(KEYINPUT46), .A2(n1186), .ZN(n1157) );
XOR2_X1 U845 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U846 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U847 ( .A1(KEYINPUT4), .A2(n1191), .ZN(n1190) );
NOR2_X1 U848 ( .A1(KEYINPUT15), .A2(n1192), .ZN(n1189) );
NOR2_X1 U849 ( .A1(n1193), .A2(G952), .ZN(n1107) );
XOR2_X1 U850 ( .A(G953), .B(KEYINPUT57), .Z(n1193) );
XNOR2_X1 U851 ( .A(n1166), .B(n1194), .ZN(G48) );
NAND2_X1 U852 ( .A1(KEYINPUT19), .A2(G146), .ZN(n1194) );
NOR3_X1 U853 ( .A1(n1053), .A2(n1063), .A3(n1169), .ZN(n1166) );
XOR2_X1 U854 ( .A(G143), .B(n1165), .Z(G45) );
AND3_X1 U855 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1165) );
AND3_X1 U856 ( .A1(n1198), .A2(n1199), .A3(n1022), .ZN(n1197) );
XOR2_X1 U857 ( .A(n1152), .B(n1174), .Z(G42) );
NAND2_X1 U858 ( .A1(n1200), .A2(n1201), .ZN(n1174) );
XNOR2_X1 U859 ( .A(G137), .B(n1173), .ZN(G39) );
NAND3_X1 U860 ( .A1(n1202), .A2(n1044), .A3(n1200), .ZN(n1173) );
XNOR2_X1 U861 ( .A(G134), .B(n1161), .ZN(G36) );
NAND3_X1 U862 ( .A1(n1183), .A2(n1050), .A3(n1200), .ZN(n1161) );
INV_X1 U863 ( .A(n1171), .ZN(n1200) );
NAND4_X1 U864 ( .A1(n1037), .A2(n1203), .A3(n1036), .A4(n1199), .ZN(n1171) );
XOR2_X1 U865 ( .A(n1204), .B(n1205), .Z(G33) );
NAND2_X1 U866 ( .A1(G131), .A2(n1206), .ZN(n1205) );
XOR2_X1 U867 ( .A(KEYINPUT2), .B(KEYINPUT0), .Z(n1206) );
NAND4_X1 U868 ( .A1(n1207), .A2(n1196), .A3(n1037), .A4(n1185), .ZN(n1204) );
AND3_X1 U869 ( .A1(n1036), .A2(n1203), .A3(n1050), .ZN(n1196) );
XOR2_X1 U870 ( .A(n1199), .B(KEYINPUT49), .Z(n1207) );
XOR2_X1 U871 ( .A(G128), .B(n1208), .Z(G30) );
NOR3_X1 U872 ( .A1(n1209), .A2(n1170), .A3(n1169), .ZN(n1208) );
NAND4_X1 U873 ( .A1(n1202), .A2(n1058), .A3(n1210), .A4(n1199), .ZN(n1169) );
XOR2_X1 U874 ( .A(KEYINPUT22), .B(n1183), .Z(n1209) );
XOR2_X1 U875 ( .A(n1141), .B(n1184), .Z(G3) );
NAND3_X1 U876 ( .A1(n1182), .A2(n1050), .A3(n1049), .ZN(n1184) );
NAND3_X1 U877 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(G27) );
NAND2_X1 U878 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND3_X1 U879 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
NAND2_X1 U880 ( .A1(KEYINPUT10), .A2(n1219), .ZN(n1218) );
NAND2_X1 U881 ( .A1(G125), .A2(n1220), .ZN(n1217) );
INV_X1 U882 ( .A(KEYINPUT36), .ZN(n1220) );
NAND2_X1 U883 ( .A1(KEYINPUT36), .A2(n1221), .ZN(n1216) );
NAND2_X1 U884 ( .A1(G125), .A2(n1222), .ZN(n1221) );
NAND2_X1 U885 ( .A1(KEYINPUT13), .A2(n1223), .ZN(n1222) );
INV_X1 U886 ( .A(n1162), .ZN(n1214) );
NAND4_X1 U887 ( .A1(n1162), .A2(n1219), .A3(G125), .A4(n1223), .ZN(n1212) );
INV_X1 U888 ( .A(KEYINPUT10), .ZN(n1223) );
INV_X1 U889 ( .A(KEYINPUT13), .ZN(n1219) );
NAND2_X1 U890 ( .A1(KEYINPUT10), .A2(n1224), .ZN(n1211) );
NAND2_X1 U891 ( .A1(G125), .A2(n1225), .ZN(n1224) );
NAND2_X1 U892 ( .A1(KEYINPUT13), .A2(n1162), .ZN(n1225) );
NAND4_X1 U893 ( .A1(n1201), .A2(n1048), .A3(n1058), .A4(n1199), .ZN(n1162) );
NAND2_X1 U894 ( .A1(n1066), .A2(n1226), .ZN(n1199) );
NAND3_X1 U895 ( .A1(G902), .A2(n1227), .A3(n1077), .ZN(n1226) );
NOR2_X1 U896 ( .A1(n1011), .A2(G900), .ZN(n1077) );
INV_X1 U897 ( .A(n1041), .ZN(n1048) );
NOR3_X1 U898 ( .A1(n1228), .A2(n1202), .A3(n1053), .ZN(n1201) );
INV_X1 U899 ( .A(n1185), .ZN(n1053) );
XNOR2_X1 U900 ( .A(n1175), .B(n1229), .ZN(G24) );
NOR2_X1 U901 ( .A1(KEYINPUT20), .A2(n1230), .ZN(n1229) );
NAND4_X1 U902 ( .A1(n1195), .A2(n1231), .A3(n1198), .A4(n1051), .ZN(n1175) );
NAND2_X1 U903 ( .A1(n1232), .A2(n1233), .ZN(n1051) );
OR2_X1 U904 ( .A1(n1172), .A2(KEYINPUT34), .ZN(n1233) );
NAND3_X1 U905 ( .A1(n1042), .A2(n1228), .A3(KEYINPUT34), .ZN(n1232) );
XOR2_X1 U906 ( .A(n1234), .B(n1176), .Z(G21) );
NAND3_X1 U907 ( .A1(n1202), .A2(n1044), .A3(n1231), .ZN(n1176) );
XOR2_X1 U908 ( .A(n1235), .B(n1181), .Z(G18) );
NAND3_X1 U909 ( .A1(n1183), .A2(n1050), .A3(n1231), .ZN(n1181) );
INV_X1 U910 ( .A(n1054), .ZN(n1183) );
NAND2_X1 U911 ( .A1(n1198), .A2(n1236), .ZN(n1054) );
XNOR2_X1 U912 ( .A(G113), .B(n1180), .ZN(G15) );
NAND3_X1 U913 ( .A1(n1231), .A2(n1050), .A3(n1185), .ZN(n1180) );
NOR2_X1 U914 ( .A1(n1236), .A2(n1198), .ZN(n1185) );
INV_X1 U915 ( .A(n1195), .ZN(n1236) );
INV_X1 U916 ( .A(n1172), .ZN(n1050) );
NAND2_X1 U917 ( .A1(n1202), .A2(n1228), .ZN(n1172) );
INV_X1 U918 ( .A(n1210), .ZN(n1228) );
NOR2_X1 U919 ( .A1(n1041), .A2(n1237), .ZN(n1231) );
NAND2_X1 U920 ( .A1(n1065), .A2(n1238), .ZN(n1041) );
XNOR2_X1 U921 ( .A(G110), .B(n1179), .ZN(G12) );
NAND3_X1 U922 ( .A1(n1182), .A2(n1042), .A3(n1044), .ZN(n1179) );
AND2_X1 U923 ( .A1(n1049), .A2(n1210), .ZN(n1044) );
XOR2_X1 U924 ( .A(n1024), .B(n1026), .Z(n1210) );
NAND2_X1 U925 ( .A1(n1239), .A2(n1240), .ZN(n1026) );
XOR2_X1 U926 ( .A(KEYINPUT35), .B(G217), .Z(n1239) );
NAND2_X1 U927 ( .A1(n1241), .A2(n1109), .ZN(n1024) );
XNOR2_X1 U928 ( .A(n1242), .B(n1243), .ZN(n1109) );
XOR2_X1 U929 ( .A(n1244), .B(n1245), .Z(n1242) );
XOR2_X1 U930 ( .A(n1246), .B(n1247), .Z(n1245) );
XNOR2_X1 U931 ( .A(n1248), .B(n1249), .ZN(n1247) );
AND4_X1 U932 ( .A1(n1250), .A2(n1011), .A3(G234), .A4(G221), .ZN(n1249) );
INV_X1 U933 ( .A(KEYINPUT25), .ZN(n1250) );
NAND2_X1 U934 ( .A1(KEYINPUT58), .A2(n1251), .ZN(n1248) );
XOR2_X1 U935 ( .A(G119), .B(G110), .Z(n1246) );
XOR2_X1 U936 ( .A(n1252), .B(n1253), .Z(n1244) );
XOR2_X1 U937 ( .A(G137), .B(G128), .Z(n1253) );
XNOR2_X1 U938 ( .A(KEYINPUT47), .B(KEYINPUT29), .ZN(n1252) );
XNOR2_X1 U939 ( .A(n1254), .B(KEYINPUT55), .ZN(n1241) );
NOR2_X1 U940 ( .A1(n1198), .A2(n1195), .ZN(n1049) );
XNOR2_X1 U941 ( .A(n1019), .B(KEYINPUT5), .ZN(n1195) );
XNOR2_X1 U942 ( .A(n1255), .B(G475), .ZN(n1019) );
OR2_X1 U943 ( .A1(n1119), .A2(n1254), .ZN(n1255) );
XNOR2_X1 U944 ( .A(n1256), .B(n1257), .ZN(n1119) );
XNOR2_X1 U945 ( .A(n1258), .B(n1259), .ZN(n1257) );
XOR2_X1 U946 ( .A(n1260), .B(n1261), .Z(n1259) );
NOR2_X1 U947 ( .A1(KEYINPUT21), .A2(n1262), .ZN(n1261) );
XOR2_X1 U948 ( .A(G146), .B(n1243), .Z(n1262) );
INV_X1 U949 ( .A(n1083), .ZN(n1243) );
XOR2_X1 U950 ( .A(n1152), .B(n1191), .Z(n1083) );
NAND2_X1 U951 ( .A1(G214), .A2(n1263), .ZN(n1260) );
XOR2_X1 U952 ( .A(n1264), .B(n1265), .Z(n1256) );
XOR2_X1 U953 ( .A(G131), .B(G122), .Z(n1265) );
XNOR2_X1 U954 ( .A(G104), .B(G113), .ZN(n1264) );
XOR2_X1 U955 ( .A(n1266), .B(n1030), .Z(n1198) );
NOR2_X1 U956 ( .A1(n1114), .A2(n1254), .ZN(n1030) );
INV_X1 U957 ( .A(n1267), .ZN(n1254) );
XNOR2_X1 U958 ( .A(n1268), .B(n1269), .ZN(n1114) );
XOR2_X1 U959 ( .A(n1270), .B(n1271), .Z(n1269) );
NAND3_X1 U960 ( .A1(G217), .A2(n1011), .A3(G234), .ZN(n1271) );
NAND2_X1 U961 ( .A1(KEYINPUT26), .A2(n1272), .ZN(n1270) );
XOR2_X1 U962 ( .A(n1273), .B(n1274), .Z(n1272) );
XOR2_X1 U963 ( .A(n1275), .B(G116), .Z(n1274) );
NAND2_X1 U964 ( .A1(KEYINPUT51), .A2(n1006), .ZN(n1275) );
INV_X1 U965 ( .A(G107), .ZN(n1006) );
XOR2_X1 U966 ( .A(n1230), .B(KEYINPUT62), .Z(n1273) );
XOR2_X1 U967 ( .A(n1276), .B(G134), .Z(n1268) );
NAND2_X1 U968 ( .A1(KEYINPUT39), .A2(n1277), .ZN(n1276) );
NAND2_X1 U969 ( .A1(KEYINPUT60), .A2(n1031), .ZN(n1266) );
INV_X1 U970 ( .A(G478), .ZN(n1031) );
INV_X1 U971 ( .A(n1202), .ZN(n1042) );
XNOR2_X1 U972 ( .A(n1021), .B(n1278), .ZN(n1202) );
NOR2_X1 U973 ( .A1(G472), .A2(KEYINPUT28), .ZN(n1278) );
AND2_X1 U974 ( .A1(n1267), .A2(n1279), .ZN(n1021) );
XOR2_X1 U975 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U976 ( .A(n1135), .B(n1082), .ZN(n1281) );
XOR2_X1 U977 ( .A(n1282), .B(n1132), .Z(n1082) );
XNOR2_X1 U978 ( .A(n1283), .B(n1284), .ZN(n1135) );
NOR2_X1 U979 ( .A1(KEYINPUT48), .A2(n1285), .ZN(n1284) );
XOR2_X1 U980 ( .A(n1235), .B(KEYINPUT31), .Z(n1285) );
INV_X1 U981 ( .A(G116), .ZN(n1235) );
XOR2_X1 U982 ( .A(G113), .B(n1234), .Z(n1283) );
INV_X1 U983 ( .A(G119), .ZN(n1234) );
XOR2_X1 U984 ( .A(n1286), .B(KEYINPUT37), .Z(n1280) );
NAND2_X1 U985 ( .A1(n1287), .A2(n1138), .ZN(n1286) );
NAND3_X1 U986 ( .A1(G101), .A2(n1263), .A3(G210), .ZN(n1138) );
NAND2_X1 U987 ( .A1(n1288), .A2(n1140), .ZN(n1287) );
NAND2_X1 U988 ( .A1(G210), .A2(n1263), .ZN(n1140) );
NOR2_X1 U989 ( .A1(G953), .A2(G237), .ZN(n1263) );
XOR2_X1 U990 ( .A(KEYINPUT43), .B(G101), .Z(n1288) );
NOR2_X1 U991 ( .A1(n1237), .A2(n1170), .ZN(n1182) );
XOR2_X1 U992 ( .A(n1063), .B(KEYINPUT9), .Z(n1170) );
INV_X1 U993 ( .A(n1203), .ZN(n1063) );
NOR2_X1 U994 ( .A1(n1065), .A2(n1017), .ZN(n1203) );
INV_X1 U995 ( .A(n1238), .ZN(n1017) );
NAND2_X1 U996 ( .A1(G221), .A2(n1240), .ZN(n1238) );
NAND2_X1 U997 ( .A1(G234), .A2(n1160), .ZN(n1240) );
XOR2_X1 U998 ( .A(n1029), .B(G469), .Z(n1065) );
NAND2_X1 U999 ( .A1(n1289), .A2(n1267), .ZN(n1029) );
XOR2_X1 U1000 ( .A(n1290), .B(n1136), .Z(n1289) );
INV_X1 U1001 ( .A(n1282), .ZN(n1136) );
XNOR2_X1 U1002 ( .A(G131), .B(n1291), .ZN(n1282) );
XOR2_X1 U1003 ( .A(G137), .B(G134), .Z(n1291) );
XNOR2_X1 U1004 ( .A(n1292), .B(n1293), .ZN(n1290) );
NAND2_X1 U1005 ( .A1(n1294), .A2(KEYINPUT14), .ZN(n1293) );
XOR2_X1 U1006 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1007 ( .A(G110), .B(n1153), .Z(n1296) );
NOR2_X1 U1008 ( .A1(n1076), .A2(G953), .ZN(n1153) );
INV_X1 U1009 ( .A(G227), .ZN(n1076) );
NAND2_X1 U1010 ( .A1(KEYINPUT8), .A2(n1152), .ZN(n1295) );
INV_X1 U1011 ( .A(G140), .ZN(n1152) );
NAND2_X1 U1012 ( .A1(KEYINPUT63), .A2(n1297), .ZN(n1292) );
XOR2_X1 U1013 ( .A(n1187), .B(n1147), .Z(n1297) );
XNOR2_X1 U1014 ( .A(n1298), .B(n1299), .ZN(n1147) );
XNOR2_X1 U1015 ( .A(KEYINPUT44), .B(n1300), .ZN(n1298) );
NOR2_X1 U1016 ( .A1(KEYINPUT11), .A2(n1301), .ZN(n1300) );
XOR2_X1 U1017 ( .A(KEYINPUT23), .B(G101), .Z(n1301) );
INV_X1 U1018 ( .A(n1132), .ZN(n1187) );
NAND2_X1 U1019 ( .A1(n1058), .A2(n1302), .ZN(n1237) );
NAND2_X1 U1020 ( .A1(n1066), .A2(n1303), .ZN(n1302) );
NAND4_X1 U1021 ( .A1(G953), .A2(G902), .A3(n1227), .A4(n1103), .ZN(n1303) );
INV_X1 U1022 ( .A(G898), .ZN(n1103) );
NAND3_X1 U1023 ( .A1(n1227), .A2(n1011), .A3(G952), .ZN(n1066) );
NAND2_X1 U1024 ( .A1(G237), .A2(G234), .ZN(n1227) );
AND2_X1 U1025 ( .A1(n1036), .A2(n1022), .ZN(n1058) );
INV_X1 U1026 ( .A(n1037), .ZN(n1022) );
XNOR2_X1 U1027 ( .A(n1304), .B(n1159), .ZN(n1037) );
NAND2_X1 U1028 ( .A1(G210), .A2(n1305), .ZN(n1159) );
NAND2_X1 U1029 ( .A1(n1267), .A2(n1306), .ZN(n1304) );
XOR2_X1 U1030 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U1031 ( .A(n1191), .B(n1156), .ZN(n1308) );
XOR2_X1 U1032 ( .A(n1309), .B(n1100), .Z(n1156) );
NAND3_X1 U1033 ( .A1(n1310), .A2(n1311), .A3(n1312), .ZN(n1100) );
NAND2_X1 U1034 ( .A1(KEYINPUT12), .A2(G110), .ZN(n1312) );
NAND3_X1 U1035 ( .A1(n1313), .A2(n1314), .A3(n1230), .ZN(n1311) );
INV_X1 U1036 ( .A(KEYINPUT12), .ZN(n1314) );
OR2_X1 U1037 ( .A1(n1230), .A2(n1313), .ZN(n1310) );
NOR2_X1 U1038 ( .A1(G110), .A2(KEYINPUT6), .ZN(n1313) );
INV_X1 U1039 ( .A(G122), .ZN(n1230) );
NAND2_X1 U1040 ( .A1(n1315), .A2(n1105), .ZN(n1309) );
NAND2_X1 U1041 ( .A1(n1316), .A2(n1317), .ZN(n1105) );
XOR2_X1 U1042 ( .A(G101), .B(n1299), .Z(n1317) );
XNOR2_X1 U1043 ( .A(G113), .B(n1318), .ZN(n1316) );
XOR2_X1 U1044 ( .A(n1104), .B(KEYINPUT53), .Z(n1315) );
NAND2_X1 U1045 ( .A1(n1319), .A2(n1320), .ZN(n1104) );
XOR2_X1 U1046 ( .A(n1141), .B(n1299), .Z(n1320) );
XOR2_X1 U1047 ( .A(G104), .B(G107), .Z(n1299) );
INV_X1 U1048 ( .A(G101), .ZN(n1141) );
XOR2_X1 U1049 ( .A(n1318), .B(G113), .Z(n1319) );
NAND2_X1 U1050 ( .A1(KEYINPUT24), .A2(n1321), .ZN(n1318) );
XOR2_X1 U1051 ( .A(G119), .B(G116), .Z(n1321) );
XOR2_X1 U1052 ( .A(G125), .B(KEYINPUT1), .Z(n1191) );
XOR2_X1 U1053 ( .A(n1192), .B(n1132), .Z(n1307) );
XOR2_X1 U1054 ( .A(n1251), .B(n1277), .Z(n1132) );
XOR2_X1 U1055 ( .A(G128), .B(n1258), .Z(n1277) );
XOR2_X1 U1056 ( .A(G143), .B(KEYINPUT56), .Z(n1258) );
INV_X1 U1057 ( .A(G146), .ZN(n1251) );
AND2_X1 U1058 ( .A1(G224), .A2(n1011), .ZN(n1192) );
INV_X1 U1059 ( .A(G953), .ZN(n1011) );
XOR2_X1 U1060 ( .A(n1160), .B(KEYINPUT30), .Z(n1267) );
XNOR2_X1 U1061 ( .A(n1016), .B(KEYINPUT38), .ZN(n1036) );
AND2_X1 U1062 ( .A1(G214), .A2(n1305), .ZN(n1016) );
NAND2_X1 U1063 ( .A1(n1322), .A2(n1160), .ZN(n1305) );
INV_X1 U1064 ( .A(G902), .ZN(n1160) );
INV_X1 U1065 ( .A(G237), .ZN(n1322) );
endmodule


