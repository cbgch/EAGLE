//Key = 0000011110001001100000000011010111010000100001011000100100101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
n1440, n1441, n1442;

XNOR2_X1 U794 ( .A(G107), .B(n1090), .ZN(G9) );
NAND3_X1 U795 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
NOR2_X1 U796 ( .A1(n1094), .A2(n1095), .ZN(G75) );
NOR4_X1 U797 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1095) );
NOR2_X1 U798 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NOR3_X1 U799 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1100) );
NOR2_X1 U800 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NOR2_X1 U801 ( .A1(n1107), .A2(n1108), .ZN(n1103) );
XOR2_X1 U802 ( .A(KEYINPUT32), .B(n1109), .Z(n1108) );
INV_X1 U803 ( .A(n1110), .ZN(n1107) );
NOR2_X1 U804 ( .A1(n1111), .A2(n1112), .ZN(n1102) );
XOR2_X1 U805 ( .A(KEYINPUT49), .B(n1113), .Z(n1097) );
NOR4_X1 U806 ( .A1(n1112), .A2(n1114), .A3(n1101), .A4(n1115), .ZN(n1113) );
OR3_X1 U807 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1101) );
NAND3_X1 U808 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1096) );
NAND4_X1 U809 ( .A1(n1122), .A2(n1109), .A3(n1123), .A4(n1124), .ZN(n1121) );
NAND2_X1 U810 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND3_X1 U811 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1126) );
NAND3_X1 U812 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1128) );
NAND2_X1 U813 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
OR2_X1 U814 ( .A1(n1117), .A2(KEYINPUT16), .ZN(n1130) );
NAND3_X1 U815 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1127) );
NAND2_X1 U816 ( .A1(KEYINPUT24), .A2(n1133), .ZN(n1136) );
NAND2_X1 U817 ( .A1(n1138), .A2(n1139), .ZN(n1133) );
NAND2_X1 U818 ( .A1(KEYINPUT16), .A2(n1091), .ZN(n1135) );
NAND2_X1 U819 ( .A1(n1091), .A2(n1140), .ZN(n1125) );
INV_X1 U820 ( .A(n1118), .ZN(n1122) );
NOR3_X1 U821 ( .A1(n1141), .A2(G953), .A3(G952), .ZN(n1094) );
INV_X1 U822 ( .A(n1119), .ZN(n1141) );
NAND4_X1 U823 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1119) );
NOR4_X1 U824 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1145) );
NOR2_X1 U825 ( .A1(G478), .A2(n1150), .ZN(n1149) );
NOR3_X1 U826 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
NOR2_X1 U827 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NOR2_X1 U828 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NOR2_X1 U829 ( .A1(KEYINPUT53), .A2(KEYINPUT45), .ZN(n1156) );
NOR2_X1 U830 ( .A1(n1157), .A2(n1158), .ZN(n1152) );
INV_X1 U831 ( .A(KEYINPUT47), .ZN(n1157) );
AND2_X1 U832 ( .A1(KEYINPUT45), .A2(KEYINPUT53), .ZN(n1151) );
NOR4_X1 U833 ( .A1(n1159), .A2(n1160), .A3(KEYINPUT53), .A4(n1154), .ZN(n1148) );
NAND3_X1 U834 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1146) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(n1162) );
NAND2_X1 U836 ( .A1(KEYINPUT35), .A2(n1166), .ZN(n1165) );
NAND2_X1 U837 ( .A1(KEYINPUT53), .A2(n1167), .ZN(n1161) );
NAND2_X1 U838 ( .A1(n1158), .A2(n1168), .ZN(n1167) );
NAND2_X1 U839 ( .A1(G478), .A2(n1160), .ZN(n1168) );
INV_X1 U840 ( .A(KEYINPUT45), .ZN(n1160) );
NOR3_X1 U841 ( .A1(n1169), .A2(n1170), .A3(n1137), .ZN(n1144) );
INV_X1 U842 ( .A(n1115), .ZN(n1169) );
NAND2_X1 U843 ( .A1(n1171), .A2(n1172), .ZN(n1143) );
XOR2_X1 U844 ( .A(KEYINPUT22), .B(n1173), .Z(n1171) );
XOR2_X1 U845 ( .A(n1174), .B(n1175), .Z(n1142) );
XOR2_X1 U846 ( .A(KEYINPUT42), .B(n1176), .Z(n1175) );
NOR2_X1 U847 ( .A1(KEYINPUT1), .A2(n1177), .ZN(n1174) );
INV_X1 U848 ( .A(n1178), .ZN(n1177) );
NAND3_X1 U849 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(G72) );
OR2_X1 U850 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND2_X1 U851 ( .A1(n1184), .A2(n1185), .ZN(n1180) );
INV_X1 U852 ( .A(KEYINPUT48), .ZN(n1185) );
NAND2_X1 U853 ( .A1(n1186), .A2(n1183), .ZN(n1184) );
XNOR2_X1 U854 ( .A(KEYINPUT5), .B(n1182), .ZN(n1186) );
NAND2_X1 U855 ( .A1(KEYINPUT48), .A2(n1187), .ZN(n1179) );
NAND2_X1 U856 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NAND3_X1 U857 ( .A1(KEYINPUT5), .A2(n1183), .A3(n1182), .ZN(n1189) );
XNOR2_X1 U858 ( .A(n1190), .B(n1191), .ZN(n1183) );
NOR2_X1 U859 ( .A1(n1192), .A2(G953), .ZN(n1191) );
NOR3_X1 U860 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1192) );
NAND2_X1 U861 ( .A1(n1196), .A2(n1197), .ZN(n1190) );
NAND2_X1 U862 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U863 ( .A(n1200), .B(n1201), .Z(n1196) );
XOR2_X1 U864 ( .A(G128), .B(G125), .Z(n1201) );
XOR2_X1 U865 ( .A(n1202), .B(n1203), .Z(n1200) );
NAND2_X1 U866 ( .A1(n1204), .A2(KEYINPUT33), .ZN(n1202) );
XNOR2_X1 U867 ( .A(G134), .B(n1205), .ZN(n1204) );
NOR2_X1 U868 ( .A1(G137), .A2(KEYINPUT56), .ZN(n1205) );
OR2_X1 U869 ( .A1(n1182), .A2(KEYINPUT5), .ZN(n1188) );
NAND2_X1 U870 ( .A1(G953), .A2(n1206), .ZN(n1182) );
NAND2_X1 U871 ( .A1(G900), .A2(G227), .ZN(n1206) );
XOR2_X1 U872 ( .A(n1207), .B(n1208), .Z(G69) );
NOR2_X1 U873 ( .A1(n1209), .A2(n1120), .ZN(n1208) );
NOR2_X1 U874 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND2_X1 U875 ( .A1(n1212), .A2(KEYINPUT40), .ZN(n1207) );
XOR2_X1 U876 ( .A(n1213), .B(n1214), .Z(n1212) );
NOR3_X1 U877 ( .A1(n1215), .A2(KEYINPUT18), .A3(G953), .ZN(n1214) );
NAND2_X1 U878 ( .A1(n1216), .A2(n1217), .ZN(n1213) );
NAND2_X1 U879 ( .A1(n1198), .A2(n1211), .ZN(n1217) );
XOR2_X1 U880 ( .A(n1218), .B(n1219), .Z(n1216) );
XNOR2_X1 U881 ( .A(n1220), .B(n1221), .ZN(n1219) );
NOR2_X1 U882 ( .A1(n1222), .A2(n1223), .ZN(G66) );
NOR2_X1 U883 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
XOR2_X1 U884 ( .A(n1226), .B(n1227), .Z(n1225) );
NOR2_X1 U885 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND2_X1 U886 ( .A1(n1230), .A2(n1231), .ZN(n1226) );
NOR2_X1 U887 ( .A1(n1230), .A2(n1231), .ZN(n1224) );
INV_X1 U888 ( .A(KEYINPUT30), .ZN(n1231) );
NOR2_X1 U889 ( .A1(n1222), .A2(n1232), .ZN(G63) );
NOR3_X1 U890 ( .A1(n1154), .A2(n1233), .A3(n1234), .ZN(n1232) );
NOR3_X1 U891 ( .A1(n1235), .A2(n1159), .A3(n1229), .ZN(n1234) );
NOR2_X1 U892 ( .A1(n1236), .A2(n1237), .ZN(n1233) );
INV_X1 U893 ( .A(n1235), .ZN(n1237) );
NOR2_X1 U894 ( .A1(n1238), .A2(n1159), .ZN(n1236) );
INV_X1 U895 ( .A(G478), .ZN(n1159) );
INV_X1 U896 ( .A(n1158), .ZN(n1154) );
NOR2_X1 U897 ( .A1(n1222), .A2(n1239), .ZN(G60) );
XOR2_X1 U898 ( .A(n1240), .B(n1241), .Z(n1239) );
NOR2_X1 U899 ( .A1(n1242), .A2(n1229), .ZN(n1241) );
XOR2_X1 U900 ( .A(n1243), .B(n1244), .Z(G6) );
XOR2_X1 U901 ( .A(n1245), .B(KEYINPUT2), .Z(n1244) );
NOR2_X1 U902 ( .A1(n1222), .A2(n1246), .ZN(G57) );
XOR2_X1 U903 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U904 ( .A(n1249), .B(n1250), .Z(n1248) );
XOR2_X1 U905 ( .A(KEYINPUT58), .B(n1251), .Z(n1247) );
NOR2_X1 U906 ( .A1(n1252), .A2(n1229), .ZN(n1251) );
INV_X1 U907 ( .A(G472), .ZN(n1252) );
NOR2_X1 U908 ( .A1(n1222), .A2(n1253), .ZN(G54) );
XOR2_X1 U909 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U910 ( .A(KEYINPUT11), .B(n1256), .Z(n1255) );
NOR2_X1 U911 ( .A1(n1166), .A2(n1229), .ZN(n1256) );
INV_X1 U912 ( .A(G469), .ZN(n1166) );
NOR2_X1 U913 ( .A1(n1222), .A2(n1257), .ZN(G51) );
NOR3_X1 U914 ( .A1(n1176), .A2(n1258), .A3(n1259), .ZN(n1257) );
NOR4_X1 U915 ( .A1(n1260), .A2(n1261), .A3(n1178), .A4(n1229), .ZN(n1259) );
NAND2_X1 U916 ( .A1(G902), .A2(n1099), .ZN(n1229) );
NOR2_X1 U917 ( .A1(n1262), .A2(n1263), .ZN(n1258) );
NOR3_X1 U918 ( .A1(n1261), .A2(n1238), .A3(n1178), .ZN(n1262) );
INV_X1 U919 ( .A(n1099), .ZN(n1238) );
NAND4_X1 U920 ( .A1(n1264), .A2(n1215), .A3(n1265), .A4(n1266), .ZN(n1099) );
XOR2_X1 U921 ( .A(KEYINPUT55), .B(n1194), .Z(n1266) );
INV_X1 U922 ( .A(n1193), .ZN(n1265) );
NAND3_X1 U923 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(n1193) );
AND2_X1 U924 ( .A1(n1270), .A2(n1271), .ZN(n1215) );
AND4_X1 U925 ( .A1(n1272), .A2(n1273), .A3(n1274), .A4(n1243), .ZN(n1271) );
NAND3_X1 U926 ( .A1(n1091), .A2(n1092), .A3(n1110), .ZN(n1243) );
OR4_X1 U927 ( .A1(n1275), .A2(n1117), .A3(n1105), .A4(n1276), .ZN(n1274) );
XOR2_X1 U928 ( .A(KEYINPUT59), .B(n1277), .Z(n1276) );
NOR4_X1 U929 ( .A1(n1278), .A2(n1279), .A3(n1280), .A4(n1281), .ZN(n1270) );
NOR3_X1 U930 ( .A1(n1282), .A2(n1112), .A3(n1283), .ZN(n1281) );
INV_X1 U931 ( .A(n1284), .ZN(n1280) );
NOR3_X1 U932 ( .A1(n1285), .A2(n1277), .A3(n1138), .ZN(n1278) );
NAND3_X1 U933 ( .A1(n1286), .A2(n1287), .A3(n1123), .ZN(n1285) );
OR2_X1 U934 ( .A1(n1288), .A2(KEYINPUT36), .ZN(n1287) );
NAND2_X1 U935 ( .A1(KEYINPUT36), .A2(n1289), .ZN(n1286) );
NAND2_X1 U936 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
XOR2_X1 U937 ( .A(n1195), .B(KEYINPUT8), .Z(n1264) );
NAND4_X1 U938 ( .A1(n1292), .A2(n1293), .A3(n1294), .A4(n1295), .ZN(n1195) );
NAND3_X1 U939 ( .A1(n1296), .A2(n1297), .A3(n1298), .ZN(n1293) );
INV_X1 U940 ( .A(KEYINPUT54), .ZN(n1297) );
NAND2_X1 U941 ( .A1(n1299), .A2(n1300), .ZN(n1292) );
NAND2_X1 U942 ( .A1(n1301), .A2(n1302), .ZN(n1299) );
NAND4_X1 U943 ( .A1(KEYINPUT54), .A2(n1296), .A3(n1290), .A4(n1116), .ZN(n1302) );
NAND3_X1 U944 ( .A1(n1093), .A2(n1288), .A3(n1303), .ZN(n1301) );
INV_X1 U945 ( .A(KEYINPUT63), .ZN(n1261) );
NOR2_X1 U946 ( .A1(n1120), .A2(G952), .ZN(n1222) );
XNOR2_X1 U947 ( .A(G146), .B(n1269), .ZN(G48) );
NAND4_X1 U948 ( .A1(n1303), .A2(n1110), .A3(n1288), .A4(n1300), .ZN(n1269) );
INV_X1 U949 ( .A(n1275), .ZN(n1288) );
XOR2_X1 U950 ( .A(n1304), .B(G143), .Z(G45) );
NAND2_X1 U951 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
OR2_X1 U952 ( .A1(n1268), .A2(KEYINPUT14), .ZN(n1306) );
NAND2_X1 U953 ( .A1(n1307), .A2(n1308), .ZN(n1268) );
NAND3_X1 U954 ( .A1(n1307), .A2(n1138), .A3(KEYINPUT14), .ZN(n1305) );
NOR4_X1 U955 ( .A1(n1275), .A2(n1309), .A3(n1310), .A4(n1311), .ZN(n1307) );
XOR2_X1 U956 ( .A(G140), .B(n1194), .Z(G42) );
AND3_X1 U957 ( .A1(n1110), .A2(n1312), .A3(n1298), .ZN(n1194) );
XNOR2_X1 U958 ( .A(G137), .B(n1267), .ZN(G39) );
NAND3_X1 U959 ( .A1(n1303), .A2(n1123), .A3(n1298), .ZN(n1267) );
XNOR2_X1 U960 ( .A(G134), .B(n1313), .ZN(G36) );
NAND2_X1 U961 ( .A1(n1298), .A2(n1296), .ZN(n1313) );
XNOR2_X1 U962 ( .A(G131), .B(n1294), .ZN(G33) );
NAND3_X1 U963 ( .A1(n1110), .A2(n1308), .A3(n1298), .ZN(n1294) );
NOR3_X1 U964 ( .A1(n1111), .A2(n1310), .A3(n1116), .ZN(n1298) );
NAND2_X1 U965 ( .A1(n1314), .A2(n1129), .ZN(n1116) );
XOR2_X1 U966 ( .A(n1134), .B(n1137), .Z(n1314) );
INV_X1 U967 ( .A(KEYINPUT24), .ZN(n1134) );
NAND2_X1 U968 ( .A1(n1315), .A2(n1316), .ZN(G30) );
NAND2_X1 U969 ( .A1(G128), .A2(n1317), .ZN(n1316) );
XOR2_X1 U970 ( .A(n1318), .B(KEYINPUT39), .Z(n1315) );
OR2_X1 U971 ( .A1(n1317), .A2(G128), .ZN(n1318) );
NAND4_X1 U972 ( .A1(n1319), .A2(n1303), .A3(n1320), .A4(n1093), .ZN(n1317) );
INV_X1 U973 ( .A(n1105), .ZN(n1093) );
NOR2_X1 U974 ( .A1(n1321), .A2(n1111), .ZN(n1320) );
XOR2_X1 U975 ( .A(n1291), .B(KEYINPUT19), .Z(n1321) );
XOR2_X1 U976 ( .A(n1300), .B(KEYINPUT38), .Z(n1319) );
NAND2_X1 U977 ( .A1(n1322), .A2(n1323), .ZN(G3) );
NAND2_X1 U978 ( .A1(G101), .A2(n1324), .ZN(n1323) );
XOR2_X1 U979 ( .A(n1325), .B(KEYINPUT37), .Z(n1322) );
OR2_X1 U980 ( .A1(n1324), .A2(G101), .ZN(n1325) );
NAND3_X1 U981 ( .A1(n1092), .A2(n1308), .A3(n1123), .ZN(n1324) );
NAND2_X1 U982 ( .A1(n1326), .A2(n1327), .ZN(G27) );
NAND2_X1 U983 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
XOR2_X1 U984 ( .A(KEYINPUT27), .B(n1330), .Z(n1326) );
NOR2_X1 U985 ( .A1(n1328), .A2(n1329), .ZN(n1330) );
INV_X1 U986 ( .A(n1295), .ZN(n1328) );
NAND4_X1 U987 ( .A1(n1110), .A2(n1109), .A3(n1331), .A4(n1312), .ZN(n1295) );
NOR2_X1 U988 ( .A1(n1310), .A2(n1291), .ZN(n1331) );
INV_X1 U989 ( .A(n1140), .ZN(n1291) );
INV_X1 U990 ( .A(n1300), .ZN(n1310) );
NAND2_X1 U991 ( .A1(n1118), .A2(n1332), .ZN(n1300) );
NAND2_X1 U992 ( .A1(n1333), .A2(n1199), .ZN(n1332) );
INV_X1 U993 ( .A(G900), .ZN(n1199) );
XOR2_X1 U994 ( .A(n1334), .B(n1273), .Z(G24) );
OR4_X1 U995 ( .A1(n1283), .A2(n1117), .A3(n1309), .A4(n1311), .ZN(n1273) );
INV_X1 U996 ( .A(n1091), .ZN(n1117) );
XNOR2_X1 U997 ( .A(G119), .B(n1335), .ZN(G21) );
NAND3_X1 U998 ( .A1(n1303), .A2(n1336), .A3(n1337), .ZN(n1335) );
XOR2_X1 U999 ( .A(n1112), .B(KEYINPUT29), .Z(n1337) );
INV_X1 U1000 ( .A(n1282), .ZN(n1303) );
NAND2_X1 U1001 ( .A1(n1338), .A2(n1147), .ZN(n1282) );
XOR2_X1 U1002 ( .A(n1339), .B(n1284), .Z(G18) );
NAND2_X1 U1003 ( .A1(n1296), .A2(n1336), .ZN(n1284) );
NOR2_X1 U1004 ( .A1(n1105), .A2(n1138), .ZN(n1296) );
INV_X1 U1005 ( .A(n1308), .ZN(n1138) );
NAND2_X1 U1006 ( .A1(n1311), .A2(n1340), .ZN(n1105) );
NAND3_X1 U1007 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(G15) );
NAND2_X1 U1008 ( .A1(G113), .A2(n1344), .ZN(n1343) );
NAND2_X1 U1009 ( .A1(n1345), .A2(n1346), .ZN(n1342) );
INV_X1 U1010 ( .A(KEYINPUT26), .ZN(n1346) );
NAND2_X1 U1011 ( .A1(n1347), .A2(n1279), .ZN(n1345) );
INV_X1 U1012 ( .A(n1344), .ZN(n1279) );
XNOR2_X1 U1013 ( .A(KEYINPUT9), .B(G113), .ZN(n1347) );
NAND2_X1 U1014 ( .A1(KEYINPUT26), .A2(n1348), .ZN(n1341) );
NAND2_X1 U1015 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
OR3_X1 U1016 ( .A1(n1344), .A2(G113), .A3(KEYINPUT9), .ZN(n1350) );
NAND3_X1 U1017 ( .A1(n1336), .A2(n1308), .A3(n1110), .ZN(n1344) );
NOR2_X1 U1018 ( .A1(n1340), .A2(n1311), .ZN(n1110) );
NAND2_X1 U1019 ( .A1(n1351), .A2(n1352), .ZN(n1308) );
OR3_X1 U1020 ( .A1(n1147), .A2(n1353), .A3(KEYINPUT21), .ZN(n1352) );
NAND2_X1 U1021 ( .A1(KEYINPUT21), .A2(n1091), .ZN(n1351) );
NOR2_X1 U1022 ( .A1(n1147), .A2(n1338), .ZN(n1091) );
INV_X1 U1023 ( .A(n1283), .ZN(n1336) );
NAND3_X1 U1024 ( .A1(n1140), .A2(n1354), .A3(n1109), .ZN(n1283) );
INV_X1 U1025 ( .A(n1106), .ZN(n1109) );
NAND2_X1 U1026 ( .A1(n1355), .A2(n1115), .ZN(n1106) );
NAND2_X1 U1027 ( .A1(KEYINPUT9), .A2(G113), .ZN(n1349) );
XNOR2_X1 U1028 ( .A(G110), .B(n1272), .ZN(G12) );
NAND3_X1 U1029 ( .A1(n1312), .A2(n1092), .A3(n1123), .ZN(n1272) );
INV_X1 U1030 ( .A(n1112), .ZN(n1123) );
NAND2_X1 U1031 ( .A1(n1309), .A2(n1311), .ZN(n1112) );
NOR2_X1 U1032 ( .A1(n1356), .A2(n1170), .ZN(n1311) );
NOR2_X1 U1033 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
AND2_X1 U1034 ( .A1(n1173), .A2(n1172), .ZN(n1356) );
NAND2_X1 U1035 ( .A1(n1357), .A2(n1358), .ZN(n1172) );
XOR2_X1 U1036 ( .A(KEYINPUT23), .B(n1359), .Z(n1357) );
INV_X1 U1037 ( .A(n1240), .ZN(n1359) );
XOR2_X1 U1038 ( .A(n1360), .B(n1361), .Z(n1240) );
XOR2_X1 U1039 ( .A(n1362), .B(n1363), .Z(n1361) );
XOR2_X1 U1040 ( .A(n1364), .B(G122), .Z(n1363) );
NAND2_X1 U1041 ( .A1(G214), .A2(n1365), .ZN(n1364) );
XNOR2_X1 U1042 ( .A(KEYINPUT43), .B(KEYINPUT60), .ZN(n1362) );
XOR2_X1 U1043 ( .A(n1366), .B(n1367), .Z(n1360) );
XOR2_X1 U1044 ( .A(n1368), .B(n1369), .Z(n1367) );
NAND2_X1 U1045 ( .A1(KEYINPUT6), .A2(n1245), .ZN(n1368) );
INV_X1 U1046 ( .A(G104), .ZN(n1245) );
XNOR2_X1 U1047 ( .A(n1242), .B(KEYINPUT57), .ZN(n1173) );
INV_X1 U1048 ( .A(G475), .ZN(n1242) );
INV_X1 U1049 ( .A(n1340), .ZN(n1309) );
XNOR2_X1 U1050 ( .A(n1158), .B(G478), .ZN(n1340) );
NAND2_X1 U1051 ( .A1(n1235), .A2(n1358), .ZN(n1158) );
XOR2_X1 U1052 ( .A(n1370), .B(n1371), .Z(n1235) );
XOR2_X1 U1053 ( .A(n1372), .B(n1373), .Z(n1371) );
XNOR2_X1 U1054 ( .A(n1374), .B(n1375), .ZN(n1373) );
NOR2_X1 U1055 ( .A1(G134), .A2(KEYINPUT3), .ZN(n1375) );
NOR3_X1 U1056 ( .A1(KEYINPUT17), .A2(n1376), .A3(n1377), .ZN(n1374) );
AND3_X1 U1057 ( .A1(KEYINPUT41), .A2(n1339), .A3(G122), .ZN(n1377) );
NOR2_X1 U1058 ( .A1(KEYINPUT41), .A2(n1378), .ZN(n1376) );
XOR2_X1 U1059 ( .A(G122), .B(G116), .Z(n1378) );
NAND2_X1 U1060 ( .A1(G217), .A2(n1379), .ZN(n1372) );
XNOR2_X1 U1061 ( .A(G107), .B(n1380), .ZN(n1370) );
XOR2_X1 U1062 ( .A(G143), .B(G128), .Z(n1380) );
NOR2_X1 U1063 ( .A1(n1275), .A2(n1277), .ZN(n1092) );
INV_X1 U1064 ( .A(n1354), .ZN(n1277) );
NAND2_X1 U1065 ( .A1(n1118), .A2(n1381), .ZN(n1354) );
NAND2_X1 U1066 ( .A1(n1333), .A2(n1211), .ZN(n1381) );
INV_X1 U1067 ( .A(G898), .ZN(n1211) );
AND3_X1 U1068 ( .A1(n1198), .A2(n1382), .A3(G902), .ZN(n1333) );
XOR2_X1 U1069 ( .A(G953), .B(KEYINPUT25), .Z(n1198) );
NAND3_X1 U1070 ( .A1(n1382), .A2(n1120), .A3(G952), .ZN(n1118) );
NAND2_X1 U1071 ( .A1(G237), .A2(G234), .ZN(n1382) );
NAND2_X1 U1072 ( .A1(n1140), .A2(n1290), .ZN(n1275) );
INV_X1 U1073 ( .A(n1111), .ZN(n1290) );
NAND2_X1 U1074 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
NAND2_X1 U1075 ( .A1(G221), .A2(n1383), .ZN(n1115) );
INV_X1 U1076 ( .A(n1355), .ZN(n1114) );
XOR2_X1 U1077 ( .A(n1164), .B(G469), .Z(n1355) );
NAND2_X1 U1078 ( .A1(n1384), .A2(n1358), .ZN(n1164) );
XOR2_X1 U1079 ( .A(KEYINPUT10), .B(n1385), .Z(n1384) );
INV_X1 U1080 ( .A(n1254), .ZN(n1385) );
XOR2_X1 U1081 ( .A(n1386), .B(n1387), .Z(n1254) );
XOR2_X1 U1082 ( .A(n1388), .B(n1389), .Z(n1387) );
XOR2_X1 U1083 ( .A(G110), .B(n1390), .Z(n1389) );
NOR2_X1 U1084 ( .A1(KEYINPUT4), .A2(n1391), .ZN(n1390) );
XOR2_X1 U1085 ( .A(KEYINPUT0), .B(G101), .Z(n1391) );
AND2_X1 U1086 ( .A1(n1120), .A2(G227), .ZN(n1388) );
XOR2_X1 U1087 ( .A(n1392), .B(n1393), .Z(n1386) );
XNOR2_X1 U1088 ( .A(n1203), .B(n1394), .ZN(n1392) );
XNOR2_X1 U1089 ( .A(n1369), .B(n1395), .ZN(n1203) );
NOR2_X1 U1090 ( .A1(KEYINPUT20), .A2(n1396), .ZN(n1395) );
XNOR2_X1 U1091 ( .A(G131), .B(G140), .ZN(n1369) );
NOR2_X1 U1092 ( .A1(n1129), .A2(n1137), .ZN(n1140) );
INV_X1 U1093 ( .A(n1132), .ZN(n1137) );
NAND2_X1 U1094 ( .A1(G214), .A2(n1397), .ZN(n1132) );
XOR2_X1 U1095 ( .A(n1176), .B(n1178), .Z(n1129) );
NAND2_X1 U1096 ( .A1(G210), .A2(n1397), .ZN(n1178) );
NAND2_X1 U1097 ( .A1(n1358), .A2(n1398), .ZN(n1397) );
INV_X1 U1098 ( .A(G237), .ZN(n1398) );
NOR2_X1 U1099 ( .A1(n1263), .A2(G902), .ZN(n1176) );
INV_X1 U1100 ( .A(n1260), .ZN(n1263) );
XOR2_X1 U1101 ( .A(n1399), .B(n1400), .Z(n1260) );
XOR2_X1 U1102 ( .A(n1401), .B(n1402), .Z(n1400) );
XOR2_X1 U1103 ( .A(n1403), .B(n1404), .Z(n1402) );
NOR2_X1 U1104 ( .A1(G953), .A2(n1210), .ZN(n1404) );
INV_X1 U1105 ( .A(G224), .ZN(n1210) );
NAND2_X1 U1106 ( .A1(KEYINPUT31), .A2(n1220), .ZN(n1401) );
XOR2_X1 U1107 ( .A(n1334), .B(n1405), .Z(n1220) );
NOR2_X1 U1108 ( .A1(G110), .A2(KEYINPUT51), .ZN(n1405) );
INV_X1 U1109 ( .A(G122), .ZN(n1334) );
XOR2_X1 U1110 ( .A(n1366), .B(n1406), .Z(n1399) );
INV_X1 U1111 ( .A(n1218), .ZN(n1406) );
XOR2_X1 U1112 ( .A(n1407), .B(n1408), .Z(n1218) );
XOR2_X1 U1113 ( .A(G116), .B(n1409), .Z(n1408) );
XOR2_X1 U1114 ( .A(KEYINPUT7), .B(G119), .Z(n1409) );
XOR2_X1 U1115 ( .A(n1410), .B(n1393), .Z(n1407) );
XOR2_X1 U1116 ( .A(G104), .B(G107), .Z(n1393) );
INV_X1 U1117 ( .A(G101), .ZN(n1410) );
XOR2_X1 U1118 ( .A(n1329), .B(n1411), .Z(n1366) );
INV_X1 U1119 ( .A(n1139), .ZN(n1312) );
NAND2_X1 U1120 ( .A1(n1353), .A2(n1147), .ZN(n1139) );
XOR2_X1 U1121 ( .A(n1412), .B(n1228), .Z(n1147) );
NAND2_X1 U1122 ( .A1(G217), .A2(n1383), .ZN(n1228) );
NAND2_X1 U1123 ( .A1(n1413), .A2(n1358), .ZN(n1383) );
XNOR2_X1 U1124 ( .A(G234), .B(KEYINPUT15), .ZN(n1413) );
OR2_X1 U1125 ( .A1(n1230), .A2(G902), .ZN(n1412) );
XNOR2_X1 U1126 ( .A(n1414), .B(n1415), .ZN(n1230) );
XOR2_X1 U1127 ( .A(n1416), .B(n1417), .Z(n1415) );
XOR2_X1 U1128 ( .A(G137), .B(G110), .Z(n1417) );
NOR2_X1 U1129 ( .A1(KEYINPUT50), .A2(n1418), .ZN(n1416) );
XOR2_X1 U1130 ( .A(G128), .B(G119), .Z(n1418) );
XOR2_X1 U1131 ( .A(n1419), .B(n1420), .Z(n1414) );
AND2_X1 U1132 ( .A1(n1379), .A2(G221), .ZN(n1420) );
AND2_X1 U1133 ( .A1(G234), .A2(n1120), .ZN(n1379) );
INV_X1 U1134 ( .A(G953), .ZN(n1120) );
NAND3_X1 U1135 ( .A1(KEYINPUT12), .A2(n1421), .A3(n1422), .ZN(n1419) );
XOR2_X1 U1136 ( .A(n1423), .B(KEYINPUT44), .Z(n1422) );
NAND2_X1 U1137 ( .A1(n1424), .A2(n1425), .ZN(n1423) );
OR2_X1 U1138 ( .A1(n1425), .A2(n1424), .ZN(n1421) );
AND3_X1 U1139 ( .A1(n1426), .A2(n1427), .A3(n1428), .ZN(n1424) );
OR2_X1 U1140 ( .A1(n1429), .A2(KEYINPUT62), .ZN(n1428) );
NAND4_X1 U1141 ( .A1(n1429), .A2(n1430), .A3(KEYINPUT62), .A4(n1329), .ZN(n1427) );
INV_X1 U1142 ( .A(G125), .ZN(n1329) );
NAND2_X1 U1143 ( .A1(G125), .A2(n1431), .ZN(n1426) );
NAND2_X1 U1144 ( .A1(n1429), .A2(n1430), .ZN(n1431) );
INV_X1 U1145 ( .A(KEYINPUT46), .ZN(n1430) );
XOR2_X1 U1146 ( .A(G140), .B(KEYINPUT60), .Z(n1429) );
XOR2_X1 U1147 ( .A(G146), .B(KEYINPUT43), .Z(n1425) );
INV_X1 U1148 ( .A(n1338), .ZN(n1353) );
XOR2_X1 U1149 ( .A(n1163), .B(KEYINPUT52), .Z(n1338) );
XOR2_X1 U1150 ( .A(n1432), .B(G472), .Z(n1163) );
NAND2_X1 U1151 ( .A1(n1433), .A2(n1358), .ZN(n1432) );
INV_X1 U1152 ( .A(G902), .ZN(n1358) );
XOR2_X1 U1153 ( .A(n1434), .B(n1435), .Z(n1433) );
INV_X1 U1154 ( .A(n1249), .ZN(n1435) );
XOR2_X1 U1155 ( .A(n1436), .B(n1437), .Z(n1249) );
XOR2_X1 U1156 ( .A(n1394), .B(n1411), .Z(n1437) );
XNOR2_X1 U1157 ( .A(n1396), .B(n1221), .ZN(n1411) );
XOR2_X1 U1158 ( .A(G113), .B(KEYINPUT34), .Z(n1221) );
XNOR2_X1 U1159 ( .A(G143), .B(G146), .ZN(n1396) );
XNOR2_X1 U1160 ( .A(n1438), .B(n1439), .ZN(n1394) );
NOR2_X1 U1161 ( .A1(KEYINPUT28), .A2(G134), .ZN(n1439) );
XOR2_X1 U1162 ( .A(G137), .B(n1403), .Z(n1438) );
INV_X1 U1163 ( .A(G128), .ZN(n1403) );
XOR2_X1 U1164 ( .A(n1440), .B(n1441), .Z(n1436) );
NOR2_X1 U1165 ( .A1(KEYINPUT13), .A2(G119), .ZN(n1441) );
XOR2_X1 U1166 ( .A(G131), .B(n1339), .Z(n1440) );
INV_X1 U1167 ( .A(G116), .ZN(n1339) );
NOR2_X1 U1168 ( .A1(KEYINPUT61), .A2(n1250), .ZN(n1434) );
XOR2_X1 U1169 ( .A(n1442), .B(G101), .Z(n1250) );
NAND2_X1 U1170 ( .A1(G210), .A2(n1365), .ZN(n1442) );
NOR2_X1 U1171 ( .A1(G953), .A2(G237), .ZN(n1365) );
endmodule


