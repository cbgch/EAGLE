//Key = 0110111111001110111110111000010010011111111101001101010100100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295;

XOR2_X1 U709 ( .A(G107), .B(n978), .Z(G9) );
NOR2_X1 U710 ( .A1(n979), .A2(n980), .ZN(G75) );
NOR4_X1 U711 ( .A1(G953), .A2(n981), .A3(n982), .A4(n983), .ZN(n980) );
INV_X1 U712 ( .A(n984), .ZN(n983) );
NOR2_X1 U713 ( .A1(n985), .A2(n986), .ZN(n982) );
NOR2_X1 U714 ( .A1(n987), .A2(n988), .ZN(n985) );
NOR4_X1 U715 ( .A1(n989), .A2(n990), .A3(n991), .A4(n992), .ZN(n988) );
NOR4_X1 U716 ( .A1(n993), .A2(n994), .A3(n995), .A4(n996), .ZN(n990) );
NOR2_X1 U717 ( .A1(n997), .A2(n998), .ZN(n996) );
XNOR2_X1 U718 ( .A(KEYINPUT38), .B(n999), .ZN(n998) );
INV_X1 U719 ( .A(n1000), .ZN(n997) );
NOR2_X1 U720 ( .A1(n1001), .A2(n1002), .ZN(n995) );
NOR2_X1 U721 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
AND2_X1 U722 ( .A1(n1005), .A2(n1006), .ZN(n994) );
NOR2_X1 U723 ( .A1(n1007), .A2(n1008), .ZN(n989) );
NOR3_X1 U724 ( .A1(n999), .A2(n1009), .A3(n1002), .ZN(n1008) );
NOR2_X1 U725 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
INV_X1 U726 ( .A(n993), .ZN(n1007) );
NOR3_X1 U727 ( .A1(n999), .A2(n1012), .A3(n1002), .ZN(n987) );
INV_X1 U728 ( .A(n1013), .ZN(n1002) );
NOR2_X1 U729 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR3_X1 U730 ( .A1(n981), .A2(G953), .A3(G952), .ZN(n979) );
AND4_X1 U731 ( .A1(n1016), .A2(n1017), .A3(n1018), .A4(n1019), .ZN(n981) );
NOR4_X1 U732 ( .A1(n1020), .A2(n993), .A3(n1021), .A4(n1022), .ZN(n1019) );
XNOR2_X1 U733 ( .A(G475), .B(n1023), .ZN(n1022) );
XNOR2_X1 U734 ( .A(n1024), .B(n1025), .ZN(n1021) );
NOR2_X1 U735 ( .A1(KEYINPUT61), .A2(n1026), .ZN(n1025) );
INV_X1 U736 ( .A(G469), .ZN(n1026) );
XOR2_X1 U737 ( .A(n1027), .B(n1028), .Z(n1020) );
XNOR2_X1 U738 ( .A(KEYINPUT31), .B(n1029), .ZN(n1028) );
NAND2_X1 U739 ( .A1(n1030), .A2(n1031), .ZN(n1027) );
XNOR2_X1 U740 ( .A(KEYINPUT5), .B(KEYINPUT2), .ZN(n1030) );
NOR3_X1 U741 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1018) );
INV_X1 U742 ( .A(n1035), .ZN(n1032) );
NAND2_X1 U743 ( .A1(G478), .A2(n1036), .ZN(n1017) );
XNOR2_X1 U744 ( .A(KEYINPUT13), .B(n1037), .ZN(n1036) );
XOR2_X1 U745 ( .A(n1038), .B(n1039), .Z(n1016) );
NOR2_X1 U746 ( .A1(n1040), .A2(KEYINPUT30), .ZN(n1039) );
XOR2_X1 U747 ( .A(n1041), .B(n1042), .Z(G72) );
NOR2_X1 U748 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
AND2_X1 U749 ( .A1(G227), .A2(G900), .ZN(n1043) );
NAND2_X1 U750 ( .A1(n1045), .A2(n1046), .ZN(n1041) );
NAND2_X1 U751 ( .A1(n1047), .A2(n1044), .ZN(n1046) );
XOR2_X1 U752 ( .A(n1048), .B(n1049), .Z(n1047) );
NAND3_X1 U753 ( .A1(n1049), .A2(G900), .A3(G953), .ZN(n1045) );
NOR2_X1 U754 ( .A1(KEYINPUT0), .A2(n1050), .ZN(n1049) );
XOR2_X1 U755 ( .A(n1051), .B(n1052), .Z(n1050) );
XOR2_X1 U756 ( .A(n1053), .B(n1054), .Z(n1052) );
XNOR2_X1 U757 ( .A(G134), .B(KEYINPUT1), .ZN(n1054) );
NAND2_X1 U758 ( .A1(KEYINPUT48), .A2(n1055), .ZN(n1053) );
XOR2_X1 U759 ( .A(KEYINPUT58), .B(G137), .Z(n1055) );
XOR2_X1 U760 ( .A(n1056), .B(n1057), .Z(n1051) );
XNOR2_X1 U761 ( .A(n1058), .B(n1059), .ZN(n1057) );
XOR2_X1 U762 ( .A(n1060), .B(n1061), .Z(G69) );
XOR2_X1 U763 ( .A(n1062), .B(n1063), .Z(n1061) );
NOR2_X1 U764 ( .A1(n1064), .A2(G953), .ZN(n1063) );
NOR2_X1 U765 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
INV_X1 U766 ( .A(n1067), .ZN(n1065) );
NOR3_X1 U767 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1062) );
XNOR2_X1 U768 ( .A(n1071), .B(KEYINPUT6), .ZN(n1070) );
NOR2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1069) );
XOR2_X1 U770 ( .A(KEYINPUT52), .B(n1074), .Z(n1068) );
NOR2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
XNOR2_X1 U772 ( .A(KEYINPUT34), .B(n1072), .ZN(n1076) );
XNOR2_X1 U773 ( .A(n1073), .B(KEYINPUT25), .ZN(n1075) );
XOR2_X1 U774 ( .A(n1077), .B(n1078), .Z(n1073) );
NOR2_X1 U775 ( .A1(KEYINPUT11), .A2(n1079), .ZN(n1078) );
NOR2_X1 U776 ( .A1(n1080), .A2(n1044), .ZN(n1060) );
AND2_X1 U777 ( .A1(G224), .A2(G898), .ZN(n1080) );
NOR2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(G66) );
NOR3_X1 U779 ( .A1(n1038), .A2(n1083), .A3(n1084), .ZN(n1082) );
AND3_X1 U780 ( .A1(n1085), .A2(n1040), .A3(n1086), .ZN(n1084) );
INV_X1 U781 ( .A(n1087), .ZN(n1040) );
NOR2_X1 U782 ( .A1(n1088), .A2(n1085), .ZN(n1083) );
NOR2_X1 U783 ( .A1(n984), .A2(n1087), .ZN(n1088) );
NOR2_X1 U784 ( .A1(n1081), .A2(n1089), .ZN(G63) );
XOR2_X1 U785 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND3_X1 U786 ( .A1(n1086), .A2(G478), .A3(KEYINPUT32), .ZN(n1090) );
NOR2_X1 U787 ( .A1(n1081), .A2(n1092), .ZN(G60) );
XOR2_X1 U788 ( .A(n1093), .B(n1094), .Z(n1092) );
XNOR2_X1 U789 ( .A(KEYINPUT35), .B(n1095), .ZN(n1094) );
NAND2_X1 U790 ( .A1(n1086), .A2(G475), .ZN(n1093) );
XOR2_X1 U791 ( .A(n1096), .B(n1097), .Z(G6) );
NOR2_X1 U792 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U793 ( .A1(KEYINPUT47), .A2(n1100), .ZN(n1096) );
NOR2_X1 U794 ( .A1(n1081), .A2(n1101), .ZN(G57) );
XOR2_X1 U795 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U796 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U797 ( .A1(n1086), .A2(G472), .ZN(n1105) );
NAND2_X1 U798 ( .A1(n1106), .A2(KEYINPUT16), .ZN(n1104) );
XOR2_X1 U799 ( .A(n1107), .B(n1108), .Z(n1106) );
XNOR2_X1 U800 ( .A(G101), .B(n1109), .ZN(n1102) );
NOR2_X1 U801 ( .A1(n1081), .A2(n1110), .ZN(G54) );
XOR2_X1 U802 ( .A(n1111), .B(n1112), .Z(n1110) );
NAND2_X1 U803 ( .A1(n1086), .A2(G469), .ZN(n1112) );
NAND3_X1 U804 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1111) );
OR2_X1 U805 ( .A1(n1116), .A2(KEYINPUT23), .ZN(n1115) );
NAND3_X1 U806 ( .A1(KEYINPUT23), .A2(n1116), .A3(n1117), .ZN(n1114) );
NAND2_X1 U807 ( .A1(n1118), .A2(n1119), .ZN(n1113) );
NAND2_X1 U808 ( .A1(KEYINPUT23), .A2(n1120), .ZN(n1119) );
XNOR2_X1 U809 ( .A(KEYINPUT22), .B(n1116), .ZN(n1120) );
INV_X1 U810 ( .A(n1117), .ZN(n1118) );
XNOR2_X1 U811 ( .A(n1121), .B(n1122), .ZN(n1117) );
XNOR2_X1 U812 ( .A(G140), .B(n1123), .ZN(n1122) );
NOR2_X1 U813 ( .A1(n1044), .A2(G952), .ZN(n1081) );
NOR2_X1 U814 ( .A1(n1124), .A2(n1125), .ZN(G51) );
XOR2_X1 U815 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U816 ( .A1(n1086), .A2(n1128), .ZN(n1127) );
INV_X1 U817 ( .A(n1029), .ZN(n1128) );
NOR2_X1 U818 ( .A1(n1129), .A2(n984), .ZN(n1086) );
NOR3_X1 U819 ( .A1(n1048), .A2(n1066), .A3(n1130), .ZN(n984) );
XNOR2_X1 U820 ( .A(n1067), .B(KEYINPUT56), .ZN(n1130) );
NAND4_X1 U821 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1066) );
NOR3_X1 U822 ( .A1(n978), .A2(n1135), .A3(n1136), .ZN(n1134) );
INV_X1 U823 ( .A(n1137), .ZN(n1136) );
NOR2_X1 U824 ( .A1(n1138), .A2(n1098), .ZN(n978) );
NAND3_X1 U825 ( .A1(n1013), .A2(n1139), .A3(n1140), .ZN(n1098) );
NAND3_X1 U826 ( .A1(n1141), .A2(n1139), .A3(n1013), .ZN(n1133) );
NAND2_X1 U827 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U828 ( .A1(n1140), .A2(n1144), .ZN(n1143) );
XNOR2_X1 U829 ( .A(KEYINPUT63), .B(n1099), .ZN(n1144) );
NAND2_X1 U830 ( .A1(n1015), .A2(n1145), .ZN(n1142) );
NAND4_X1 U831 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1048) );
NOR4_X1 U832 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1149) );
INV_X1 U833 ( .A(n1154), .ZN(n1151) );
NAND3_X1 U834 ( .A1(n1155), .A2(n1156), .A3(n1000), .ZN(n1148) );
NAND2_X1 U835 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND3_X1 U836 ( .A1(n1145), .A2(n1159), .A3(n1140), .ZN(n1158) );
INV_X1 U837 ( .A(KEYINPUT36), .ZN(n1159) );
NAND3_X1 U838 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1155) );
NAND3_X1 U839 ( .A1(n1140), .A2(n1145), .A3(KEYINPUT36), .ZN(n1161) );
NAND2_X1 U840 ( .A1(n1014), .A2(n1163), .ZN(n1160) );
XNOR2_X1 U841 ( .A(KEYINPUT44), .B(n1099), .ZN(n1163) );
NAND4_X1 U842 ( .A1(n1006), .A2(n1014), .A3(n1162), .A4(n1164), .ZN(n1146) );
NAND2_X1 U843 ( .A1(n1165), .A2(n1166), .ZN(n1126) );
OR2_X1 U844 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U845 ( .A(n1169), .B(KEYINPUT3), .Z(n1165) );
NAND2_X1 U846 ( .A1(n1168), .A2(n1167), .ZN(n1169) );
XOR2_X1 U847 ( .A(n1170), .B(KEYINPUT33), .Z(n1167) );
NOR2_X1 U848 ( .A1(G952), .A2(n1171), .ZN(n1124) );
XNOR2_X1 U849 ( .A(G953), .B(KEYINPUT54), .ZN(n1171) );
XNOR2_X1 U850 ( .A(G146), .B(n1147), .ZN(G48) );
NAND2_X1 U851 ( .A1(n1172), .A2(n1173), .ZN(n1147) );
XNOR2_X1 U852 ( .A(G143), .B(n1174), .ZN(G45) );
NAND4_X1 U853 ( .A1(n1000), .A2(n1140), .A3(n1145), .A4(n1162), .ZN(n1174) );
XOR2_X1 U854 ( .A(G140), .B(n1153), .Z(G42) );
AND2_X1 U855 ( .A1(n1014), .A2(n1175), .ZN(n1153) );
XNOR2_X1 U856 ( .A(G137), .B(n1176), .ZN(G39) );
NAND4_X1 U857 ( .A1(n1177), .A2(n1006), .A3(n1014), .A4(n1164), .ZN(n1176) );
XNOR2_X1 U858 ( .A(n1157), .B(KEYINPUT57), .ZN(n1177) );
XOR2_X1 U859 ( .A(G134), .B(n1152), .Z(G36) );
NOR3_X1 U860 ( .A1(n1138), .A2(n1157), .A3(n1178), .ZN(n1152) );
XOR2_X1 U861 ( .A(G131), .B(n1179), .Z(G33) );
NOR2_X1 U862 ( .A1(n1180), .A2(n1178), .ZN(n1179) );
NAND2_X1 U863 ( .A1(n1000), .A2(n1014), .ZN(n1178) );
NOR3_X1 U864 ( .A1(n1181), .A2(n991), .A3(n993), .ZN(n1014) );
XNOR2_X1 U865 ( .A(G128), .B(n1154), .ZN(G30) );
NAND3_X1 U866 ( .A1(n1003), .A2(n1162), .A3(n1172), .ZN(n1154) );
AND3_X1 U867 ( .A1(n1140), .A2(n1164), .A3(n1182), .ZN(n1172) );
XNOR2_X1 U868 ( .A(G101), .B(n1137), .ZN(G3) );
NAND4_X1 U869 ( .A1(n1183), .A2(n1000), .A3(n1140), .A4(n1139), .ZN(n1137) );
XNOR2_X1 U870 ( .A(n1184), .B(n1150), .ZN(G27) );
AND2_X1 U871 ( .A1(n1015), .A2(n1175), .ZN(n1150) );
NOR3_X1 U872 ( .A1(n1185), .A2(n1164), .A3(n1180), .ZN(n1175) );
INV_X1 U873 ( .A(n1173), .ZN(n1180) );
NOR2_X1 U874 ( .A1(n1099), .A2(n1157), .ZN(n1173) );
INV_X1 U875 ( .A(n1162), .ZN(n1157) );
NAND2_X1 U876 ( .A1(n986), .A2(n1186), .ZN(n1162) );
NAND4_X1 U877 ( .A1(G902), .A2(G953), .A3(n1187), .A4(n1188), .ZN(n1186) );
INV_X1 U878 ( .A(G900), .ZN(n1188) );
XOR2_X1 U879 ( .A(n1189), .B(n1190), .Z(G24) );
XOR2_X1 U880 ( .A(KEYINPUT41), .B(G122), .Z(n1190) );
NAND4_X1 U881 ( .A1(n1191), .A2(n1145), .A3(n1013), .A4(n1192), .ZN(n1189) );
AND3_X1 U882 ( .A1(n1181), .A2(n1011), .A3(n1139), .ZN(n1192) );
NOR2_X1 U883 ( .A1(n1164), .A2(n1182), .ZN(n1013) );
NAND2_X1 U884 ( .A1(n1193), .A2(n1194), .ZN(n1145) );
OR2_X1 U885 ( .A1(n1138), .A2(KEYINPUT17), .ZN(n1194) );
INV_X1 U886 ( .A(n1003), .ZN(n1138) );
NAND3_X1 U887 ( .A1(n1195), .A2(n1196), .A3(KEYINPUT17), .ZN(n1193) );
XOR2_X1 U888 ( .A(KEYINPUT28), .B(n1197), .Z(n1191) );
AND2_X1 U889 ( .A1(n1010), .A2(n991), .ZN(n1197) );
INV_X1 U890 ( .A(n1198), .ZN(n991) );
XNOR2_X1 U891 ( .A(G119), .B(n1131), .ZN(G21) );
NAND4_X1 U892 ( .A1(n1006), .A2(n1015), .A3(n1164), .A4(n1139), .ZN(n1131) );
XOR2_X1 U893 ( .A(G116), .B(n1199), .Z(G18) );
NOR2_X1 U894 ( .A1(KEYINPUT15), .A2(n1067), .ZN(n1199) );
NAND2_X1 U895 ( .A1(n1200), .A2(n1003), .ZN(n1067) );
NOR2_X1 U896 ( .A1(n1195), .A2(n1201), .ZN(n1003) );
XNOR2_X1 U897 ( .A(G113), .B(n1132), .ZN(G15) );
NAND2_X1 U898 ( .A1(n1200), .A2(n1004), .ZN(n1132) );
INV_X1 U899 ( .A(n1099), .ZN(n1004) );
NAND2_X1 U900 ( .A1(n1201), .A2(n1202), .ZN(n1099) );
XNOR2_X1 U901 ( .A(KEYINPUT17), .B(n1195), .ZN(n1202) );
AND3_X1 U902 ( .A1(n1015), .A2(n1139), .A3(n1000), .ZN(n1200) );
NOR2_X1 U903 ( .A1(n1182), .A2(n1005), .ZN(n1000) );
INV_X1 U904 ( .A(n1185), .ZN(n1182) );
NOR3_X1 U905 ( .A1(n1198), .A2(n992), .A3(n993), .ZN(n1015) );
INV_X1 U906 ( .A(n1181), .ZN(n992) );
XOR2_X1 U907 ( .A(n1203), .B(n1204), .Z(G12) );
XNOR2_X1 U908 ( .A(KEYINPUT9), .B(n1123), .ZN(n1204) );
NAND2_X1 U909 ( .A1(KEYINPUT7), .A2(n1135), .ZN(n1203) );
AND4_X1 U910 ( .A1(n1006), .A2(n1140), .A3(n1005), .A4(n1139), .ZN(n1135) );
NAND2_X1 U911 ( .A1(n986), .A2(n1205), .ZN(n1139) );
NAND3_X1 U912 ( .A1(n1071), .A2(n1187), .A3(G902), .ZN(n1205) );
AND2_X1 U913 ( .A1(G953), .A2(n1206), .ZN(n1071) );
XOR2_X1 U914 ( .A(KEYINPUT4), .B(G898), .Z(n1206) );
NAND3_X1 U915 ( .A1(n1187), .A2(n1044), .A3(G952), .ZN(n986) );
NAND2_X1 U916 ( .A1(G237), .A2(G234), .ZN(n1187) );
INV_X1 U917 ( .A(n1164), .ZN(n1005) );
NAND2_X1 U918 ( .A1(n1207), .A2(n1035), .ZN(n1164) );
NAND2_X1 U919 ( .A1(G472), .A2(n1208), .ZN(n1035) );
OR2_X1 U920 ( .A1(n1209), .A2(G902), .ZN(n1208) );
XOR2_X1 U921 ( .A(KEYINPUT14), .B(n1033), .Z(n1207) );
NOR3_X1 U922 ( .A1(G472), .A2(G902), .A3(n1209), .ZN(n1033) );
XOR2_X1 U923 ( .A(n1210), .B(n1107), .Z(n1209) );
XOR2_X1 U924 ( .A(n1211), .B(n1212), .Z(n1107) );
INV_X1 U925 ( .A(n1213), .ZN(n1212) );
XOR2_X1 U926 ( .A(n1214), .B(n1215), .Z(n1210) );
NOR2_X1 U927 ( .A1(KEYINPUT60), .A2(n1108), .ZN(n1215) );
XNOR2_X1 U928 ( .A(n1216), .B(KEYINPUT45), .ZN(n1108) );
NAND3_X1 U929 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1214) );
OR2_X1 U930 ( .A1(n1109), .A2(KEYINPUT42), .ZN(n1219) );
NAND3_X1 U931 ( .A1(KEYINPUT42), .A2(n1109), .A3(n1220), .ZN(n1218) );
INV_X1 U932 ( .A(G101), .ZN(n1220) );
NAND2_X1 U933 ( .A1(G101), .A2(n1221), .ZN(n1217) );
NAND2_X1 U934 ( .A1(KEYINPUT42), .A2(n1222), .ZN(n1221) );
XNOR2_X1 U935 ( .A(KEYINPUT24), .B(n1109), .ZN(n1222) );
NAND2_X1 U936 ( .A1(G210), .A2(n1223), .ZN(n1109) );
NOR3_X1 U937 ( .A1(n1198), .A2(n1181), .A3(n993), .ZN(n1140) );
NAND2_X1 U938 ( .A1(n1011), .A2(n1010), .ZN(n993) );
NAND2_X1 U939 ( .A1(G214), .A2(n1224), .ZN(n1010) );
NAND2_X1 U940 ( .A1(G221), .A2(n1225), .ZN(n1011) );
XNOR2_X1 U941 ( .A(n1024), .B(n1226), .ZN(n1181) );
NOR2_X1 U942 ( .A1(G469), .A2(KEYINPUT26), .ZN(n1226) );
NAND3_X1 U943 ( .A1(n1227), .A2(n1228), .A3(n1129), .ZN(n1024) );
NAND3_X1 U944 ( .A1(n1229), .A2(n1116), .A3(n1230), .ZN(n1228) );
INV_X1 U945 ( .A(KEYINPUT20), .ZN(n1230) );
NAND2_X1 U946 ( .A1(n1231), .A2(KEYINPUT20), .ZN(n1227) );
XOR2_X1 U947 ( .A(n1116), .B(n1229), .Z(n1231) );
XOR2_X1 U948 ( .A(n1232), .B(n1233), .Z(n1229) );
NOR2_X1 U949 ( .A1(KEYINPUT62), .A2(n1121), .ZN(n1233) );
NAND2_X1 U950 ( .A1(G227), .A2(n1044), .ZN(n1121) );
XNOR2_X1 U951 ( .A(G110), .B(n1234), .ZN(n1232) );
NOR2_X1 U952 ( .A1(G140), .A2(KEYINPUT46), .ZN(n1234) );
XOR2_X1 U953 ( .A(n1235), .B(n1236), .Z(n1116) );
XNOR2_X1 U954 ( .A(n1213), .B(n1237), .ZN(n1236) );
XNOR2_X1 U955 ( .A(G101), .B(KEYINPUT8), .ZN(n1237) );
XNOR2_X1 U956 ( .A(n1238), .B(n1239), .ZN(n1213) );
XOR2_X1 U957 ( .A(G137), .B(G134), .Z(n1239) );
NAND2_X1 U958 ( .A1(KEYINPUT29), .A2(n1240), .ZN(n1238) );
XOR2_X1 U959 ( .A(n1056), .B(n1241), .Z(n1235) );
XNOR2_X1 U960 ( .A(G128), .B(n1242), .ZN(n1056) );
XOR2_X1 U961 ( .A(n1243), .B(n1031), .Z(n1198) );
NAND2_X1 U962 ( .A1(n1244), .A2(n1129), .ZN(n1031) );
XNOR2_X1 U963 ( .A(n1168), .B(n1170), .ZN(n1244) );
XNOR2_X1 U964 ( .A(n1245), .B(n1216), .ZN(n1170) );
XOR2_X1 U965 ( .A(n1242), .B(n1246), .Z(n1216) );
NOR2_X1 U966 ( .A1(KEYINPUT50), .A2(n1247), .ZN(n1246) );
XNOR2_X1 U967 ( .A(G146), .B(n1248), .ZN(n1242) );
XNOR2_X1 U968 ( .A(G125), .B(n1249), .ZN(n1245) );
AND2_X1 U969 ( .A1(n1044), .A2(G224), .ZN(n1249) );
AND2_X1 U970 ( .A1(n1250), .A2(n1251), .ZN(n1168) );
NAND2_X1 U971 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
XNOR2_X1 U972 ( .A(n1254), .B(n1079), .ZN(n1252) );
NAND2_X1 U973 ( .A1(n1255), .A2(n1256), .ZN(n1250) );
XNOR2_X1 U974 ( .A(KEYINPUT40), .B(n1072), .ZN(n1256) );
INV_X1 U975 ( .A(n1253), .ZN(n1072) );
XOR2_X1 U976 ( .A(G110), .B(n1257), .Z(n1253) );
XOR2_X1 U977 ( .A(KEYINPUT18), .B(G122), .Z(n1257) );
XOR2_X1 U978 ( .A(n1254), .B(n1079), .Z(n1255) );
XOR2_X1 U979 ( .A(n1211), .B(KEYINPUT19), .Z(n1079) );
XNOR2_X1 U980 ( .A(G113), .B(n1258), .ZN(n1211) );
XOR2_X1 U981 ( .A(G119), .B(G116), .Z(n1258) );
NAND2_X1 U982 ( .A1(KEYINPUT39), .A2(n1077), .ZN(n1254) );
XOR2_X1 U983 ( .A(G101), .B(n1259), .Z(n1077) );
NOR2_X1 U984 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NOR3_X1 U985 ( .A1(KEYINPUT55), .A2(G107), .A3(n1100), .ZN(n1261) );
NOR2_X1 U986 ( .A1(n1241), .A2(n1262), .ZN(n1260) );
INV_X1 U987 ( .A(KEYINPUT55), .ZN(n1262) );
XNOR2_X1 U988 ( .A(n1100), .B(G107), .ZN(n1241) );
INV_X1 U989 ( .A(G104), .ZN(n1100) );
NAND2_X1 U990 ( .A1(KEYINPUT53), .A2(n1029), .ZN(n1243) );
NAND2_X1 U991 ( .A1(G210), .A2(n1224), .ZN(n1029) );
NAND2_X1 U992 ( .A1(n1263), .A2(n1129), .ZN(n1224) );
INV_X1 U993 ( .A(G237), .ZN(n1263) );
NOR2_X1 U994 ( .A1(n999), .A2(n1185), .ZN(n1006) );
XOR2_X1 U995 ( .A(n1264), .B(n1087), .Z(n1185) );
NAND2_X1 U996 ( .A1(G217), .A2(n1225), .ZN(n1087) );
NAND2_X1 U997 ( .A1(G234), .A2(n1129), .ZN(n1225) );
XNOR2_X1 U998 ( .A(n1038), .B(KEYINPUT49), .ZN(n1264) );
NOR2_X1 U999 ( .A1(n1085), .A2(G902), .ZN(n1038) );
XOR2_X1 U1000 ( .A(n1265), .B(n1266), .Z(n1085) );
XOR2_X1 U1001 ( .A(G119), .B(n1267), .Z(n1266) );
XNOR2_X1 U1002 ( .A(G137), .B(n1247), .ZN(n1267) );
XOR2_X1 U1003 ( .A(n1268), .B(n1269), .Z(n1265) );
XNOR2_X1 U1004 ( .A(n1270), .B(n1123), .ZN(n1268) );
INV_X1 U1005 ( .A(G110), .ZN(n1123) );
NAND2_X1 U1006 ( .A1(G221), .A2(n1271), .ZN(n1270) );
INV_X1 U1007 ( .A(n1183), .ZN(n999) );
NOR2_X1 U1008 ( .A1(n1196), .A2(n1195), .ZN(n1183) );
NAND2_X1 U1009 ( .A1(n1272), .A2(n1273), .ZN(n1195) );
NAND2_X1 U1010 ( .A1(n1274), .A2(G475), .ZN(n1273) );
XOR2_X1 U1011 ( .A(KEYINPUT12), .B(n1275), .Z(n1272) );
NOR2_X1 U1012 ( .A1(G475), .A2(n1274), .ZN(n1275) );
XOR2_X1 U1013 ( .A(n1023), .B(KEYINPUT10), .Z(n1274) );
NAND2_X1 U1014 ( .A1(n1129), .A2(n1095), .ZN(n1023) );
NAND2_X1 U1015 ( .A1(n1276), .A2(n1277), .ZN(n1095) );
OR2_X1 U1016 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
XOR2_X1 U1017 ( .A(n1280), .B(KEYINPUT27), .Z(n1276) );
NAND2_X1 U1018 ( .A1(n1279), .A2(n1278), .ZN(n1280) );
XOR2_X1 U1019 ( .A(G104), .B(n1281), .Z(n1278) );
XOR2_X1 U1020 ( .A(G122), .B(G113), .Z(n1281) );
XNOR2_X1 U1021 ( .A(n1282), .B(n1269), .ZN(n1279) );
XOR2_X1 U1022 ( .A(G146), .B(n1058), .Z(n1269) );
XNOR2_X1 U1023 ( .A(n1184), .B(G140), .ZN(n1058) );
INV_X1 U1024 ( .A(G125), .ZN(n1184) );
NAND2_X1 U1025 ( .A1(KEYINPUT51), .A2(n1283), .ZN(n1282) );
XOR2_X1 U1026 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U1027 ( .A(G143), .B(n1286), .ZN(n1285) );
NAND2_X1 U1028 ( .A1(G214), .A2(n1223), .ZN(n1286) );
NOR2_X1 U1029 ( .A1(G953), .A2(G237), .ZN(n1223) );
NOR2_X1 U1030 ( .A1(KEYINPUT21), .A2(n1059), .ZN(n1284) );
INV_X1 U1031 ( .A(n1240), .ZN(n1059) );
XOR2_X1 U1032 ( .A(G131), .B(KEYINPUT43), .Z(n1240) );
INV_X1 U1033 ( .A(n1201), .ZN(n1196) );
NOR2_X1 U1034 ( .A1(n1287), .A2(n1034), .ZN(n1201) );
NOR2_X1 U1035 ( .A1(n1037), .A2(G478), .ZN(n1034) );
AND2_X1 U1036 ( .A1(G478), .A2(n1037), .ZN(n1287) );
NAND2_X1 U1037 ( .A1(n1091), .A2(n1129), .ZN(n1037) );
INV_X1 U1038 ( .A(G902), .ZN(n1129) );
XNOR2_X1 U1039 ( .A(n1288), .B(n1289), .ZN(n1091) );
AND2_X1 U1040 ( .A1(n1271), .A2(G217), .ZN(n1289) );
AND2_X1 U1041 ( .A1(G234), .A2(n1044), .ZN(n1271) );
INV_X1 U1042 ( .A(G953), .ZN(n1044) );
NAND2_X1 U1043 ( .A1(n1290), .A2(KEYINPUT37), .ZN(n1288) );
XOR2_X1 U1044 ( .A(n1291), .B(n1292), .Z(n1290) );
XNOR2_X1 U1045 ( .A(n1247), .B(n1293), .ZN(n1292) );
XNOR2_X1 U1046 ( .A(n1248), .B(G134), .ZN(n1293) );
INV_X1 U1047 ( .A(G143), .ZN(n1248) );
INV_X1 U1048 ( .A(G128), .ZN(n1247) );
XOR2_X1 U1049 ( .A(n1294), .B(n1295), .Z(n1291) );
NOR2_X1 U1050 ( .A1(KEYINPUT59), .A2(G107), .ZN(n1295) );
XNOR2_X1 U1051 ( .A(G116), .B(G122), .ZN(n1294) );
endmodule


