//Key = 1011001001010111000011111000001011100001110110101011000101001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;

XNOR2_X1 U755 ( .A(G107), .B(n1046), .ZN(G9) );
NAND4_X1 U756 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
NOR2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
XOR2_X1 U758 ( .A(n1053), .B(KEYINPUT39), .Z(n1052) );
INV_X1 U759 ( .A(n1054), .ZN(n1051) );
NAND3_X1 U760 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(G75) );
NAND2_X1 U761 ( .A1(G952), .A2(n1058), .ZN(n1057) );
NAND3_X1 U762 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
NAND2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NAND2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND3_X1 U765 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
NAND2_X1 U766 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NAND2_X1 U767 ( .A1(n1048), .A2(n1071), .ZN(n1070) );
NAND2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1069) );
NAND2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U771 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND3_X1 U772 ( .A1(n1074), .A2(n1080), .A3(n1048), .ZN(n1064) );
NAND2_X1 U773 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U774 ( .A1(n1066), .A2(n1083), .ZN(n1082) );
NAND2_X1 U775 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U776 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U777 ( .A(KEYINPUT27), .B(n1088), .Z(n1087) );
INV_X1 U778 ( .A(n1047), .ZN(n1084) );
NAND2_X1 U779 ( .A1(n1068), .A2(n1089), .ZN(n1081) );
NAND2_X1 U780 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U781 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U782 ( .A(n1094), .B(KEYINPUT37), .Z(n1062) );
NAND4_X1 U783 ( .A1(n1066), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1055) );
NOR3_X1 U784 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1097) );
XOR2_X1 U785 ( .A(n1101), .B(n1102), .Z(n1100) );
XNOR2_X1 U786 ( .A(G475), .B(n1103), .ZN(n1099) );
NAND4_X1 U787 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1098) );
NAND2_X1 U788 ( .A1(KEYINPUT31), .A2(n1108), .ZN(n1107) );
NAND2_X1 U789 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XNOR2_X1 U790 ( .A(KEYINPUT41), .B(n1111), .ZN(n1109) );
NAND2_X1 U791 ( .A1(n1112), .A2(n1113), .ZN(n1106) );
INV_X1 U792 ( .A(KEYINPUT31), .ZN(n1113) );
NAND2_X1 U793 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NAND3_X1 U794 ( .A1(KEYINPUT41), .A2(n1110), .A3(n1111), .ZN(n1115) );
OR2_X1 U795 ( .A1(n1111), .A2(KEYINPUT41), .ZN(n1114) );
NAND2_X1 U796 ( .A1(KEYINPUT4), .A2(n1116), .ZN(n1105) );
OR2_X1 U797 ( .A1(n1117), .A2(KEYINPUT4), .ZN(n1104) );
NOR3_X1 U798 ( .A1(n1118), .A2(n1119), .A3(n1086), .ZN(n1096) );
INV_X1 U799 ( .A(n1120), .ZN(n1119) );
NOR2_X1 U800 ( .A1(n1111), .A2(n1110), .ZN(n1118) );
XNOR2_X1 U801 ( .A(G472), .B(n1121), .ZN(n1095) );
NAND2_X1 U802 ( .A1(KEYINPUT62), .A2(n1122), .ZN(n1121) );
NAND2_X1 U803 ( .A1(n1123), .A2(n1124), .ZN(G72) );
NAND2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
NAND3_X1 U806 ( .A1(n1129), .A2(n1056), .A3(KEYINPUT46), .ZN(n1128) );
NAND2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1127) );
NAND4_X1 U808 ( .A1(n1132), .A2(n1133), .A3(n1059), .A4(n1134), .ZN(n1123) );
INV_X1 U809 ( .A(n1126), .ZN(n1134) );
NAND2_X1 U810 ( .A1(n1135), .A2(n1136), .ZN(n1126) );
NAND2_X1 U811 ( .A1(G953), .A2(n1137), .ZN(n1136) );
XOR2_X1 U812 ( .A(n1138), .B(n1139), .Z(n1135) );
XNOR2_X1 U813 ( .A(G125), .B(G140), .ZN(n1139) );
NAND2_X1 U814 ( .A1(n1140), .A2(n1141), .ZN(n1138) );
NAND4_X1 U815 ( .A1(G137), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1141) );
NAND2_X1 U816 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U817 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
NAND3_X1 U818 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1140) );
NAND2_X1 U819 ( .A1(G137), .A2(n1142), .ZN(n1151) );
INV_X1 U820 ( .A(KEYINPUT45), .ZN(n1142) );
NAND2_X1 U821 ( .A1(n1148), .A2(n1146), .ZN(n1150) );
INV_X1 U822 ( .A(n1147), .ZN(n1146) );
XNOR2_X1 U823 ( .A(KEYINPUT13), .B(n1152), .ZN(n1148) );
NAND2_X1 U824 ( .A1(n1145), .A2(n1147), .ZN(n1149) );
XNOR2_X1 U825 ( .A(KEYINPUT15), .B(n1153), .ZN(n1145) );
OR2_X1 U826 ( .A1(n1130), .A2(KEYINPUT46), .ZN(n1133) );
NAND3_X1 U827 ( .A1(n1130), .A2(n1131), .A3(KEYINPUT46), .ZN(n1132) );
INV_X1 U828 ( .A(KEYINPUT26), .ZN(n1131) );
AND2_X1 U829 ( .A1(G953), .A2(n1154), .ZN(n1130) );
NAND2_X1 U830 ( .A1(G900), .A2(G227), .ZN(n1154) );
XOR2_X1 U831 ( .A(n1155), .B(n1156), .Z(G69) );
XOR2_X1 U832 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U833 ( .A1(n1056), .A2(n1159), .ZN(n1158) );
NAND3_X1 U834 ( .A1(n1160), .A2(n1161), .A3(KEYINPUT51), .ZN(n1157) );
NAND2_X1 U835 ( .A1(G953), .A2(n1162), .ZN(n1161) );
XOR2_X1 U836 ( .A(n1163), .B(n1164), .Z(n1160) );
XOR2_X1 U837 ( .A(n1165), .B(KEYINPUT43), .Z(n1164) );
NOR2_X1 U838 ( .A1(n1166), .A2(n1056), .ZN(n1155) );
NOR2_X1 U839 ( .A1(n1167), .A2(n1162), .ZN(n1166) );
NOR2_X1 U840 ( .A1(n1168), .A2(n1169), .ZN(G66) );
NOR2_X1 U841 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U842 ( .A(KEYINPUT47), .B(n1172), .Z(n1171) );
NOR2_X1 U843 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U844 ( .A(KEYINPUT9), .B(n1175), .Z(n1174) );
NOR2_X1 U845 ( .A1(n1175), .A2(n1176), .ZN(n1170) );
INV_X1 U846 ( .A(n1173), .ZN(n1176) );
NOR2_X1 U847 ( .A1(n1177), .A2(n1102), .ZN(n1173) );
NOR2_X1 U848 ( .A1(n1168), .A2(n1178), .ZN(G63) );
XOR2_X1 U849 ( .A(n1179), .B(n1180), .Z(n1178) );
NAND2_X1 U850 ( .A1(n1181), .A2(G478), .ZN(n1179) );
NOR2_X1 U851 ( .A1(n1168), .A2(n1182), .ZN(G60) );
NOR3_X1 U852 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1182) );
NOR3_X1 U853 ( .A1(n1186), .A2(n1187), .A3(n1177), .ZN(n1185) );
NOR2_X1 U854 ( .A1(n1188), .A2(n1189), .ZN(n1184) );
NOR2_X1 U855 ( .A1(n1190), .A2(n1187), .ZN(n1188) );
NOR2_X1 U856 ( .A1(n1129), .A2(n1159), .ZN(n1190) );
XOR2_X1 U857 ( .A(G104), .B(n1191), .Z(G6) );
NOR2_X1 U858 ( .A1(n1168), .A2(n1192), .ZN(G57) );
XOR2_X1 U859 ( .A(n1193), .B(n1194), .Z(n1192) );
NAND2_X1 U860 ( .A1(KEYINPUT33), .A2(n1195), .ZN(n1194) );
NAND2_X1 U861 ( .A1(n1196), .A2(n1197), .ZN(n1193) );
NAND2_X1 U862 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U863 ( .A(n1200), .B(n1201), .Z(n1196) );
NOR2_X1 U864 ( .A1(n1198), .A2(n1199), .ZN(n1201) );
INV_X1 U865 ( .A(KEYINPUT40), .ZN(n1199) );
XNOR2_X1 U866 ( .A(n1202), .B(n1203), .ZN(n1198) );
NAND2_X1 U867 ( .A1(KEYINPUT14), .A2(n1204), .ZN(n1202) );
NAND2_X1 U868 ( .A1(n1181), .A2(G472), .ZN(n1200) );
NOR2_X1 U869 ( .A1(n1168), .A2(n1205), .ZN(G54) );
XOR2_X1 U870 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U871 ( .A(n1208), .B(n1209), .Z(n1207) );
NAND2_X1 U872 ( .A1(KEYINPUT61), .A2(n1153), .ZN(n1208) );
XNOR2_X1 U873 ( .A(KEYINPUT12), .B(n1210), .ZN(n1206) );
NOR3_X1 U874 ( .A1(n1177), .A2(KEYINPUT19), .A3(n1211), .ZN(n1210) );
NOR2_X1 U875 ( .A1(n1168), .A2(n1212), .ZN(G51) );
NOR2_X1 U876 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XOR2_X1 U877 ( .A(n1215), .B(n1216), .Z(n1214) );
NAND2_X1 U878 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NAND2_X1 U879 ( .A1(n1181), .A2(n1219), .ZN(n1215) );
INV_X1 U880 ( .A(n1177), .ZN(n1181) );
NAND2_X1 U881 ( .A1(G902), .A2(n1220), .ZN(n1177) );
NAND2_X1 U882 ( .A1(n1061), .A2(n1059), .ZN(n1220) );
INV_X1 U883 ( .A(n1129), .ZN(n1059) );
NAND4_X1 U884 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1129) );
AND4_X1 U885 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1224) );
NAND4_X1 U886 ( .A1(n1229), .A2(n1230), .A3(n1068), .A4(n1231), .ZN(n1228) );
NOR2_X1 U887 ( .A1(n1232), .A2(n1233), .ZN(n1223) );
INV_X1 U888 ( .A(n1159), .ZN(n1061) );
NAND4_X1 U889 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1159) );
NOR4_X1 U890 ( .A1(n1238), .A2(n1239), .A3(n1191), .A4(n1240), .ZN(n1237) );
INV_X1 U891 ( .A(n1241), .ZN(n1240) );
AND3_X1 U892 ( .A1(n1242), .A2(n1048), .A3(n1243), .ZN(n1191) );
NAND2_X1 U893 ( .A1(n1050), .A2(n1244), .ZN(n1236) );
NAND2_X1 U894 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND3_X1 U895 ( .A1(n1247), .A2(n1230), .A3(n1248), .ZN(n1246) );
NAND2_X1 U896 ( .A1(n1243), .A2(n1048), .ZN(n1245) );
NOR2_X1 U897 ( .A1(n1217), .A2(n1218), .ZN(n1213) );
INV_X1 U898 ( .A(KEYINPUT25), .ZN(n1218) );
XNOR2_X1 U899 ( .A(n1249), .B(n1250), .ZN(n1217) );
NAND2_X1 U900 ( .A1(KEYINPUT63), .A2(n1251), .ZN(n1249) );
NOR2_X1 U901 ( .A1(n1056), .A2(G952), .ZN(n1168) );
XNOR2_X1 U902 ( .A(G146), .B(n1227), .ZN(G48) );
NAND3_X1 U903 ( .A1(n1252), .A2(n1242), .A3(n1253), .ZN(n1227) );
XNOR2_X1 U904 ( .A(G143), .B(n1226), .ZN(G45) );
NAND3_X1 U905 ( .A1(n1254), .A2(n1247), .A3(n1253), .ZN(n1226) );
NAND2_X1 U906 ( .A1(n1255), .A2(n1256), .ZN(G42) );
NAND2_X1 U907 ( .A1(G140), .A2(n1225), .ZN(n1256) );
XOR2_X1 U908 ( .A(n1257), .B(KEYINPUT56), .Z(n1255) );
OR2_X1 U909 ( .A1(n1225), .A2(G140), .ZN(n1257) );
NAND2_X1 U910 ( .A1(n1231), .A2(n1258), .ZN(n1225) );
XNOR2_X1 U911 ( .A(G137), .B(n1221), .ZN(G39) );
NAND4_X1 U912 ( .A1(n1078), .A2(n1258), .A3(n1074), .A4(n1259), .ZN(n1221) );
XNOR2_X1 U913 ( .A(G134), .B(n1222), .ZN(G36) );
NAND3_X1 U914 ( .A1(n1247), .A2(n1050), .A3(n1258), .ZN(n1222) );
XOR2_X1 U915 ( .A(G131), .B(n1233), .Z(G33) );
AND3_X1 U916 ( .A1(n1247), .A2(n1242), .A3(n1258), .ZN(n1233) );
AND2_X1 U917 ( .A1(n1253), .A2(n1066), .ZN(n1258) );
NOR2_X1 U918 ( .A1(n1260), .A2(n1092), .ZN(n1066) );
XNOR2_X1 U919 ( .A(G128), .B(n1261), .ZN(G30) );
NOR2_X1 U920 ( .A1(n1232), .A2(KEYINPUT10), .ZN(n1261) );
AND3_X1 U921 ( .A1(n1252), .A2(n1050), .A3(n1253), .ZN(n1232) );
AND2_X1 U922 ( .A1(n1047), .A2(n1229), .ZN(n1253) );
XOR2_X1 U923 ( .A(n1239), .B(n1262), .Z(G3) );
XOR2_X1 U924 ( .A(KEYINPUT42), .B(G101), .Z(n1262) );
AND3_X1 U925 ( .A1(n1243), .A2(n1074), .A3(n1247), .ZN(n1239) );
XOR2_X1 U926 ( .A(n1263), .B(n1264), .Z(G27) );
NAND2_X1 U927 ( .A1(KEYINPUT22), .A2(G125), .ZN(n1264) );
NAND4_X1 U928 ( .A1(n1265), .A2(n1231), .A3(n1068), .A4(n1229), .ZN(n1263) );
NAND2_X1 U929 ( .A1(n1266), .A2(n1267), .ZN(n1229) );
NAND2_X1 U930 ( .A1(n1268), .A2(n1137), .ZN(n1267) );
INV_X1 U931 ( .A(G900), .ZN(n1137) );
NOR3_X1 U932 ( .A1(n1259), .A2(n1072), .A3(n1269), .ZN(n1231) );
INV_X1 U933 ( .A(n1242), .ZN(n1072) );
XNOR2_X1 U934 ( .A(n1230), .B(KEYINPUT11), .ZN(n1265) );
XNOR2_X1 U935 ( .A(G122), .B(n1234), .ZN(G24) );
NAND3_X1 U936 ( .A1(n1248), .A2(n1048), .A3(n1254), .ZN(n1234) );
AND3_X1 U937 ( .A1(n1270), .A2(n1271), .A3(n1230), .ZN(n1254) );
NOR2_X1 U938 ( .A1(n1259), .A2(n1078), .ZN(n1048) );
XNOR2_X1 U939 ( .A(G119), .B(n1235), .ZN(G21) );
NAND3_X1 U940 ( .A1(n1248), .A2(n1074), .A3(n1252), .ZN(n1235) );
NOR3_X1 U941 ( .A1(n1090), .A2(n1079), .A3(n1269), .ZN(n1252) );
XOR2_X1 U942 ( .A(n1272), .B(n1273), .Z(G18) );
NOR4_X1 U943 ( .A1(n1274), .A2(n1090), .A3(n1076), .A4(n1275), .ZN(n1273) );
INV_X1 U944 ( .A(n1247), .ZN(n1076) );
INV_X1 U945 ( .A(n1230), .ZN(n1090) );
XNOR2_X1 U946 ( .A(n1050), .B(KEYINPUT36), .ZN(n1274) );
INV_X1 U947 ( .A(n1073), .ZN(n1050) );
NAND2_X1 U948 ( .A1(n1270), .A2(n1276), .ZN(n1073) );
XNOR2_X1 U949 ( .A(KEYINPUT53), .B(n1271), .ZN(n1276) );
XOR2_X1 U950 ( .A(n1277), .B(KEYINPUT5), .Z(n1270) );
NAND2_X1 U951 ( .A1(KEYINPUT44), .A2(n1278), .ZN(n1272) );
XNOR2_X1 U952 ( .A(G113), .B(n1241), .ZN(G15) );
NAND4_X1 U953 ( .A1(n1248), .A2(n1247), .A3(n1053), .A4(n1242), .ZN(n1241) );
NOR2_X1 U954 ( .A1(n1079), .A2(n1078), .ZN(n1247) );
INV_X1 U955 ( .A(n1275), .ZN(n1248) );
NAND2_X1 U956 ( .A1(n1068), .A2(n1054), .ZN(n1275) );
AND2_X1 U957 ( .A1(n1279), .A2(n1280), .ZN(n1068) );
XNOR2_X1 U958 ( .A(n1088), .B(KEYINPUT32), .ZN(n1279) );
XNOR2_X1 U959 ( .A(n1238), .B(n1281), .ZN(G12) );
NAND2_X1 U960 ( .A1(KEYINPUT57), .A2(G110), .ZN(n1281) );
AND4_X1 U961 ( .A1(n1078), .A2(n1243), .A3(n1079), .A4(n1074), .ZN(n1238) );
NAND2_X1 U962 ( .A1(n1282), .A2(n1283), .ZN(n1074) );
OR3_X1 U963 ( .A1(n1277), .A2(n1271), .A3(KEYINPUT53), .ZN(n1283) );
INV_X1 U964 ( .A(n1284), .ZN(n1271) );
NAND2_X1 U965 ( .A1(KEYINPUT53), .A2(n1242), .ZN(n1282) );
NOR2_X1 U966 ( .A1(n1284), .A2(n1277), .ZN(n1242) );
NAND2_X1 U967 ( .A1(n1285), .A2(n1120), .ZN(n1277) );
NAND3_X1 U968 ( .A1(n1116), .A2(n1286), .A3(n1180), .ZN(n1120) );
INV_X1 U969 ( .A(G478), .ZN(n1116) );
XOR2_X1 U970 ( .A(n1117), .B(KEYINPUT8), .Z(n1285) );
NAND2_X1 U971 ( .A1(G478), .A2(n1287), .ZN(n1117) );
NAND2_X1 U972 ( .A1(n1180), .A2(n1286), .ZN(n1287) );
XOR2_X1 U973 ( .A(n1288), .B(n1289), .Z(n1180) );
XOR2_X1 U974 ( .A(n1290), .B(n1291), .Z(n1289) );
XNOR2_X1 U975 ( .A(n1278), .B(n1292), .ZN(n1291) );
AND4_X1 U976 ( .A1(n1293), .A2(n1056), .A3(G234), .A4(G217), .ZN(n1292) );
INV_X1 U977 ( .A(KEYINPUT17), .ZN(n1293) );
INV_X1 U978 ( .A(G116), .ZN(n1278) );
XNOR2_X1 U979 ( .A(G134), .B(n1294), .ZN(n1290) );
XNOR2_X1 U980 ( .A(n1295), .B(n1296), .ZN(n1288) );
XNOR2_X1 U981 ( .A(n1297), .B(n1298), .ZN(n1296) );
NOR2_X1 U982 ( .A1(G143), .A2(KEYINPUT49), .ZN(n1298) );
NAND2_X1 U983 ( .A1(KEYINPUT30), .A2(n1299), .ZN(n1297) );
XOR2_X1 U984 ( .A(n1300), .B(n1103), .Z(n1284) );
INV_X1 U985 ( .A(n1183), .ZN(n1103) );
NOR2_X1 U986 ( .A1(n1189), .A2(G902), .ZN(n1183) );
INV_X1 U987 ( .A(n1186), .ZN(n1189) );
XNOR2_X1 U988 ( .A(n1301), .B(G104), .ZN(n1186) );
XOR2_X1 U989 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U990 ( .A(n1304), .B(n1305), .Z(n1303) );
XOR2_X1 U991 ( .A(G140), .B(G131), .Z(n1305) );
XOR2_X1 U992 ( .A(KEYINPUT0), .B(G146), .Z(n1304) );
XOR2_X1 U993 ( .A(n1306), .B(n1307), .Z(n1302) );
XOR2_X1 U994 ( .A(n1295), .B(n1308), .Z(n1307) );
XOR2_X1 U995 ( .A(n1309), .B(n1310), .Z(n1306) );
NOR2_X1 U996 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U997 ( .A(KEYINPUT58), .B(n1313), .Z(n1312) );
NOR2_X1 U998 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
XOR2_X1 U999 ( .A(n1316), .B(KEYINPUT1), .Z(n1314) );
AND2_X1 U1000 ( .A1(n1316), .A2(n1315), .ZN(n1311) );
NAND2_X1 U1001 ( .A1(G214), .A2(n1317), .ZN(n1316) );
NAND2_X1 U1002 ( .A1(KEYINPUT20), .A2(n1318), .ZN(n1309) );
NAND2_X1 U1003 ( .A1(KEYINPUT24), .A2(n1187), .ZN(n1300) );
INV_X1 U1004 ( .A(G475), .ZN(n1187) );
INV_X1 U1005 ( .A(n1259), .ZN(n1079) );
XNOR2_X1 U1006 ( .A(n1122), .B(G472), .ZN(n1259) );
NAND2_X1 U1007 ( .A1(n1319), .A2(n1286), .ZN(n1122) );
XOR2_X1 U1008 ( .A(n1195), .B(n1320), .Z(n1319) );
NOR2_X1 U1009 ( .A1(KEYINPUT29), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1010 ( .A(n1204), .B(n1203), .Z(n1321) );
XNOR2_X1 U1011 ( .A(n1322), .B(n1323), .ZN(n1203) );
XOR2_X1 U1012 ( .A(KEYINPUT54), .B(KEYINPUT16), .Z(n1323) );
XNOR2_X1 U1013 ( .A(n1324), .B(n1318), .ZN(n1322) );
INV_X1 U1014 ( .A(G113), .ZN(n1318) );
XNOR2_X1 U1015 ( .A(n1325), .B(n1326), .ZN(n1204) );
INV_X1 U1016 ( .A(n1327), .ZN(n1326) );
XOR2_X1 U1017 ( .A(n1328), .B(G101), .Z(n1195) );
NAND2_X1 U1018 ( .A1(G210), .A2(n1317), .ZN(n1328) );
NOR2_X1 U1019 ( .A1(G953), .A2(G237), .ZN(n1317) );
AND3_X1 U1020 ( .A1(n1053), .A2(n1054), .A3(n1047), .ZN(n1243) );
NOR2_X1 U1021 ( .A1(n1088), .A2(n1086), .ZN(n1047) );
INV_X1 U1022 ( .A(n1280), .ZN(n1086) );
NAND2_X1 U1023 ( .A1(G221), .A2(n1329), .ZN(n1280) );
XOR2_X1 U1024 ( .A(n1110), .B(n1111), .Z(n1088) );
XOR2_X1 U1025 ( .A(n1211), .B(KEYINPUT50), .Z(n1111) );
INV_X1 U1026 ( .A(G469), .ZN(n1211) );
NAND2_X1 U1027 ( .A1(n1330), .A2(n1286), .ZN(n1110) );
XNOR2_X1 U1028 ( .A(n1209), .B(n1153), .ZN(n1330) );
INV_X1 U1029 ( .A(n1152), .ZN(n1153) );
XOR2_X1 U1030 ( .A(G128), .B(n1331), .Z(n1152) );
NOR2_X1 U1031 ( .A1(KEYINPUT38), .A2(n1332), .ZN(n1331) );
XNOR2_X1 U1032 ( .A(G146), .B(n1315), .ZN(n1332) );
INV_X1 U1033 ( .A(G143), .ZN(n1315) );
XOR2_X1 U1034 ( .A(n1333), .B(n1334), .Z(n1209) );
XOR2_X1 U1035 ( .A(n1335), .B(n1336), .Z(n1334) );
XNOR2_X1 U1036 ( .A(G101), .B(n1337), .ZN(n1336) );
NOR2_X1 U1037 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
XNOR2_X1 U1038 ( .A(KEYINPUT7), .B(n1056), .ZN(n1339) );
INV_X1 U1039 ( .A(G227), .ZN(n1338) );
NAND2_X1 U1040 ( .A1(n1340), .A2(KEYINPUT34), .ZN(n1335) );
XNOR2_X1 U1041 ( .A(G107), .B(n1341), .ZN(n1340) );
XOR2_X1 U1042 ( .A(n1325), .B(n1342), .Z(n1333) );
XNOR2_X1 U1043 ( .A(n1147), .B(G137), .ZN(n1325) );
XOR2_X1 U1044 ( .A(G131), .B(n1343), .Z(n1147) );
XOR2_X1 U1045 ( .A(KEYINPUT18), .B(G134), .Z(n1343) );
NAND2_X1 U1046 ( .A1(n1266), .A2(n1344), .ZN(n1054) );
NAND2_X1 U1047 ( .A1(n1268), .A2(n1162), .ZN(n1344) );
INV_X1 U1048 ( .A(G898), .ZN(n1162) );
AND3_X1 U1049 ( .A1(G953), .A2(n1094), .A3(G902), .ZN(n1268) );
NAND3_X1 U1050 ( .A1(n1094), .A2(n1056), .A3(G952), .ZN(n1266) );
NAND2_X1 U1051 ( .A1(G237), .A2(G234), .ZN(n1094) );
XNOR2_X1 U1052 ( .A(n1230), .B(KEYINPUT3), .ZN(n1053) );
NOR2_X1 U1053 ( .A1(n1093), .A2(n1092), .ZN(n1230) );
AND2_X1 U1054 ( .A1(G214), .A2(n1345), .ZN(n1092) );
INV_X1 U1055 ( .A(n1260), .ZN(n1093) );
XNOR2_X1 U1056 ( .A(n1346), .B(n1219), .ZN(n1260) );
AND2_X1 U1057 ( .A1(G210), .A2(n1345), .ZN(n1219) );
NAND2_X1 U1058 ( .A1(n1347), .A2(n1286), .ZN(n1345) );
INV_X1 U1059 ( .A(G237), .ZN(n1347) );
NAND2_X1 U1060 ( .A1(n1348), .A2(n1286), .ZN(n1346) );
XOR2_X1 U1061 ( .A(n1251), .B(n1250), .Z(n1348) );
XNOR2_X1 U1062 ( .A(n1165), .B(n1349), .ZN(n1250) );
NOR2_X1 U1063 ( .A1(KEYINPUT59), .A2(n1163), .ZN(n1349) );
XOR2_X1 U1064 ( .A(n1350), .B(n1351), .Z(n1163) );
NOR3_X1 U1065 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1351) );
NOR2_X1 U1066 ( .A1(KEYINPUT6), .A2(n1355), .ZN(n1354) );
NOR3_X1 U1067 ( .A1(n1341), .A2(G107), .A3(n1356), .ZN(n1353) );
NOR2_X1 U1068 ( .A1(n1357), .A2(n1299), .ZN(n1352) );
INV_X1 U1069 ( .A(G107), .ZN(n1299) );
NOR2_X1 U1070 ( .A1(n1356), .A2(n1358), .ZN(n1357) );
XNOR2_X1 U1071 ( .A(KEYINPUT28), .B(n1355), .ZN(n1358) );
INV_X1 U1072 ( .A(n1341), .ZN(n1355) );
XOR2_X1 U1073 ( .A(G104), .B(KEYINPUT2), .Z(n1341) );
INV_X1 U1074 ( .A(KEYINPUT6), .ZN(n1356) );
XOR2_X1 U1075 ( .A(n1359), .B(G101), .Z(n1350) );
NAND2_X1 U1076 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
OR2_X1 U1077 ( .A1(n1362), .A2(G113), .ZN(n1361) );
XOR2_X1 U1078 ( .A(n1363), .B(KEYINPUT35), .Z(n1360) );
NAND2_X1 U1079 ( .A1(G113), .A2(n1362), .ZN(n1363) );
XNOR2_X1 U1080 ( .A(n1324), .B(KEYINPUT55), .ZN(n1362) );
XNOR2_X1 U1081 ( .A(G116), .B(n1364), .ZN(n1324) );
XOR2_X1 U1082 ( .A(KEYINPUT21), .B(G119), .Z(n1364) );
XNOR2_X1 U1083 ( .A(G110), .B(n1295), .ZN(n1165) );
XOR2_X1 U1084 ( .A(G122), .B(KEYINPUT60), .Z(n1295) );
XOR2_X1 U1085 ( .A(n1327), .B(n1365), .Z(n1251) );
XOR2_X1 U1086 ( .A(G125), .B(n1366), .Z(n1365) );
NOR2_X1 U1087 ( .A1(G953), .A2(n1167), .ZN(n1366) );
INV_X1 U1088 ( .A(G224), .ZN(n1167) );
XOR2_X1 U1089 ( .A(G143), .B(n1367), .Z(n1327) );
INV_X1 U1090 ( .A(n1269), .ZN(n1078) );
XOR2_X1 U1091 ( .A(n1368), .B(n1101), .Z(n1269) );
NAND2_X1 U1092 ( .A1(n1175), .A2(n1286), .ZN(n1101) );
XNOR2_X1 U1093 ( .A(n1369), .B(n1370), .ZN(n1175) );
XOR2_X1 U1094 ( .A(n1371), .B(n1372), .Z(n1370) );
XNOR2_X1 U1095 ( .A(G137), .B(n1373), .ZN(n1372) );
NOR2_X1 U1096 ( .A1(G119), .A2(KEYINPUT52), .ZN(n1373) );
NAND3_X1 U1097 ( .A1(G234), .A2(n1056), .A3(G221), .ZN(n1371) );
INV_X1 U1098 ( .A(G953), .ZN(n1056) );
XNOR2_X1 U1099 ( .A(n1342), .B(n1374), .ZN(n1369) );
XOR2_X1 U1100 ( .A(n1367), .B(n1308), .Z(n1374) );
XOR2_X1 U1101 ( .A(G125), .B(KEYINPUT23), .Z(n1308) );
XNOR2_X1 U1102 ( .A(n1294), .B(G146), .ZN(n1367) );
INV_X1 U1103 ( .A(G128), .ZN(n1294) );
XOR2_X1 U1104 ( .A(G110), .B(G140), .Z(n1342) );
NAND2_X1 U1105 ( .A1(KEYINPUT48), .A2(n1102), .ZN(n1368) );
NAND2_X1 U1106 ( .A1(G217), .A2(n1329), .ZN(n1102) );
NAND2_X1 U1107 ( .A1(G234), .A2(n1286), .ZN(n1329) );
INV_X1 U1108 ( .A(G902), .ZN(n1286) );
endmodule


