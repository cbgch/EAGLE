//Key = 0111101011110110010010000001100101100111101011011101110000100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298;

XOR2_X1 U705 ( .A(n981), .B(n982), .Z(G9) );
NAND2_X1 U706 ( .A1(KEYINPUT52), .A2(G107), .ZN(n982) );
NOR2_X1 U707 ( .A1(n983), .A2(n984), .ZN(G75) );
NOR3_X1 U708 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n984) );
NAND3_X1 U709 ( .A1(n988), .A2(n989), .A3(n990), .ZN(n985) );
NAND2_X1 U710 ( .A1(n991), .A2(n992), .ZN(n990) );
NAND2_X1 U711 ( .A1(n993), .A2(n994), .ZN(n992) );
NAND3_X1 U712 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n994) );
NAND2_X1 U713 ( .A1(n998), .A2(n999), .ZN(n996) );
NAND2_X1 U714 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NAND2_X1 U715 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NAND2_X1 U716 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NAND2_X1 U717 ( .A1(n1006), .A2(n1007), .ZN(n998) );
XNOR2_X1 U718 ( .A(n1008), .B(KEYINPUT53), .ZN(n1006) );
NAND2_X1 U719 ( .A1(n1008), .A2(n1009), .ZN(n993) );
NAND2_X1 U720 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND3_X1 U721 ( .A1(n1012), .A2(n995), .A3(n997), .ZN(n1011) );
NAND2_X1 U722 ( .A1(n1000), .A2(n1013), .ZN(n1010) );
NAND3_X1 U723 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NAND2_X1 U724 ( .A1(n997), .A2(n1017), .ZN(n1016) );
NAND2_X1 U725 ( .A1(n1018), .A2(n1019), .ZN(n1015) );
XOR2_X1 U726 ( .A(KEYINPUT57), .B(n997), .Z(n1019) );
NAND2_X1 U727 ( .A1(n995), .A2(n1020), .ZN(n1014) );
NAND2_X1 U728 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U729 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
XNOR2_X1 U730 ( .A(KEYINPUT21), .B(n1025), .ZN(n1021) );
INV_X1 U731 ( .A(n1026), .ZN(n991) );
NOR3_X1 U732 ( .A1(n1027), .A2(G953), .A3(G952), .ZN(n983) );
INV_X1 U733 ( .A(n988), .ZN(n1027) );
NAND4_X1 U734 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n988) );
NOR4_X1 U735 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
NOR3_X1 U736 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1030) );
XOR2_X1 U737 ( .A(n1039), .B(n1040), .Z(G72) );
NOR2_X1 U738 ( .A1(n1041), .A2(n989), .ZN(n1040) );
AND2_X1 U739 ( .A1(G227), .A2(G900), .ZN(n1041) );
NAND2_X1 U740 ( .A1(n1042), .A2(n1043), .ZN(n1039) );
OR3_X1 U741 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
XOR2_X1 U742 ( .A(KEYINPUT51), .B(n1047), .Z(n1042) );
NOR2_X1 U743 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XOR2_X1 U744 ( .A(KEYINPUT33), .B(n1050), .Z(n1049) );
AND2_X1 U745 ( .A1(n1046), .A2(n989), .ZN(n1050) );
NAND2_X1 U746 ( .A1(n1051), .A2(n1052), .ZN(n1046) );
NOR2_X1 U747 ( .A1(n1045), .A2(n1044), .ZN(n1048) );
XNOR2_X1 U748 ( .A(n1053), .B(n1054), .ZN(n1044) );
XOR2_X1 U749 ( .A(n1055), .B(n1056), .Z(n1054) );
XNOR2_X1 U750 ( .A(G131), .B(G137), .ZN(n1056) );
NAND2_X1 U751 ( .A1(KEYINPUT14), .A2(n1057), .ZN(n1055) );
XNOR2_X1 U752 ( .A(KEYINPUT41), .B(n1058), .ZN(n1057) );
XOR2_X1 U753 ( .A(n1059), .B(n1060), .Z(n1053) );
NAND2_X1 U754 ( .A1(n1061), .A2(n1062), .ZN(G69) );
NAND2_X1 U755 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U756 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
OR2_X1 U757 ( .A1(n989), .A2(G224), .ZN(n1066) );
INV_X1 U758 ( .A(n1067), .ZN(n1063) );
NAND2_X1 U759 ( .A1(n1068), .A2(n1067), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NAND3_X1 U761 ( .A1(n1071), .A2(n1065), .A3(n1072), .ZN(n1070) );
INV_X1 U762 ( .A(n1073), .ZN(n1065) );
NAND2_X1 U763 ( .A1(KEYINPUT11), .A2(n987), .ZN(n1071) );
NAND3_X1 U764 ( .A1(n1074), .A2(n1075), .A3(n987), .ZN(n1069) );
NAND2_X1 U765 ( .A1(KEYINPUT11), .A2(G953), .ZN(n1075) );
NAND2_X1 U766 ( .A1(n1076), .A2(n989), .ZN(n1074) );
NAND2_X1 U767 ( .A1(n1077), .A2(KEYINPUT11), .ZN(n1076) );
INV_X1 U768 ( .A(n1072), .ZN(n1077) );
XNOR2_X1 U769 ( .A(n1078), .B(KEYINPUT12), .ZN(n1072) );
NAND3_X1 U770 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NAND2_X1 U771 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U772 ( .A1(n1084), .A2(KEYINPUT44), .ZN(n1083) );
XNOR2_X1 U773 ( .A(n1085), .B(KEYINPUT2), .ZN(n1084) );
INV_X1 U774 ( .A(n1086), .ZN(n1082) );
NAND3_X1 U775 ( .A1(KEYINPUT44), .A2(n1086), .A3(n1085), .ZN(n1080) );
XNOR2_X1 U776 ( .A(n1087), .B(n1088), .ZN(n1086) );
NAND2_X1 U777 ( .A1(KEYINPUT42), .A2(n1089), .ZN(n1087) );
XOR2_X1 U778 ( .A(KEYINPUT30), .B(n1090), .Z(n1089) );
OR2_X1 U779 ( .A1(n1085), .A2(KEYINPUT44), .ZN(n1079) );
NAND2_X1 U780 ( .A1(G953), .A2(n1091), .ZN(n1068) );
NAND2_X1 U781 ( .A1(G898), .A2(G224), .ZN(n1091) );
NOR3_X1 U782 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(G66) );
NOR2_X1 U783 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XOR2_X1 U784 ( .A(KEYINPUT37), .B(n1097), .Z(n1096) );
INV_X1 U785 ( .A(n1098), .ZN(n1095) );
NOR2_X1 U786 ( .A1(n1098), .A2(n1099), .ZN(n1093) );
XNOR2_X1 U787 ( .A(n1097), .B(KEYINPUT38), .ZN(n1099) );
NOR2_X1 U788 ( .A1(n1100), .A2(n1101), .ZN(n1097) );
NOR2_X1 U789 ( .A1(n1092), .A2(n1102), .ZN(G63) );
XOR2_X1 U790 ( .A(n1103), .B(n1104), .Z(n1102) );
AND2_X1 U791 ( .A1(G478), .A2(n1105), .ZN(n1104) );
NAND2_X1 U792 ( .A1(KEYINPUT9), .A2(n1106), .ZN(n1103) );
NOR2_X1 U793 ( .A1(n1092), .A2(n1107), .ZN(G60) );
XOR2_X1 U794 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U795 ( .A1(n1105), .A2(G475), .ZN(n1108) );
XNOR2_X1 U796 ( .A(n1110), .B(n1111), .ZN(G6) );
XOR2_X1 U797 ( .A(KEYINPUT47), .B(G104), .Z(n1111) );
NOR2_X1 U798 ( .A1(n1112), .A2(n1113), .ZN(G57) );
XOR2_X1 U799 ( .A(n1114), .B(n1115), .Z(n1113) );
XNOR2_X1 U800 ( .A(n1116), .B(n1117), .ZN(n1115) );
XOR2_X1 U801 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U802 ( .A(n1120), .B(n1121), .Z(n1114) );
XOR2_X1 U803 ( .A(n1122), .B(n1123), .Z(n1121) );
AND2_X1 U804 ( .A1(G472), .A2(n1105), .ZN(n1123) );
NOR2_X1 U805 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
XOR2_X1 U806 ( .A(KEYINPUT50), .B(KEYINPUT31), .Z(n1120) );
NOR2_X1 U807 ( .A1(n1126), .A2(n989), .ZN(n1112) );
XNOR2_X1 U808 ( .A(G952), .B(KEYINPUT1), .ZN(n1126) );
NOR2_X1 U809 ( .A1(n1092), .A2(n1127), .ZN(G54) );
XOR2_X1 U810 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U811 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U812 ( .A1(KEYINPUT48), .A2(n1132), .ZN(n1130) );
XOR2_X1 U813 ( .A(n1133), .B(n1134), .Z(n1128) );
XOR2_X1 U814 ( .A(n1135), .B(G140), .Z(n1134) );
NAND2_X1 U815 ( .A1(n1105), .A2(G469), .ZN(n1133) );
INV_X1 U816 ( .A(n1100), .ZN(n1105) );
NOR2_X1 U817 ( .A1(n1092), .A2(n1136), .ZN(G51) );
XOR2_X1 U818 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U819 ( .A1(n1100), .A2(n1139), .ZN(n1138) );
XOR2_X1 U820 ( .A(KEYINPUT39), .B(n1140), .Z(n1139) );
NAND2_X1 U821 ( .A1(G902), .A2(n1141), .ZN(n1100) );
NAND2_X1 U822 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XNOR2_X1 U823 ( .A(KEYINPUT46), .B(n987), .ZN(n1143) );
NAND4_X1 U824 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n987) );
AND4_X1 U825 ( .A1(n981), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1147) );
NAND3_X1 U826 ( .A1(n1000), .A2(n1151), .A3(n1017), .ZN(n981) );
NOR2_X1 U827 ( .A1(n1110), .A2(n1152), .ZN(n1146) );
NOR2_X1 U828 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
AND3_X1 U829 ( .A1(n1000), .A2(n1151), .A3(n1018), .ZN(n1110) );
INV_X1 U830 ( .A(n986), .ZN(n1142) );
NAND2_X1 U831 ( .A1(n1155), .A2(n1051), .ZN(n986) );
AND4_X1 U832 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1051) );
AND4_X1 U833 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1159) );
NAND4_X1 U834 ( .A1(n1164), .A2(n1018), .A3(n1012), .A4(n1165), .ZN(n1158) );
XOR2_X1 U835 ( .A(KEYINPUT19), .B(n997), .Z(n1165) );
XOR2_X1 U836 ( .A(n1052), .B(KEYINPUT54), .Z(n1155) );
NOR2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(n1137) );
XOR2_X1 U838 ( .A(KEYINPUT26), .B(n1168), .Z(n1167) );
NOR2_X1 U839 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
AND2_X1 U840 ( .A1(n1170), .A2(n1169), .ZN(n1166) );
XOR2_X1 U841 ( .A(n1171), .B(n1172), .Z(n1169) );
XOR2_X1 U842 ( .A(n1173), .B(KEYINPUT24), .Z(n1170) );
NOR2_X1 U843 ( .A1(n989), .A2(G952), .ZN(n1092) );
XNOR2_X1 U844 ( .A(G146), .B(n1156), .ZN(G48) );
NAND4_X1 U845 ( .A1(n1164), .A2(n1174), .A3(n1025), .A4(n1018), .ZN(n1156) );
XOR2_X1 U846 ( .A(n1157), .B(n1175), .Z(G45) );
NAND2_X1 U847 ( .A1(KEYINPUT34), .A2(G143), .ZN(n1175) );
NAND4_X1 U848 ( .A1(n1025), .A2(n1164), .A3(n1176), .A4(n1007), .ZN(n1157) );
NOR2_X1 U849 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XOR2_X1 U850 ( .A(G140), .B(n1179), .Z(G42) );
AND2_X1 U851 ( .A1(n1012), .A2(n1180), .ZN(n1179) );
XNOR2_X1 U852 ( .A(G137), .B(n1163), .ZN(G39) );
NAND3_X1 U853 ( .A1(n1174), .A2(n995), .A3(n1181), .ZN(n1163) );
XNOR2_X1 U854 ( .A(G134), .B(n1162), .ZN(G36) );
NAND3_X1 U855 ( .A1(n1007), .A2(n1017), .A3(n1181), .ZN(n1162) );
XOR2_X1 U856 ( .A(n1052), .B(n1182), .Z(G33) );
NAND2_X1 U857 ( .A1(KEYINPUT28), .A2(G131), .ZN(n1182) );
NAND2_X1 U858 ( .A1(n1180), .A2(n1007), .ZN(n1052) );
AND2_X1 U859 ( .A1(n1181), .A2(n1018), .ZN(n1180) );
AND2_X1 U860 ( .A1(n1164), .A2(n997), .ZN(n1181) );
AND2_X1 U861 ( .A1(n1023), .A2(n1029), .ZN(n997) );
XNOR2_X1 U862 ( .A(n1035), .B(KEYINPUT59), .ZN(n1023) );
AND2_X1 U863 ( .A1(n1183), .A2(n1184), .ZN(n1164) );
NAND2_X1 U864 ( .A1(n1185), .A2(n1186), .ZN(G30) );
OR2_X1 U865 ( .A1(n1161), .A2(G128), .ZN(n1186) );
XOR2_X1 U866 ( .A(n1187), .B(KEYINPUT16), .Z(n1185) );
NAND2_X1 U867 ( .A1(G128), .A2(n1161), .ZN(n1187) );
NAND4_X1 U868 ( .A1(n1188), .A2(n1174), .A3(n1017), .A4(n1189), .ZN(n1161) );
XOR2_X1 U869 ( .A(n1190), .B(n1191), .Z(G3) );
NOR2_X1 U870 ( .A1(KEYINPUT23), .A2(n1192), .ZN(n1191) );
NOR2_X1 U871 ( .A1(n1153), .A2(n1193), .ZN(n1190) );
XNOR2_X1 U872 ( .A(KEYINPUT62), .B(n1154), .ZN(n1193) );
NAND4_X1 U873 ( .A1(n1007), .A2(n995), .A3(n1189), .A4(n1194), .ZN(n1154) );
XNOR2_X1 U874 ( .A(G125), .B(n1160), .ZN(G27) );
NAND4_X1 U875 ( .A1(n1188), .A2(n1018), .A3(n1012), .A4(n1008), .ZN(n1160) );
INV_X1 U876 ( .A(n1034), .ZN(n1008) );
AND2_X1 U877 ( .A1(n1025), .A2(n1184), .ZN(n1188) );
NAND2_X1 U878 ( .A1(n1026), .A2(n1195), .ZN(n1184) );
NAND2_X1 U879 ( .A1(n1045), .A2(n1196), .ZN(n1195) );
NOR2_X1 U880 ( .A1(n989), .A2(G900), .ZN(n1045) );
INV_X1 U881 ( .A(n1197), .ZN(n1025) );
XOR2_X1 U882 ( .A(n1144), .B(n1198), .Z(G24) );
NAND2_X1 U883 ( .A1(KEYINPUT3), .A2(G122), .ZN(n1198) );
NAND4_X1 U884 ( .A1(n1199), .A2(n1000), .A3(n1200), .A4(n1033), .ZN(n1144) );
INV_X1 U885 ( .A(n1178), .ZN(n1200) );
NOR2_X1 U886 ( .A1(n1201), .A2(n1032), .ZN(n1000) );
XNOR2_X1 U887 ( .A(n1145), .B(n1202), .ZN(G21) );
NOR2_X1 U888 ( .A1(KEYINPUT36), .A2(n1203), .ZN(n1202) );
NAND3_X1 U889 ( .A1(n1199), .A2(n995), .A3(n1174), .ZN(n1145) );
AND2_X1 U890 ( .A1(n1032), .A2(n1201), .ZN(n1174) );
XNOR2_X1 U891 ( .A(G116), .B(n1150), .ZN(G18) );
NAND3_X1 U892 ( .A1(n1007), .A2(n1017), .A3(n1199), .ZN(n1150) );
NOR3_X1 U893 ( .A1(n1034), .A2(n1204), .A3(n1197), .ZN(n1199) );
XOR2_X1 U894 ( .A(n1205), .B(KEYINPUT49), .Z(n1197) );
NOR2_X1 U895 ( .A1(n1033), .A2(n1178), .ZN(n1017) );
XOR2_X1 U896 ( .A(n1206), .B(KEYINPUT60), .Z(n1178) );
XNOR2_X1 U897 ( .A(G113), .B(n1149), .ZN(G15) );
NAND3_X1 U898 ( .A1(n1007), .A2(n1018), .A3(n1207), .ZN(n1149) );
NOR3_X1 U899 ( .A1(n1034), .A2(n1204), .A3(n1153), .ZN(n1207) );
INV_X1 U900 ( .A(n1205), .ZN(n1153) );
INV_X1 U901 ( .A(n1194), .ZN(n1204) );
NAND2_X1 U902 ( .A1(n1005), .A2(n1208), .ZN(n1034) );
AND2_X1 U903 ( .A1(n1206), .A2(n1033), .ZN(n1018) );
AND2_X1 U904 ( .A1(n1209), .A2(n1032), .ZN(n1007) );
XNOR2_X1 U905 ( .A(n1132), .B(n1210), .ZN(G12) );
NOR2_X1 U906 ( .A1(KEYINPUT18), .A2(n1148), .ZN(n1210) );
NAND3_X1 U907 ( .A1(n995), .A2(n1151), .A3(n1012), .ZN(n1148) );
NOR2_X1 U908 ( .A1(n1032), .A2(n1209), .ZN(n1012) );
INV_X1 U909 ( .A(n1201), .ZN(n1209) );
NAND2_X1 U910 ( .A1(n1211), .A2(n1028), .ZN(n1201) );
NAND2_X1 U911 ( .A1(n1212), .A2(n1213), .ZN(n1028) );
XOR2_X1 U912 ( .A(KEYINPUT20), .B(n1037), .Z(n1211) );
NOR2_X1 U913 ( .A1(n1213), .A2(n1212), .ZN(n1037) );
INV_X1 U914 ( .A(n1101), .ZN(n1212) );
NAND2_X1 U915 ( .A1(G217), .A2(n1214), .ZN(n1101) );
NAND2_X1 U916 ( .A1(n1098), .A2(n1215), .ZN(n1213) );
XNOR2_X1 U917 ( .A(n1216), .B(n1217), .ZN(n1098) );
NOR2_X1 U918 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
INV_X1 U919 ( .A(G221), .ZN(n1219) );
XOR2_X1 U920 ( .A(n1220), .B(G137), .Z(n1216) );
NAND2_X1 U921 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NAND2_X1 U922 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
NAND2_X1 U923 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
NAND2_X1 U924 ( .A1(KEYINPUT4), .A2(n1227), .ZN(n1226) );
INV_X1 U925 ( .A(n1228), .ZN(n1227) );
INV_X1 U926 ( .A(KEYINPUT29), .ZN(n1225) );
NAND2_X1 U927 ( .A1(n1228), .A2(n1229), .ZN(n1221) );
NAND2_X1 U928 ( .A1(KEYINPUT4), .A2(n1230), .ZN(n1229) );
OR2_X1 U929 ( .A1(n1223), .A2(KEYINPUT29), .ZN(n1230) );
XOR2_X1 U930 ( .A(n1231), .B(KEYINPUT17), .Z(n1223) );
XOR2_X1 U931 ( .A(G110), .B(n1232), .Z(n1228) );
XNOR2_X1 U932 ( .A(G128), .B(n1203), .ZN(n1232) );
XNOR2_X1 U933 ( .A(n1233), .B(G472), .ZN(n1032) );
NAND2_X1 U934 ( .A1(n1234), .A2(n1215), .ZN(n1233) );
XOR2_X1 U935 ( .A(n1235), .B(n1236), .Z(n1234) );
XOR2_X1 U936 ( .A(KEYINPUT61), .B(n1237), .Z(n1236) );
NOR2_X1 U937 ( .A1(n1124), .A2(n1238), .ZN(n1237) );
XNOR2_X1 U938 ( .A(n1125), .B(KEYINPUT27), .ZN(n1238) );
AND2_X1 U939 ( .A1(n1192), .A2(n1239), .ZN(n1125) );
NAND2_X1 U940 ( .A1(G210), .A2(n1240), .ZN(n1239) );
AND3_X1 U941 ( .A1(G101), .A2(n1240), .A3(G210), .ZN(n1124) );
XNOR2_X1 U942 ( .A(n1241), .B(n1242), .ZN(n1235) );
INV_X1 U943 ( .A(n1116), .ZN(n1242) );
XOR2_X1 U944 ( .A(n1090), .B(KEYINPUT32), .Z(n1116) );
NAND2_X1 U945 ( .A1(n1243), .A2(n1244), .ZN(n1241) );
NAND2_X1 U946 ( .A1(n1118), .A2(n1119), .ZN(n1244) );
XOR2_X1 U947 ( .A(KEYINPUT10), .B(n1245), .Z(n1243) );
NOR2_X1 U948 ( .A1(n1118), .A2(n1119), .ZN(n1245) );
AND3_X1 U949 ( .A1(n1189), .A2(n1194), .A3(n1205), .ZN(n1151) );
NOR2_X1 U950 ( .A1(n1246), .A2(n1024), .ZN(n1205) );
INV_X1 U951 ( .A(n1029), .ZN(n1024) );
NAND2_X1 U952 ( .A1(G214), .A2(n1247), .ZN(n1029) );
INV_X1 U953 ( .A(n1035), .ZN(n1246) );
XNOR2_X1 U954 ( .A(n1248), .B(n1140), .ZN(n1035) );
AND2_X1 U955 ( .A1(G210), .A2(n1247), .ZN(n1140) );
NAND2_X1 U956 ( .A1(n1249), .A2(n1215), .ZN(n1247) );
INV_X1 U957 ( .A(G237), .ZN(n1249) );
NAND2_X1 U958 ( .A1(n1250), .A2(n1215), .ZN(n1248) );
XNOR2_X1 U959 ( .A(n1251), .B(n1252), .ZN(n1250) );
XOR2_X1 U960 ( .A(n1171), .B(n1253), .Z(n1252) );
NOR2_X1 U961 ( .A1(KEYINPUT35), .A2(n1172), .ZN(n1253) );
XOR2_X1 U962 ( .A(G125), .B(n1118), .Z(n1172) );
XOR2_X1 U963 ( .A(n1059), .B(KEYINPUT8), .Z(n1118) );
AND2_X1 U964 ( .A1(G224), .A2(n989), .ZN(n1171) );
INV_X1 U965 ( .A(n1173), .ZN(n1251) );
XOR2_X1 U966 ( .A(n1085), .B(n1254), .Z(n1173) );
XOR2_X1 U967 ( .A(n1088), .B(n1090), .Z(n1254) );
XNOR2_X1 U968 ( .A(n1255), .B(n1256), .ZN(n1090) );
XNOR2_X1 U969 ( .A(KEYINPUT58), .B(n1203), .ZN(n1256) );
INV_X1 U970 ( .A(G119), .ZN(n1203) );
XNOR2_X1 U971 ( .A(G113), .B(G116), .ZN(n1255) );
XNOR2_X1 U972 ( .A(n1257), .B(n1258), .ZN(n1088) );
NOR2_X1 U973 ( .A1(KEYINPUT43), .A2(G104), .ZN(n1258) );
XNOR2_X1 U974 ( .A(G101), .B(G107), .ZN(n1257) );
XNOR2_X1 U975 ( .A(n1259), .B(n1260), .ZN(n1085) );
XNOR2_X1 U976 ( .A(G122), .B(n1132), .ZN(n1260) );
XNOR2_X1 U977 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n1259) );
NAND2_X1 U978 ( .A1(n1026), .A2(n1261), .ZN(n1194) );
NAND2_X1 U979 ( .A1(n1073), .A2(n1196), .ZN(n1261) );
AND2_X1 U980 ( .A1(n1262), .A2(n1263), .ZN(n1196) );
XNOR2_X1 U981 ( .A(G902), .B(KEYINPUT45), .ZN(n1262) );
NOR2_X1 U982 ( .A1(n989), .A2(G898), .ZN(n1073) );
NAND3_X1 U983 ( .A1(n1263), .A2(n989), .A3(G952), .ZN(n1026) );
NAND2_X1 U984 ( .A1(G237), .A2(G234), .ZN(n1263) );
XNOR2_X1 U985 ( .A(n1002), .B(KEYINPUT22), .ZN(n1189) );
INV_X1 U986 ( .A(n1183), .ZN(n1002) );
NOR2_X1 U987 ( .A1(n1005), .A2(n1004), .ZN(n1183) );
INV_X1 U988 ( .A(n1208), .ZN(n1004) );
NAND2_X1 U989 ( .A1(G221), .A2(n1214), .ZN(n1208) );
NAND2_X1 U990 ( .A1(G234), .A2(n1215), .ZN(n1214) );
XOR2_X1 U991 ( .A(n1264), .B(G469), .Z(n1005) );
NAND2_X1 U992 ( .A1(n1265), .A2(n1215), .ZN(n1264) );
XOR2_X1 U993 ( .A(n1266), .B(n1267), .Z(n1265) );
XNOR2_X1 U994 ( .A(n1132), .B(n1268), .ZN(n1267) );
NOR2_X1 U995 ( .A1(G140), .A2(KEYINPUT0), .ZN(n1268) );
XOR2_X1 U996 ( .A(n1135), .B(n1269), .Z(n1266) );
NOR2_X1 U997 ( .A1(KEYINPUT63), .A2(n1131), .ZN(n1269) );
XOR2_X1 U998 ( .A(n1270), .B(n1271), .Z(n1131) );
XOR2_X1 U999 ( .A(n1272), .B(n1273), .Z(n1271) );
XNOR2_X1 U1000 ( .A(G104), .B(n1192), .ZN(n1273) );
INV_X1 U1001 ( .A(G101), .ZN(n1192) );
NOR2_X1 U1002 ( .A1(KEYINPUT15), .A2(n1274), .ZN(n1272) );
INV_X1 U1003 ( .A(G107), .ZN(n1274) );
XOR2_X1 U1004 ( .A(n1059), .B(n1119), .Z(n1270) );
XNOR2_X1 U1005 ( .A(n1275), .B(n1276), .ZN(n1119) );
NOR2_X1 U1006 ( .A1(KEYINPUT56), .A2(n1277), .ZN(n1276) );
XNOR2_X1 U1007 ( .A(G134), .B(G137), .ZN(n1275) );
XOR2_X1 U1008 ( .A(G146), .B(n1278), .Z(n1059) );
NAND2_X1 U1009 ( .A1(n1279), .A2(n989), .ZN(n1135) );
XOR2_X1 U1010 ( .A(KEYINPUT7), .B(G227), .Z(n1279) );
AND2_X1 U1011 ( .A1(n1177), .A2(n1206), .ZN(n995) );
NOR2_X1 U1012 ( .A1(n1280), .A2(n1038), .ZN(n1206) );
NOR2_X1 U1013 ( .A1(n1281), .A2(G478), .ZN(n1038) );
XNOR2_X1 U1014 ( .A(KEYINPUT40), .B(n1036), .ZN(n1280) );
AND2_X1 U1015 ( .A1(G478), .A2(n1281), .ZN(n1036) );
NAND2_X1 U1016 ( .A1(n1106), .A2(n1215), .ZN(n1281) );
XNOR2_X1 U1017 ( .A(n1282), .B(n1283), .ZN(n1106) );
XOR2_X1 U1018 ( .A(G116), .B(n1284), .Z(n1283) );
XNOR2_X1 U1019 ( .A(n1058), .B(G122), .ZN(n1284) );
INV_X1 U1020 ( .A(G134), .ZN(n1058) );
XOR2_X1 U1021 ( .A(n1285), .B(n1286), .Z(n1282) );
NOR2_X1 U1022 ( .A1(n1218), .A2(n1287), .ZN(n1286) );
INV_X1 U1023 ( .A(G217), .ZN(n1287) );
NAND2_X1 U1024 ( .A1(G234), .A2(n989), .ZN(n1218) );
INV_X1 U1025 ( .A(G953), .ZN(n989) );
XNOR2_X1 U1026 ( .A(G107), .B(n1288), .ZN(n1285) );
NOR2_X1 U1027 ( .A1(KEYINPUT55), .A2(n1278), .ZN(n1288) );
XNOR2_X1 U1028 ( .A(G143), .B(G128), .ZN(n1278) );
INV_X1 U1029 ( .A(n1033), .ZN(n1177) );
XNOR2_X1 U1030 ( .A(n1289), .B(G475), .ZN(n1033) );
NAND2_X1 U1031 ( .A1(n1109), .A2(n1215), .ZN(n1289) );
INV_X1 U1032 ( .A(G902), .ZN(n1215) );
XOR2_X1 U1033 ( .A(n1290), .B(n1291), .Z(n1109) );
XNOR2_X1 U1034 ( .A(G122), .B(n1292), .ZN(n1291) );
INV_X1 U1035 ( .A(G113), .ZN(n1292) );
XOR2_X1 U1036 ( .A(n1293), .B(G104), .Z(n1290) );
NAND2_X1 U1037 ( .A1(KEYINPUT13), .A2(n1294), .ZN(n1293) );
XOR2_X1 U1038 ( .A(n1231), .B(n1295), .Z(n1294) );
XNOR2_X1 U1039 ( .A(n1277), .B(n1296), .ZN(n1295) );
NOR2_X1 U1040 ( .A1(KEYINPUT25), .A2(n1297), .ZN(n1296) );
XNOR2_X1 U1041 ( .A(G143), .B(n1298), .ZN(n1297) );
NAND2_X1 U1042 ( .A1(G214), .A2(n1240), .ZN(n1298) );
NOR2_X1 U1043 ( .A1(G953), .A2(G237), .ZN(n1240) );
INV_X1 U1044 ( .A(G131), .ZN(n1277) );
XOR2_X1 U1045 ( .A(G146), .B(n1060), .Z(n1231) );
XOR2_X1 U1046 ( .A(G125), .B(G140), .Z(n1060) );
INV_X1 U1047 ( .A(G110), .ZN(n1132) );
endmodule


