//Key = 0111011100110001101100010011010100110100010000100000000100010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435;

XNOR2_X1 U758 ( .A(n1076), .B(n1077), .ZN(G9) );
NOR2_X1 U759 ( .A1(n1078), .A2(n1079), .ZN(G75) );
NOR3_X1 U760 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NOR2_X1 U761 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
INV_X1 U762 ( .A(n1085), .ZN(n1084) );
NOR2_X1 U763 ( .A1(n1086), .A2(n1087), .ZN(n1083) );
NOR2_X1 U764 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
INV_X1 U765 ( .A(KEYINPUT42), .ZN(n1089) );
NOR4_X1 U766 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1088) );
NOR2_X1 U767 ( .A1(n1094), .A2(n1093), .ZN(n1086) );
NOR2_X1 U768 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U769 ( .A1(n1097), .A2(n1092), .ZN(n1096) );
NOR2_X1 U770 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U771 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U772 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR3_X1 U773 ( .A1(n1091), .A2(KEYINPUT42), .A3(n1090), .ZN(n1098) );
INV_X1 U774 ( .A(n1104), .ZN(n1090) );
NOR3_X1 U775 ( .A1(n1091), .A2(n1105), .A3(n1101), .ZN(n1095) );
INV_X1 U776 ( .A(n1106), .ZN(n1101) );
INV_X1 U777 ( .A(n1107), .ZN(n1091) );
NAND3_X1 U778 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1080) );
NAND3_X1 U779 ( .A1(n1111), .A2(n1112), .A3(n1107), .ZN(n1110) );
NAND2_X1 U780 ( .A1(n1113), .A2(n1093), .ZN(n1112) );
NAND2_X1 U781 ( .A1(KEYINPUT58), .A2(n1114), .ZN(n1113) );
NAND3_X1 U782 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1111) );
INV_X1 U783 ( .A(n1093), .ZN(n1117) );
NAND2_X1 U784 ( .A1(n1114), .A2(n1118), .ZN(n1116) );
INV_X1 U785 ( .A(KEYINPUT58), .ZN(n1118) );
AND4_X1 U786 ( .A1(n1119), .A2(n1085), .A3(n1106), .A4(n1120), .ZN(n1114) );
NAND2_X1 U787 ( .A1(n1121), .A2(n1122), .ZN(n1115) );
NAND2_X1 U788 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U789 ( .A1(n1106), .A2(n1125), .ZN(n1124) );
NAND2_X1 U790 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U791 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U792 ( .A1(n1130), .A2(n1085), .ZN(n1123) );
NOR3_X1 U793 ( .A1(n1131), .A2(G953), .A3(G952), .ZN(n1078) );
INV_X1 U794 ( .A(n1108), .ZN(n1131) );
NAND4_X1 U795 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1108) );
NOR4_X1 U796 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1135) );
XNOR2_X1 U797 ( .A(n1140), .B(n1141), .ZN(n1139) );
XNOR2_X1 U798 ( .A(G472), .B(n1142), .ZN(n1138) );
XOR2_X1 U799 ( .A(KEYINPUT43), .B(n1143), .Z(n1137) );
AND2_X1 U800 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NOR3_X1 U801 ( .A1(n1146), .A2(n1120), .A3(n1129), .ZN(n1134) );
NOR2_X1 U802 ( .A1(n1145), .A2(n1144), .ZN(n1146) );
XNOR2_X1 U803 ( .A(n1147), .B(n1148), .ZN(n1133) );
XNOR2_X1 U804 ( .A(G475), .B(KEYINPUT61), .ZN(n1148) );
XNOR2_X1 U805 ( .A(KEYINPUT63), .B(n1128), .ZN(n1132) );
INV_X1 U806 ( .A(n1149), .ZN(n1128) );
XOR2_X1 U807 ( .A(n1150), .B(n1151), .Z(G72) );
XOR2_X1 U808 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U809 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U810 ( .A1(G953), .A2(n1156), .ZN(n1155) );
XOR2_X1 U811 ( .A(n1157), .B(n1158), .Z(n1154) );
XOR2_X1 U812 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR3_X1 U813 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1160) );
NOR2_X1 U814 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XNOR2_X1 U815 ( .A(G131), .B(n1166), .ZN(n1165) );
NOR3_X1 U816 ( .A1(G140), .A2(G131), .A3(n1166), .ZN(n1162) );
AND2_X1 U817 ( .A1(G131), .A2(n1167), .ZN(n1161) );
XNOR2_X1 U818 ( .A(G134), .B(n1168), .ZN(n1157) );
XNOR2_X1 U819 ( .A(KEYINPUT49), .B(n1169), .ZN(n1168) );
NAND2_X1 U820 ( .A1(n1170), .A2(n1171), .ZN(n1152) );
NAND2_X1 U821 ( .A1(G900), .A2(G227), .ZN(n1171) );
NOR2_X1 U822 ( .A1(n1172), .A2(G953), .ZN(n1150) );
AND2_X1 U823 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U824 ( .A(n1175), .B(n1176), .Z(G69) );
NAND2_X1 U825 ( .A1(KEYINPUT27), .A2(n1177), .ZN(n1176) );
XOR2_X1 U826 ( .A(n1178), .B(n1179), .Z(n1177) );
NOR2_X1 U827 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XNOR2_X1 U828 ( .A(KEYINPUT8), .B(n1109), .ZN(n1181) );
NOR2_X1 U829 ( .A1(n1182), .A2(n1183), .ZN(n1178) );
XOR2_X1 U830 ( .A(n1184), .B(n1185), .Z(n1183) );
NAND2_X1 U831 ( .A1(n1170), .A2(n1186), .ZN(n1175) );
XOR2_X1 U832 ( .A(KEYINPUT11), .B(n1187), .Z(n1186) );
AND2_X1 U833 ( .A1(G224), .A2(G898), .ZN(n1187) );
XNOR2_X1 U834 ( .A(G953), .B(KEYINPUT1), .ZN(n1170) );
NOR2_X1 U835 ( .A1(n1188), .A2(n1189), .ZN(G66) );
NOR3_X1 U836 ( .A1(n1145), .A2(n1190), .A3(n1191), .ZN(n1189) );
NOR2_X1 U837 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NOR2_X1 U838 ( .A1(n1194), .A2(n1144), .ZN(n1192) );
NOR3_X1 U839 ( .A1(n1195), .A2(n1144), .A3(n1196), .ZN(n1190) );
INV_X1 U840 ( .A(n1193), .ZN(n1195) );
NOR2_X1 U841 ( .A1(n1188), .A2(n1197), .ZN(G63) );
NOR3_X1 U842 ( .A1(n1141), .A2(n1198), .A3(n1199), .ZN(n1197) );
NOR3_X1 U843 ( .A1(n1200), .A2(n1140), .A3(n1196), .ZN(n1199) );
INV_X1 U844 ( .A(n1201), .ZN(n1200) );
NOR2_X1 U845 ( .A1(n1202), .A2(n1201), .ZN(n1198) );
NOR2_X1 U846 ( .A1(n1194), .A2(n1140), .ZN(n1202) );
NOR2_X1 U847 ( .A1(n1188), .A2(n1203), .ZN(G60) );
NOR3_X1 U848 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1203) );
NOR2_X1 U849 ( .A1(KEYINPUT23), .A2(n1207), .ZN(n1206) );
NOR2_X1 U850 ( .A1(n1208), .A2(n1209), .ZN(n1205) );
NOR2_X1 U851 ( .A1(n1210), .A2(n1147), .ZN(n1208) );
NOR2_X1 U852 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NOR2_X1 U853 ( .A1(n1194), .A2(n1213), .ZN(n1211) );
INV_X1 U854 ( .A(n1082), .ZN(n1194) );
NOR3_X1 U855 ( .A1(n1196), .A2(n1214), .A3(n1213), .ZN(n1204) );
NOR2_X1 U856 ( .A1(n1212), .A2(n1209), .ZN(n1214) );
INV_X1 U857 ( .A(KEYINPUT23), .ZN(n1209) );
XNOR2_X1 U858 ( .A(G104), .B(n1215), .ZN(G6) );
NOR2_X1 U859 ( .A1(n1216), .A2(KEYINPUT48), .ZN(n1215) );
NOR2_X1 U860 ( .A1(n1188), .A2(n1217), .ZN(G57) );
XOR2_X1 U861 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U862 ( .A(n1220), .B(n1221), .Z(n1219) );
NAND2_X1 U863 ( .A1(KEYINPUT62), .A2(n1222), .ZN(n1220) );
XOR2_X1 U864 ( .A(KEYINPUT14), .B(n1223), .Z(n1218) );
NOR2_X1 U865 ( .A1(n1224), .A2(n1196), .ZN(n1223) );
INV_X1 U866 ( .A(G472), .ZN(n1224) );
NOR2_X1 U867 ( .A1(n1188), .A2(n1225), .ZN(G54) );
XOR2_X1 U868 ( .A(n1226), .B(n1227), .Z(n1225) );
NOR2_X1 U869 ( .A1(n1228), .A2(n1196), .ZN(n1227) );
NOR2_X1 U870 ( .A1(KEYINPUT30), .A2(n1229), .ZN(n1226) );
XOR2_X1 U871 ( .A(n1230), .B(n1231), .Z(n1229) );
NOR2_X1 U872 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NOR3_X1 U873 ( .A1(n1234), .A2(KEYINPUT45), .A3(n1235), .ZN(n1233) );
INV_X1 U874 ( .A(n1236), .ZN(n1234) );
NOR2_X1 U875 ( .A1(n1236), .A2(n1237), .ZN(n1232) );
NOR2_X1 U876 ( .A1(n1238), .A2(n1235), .ZN(n1237) );
AND2_X1 U877 ( .A1(n1239), .A2(KEYINPUT45), .ZN(n1238) );
NOR2_X1 U878 ( .A1(KEYINPUT52), .A2(n1239), .ZN(n1236) );
XNOR2_X1 U879 ( .A(n1240), .B(n1164), .ZN(n1239) );
XNOR2_X1 U880 ( .A(n1241), .B(n1242), .ZN(n1230) );
NOR2_X1 U881 ( .A1(KEYINPUT39), .A2(n1243), .ZN(n1242) );
XOR2_X1 U882 ( .A(n1244), .B(n1245), .Z(n1243) );
NOR2_X1 U883 ( .A1(n1188), .A2(n1246), .ZN(G51) );
XOR2_X1 U884 ( .A(n1247), .B(n1248), .Z(n1246) );
NOR2_X1 U885 ( .A1(n1249), .A2(n1196), .ZN(n1248) );
NAND2_X1 U886 ( .A1(G902), .A2(n1082), .ZN(n1196) );
NAND4_X1 U887 ( .A1(n1174), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1082) );
OR2_X1 U888 ( .A1(n1180), .A2(KEYINPUT17), .ZN(n1252) );
AND2_X1 U889 ( .A1(n1253), .A2(n1254), .ZN(n1180) );
NAND2_X1 U890 ( .A1(KEYINPUT17), .A2(n1255), .ZN(n1251) );
NAND2_X1 U891 ( .A1(n1256), .A2(n1253), .ZN(n1255) );
AND4_X1 U892 ( .A1(n1257), .A2(n1258), .A3(n1259), .A4(n1260), .ZN(n1253) );
NOR4_X1 U893 ( .A1(n1261), .A2(n1216), .A3(n1077), .A4(n1262), .ZN(n1260) );
INV_X1 U894 ( .A(n1263), .ZN(n1262) );
AND3_X1 U895 ( .A1(n1102), .A2(n1106), .A3(n1264), .ZN(n1077) );
AND3_X1 U896 ( .A1(n1264), .A2(n1106), .A3(n1103), .ZN(n1216) );
OR2_X1 U897 ( .A1(n1265), .A2(KEYINPUT21), .ZN(n1259) );
NAND3_X1 U898 ( .A1(n1266), .A2(n1267), .A3(n1121), .ZN(n1258) );
NAND2_X1 U899 ( .A1(n1268), .A2(n1269), .ZN(n1266) );
NAND3_X1 U900 ( .A1(KEYINPUT21), .A2(n1107), .A3(n1270), .ZN(n1269) );
NOR3_X1 U901 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1270) );
NAND2_X1 U902 ( .A1(n1272), .A2(n1274), .ZN(n1257) );
XNOR2_X1 U903 ( .A(KEYINPUT57), .B(n1275), .ZN(n1274) );
INV_X1 U904 ( .A(n1254), .ZN(n1256) );
XNOR2_X1 U905 ( .A(KEYINPUT41), .B(n1173), .ZN(n1250) );
AND4_X1 U906 ( .A1(n1276), .A2(n1277), .A3(n1278), .A4(n1279), .ZN(n1174) );
AND4_X1 U907 ( .A1(n1280), .A2(n1281), .A3(n1282), .A4(n1283), .ZN(n1279) );
NAND3_X1 U908 ( .A1(n1284), .A2(n1272), .A3(n1103), .ZN(n1278) );
NAND4_X1 U909 ( .A1(n1104), .A2(n1085), .A3(n1285), .A4(n1102), .ZN(n1276) );
NOR2_X1 U910 ( .A1(KEYINPUT20), .A2(n1286), .ZN(n1247) );
XOR2_X1 U911 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U912 ( .A(n1289), .B(n1290), .Z(n1288) );
XNOR2_X1 U913 ( .A(KEYINPUT9), .B(n1166), .ZN(n1290) );
XOR2_X1 U914 ( .A(n1291), .B(n1292), .Z(n1287) );
XNOR2_X1 U915 ( .A(n1293), .B(n1244), .ZN(n1292) );
NOR2_X1 U916 ( .A1(n1109), .A2(G952), .ZN(n1188) );
XNOR2_X1 U917 ( .A(G146), .B(n1294), .ZN(G48) );
NAND3_X1 U918 ( .A1(n1103), .A2(n1284), .A3(n1295), .ZN(n1294) );
XNOR2_X1 U919 ( .A(n1272), .B(KEYINPUT19), .ZN(n1295) );
XNOR2_X1 U920 ( .A(G143), .B(n1277), .ZN(G45) );
NAND4_X1 U921 ( .A1(n1296), .A2(n1104), .A3(n1297), .A4(n1285), .ZN(n1277) );
NOR2_X1 U922 ( .A1(n1298), .A2(n1126), .ZN(n1297) );
NAND2_X1 U923 ( .A1(n1299), .A2(n1300), .ZN(G42) );
OR2_X1 U924 ( .A1(n1283), .A2(G140), .ZN(n1300) );
XOR2_X1 U925 ( .A(n1301), .B(KEYINPUT40), .Z(n1299) );
NAND2_X1 U926 ( .A1(G140), .A2(n1283), .ZN(n1301) );
NAND2_X1 U927 ( .A1(n1130), .A2(n1302), .ZN(n1283) );
XNOR2_X1 U928 ( .A(G137), .B(n1282), .ZN(G39) );
NAND3_X1 U929 ( .A1(n1085), .A2(n1284), .A3(n1107), .ZN(n1282) );
XNOR2_X1 U930 ( .A(G134), .B(n1303), .ZN(G36) );
NAND4_X1 U931 ( .A1(n1304), .A2(n1104), .A3(n1305), .A4(n1085), .ZN(n1303) );
NOR2_X1 U932 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
INV_X1 U933 ( .A(n1102), .ZN(n1307) );
XOR2_X1 U934 ( .A(n1105), .B(KEYINPUT55), .Z(n1304) );
XNOR2_X1 U935 ( .A(G131), .B(n1281), .ZN(G33) );
NAND2_X1 U936 ( .A1(n1104), .A2(n1302), .ZN(n1281) );
AND3_X1 U937 ( .A1(n1085), .A2(n1285), .A3(n1103), .ZN(n1302) );
NOR2_X1 U938 ( .A1(n1149), .A2(n1129), .ZN(n1085) );
INV_X1 U939 ( .A(n1308), .ZN(n1129) );
NAND3_X1 U940 ( .A1(n1309), .A2(n1310), .A3(n1311), .ZN(G30) );
NAND2_X1 U941 ( .A1(n1280), .A2(n1312), .ZN(n1311) );
OR3_X1 U942 ( .A1(n1312), .A2(n1280), .A3(G128), .ZN(n1310) );
INV_X1 U943 ( .A(KEYINPUT2), .ZN(n1312) );
NAND2_X1 U944 ( .A1(G128), .A2(n1313), .ZN(n1309) );
NAND2_X1 U945 ( .A1(KEYINPUT2), .A2(n1314), .ZN(n1313) );
XNOR2_X1 U946 ( .A(KEYINPUT33), .B(n1280), .ZN(n1314) );
NAND3_X1 U947 ( .A1(n1102), .A2(n1272), .A3(n1284), .ZN(n1280) );
AND3_X1 U948 ( .A1(n1315), .A2(n1316), .A3(n1285), .ZN(n1284) );
NOR2_X1 U949 ( .A1(n1105), .A2(n1306), .ZN(n1285) );
XNOR2_X1 U950 ( .A(G101), .B(n1254), .ZN(G3) );
NAND3_X1 U951 ( .A1(n1104), .A2(n1264), .A3(n1107), .ZN(n1254) );
XNOR2_X1 U952 ( .A(G125), .B(n1173), .ZN(G27) );
NAND4_X1 U953 ( .A1(n1121), .A2(n1130), .A3(n1317), .A4(n1103), .ZN(n1173) );
NOR2_X1 U954 ( .A1(n1306), .A2(n1126), .ZN(n1317) );
AND2_X1 U955 ( .A1(n1093), .A2(n1318), .ZN(n1306) );
NAND4_X1 U956 ( .A1(G902), .A2(G953), .A3(n1319), .A4(n1156), .ZN(n1318) );
INV_X1 U957 ( .A(G900), .ZN(n1156) );
XOR2_X1 U958 ( .A(G122), .B(n1320), .Z(G24) );
NOR3_X1 U959 ( .A1(n1268), .A2(n1321), .A3(n1322), .ZN(n1320) );
XNOR2_X1 U960 ( .A(n1121), .B(KEYINPUT53), .ZN(n1322) );
NAND4_X1 U961 ( .A1(n1296), .A2(n1106), .A3(n1272), .A4(n1323), .ZN(n1268) );
INV_X1 U962 ( .A(n1126), .ZN(n1272) );
NOR2_X1 U963 ( .A1(n1316), .A2(n1315), .ZN(n1106) );
XNOR2_X1 U964 ( .A(G119), .B(n1265), .ZN(G21) );
NAND4_X1 U965 ( .A1(n1324), .A2(n1107), .A3(n1315), .A4(n1316), .ZN(n1265) );
XOR2_X1 U966 ( .A(G116), .B(n1325), .Z(G18) );
NOR2_X1 U967 ( .A1(n1126), .A2(n1275), .ZN(n1325) );
NAND4_X1 U968 ( .A1(n1121), .A2(n1104), .A3(n1102), .A4(n1267), .ZN(n1275) );
NOR2_X1 U969 ( .A1(n1296), .A2(n1298), .ZN(n1102) );
INV_X1 U970 ( .A(n1323), .ZN(n1298) );
INV_X1 U971 ( .A(n1092), .ZN(n1121) );
XNOR2_X1 U972 ( .A(G113), .B(n1263), .ZN(G15) );
NAND3_X1 U973 ( .A1(n1104), .A2(n1103), .A3(n1324), .ZN(n1263) );
NOR3_X1 U974 ( .A1(n1126), .A2(n1321), .A3(n1092), .ZN(n1324) );
NAND2_X1 U975 ( .A1(n1326), .A2(n1119), .ZN(n1092) );
INV_X1 U976 ( .A(n1136), .ZN(n1119) );
NOR2_X1 U977 ( .A1(n1323), .A2(n1327), .ZN(n1103) );
NOR2_X1 U978 ( .A1(n1271), .A2(n1316), .ZN(n1104) );
NAND2_X1 U979 ( .A1(n1328), .A2(n1329), .ZN(G12) );
NAND2_X1 U980 ( .A1(n1261), .A2(n1240), .ZN(n1329) );
XOR2_X1 U981 ( .A(KEYINPUT3), .B(n1330), .Z(n1328) );
NOR2_X1 U982 ( .A1(n1261), .A2(n1240), .ZN(n1330) );
AND3_X1 U983 ( .A1(n1107), .A2(n1264), .A3(n1130), .ZN(n1261) );
NOR2_X1 U984 ( .A1(n1315), .A2(n1273), .ZN(n1130) );
INV_X1 U985 ( .A(n1316), .ZN(n1273) );
XOR2_X1 U986 ( .A(n1331), .B(n1144), .Z(n1316) );
NAND2_X1 U987 ( .A1(G217), .A2(n1332), .ZN(n1144) );
XNOR2_X1 U988 ( .A(n1145), .B(KEYINPUT4), .ZN(n1331) );
NOR2_X1 U989 ( .A1(n1193), .A2(G902), .ZN(n1145) );
XNOR2_X1 U990 ( .A(n1333), .B(n1334), .ZN(n1193) );
XOR2_X1 U991 ( .A(n1335), .B(n1336), .Z(n1334) );
XOR2_X1 U992 ( .A(n1337), .B(n1338), .Z(n1336) );
NOR2_X1 U993 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
NOR2_X1 U994 ( .A1(n1341), .A2(n1164), .ZN(n1340) );
NOR2_X1 U995 ( .A1(KEYINPUT54), .A2(G125), .ZN(n1341) );
NOR2_X1 U996 ( .A1(KEYINPUT54), .A2(n1342), .ZN(n1339) );
INV_X1 U997 ( .A(n1167), .ZN(n1342) );
NAND2_X1 U998 ( .A1(KEYINPUT34), .A2(n1343), .ZN(n1337) );
XOR2_X1 U999 ( .A(n1344), .B(n1345), .Z(n1343) );
XNOR2_X1 U1000 ( .A(G110), .B(n1346), .ZN(n1345) );
NOR2_X1 U1001 ( .A1(G128), .A2(KEYINPUT22), .ZN(n1346) );
XNOR2_X1 U1002 ( .A(G119), .B(KEYINPUT44), .ZN(n1344) );
NAND2_X1 U1003 ( .A1(n1347), .A2(n1348), .ZN(n1335) );
NAND2_X1 U1004 ( .A1(KEYINPUT25), .A2(n1349), .ZN(n1348) );
NAND2_X1 U1005 ( .A1(KEYINPUT46), .A2(n1350), .ZN(n1347) );
INV_X1 U1006 ( .A(n1349), .ZN(n1350) );
NAND2_X1 U1007 ( .A1(n1351), .A2(G221), .ZN(n1349) );
XNOR2_X1 U1008 ( .A(G137), .B(n1352), .ZN(n1333) );
XOR2_X1 U1009 ( .A(KEYINPUT18), .B(G146), .Z(n1352) );
INV_X1 U1010 ( .A(n1271), .ZN(n1315) );
XNOR2_X1 U1011 ( .A(n1142), .B(n1353), .ZN(n1271) );
NOR2_X1 U1012 ( .A1(G472), .A2(KEYINPUT50), .ZN(n1353) );
NAND2_X1 U1013 ( .A1(n1354), .A2(n1355), .ZN(n1142) );
XOR2_X1 U1014 ( .A(n1222), .B(n1221), .Z(n1354) );
XOR2_X1 U1015 ( .A(n1356), .B(n1357), .Z(n1221) );
AND2_X1 U1016 ( .A1(G210), .A2(n1358), .ZN(n1357) );
NAND3_X1 U1017 ( .A1(n1359), .A2(n1360), .A3(n1361), .ZN(n1222) );
NAND2_X1 U1018 ( .A1(KEYINPUT38), .A2(n1362), .ZN(n1361) );
NAND3_X1 U1019 ( .A1(n1363), .A2(n1364), .A3(n1365), .ZN(n1360) );
INV_X1 U1020 ( .A(KEYINPUT38), .ZN(n1364) );
OR2_X1 U1021 ( .A1(n1365), .A2(n1363), .ZN(n1359) );
NOR2_X1 U1022 ( .A1(KEYINPUT24), .A2(n1362), .ZN(n1363) );
NOR3_X1 U1023 ( .A1(n1126), .A2(n1321), .A3(n1105), .ZN(n1264) );
NAND2_X1 U1024 ( .A1(n1326), .A2(n1136), .ZN(n1105) );
XOR2_X1 U1025 ( .A(n1366), .B(n1228), .Z(n1136) );
INV_X1 U1026 ( .A(G469), .ZN(n1228) );
NAND2_X1 U1027 ( .A1(n1367), .A2(n1355), .ZN(n1366) );
XOR2_X1 U1028 ( .A(n1368), .B(n1369), .Z(n1367) );
XNOR2_X1 U1029 ( .A(n1356), .B(n1245), .ZN(n1369) );
XNOR2_X1 U1030 ( .A(n1370), .B(n1371), .ZN(n1245) );
XNOR2_X1 U1031 ( .A(G107), .B(KEYINPUT51), .ZN(n1370) );
XNOR2_X1 U1032 ( .A(n1244), .B(n1372), .ZN(n1356) );
INV_X1 U1033 ( .A(n1241), .ZN(n1372) );
XNOR2_X1 U1034 ( .A(n1373), .B(n1374), .ZN(n1241) );
XNOR2_X1 U1035 ( .A(n1169), .B(G131), .ZN(n1374) );
INV_X1 U1036 ( .A(G137), .ZN(n1169) );
NAND2_X1 U1037 ( .A1(KEYINPUT16), .A2(n1375), .ZN(n1373) );
INV_X1 U1038 ( .A(G134), .ZN(n1375) );
XOR2_X1 U1039 ( .A(n1159), .B(G101), .Z(n1244) );
XOR2_X1 U1040 ( .A(n1235), .B(n1376), .Z(n1368) );
XNOR2_X1 U1041 ( .A(n1377), .B(n1240), .ZN(n1376) );
NAND2_X1 U1042 ( .A1(KEYINPUT35), .A2(n1164), .ZN(n1377) );
INV_X1 U1043 ( .A(G140), .ZN(n1164) );
NAND2_X1 U1044 ( .A1(G227), .A2(n1109), .ZN(n1235) );
XNOR2_X1 U1045 ( .A(KEYINPUT56), .B(n1120), .ZN(n1326) );
AND2_X1 U1046 ( .A1(G221), .A2(n1332), .ZN(n1120) );
NAND2_X1 U1047 ( .A1(G234), .A2(n1355), .ZN(n1332) );
INV_X1 U1048 ( .A(n1267), .ZN(n1321) );
NAND2_X1 U1049 ( .A1(n1093), .A2(n1378), .ZN(n1267) );
NAND3_X1 U1050 ( .A1(n1182), .A2(n1319), .A3(G902), .ZN(n1378) );
NOR2_X1 U1051 ( .A1(n1109), .A2(G898), .ZN(n1182) );
NAND3_X1 U1052 ( .A1(n1319), .A2(n1109), .A3(G952), .ZN(n1093) );
NAND2_X1 U1053 ( .A1(G237), .A2(G234), .ZN(n1319) );
NAND2_X1 U1054 ( .A1(n1379), .A2(n1149), .ZN(n1126) );
XOR2_X1 U1055 ( .A(n1380), .B(n1249), .Z(n1149) );
NAND2_X1 U1056 ( .A1(G210), .A2(n1381), .ZN(n1249) );
NAND2_X1 U1057 ( .A1(n1382), .A2(n1355), .ZN(n1380) );
XNOR2_X1 U1058 ( .A(n1184), .B(n1383), .ZN(n1382) );
XOR2_X1 U1059 ( .A(n1384), .B(n1289), .Z(n1383) );
NOR2_X1 U1060 ( .A1(KEYINPUT13), .A2(n1185), .ZN(n1289) );
XNOR2_X1 U1061 ( .A(G122), .B(n1240), .ZN(n1185) );
INV_X1 U1062 ( .A(G110), .ZN(n1240) );
NAND2_X1 U1063 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
OR2_X1 U1064 ( .A1(n1387), .A2(n1293), .ZN(n1386) );
XOR2_X1 U1065 ( .A(n1388), .B(KEYINPUT36), .Z(n1385) );
NAND2_X1 U1066 ( .A1(n1293), .A2(n1387), .ZN(n1388) );
XNOR2_X1 U1067 ( .A(n1159), .B(n1389), .ZN(n1387) );
XNOR2_X1 U1068 ( .A(KEYINPUT15), .B(n1166), .ZN(n1389) );
XNOR2_X1 U1069 ( .A(G146), .B(n1390), .ZN(n1159) );
AND2_X1 U1070 ( .A1(G224), .A2(n1109), .ZN(n1293) );
XNOR2_X1 U1071 ( .A(n1291), .B(G101), .ZN(n1184) );
XOR2_X1 U1072 ( .A(n1391), .B(n1392), .Z(n1291) );
XNOR2_X1 U1073 ( .A(KEYINPUT28), .B(n1365), .ZN(n1392) );
INV_X1 U1074 ( .A(G113), .ZN(n1365) );
XNOR2_X1 U1075 ( .A(n1393), .B(n1362), .ZN(n1391) );
XNOR2_X1 U1076 ( .A(G116), .B(G119), .ZN(n1362) );
NAND3_X1 U1077 ( .A1(n1394), .A2(n1395), .A3(n1396), .ZN(n1393) );
OR2_X1 U1078 ( .A1(n1371), .A2(KEYINPUT10), .ZN(n1396) );
NAND3_X1 U1079 ( .A1(KEYINPUT10), .A2(n1397), .A3(G107), .ZN(n1395) );
INV_X1 U1080 ( .A(n1398), .ZN(n1397) );
NAND2_X1 U1081 ( .A1(n1398), .A2(n1076), .ZN(n1394) );
NAND2_X1 U1082 ( .A1(KEYINPUT37), .A2(n1371), .ZN(n1398) );
XOR2_X1 U1083 ( .A(G104), .B(KEYINPUT47), .Z(n1371) );
XNOR2_X1 U1084 ( .A(KEYINPUT7), .B(n1308), .ZN(n1379) );
NAND2_X1 U1085 ( .A1(G214), .A2(n1381), .ZN(n1308) );
NAND2_X1 U1086 ( .A1(n1399), .A2(n1355), .ZN(n1381) );
INV_X1 U1087 ( .A(G902), .ZN(n1355) );
INV_X1 U1088 ( .A(G237), .ZN(n1399) );
NOR2_X1 U1089 ( .A1(n1323), .A2(n1296), .ZN(n1107) );
INV_X1 U1090 ( .A(n1327), .ZN(n1296) );
XOR2_X1 U1091 ( .A(n1400), .B(n1401), .Z(n1327) );
INV_X1 U1092 ( .A(n1147), .ZN(n1401) );
NOR2_X1 U1093 ( .A1(n1212), .A2(G902), .ZN(n1147) );
INV_X1 U1094 ( .A(n1207), .ZN(n1212) );
XNOR2_X1 U1095 ( .A(n1402), .B(n1403), .ZN(n1207) );
XOR2_X1 U1096 ( .A(n1404), .B(n1405), .Z(n1403) );
XOR2_X1 U1097 ( .A(n1406), .B(n1407), .Z(n1405) );
NAND2_X1 U1098 ( .A1(n1408), .A2(KEYINPUT6), .ZN(n1407) );
XOR2_X1 U1099 ( .A(n1409), .B(n1410), .Z(n1408) );
XOR2_X1 U1100 ( .A(G143), .B(G131), .Z(n1410) );
NAND2_X1 U1101 ( .A1(n1358), .A2(G214), .ZN(n1409) );
NOR2_X1 U1102 ( .A1(G953), .A2(G237), .ZN(n1358) );
NAND2_X1 U1103 ( .A1(n1411), .A2(n1412), .ZN(n1406) );
NAND2_X1 U1104 ( .A1(G140), .A2(n1413), .ZN(n1412) );
NAND2_X1 U1105 ( .A1(n1414), .A2(n1166), .ZN(n1413) );
INV_X1 U1106 ( .A(G125), .ZN(n1166) );
NAND2_X1 U1107 ( .A1(n1167), .A2(n1414), .ZN(n1411) );
INV_X1 U1108 ( .A(KEYINPUT32), .ZN(n1414) );
NOR2_X1 U1109 ( .A1(G125), .A2(G140), .ZN(n1167) );
NOR2_X1 U1110 ( .A1(G113), .A2(KEYINPUT0), .ZN(n1404) );
XNOR2_X1 U1111 ( .A(G104), .B(n1415), .ZN(n1402) );
XOR2_X1 U1112 ( .A(G146), .B(G122), .Z(n1415) );
NAND2_X1 U1113 ( .A1(KEYINPUT59), .A2(n1213), .ZN(n1400) );
INV_X1 U1114 ( .A(G475), .ZN(n1213) );
NAND3_X1 U1115 ( .A1(n1416), .A2(n1417), .A3(n1418), .ZN(n1323) );
NAND2_X1 U1116 ( .A1(KEYINPUT12), .A2(n1419), .ZN(n1418) );
NAND3_X1 U1117 ( .A1(n1420), .A2(n1421), .A3(G478), .ZN(n1417) );
NAND2_X1 U1118 ( .A1(n1422), .A2(n1140), .ZN(n1416) );
INV_X1 U1119 ( .A(G478), .ZN(n1140) );
NAND2_X1 U1120 ( .A1(n1423), .A2(n1421), .ZN(n1422) );
INV_X1 U1121 ( .A(KEYINPUT12), .ZN(n1421) );
XNOR2_X1 U1122 ( .A(KEYINPUT60), .B(n1419), .ZN(n1423) );
INV_X1 U1123 ( .A(n1420), .ZN(n1419) );
XOR2_X1 U1124 ( .A(n1141), .B(KEYINPUT31), .Z(n1420) );
NOR2_X1 U1125 ( .A1(n1201), .A2(G902), .ZN(n1141) );
XNOR2_X1 U1126 ( .A(n1424), .B(n1425), .ZN(n1201) );
AND2_X1 U1127 ( .A1(n1351), .A2(G217), .ZN(n1425) );
AND2_X1 U1128 ( .A1(G234), .A2(n1109), .ZN(n1351) );
INV_X1 U1129 ( .A(G953), .ZN(n1109) );
NAND3_X1 U1130 ( .A1(n1426), .A2(n1427), .A3(KEYINPUT29), .ZN(n1424) );
NAND2_X1 U1131 ( .A1(n1428), .A2(n1429), .ZN(n1427) );
NAND2_X1 U1132 ( .A1(n1430), .A2(n1431), .ZN(n1428) );
NAND2_X1 U1133 ( .A1(KEYINPUT5), .A2(n1432), .ZN(n1431) );
NAND2_X1 U1134 ( .A1(n1433), .A2(n1434), .ZN(n1430) );
INV_X1 U1135 ( .A(KEYINPUT5), .ZN(n1434) );
OR2_X1 U1136 ( .A1(n1429), .A2(n1432), .ZN(n1426) );
NAND2_X1 U1137 ( .A1(KEYINPUT26), .A2(n1433), .ZN(n1432) );
XNOR2_X1 U1138 ( .A(G134), .B(n1390), .ZN(n1433) );
XOR2_X1 U1139 ( .A(G143), .B(G128), .Z(n1390) );
XOR2_X1 U1140 ( .A(n1076), .B(n1435), .Z(n1429) );
XOR2_X1 U1141 ( .A(G122), .B(G116), .Z(n1435) );
INV_X1 U1142 ( .A(G107), .ZN(n1076) );
endmodule


