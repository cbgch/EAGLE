//Key = 1000011100111010110101101101000010111111010000110011110001011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;

XOR2_X1 U732 ( .A(n1019), .B(n1020), .Z(G9) );
NAND2_X1 U733 ( .A1(KEYINPUT61), .A2(G107), .ZN(n1020) );
NOR2_X1 U734 ( .A1(n1021), .A2(n1022), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1022) );
XOR2_X1 U736 ( .A(n1027), .B(KEYINPUT54), .Z(n1025) );
NAND3_X1 U737 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1023) );
NAND2_X1 U738 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U739 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND4_X1 U740 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1034) );
NAND3_X1 U741 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NAND2_X1 U742 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U743 ( .A1(n1044), .A2(n1045), .ZN(n1039) );
NAND2_X1 U744 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U745 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND3_X1 U746 ( .A1(n1044), .A2(n1050), .A3(n1042), .ZN(n1033) );
NAND2_X1 U747 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U748 ( .A1(n1035), .A2(n1053), .ZN(n1052) );
NAND2_X1 U749 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U750 ( .A1(n1037), .A2(n1056), .ZN(n1055) );
OR2_X1 U751 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U752 ( .A1(n1036), .A2(n1059), .ZN(n1054) );
NAND2_X1 U753 ( .A1(n1036), .A2(n1060), .ZN(n1051) );
INV_X1 U754 ( .A(n1061), .ZN(n1031) );
NOR3_X1 U755 ( .A1(n1062), .A2(G953), .A3(G952), .ZN(n1021) );
INV_X1 U756 ( .A(n1028), .ZN(n1062) );
NAND4_X1 U757 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1028) );
NOR4_X1 U758 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
XOR2_X1 U759 ( .A(n1071), .B(n1072), .Z(n1070) );
XNOR2_X1 U760 ( .A(KEYINPUT42), .B(n1035), .ZN(n1069) );
NOR2_X1 U761 ( .A1(n1059), .A2(n1048), .ZN(n1065) );
XNOR2_X1 U762 ( .A(n1073), .B(n1074), .ZN(n1064) );
XNOR2_X1 U763 ( .A(n1075), .B(KEYINPUT10), .ZN(n1074) );
INV_X1 U764 ( .A(n1076), .ZN(n1075) );
XOR2_X1 U765 ( .A(KEYINPUT20), .B(n1077), .Z(n1063) );
XOR2_X1 U766 ( .A(n1078), .B(n1079), .Z(G72) );
XOR2_X1 U767 ( .A(n1080), .B(n1081), .Z(n1079) );
NAND2_X1 U768 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U769 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
INV_X1 U770 ( .A(n1026), .ZN(n1085) );
XOR2_X1 U771 ( .A(n1024), .B(KEYINPUT37), .Z(n1084) );
XNOR2_X1 U772 ( .A(KEYINPUT22), .B(n1029), .ZN(n1082) );
NAND3_X1 U773 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1080) );
NAND2_X1 U774 ( .A1(G953), .A2(n1089), .ZN(n1088) );
NAND2_X1 U775 ( .A1(n1090), .A2(n1091), .ZN(n1087) );
NAND2_X1 U776 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NAND2_X1 U777 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
INV_X1 U778 ( .A(n1096), .ZN(n1095) );
NAND2_X1 U779 ( .A1(n1096), .A2(n1097), .ZN(n1092) );
XNOR2_X1 U780 ( .A(n1098), .B(KEYINPUT7), .ZN(n1096) );
NAND2_X1 U781 ( .A1(G140), .A2(n1099), .ZN(n1086) );
NAND2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U783 ( .A1(n1102), .A2(n1094), .ZN(n1101) );
NAND2_X1 U784 ( .A1(n1097), .A2(n1103), .ZN(n1100) );
INV_X1 U785 ( .A(n1102), .ZN(n1103) );
XNOR2_X1 U786 ( .A(n1098), .B(KEYINPUT51), .ZN(n1102) );
XNOR2_X1 U787 ( .A(n1104), .B(KEYINPUT18), .ZN(n1098) );
XNOR2_X1 U788 ( .A(n1094), .B(KEYINPUT30), .ZN(n1097) );
XOR2_X1 U789 ( .A(n1105), .B(n1106), .Z(n1094) );
XNOR2_X1 U790 ( .A(n1107), .B(KEYINPUT58), .ZN(n1106) );
NAND2_X1 U791 ( .A1(KEYINPUT60), .A2(n1108), .ZN(n1107) );
NOR2_X1 U792 ( .A1(n1109), .A2(n1029), .ZN(n1078) );
AND2_X1 U793 ( .A1(G227), .A2(G900), .ZN(n1109) );
XOR2_X1 U794 ( .A(n1110), .B(n1111), .Z(G69) );
NOR2_X1 U795 ( .A1(n1112), .A2(n1029), .ZN(n1111) );
NOR2_X1 U796 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND2_X1 U797 ( .A1(n1115), .A2(n1116), .ZN(n1110) );
NAND3_X1 U798 ( .A1(n1117), .A2(n1027), .A3(n1118), .ZN(n1116) );
NAND2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1115) );
NAND2_X1 U800 ( .A1(n1118), .A2(n1027), .ZN(n1120) );
XNOR2_X1 U801 ( .A(n1029), .B(KEYINPUT0), .ZN(n1118) );
XNOR2_X1 U802 ( .A(KEYINPUT8), .B(n1117), .ZN(n1119) );
NAND2_X1 U803 ( .A1(n1121), .A2(n1122), .ZN(n1117) );
NAND2_X1 U804 ( .A1(G953), .A2(n1114), .ZN(n1122) );
NOR2_X1 U805 ( .A1(n1123), .A2(n1124), .ZN(G66) );
XOR2_X1 U806 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND2_X1 U807 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
XNOR2_X1 U808 ( .A(KEYINPUT29), .B(n1076), .ZN(n1128) );
NOR2_X1 U809 ( .A1(n1123), .A2(n1129), .ZN(G63) );
XOR2_X1 U810 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U811 ( .A1(n1127), .A2(G478), .ZN(n1130) );
NOR2_X1 U812 ( .A1(n1123), .A2(n1132), .ZN(G60) );
XOR2_X1 U813 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U814 ( .A1(n1127), .A2(G475), .ZN(n1133) );
XOR2_X1 U815 ( .A(G104), .B(n1135), .Z(G6) );
NOR2_X1 U816 ( .A1(n1046), .A2(n1136), .ZN(n1135) );
NOR2_X1 U817 ( .A1(n1123), .A2(n1137), .ZN(G57) );
XOR2_X1 U818 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U819 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U820 ( .A(n1142), .B(n1143), .ZN(n1141) );
NAND2_X1 U821 ( .A1(n1127), .A2(G472), .ZN(n1142) );
XOR2_X1 U822 ( .A(n1144), .B(n1145), .Z(n1138) );
XOR2_X1 U823 ( .A(n1146), .B(KEYINPUT4), .Z(n1145) );
NAND2_X1 U824 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U825 ( .A1(KEYINPUT62), .A2(n1149), .ZN(n1144) );
NOR2_X1 U826 ( .A1(n1123), .A2(n1150), .ZN(G54) );
XOR2_X1 U827 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U828 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U829 ( .A1(n1127), .A2(G469), .ZN(n1153) );
NOR2_X1 U830 ( .A1(n1155), .A2(n1156), .ZN(n1151) );
NOR2_X1 U831 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XOR2_X1 U832 ( .A(KEYINPUT25), .B(n1159), .Z(n1158) );
NOR2_X1 U833 ( .A1(n1160), .A2(n1159), .ZN(n1155) );
XNOR2_X1 U834 ( .A(n1091), .B(n1161), .ZN(n1159) );
NOR2_X1 U835 ( .A1(G110), .A2(KEYINPUT15), .ZN(n1161) );
INV_X1 U836 ( .A(n1157), .ZN(n1160) );
NOR2_X1 U837 ( .A1(n1029), .A2(G952), .ZN(n1123) );
NOR2_X1 U838 ( .A1(n1162), .A2(n1163), .ZN(G51) );
XOR2_X1 U839 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U840 ( .A1(n1127), .A2(n1072), .ZN(n1164) );
AND2_X1 U841 ( .A1(G902), .A2(n1166), .ZN(n1127) );
OR3_X1 U842 ( .A1(n1026), .A2(n1027), .A3(n1024), .ZN(n1166) );
NAND4_X1 U843 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1024) );
NAND3_X1 U844 ( .A1(n1171), .A2(n1057), .A3(n1172), .ZN(n1168) );
NAND2_X1 U845 ( .A1(n1173), .A2(n1174), .ZN(n1167) );
XOR2_X1 U846 ( .A(KEYINPUT3), .B(n1175), .Z(n1174) );
NAND3_X1 U847 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1027) );
AND3_X1 U848 ( .A1(n1179), .A2(n1019), .A3(n1180), .ZN(n1178) );
NAND4_X1 U849 ( .A1(n1173), .A2(n1058), .A3(n1044), .A4(n1181), .ZN(n1019) );
NAND2_X1 U850 ( .A1(n1173), .A2(n1182), .ZN(n1176) );
NAND4_X1 U851 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1182) );
NAND3_X1 U852 ( .A1(n1187), .A2(n1044), .A3(n1188), .ZN(n1186) );
XNOR2_X1 U853 ( .A(n1189), .B(KEYINPUT57), .ZN(n1188) );
NAND3_X1 U854 ( .A1(n1043), .A2(n1181), .A3(n1036), .ZN(n1185) );
XNOR2_X1 U855 ( .A(KEYINPUT47), .B(n1136), .ZN(n1184) );
NAND3_X1 U856 ( .A1(n1044), .A2(n1181), .A3(n1057), .ZN(n1136) );
XNOR2_X1 U857 ( .A(KEYINPUT14), .B(n1190), .ZN(n1183) );
NAND4_X1 U858 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1026) );
NAND3_X1 U859 ( .A1(n1195), .A2(n1042), .A3(n1036), .ZN(n1191) );
NOR2_X1 U860 ( .A1(G952), .A2(n1196), .ZN(n1162) );
XNOR2_X1 U861 ( .A(G953), .B(KEYINPUT56), .ZN(n1196) );
XOR2_X1 U862 ( .A(n1192), .B(n1197), .Z(G48) );
NAND2_X1 U863 ( .A1(KEYINPUT41), .A2(G146), .ZN(n1197) );
NAND3_X1 U864 ( .A1(n1057), .A2(n1173), .A3(n1195), .ZN(n1192) );
XNOR2_X1 U865 ( .A(G143), .B(n1193), .ZN(G45) );
NAND3_X1 U866 ( .A1(n1189), .A2(n1172), .A3(n1198), .ZN(n1193) );
XNOR2_X1 U867 ( .A(G140), .B(n1199), .ZN(G42) );
NOR2_X1 U868 ( .A1(n1200), .A2(KEYINPUT63), .ZN(n1199) );
INV_X1 U869 ( .A(n1194), .ZN(n1200) );
NAND4_X1 U870 ( .A1(n1172), .A2(n1042), .A3(n1057), .A4(n1043), .ZN(n1194) );
XOR2_X1 U871 ( .A(G137), .B(n1201), .Z(G39) );
NOR3_X1 U872 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1201) );
XOR2_X1 U873 ( .A(KEYINPUT52), .B(n1042), .Z(n1202) );
XNOR2_X1 U874 ( .A(G134), .B(n1169), .ZN(G36) );
NAND3_X1 U875 ( .A1(n1171), .A2(n1058), .A3(n1172), .ZN(n1169) );
XNOR2_X1 U876 ( .A(G131), .B(n1205), .ZN(G33) );
NAND4_X1 U877 ( .A1(n1206), .A2(n1171), .A3(n1057), .A4(n1207), .ZN(n1205) );
INV_X1 U878 ( .A(n1040), .ZN(n1171) );
NAND3_X1 U879 ( .A1(n1208), .A2(n1067), .A3(n1042), .ZN(n1040) );
NOR2_X1 U880 ( .A1(n1209), .A2(n1048), .ZN(n1042) );
XNOR2_X1 U881 ( .A(n1060), .B(KEYINPUT16), .ZN(n1206) );
NAND2_X1 U882 ( .A1(n1210), .A2(n1211), .ZN(G30) );
NAND4_X1 U883 ( .A1(n1175), .A2(n1173), .A3(n1212), .A4(n1213), .ZN(n1211) );
NAND2_X1 U884 ( .A1(G128), .A2(n1214), .ZN(n1213) );
OR2_X1 U885 ( .A1(G128), .A2(KEYINPUT5), .ZN(n1212) );
NAND3_X1 U886 ( .A1(n1215), .A2(n1214), .A3(G128), .ZN(n1210) );
INV_X1 U887 ( .A(KEYINPUT13), .ZN(n1214) );
NAND3_X1 U888 ( .A1(n1175), .A2(n1173), .A3(KEYINPUT5), .ZN(n1215) );
AND2_X1 U889 ( .A1(n1195), .A2(n1058), .ZN(n1175) );
INV_X1 U890 ( .A(n1203), .ZN(n1195) );
NAND3_X1 U891 ( .A1(n1172), .A2(n1067), .A3(n1216), .ZN(n1203) );
AND2_X1 U892 ( .A1(n1060), .A2(n1207), .ZN(n1172) );
XNOR2_X1 U893 ( .A(G101), .B(n1177), .ZN(G3) );
NAND3_X1 U894 ( .A1(n1198), .A2(n1181), .A3(n1036), .ZN(n1177) );
XNOR2_X1 U895 ( .A(G125), .B(n1170), .ZN(G27) );
NAND4_X1 U896 ( .A1(n1035), .A2(n1043), .A3(n1057), .A4(n1217), .ZN(n1170) );
AND3_X1 U897 ( .A1(n1173), .A2(n1207), .A3(n1037), .ZN(n1217) );
NAND2_X1 U898 ( .A1(n1061), .A2(n1218), .ZN(n1207) );
NAND4_X1 U899 ( .A1(G953), .A2(G902), .A3(n1219), .A4(n1089), .ZN(n1218) );
INV_X1 U900 ( .A(G900), .ZN(n1089) );
XNOR2_X1 U901 ( .A(G122), .B(n1220), .ZN(G24) );
NAND3_X1 U902 ( .A1(n1221), .A2(n1187), .A3(n1222), .ZN(n1220) );
AND3_X1 U903 ( .A1(n1189), .A2(n1223), .A3(n1044), .ZN(n1222) );
NOR2_X1 U904 ( .A1(n1067), .A2(n1224), .ZN(n1044) );
INV_X1 U905 ( .A(KEYINPUT31), .ZN(n1223) );
NOR2_X1 U906 ( .A1(n1077), .A2(n1225), .ZN(n1189) );
XNOR2_X1 U907 ( .A(n1173), .B(KEYINPUT21), .ZN(n1221) );
XOR2_X1 U908 ( .A(G119), .B(n1226), .Z(G21) );
NOR2_X1 U909 ( .A1(n1046), .A2(n1190), .ZN(n1226) );
NAND4_X1 U910 ( .A1(n1187), .A2(n1036), .A3(n1216), .A4(n1067), .ZN(n1190) );
XNOR2_X1 U911 ( .A(n1224), .B(KEYINPUT32), .ZN(n1216) );
INV_X1 U912 ( .A(n1173), .ZN(n1046) );
XNOR2_X1 U913 ( .A(G116), .B(n1179), .ZN(G18) );
NAND3_X1 U914 ( .A1(n1198), .A2(n1058), .A3(n1187), .ZN(n1179) );
AND2_X1 U915 ( .A1(n1077), .A2(n1068), .ZN(n1058) );
XNOR2_X1 U916 ( .A(G113), .B(n1180), .ZN(G15) );
NAND3_X1 U917 ( .A1(n1198), .A2(n1057), .A3(n1187), .ZN(n1180) );
AND3_X1 U918 ( .A1(n1037), .A2(n1227), .A3(n1035), .ZN(n1187) );
NOR2_X1 U919 ( .A1(n1068), .A2(n1077), .ZN(n1057) );
AND3_X1 U920 ( .A1(n1208), .A2(n1067), .A3(n1173), .ZN(n1198) );
XOR2_X1 U921 ( .A(n1228), .B(n1229), .Z(G12) );
NOR2_X1 U922 ( .A1(G110), .A2(KEYINPUT43), .ZN(n1229) );
NAND4_X1 U923 ( .A1(n1230), .A2(n1036), .A3(n1043), .A4(n1181), .ZN(n1228) );
AND2_X1 U924 ( .A1(n1060), .A2(n1227), .ZN(n1181) );
NAND2_X1 U925 ( .A1(n1061), .A2(n1231), .ZN(n1227) );
NAND4_X1 U926 ( .A1(G953), .A2(G902), .A3(n1219), .A4(n1114), .ZN(n1231) );
INV_X1 U927 ( .A(G898), .ZN(n1114) );
NAND3_X1 U928 ( .A1(n1219), .A2(n1029), .A3(G952), .ZN(n1061) );
NAND2_X1 U929 ( .A1(G237), .A2(G234), .ZN(n1219) );
NOR2_X1 U930 ( .A1(n1232), .A2(n1035), .ZN(n1060) );
XOR2_X1 U931 ( .A(n1233), .B(G469), .Z(n1035) );
NAND2_X1 U932 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U933 ( .A(n1236), .B(n1237), .Z(n1234) );
XNOR2_X1 U934 ( .A(n1091), .B(n1238), .ZN(n1237) );
NOR2_X1 U935 ( .A1(G110), .A2(KEYINPUT23), .ZN(n1238) );
XOR2_X1 U936 ( .A(n1154), .B(n1239), .Z(n1236) );
NOR2_X1 U937 ( .A1(KEYINPUT9), .A2(n1157), .ZN(n1239) );
NAND2_X1 U938 ( .A1(G227), .A2(n1029), .ZN(n1157) );
XOR2_X1 U939 ( .A(n1240), .B(n1241), .Z(n1154) );
XNOR2_X1 U940 ( .A(n1108), .B(n1105), .ZN(n1240) );
XOR2_X1 U941 ( .A(G128), .B(n1242), .Z(n1108) );
XOR2_X1 U942 ( .A(n1037), .B(KEYINPUT17), .Z(n1232) );
XOR2_X1 U943 ( .A(n1059), .B(KEYINPUT6), .Z(n1037) );
AND2_X1 U944 ( .A1(G221), .A2(n1243), .ZN(n1059) );
NOR2_X1 U945 ( .A1(n1067), .A2(n1208), .ZN(n1043) );
INV_X1 U946 ( .A(n1224), .ZN(n1208) );
XOR2_X1 U947 ( .A(n1244), .B(n1076), .Z(n1224) );
NAND2_X1 U948 ( .A1(G217), .A2(n1243), .ZN(n1076) );
NAND2_X1 U949 ( .A1(G234), .A2(n1235), .ZN(n1243) );
NAND2_X1 U950 ( .A1(KEYINPUT19), .A2(n1073), .ZN(n1244) );
AND2_X1 U951 ( .A1(n1126), .A2(n1235), .ZN(n1073) );
XNOR2_X1 U952 ( .A(n1245), .B(n1246), .ZN(n1126) );
XNOR2_X1 U953 ( .A(n1247), .B(n1248), .ZN(n1246) );
XOR2_X1 U954 ( .A(KEYINPUT24), .B(G137), .Z(n1248) );
XOR2_X1 U955 ( .A(n1249), .B(n1250), .Z(n1245) );
XOR2_X1 U956 ( .A(n1251), .B(n1252), .Z(n1250) );
NAND2_X1 U957 ( .A1(KEYINPUT11), .A2(n1253), .ZN(n1252) );
XOR2_X1 U958 ( .A(G119), .B(n1254), .Z(n1253) );
XOR2_X1 U959 ( .A(KEYINPUT33), .B(G128), .Z(n1254) );
NAND3_X1 U960 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1251) );
NAND2_X1 U961 ( .A1(KEYINPUT55), .A2(n1258), .ZN(n1257) );
NAND3_X1 U962 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1256) );
INV_X1 U963 ( .A(KEYINPUT55), .ZN(n1260) );
OR2_X1 U964 ( .A1(n1261), .A2(n1259), .ZN(n1255) );
NOR2_X1 U965 ( .A1(KEYINPUT49), .A2(n1258), .ZN(n1259) );
NAND2_X1 U966 ( .A1(G221), .A2(n1262), .ZN(n1249) );
XNOR2_X1 U967 ( .A(n1263), .B(G472), .ZN(n1067) );
NAND2_X1 U968 ( .A1(n1264), .A2(n1235), .ZN(n1263) );
XOR2_X1 U969 ( .A(n1265), .B(n1266), .Z(n1264) );
NAND2_X1 U970 ( .A1(KEYINPUT36), .A2(n1267), .ZN(n1266) );
XOR2_X1 U971 ( .A(n1140), .B(n1268), .Z(n1267) );
XNOR2_X1 U972 ( .A(n1149), .B(n1143), .ZN(n1268) );
XNOR2_X1 U973 ( .A(n1269), .B(n1270), .ZN(n1143) );
XOR2_X1 U974 ( .A(KEYINPUT40), .B(G119), .Z(n1270) );
XNOR2_X1 U975 ( .A(G113), .B(G116), .ZN(n1269) );
INV_X1 U976 ( .A(n1105), .ZN(n1149) );
XNOR2_X1 U977 ( .A(n1271), .B(n1272), .ZN(n1105) );
XNOR2_X1 U978 ( .A(G137), .B(G134), .ZN(n1271) );
NAND2_X1 U979 ( .A1(n1273), .A2(n1148), .ZN(n1265) );
NAND2_X1 U980 ( .A1(n1274), .A2(n1275), .ZN(n1148) );
NAND2_X1 U981 ( .A1(n1276), .A2(G210), .ZN(n1275) );
XOR2_X1 U982 ( .A(n1147), .B(KEYINPUT44), .Z(n1273) );
NAND3_X1 U983 ( .A1(n1277), .A2(G210), .A3(n1276), .ZN(n1147) );
INV_X1 U984 ( .A(n1274), .ZN(n1277) );
INV_X1 U985 ( .A(n1204), .ZN(n1036) );
NAND2_X1 U986 ( .A1(n1225), .A2(n1077), .ZN(n1204) );
XNOR2_X1 U987 ( .A(n1278), .B(n1279), .ZN(n1077) );
XOR2_X1 U988 ( .A(KEYINPUT53), .B(G475), .Z(n1279) );
NAND2_X1 U989 ( .A1(n1134), .A2(n1235), .ZN(n1278) );
XNOR2_X1 U990 ( .A(n1280), .B(n1281), .ZN(n1134) );
XNOR2_X1 U991 ( .A(n1242), .B(n1258), .ZN(n1281) );
XNOR2_X1 U992 ( .A(n1091), .B(n1282), .ZN(n1258) );
INV_X1 U993 ( .A(G140), .ZN(n1091) );
XOR2_X1 U994 ( .A(n1283), .B(n1272), .Z(n1280) );
XOR2_X1 U995 ( .A(G131), .B(KEYINPUT27), .Z(n1272) );
XOR2_X1 U996 ( .A(n1284), .B(n1285), .Z(n1283) );
AND2_X1 U997 ( .A1(G214), .A2(n1276), .ZN(n1285) );
AND2_X1 U998 ( .A1(n1286), .A2(n1029), .ZN(n1276) );
XNOR2_X1 U999 ( .A(G237), .B(KEYINPUT48), .ZN(n1286) );
NAND2_X1 U1000 ( .A1(KEYINPUT35), .A2(n1287), .ZN(n1284) );
XNOR2_X1 U1001 ( .A(G104), .B(n1288), .ZN(n1287) );
NOR2_X1 U1002 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
AND2_X1 U1003 ( .A1(KEYINPUT26), .A2(n1291), .ZN(n1290) );
NOR2_X1 U1004 ( .A1(KEYINPUT2), .A2(n1291), .ZN(n1289) );
INV_X1 U1005 ( .A(n1068), .ZN(n1225) );
XNOR2_X1 U1006 ( .A(n1292), .B(G478), .ZN(n1068) );
NAND2_X1 U1007 ( .A1(n1131), .A2(n1235), .ZN(n1292) );
XOR2_X1 U1008 ( .A(n1293), .B(n1294), .Z(n1131) );
XNOR2_X1 U1009 ( .A(n1295), .B(n1296), .ZN(n1294) );
NAND2_X1 U1010 ( .A1(G217), .A2(n1262), .ZN(n1295) );
AND2_X1 U1011 ( .A1(G234), .A2(n1029), .ZN(n1262) );
INV_X1 U1012 ( .A(G953), .ZN(n1029) );
XOR2_X1 U1013 ( .A(n1297), .B(n1298), .Z(n1293) );
XNOR2_X1 U1014 ( .A(n1299), .B(G107), .ZN(n1298) );
NAND2_X1 U1015 ( .A1(n1300), .A2(n1301), .ZN(n1297) );
NAND2_X1 U1016 ( .A1(G134), .A2(n1302), .ZN(n1301) );
XOR2_X1 U1017 ( .A(KEYINPUT50), .B(n1303), .Z(n1300) );
NOR2_X1 U1018 ( .A1(G134), .A2(n1302), .ZN(n1303) );
XNOR2_X1 U1019 ( .A(n1304), .B(G128), .ZN(n1302) );
INV_X1 U1020 ( .A(G143), .ZN(n1304) );
XNOR2_X1 U1021 ( .A(n1173), .B(KEYINPUT46), .ZN(n1230) );
NOR2_X1 U1022 ( .A1(n1049), .A2(n1048), .ZN(n1173) );
AND2_X1 U1023 ( .A1(G214), .A2(n1305), .ZN(n1048) );
INV_X1 U1024 ( .A(n1209), .ZN(n1049) );
XNOR2_X1 U1025 ( .A(n1306), .B(n1072), .ZN(n1209) );
AND2_X1 U1026 ( .A1(G210), .A2(n1305), .ZN(n1072) );
NAND2_X1 U1027 ( .A1(n1307), .A2(n1235), .ZN(n1305) );
INV_X1 U1028 ( .A(G237), .ZN(n1307) );
NAND2_X1 U1029 ( .A1(KEYINPUT39), .A2(n1071), .ZN(n1306) );
AND2_X1 U1030 ( .A1(n1308), .A2(n1235), .ZN(n1071) );
INV_X1 U1031 ( .A(G902), .ZN(n1235) );
XNOR2_X1 U1032 ( .A(n1165), .B(KEYINPUT38), .ZN(n1308) );
XNOR2_X1 U1033 ( .A(n1309), .B(n1310), .ZN(n1165) );
XNOR2_X1 U1034 ( .A(n1311), .B(n1282), .ZN(n1310) );
INV_X1 U1035 ( .A(n1104), .ZN(n1282) );
XOR2_X1 U1036 ( .A(G125), .B(KEYINPUT45), .Z(n1104) );
NOR2_X1 U1037 ( .A1(G953), .A2(n1113), .ZN(n1311) );
INV_X1 U1038 ( .A(G224), .ZN(n1113) );
XNOR2_X1 U1039 ( .A(n1121), .B(n1140), .ZN(n1309) );
XOR2_X1 U1040 ( .A(n1242), .B(n1312), .Z(n1140) );
NOR2_X1 U1041 ( .A1(G128), .A2(KEYINPUT28), .ZN(n1312) );
XNOR2_X1 U1042 ( .A(G143), .B(n1261), .ZN(n1242) );
INV_X1 U1043 ( .A(G146), .ZN(n1261) );
XNOR2_X1 U1044 ( .A(n1313), .B(n1314), .ZN(n1121) );
XOR2_X1 U1045 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1046 ( .A(G119), .B(n1317), .ZN(n1316) );
NAND2_X1 U1047 ( .A1(KEYINPUT59), .A2(n1247), .ZN(n1317) );
INV_X1 U1048 ( .A(G110), .ZN(n1247) );
NOR2_X1 U1049 ( .A1(KEYINPUT1), .A2(n1299), .ZN(n1315) );
INV_X1 U1050 ( .A(G116), .ZN(n1299) );
XOR2_X1 U1051 ( .A(n1291), .B(n1241), .Z(n1313) );
XNOR2_X1 U1052 ( .A(n1318), .B(n1274), .ZN(n1241) );
XOR2_X1 U1053 ( .A(G101), .B(KEYINPUT12), .Z(n1274) );
XNOR2_X1 U1054 ( .A(G104), .B(G107), .ZN(n1318) );
XNOR2_X1 U1055 ( .A(G113), .B(n1296), .ZN(n1291) );
XOR2_X1 U1056 ( .A(G122), .B(KEYINPUT34), .Z(n1296) );
endmodule


