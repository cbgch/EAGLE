//Key = 0111100000011000111010100110100000100001010110100011110100110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336;

XNOR2_X1 U733 ( .A(G107), .B(n1015), .ZN(G9) );
NOR2_X1 U734 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR3_X1 U735 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1017) );
AND4_X1 U736 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1019) );
INV_X1 U737 ( .A(KEYINPUT32), .ZN(n1018) );
NOR2_X1 U738 ( .A1(KEYINPUT32), .A2(n1025), .ZN(n1016) );
NOR2_X1 U739 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR4_X1 U740 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1027) );
NAND3_X1 U741 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1028) );
NAND4_X1 U742 ( .A1(n1035), .A2(n1022), .A3(n1036), .A4(n1037), .ZN(n1034) );
NAND2_X1 U743 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND3_X1 U744 ( .A1(n1040), .A2(n1041), .A3(KEYINPUT21), .ZN(n1038) );
NAND3_X1 U745 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1036) );
NAND2_X1 U746 ( .A1(n1041), .A2(n1045), .ZN(n1043) );
NAND2_X1 U747 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND3_X1 U748 ( .A1(G214), .A2(n1048), .A3(n1049), .ZN(n1047) );
NAND2_X1 U749 ( .A1(n1040), .A2(n1050), .ZN(n1046) );
INV_X1 U750 ( .A(KEYINPUT21), .ZN(n1050) );
XNOR2_X1 U751 ( .A(n1051), .B(KEYINPUT2), .ZN(n1040) );
NAND2_X1 U752 ( .A1(n1052), .A2(n1053), .ZN(n1042) );
NAND2_X1 U753 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U754 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
INV_X1 U755 ( .A(n1024), .ZN(n1054) );
NAND4_X1 U756 ( .A1(n1044), .A2(n1041), .A3(n1052), .A4(n1058), .ZN(n1032) );
NAND2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U758 ( .A1(n1022), .A2(n1061), .ZN(n1060) );
OR2_X1 U759 ( .A1(n1062), .A2(n1023), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1035), .A2(n1063), .ZN(n1059) );
NAND2_X1 U761 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
XNOR2_X1 U762 ( .A(n1066), .B(KEYINPUT6), .ZN(n1064) );
NOR3_X1 U763 ( .A1(n1067), .A2(n1068), .A3(n1031), .ZN(n1026) );
INV_X1 U764 ( .A(n1033), .ZN(n1068) );
NAND4_X1 U765 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1033) );
NOR4_X1 U766 ( .A1(n1056), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1072) );
XNOR2_X1 U767 ( .A(n1076), .B(n1077), .ZN(n1071) );
XNOR2_X1 U768 ( .A(n1078), .B(G475), .ZN(n1070) );
XNOR2_X1 U769 ( .A(n1079), .B(n1080), .ZN(n1069) );
NAND2_X1 U770 ( .A1(KEYINPUT44), .A2(n1081), .ZN(n1079) );
XNOR2_X1 U771 ( .A(KEYINPUT24), .B(n1030), .ZN(n1067) );
XOR2_X1 U772 ( .A(n1082), .B(n1083), .Z(G72) );
NOR2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
AND2_X1 U774 ( .A1(G227), .A2(G900), .ZN(n1084) );
NAND2_X1 U775 ( .A1(n1086), .A2(n1087), .ZN(n1082) );
NAND3_X1 U776 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1087) );
INV_X1 U777 ( .A(n1091), .ZN(n1089) );
OR2_X1 U778 ( .A1(n1090), .A2(n1088), .ZN(n1086) );
XNOR2_X1 U779 ( .A(n1092), .B(n1093), .ZN(n1088) );
XNOR2_X1 U780 ( .A(n1094), .B(n1095), .ZN(n1093) );
NAND2_X1 U781 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NAND2_X1 U782 ( .A1(G131), .A2(n1098), .ZN(n1097) );
XOR2_X1 U783 ( .A(n1099), .B(KEYINPUT15), .Z(n1096) );
OR2_X1 U784 ( .A1(n1098), .A2(G131), .ZN(n1099) );
XNOR2_X1 U785 ( .A(G140), .B(n1100), .ZN(n1092) );
NOR2_X1 U786 ( .A1(G125), .A2(KEYINPUT29), .ZN(n1100) );
OR2_X1 U787 ( .A1(G953), .A2(n1101), .ZN(n1090) );
XOR2_X1 U788 ( .A(n1102), .B(n1103), .Z(G69) );
XOR2_X1 U789 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U791 ( .A1(G953), .A2(n1108), .ZN(n1107) );
XNOR2_X1 U792 ( .A(n1109), .B(n1110), .ZN(n1106) );
XNOR2_X1 U793 ( .A(n1111), .B(n1112), .ZN(n1109) );
NAND2_X1 U794 ( .A1(n1113), .A2(n1085), .ZN(n1104) );
XOR2_X1 U795 ( .A(n1114), .B(KEYINPUT57), .Z(n1113) );
NAND2_X1 U796 ( .A1(n1115), .A2(n1025), .ZN(n1114) );
NOR2_X1 U797 ( .A1(n1116), .A2(n1085), .ZN(n1102) );
NOR2_X1 U798 ( .A1(n1117), .A2(n1108), .ZN(n1116) );
NOR2_X1 U799 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XOR2_X1 U800 ( .A(n1120), .B(n1121), .Z(n1119) );
XOR2_X1 U801 ( .A(KEYINPUT22), .B(n1122), .Z(n1121) );
NOR2_X1 U802 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U803 ( .A1(n1118), .A2(n1125), .ZN(G63) );
XOR2_X1 U804 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND3_X1 U805 ( .A1(n1128), .A2(n1029), .A3(G478), .ZN(n1126) );
XNOR2_X1 U806 ( .A(KEYINPUT49), .B(n1129), .ZN(n1128) );
NOR2_X1 U807 ( .A1(n1118), .A2(n1130), .ZN(G60) );
NOR3_X1 U808 ( .A1(n1078), .A2(n1131), .A3(n1132), .ZN(n1130) );
NOR3_X1 U809 ( .A1(n1133), .A2(n1134), .A3(n1124), .ZN(n1132) );
INV_X1 U810 ( .A(G475), .ZN(n1134) );
NOR2_X1 U811 ( .A1(n1135), .A2(n1136), .ZN(n1131) );
AND2_X1 U812 ( .A1(n1029), .A2(G475), .ZN(n1135) );
XNOR2_X1 U813 ( .A(G104), .B(n1137), .ZN(G6) );
NOR2_X1 U814 ( .A1(n1118), .A2(n1138), .ZN(G57) );
XOR2_X1 U815 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U816 ( .A1(KEYINPUT7), .A2(n1141), .ZN(n1139) );
XOR2_X1 U817 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U818 ( .A(KEYINPUT61), .B(n1144), .Z(n1143) );
NOR2_X1 U819 ( .A1(n1080), .A2(n1124), .ZN(n1144) );
NOR2_X1 U820 ( .A1(n1118), .A2(n1145), .ZN(G54) );
XOR2_X1 U821 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U822 ( .A1(n1077), .A2(n1124), .ZN(n1147) );
NOR2_X1 U823 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
XOR2_X1 U824 ( .A(KEYINPUT27), .B(n1150), .Z(n1149) );
NOR2_X1 U825 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
AND2_X1 U826 ( .A1(n1151), .A2(n1152), .ZN(n1148) );
XOR2_X1 U827 ( .A(n1153), .B(n1154), .Z(n1152) );
XNOR2_X1 U828 ( .A(KEYINPUT62), .B(n1155), .ZN(n1153) );
NOR2_X1 U829 ( .A1(KEYINPUT0), .A2(n1156), .ZN(n1155) );
XNOR2_X1 U830 ( .A(G110), .B(G140), .ZN(n1156) );
NOR2_X1 U831 ( .A1(n1118), .A2(n1157), .ZN(G51) );
XOR2_X1 U832 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U833 ( .A1(n1160), .A2(n1124), .ZN(n1159) );
NAND2_X1 U834 ( .A1(G902), .A2(n1029), .ZN(n1124) );
NAND3_X1 U835 ( .A1(n1101), .A2(n1161), .A3(n1115), .ZN(n1029) );
AND4_X1 U836 ( .A1(n1137), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1115) );
AND4_X1 U837 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
NAND3_X1 U838 ( .A1(n1169), .A2(n1022), .A3(n1062), .ZN(n1137) );
XNOR2_X1 U839 ( .A(KEYINPUT17), .B(n1025), .ZN(n1161) );
NAND3_X1 U840 ( .A1(n1023), .A2(n1022), .A3(n1169), .ZN(n1025) );
AND4_X1 U841 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1101) );
NOR4_X1 U842 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1173) );
INV_X1 U843 ( .A(n1178), .ZN(n1174) );
AND2_X1 U844 ( .A1(n1179), .A2(n1180), .ZN(n1172) );
NOR2_X1 U845 ( .A1(n1181), .A2(n1182), .ZN(n1158) );
XOR2_X1 U846 ( .A(n1183), .B(KEYINPUT39), .Z(n1182) );
NAND2_X1 U847 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
XNOR2_X1 U848 ( .A(n1186), .B(KEYINPUT26), .ZN(n1184) );
NOR2_X1 U849 ( .A1(n1186), .A2(n1185), .ZN(n1181) );
AND2_X1 U850 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
OR2_X1 U851 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U852 ( .A1(n1191), .A2(n1189), .ZN(n1187) );
XOR2_X1 U853 ( .A(n1192), .B(n1193), .Z(n1189) );
NOR2_X1 U854 ( .A1(KEYINPUT54), .A2(n1095), .ZN(n1193) );
XNOR2_X1 U855 ( .A(G125), .B(KEYINPUT28), .ZN(n1192) );
XNOR2_X1 U856 ( .A(n1190), .B(KEYINPUT50), .ZN(n1191) );
NOR2_X1 U857 ( .A1(n1085), .A2(G952), .ZN(n1118) );
XNOR2_X1 U858 ( .A(n1194), .B(n1176), .ZN(G48) );
AND3_X1 U859 ( .A1(n1062), .A2(n1051), .A3(n1195), .ZN(n1176) );
XNOR2_X1 U860 ( .A(G143), .B(n1171), .ZN(G45) );
NAND4_X1 U861 ( .A1(n1196), .A2(n1066), .A3(n1197), .A4(n1198), .ZN(n1171) );
NOR2_X1 U862 ( .A1(n1199), .A2(n1020), .ZN(n1197) );
XOR2_X1 U863 ( .A(G140), .B(n1175), .Z(G42) );
AND2_X1 U864 ( .A1(n1200), .A2(n1201), .ZN(n1175) );
XNOR2_X1 U865 ( .A(G137), .B(n1180), .ZN(G39) );
NAND3_X1 U866 ( .A1(n1035), .A2(n1052), .A3(n1195), .ZN(n1180) );
XNOR2_X1 U867 ( .A(G134), .B(n1179), .ZN(G36) );
NAND4_X1 U868 ( .A1(n1196), .A2(n1066), .A3(n1052), .A4(n1023), .ZN(n1179) );
XNOR2_X1 U869 ( .A(G131), .B(n1178), .ZN(G33) );
NAND2_X1 U870 ( .A1(n1200), .A2(n1066), .ZN(n1178) );
AND3_X1 U871 ( .A1(n1062), .A2(n1052), .A3(n1196), .ZN(n1200) );
INV_X1 U872 ( .A(n1074), .ZN(n1052) );
NAND2_X1 U873 ( .A1(n1049), .A2(n1202), .ZN(n1074) );
NAND2_X1 U874 ( .A1(G214), .A2(n1048), .ZN(n1202) );
XOR2_X1 U875 ( .A(n1203), .B(G128), .Z(G30) );
NAND2_X1 U876 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NAND3_X1 U877 ( .A1(n1051), .A2(n1206), .A3(n1207), .ZN(n1205) );
INV_X1 U878 ( .A(KEYINPUT34), .ZN(n1207) );
NAND2_X1 U879 ( .A1(n1177), .A2(KEYINPUT34), .ZN(n1204) );
NOR2_X1 U880 ( .A1(n1206), .A2(n1020), .ZN(n1177) );
INV_X1 U881 ( .A(n1051), .ZN(n1020) );
NAND2_X1 U882 ( .A1(n1195), .A2(n1023), .ZN(n1206) );
AND3_X1 U883 ( .A1(n1073), .A2(n1208), .A3(n1196), .ZN(n1195) );
AND2_X1 U884 ( .A1(n1024), .A2(n1209), .ZN(n1196) );
XNOR2_X1 U885 ( .A(n1210), .B(n1211), .ZN(G3) );
NAND2_X1 U886 ( .A1(n1212), .A2(n1213), .ZN(n1210) );
OR2_X1 U887 ( .A1(n1163), .A2(KEYINPUT14), .ZN(n1213) );
NAND3_X1 U888 ( .A1(n1035), .A2(n1169), .A3(n1066), .ZN(n1163) );
NAND4_X1 U889 ( .A1(n1169), .A2(n1214), .A3(n1066), .A4(KEYINPUT14), .ZN(n1212) );
INV_X1 U890 ( .A(n1035), .ZN(n1214) );
XNOR2_X1 U891 ( .A(G125), .B(n1170), .ZN(G27) );
NAND4_X1 U892 ( .A1(n1062), .A2(n1041), .A3(n1215), .A4(n1201), .ZN(n1170) );
AND2_X1 U893 ( .A1(n1209), .A2(n1051), .ZN(n1215) );
NAND2_X1 U894 ( .A1(n1039), .A2(n1216), .ZN(n1209) );
NAND3_X1 U895 ( .A1(G902), .A2(n1217), .A3(n1091), .ZN(n1216) );
NOR2_X1 U896 ( .A1(n1085), .A2(G900), .ZN(n1091) );
XOR2_X1 U897 ( .A(n1218), .B(n1219), .Z(G24) );
XNOR2_X1 U898 ( .A(KEYINPUT40), .B(n1220), .ZN(n1219) );
NOR2_X1 U899 ( .A1(KEYINPUT8), .A2(n1162), .ZN(n1218) );
NAND4_X1 U900 ( .A1(n1198), .A2(n1221), .A3(n1022), .A4(n1075), .ZN(n1162) );
NOR2_X1 U901 ( .A1(n1208), .A2(n1073), .ZN(n1022) );
XNOR2_X1 U902 ( .A(G119), .B(n1168), .ZN(G21) );
NAND4_X1 U903 ( .A1(n1221), .A2(n1035), .A3(n1073), .A4(n1208), .ZN(n1168) );
INV_X1 U904 ( .A(n1222), .ZN(n1208) );
XOR2_X1 U905 ( .A(G116), .B(n1223), .Z(G18) );
NOR2_X1 U906 ( .A1(KEYINPUT47), .A2(n1167), .ZN(n1223) );
NAND3_X1 U907 ( .A1(n1066), .A2(n1023), .A3(n1221), .ZN(n1167) );
NOR2_X1 U908 ( .A1(n1198), .A2(n1199), .ZN(n1023) );
INV_X1 U909 ( .A(n1075), .ZN(n1199) );
NAND2_X1 U910 ( .A1(n1224), .A2(n1225), .ZN(G15) );
NAND2_X1 U911 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
INV_X1 U912 ( .A(n1166), .ZN(n1227) );
XNOR2_X1 U913 ( .A(G113), .B(KEYINPUT37), .ZN(n1226) );
XOR2_X1 U914 ( .A(n1228), .B(KEYINPUT45), .Z(n1224) );
NAND2_X1 U915 ( .A1(n1229), .A2(n1166), .ZN(n1228) );
NAND3_X1 U916 ( .A1(n1221), .A2(n1066), .A3(n1062), .ZN(n1166) );
NOR2_X1 U917 ( .A1(n1230), .A2(n1075), .ZN(n1062) );
NOR2_X1 U918 ( .A1(n1073), .A2(n1222), .ZN(n1066) );
AND3_X1 U919 ( .A1(n1051), .A2(n1021), .A3(n1041), .ZN(n1221) );
AND2_X1 U920 ( .A1(n1057), .A2(n1231), .ZN(n1041) );
XNOR2_X1 U921 ( .A(KEYINPUT33), .B(n1232), .ZN(n1229) );
INV_X1 U922 ( .A(G113), .ZN(n1232) );
XNOR2_X1 U923 ( .A(n1233), .B(n1165), .ZN(G12) );
NAND3_X1 U924 ( .A1(n1201), .A2(n1169), .A3(n1035), .ZN(n1165) );
NOR2_X1 U925 ( .A1(n1075), .A2(n1198), .ZN(n1035) );
INV_X1 U926 ( .A(n1230), .ZN(n1198) );
XOR2_X1 U927 ( .A(n1078), .B(n1234), .Z(n1230) );
NOR2_X1 U928 ( .A1(G475), .A2(KEYINPUT48), .ZN(n1234) );
NOR2_X1 U929 ( .A1(n1136), .A2(G902), .ZN(n1078) );
INV_X1 U930 ( .A(n1133), .ZN(n1136) );
XNOR2_X1 U931 ( .A(n1235), .B(n1236), .ZN(n1133) );
XOR2_X1 U932 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U933 ( .A(n1239), .B(n1240), .Z(n1238) );
NOR2_X1 U934 ( .A1(KEYINPUT38), .A2(n1241), .ZN(n1240) );
XOR2_X1 U935 ( .A(n1242), .B(n1243), .Z(n1241) );
NOR2_X1 U936 ( .A1(KEYINPUT23), .A2(G104), .ZN(n1243) );
XNOR2_X1 U937 ( .A(G113), .B(G122), .ZN(n1242) );
NAND2_X1 U938 ( .A1(n1244), .A2(G214), .ZN(n1239) );
XNOR2_X1 U939 ( .A(G131), .B(G125), .ZN(n1237) );
XOR2_X1 U940 ( .A(n1245), .B(n1246), .Z(n1235) );
XNOR2_X1 U941 ( .A(KEYINPUT43), .B(n1194), .ZN(n1246) );
XNOR2_X1 U942 ( .A(G143), .B(G140), .ZN(n1245) );
XNOR2_X1 U943 ( .A(n1247), .B(G478), .ZN(n1075) );
NAND2_X1 U944 ( .A1(n1127), .A2(n1129), .ZN(n1247) );
XNOR2_X1 U945 ( .A(n1248), .B(n1249), .ZN(n1127) );
XOR2_X1 U946 ( .A(n1250), .B(n1251), .Z(n1249) );
NOR2_X1 U947 ( .A1(KEYINPUT36), .A2(n1220), .ZN(n1251) );
AND2_X1 U948 ( .A1(n1252), .A2(G217), .ZN(n1250) );
XOR2_X1 U949 ( .A(n1253), .B(n1254), .Z(n1248) );
XNOR2_X1 U950 ( .A(G116), .B(n1255), .ZN(n1254) );
NAND3_X1 U951 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1253) );
NAND2_X1 U952 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NAND2_X1 U953 ( .A1(n1261), .A2(n1262), .ZN(n1257) );
INV_X1 U954 ( .A(KEYINPUT25), .ZN(n1262) );
NAND2_X1 U955 ( .A1(n1263), .A2(G134), .ZN(n1261) );
XNOR2_X1 U956 ( .A(KEYINPUT11), .B(n1264), .ZN(n1263) );
NAND2_X1 U957 ( .A1(KEYINPUT25), .A2(n1265), .ZN(n1256) );
NAND2_X1 U958 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
OR2_X1 U959 ( .A1(n1264), .A2(KEYINPUT11), .ZN(n1267) );
NAND3_X1 U960 ( .A1(G134), .A2(n1264), .A3(KEYINPUT11), .ZN(n1266) );
AND3_X1 U961 ( .A1(n1024), .A2(n1021), .A3(n1051), .ZN(n1169) );
NOR2_X1 U962 ( .A1(n1049), .A2(n1268), .ZN(n1051) );
AND2_X1 U963 ( .A1(G214), .A2(n1048), .ZN(n1268) );
XNOR2_X1 U964 ( .A(n1269), .B(n1160), .ZN(n1049) );
NAND2_X1 U965 ( .A1(G210), .A2(n1048), .ZN(n1160) );
NAND2_X1 U966 ( .A1(n1270), .A2(n1129), .ZN(n1048) );
XNOR2_X1 U967 ( .A(G237), .B(KEYINPUT31), .ZN(n1270) );
NAND2_X1 U968 ( .A1(n1271), .A2(n1129), .ZN(n1269) );
XOR2_X1 U969 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U970 ( .A(n1095), .B(n1274), .Z(n1273) );
XOR2_X1 U971 ( .A(n1185), .B(n1275), .Z(n1274) );
NAND2_X1 U972 ( .A1(KEYINPUT3), .A2(n1190), .ZN(n1275) );
NOR2_X1 U973 ( .A1(n1117), .A2(G953), .ZN(n1190) );
INV_X1 U974 ( .A(G224), .ZN(n1117) );
NAND2_X1 U975 ( .A1(n1276), .A2(n1277), .ZN(n1185) );
NAND2_X1 U976 ( .A1(n1278), .A2(n1111), .ZN(n1277) );
XOR2_X1 U977 ( .A(n1279), .B(KEYINPUT10), .Z(n1276) );
NAND2_X1 U978 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
XNOR2_X1 U979 ( .A(KEYINPUT58), .B(n1282), .ZN(n1281) );
INV_X1 U980 ( .A(n1111), .ZN(n1282) );
XOR2_X1 U981 ( .A(G110), .B(n1283), .Z(n1111) );
XNOR2_X1 U982 ( .A(KEYINPUT9), .B(n1220), .ZN(n1283) );
INV_X1 U983 ( .A(G122), .ZN(n1220) );
XOR2_X1 U984 ( .A(n1278), .B(KEYINPUT4), .Z(n1280) );
XNOR2_X1 U985 ( .A(n1112), .B(n1284), .ZN(n1278) );
NOR2_X1 U986 ( .A1(KEYINPUT30), .A2(n1110), .ZN(n1284) );
XOR2_X1 U987 ( .A(n1255), .B(n1285), .Z(n1110) );
XOR2_X1 U988 ( .A(n1286), .B(n1287), .Z(n1272) );
XOR2_X1 U989 ( .A(KEYINPUT53), .B(G125), .Z(n1287) );
XOR2_X1 U990 ( .A(KEYINPUT63), .B(KEYINPUT55), .Z(n1286) );
NAND2_X1 U991 ( .A1(n1039), .A2(n1288), .ZN(n1021) );
NAND4_X1 U992 ( .A1(G953), .A2(G902), .A3(n1217), .A4(n1108), .ZN(n1288) );
INV_X1 U993 ( .A(G898), .ZN(n1108) );
INV_X1 U994 ( .A(n1044), .ZN(n1039) );
NOR3_X1 U995 ( .A1(n1031), .A2(n1289), .A3(n1030), .ZN(n1044) );
INV_X1 U996 ( .A(G952), .ZN(n1030) );
INV_X1 U997 ( .A(n1217), .ZN(n1289) );
NAND2_X1 U998 ( .A1(G234), .A2(G237), .ZN(n1217) );
XOR2_X1 U999 ( .A(G953), .B(KEYINPUT13), .Z(n1031) );
NOR2_X1 U1000 ( .A1(n1057), .A2(n1056), .ZN(n1024) );
INV_X1 U1001 ( .A(n1231), .ZN(n1056) );
NAND2_X1 U1002 ( .A1(G221), .A2(n1290), .ZN(n1231) );
XOR2_X1 U1003 ( .A(n1291), .B(n1076), .Z(n1057) );
NAND3_X1 U1004 ( .A1(n1292), .A2(n1293), .A3(n1129), .ZN(n1076) );
NAND2_X1 U1005 ( .A1(n1294), .A2(n1154), .ZN(n1293) );
XOR2_X1 U1006 ( .A(n1151), .B(n1295), .Z(n1294) );
NOR2_X1 U1007 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
NAND2_X1 U1008 ( .A1(n1298), .A2(n1299), .ZN(n1292) );
INV_X1 U1009 ( .A(n1154), .ZN(n1299) );
NAND2_X1 U1010 ( .A1(G227), .A2(n1085), .ZN(n1154) );
XOR2_X1 U1011 ( .A(n1151), .B(n1300), .Z(n1298) );
NOR2_X1 U1012 ( .A1(n1301), .A2(n1297), .ZN(n1300) );
INV_X1 U1013 ( .A(KEYINPUT51), .ZN(n1297) );
XOR2_X1 U1014 ( .A(n1296), .B(KEYINPUT52), .Z(n1301) );
NAND2_X1 U1015 ( .A1(n1302), .A2(n1303), .ZN(n1296) );
NAND2_X1 U1016 ( .A1(G110), .A2(n1304), .ZN(n1303) );
XOR2_X1 U1017 ( .A(KEYINPUT41), .B(n1305), .Z(n1302) );
NOR2_X1 U1018 ( .A1(G110), .A2(n1304), .ZN(n1305) );
XOR2_X1 U1019 ( .A(KEYINPUT16), .B(G140), .Z(n1304) );
XOR2_X1 U1020 ( .A(n1306), .B(n1307), .Z(n1151) );
NAND2_X1 U1021 ( .A1(n1308), .A2(n1309), .ZN(n1306) );
NAND2_X1 U1022 ( .A1(n1285), .A2(G107), .ZN(n1309) );
NAND2_X1 U1023 ( .A1(n1310), .A2(n1255), .ZN(n1308) );
INV_X1 U1024 ( .A(G107), .ZN(n1255) );
XNOR2_X1 U1025 ( .A(n1285), .B(KEYINPUT60), .ZN(n1310) );
XNOR2_X1 U1026 ( .A(G104), .B(n1211), .ZN(n1285) );
NAND2_X1 U1027 ( .A1(KEYINPUT20), .A2(n1077), .ZN(n1291) );
INV_X1 U1028 ( .A(G469), .ZN(n1077) );
INV_X1 U1029 ( .A(n1065), .ZN(n1201) );
NAND2_X1 U1030 ( .A1(n1222), .A2(n1073), .ZN(n1065) );
XOR2_X1 U1031 ( .A(n1311), .B(n1123), .Z(n1073) );
NAND2_X1 U1032 ( .A1(G217), .A2(n1290), .ZN(n1123) );
NAND2_X1 U1033 ( .A1(G234), .A2(n1129), .ZN(n1290) );
NAND2_X1 U1034 ( .A1(n1120), .A2(n1129), .ZN(n1311) );
XOR2_X1 U1035 ( .A(n1312), .B(n1313), .Z(n1120) );
XOR2_X1 U1036 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1037 ( .A(n1316), .B(n1317), .Z(n1315) );
NOR2_X1 U1038 ( .A1(G125), .A2(n1318), .ZN(n1317) );
XNOR2_X1 U1039 ( .A(KEYINPUT19), .B(KEYINPUT1), .ZN(n1318) );
NAND2_X1 U1040 ( .A1(n1252), .A2(G221), .ZN(n1316) );
AND2_X1 U1041 ( .A1(G234), .A2(n1085), .ZN(n1252) );
INV_X1 U1042 ( .A(G953), .ZN(n1085) );
XNOR2_X1 U1043 ( .A(n1319), .B(n1320), .ZN(n1314) );
NOR2_X1 U1044 ( .A1(KEYINPUT42), .A2(G137), .ZN(n1320) );
NOR2_X1 U1045 ( .A1(KEYINPUT5), .A2(n1321), .ZN(n1319) );
XNOR2_X1 U1046 ( .A(KEYINPUT56), .B(n1194), .ZN(n1321) );
INV_X1 U1047 ( .A(G146), .ZN(n1194) );
XOR2_X1 U1048 ( .A(n1322), .B(n1323), .Z(n1312) );
XOR2_X1 U1049 ( .A(G140), .B(G128), .Z(n1323) );
XNOR2_X1 U1050 ( .A(G119), .B(G110), .ZN(n1322) );
XOR2_X1 U1051 ( .A(n1081), .B(n1080), .Z(n1222) );
INV_X1 U1052 ( .A(G472), .ZN(n1080) );
AND2_X1 U1053 ( .A1(n1324), .A2(n1129), .ZN(n1081) );
INV_X1 U1054 ( .A(G902), .ZN(n1129) );
XOR2_X1 U1055 ( .A(n1325), .B(n1140), .Z(n1324) );
AND2_X1 U1056 ( .A1(n1326), .A2(n1327), .ZN(n1140) );
NAND2_X1 U1057 ( .A1(n1328), .A2(n1211), .ZN(n1327) );
INV_X1 U1058 ( .A(G101), .ZN(n1211) );
NAND2_X1 U1059 ( .A1(n1244), .A2(G210), .ZN(n1328) );
NAND3_X1 U1060 ( .A1(n1244), .A2(G210), .A3(G101), .ZN(n1326) );
NOR2_X1 U1061 ( .A1(G953), .A2(G237), .ZN(n1244) );
NAND2_X1 U1062 ( .A1(n1329), .A2(KEYINPUT59), .ZN(n1325) );
XOR2_X1 U1063 ( .A(n1142), .B(KEYINPUT18), .Z(n1329) );
XNOR2_X1 U1064 ( .A(n1307), .B(n1112), .ZN(n1142) );
XOR2_X1 U1065 ( .A(G113), .B(n1330), .Z(n1112) );
XOR2_X1 U1066 ( .A(G119), .B(G116), .Z(n1330) );
XNOR2_X1 U1067 ( .A(n1331), .B(n1332), .ZN(n1307) );
XOR2_X1 U1068 ( .A(n1098), .B(n1095), .Z(n1332) );
XOR2_X1 U1069 ( .A(G146), .B(n1264), .Z(n1095) );
INV_X1 U1070 ( .A(n1259), .ZN(n1264) );
XOR2_X1 U1071 ( .A(G128), .B(n1333), .Z(n1259) );
INV_X1 U1072 ( .A(G143), .ZN(n1333) );
XNOR2_X1 U1073 ( .A(G137), .B(n1260), .ZN(n1098) );
INV_X1 U1074 ( .A(G134), .ZN(n1260) );
XNOR2_X1 U1075 ( .A(n1334), .B(n1335), .ZN(n1331) );
INV_X1 U1076 ( .A(G131), .ZN(n1335) );
XNOR2_X1 U1077 ( .A(KEYINPUT35), .B(KEYINPUT12), .ZN(n1334) );
NAND2_X1 U1078 ( .A1(KEYINPUT46), .A2(n1336), .ZN(n1233) );
INV_X1 U1079 ( .A(G110), .ZN(n1336) );
endmodule


