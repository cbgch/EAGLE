//Key = 0010111000011100011001011100000111001000011000000110010000001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457;

XNOR2_X1 U783 ( .A(G107), .B(n1098), .ZN(G9) );
NOR2_X1 U784 ( .A1(n1099), .A2(n1100), .ZN(G75) );
NOR4_X1 U785 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1100) );
NOR4_X1 U786 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1102) );
INV_X1 U787 ( .A(n1109), .ZN(n1108) );
NOR3_X1 U788 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1106) );
NOR2_X1 U789 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U790 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NOR2_X1 U791 ( .A1(KEYINPUT22), .A2(n1117), .ZN(n1115) );
NOR2_X1 U792 ( .A1(n1118), .A2(n1119), .ZN(n1111) );
NOR2_X1 U793 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
NOR2_X1 U794 ( .A1(n1122), .A2(n1123), .ZN(n1105) );
AND3_X1 U795 ( .A1(KEYINPUT22), .A2(n1124), .A3(n1125), .ZN(n1123) );
INV_X1 U796 ( .A(n1110), .ZN(n1122) );
NOR4_X1 U797 ( .A1(n1126), .A2(n1119), .A3(n1114), .A4(n1110), .ZN(n1101) );
NOR2_X1 U798 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U799 ( .A1(n1129), .A2(n1107), .ZN(n1128) );
NOR2_X1 U800 ( .A1(n1130), .A2(n1131), .ZN(n1127) );
NOR2_X1 U801 ( .A1(n1132), .A2(n1133), .ZN(n1130) );
NOR2_X1 U802 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NOR2_X1 U803 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NOR3_X1 U804 ( .A1(n1138), .A2(KEYINPUT54), .A3(n1139), .ZN(n1136) );
NOR2_X1 U805 ( .A1(n1140), .A2(n1107), .ZN(n1132) );
NOR2_X1 U806 ( .A1(n1134), .A2(KEYINPUT54), .ZN(n1140) );
NOR2_X1 U807 ( .A1(G952), .A2(n1103), .ZN(n1099) );
NAND2_X1 U808 ( .A1(n1141), .A2(n1142), .ZN(n1103) );
NAND4_X1 U809 ( .A1(n1143), .A2(n1144), .A3(n1109), .A4(n1145), .ZN(n1142) );
NOR4_X1 U810 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1145) );
XOR2_X1 U811 ( .A(n1150), .B(n1151), .Z(n1149) );
XNOR2_X1 U812 ( .A(KEYINPUT57), .B(KEYINPUT18), .ZN(n1150) );
NOR2_X1 U813 ( .A1(n1152), .A2(n1153), .ZN(n1148) );
XNOR2_X1 U814 ( .A(G475), .B(n1154), .ZN(n1153) );
XNOR2_X1 U815 ( .A(KEYINPUT44), .B(KEYINPUT4), .ZN(n1154) );
INV_X1 U816 ( .A(n1155), .ZN(n1152) );
NOR3_X1 U817 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1147) );
NOR2_X1 U818 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
AND3_X1 U819 ( .A1(n1160), .A2(n1159), .A3(KEYINPUT49), .ZN(n1157) );
NOR2_X1 U820 ( .A1(n1161), .A2(KEYINPUT8), .ZN(n1159) );
NOR2_X1 U821 ( .A1(KEYINPUT49), .A2(n1162), .ZN(n1156) );
INV_X1 U822 ( .A(n1161), .ZN(n1162) );
XOR2_X1 U823 ( .A(n1163), .B(n1164), .Z(G72) );
NOR2_X1 U824 ( .A1(n1165), .A2(n1141), .ZN(n1164) );
NOR2_X1 U825 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NAND2_X1 U826 ( .A1(n1168), .A2(n1169), .ZN(n1163) );
NAND3_X1 U827 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1169) );
NAND2_X1 U828 ( .A1(G953), .A2(n1167), .ZN(n1171) );
NAND2_X1 U829 ( .A1(n1173), .A2(n1141), .ZN(n1170) );
XOR2_X1 U830 ( .A(n1174), .B(KEYINPUT3), .Z(n1168) );
NAND3_X1 U831 ( .A1(n1173), .A2(n1141), .A3(n1175), .ZN(n1174) );
INV_X1 U832 ( .A(n1172), .ZN(n1175) );
XOR2_X1 U833 ( .A(n1176), .B(n1177), .Z(n1172) );
XOR2_X1 U834 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U835 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U836 ( .A(n1182), .B(G131), .Z(n1176) );
XNOR2_X1 U837 ( .A(KEYINPUT15), .B(KEYINPUT1), .ZN(n1182) );
NAND2_X1 U838 ( .A1(n1183), .A2(n1184), .ZN(n1173) );
XOR2_X1 U839 ( .A(KEYINPUT51), .B(n1185), .Z(n1184) );
NAND2_X1 U840 ( .A1(n1186), .A2(n1187), .ZN(G69) );
NAND4_X1 U841 ( .A1(G953), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1187) );
INV_X1 U842 ( .A(KEYINPUT61), .ZN(n1190) );
NAND4_X1 U843 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1186) );
NAND3_X1 U844 ( .A1(n1195), .A2(n1196), .A3(n1141), .ZN(n1194) );
NAND2_X1 U845 ( .A1(G953), .A2(n1197), .ZN(n1193) );
NAND2_X1 U846 ( .A1(n1195), .A2(n1198), .ZN(n1197) );
NAND2_X1 U847 ( .A1(n1199), .A2(n1188), .ZN(n1198) );
NAND2_X1 U848 ( .A1(KEYINPUT48), .A2(n1199), .ZN(n1192) );
NAND3_X1 U849 ( .A1(n1200), .A2(n1188), .A3(G953), .ZN(n1199) );
NAND2_X1 U850 ( .A1(G898), .A2(G224), .ZN(n1188) );
OR2_X1 U851 ( .A1(KEYINPUT48), .A2(KEYINPUT61), .ZN(n1200) );
OR2_X1 U852 ( .A1(n1196), .A2(n1195), .ZN(n1191) );
INV_X1 U853 ( .A(n1189), .ZN(n1195) );
NAND2_X1 U854 ( .A1(n1201), .A2(n1202), .ZN(n1189) );
NAND2_X1 U855 ( .A1(G953), .A2(n1203), .ZN(n1202) );
XNOR2_X1 U856 ( .A(n1204), .B(n1205), .ZN(n1201) );
XNOR2_X1 U857 ( .A(n1206), .B(n1207), .ZN(n1205) );
NOR2_X1 U858 ( .A1(KEYINPUT52), .A2(n1208), .ZN(n1207) );
NAND2_X1 U859 ( .A1(KEYINPUT42), .A2(n1209), .ZN(n1206) );
NAND3_X1 U860 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1196) );
XOR2_X1 U861 ( .A(n1213), .B(KEYINPUT12), .Z(n1212) );
NAND2_X1 U862 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U863 ( .A(n1216), .B(KEYINPUT19), .Z(n1214) );
XOR2_X1 U864 ( .A(n1217), .B(KEYINPUT43), .Z(n1210) );
NOR2_X1 U865 ( .A1(n1218), .A2(n1219), .ZN(G66) );
NOR3_X1 U866 ( .A1(n1161), .A2(n1220), .A3(n1221), .ZN(n1219) );
NOR3_X1 U867 ( .A1(n1222), .A2(n1160), .A3(n1223), .ZN(n1221) );
NOR2_X1 U868 ( .A1(n1224), .A2(n1225), .ZN(n1220) );
NOR2_X1 U869 ( .A1(n1226), .A2(n1160), .ZN(n1224) );
INV_X1 U870 ( .A(n1104), .ZN(n1226) );
NOR2_X1 U871 ( .A1(n1218), .A2(n1227), .ZN(G63) );
XOR2_X1 U872 ( .A(n1228), .B(n1229), .Z(n1227) );
AND2_X1 U873 ( .A1(G478), .A2(n1230), .ZN(n1229) );
NOR2_X1 U874 ( .A1(n1218), .A2(n1231), .ZN(G60) );
XOR2_X1 U875 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U876 ( .A(KEYINPUT5), .B(n1234), .Z(n1233) );
AND2_X1 U877 ( .A1(G475), .A2(n1230), .ZN(n1234) );
XNOR2_X1 U878 ( .A(G104), .B(n1216), .ZN(G6) );
NOR2_X1 U879 ( .A1(n1218), .A2(n1235), .ZN(G57) );
XOR2_X1 U880 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U881 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U882 ( .A(G101), .B(n1240), .Z(n1239) );
NOR2_X1 U883 ( .A1(KEYINPUT59), .A2(n1241), .ZN(n1240) );
NOR2_X1 U884 ( .A1(n1242), .A2(KEYINPUT29), .ZN(n1238) );
AND2_X1 U885 ( .A1(G472), .A2(n1230), .ZN(n1242) );
XOR2_X1 U886 ( .A(n1243), .B(n1244), .Z(n1236) );
XOR2_X1 U887 ( .A(n1209), .B(n1245), .Z(n1243) );
NOR2_X1 U888 ( .A1(n1218), .A2(n1246), .ZN(G54) );
XOR2_X1 U889 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U890 ( .A(n1249), .B(n1250), .Z(n1248) );
NOR2_X1 U891 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NOR2_X1 U892 ( .A1(n1253), .A2(n1254), .ZN(n1251) );
XNOR2_X1 U893 ( .A(n1255), .B(n1256), .ZN(n1247) );
AND2_X1 U894 ( .A1(G469), .A2(n1230), .ZN(n1256) );
NOR2_X1 U895 ( .A1(n1218), .A2(n1257), .ZN(G51) );
XOR2_X1 U896 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U897 ( .A(n1260), .B(n1261), .Z(n1259) );
NOR2_X1 U898 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XOR2_X1 U899 ( .A(n1264), .B(KEYINPUT31), .Z(n1263) );
NAND2_X1 U900 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NOR2_X1 U901 ( .A1(n1265), .A2(n1266), .ZN(n1262) );
XOR2_X1 U902 ( .A(G125), .B(n1267), .Z(n1266) );
NOR2_X1 U903 ( .A1(KEYINPUT45), .A2(n1244), .ZN(n1267) );
NAND3_X1 U904 ( .A1(n1230), .A2(G210), .A3(KEYINPUT25), .ZN(n1258) );
INV_X1 U905 ( .A(n1223), .ZN(n1230) );
NAND2_X1 U906 ( .A1(G902), .A2(n1104), .ZN(n1223) );
NAND4_X1 U907 ( .A1(n1216), .A2(n1217), .A3(n1215), .A4(n1268), .ZN(n1104) );
AND3_X1 U908 ( .A1(n1185), .A2(n1211), .A3(n1183), .ZN(n1268) );
AND3_X1 U909 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1183) );
NAND2_X1 U910 ( .A1(n1121), .A2(n1272), .ZN(n1271) );
NAND2_X1 U911 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND3_X1 U912 ( .A1(n1125), .A2(n1144), .A3(n1275), .ZN(n1274) );
NAND2_X1 U913 ( .A1(n1116), .A2(n1276), .ZN(n1273) );
NAND2_X1 U914 ( .A1(n1277), .A2(n1278), .ZN(n1269) );
INV_X1 U915 ( .A(n1279), .ZN(n1278) );
XOR2_X1 U916 ( .A(n1280), .B(KEYINPUT11), .Z(n1277) );
NOR3_X1 U917 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1211) );
NOR4_X1 U918 ( .A1(n1284), .A2(n1285), .A3(n1286), .A4(n1287), .ZN(n1185) );
INV_X1 U919 ( .A(n1288), .ZN(n1285) );
INV_X1 U920 ( .A(n1289), .ZN(n1284) );
AND3_X1 U921 ( .A1(n1290), .A2(n1098), .A3(n1291), .ZN(n1215) );
NAND3_X1 U922 ( .A1(n1125), .A2(n1124), .A3(n1292), .ZN(n1291) );
NOR3_X1 U923 ( .A1(n1129), .A2(n1293), .A3(n1294), .ZN(n1292) );
XOR2_X1 U924 ( .A(n1295), .B(KEYINPUT53), .Z(n1294) );
INV_X1 U925 ( .A(n1117), .ZN(n1125) );
NAND3_X1 U926 ( .A1(n1296), .A2(n1297), .A3(n1120), .ZN(n1098) );
NAND3_X1 U927 ( .A1(n1296), .A2(n1297), .A3(n1121), .ZN(n1216) );
INV_X1 U928 ( .A(n1119), .ZN(n1296) );
NOR2_X1 U929 ( .A1(n1141), .A2(G952), .ZN(n1218) );
XOR2_X1 U930 ( .A(n1298), .B(n1299), .Z(G48) );
NOR2_X1 U931 ( .A1(KEYINPUT28), .A2(n1300), .ZN(n1299) );
XOR2_X1 U932 ( .A(n1301), .B(KEYINPUT16), .Z(n1300) );
NAND2_X1 U933 ( .A1(n1302), .A2(n1303), .ZN(n1298) );
OR2_X1 U934 ( .A1(n1288), .A2(KEYINPUT63), .ZN(n1303) );
NAND2_X1 U935 ( .A1(n1275), .A2(n1304), .ZN(n1288) );
NAND4_X1 U936 ( .A1(n1305), .A2(n1129), .A3(n1304), .A4(KEYINPUT63), .ZN(n1302) );
NOR3_X1 U937 ( .A1(n1280), .A2(n1306), .A3(n1307), .ZN(n1304) );
XOR2_X1 U938 ( .A(n1308), .B(n1289), .Z(G45) );
NAND3_X1 U939 ( .A1(n1116), .A2(n1275), .A3(n1309), .ZN(n1289) );
NOR3_X1 U940 ( .A1(n1306), .A2(n1310), .A3(n1143), .ZN(n1309) );
XOR2_X1 U941 ( .A(G140), .B(n1286), .Z(G42) );
NOR3_X1 U942 ( .A1(n1307), .A2(n1311), .A3(n1117), .ZN(n1286) );
XOR2_X1 U943 ( .A(n1287), .B(n1312), .Z(G39) );
NOR2_X1 U944 ( .A1(KEYINPUT7), .A2(n1313), .ZN(n1312) );
INV_X1 U945 ( .A(G137), .ZN(n1313) );
NOR3_X1 U946 ( .A1(n1311), .A2(n1280), .A3(n1114), .ZN(n1287) );
NAND2_X1 U947 ( .A1(n1314), .A2(n1315), .ZN(G36) );
OR2_X1 U948 ( .A1(n1270), .A2(G134), .ZN(n1315) );
XOR2_X1 U949 ( .A(n1316), .B(KEYINPUT58), .Z(n1314) );
NAND2_X1 U950 ( .A1(G134), .A2(n1270), .ZN(n1316) );
NAND3_X1 U951 ( .A1(n1276), .A2(n1120), .A3(n1116), .ZN(n1270) );
INV_X1 U952 ( .A(n1311), .ZN(n1276) );
XOR2_X1 U953 ( .A(G131), .B(n1317), .Z(G33) );
NOR3_X1 U954 ( .A1(n1318), .A2(n1311), .A3(n1319), .ZN(n1317) );
NAND3_X1 U955 ( .A1(n1137), .A2(n1305), .A3(n1109), .ZN(n1311) );
NOR2_X1 U956 ( .A1(n1131), .A2(n1134), .ZN(n1109) );
INV_X1 U957 ( .A(n1320), .ZN(n1134) );
INV_X1 U958 ( .A(n1306), .ZN(n1137) );
XOR2_X1 U959 ( .A(KEYINPUT24), .B(n1121), .Z(n1318) );
INV_X1 U960 ( .A(n1307), .ZN(n1121) );
XOR2_X1 U961 ( .A(G128), .B(n1321), .Z(G30) );
NOR2_X1 U962 ( .A1(n1280), .A2(n1279), .ZN(n1321) );
NAND3_X1 U963 ( .A1(n1120), .A2(n1322), .A3(n1275), .ZN(n1279) );
XNOR2_X1 U964 ( .A(G101), .B(n1290), .ZN(G3) );
OR2_X1 U965 ( .A1(n1323), .A2(n1319), .ZN(n1290) );
XNOR2_X1 U966 ( .A(G125), .B(n1324), .ZN(G27) );
NAND3_X1 U967 ( .A1(KEYINPUT50), .A2(n1275), .A3(n1325), .ZN(n1324) );
NOR3_X1 U968 ( .A1(n1117), .A2(n1107), .A3(n1307), .ZN(n1325) );
AND2_X1 U969 ( .A1(n1326), .A2(n1305), .ZN(n1275) );
NAND2_X1 U970 ( .A1(n1327), .A2(n1110), .ZN(n1305) );
NAND4_X1 U971 ( .A1(G953), .A2(G902), .A3(n1328), .A4(n1167), .ZN(n1327) );
INV_X1 U972 ( .A(G900), .ZN(n1167) );
NAND2_X1 U973 ( .A1(n1329), .A2(n1330), .ZN(G24) );
NAND2_X1 U974 ( .A1(n1283), .A2(n1331), .ZN(n1330) );
XOR2_X1 U975 ( .A(KEYINPUT60), .B(n1332), .Z(n1329) );
NOR2_X1 U976 ( .A1(n1283), .A2(n1331), .ZN(n1332) );
NOR4_X1 U977 ( .A1(n1333), .A2(n1119), .A3(n1143), .A4(n1310), .ZN(n1283) );
NAND2_X1 U978 ( .A1(n1334), .A2(n1335), .ZN(n1119) );
XOR2_X1 U979 ( .A(G119), .B(n1281), .Z(G21) );
NOR3_X1 U980 ( .A1(n1114), .A2(n1280), .A3(n1333), .ZN(n1281) );
NAND2_X1 U981 ( .A1(n1336), .A2(n1151), .ZN(n1280) );
XNOR2_X1 U982 ( .A(G116), .B(n1217), .ZN(G18) );
NAND3_X1 U983 ( .A1(n1116), .A2(n1120), .A3(n1337), .ZN(n1217) );
INV_X1 U984 ( .A(n1333), .ZN(n1337) );
NOR2_X1 U985 ( .A1(n1338), .A2(n1143), .ZN(n1120) );
INV_X1 U986 ( .A(n1319), .ZN(n1116) );
NAND2_X1 U987 ( .A1(n1339), .A2(n1340), .ZN(G15) );
NAND2_X1 U988 ( .A1(n1282), .A2(n1341), .ZN(n1340) );
XOR2_X1 U989 ( .A(KEYINPUT17), .B(n1342), .Z(n1339) );
NOR2_X1 U990 ( .A1(n1282), .A2(n1341), .ZN(n1342) );
NOR3_X1 U991 ( .A1(n1319), .A2(n1307), .A3(n1333), .ZN(n1282) );
NAND3_X1 U992 ( .A1(n1326), .A2(n1295), .A3(n1144), .ZN(n1333) );
INV_X1 U993 ( .A(n1107), .ZN(n1144) );
NAND2_X1 U994 ( .A1(n1343), .A2(n1138), .ZN(n1107) );
NAND2_X1 U995 ( .A1(n1143), .A2(n1338), .ZN(n1307) );
INV_X1 U996 ( .A(n1310), .ZN(n1338) );
NAND2_X1 U997 ( .A1(n1335), .A2(n1151), .ZN(n1319) );
INV_X1 U998 ( .A(n1334), .ZN(n1151) );
XOR2_X1 U999 ( .A(G110), .B(n1344), .Z(G12) );
NOR2_X1 U1000 ( .A1(n1117), .A2(n1323), .ZN(n1344) );
NAND2_X1 U1001 ( .A1(n1124), .A2(n1297), .ZN(n1323) );
AND3_X1 U1002 ( .A1(n1322), .A2(n1295), .A3(n1326), .ZN(n1297) );
INV_X1 U1003 ( .A(n1129), .ZN(n1326) );
NAND2_X1 U1004 ( .A1(n1320), .A2(n1131), .ZN(n1129) );
NAND2_X1 U1005 ( .A1(n1345), .A2(n1346), .ZN(n1131) );
NAND3_X1 U1006 ( .A1(n1347), .A2(n1348), .A3(n1349), .ZN(n1346) );
NAND2_X1 U1007 ( .A1(KEYINPUT36), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1008 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
NAND2_X1 U1009 ( .A1(G237), .A2(G210), .ZN(n1351) );
NAND2_X1 U1010 ( .A1(n1353), .A2(n1354), .ZN(n1347) );
NAND2_X1 U1011 ( .A1(G902), .A2(n1355), .ZN(n1353) );
NAND2_X1 U1012 ( .A1(G210), .A2(n1356), .ZN(n1345) );
NAND2_X1 U1013 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
NAND2_X1 U1014 ( .A1(G237), .A2(n1359), .ZN(n1358) );
NAND2_X1 U1015 ( .A1(n1349), .A2(n1360), .ZN(n1359) );
NAND2_X1 U1016 ( .A1(n1352), .A2(n1354), .ZN(n1360) );
NAND2_X1 U1017 ( .A1(G902), .A2(n1361), .ZN(n1357) );
NAND2_X1 U1018 ( .A1(n1349), .A2(n1354), .ZN(n1361) );
INV_X1 U1019 ( .A(KEYINPUT36), .ZN(n1354) );
XNOR2_X1 U1020 ( .A(n1362), .B(n1363), .ZN(n1349) );
XOR2_X1 U1021 ( .A(n1364), .B(n1265), .Z(n1363) );
AND2_X1 U1022 ( .A1(G224), .A2(n1141), .ZN(n1265) );
NOR2_X1 U1023 ( .A1(KEYINPUT26), .A2(n1365), .ZN(n1364) );
XOR2_X1 U1024 ( .A(n1260), .B(G125), .Z(n1362) );
NAND3_X1 U1025 ( .A1(n1366), .A2(n1367), .A3(n1368), .ZN(n1260) );
NAND2_X1 U1026 ( .A1(KEYINPUT27), .A2(n1369), .ZN(n1368) );
NAND3_X1 U1027 ( .A1(n1370), .A2(n1371), .A3(n1372), .ZN(n1367) );
INV_X1 U1028 ( .A(KEYINPUT27), .ZN(n1371) );
OR2_X1 U1029 ( .A1(n1372), .A2(n1370), .ZN(n1366) );
NOR2_X1 U1030 ( .A1(KEYINPUT14), .A2(n1369), .ZN(n1370) );
XNOR2_X1 U1031 ( .A(n1209), .B(n1204), .ZN(n1369) );
XNOR2_X1 U1032 ( .A(n1373), .B(n1374), .ZN(n1204) );
XOR2_X1 U1033 ( .A(KEYINPUT2), .B(n1375), .Z(n1374) );
NOR2_X1 U1034 ( .A1(G104), .A2(n1376), .ZN(n1375) );
XNOR2_X1 U1035 ( .A(KEYINPUT46), .B(KEYINPUT23), .ZN(n1376) );
INV_X1 U1036 ( .A(n1208), .ZN(n1372) );
XNOR2_X1 U1037 ( .A(n1377), .B(G122), .ZN(n1208) );
NAND2_X1 U1038 ( .A1(G214), .A2(n1378), .ZN(n1320) );
OR2_X1 U1039 ( .A1(G237), .A2(G902), .ZN(n1378) );
NAND2_X1 U1040 ( .A1(n1110), .A2(n1379), .ZN(n1295) );
NAND4_X1 U1041 ( .A1(G953), .A2(G902), .A3(n1328), .A4(n1203), .ZN(n1379) );
INV_X1 U1042 ( .A(G898), .ZN(n1203) );
NAND3_X1 U1043 ( .A1(n1328), .A2(n1141), .A3(n1380), .ZN(n1110) );
XOR2_X1 U1044 ( .A(KEYINPUT39), .B(G952), .Z(n1380) );
NAND2_X1 U1045 ( .A1(G237), .A2(G234), .ZN(n1328) );
INV_X1 U1046 ( .A(n1293), .ZN(n1322) );
XOR2_X1 U1047 ( .A(n1306), .B(KEYINPUT35), .Z(n1293) );
NAND2_X1 U1048 ( .A1(n1139), .A2(n1138), .ZN(n1306) );
NAND2_X1 U1049 ( .A1(G221), .A2(n1381), .ZN(n1138) );
INV_X1 U1050 ( .A(n1343), .ZN(n1139) );
XOR2_X1 U1051 ( .A(n1382), .B(G469), .Z(n1343) );
NAND2_X1 U1052 ( .A1(n1383), .A2(n1352), .ZN(n1382) );
XOR2_X1 U1053 ( .A(n1384), .B(n1385), .Z(n1383) );
NAND2_X1 U1054 ( .A1(KEYINPUT41), .A2(n1386), .ZN(n1385) );
XNOR2_X1 U1055 ( .A(n1249), .B(n1387), .ZN(n1386) );
NAND2_X1 U1056 ( .A1(KEYINPUT13), .A2(n1255), .ZN(n1387) );
XOR2_X1 U1057 ( .A(G140), .B(G110), .Z(n1255) );
NOR2_X1 U1058 ( .A1(n1166), .A2(G953), .ZN(n1249) );
INV_X1 U1059 ( .A(G227), .ZN(n1166) );
NAND3_X1 U1060 ( .A1(n1388), .A2(n1389), .A3(n1390), .ZN(n1384) );
NAND2_X1 U1061 ( .A1(n1391), .A2(n1392), .ZN(n1390) );
NAND2_X1 U1062 ( .A1(KEYINPUT30), .A2(n1393), .ZN(n1389) );
NAND3_X1 U1063 ( .A1(n1394), .A2(n1395), .A3(n1254), .ZN(n1393) );
INV_X1 U1064 ( .A(n1391), .ZN(n1254) );
NOR2_X1 U1065 ( .A1(n1396), .A2(n1397), .ZN(n1391) );
NAND2_X1 U1066 ( .A1(n1392), .A2(n1245), .ZN(n1395) );
NAND3_X1 U1067 ( .A1(n1253), .A2(n1396), .A3(n1397), .ZN(n1394) );
NAND2_X1 U1068 ( .A1(n1252), .A2(n1398), .ZN(n1388) );
INV_X1 U1069 ( .A(KEYINPUT30), .ZN(n1398) );
NAND2_X1 U1070 ( .A1(n1399), .A2(n1400), .ZN(n1252) );
NAND2_X1 U1071 ( .A1(n1401), .A2(n1396), .ZN(n1400) );
XOR2_X1 U1072 ( .A(n1397), .B(n1253), .Z(n1401) );
INV_X1 U1073 ( .A(n1392), .ZN(n1253) );
OR3_X1 U1074 ( .A1(n1392), .A2(n1245), .A3(n1396), .ZN(n1399) );
XOR2_X1 U1075 ( .A(G104), .B(n1402), .Z(n1396) );
INV_X1 U1076 ( .A(n1373), .ZN(n1402) );
XNOR2_X1 U1077 ( .A(G107), .B(G101), .ZN(n1373) );
XNOR2_X1 U1078 ( .A(n1180), .B(KEYINPUT40), .ZN(n1392) );
XNOR2_X1 U1079 ( .A(n1403), .B(G128), .ZN(n1180) );
NAND2_X1 U1080 ( .A1(n1404), .A2(n1405), .ZN(n1403) );
NAND2_X1 U1081 ( .A1(n1406), .A2(n1308), .ZN(n1405) );
NAND2_X1 U1082 ( .A1(n1407), .A2(n1408), .ZN(n1406) );
NAND2_X1 U1083 ( .A1(KEYINPUT33), .A2(n1301), .ZN(n1408) );
NAND2_X1 U1084 ( .A1(G146), .A2(n1409), .ZN(n1404) );
NAND2_X1 U1085 ( .A1(KEYINPUT33), .A2(n1410), .ZN(n1409) );
NAND2_X1 U1086 ( .A1(G143), .A2(n1407), .ZN(n1410) );
INV_X1 U1087 ( .A(KEYINPUT34), .ZN(n1407) );
INV_X1 U1088 ( .A(n1114), .ZN(n1124) );
NAND2_X1 U1089 ( .A1(n1143), .A2(n1310), .ZN(n1114) );
NOR2_X1 U1090 ( .A1(n1411), .A2(n1146), .ZN(n1310) );
NOR2_X1 U1091 ( .A1(n1155), .A2(G475), .ZN(n1146) );
AND2_X1 U1092 ( .A1(G475), .A2(n1155), .ZN(n1411) );
NAND2_X1 U1093 ( .A1(n1232), .A2(n1352), .ZN(n1155) );
XOR2_X1 U1094 ( .A(n1412), .B(n1413), .Z(n1232) );
XOR2_X1 U1095 ( .A(n1414), .B(n1415), .Z(n1413) );
XNOR2_X1 U1096 ( .A(n1416), .B(n1417), .ZN(n1415) );
NOR2_X1 U1097 ( .A1(G113), .A2(KEYINPUT62), .ZN(n1417) );
NOR2_X1 U1098 ( .A1(KEYINPUT37), .A2(n1418), .ZN(n1416) );
XOR2_X1 U1099 ( .A(n1419), .B(n1420), .Z(n1418) );
NOR3_X1 U1100 ( .A1(n1421), .A2(G953), .A3(G237), .ZN(n1420) );
INV_X1 U1101 ( .A(G214), .ZN(n1421) );
XOR2_X1 U1102 ( .A(G131), .B(n1308), .Z(n1419) );
XOR2_X1 U1103 ( .A(n1422), .B(n1423), .Z(n1412) );
XOR2_X1 U1104 ( .A(KEYINPUT38), .B(G146), .Z(n1423) );
XOR2_X1 U1105 ( .A(G104), .B(n1331), .Z(n1422) );
INV_X1 U1106 ( .A(G122), .ZN(n1331) );
XNOR2_X1 U1107 ( .A(G478), .B(n1424), .ZN(n1143) );
NOR2_X1 U1108 ( .A1(n1228), .A2(G902), .ZN(n1424) );
AND2_X1 U1109 ( .A1(n1425), .A2(n1426), .ZN(n1228) );
NAND2_X1 U1110 ( .A1(n1427), .A2(n1428), .ZN(n1426) );
XOR2_X1 U1111 ( .A(KEYINPUT21), .B(n1429), .Z(n1425) );
NOR2_X1 U1112 ( .A1(n1427), .A2(n1428), .ZN(n1429) );
XOR2_X1 U1113 ( .A(n1430), .B(n1431), .Z(n1428) );
XOR2_X1 U1114 ( .A(n1432), .B(n1433), .Z(n1431) );
XOR2_X1 U1115 ( .A(G134), .B(G128), .Z(n1433) );
XOR2_X1 U1116 ( .A(KEYINPUT47), .B(G143), .Z(n1432) );
XNOR2_X1 U1117 ( .A(G107), .B(n1434), .ZN(n1430) );
XOR2_X1 U1118 ( .A(G122), .B(G116), .Z(n1434) );
AND3_X1 U1119 ( .A1(G217), .A2(n1141), .A3(G234), .ZN(n1427) );
NAND2_X1 U1120 ( .A1(n1334), .A2(n1336), .ZN(n1117) );
INV_X1 U1121 ( .A(n1335), .ZN(n1336) );
XOR2_X1 U1122 ( .A(n1161), .B(n1160), .Z(n1335) );
NAND2_X1 U1123 ( .A1(G217), .A2(n1381), .ZN(n1160) );
NAND2_X1 U1124 ( .A1(G234), .A2(n1352), .ZN(n1381) );
NOR2_X1 U1125 ( .A1(n1225), .A2(G902), .ZN(n1161) );
INV_X1 U1126 ( .A(n1222), .ZN(n1225) );
XOR2_X1 U1127 ( .A(n1435), .B(n1436), .Z(n1222) );
XOR2_X1 U1128 ( .A(n1437), .B(n1438), .Z(n1436) );
XOR2_X1 U1129 ( .A(n1439), .B(n1440), .Z(n1438) );
NOR2_X1 U1130 ( .A1(G119), .A2(KEYINPUT56), .ZN(n1440) );
NAND2_X1 U1131 ( .A1(n1441), .A2(n1442), .ZN(n1439) );
NAND2_X1 U1132 ( .A1(G146), .A2(n1178), .ZN(n1442) );
XOR2_X1 U1133 ( .A(n1443), .B(KEYINPUT10), .Z(n1441) );
NAND2_X1 U1134 ( .A1(n1414), .A2(n1301), .ZN(n1443) );
INV_X1 U1135 ( .A(G146), .ZN(n1301) );
INV_X1 U1136 ( .A(n1178), .ZN(n1414) );
XOR2_X1 U1137 ( .A(G140), .B(G125), .Z(n1178) );
NAND3_X1 U1138 ( .A1(G234), .A2(n1141), .A3(G221), .ZN(n1437) );
INV_X1 U1139 ( .A(G953), .ZN(n1141) );
XOR2_X1 U1140 ( .A(n1377), .B(n1444), .Z(n1435) );
XOR2_X1 U1141 ( .A(G137), .B(G128), .Z(n1444) );
INV_X1 U1142 ( .A(G110), .ZN(n1377) );
XOR2_X1 U1143 ( .A(n1445), .B(G472), .Z(n1334) );
NAND2_X1 U1144 ( .A1(n1446), .A2(n1352), .ZN(n1445) );
INV_X1 U1145 ( .A(G902), .ZN(n1352) );
XOR2_X1 U1146 ( .A(n1447), .B(n1448), .Z(n1446) );
XOR2_X1 U1147 ( .A(n1449), .B(n1450), .Z(n1448) );
XNOR2_X1 U1148 ( .A(G101), .B(n1241), .ZN(n1450) );
OR3_X1 U1149 ( .A1(G237), .A2(G953), .A3(n1355), .ZN(n1241) );
INV_X1 U1150 ( .A(G210), .ZN(n1355) );
NOR2_X1 U1151 ( .A1(KEYINPUT9), .A2(n1209), .ZN(n1449) );
XOR2_X1 U1152 ( .A(n1341), .B(n1451), .Z(n1209) );
XOR2_X1 U1153 ( .A(G119), .B(G116), .Z(n1451) );
INV_X1 U1154 ( .A(G113), .ZN(n1341) );
XOR2_X1 U1155 ( .A(n1452), .B(n1244), .Z(n1447) );
INV_X1 U1156 ( .A(n1365), .ZN(n1244) );
XNOR2_X1 U1157 ( .A(G128), .B(n1453), .ZN(n1365) );
NOR2_X1 U1158 ( .A1(KEYINPUT0), .A2(n1454), .ZN(n1453) );
XOR2_X1 U1159 ( .A(n1308), .B(G146), .Z(n1454) );
INV_X1 U1160 ( .A(G143), .ZN(n1308) );
NAND2_X1 U1161 ( .A1(KEYINPUT32), .A2(n1245), .ZN(n1452) );
INV_X1 U1162 ( .A(n1397), .ZN(n1245) );
XOR2_X1 U1163 ( .A(n1455), .B(n1181), .Z(n1397) );
XOR2_X1 U1164 ( .A(G137), .B(G134), .Z(n1181) );
NAND2_X1 U1165 ( .A1(n1456), .A2(n1457), .ZN(n1455) );
XOR2_X1 U1166 ( .A(KEYINPUT6), .B(KEYINPUT55), .Z(n1457) );
XNOR2_X1 U1167 ( .A(G131), .B(KEYINPUT20), .ZN(n1456) );
endmodule


