//Key = 0100010110011110101111100011111001100011111010111001010000110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381;

XOR2_X1 U756 ( .A(G107), .B(n1045), .Z(G9) );
NOR2_X1 U757 ( .A1(n1046), .A2(n1047), .ZN(G75) );
NOR4_X1 U758 ( .A1(n1048), .A2(n1049), .A3(KEYINPUT36), .A4(G953), .ZN(n1047) );
NAND3_X1 U759 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1048) );
NAND2_X1 U760 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NAND2_X1 U761 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND3_X1 U762 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
NAND3_X1 U763 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1058) );
INV_X1 U764 ( .A(n1063), .ZN(n1062) );
NAND2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1061) );
NAND2_X1 U766 ( .A1(n1066), .A2(n1067), .ZN(n1060) );
NAND3_X1 U767 ( .A1(n1065), .A2(n1068), .A3(n1066), .ZN(n1055) );
NAND2_X1 U768 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U769 ( .A1(n1059), .A2(n1071), .ZN(n1070) );
NAND2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U771 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U772 ( .A1(n1057), .A2(n1076), .ZN(n1069) );
NAND2_X1 U773 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
INV_X1 U775 ( .A(n1081), .ZN(n1053) );
NOR3_X1 U776 ( .A1(n1049), .A2(G953), .A3(G952), .ZN(n1046) );
AND4_X1 U777 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1049) );
NOR4_X1 U778 ( .A1(n1074), .A2(n1079), .A3(n1086), .A4(n1087), .ZN(n1085) );
NOR3_X1 U779 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1086) );
AND2_X1 U780 ( .A1(n1091), .A2(G478), .ZN(n1090) );
NOR3_X1 U781 ( .A1(G478), .A2(KEYINPUT50), .A3(n1091), .ZN(n1089) );
NAND2_X1 U782 ( .A1(KEYINPUT7), .A2(n1092), .ZN(n1091) );
INV_X1 U783 ( .A(n1093), .ZN(n1092) );
AND2_X1 U784 ( .A1(n1093), .A2(KEYINPUT50), .ZN(n1088) );
NOR2_X1 U785 ( .A1(n1094), .A2(n1095), .ZN(n1084) );
XOR2_X1 U786 ( .A(n1096), .B(n1097), .Z(n1095) );
XOR2_X1 U787 ( .A(n1098), .B(n1099), .Z(n1094) );
XOR2_X1 U788 ( .A(n1075), .B(KEYINPUT54), .Z(n1082) );
XOR2_X1 U789 ( .A(n1100), .B(n1101), .Z(G72) );
NOR2_X1 U790 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U791 ( .A(KEYINPUT25), .B(n1104), .Z(n1103) );
NOR2_X1 U792 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XNOR2_X1 U793 ( .A(KEYINPUT43), .B(n1107), .ZN(n1106) );
INV_X1 U794 ( .A(n1108), .ZN(n1105) );
NOR2_X1 U795 ( .A1(n1108), .A2(n1107), .ZN(n1102) );
NAND2_X1 U796 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
XOR2_X1 U797 ( .A(n1111), .B(n1112), .Z(n1109) );
XOR2_X1 U798 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U799 ( .A(n1115), .B(n1116), .Z(n1111) );
XOR2_X1 U800 ( .A(G125), .B(n1117), .Z(n1116) );
NAND2_X1 U801 ( .A1(KEYINPUT14), .A2(G140), .ZN(n1115) );
NOR2_X1 U802 ( .A1(G953), .A2(n1050), .ZN(n1108) );
NAND2_X1 U803 ( .A1(G953), .A2(n1118), .ZN(n1100) );
NAND2_X1 U804 ( .A1(G900), .A2(G227), .ZN(n1118) );
NAND2_X1 U805 ( .A1(n1119), .A2(n1120), .ZN(G69) );
NAND2_X1 U806 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U807 ( .A1(G953), .A2(n1123), .ZN(n1122) );
NAND2_X1 U808 ( .A1(n1124), .A2(n1125), .ZN(n1121) );
NAND2_X1 U809 ( .A1(n1126), .A2(n1127), .ZN(n1124) );
XOR2_X1 U810 ( .A(n1128), .B(KEYINPUT63), .Z(n1126) );
XOR2_X1 U811 ( .A(n1129), .B(KEYINPUT6), .Z(n1119) );
NAND3_X1 U812 ( .A1(n1123), .A2(n1125), .A3(G953), .ZN(n1129) );
NAND3_X1 U813 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1125) );
XOR2_X1 U814 ( .A(n1127), .B(KEYINPUT19), .Z(n1132) );
NAND2_X1 U815 ( .A1(G953), .A2(n1133), .ZN(n1131) );
XNOR2_X1 U816 ( .A(KEYINPUT63), .B(n1128), .ZN(n1130) );
XOR2_X1 U817 ( .A(n1134), .B(KEYINPUT21), .Z(n1128) );
NAND2_X1 U818 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U819 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U820 ( .A1(G898), .A2(G224), .ZN(n1123) );
NOR2_X1 U821 ( .A1(n1139), .A2(n1140), .ZN(G66) );
XOR2_X1 U822 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U823 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
NOR2_X1 U824 ( .A1(n1145), .A2(n1146), .ZN(G63) );
XOR2_X1 U825 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR3_X1 U826 ( .A1(n1149), .A2(KEYINPUT55), .A3(n1150), .ZN(n1148) );
NOR2_X1 U827 ( .A1(n1151), .A2(n1152), .ZN(n1145) );
XNOR2_X1 U828 ( .A(G952), .B(KEYINPUT46), .ZN(n1151) );
NOR2_X1 U829 ( .A1(n1139), .A2(n1153), .ZN(G60) );
XOR2_X1 U830 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U831 ( .A1(n1156), .A2(KEYINPUT60), .ZN(n1155) );
INV_X1 U832 ( .A(n1157), .ZN(n1156) );
NAND2_X1 U833 ( .A1(n1143), .A2(G475), .ZN(n1154) );
XNOR2_X1 U834 ( .A(G104), .B(n1158), .ZN(G6) );
NAND4_X1 U835 ( .A1(KEYINPUT8), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1158) );
XOR2_X1 U836 ( .A(n1065), .B(KEYINPUT57), .Z(n1160) );
NOR2_X1 U837 ( .A1(n1139), .A2(n1162), .ZN(G57) );
XOR2_X1 U838 ( .A(n1163), .B(n1164), .Z(n1162) );
XNOR2_X1 U839 ( .A(n1165), .B(n1166), .ZN(n1164) );
NAND2_X1 U840 ( .A1(KEYINPUT27), .A2(n1167), .ZN(n1166) );
XOR2_X1 U841 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U842 ( .A1(KEYINPUT15), .A2(n1170), .ZN(n1169) );
AND2_X1 U843 ( .A1(G472), .A2(n1143), .ZN(n1168) );
XOR2_X1 U844 ( .A(n1171), .B(KEYINPUT41), .Z(n1163) );
INV_X1 U845 ( .A(G101), .ZN(n1171) );
NOR2_X1 U846 ( .A1(n1139), .A2(n1172), .ZN(G54) );
XOR2_X1 U847 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U848 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U849 ( .A(n1177), .B(n1178), .Z(n1176) );
XNOR2_X1 U850 ( .A(n1179), .B(n1180), .ZN(n1175) );
NAND2_X1 U851 ( .A1(n1143), .A2(G469), .ZN(n1179) );
INV_X1 U852 ( .A(n1149), .ZN(n1143) );
XOR2_X1 U853 ( .A(n1181), .B(n1182), .Z(n1173) );
XOR2_X1 U854 ( .A(KEYINPUT37), .B(n1183), .Z(n1182) );
XOR2_X1 U855 ( .A(KEYINPUT61), .B(KEYINPUT52), .Z(n1181) );
NOR2_X1 U856 ( .A1(n1139), .A2(n1184), .ZN(G51) );
XOR2_X1 U857 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U858 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND2_X1 U859 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U860 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U861 ( .A(KEYINPUT22), .B(n1193), .Z(n1189) );
NOR2_X1 U862 ( .A1(n1191), .A2(n1194), .ZN(n1193) );
XOR2_X1 U863 ( .A(n1192), .B(KEYINPUT32), .Z(n1194) );
OR2_X1 U864 ( .A1(n1149), .A2(n1099), .ZN(n1185) );
NAND2_X1 U865 ( .A1(n1195), .A2(n1196), .ZN(n1149) );
NAND2_X1 U866 ( .A1(n1052), .A2(n1050), .ZN(n1196) );
AND4_X1 U867 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1050) );
AND4_X1 U868 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
NOR2_X1 U869 ( .A1(n1205), .A2(n1206), .ZN(n1199) );
NAND2_X1 U870 ( .A1(n1207), .A2(n1208), .ZN(n1198) );
NAND3_X1 U871 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1208) );
NAND4_X1 U872 ( .A1(KEYINPUT45), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1211) );
AND2_X1 U873 ( .A1(n1161), .A2(n1057), .ZN(n1213) );
OR3_X1 U874 ( .A1(n1215), .A2(n1216), .A3(KEYINPUT59), .ZN(n1210) );
NAND2_X1 U875 ( .A1(n1217), .A2(KEYINPUT59), .ZN(n1209) );
OR2_X1 U876 ( .A1(n1218), .A2(KEYINPUT45), .ZN(n1197) );
INV_X1 U877 ( .A(n1127), .ZN(n1052) );
NAND4_X1 U878 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1127) );
NOR4_X1 U879 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1045), .ZN(n1222) );
AND3_X1 U880 ( .A1(n1064), .A2(n1065), .A3(n1159), .ZN(n1045) );
NAND2_X1 U881 ( .A1(n1159), .A2(n1063), .ZN(n1221) );
NAND2_X1 U882 ( .A1(n1226), .A2(n1227), .ZN(n1063) );
NAND2_X1 U883 ( .A1(n1161), .A2(n1065), .ZN(n1227) );
NAND2_X1 U884 ( .A1(n1214), .A2(n1066), .ZN(n1226) );
NAND4_X1 U885 ( .A1(n1228), .A2(n1066), .A3(n1087), .A4(n1229), .ZN(n1219) );
XOR2_X1 U886 ( .A(n1230), .B(KEYINPUT58), .Z(n1195) );
NOR2_X1 U887 ( .A1(n1152), .A2(G952), .ZN(n1139) );
XOR2_X1 U888 ( .A(G146), .B(n1206), .Z(G48) );
AND3_X1 U889 ( .A1(n1207), .A2(n1161), .A3(n1231), .ZN(n1206) );
XOR2_X1 U890 ( .A(G143), .B(n1232), .Z(G45) );
NOR2_X1 U891 ( .A1(n1077), .A2(n1233), .ZN(n1232) );
XOR2_X1 U892 ( .A(KEYINPUT40), .B(n1217), .Z(n1233) );
AND2_X1 U893 ( .A1(n1234), .A2(n1216), .ZN(n1217) );
XOR2_X1 U894 ( .A(G140), .B(n1205), .Z(G42) );
AND4_X1 U895 ( .A1(n1059), .A2(n1235), .A3(n1214), .A4(n1161), .ZN(n1205) );
XNOR2_X1 U896 ( .A(G137), .B(n1204), .ZN(G39) );
NAND3_X1 U897 ( .A1(n1231), .A2(n1066), .A3(n1059), .ZN(n1204) );
XNOR2_X1 U898 ( .A(G134), .B(n1203), .ZN(G36) );
NAND3_X1 U899 ( .A1(n1234), .A2(n1064), .A3(n1059), .ZN(n1203) );
XOR2_X1 U900 ( .A(n1117), .B(n1202), .Z(G33) );
NAND3_X1 U901 ( .A1(n1234), .A2(n1161), .A3(n1059), .ZN(n1202) );
NOR2_X1 U902 ( .A1(n1236), .A2(n1079), .ZN(n1059) );
INV_X1 U903 ( .A(n1080), .ZN(n1236) );
INV_X1 U904 ( .A(n1215), .ZN(n1234) );
NAND2_X1 U905 ( .A1(n1235), .A2(n1067), .ZN(n1215) );
XNOR2_X1 U906 ( .A(G128), .B(n1201), .ZN(G30) );
NAND3_X1 U907 ( .A1(n1064), .A2(n1207), .A3(n1231), .ZN(n1201) );
AND3_X1 U908 ( .A1(n1087), .A2(n1229), .A3(n1235), .ZN(n1231) );
NOR2_X1 U909 ( .A1(n1072), .A2(n1212), .ZN(n1235) );
INV_X1 U910 ( .A(n1237), .ZN(n1072) );
XOR2_X1 U911 ( .A(G101), .B(n1225), .Z(G3) );
AND3_X1 U912 ( .A1(n1159), .A2(n1067), .A3(n1066), .ZN(n1225) );
INV_X1 U913 ( .A(n1238), .ZN(n1159) );
XOR2_X1 U914 ( .A(n1218), .B(n1239), .Z(G27) );
XOR2_X1 U915 ( .A(KEYINPUT30), .B(G125), .Z(n1239) );
NAND4_X1 U916 ( .A1(n1214), .A2(n1057), .A3(n1240), .A4(n1207), .ZN(n1218) );
NOR2_X1 U917 ( .A1(n1212), .A2(n1241), .ZN(n1240) );
INV_X1 U918 ( .A(n1161), .ZN(n1241) );
AND2_X1 U919 ( .A1(n1242), .A2(n1081), .ZN(n1212) );
NAND2_X1 U920 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
INV_X1 U921 ( .A(n1110), .ZN(n1243) );
NAND2_X1 U922 ( .A1(G953), .A2(n1245), .ZN(n1110) );
XOR2_X1 U923 ( .A(KEYINPUT26), .B(G900), .Z(n1245) );
INV_X1 U924 ( .A(n1246), .ZN(n1214) );
NAND2_X1 U925 ( .A1(n1247), .A2(n1248), .ZN(G24) );
NAND2_X1 U926 ( .A1(G122), .A2(n1220), .ZN(n1248) );
XOR2_X1 U927 ( .A(KEYINPUT51), .B(n1249), .Z(n1247) );
NOR2_X1 U928 ( .A1(G122), .A2(n1220), .ZN(n1249) );
NAND3_X1 U929 ( .A1(n1216), .A2(n1065), .A3(n1228), .ZN(n1220) );
NAND2_X1 U930 ( .A1(n1250), .A2(n1251), .ZN(n1065) );
NAND2_X1 U931 ( .A1(n1067), .A2(n1252), .ZN(n1251) );
INV_X1 U932 ( .A(KEYINPUT28), .ZN(n1252) );
NAND3_X1 U933 ( .A1(n1083), .A2(n1253), .A3(KEYINPUT28), .ZN(n1250) );
NAND2_X1 U934 ( .A1(n1254), .A2(n1255), .ZN(n1216) );
NAND3_X1 U935 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1255) );
INV_X1 U936 ( .A(KEYINPUT2), .ZN(n1258) );
NAND2_X1 U937 ( .A1(KEYINPUT2), .A2(n1064), .ZN(n1254) );
XOR2_X1 U938 ( .A(n1259), .B(n1260), .Z(G21) );
NOR2_X1 U939 ( .A1(KEYINPUT49), .A2(n1261), .ZN(n1260) );
INV_X1 U940 ( .A(G119), .ZN(n1261) );
NOR3_X1 U941 ( .A1(n1262), .A2(n1083), .A3(n1253), .ZN(n1259) );
NAND3_X1 U942 ( .A1(n1263), .A2(n1264), .A3(n1066), .ZN(n1262) );
NAND2_X1 U943 ( .A1(KEYINPUT39), .A2(n1265), .ZN(n1264) );
NAND2_X1 U944 ( .A1(n1266), .A2(n1267), .ZN(n1263) );
INV_X1 U945 ( .A(KEYINPUT39), .ZN(n1267) );
NAND3_X1 U946 ( .A1(n1077), .A2(n1268), .A3(n1057), .ZN(n1266) );
INV_X1 U947 ( .A(n1207), .ZN(n1077) );
XNOR2_X1 U948 ( .A(n1224), .B(n1269), .ZN(G18) );
NAND2_X1 U949 ( .A1(KEYINPUT42), .A2(G116), .ZN(n1269) );
AND3_X1 U950 ( .A1(n1064), .A2(n1067), .A3(n1228), .ZN(n1224) );
NOR2_X1 U951 ( .A1(n1256), .A2(n1270), .ZN(n1064) );
XOR2_X1 U952 ( .A(G113), .B(n1223), .Z(G15) );
AND3_X1 U953 ( .A1(n1067), .A2(n1161), .A3(n1228), .ZN(n1223) );
INV_X1 U954 ( .A(n1265), .ZN(n1228) );
NAND3_X1 U955 ( .A1(n1207), .A2(n1268), .A3(n1057), .ZN(n1265) );
NOR2_X1 U956 ( .A1(n1271), .A2(n1074), .ZN(n1057) );
INV_X1 U957 ( .A(n1075), .ZN(n1271) );
NAND2_X1 U958 ( .A1(n1272), .A2(n1273), .ZN(n1161) );
NAND3_X1 U959 ( .A1(n1270), .A2(n1256), .A3(n1274), .ZN(n1273) );
INV_X1 U960 ( .A(KEYINPUT56), .ZN(n1274) );
INV_X1 U961 ( .A(n1257), .ZN(n1270) );
NAND2_X1 U962 ( .A1(KEYINPUT56), .A2(n1066), .ZN(n1272) );
NOR2_X1 U963 ( .A1(n1087), .A2(n1083), .ZN(n1067) );
INV_X1 U964 ( .A(n1253), .ZN(n1087) );
XOR2_X1 U965 ( .A(G110), .B(n1275), .Z(G12) );
NOR4_X1 U966 ( .A1(KEYINPUT62), .A2(n1238), .A3(n1246), .A4(n1276), .ZN(n1275) );
XOR2_X1 U967 ( .A(KEYINPUT5), .B(n1066), .Z(n1276) );
NOR2_X1 U968 ( .A1(n1256), .A2(n1257), .ZN(n1066) );
XOR2_X1 U969 ( .A(n1150), .B(n1277), .Z(n1257) );
NOR2_X1 U970 ( .A1(n1093), .A2(KEYINPUT4), .ZN(n1277) );
NOR2_X1 U971 ( .A1(n1147), .A2(G902), .ZN(n1093) );
XOR2_X1 U972 ( .A(n1278), .B(n1279), .Z(n1147) );
XOR2_X1 U973 ( .A(G107), .B(n1280), .Z(n1279) );
XOR2_X1 U974 ( .A(G134), .B(G128), .Z(n1280) );
XNOR2_X1 U975 ( .A(n1281), .B(n1282), .ZN(n1278) );
XOR2_X1 U976 ( .A(n1283), .B(n1284), .Z(n1281) );
AND2_X1 U977 ( .A1(n1285), .A2(G217), .ZN(n1284) );
NAND2_X1 U978 ( .A1(n1286), .A2(n1287), .ZN(n1283) );
NAND2_X1 U979 ( .A1(G122), .A2(n1288), .ZN(n1287) );
XOR2_X1 U980 ( .A(KEYINPUT1), .B(n1289), .Z(n1286) );
NOR2_X1 U981 ( .A1(G122), .A2(n1288), .ZN(n1289) );
INV_X1 U982 ( .A(G116), .ZN(n1288) );
INV_X1 U983 ( .A(G478), .ZN(n1150) );
XNOR2_X1 U984 ( .A(n1096), .B(n1290), .ZN(n1256) );
NOR2_X1 U985 ( .A1(KEYINPUT17), .A2(n1097), .ZN(n1290) );
XNOR2_X1 U986 ( .A(G475), .B(KEYINPUT35), .ZN(n1097) );
NAND2_X1 U987 ( .A1(n1230), .A2(n1157), .ZN(n1096) );
NAND3_X1 U988 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n1157) );
OR2_X1 U989 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
NAND2_X1 U990 ( .A1(KEYINPUT24), .A2(n1296), .ZN(n1292) );
NAND2_X1 U991 ( .A1(n1297), .A2(n1295), .ZN(n1296) );
XNOR2_X1 U992 ( .A(n1294), .B(KEYINPUT20), .ZN(n1297) );
NAND2_X1 U993 ( .A1(n1298), .A2(n1299), .ZN(n1291) );
INV_X1 U994 ( .A(KEYINPUT24), .ZN(n1299) );
NAND2_X1 U995 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
OR2_X1 U996 ( .A1(n1294), .A2(KEYINPUT20), .ZN(n1301) );
NAND3_X1 U997 ( .A1(n1294), .A2(n1295), .A3(KEYINPUT20), .ZN(n1300) );
XNOR2_X1 U998 ( .A(G104), .B(n1302), .ZN(n1295) );
XOR2_X1 U999 ( .A(G122), .B(G113), .Z(n1302) );
XNOR2_X1 U1000 ( .A(n1303), .B(n1304), .ZN(n1294) );
XNOR2_X1 U1001 ( .A(G125), .B(n1305), .ZN(n1304) );
NAND3_X1 U1002 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1305) );
OR2_X1 U1003 ( .A1(n1309), .A2(KEYINPUT47), .ZN(n1308) );
NAND3_X1 U1004 ( .A1(KEYINPUT47), .A2(n1310), .A3(n1117), .ZN(n1307) );
INV_X1 U1005 ( .A(n1311), .ZN(n1310) );
NAND2_X1 U1006 ( .A1(G131), .A2(n1311), .ZN(n1306) );
NAND2_X1 U1007 ( .A1(KEYINPUT44), .A2(n1309), .ZN(n1311) );
XOR2_X1 U1008 ( .A(n1312), .B(n1282), .Z(n1309) );
NAND3_X1 U1009 ( .A1(n1313), .A2(n1152), .A3(G214), .ZN(n1312) );
XOR2_X1 U1010 ( .A(G146), .B(n1314), .Z(n1303) );
NAND2_X1 U1011 ( .A1(n1315), .A2(n1316), .ZN(n1246) );
XOR2_X1 U1012 ( .A(KEYINPUT28), .B(n1229), .Z(n1316) );
INV_X1 U1013 ( .A(n1083), .ZN(n1229) );
XOR2_X1 U1014 ( .A(n1317), .B(G472), .Z(n1083) );
NAND2_X1 U1015 ( .A1(n1318), .A2(n1230), .ZN(n1317) );
XOR2_X1 U1016 ( .A(n1319), .B(n1320), .Z(n1318) );
XOR2_X1 U1017 ( .A(G101), .B(n1321), .Z(n1320) );
NOR2_X1 U1018 ( .A1(n1165), .A2(KEYINPUT31), .ZN(n1321) );
AND3_X1 U1019 ( .A1(n1313), .A2(n1152), .A3(G210), .ZN(n1165) );
NAND2_X1 U1020 ( .A1(KEYINPUT53), .A2(n1170), .ZN(n1319) );
XOR2_X1 U1021 ( .A(n1322), .B(n1113), .Z(n1170) );
XNOR2_X1 U1022 ( .A(n1180), .B(n1323), .ZN(n1322) );
XOR2_X1 U1023 ( .A(n1253), .B(KEYINPUT33), .Z(n1315) );
XOR2_X1 U1024 ( .A(n1324), .B(n1144), .Z(n1253) );
AND2_X1 U1025 ( .A1(G217), .A2(n1325), .ZN(n1144) );
NAND2_X1 U1026 ( .A1(n1142), .A2(n1230), .ZN(n1324) );
XOR2_X1 U1027 ( .A(n1326), .B(n1327), .Z(n1142) );
XOR2_X1 U1028 ( .A(n1328), .B(n1329), .Z(n1327) );
XOR2_X1 U1029 ( .A(G119), .B(G110), .Z(n1329) );
XOR2_X1 U1030 ( .A(G137), .B(G125), .Z(n1328) );
XNOR2_X1 U1031 ( .A(n1330), .B(n1331), .ZN(n1326) );
XOR2_X1 U1032 ( .A(n1332), .B(n1333), .Z(n1331) );
NAND2_X1 U1033 ( .A1(n1285), .A2(G221), .ZN(n1333) );
AND2_X1 U1034 ( .A1(G234), .A2(n1152), .ZN(n1285) );
NAND2_X1 U1035 ( .A1(KEYINPUT18), .A2(n1314), .ZN(n1332) );
INV_X1 U1036 ( .A(G140), .ZN(n1314) );
NAND3_X1 U1037 ( .A1(n1237), .A2(n1268), .A3(n1207), .ZN(n1238) );
NOR2_X1 U1038 ( .A1(n1080), .A2(n1079), .ZN(n1207) );
AND2_X1 U1039 ( .A1(G214), .A2(n1334), .ZN(n1079) );
XOR2_X1 U1040 ( .A(n1098), .B(n1335), .Z(n1080) );
NOR2_X1 U1041 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
AND2_X1 U1042 ( .A1(KEYINPUT29), .A2(n1099), .ZN(n1337) );
NOR2_X1 U1043 ( .A1(KEYINPUT16), .A2(n1099), .ZN(n1336) );
NAND2_X1 U1044 ( .A1(G210), .A2(n1334), .ZN(n1099) );
NAND2_X1 U1045 ( .A1(n1230), .A2(n1313), .ZN(n1334) );
INV_X1 U1046 ( .A(G237), .ZN(n1313) );
NAND2_X1 U1047 ( .A1(n1338), .A2(n1230), .ZN(n1098) );
XOR2_X1 U1048 ( .A(n1191), .B(n1339), .Z(n1338) );
XOR2_X1 U1049 ( .A(n1187), .B(n1340), .Z(n1339) );
NOR2_X1 U1050 ( .A1(KEYINPUT0), .A2(n1192), .ZN(n1340) );
NAND2_X1 U1051 ( .A1(G224), .A2(n1152), .ZN(n1192) );
NAND3_X1 U1052 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1187) );
OR2_X1 U1053 ( .A1(n1135), .A2(KEYINPUT23), .ZN(n1343) );
OR2_X1 U1054 ( .A1(n1138), .A2(n1137), .ZN(n1135) );
OR2_X1 U1055 ( .A1(n1344), .A2(n1345), .ZN(n1138) );
AND2_X1 U1056 ( .A1(n1323), .A2(n1346), .ZN(n1345) );
NAND3_X1 U1057 ( .A1(n1344), .A2(KEYINPUT23), .A3(n1347), .ZN(n1342) );
NAND2_X1 U1058 ( .A1(n1137), .A2(n1348), .ZN(n1341) );
NAND2_X1 U1059 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1060 ( .A1(n1323), .A2(n1346), .ZN(n1350) );
XNOR2_X1 U1061 ( .A(KEYINPUT23), .B(n1344), .ZN(n1349) );
NOR2_X1 U1062 ( .A1(n1346), .A2(n1323), .ZN(n1344) );
XOR2_X1 U1063 ( .A(n1351), .B(n1352), .Z(n1323) );
XOR2_X1 U1064 ( .A(G119), .B(G116), .Z(n1352) );
INV_X1 U1065 ( .A(G113), .ZN(n1351) );
NAND2_X1 U1066 ( .A1(n1353), .A2(n1354), .ZN(n1346) );
NAND2_X1 U1067 ( .A1(G101), .A2(n1355), .ZN(n1354) );
XOR2_X1 U1068 ( .A(n1356), .B(KEYINPUT10), .Z(n1353) );
OR2_X1 U1069 ( .A1(n1355), .A2(G101), .ZN(n1356) );
INV_X1 U1070 ( .A(n1347), .ZN(n1137) );
XOR2_X1 U1071 ( .A(n1357), .B(G122), .Z(n1347) );
INV_X1 U1072 ( .A(G110), .ZN(n1357) );
XOR2_X1 U1073 ( .A(n1358), .B(n1113), .Z(n1191) );
XNOR2_X1 U1074 ( .A(G125), .B(KEYINPUT3), .ZN(n1358) );
NAND2_X1 U1075 ( .A1(n1359), .A2(n1081), .ZN(n1268) );
NAND3_X1 U1076 ( .A1(n1360), .A2(n1152), .A3(G952), .ZN(n1081) );
NAND3_X1 U1077 ( .A1(n1244), .A2(n1133), .A3(G953), .ZN(n1359) );
INV_X1 U1078 ( .A(G898), .ZN(n1133) );
AND2_X1 U1079 ( .A1(G902), .A2(n1360), .ZN(n1244) );
NAND2_X1 U1080 ( .A1(G237), .A2(G234), .ZN(n1360) );
NOR2_X1 U1081 ( .A1(n1075), .A2(n1074), .ZN(n1237) );
AND2_X1 U1082 ( .A1(G221), .A2(n1325), .ZN(n1074) );
NAND2_X1 U1083 ( .A1(G234), .A2(n1230), .ZN(n1325) );
XOR2_X1 U1084 ( .A(n1361), .B(G469), .Z(n1075) );
NAND2_X1 U1085 ( .A1(n1362), .A2(n1230), .ZN(n1361) );
INV_X1 U1086 ( .A(G902), .ZN(n1230) );
XOR2_X1 U1087 ( .A(n1363), .B(n1364), .Z(n1362) );
XOR2_X1 U1088 ( .A(n1365), .B(n1183), .Z(n1364) );
AND2_X1 U1089 ( .A1(G227), .A2(n1152), .ZN(n1183) );
INV_X1 U1090 ( .A(G953), .ZN(n1152) );
NAND2_X1 U1091 ( .A1(n1366), .A2(n1367), .ZN(n1365) );
NAND2_X1 U1092 ( .A1(n1177), .A2(n1180), .ZN(n1367) );
XOR2_X1 U1093 ( .A(KEYINPUT12), .B(n1368), .Z(n1366) );
NOR2_X1 U1094 ( .A1(n1177), .A2(n1180), .ZN(n1368) );
NAND3_X1 U1095 ( .A1(n1369), .A2(n1370), .A3(n1371), .ZN(n1180) );
NAND2_X1 U1096 ( .A1(G131), .A2(n1372), .ZN(n1371) );
NAND2_X1 U1097 ( .A1(n1373), .A2(n1374), .ZN(n1370) );
INV_X1 U1098 ( .A(KEYINPUT13), .ZN(n1374) );
NAND2_X1 U1099 ( .A1(n1375), .A2(n1117), .ZN(n1373) );
INV_X1 U1100 ( .A(G131), .ZN(n1117) );
XOR2_X1 U1101 ( .A(KEYINPUT38), .B(n1372), .Z(n1375) );
NAND2_X1 U1102 ( .A1(KEYINPUT13), .A2(n1376), .ZN(n1369) );
NAND2_X1 U1103 ( .A1(n1377), .A2(n1378), .ZN(n1376) );
NAND2_X1 U1104 ( .A1(n1372), .A2(n1379), .ZN(n1378) );
OR3_X1 U1105 ( .A1(n1372), .A2(G131), .A3(n1379), .ZN(n1377) );
INV_X1 U1106 ( .A(KEYINPUT38), .ZN(n1379) );
XOR2_X1 U1107 ( .A(n1114), .B(KEYINPUT9), .Z(n1372) );
XOR2_X1 U1108 ( .A(G134), .B(G137), .Z(n1114) );
XOR2_X1 U1109 ( .A(n1380), .B(n1381), .Z(n1177) );
XOR2_X1 U1110 ( .A(KEYINPUT11), .B(G101), .Z(n1381) );
XNOR2_X1 U1111 ( .A(n1355), .B(n1113), .ZN(n1380) );
XNOR2_X1 U1112 ( .A(n1282), .B(n1330), .ZN(n1113) );
XOR2_X1 U1113 ( .A(G128), .B(G146), .Z(n1330) );
XNOR2_X1 U1114 ( .A(G143), .B(KEYINPUT48), .ZN(n1282) );
XOR2_X1 U1115 ( .A(G104), .B(G107), .Z(n1355) );
NAND2_X1 U1116 ( .A1(KEYINPUT34), .A2(n1178), .ZN(n1363) );
XOR2_X1 U1117 ( .A(G110), .B(G140), .Z(n1178) );
endmodule


