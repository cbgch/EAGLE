//Key = 0001001101101000101010101000111010001010001100111111100010100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398;

XOR2_X1 U756 ( .A(G107), .B(n1058), .Z(G9) );
NOR2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(G75) );
NOR4_X1 U758 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1060) );
NAND3_X1 U759 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U761 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U762 ( .A1(KEYINPUT23), .A2(n1072), .ZN(n1071) );
NAND2_X1 U763 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U764 ( .A1(n1075), .A2(n1076), .ZN(n1070) );
NAND2_X1 U765 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND4_X1 U766 ( .A1(n1079), .A2(n1080), .A3(n1074), .A4(n1081), .ZN(n1078) );
INV_X1 U767 ( .A(KEYINPUT23), .ZN(n1081) );
NAND3_X1 U768 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1077) );
NAND2_X1 U769 ( .A1(n1085), .A2(n1086), .ZN(n1082) );
NAND2_X1 U770 ( .A1(n1080), .A2(n1087), .ZN(n1086) );
NAND2_X1 U771 ( .A1(n1079), .A2(n1088), .ZN(n1085) );
NAND2_X1 U772 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND4_X1 U773 ( .A1(n1084), .A2(n1073), .A3(n1091), .A4(n1092), .ZN(n1065) );
NAND2_X1 U774 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND3_X1 U775 ( .A1(n1095), .A2(n1096), .A3(n1083), .ZN(n1091) );
NAND2_X1 U776 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
INV_X1 U777 ( .A(n1099), .ZN(n1097) );
AND3_X1 U778 ( .A1(n1080), .A2(n1075), .A3(n1079), .ZN(n1073) );
XNOR2_X1 U779 ( .A(KEYINPUT30), .B(n1100), .ZN(n1075) );
NOR3_X1 U780 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1059) );
NOR2_X1 U781 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
INV_X1 U782 ( .A(KEYINPUT56), .ZN(n1105) );
NOR2_X1 U783 ( .A1(G953), .A2(G952), .ZN(n1104) );
NOR2_X1 U784 ( .A1(KEYINPUT56), .A2(n1106), .ZN(n1102) );
INV_X1 U785 ( .A(n1066), .ZN(n1101) );
NAND4_X1 U786 ( .A1(n1107), .A2(n1108), .A3(n1109), .A4(n1110), .ZN(n1066) );
NOR3_X1 U787 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1110) );
NAND3_X1 U788 ( .A1(n1099), .A2(n1083), .A3(n1114), .ZN(n1111) );
NAND2_X1 U789 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR3_X1 U790 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1109) );
NOR2_X1 U791 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U792 ( .A1(G475), .A2(n1122), .ZN(n1118) );
NOR2_X1 U793 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
AND2_X1 U794 ( .A1(n1121), .A2(KEYINPUT61), .ZN(n1124) );
OR2_X1 U795 ( .A1(n1125), .A2(KEYINPUT45), .ZN(n1121) );
NOR2_X1 U796 ( .A1(KEYINPUT61), .A2(n1125), .ZN(n1123) );
XOR2_X1 U797 ( .A(KEYINPUT2), .B(n1126), .Z(n1117) );
XOR2_X1 U798 ( .A(n1127), .B(G469), .Z(n1108) );
NAND2_X1 U799 ( .A1(KEYINPUT51), .A2(n1128), .ZN(n1127) );
XOR2_X1 U800 ( .A(n1129), .B(KEYINPUT19), .Z(n1107) );
OR2_X1 U801 ( .A1(n1116), .A2(n1115), .ZN(n1129) );
XOR2_X1 U802 ( .A(n1130), .B(n1131), .Z(G72) );
XOR2_X1 U803 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U804 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND2_X1 U805 ( .A1(G900), .A2(G227), .ZN(n1135) );
XOR2_X1 U806 ( .A(KEYINPUT4), .B(G953), .Z(n1134) );
NAND2_X1 U807 ( .A1(n1136), .A2(n1062), .ZN(n1132) );
XOR2_X1 U808 ( .A(n1137), .B(KEYINPUT17), .Z(n1136) );
NOR3_X1 U809 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1130) );
NOR2_X1 U810 ( .A1(G900), .A2(n1137), .ZN(n1140) );
NOR2_X1 U811 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
NAND3_X1 U812 ( .A1(n1143), .A2(n1144), .A3(KEYINPUT48), .ZN(n1138) );
NAND2_X1 U813 ( .A1(KEYINPUT27), .A2(n1145), .ZN(n1144) );
NAND2_X1 U814 ( .A1(n1146), .A2(n1142), .ZN(n1145) );
XNOR2_X1 U815 ( .A(KEYINPUT10), .B(n1141), .ZN(n1146) );
NAND2_X1 U816 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
INV_X1 U817 ( .A(KEYINPUT27), .ZN(n1148) );
NAND2_X1 U818 ( .A1(n1149), .A2(n1150), .ZN(n1147) );
OR2_X1 U819 ( .A1(n1141), .A2(KEYINPUT10), .ZN(n1150) );
NAND3_X1 U820 ( .A1(n1142), .A2(n1141), .A3(KEYINPUT10), .ZN(n1149) );
XNOR2_X1 U821 ( .A(n1151), .B(n1152), .ZN(n1142) );
XOR2_X1 U822 ( .A(G137), .B(G131), .Z(n1152) );
XOR2_X1 U823 ( .A(n1153), .B(n1154), .Z(n1151) );
NOR2_X1 U824 ( .A1(G134), .A2(KEYINPUT26), .ZN(n1154) );
NAND2_X1 U825 ( .A1(n1155), .A2(n1156), .ZN(G69) );
NAND2_X1 U826 ( .A1(n1157), .A2(n1137), .ZN(n1156) );
XNOR2_X1 U827 ( .A(n1158), .B(n1064), .ZN(n1157) );
NAND2_X1 U828 ( .A1(n1159), .A2(G953), .ZN(n1155) );
NAND2_X1 U829 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U830 ( .A1(n1158), .A2(n1162), .ZN(n1161) );
INV_X1 U831 ( .A(G224), .ZN(n1162) );
NAND2_X1 U832 ( .A1(G224), .A2(n1163), .ZN(n1160) );
NAND2_X1 U833 ( .A1(G898), .A2(n1158), .ZN(n1163) );
NAND2_X1 U834 ( .A1(n1164), .A2(n1165), .ZN(n1158) );
NAND2_X1 U835 ( .A1(G953), .A2(n1166), .ZN(n1165) );
XOR2_X1 U836 ( .A(n1167), .B(n1168), .Z(n1164) );
NOR2_X1 U837 ( .A1(KEYINPUT34), .A2(n1169), .ZN(n1168) );
NOR2_X1 U838 ( .A1(n1106), .A2(n1170), .ZN(G66) );
XNOR2_X1 U839 ( .A(n1171), .B(n1172), .ZN(n1170) );
NOR2_X1 U840 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NOR2_X1 U841 ( .A1(n1106), .A2(n1175), .ZN(G63) );
XOR2_X1 U842 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR3_X1 U843 ( .A1(n1174), .A2(KEYINPUT40), .A3(n1178), .ZN(n1176) );
INV_X1 U844 ( .A(G478), .ZN(n1178) );
NOR2_X1 U845 ( .A1(n1106), .A2(n1179), .ZN(G60) );
NOR3_X1 U846 ( .A1(n1125), .A2(n1180), .A3(n1181), .ZN(n1179) );
NOR3_X1 U847 ( .A1(n1182), .A2(n1120), .A3(n1174), .ZN(n1181) );
NOR2_X1 U848 ( .A1(n1183), .A2(n1184), .ZN(n1180) );
NOR2_X1 U849 ( .A1(n1185), .A2(n1120), .ZN(n1183) );
NOR2_X1 U850 ( .A1(n1064), .A2(n1062), .ZN(n1185) );
XOR2_X1 U851 ( .A(G104), .B(n1186), .Z(G6) );
NOR2_X1 U852 ( .A1(n1096), .A2(n1187), .ZN(n1186) );
NOR2_X1 U853 ( .A1(n1106), .A2(n1188), .ZN(G57) );
NOR2_X1 U854 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U855 ( .A(KEYINPUT54), .B(n1191), .Z(n1190) );
NOR2_X1 U856 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XNOR2_X1 U857 ( .A(KEYINPUT42), .B(n1194), .ZN(n1193) );
NOR2_X1 U858 ( .A1(n1195), .A2(n1196), .ZN(n1189) );
INV_X1 U859 ( .A(n1192), .ZN(n1196) );
XOR2_X1 U860 ( .A(n1197), .B(n1198), .Z(n1192) );
NOR2_X1 U861 ( .A1(n1199), .A2(n1174), .ZN(n1198) );
INV_X1 U862 ( .A(G472), .ZN(n1199) );
XOR2_X1 U863 ( .A(n1194), .B(KEYINPUT42), .Z(n1195) );
XOR2_X1 U864 ( .A(n1200), .B(G101), .Z(n1194) );
NOR2_X1 U865 ( .A1(n1106), .A2(n1201), .ZN(G54) );
XOR2_X1 U866 ( .A(n1202), .B(n1203), .Z(n1201) );
XOR2_X1 U867 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U868 ( .A(KEYINPUT11), .B(n1206), .Z(n1205) );
NOR2_X1 U869 ( .A1(n1207), .A2(n1174), .ZN(n1204) );
INV_X1 U870 ( .A(G469), .ZN(n1207) );
XNOR2_X1 U871 ( .A(n1208), .B(n1209), .ZN(n1202) );
XNOR2_X1 U872 ( .A(n1210), .B(n1211), .ZN(n1209) );
NAND2_X1 U873 ( .A1(KEYINPUT36), .A2(n1212), .ZN(n1210) );
NOR2_X1 U874 ( .A1(n1106), .A2(n1213), .ZN(G51) );
XOR2_X1 U875 ( .A(n1214), .B(n1215), .Z(n1213) );
NOR2_X1 U876 ( .A1(n1116), .A2(n1174), .ZN(n1215) );
NAND2_X1 U877 ( .A1(G902), .A2(n1216), .ZN(n1174) );
OR2_X1 U878 ( .A1(n1062), .A2(n1064), .ZN(n1216) );
NAND2_X1 U879 ( .A1(n1217), .A2(n1218), .ZN(n1064) );
NOR4_X1 U880 ( .A1(n1219), .A2(n1220), .A3(n1058), .A4(n1221), .ZN(n1218) );
AND4_X1 U881 ( .A1(n1080), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1058) );
NOR2_X1 U882 ( .A1(KEYINPUT55), .A2(n1225), .ZN(n1220) );
NOR2_X1 U883 ( .A1(n1226), .A2(n1096), .ZN(n1219) );
XOR2_X1 U884 ( .A(n1187), .B(KEYINPUT59), .Z(n1226) );
NAND3_X1 U885 ( .A1(n1080), .A2(n1223), .A3(n1227), .ZN(n1187) );
NOR4_X1 U886 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1217) );
NOR3_X1 U887 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1231) );
NOR2_X1 U888 ( .A1(n1096), .A2(n1235), .ZN(n1234) );
NOR2_X1 U889 ( .A1(n1224), .A2(n1236), .ZN(n1233) );
AND2_X1 U890 ( .A1(n1237), .A2(KEYINPUT55), .ZN(n1236) );
INV_X1 U891 ( .A(n1238), .ZN(n1230) );
NAND4_X1 U892 ( .A1(n1239), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1062) );
NOR4_X1 U893 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1242) );
NAND3_X1 U894 ( .A1(n1247), .A2(n1087), .A3(n1248), .ZN(n1241) );
NAND2_X1 U895 ( .A1(n1249), .A2(n1250), .ZN(n1087) );
NAND3_X1 U896 ( .A1(n1247), .A2(n1068), .A3(n1251), .ZN(n1239) );
NAND4_X1 U897 ( .A1(KEYINPUT28), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1214) );
OR3_X1 U898 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1254) );
NAND2_X1 U899 ( .A1(n1258), .A2(n1257), .ZN(n1253) );
XOR2_X1 U900 ( .A(n1255), .B(n1256), .Z(n1258) );
NAND2_X1 U901 ( .A1(n1259), .A2(n1255), .ZN(n1252) );
NOR2_X1 U902 ( .A1(n1137), .A2(G952), .ZN(n1106) );
XOR2_X1 U903 ( .A(G146), .B(n1260), .Z(G48) );
NOR3_X1 U904 ( .A1(n1261), .A2(n1262), .A3(n1249), .ZN(n1260) );
XOR2_X1 U905 ( .A(n1096), .B(KEYINPUT25), .Z(n1262) );
XNOR2_X1 U906 ( .A(n1240), .B(n1263), .ZN(G45) );
NOR2_X1 U907 ( .A1(KEYINPUT44), .A2(n1264), .ZN(n1263) );
NAND3_X1 U908 ( .A1(n1237), .A2(n1247), .A3(n1265), .ZN(n1240) );
NOR3_X1 U909 ( .A1(n1096), .A2(n1266), .A3(n1267), .ZN(n1265) );
XOR2_X1 U910 ( .A(n1245), .B(n1268), .Z(G42) );
NOR2_X1 U911 ( .A1(KEYINPUT62), .A2(n1269), .ZN(n1268) );
XNOR2_X1 U912 ( .A(G140), .B(KEYINPUT39), .ZN(n1269) );
AND2_X1 U913 ( .A1(n1270), .A2(n1235), .ZN(n1245) );
XOR2_X1 U914 ( .A(G137), .B(n1244), .Z(G39) );
NOR3_X1 U915 ( .A1(n1271), .A2(n1094), .A3(n1261), .ZN(n1244) );
NAND3_X1 U916 ( .A1(n1247), .A2(n1126), .A3(n1272), .ZN(n1261) );
XNOR2_X1 U917 ( .A(G134), .B(n1273), .ZN(G36) );
NAND3_X1 U918 ( .A1(n1251), .A2(n1247), .A3(n1274), .ZN(n1273) );
XOR2_X1 U919 ( .A(n1094), .B(KEYINPUT6), .Z(n1274) );
XNOR2_X1 U920 ( .A(n1243), .B(n1275), .ZN(G33) );
NAND2_X1 U921 ( .A1(KEYINPUT16), .A2(G131), .ZN(n1275) );
AND2_X1 U922 ( .A1(n1237), .A2(n1270), .ZN(n1243) );
AND3_X1 U923 ( .A1(n1068), .A2(n1227), .A3(n1247), .ZN(n1270) );
AND2_X1 U924 ( .A1(n1074), .A2(n1276), .ZN(n1247) );
INV_X1 U925 ( .A(n1094), .ZN(n1068) );
NAND2_X1 U926 ( .A1(n1098), .A2(n1099), .ZN(n1094) );
XOR2_X1 U927 ( .A(n1277), .B(n1278), .Z(G30) );
XOR2_X1 U928 ( .A(KEYINPUT3), .B(G128), .Z(n1278) );
NAND4_X1 U929 ( .A1(n1279), .A2(n1248), .A3(n1222), .A4(n1276), .ZN(n1277) );
INV_X1 U930 ( .A(n1250), .ZN(n1222) );
NOR3_X1 U931 ( .A1(n1096), .A2(n1280), .A3(n1281), .ZN(n1248) );
XNOR2_X1 U932 ( .A(n1074), .B(KEYINPUT52), .ZN(n1279) );
XOR2_X1 U933 ( .A(n1282), .B(n1225), .Z(G3) );
OR3_X1 U934 ( .A1(n1090), .A2(n1096), .A3(n1232), .ZN(n1225) );
XOR2_X1 U935 ( .A(G125), .B(n1246), .Z(G27) );
AND4_X1 U936 ( .A1(n1276), .A2(n1083), .A3(n1235), .A4(n1283), .ZN(n1246) );
AND3_X1 U937 ( .A1(n1084), .A2(n1224), .A3(n1227), .ZN(n1283) );
NAND2_X1 U938 ( .A1(n1284), .A2(n1285), .ZN(n1276) );
NAND2_X1 U939 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
INV_X1 U940 ( .A(G900), .ZN(n1287) );
XOR2_X1 U941 ( .A(n1288), .B(n1238), .Z(G24) );
NAND4_X1 U942 ( .A1(n1289), .A2(n1080), .A3(n1290), .A4(n1291), .ZN(n1238) );
XOR2_X1 U943 ( .A(G119), .B(n1229), .Z(G21) );
AND4_X1 U944 ( .A1(n1289), .A2(n1079), .A3(n1272), .A4(n1126), .ZN(n1229) );
XOR2_X1 U945 ( .A(n1228), .B(n1292), .Z(G18) );
NOR2_X1 U946 ( .A1(KEYINPUT37), .A2(n1293), .ZN(n1292) );
INV_X1 U947 ( .A(G116), .ZN(n1293) );
AND2_X1 U948 ( .A1(n1289), .A2(n1251), .ZN(n1228) );
NOR2_X1 U949 ( .A1(n1090), .A2(n1250), .ZN(n1251) );
NAND2_X1 U950 ( .A1(n1266), .A2(n1290), .ZN(n1250) );
INV_X1 U951 ( .A(n1267), .ZN(n1290) );
XOR2_X1 U952 ( .A(G113), .B(n1221), .Z(G15) );
AND3_X1 U953 ( .A1(n1237), .A2(n1227), .A3(n1289), .ZN(n1221) );
AND4_X1 U954 ( .A1(n1084), .A2(n1224), .A3(n1294), .A4(n1083), .ZN(n1289) );
INV_X1 U955 ( .A(n1096), .ZN(n1224) );
INV_X1 U956 ( .A(n1249), .ZN(n1227) );
NAND2_X1 U957 ( .A1(n1267), .A2(n1291), .ZN(n1249) );
INV_X1 U958 ( .A(n1090), .ZN(n1237) );
NAND2_X1 U959 ( .A1(n1126), .A2(n1281), .ZN(n1090) );
XOR2_X1 U960 ( .A(G110), .B(n1295), .Z(G12) );
NOR3_X1 U961 ( .A1(n1232), .A2(n1089), .A3(n1296), .ZN(n1295) );
XOR2_X1 U962 ( .A(n1096), .B(KEYINPUT57), .Z(n1296) );
NAND2_X1 U963 ( .A1(n1297), .A2(n1099), .ZN(n1096) );
NAND2_X1 U964 ( .A1(G214), .A2(n1298), .ZN(n1099) );
INV_X1 U965 ( .A(n1098), .ZN(n1297) );
XOR2_X1 U966 ( .A(n1115), .B(n1116), .Z(n1098) );
NAND2_X1 U967 ( .A1(G210), .A2(n1298), .ZN(n1116) );
NAND2_X1 U968 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
INV_X1 U969 ( .A(G237), .ZN(n1299) );
AND2_X1 U970 ( .A1(n1301), .A2(n1300), .ZN(n1115) );
XOR2_X1 U971 ( .A(n1302), .B(n1303), .Z(n1301) );
INV_X1 U972 ( .A(n1255), .ZN(n1303) );
XOR2_X1 U973 ( .A(n1167), .B(n1169), .Z(n1255) );
XNOR2_X1 U974 ( .A(n1304), .B(G110), .ZN(n1169) );
NAND2_X1 U975 ( .A1(KEYINPUT58), .A2(G122), .ZN(n1304) );
XOR2_X1 U976 ( .A(n1305), .B(n1306), .Z(n1167) );
XOR2_X1 U977 ( .A(n1307), .B(n1308), .Z(n1305) );
NOR2_X1 U978 ( .A1(KEYINPUT31), .A2(n1309), .ZN(n1308) );
NOR2_X1 U979 ( .A1(n1259), .A2(n1310), .ZN(n1302) );
NOR2_X1 U980 ( .A1(n1311), .A2(n1256), .ZN(n1310) );
INV_X1 U981 ( .A(n1312), .ZN(n1256) );
XOR2_X1 U982 ( .A(n1257), .B(KEYINPUT43), .Z(n1311) );
NOR2_X1 U983 ( .A1(n1257), .A2(n1312), .ZN(n1259) );
XNOR2_X1 U984 ( .A(n1313), .B(n1314), .ZN(n1312) );
XOR2_X1 U985 ( .A(KEYINPUT18), .B(G125), .Z(n1314) );
NAND2_X1 U986 ( .A1(G224), .A2(n1137), .ZN(n1257) );
INV_X1 U987 ( .A(n1235), .ZN(n1089) );
NAND2_X1 U988 ( .A1(n1315), .A2(n1316), .ZN(n1235) );
OR3_X1 U989 ( .A1(n1126), .A2(n1281), .A3(KEYINPUT14), .ZN(n1316) );
INV_X1 U990 ( .A(n1272), .ZN(n1281) );
NAND2_X1 U991 ( .A1(KEYINPUT14), .A2(n1080), .ZN(n1315) );
NOR2_X1 U992 ( .A1(n1126), .A2(n1272), .ZN(n1080) );
XNOR2_X1 U993 ( .A(n1113), .B(KEYINPUT7), .ZN(n1272) );
XOR2_X1 U994 ( .A(n1317), .B(n1173), .Z(n1113) );
NAND2_X1 U995 ( .A1(G217), .A2(n1318), .ZN(n1173) );
NAND2_X1 U996 ( .A1(n1171), .A2(n1300), .ZN(n1317) );
XNOR2_X1 U997 ( .A(n1319), .B(n1320), .ZN(n1171) );
XOR2_X1 U998 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U999 ( .A(G137), .B(G119), .Z(n1322) );
XOR2_X1 U1000 ( .A(KEYINPUT49), .B(KEYINPUT15), .Z(n1321) );
XOR2_X1 U1001 ( .A(n1323), .B(n1324), .Z(n1319) );
XNOR2_X1 U1002 ( .A(G110), .B(n1325), .ZN(n1324) );
NAND2_X1 U1003 ( .A1(G221), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1004 ( .A(n1327), .B(n1328), .Z(n1323) );
NAND2_X1 U1005 ( .A1(KEYINPUT9), .A2(n1329), .ZN(n1327) );
XOR2_X1 U1006 ( .A(KEYINPUT32), .B(G128), .Z(n1329) );
INV_X1 U1007 ( .A(n1280), .ZN(n1126) );
XOR2_X1 U1008 ( .A(n1330), .B(G472), .Z(n1280) );
NAND2_X1 U1009 ( .A1(n1331), .A2(n1300), .ZN(n1330) );
XOR2_X1 U1010 ( .A(n1197), .B(n1332), .Z(n1331) );
XOR2_X1 U1011 ( .A(n1333), .B(KEYINPUT29), .Z(n1332) );
NAND2_X1 U1012 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
OR2_X1 U1013 ( .A1(n1282), .A2(n1200), .ZN(n1335) );
XOR2_X1 U1014 ( .A(n1336), .B(KEYINPUT41), .Z(n1334) );
NAND2_X1 U1015 ( .A1(n1282), .A2(n1200), .ZN(n1336) );
NAND2_X1 U1016 ( .A1(G210), .A2(n1337), .ZN(n1200) );
XOR2_X1 U1017 ( .A(n1338), .B(n1339), .Z(n1197) );
XOR2_X1 U1018 ( .A(KEYINPUT33), .B(n1306), .Z(n1339) );
XOR2_X1 U1019 ( .A(G113), .B(n1340), .Z(n1306) );
XOR2_X1 U1020 ( .A(G119), .B(G116), .Z(n1340) );
XNOR2_X1 U1021 ( .A(n1341), .B(n1313), .ZN(n1338) );
XOR2_X1 U1022 ( .A(G128), .B(n1342), .Z(n1313) );
XOR2_X1 U1023 ( .A(G146), .B(G143), .Z(n1342) );
NAND2_X1 U1024 ( .A1(n1079), .A2(n1223), .ZN(n1232) );
AND2_X1 U1025 ( .A1(n1074), .A2(n1294), .ZN(n1223) );
NAND2_X1 U1026 ( .A1(n1284), .A2(n1343), .ZN(n1294) );
NAND2_X1 U1027 ( .A1(n1286), .A2(n1166), .ZN(n1343) );
INV_X1 U1028 ( .A(G898), .ZN(n1166) );
AND3_X1 U1029 ( .A1(G902), .A2(n1100), .A3(G953), .ZN(n1286) );
NAND2_X1 U1030 ( .A1(n1344), .A2(n1100), .ZN(n1284) );
NAND2_X1 U1031 ( .A1(G237), .A2(G234), .ZN(n1100) );
INV_X1 U1032 ( .A(n1063), .ZN(n1344) );
NAND2_X1 U1033 ( .A1(G952), .A2(n1345), .ZN(n1063) );
XOR2_X1 U1034 ( .A(KEYINPUT56), .B(G953), .Z(n1345) );
NOR2_X1 U1035 ( .A1(n1084), .A2(n1093), .ZN(n1074) );
INV_X1 U1036 ( .A(n1083), .ZN(n1093) );
NAND2_X1 U1037 ( .A1(G221), .A2(n1318), .ZN(n1083) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1300), .ZN(n1318) );
XNOR2_X1 U1039 ( .A(n1128), .B(G469), .ZN(n1084) );
AND2_X1 U1040 ( .A1(n1346), .A2(n1300), .ZN(n1128) );
INV_X1 U1041 ( .A(G902), .ZN(n1300) );
XOR2_X1 U1042 ( .A(n1347), .B(n1348), .Z(n1346) );
XNOR2_X1 U1043 ( .A(n1212), .B(n1208), .ZN(n1348) );
XNOR2_X1 U1044 ( .A(n1153), .B(n1341), .ZN(n1208) );
XNOR2_X1 U1045 ( .A(n1349), .B(n1350), .ZN(n1341) );
XOR2_X1 U1046 ( .A(KEYINPUT0), .B(G134), .Z(n1350) );
XOR2_X1 U1047 ( .A(n1351), .B(G131), .Z(n1349) );
NAND2_X1 U1048 ( .A1(KEYINPUT22), .A2(n1352), .ZN(n1351) );
INV_X1 U1049 ( .A(G137), .ZN(n1352) );
NAND2_X1 U1050 ( .A1(n1353), .A2(n1354), .ZN(n1153) );
NAND2_X1 U1051 ( .A1(G128), .A2(n1355), .ZN(n1354) );
XOR2_X1 U1052 ( .A(n1356), .B(KEYINPUT8), .Z(n1353) );
OR2_X1 U1053 ( .A1(n1355), .A2(G128), .ZN(n1356) );
NAND2_X1 U1054 ( .A1(n1357), .A2(n1358), .ZN(n1355) );
NAND2_X1 U1055 ( .A1(G143), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1056 ( .A(n1360), .B(KEYINPUT21), .Z(n1357) );
NAND2_X1 U1057 ( .A1(G146), .A2(n1264), .ZN(n1360) );
XNOR2_X1 U1058 ( .A(n1361), .B(n1309), .ZN(n1212) );
XOR2_X1 U1059 ( .A(n1307), .B(KEYINPUT47), .Z(n1361) );
XOR2_X1 U1060 ( .A(n1282), .B(n1362), .Z(n1307) );
XOR2_X1 U1061 ( .A(KEYINPUT13), .B(G104), .Z(n1362) );
INV_X1 U1062 ( .A(G101), .ZN(n1282) );
XOR2_X1 U1063 ( .A(n1363), .B(n1364), .Z(n1347) );
XOR2_X1 U1064 ( .A(KEYINPUT63), .B(n1206), .Z(n1364) );
AND2_X1 U1065 ( .A1(n1365), .A2(n1137), .ZN(n1206) );
XNOR2_X1 U1066 ( .A(G227), .B(KEYINPUT50), .ZN(n1365) );
NAND2_X1 U1067 ( .A1(KEYINPUT12), .A2(n1211), .ZN(n1363) );
XOR2_X1 U1068 ( .A(G140), .B(G110), .Z(n1211) );
INV_X1 U1069 ( .A(n1271), .ZN(n1079) );
NAND2_X1 U1070 ( .A1(n1267), .A2(n1266), .ZN(n1271) );
INV_X1 U1071 ( .A(n1291), .ZN(n1266) );
NAND2_X1 U1072 ( .A1(n1366), .A2(n1367), .ZN(n1291) );
OR2_X1 U1073 ( .A1(n1120), .A2(n1125), .ZN(n1367) );
XOR2_X1 U1074 ( .A(n1368), .B(KEYINPUT53), .Z(n1366) );
NAND2_X1 U1075 ( .A1(n1125), .A2(n1120), .ZN(n1368) );
INV_X1 U1076 ( .A(G475), .ZN(n1120) );
NOR2_X1 U1077 ( .A1(n1184), .A2(G902), .ZN(n1125) );
INV_X1 U1078 ( .A(n1182), .ZN(n1184) );
XOR2_X1 U1079 ( .A(n1369), .B(n1370), .Z(n1182) );
XOR2_X1 U1080 ( .A(G104), .B(n1371), .Z(n1370) );
XOR2_X1 U1081 ( .A(G122), .B(G113), .Z(n1371) );
XOR2_X1 U1082 ( .A(n1372), .B(n1328), .Z(n1369) );
XNOR2_X1 U1083 ( .A(n1373), .B(n1141), .ZN(n1328) );
XOR2_X1 U1084 ( .A(G125), .B(G140), .Z(n1141) );
XOR2_X1 U1085 ( .A(n1359), .B(KEYINPUT1), .Z(n1373) );
INV_X1 U1086 ( .A(G146), .ZN(n1359) );
NAND3_X1 U1087 ( .A1(n1374), .A2(n1375), .A3(n1376), .ZN(n1372) );
OR2_X1 U1088 ( .A1(n1377), .A2(G131), .ZN(n1376) );
NAND2_X1 U1089 ( .A1(KEYINPUT35), .A2(n1378), .ZN(n1375) );
NAND2_X1 U1090 ( .A1(n1379), .A2(n1377), .ZN(n1378) );
XNOR2_X1 U1091 ( .A(KEYINPUT20), .B(G131), .ZN(n1379) );
NAND2_X1 U1092 ( .A1(n1380), .A2(n1381), .ZN(n1374) );
INV_X1 U1093 ( .A(KEYINPUT35), .ZN(n1381) );
NAND2_X1 U1094 ( .A1(n1382), .A2(n1383), .ZN(n1380) );
OR2_X1 U1095 ( .A1(G131), .A2(KEYINPUT20), .ZN(n1383) );
NAND3_X1 U1096 ( .A1(G131), .A2(n1377), .A3(KEYINPUT20), .ZN(n1382) );
XOR2_X1 U1097 ( .A(n1384), .B(G143), .Z(n1377) );
NAND2_X1 U1098 ( .A1(G214), .A2(n1337), .ZN(n1384) );
NOR2_X1 U1099 ( .A1(G953), .A2(G237), .ZN(n1337) );
XNOR2_X1 U1100 ( .A(n1112), .B(KEYINPUT5), .ZN(n1267) );
XNOR2_X1 U1101 ( .A(n1385), .B(G478), .ZN(n1112) );
OR2_X1 U1102 ( .A1(n1177), .A2(G902), .ZN(n1385) );
XNOR2_X1 U1103 ( .A(n1386), .B(n1387), .ZN(n1177) );
XNOR2_X1 U1104 ( .A(n1388), .B(n1309), .ZN(n1387) );
XOR2_X1 U1105 ( .A(G107), .B(KEYINPUT60), .Z(n1309) );
NAND2_X1 U1106 ( .A1(n1326), .A2(G217), .ZN(n1388) );
AND2_X1 U1107 ( .A1(G234), .A2(n1137), .ZN(n1326) );
INV_X1 U1108 ( .A(G953), .ZN(n1137) );
XOR2_X1 U1109 ( .A(n1389), .B(n1390), .Z(n1386) );
NOR2_X1 U1110 ( .A1(n1391), .A2(n1392), .ZN(n1390) );
XOR2_X1 U1111 ( .A(n1393), .B(KEYINPUT46), .Z(n1392) );
NAND2_X1 U1112 ( .A1(G116), .A2(n1288), .ZN(n1393) );
NOR2_X1 U1113 ( .A1(G116), .A2(n1288), .ZN(n1391) );
INV_X1 U1114 ( .A(G122), .ZN(n1288) );
NAND2_X1 U1115 ( .A1(n1394), .A2(n1395), .ZN(n1389) );
NAND2_X1 U1116 ( .A1(G134), .A2(n1396), .ZN(n1395) );
XOR2_X1 U1117 ( .A(KEYINPUT38), .B(n1397), .Z(n1394) );
NOR2_X1 U1118 ( .A1(G134), .A2(n1396), .ZN(n1397) );
XOR2_X1 U1119 ( .A(n1398), .B(n1264), .Z(n1396) );
INV_X1 U1120 ( .A(G143), .ZN(n1264) );
NAND2_X1 U1121 ( .A1(KEYINPUT24), .A2(G128), .ZN(n1398) );
endmodule


