//Key = 1111100110111111101100000001010000000010011110110111111100000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426;

NAND2_X1 U781 ( .A1(n1093), .A2(n1094), .ZN(G9) );
NAND2_X1 U782 ( .A1(G107), .A2(n1095), .ZN(n1094) );
XOR2_X1 U783 ( .A(KEYINPUT7), .B(n1096), .Z(n1093) );
NOR2_X1 U784 ( .A1(G107), .A2(n1095), .ZN(n1096) );
NAND3_X1 U785 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1095) );
XNOR2_X1 U786 ( .A(n1100), .B(KEYINPUT49), .ZN(n1099) );
NOR2_X1 U787 ( .A1(n1101), .A2(n1102), .ZN(G75) );
NOR3_X1 U788 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
NOR2_X1 U789 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NOR2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
INV_X1 U792 ( .A(n1112), .ZN(n1111) );
NOR2_X1 U793 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
NOR2_X1 U794 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NOR3_X1 U795 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1108) );
NOR2_X1 U796 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U797 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
NOR2_X1 U799 ( .A1(n1126), .A2(n1127), .ZN(n1124) );
NOR2_X1 U800 ( .A1(n1128), .A2(n1129), .ZN(n1120) );
NOR2_X1 U801 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
NAND3_X1 U802 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1103) );
NAND3_X1 U803 ( .A1(n1135), .A2(n1136), .A3(n1112), .ZN(n1134) );
NOR3_X1 U804 ( .A1(n1123), .A2(n1118), .A3(n1129), .ZN(n1112) );
INV_X1 U805 ( .A(n1137), .ZN(n1118) );
NOR3_X1 U806 ( .A1(n1138), .A2(G953), .A3(G952), .ZN(n1101) );
INV_X1 U807 ( .A(n1132), .ZN(n1138) );
NAND4_X1 U808 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1132) );
NOR3_X1 U809 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1142) );
XNOR2_X1 U810 ( .A(n1146), .B(n1147), .ZN(n1145) );
NOR2_X1 U811 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U812 ( .A(KEYINPUT16), .B(KEYINPUT11), .Z(n1149) );
XOR2_X1 U813 ( .A(n1150), .B(n1151), .Z(n1144) );
NAND2_X1 U814 ( .A1(KEYINPUT8), .A2(n1152), .ZN(n1150) );
NAND3_X1 U815 ( .A1(n1127), .A2(n1153), .A3(n1116), .ZN(n1143) );
NOR3_X1 U816 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1141) );
NOR2_X1 U817 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
INV_X1 U818 ( .A(KEYINPUT32), .ZN(n1158) );
NOR2_X1 U819 ( .A1(KEYINPUT32), .A2(n1159), .ZN(n1155) );
XNOR2_X1 U820 ( .A(G478), .B(n1160), .ZN(n1154) );
NAND2_X1 U821 ( .A1(KEYINPUT27), .A2(n1161), .ZN(n1160) );
INV_X1 U822 ( .A(n1126), .ZN(n1139) );
XOR2_X1 U823 ( .A(n1162), .B(n1163), .Z(G72) );
XOR2_X1 U824 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND3_X1 U825 ( .A1(G953), .A2(n1166), .A3(KEYINPUT41), .ZN(n1165) );
NAND2_X1 U826 ( .A1(G900), .A2(G227), .ZN(n1166) );
NAND3_X1 U827 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1164) );
XOR2_X1 U828 ( .A(n1170), .B(KEYINPUT35), .Z(n1169) );
NAND2_X1 U829 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND2_X1 U830 ( .A1(G953), .A2(n1173), .ZN(n1168) );
OR2_X1 U831 ( .A1(n1172), .A2(n1171), .ZN(n1167) );
NAND2_X1 U832 ( .A1(n1174), .A2(n1175), .ZN(n1172) );
NAND2_X1 U833 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U834 ( .A(n1178), .B(KEYINPUT39), .Z(n1174) );
OR2_X1 U835 ( .A1(n1177), .A2(n1176), .ZN(n1178) );
XOR2_X1 U836 ( .A(G134), .B(n1179), .Z(n1176) );
XOR2_X1 U837 ( .A(n1180), .B(KEYINPUT60), .Z(n1177) );
NOR2_X1 U838 ( .A1(n1181), .A2(n1182), .ZN(n1162) );
AND2_X1 U839 ( .A1(KEYINPUT14), .A2(n1183), .ZN(n1182) );
NOR2_X1 U840 ( .A1(KEYINPUT18), .A2(n1183), .ZN(n1181) );
NAND2_X1 U841 ( .A1(n1133), .A2(n1184), .ZN(n1183) );
XOR2_X1 U842 ( .A(n1185), .B(n1186), .Z(G69) );
XOR2_X1 U843 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND2_X1 U844 ( .A1(G953), .A2(n1189), .ZN(n1188) );
NAND2_X1 U845 ( .A1(G898), .A2(G224), .ZN(n1189) );
NAND2_X1 U846 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
NAND2_X1 U847 ( .A1(G953), .A2(n1192), .ZN(n1191) );
XOR2_X1 U848 ( .A(n1193), .B(n1194), .Z(n1190) );
NOR2_X1 U849 ( .A1(KEYINPUT24), .A2(n1195), .ZN(n1193) );
AND2_X1 U850 ( .A1(n1196), .A2(n1133), .ZN(n1185) );
NOR2_X1 U851 ( .A1(n1197), .A2(n1198), .ZN(G66) );
NOR3_X1 U852 ( .A1(n1146), .A2(n1199), .A3(n1200), .ZN(n1198) );
AND3_X1 U853 ( .A1(n1201), .A2(n1148), .A3(n1202), .ZN(n1200) );
INV_X1 U854 ( .A(n1203), .ZN(n1148) );
NOR2_X1 U855 ( .A1(n1204), .A2(n1201), .ZN(n1199) );
NOR2_X1 U856 ( .A1(n1205), .A2(n1203), .ZN(n1204) );
NOR2_X1 U857 ( .A1(n1197), .A2(n1206), .ZN(G63) );
XOR2_X1 U858 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR2_X1 U859 ( .A1(KEYINPUT36), .A2(n1209), .ZN(n1208) );
NAND2_X1 U860 ( .A1(n1202), .A2(G478), .ZN(n1207) );
NOR2_X1 U861 ( .A1(n1197), .A2(n1210), .ZN(G60) );
NOR3_X1 U862 ( .A1(n1151), .A2(n1211), .A3(n1212), .ZN(n1210) );
AND2_X1 U863 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NOR3_X1 U864 ( .A1(n1214), .A2(n1215), .A3(n1213), .ZN(n1211) );
NAND3_X1 U865 ( .A1(G475), .A2(n1105), .A3(KEYINPUT10), .ZN(n1213) );
XNOR2_X1 U866 ( .A(G104), .B(n1216), .ZN(G6) );
NAND3_X1 U867 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1216) );
NOR3_X1 U868 ( .A1(n1123), .A2(n1220), .A3(n1221), .ZN(n1219) );
XNOR2_X1 U869 ( .A(n1125), .B(KEYINPUT4), .ZN(n1217) );
NOR2_X1 U870 ( .A1(n1222), .A2(n1223), .ZN(G57) );
XOR2_X1 U871 ( .A(KEYINPUT20), .B(n1197), .Z(n1223) );
XOR2_X1 U872 ( .A(n1224), .B(n1225), .Z(n1222) );
XOR2_X1 U873 ( .A(n1226), .B(n1227), .Z(n1224) );
NAND2_X1 U874 ( .A1(n1202), .A2(n1228), .ZN(n1226) );
XOR2_X1 U875 ( .A(KEYINPUT31), .B(G472), .Z(n1228) );
NOR3_X1 U876 ( .A1(n1197), .A2(n1229), .A3(n1230), .ZN(G54) );
NOR2_X1 U877 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XOR2_X1 U878 ( .A(n1233), .B(n1234), .Z(n1231) );
NOR2_X1 U879 ( .A1(n1235), .A2(n1236), .ZN(n1233) );
INV_X1 U880 ( .A(KEYINPUT3), .ZN(n1236) );
NOR2_X1 U881 ( .A1(n1237), .A2(n1238), .ZN(n1229) );
XOR2_X1 U882 ( .A(n1239), .B(n1234), .Z(n1238) );
XNOR2_X1 U883 ( .A(n1240), .B(n1241), .ZN(n1234) );
XOR2_X1 U884 ( .A(n1242), .B(n1243), .Z(n1241) );
NOR2_X1 U885 ( .A1(KEYINPUT5), .A2(n1244), .ZN(n1242) );
XOR2_X1 U886 ( .A(n1245), .B(KEYINPUT15), .Z(n1240) );
NAND2_X1 U887 ( .A1(n1202), .A2(G469), .ZN(n1245) );
NOR2_X1 U888 ( .A1(n1215), .A2(n1205), .ZN(n1202) );
AND2_X1 U889 ( .A1(n1235), .A2(KEYINPUT3), .ZN(n1239) );
NAND3_X1 U890 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1235) );
NAND2_X1 U891 ( .A1(KEYINPUT58), .A2(G110), .ZN(n1248) );
OR3_X1 U892 ( .A1(n1249), .A2(KEYINPUT58), .A3(G140), .ZN(n1247) );
NAND2_X1 U893 ( .A1(G140), .A2(n1249), .ZN(n1246) );
NAND2_X1 U894 ( .A1(KEYINPUT54), .A2(n1250), .ZN(n1249) );
INV_X1 U895 ( .A(n1232), .ZN(n1237) );
NOR2_X1 U896 ( .A1(n1197), .A2(n1251), .ZN(G51) );
XOR2_X1 U897 ( .A(n1252), .B(n1253), .Z(n1251) );
XNOR2_X1 U898 ( .A(n1254), .B(n1255), .ZN(n1253) );
XOR2_X1 U899 ( .A(n1256), .B(n1257), .Z(n1252) );
XNOR2_X1 U900 ( .A(G125), .B(n1258), .ZN(n1257) );
NAND4_X1 U901 ( .A1(G210), .A2(n1259), .A3(n1260), .A4(n1105), .ZN(n1256) );
INV_X1 U902 ( .A(n1205), .ZN(n1105) );
NOR2_X1 U903 ( .A1(n1196), .A2(n1184), .ZN(n1205) );
NAND4_X1 U904 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1184) );
NOR4_X1 U905 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1264) );
INV_X1 U906 ( .A(n1269), .ZN(n1268) );
NOR2_X1 U907 ( .A1(n1270), .A2(n1271), .ZN(n1263) );
AND2_X1 U908 ( .A1(KEYINPUT2), .A2(n1272), .ZN(n1271) );
NOR3_X1 U909 ( .A1(KEYINPUT2), .A2(n1273), .A3(n1274), .ZN(n1270) );
NAND3_X1 U910 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1262) );
OR2_X1 U911 ( .A1(n1278), .A2(KEYINPUT45), .ZN(n1276) );
NAND2_X1 U912 ( .A1(KEYINPUT45), .A2(n1279), .ZN(n1275) );
NAND2_X1 U913 ( .A1(n1280), .A2(n1114), .ZN(n1279) );
INV_X1 U914 ( .A(n1221), .ZN(n1114) );
NAND2_X1 U915 ( .A1(n1125), .A2(n1281), .ZN(n1261) );
NAND2_X1 U916 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
XOR2_X1 U917 ( .A(KEYINPUT13), .B(n1284), .Z(n1282) );
NOR4_X1 U918 ( .A1(n1285), .A2(n1286), .A3(n1287), .A4(n1288), .ZN(n1284) );
NOR2_X1 U919 ( .A1(n1289), .A2(n1290), .ZN(n1286) );
INV_X1 U920 ( .A(KEYINPUT21), .ZN(n1290) );
NOR2_X1 U921 ( .A1(n1221), .A2(n1291), .ZN(n1289) );
NOR2_X1 U922 ( .A1(KEYINPUT21), .A2(n1278), .ZN(n1285) );
NAND4_X1 U923 ( .A1(n1292), .A2(n1293), .A3(n1294), .A4(n1295), .ZN(n1196) );
AND4_X1 U924 ( .A1(n1296), .A2(n1297), .A3(n1298), .A4(n1299), .ZN(n1295) );
NAND3_X1 U925 ( .A1(n1098), .A2(n1136), .A3(n1097), .ZN(n1294) );
NAND2_X1 U926 ( .A1(n1300), .A2(n1287), .ZN(n1136) );
INV_X1 U927 ( .A(n1100), .ZN(n1287) );
XNOR2_X1 U928 ( .A(KEYINPUT40), .B(n1215), .ZN(n1259) );
AND2_X1 U929 ( .A1(n1301), .A2(G953), .ZN(n1197) );
XNOR2_X1 U930 ( .A(G952), .B(KEYINPUT48), .ZN(n1301) );
XOR2_X1 U931 ( .A(G146), .B(n1302), .Z(G48) );
NOR2_X1 U932 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
XOR2_X1 U933 ( .A(n1283), .B(KEYINPUT33), .Z(n1303) );
NAND3_X1 U934 ( .A1(n1305), .A2(n1218), .A3(n1278), .ZN(n1283) );
XNOR2_X1 U935 ( .A(G143), .B(n1306), .ZN(G45) );
NOR2_X1 U936 ( .A1(n1272), .A2(KEYINPUT34), .ZN(n1306) );
NOR2_X1 U937 ( .A1(n1274), .A2(n1307), .ZN(n1272) );
INV_X1 U938 ( .A(n1273), .ZN(n1307) );
NAND3_X1 U939 ( .A1(n1131), .A2(n1125), .A3(n1278), .ZN(n1274) );
XNOR2_X1 U940 ( .A(G140), .B(n1269), .ZN(G42) );
NAND4_X1 U941 ( .A1(n1278), .A2(n1308), .A3(n1218), .A4(n1130), .ZN(n1269) );
XNOR2_X1 U942 ( .A(G137), .B(n1309), .ZN(G39) );
NAND2_X1 U943 ( .A1(n1277), .A2(n1278), .ZN(n1309) );
NOR3_X1 U944 ( .A1(n1288), .A2(n1107), .A3(n1129), .ZN(n1277) );
XNOR2_X1 U945 ( .A(n1310), .B(n1267), .ZN(G36) );
AND2_X1 U946 ( .A1(n1311), .A2(n1100), .ZN(n1267) );
XOR2_X1 U947 ( .A(G131), .B(n1266), .Z(G33) );
AND2_X1 U948 ( .A1(n1311), .A2(n1218), .ZN(n1266) );
AND3_X1 U949 ( .A1(n1308), .A2(n1131), .A3(n1278), .ZN(n1311) );
INV_X1 U950 ( .A(n1129), .ZN(n1308) );
NAND2_X1 U951 ( .A1(n1312), .A2(n1127), .ZN(n1129) );
XNOR2_X1 U952 ( .A(n1126), .B(KEYINPUT37), .ZN(n1312) );
XNOR2_X1 U953 ( .A(G128), .B(n1313), .ZN(G30) );
NAND4_X1 U954 ( .A1(n1278), .A2(n1305), .A3(n1100), .A4(n1125), .ZN(n1313) );
NOR2_X1 U955 ( .A1(n1221), .A2(n1280), .ZN(n1278) );
INV_X1 U956 ( .A(n1291), .ZN(n1280) );
XNOR2_X1 U957 ( .A(G101), .B(n1292), .ZN(G3) );
NAND3_X1 U958 ( .A1(n1131), .A2(n1097), .A3(n1314), .ZN(n1292) );
XOR2_X1 U959 ( .A(n1265), .B(n1315), .Z(G27) );
NOR2_X1 U960 ( .A1(KEYINPUT22), .A2(n1316), .ZN(n1315) );
INV_X1 U961 ( .A(G125), .ZN(n1316) );
AND4_X1 U962 ( .A1(n1125), .A2(n1291), .A3(n1135), .A4(n1317), .ZN(n1265) );
NOR2_X1 U963 ( .A1(n1318), .A2(n1300), .ZN(n1317) );
NAND2_X1 U964 ( .A1(n1319), .A2(n1320), .ZN(n1291) );
NAND4_X1 U965 ( .A1(G953), .A2(G902), .A3(n1173), .A4(n1137), .ZN(n1319) );
XOR2_X1 U966 ( .A(KEYINPUT12), .B(G900), .Z(n1173) );
INV_X1 U967 ( .A(n1304), .ZN(n1125) );
XNOR2_X1 U968 ( .A(G122), .B(n1321), .ZN(G24) );
NAND2_X1 U969 ( .A1(KEYINPUT0), .A2(n1322), .ZN(n1321) );
INV_X1 U970 ( .A(n1297), .ZN(n1322) );
NAND3_X1 U971 ( .A1(n1323), .A2(n1098), .A3(n1273), .ZN(n1297) );
NOR2_X1 U972 ( .A1(n1324), .A2(n1325), .ZN(n1273) );
INV_X1 U973 ( .A(n1123), .ZN(n1098) );
NAND2_X1 U974 ( .A1(n1140), .A2(n1326), .ZN(n1123) );
XNOR2_X1 U975 ( .A(G119), .B(n1293), .ZN(G21) );
NAND3_X1 U976 ( .A1(n1314), .A2(n1323), .A3(n1305), .ZN(n1293) );
INV_X1 U977 ( .A(n1288), .ZN(n1305) );
NAND2_X1 U978 ( .A1(n1327), .A2(n1328), .ZN(n1288) );
XNOR2_X1 U979 ( .A(G116), .B(n1296), .ZN(G18) );
NAND3_X1 U980 ( .A1(n1131), .A2(n1100), .A3(n1323), .ZN(n1296) );
NOR2_X1 U981 ( .A1(n1325), .A2(n1329), .ZN(n1100) );
XNOR2_X1 U982 ( .A(G113), .B(n1299), .ZN(G15) );
NAND3_X1 U983 ( .A1(n1323), .A2(n1131), .A3(n1218), .ZN(n1299) );
INV_X1 U984 ( .A(n1300), .ZN(n1218) );
NAND2_X1 U985 ( .A1(n1330), .A2(n1329), .ZN(n1300) );
INV_X1 U986 ( .A(n1324), .ZN(n1329) );
AND2_X1 U987 ( .A1(n1327), .A2(n1326), .ZN(n1131) );
XOR2_X1 U988 ( .A(n1140), .B(KEYINPUT1), .Z(n1327) );
NOR3_X1 U989 ( .A1(n1304), .A2(n1220), .A3(n1117), .ZN(n1323) );
INV_X1 U990 ( .A(n1135), .ZN(n1117) );
NOR2_X1 U991 ( .A1(n1115), .A2(n1331), .ZN(n1135) );
INV_X1 U992 ( .A(n1116), .ZN(n1331) );
XNOR2_X1 U993 ( .A(G110), .B(n1298), .ZN(G12) );
NAND3_X1 U994 ( .A1(n1130), .A2(n1097), .A3(n1314), .ZN(n1298) );
INV_X1 U995 ( .A(n1107), .ZN(n1314) );
NAND2_X1 U996 ( .A1(n1330), .A2(n1324), .ZN(n1107) );
XNOR2_X1 U997 ( .A(n1332), .B(n1151), .ZN(n1324) );
AND2_X1 U998 ( .A1(n1214), .A2(n1215), .ZN(n1151) );
XNOR2_X1 U999 ( .A(n1333), .B(n1334), .ZN(n1214) );
XOR2_X1 U1000 ( .A(n1335), .B(n1336), .Z(n1334) );
XNOR2_X1 U1001 ( .A(n1171), .B(n1337), .ZN(n1336) );
NOR4_X1 U1002 ( .A1(KEYINPUT17), .A2(G953), .A3(G237), .A4(n1338), .ZN(n1337) );
INV_X1 U1003 ( .A(G214), .ZN(n1338) );
XOR2_X1 U1004 ( .A(n1339), .B(n1340), .Z(n1333) );
XNOR2_X1 U1005 ( .A(G131), .B(n1341), .ZN(n1340) );
XNOR2_X1 U1006 ( .A(G104), .B(G113), .ZN(n1339) );
NAND2_X1 U1007 ( .A1(KEYINPUT47), .A2(n1152), .ZN(n1332) );
INV_X1 U1008 ( .A(G475), .ZN(n1152) );
XNOR2_X1 U1009 ( .A(n1342), .B(KEYINPUT59), .ZN(n1330) );
INV_X1 U1010 ( .A(n1325), .ZN(n1342) );
XNOR2_X1 U1011 ( .A(n1161), .B(G478), .ZN(n1325) );
NOR2_X1 U1012 ( .A1(n1209), .A2(G902), .ZN(n1161) );
XOR2_X1 U1013 ( .A(n1343), .B(n1344), .Z(n1209) );
NOR2_X1 U1014 ( .A1(KEYINPUT25), .A2(n1345), .ZN(n1344) );
XOR2_X1 U1015 ( .A(n1346), .B(n1347), .Z(n1345) );
XNOR2_X1 U1016 ( .A(G107), .B(n1348), .ZN(n1347) );
NAND2_X1 U1017 ( .A1(n1349), .A2(KEYINPUT51), .ZN(n1348) );
XNOR2_X1 U1018 ( .A(G128), .B(n1350), .ZN(n1349) );
XNOR2_X1 U1019 ( .A(n1351), .B(G134), .ZN(n1350) );
INV_X1 U1020 ( .A(G143), .ZN(n1351) );
XNOR2_X1 U1021 ( .A(n1341), .B(G116), .ZN(n1346) );
NAND3_X1 U1022 ( .A1(G234), .A2(n1133), .A3(G217), .ZN(n1343) );
NOR3_X1 U1023 ( .A1(n1304), .A2(n1220), .A3(n1221), .ZN(n1097) );
NAND2_X1 U1024 ( .A1(n1116), .A2(n1115), .ZN(n1221) );
NAND2_X1 U1025 ( .A1(n1352), .A2(n1153), .ZN(n1115) );
OR2_X1 U1026 ( .A1(n1157), .A2(G469), .ZN(n1153) );
XOR2_X1 U1027 ( .A(n1159), .B(KEYINPUT28), .Z(n1352) );
NAND2_X1 U1028 ( .A1(G469), .A2(n1157), .ZN(n1159) );
NAND3_X1 U1029 ( .A1(n1353), .A2(n1354), .A3(n1215), .ZN(n1157) );
NAND2_X1 U1030 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
INV_X1 U1031 ( .A(KEYINPUT57), .ZN(n1356) );
XOR2_X1 U1032 ( .A(n1357), .B(n1358), .Z(n1355) );
NAND3_X1 U1033 ( .A1(n1357), .A2(n1358), .A3(KEYINPUT57), .ZN(n1353) );
XOR2_X1 U1034 ( .A(n1232), .B(n1359), .Z(n1358) );
XNOR2_X1 U1035 ( .A(n1250), .B(n1360), .ZN(n1359) );
NOR2_X1 U1036 ( .A1(KEYINPUT61), .A2(n1361), .ZN(n1360) );
INV_X1 U1037 ( .A(G140), .ZN(n1361) );
INV_X1 U1038 ( .A(G110), .ZN(n1250) );
NAND2_X1 U1039 ( .A1(G227), .A2(n1133), .ZN(n1232) );
XNOR2_X1 U1040 ( .A(n1243), .B(n1244), .ZN(n1357) );
INV_X1 U1041 ( .A(n1362), .ZN(n1244) );
XOR2_X1 U1042 ( .A(n1363), .B(n1364), .Z(n1243) );
INV_X1 U1043 ( .A(n1180), .ZN(n1364) );
XNOR2_X1 U1044 ( .A(n1335), .B(n1365), .ZN(n1180) );
NOR2_X1 U1045 ( .A1(KEYINPUT26), .A2(n1366), .ZN(n1365) );
XOR2_X1 U1046 ( .A(n1367), .B(G101), .Z(n1363) );
NAND2_X1 U1047 ( .A1(KEYINPUT55), .A2(n1368), .ZN(n1367) );
NAND2_X1 U1048 ( .A1(G221), .A2(n1369), .ZN(n1116) );
AND2_X1 U1049 ( .A1(n1320), .A2(n1370), .ZN(n1220) );
NAND4_X1 U1050 ( .A1(n1371), .A2(G953), .A3(n1137), .A4(n1192), .ZN(n1370) );
INV_X1 U1051 ( .A(G898), .ZN(n1192) );
XNOR2_X1 U1052 ( .A(G902), .B(KEYINPUT53), .ZN(n1371) );
NAND3_X1 U1053 ( .A1(G952), .A2(n1137), .A3(n1372), .ZN(n1320) );
XNOR2_X1 U1054 ( .A(G953), .B(KEYINPUT56), .ZN(n1372) );
NAND2_X1 U1055 ( .A1(G237), .A2(G234), .ZN(n1137) );
NAND2_X1 U1056 ( .A1(n1126), .A2(n1127), .ZN(n1304) );
NAND2_X1 U1057 ( .A1(G214), .A2(n1260), .ZN(n1127) );
XNOR2_X1 U1058 ( .A(n1373), .B(n1374), .ZN(n1126) );
AND2_X1 U1059 ( .A1(n1260), .A2(G210), .ZN(n1374) );
NAND2_X1 U1060 ( .A1(n1375), .A2(n1215), .ZN(n1260) );
XNOR2_X1 U1061 ( .A(G237), .B(KEYINPUT63), .ZN(n1375) );
NAND2_X1 U1062 ( .A1(n1376), .A2(n1215), .ZN(n1373) );
XNOR2_X1 U1063 ( .A(n1255), .B(n1377), .ZN(n1376) );
NOR3_X1 U1064 ( .A1(n1378), .A2(n1379), .A3(n1380), .ZN(n1377) );
NOR2_X1 U1065 ( .A1(KEYINPUT46), .A2(n1258), .ZN(n1380) );
AND4_X1 U1066 ( .A1(n1258), .A2(KEYINPUT46), .A3(KEYINPUT29), .A4(n1381), .ZN(n1379) );
NOR2_X1 U1067 ( .A1(n1382), .A2(n1381), .ZN(n1378) );
XOR2_X1 U1068 ( .A(n1383), .B(G125), .Z(n1381) );
NAND2_X1 U1069 ( .A1(KEYINPUT38), .A2(n1254), .ZN(n1383) );
AND2_X1 U1070 ( .A1(n1258), .A2(KEYINPUT29), .ZN(n1382) );
AND2_X1 U1071 ( .A1(G224), .A2(n1133), .ZN(n1258) );
XNOR2_X1 U1072 ( .A(n1195), .B(n1194), .ZN(n1255) );
XNOR2_X1 U1073 ( .A(n1384), .B(G110), .ZN(n1194) );
NAND2_X1 U1074 ( .A1(KEYINPUT19), .A2(n1341), .ZN(n1384) );
INV_X1 U1075 ( .A(G122), .ZN(n1341) );
XOR2_X1 U1076 ( .A(n1385), .B(n1368), .Z(n1195) );
XOR2_X1 U1077 ( .A(G104), .B(G107), .Z(n1368) );
XOR2_X1 U1078 ( .A(n1386), .B(G101), .Z(n1385) );
NAND3_X1 U1079 ( .A1(n1387), .A2(n1388), .A3(n1389), .ZN(n1386) );
INV_X1 U1080 ( .A(n1390), .ZN(n1389) );
NAND2_X1 U1081 ( .A1(n1391), .A2(n1392), .ZN(n1388) );
INV_X1 U1082 ( .A(KEYINPUT30), .ZN(n1392) );
NAND2_X1 U1083 ( .A1(n1393), .A2(KEYINPUT30), .ZN(n1387) );
XNOR2_X1 U1084 ( .A(G113), .B(n1394), .ZN(n1393) );
NAND2_X1 U1085 ( .A1(G119), .A2(n1395), .ZN(n1394) );
INV_X1 U1086 ( .A(n1318), .ZN(n1130) );
NAND2_X1 U1087 ( .A1(n1140), .A2(n1328), .ZN(n1318) );
INV_X1 U1088 ( .A(n1326), .ZN(n1328) );
XOR2_X1 U1089 ( .A(n1146), .B(n1203), .Z(n1326) );
NAND2_X1 U1090 ( .A1(G217), .A2(n1369), .ZN(n1203) );
NAND2_X1 U1091 ( .A1(G234), .A2(n1215), .ZN(n1369) );
NOR2_X1 U1092 ( .A1(n1201), .A2(G902), .ZN(n1146) );
XOR2_X1 U1093 ( .A(n1396), .B(n1397), .Z(n1201) );
XOR2_X1 U1094 ( .A(n1398), .B(n1399), .Z(n1397) );
NAND4_X1 U1095 ( .A1(n1400), .A2(n1401), .A3(n1402), .A4(n1403), .ZN(n1399) );
NAND3_X1 U1096 ( .A1(n1404), .A2(n1405), .A3(n1406), .ZN(n1403) );
INV_X1 U1097 ( .A(KEYINPUT42), .ZN(n1406) );
OR2_X1 U1098 ( .A1(KEYINPUT52), .A2(G128), .ZN(n1404) );
NAND3_X1 U1099 ( .A1(G119), .A2(n1407), .A3(KEYINPUT42), .ZN(n1402) );
NAND2_X1 U1100 ( .A1(KEYINPUT52), .A2(n1366), .ZN(n1407) );
NAND3_X1 U1101 ( .A1(n1408), .A2(n1366), .A3(n1409), .ZN(n1401) );
INV_X1 U1102 ( .A(KEYINPUT6), .ZN(n1409) );
XNOR2_X1 U1103 ( .A(KEYINPUT52), .B(n1405), .ZN(n1408) );
NAND2_X1 U1104 ( .A1(KEYINPUT6), .A2(G128), .ZN(n1400) );
NAND2_X1 U1105 ( .A1(KEYINPUT43), .A2(n1410), .ZN(n1398) );
XOR2_X1 U1106 ( .A(G146), .B(n1171), .Z(n1410) );
XOR2_X1 U1107 ( .A(G125), .B(G140), .Z(n1171) );
XOR2_X1 U1108 ( .A(n1411), .B(n1412), .Z(n1396) );
AND3_X1 U1109 ( .A1(G221), .A2(n1133), .A3(G234), .ZN(n1412) );
INV_X1 U1110 ( .A(G953), .ZN(n1133) );
XNOR2_X1 U1111 ( .A(G137), .B(G110), .ZN(n1411) );
XOR2_X1 U1112 ( .A(n1413), .B(G472), .Z(n1140) );
NAND2_X1 U1113 ( .A1(n1414), .A2(n1215), .ZN(n1413) );
INV_X1 U1114 ( .A(G902), .ZN(n1215) );
XNOR2_X1 U1115 ( .A(n1225), .B(n1415), .ZN(n1414) );
XNOR2_X1 U1116 ( .A(n1416), .B(KEYINPUT62), .ZN(n1415) );
NAND2_X1 U1117 ( .A1(KEYINPUT50), .A2(n1227), .ZN(n1416) );
NOR3_X1 U1118 ( .A1(G237), .A2(G953), .A3(n1417), .ZN(n1227) );
INV_X1 U1119 ( .A(G210), .ZN(n1417) );
XNOR2_X1 U1120 ( .A(n1418), .B(n1419), .ZN(n1225) );
XNOR2_X1 U1121 ( .A(n1254), .B(n1362), .ZN(n1419) );
XOR2_X1 U1122 ( .A(n1179), .B(n1420), .Z(n1362) );
NOR2_X1 U1123 ( .A1(KEYINPUT23), .A2(n1310), .ZN(n1420) );
INV_X1 U1124 ( .A(G134), .ZN(n1310) );
XOR2_X1 U1125 ( .A(G131), .B(G137), .Z(n1179) );
XNOR2_X1 U1126 ( .A(n1366), .B(n1335), .ZN(n1254) );
XNOR2_X1 U1127 ( .A(G143), .B(G146), .ZN(n1335) );
INV_X1 U1128 ( .A(G128), .ZN(n1366) );
XOR2_X1 U1129 ( .A(n1421), .B(n1422), .Z(n1418) );
NOR2_X1 U1130 ( .A1(n1390), .A2(n1391), .ZN(n1422) );
NAND2_X1 U1131 ( .A1(n1423), .A2(n1424), .ZN(n1391) );
NAND2_X1 U1132 ( .A1(n1425), .A2(G119), .ZN(n1424) );
XNOR2_X1 U1133 ( .A(G113), .B(n1395), .ZN(n1425) );
NAND3_X1 U1134 ( .A1(n1395), .A2(n1426), .A3(n1405), .ZN(n1423) );
INV_X1 U1135 ( .A(G119), .ZN(n1405) );
NOR3_X1 U1136 ( .A1(n1395), .A2(G119), .A3(n1426), .ZN(n1390) );
INV_X1 U1137 ( .A(G113), .ZN(n1426) );
XOR2_X1 U1138 ( .A(G116), .B(KEYINPUT44), .Z(n1395) );
XNOR2_X1 U1139 ( .A(G101), .B(KEYINPUT9), .ZN(n1421) );
endmodule


