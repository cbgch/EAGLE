//Key = 1000010100010010100110000000110010011010101111000001101110000011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379;

XOR2_X1 U759 ( .A(G107), .B(n1046), .Z(G9) );
NAND3_X1 U760 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(G75) );
NAND2_X1 U761 ( .A1(G952), .A2(n1050), .ZN(n1049) );
NAND3_X1 U762 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1050) );
NAND2_X1 U763 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NAND2_X1 U764 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND3_X1 U765 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
NAND2_X1 U766 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NAND2_X1 U767 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U768 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1061) );
NAND2_X1 U770 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
OR3_X1 U771 ( .A1(n1071), .A2(KEYINPUT57), .A3(n1072), .ZN(n1070) );
NAND3_X1 U772 ( .A1(n1067), .A2(n1073), .A3(n1063), .ZN(n1056) );
NAND2_X1 U773 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U774 ( .A1(n1060), .A2(n1076), .ZN(n1075) );
NAND2_X1 U775 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U776 ( .A1(n1058), .A2(n1079), .ZN(n1074) );
NAND3_X1 U777 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NAND3_X1 U778 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1081) );
INV_X1 U779 ( .A(KEYINPUT39), .ZN(n1085) );
NAND2_X1 U780 ( .A1(KEYINPUT39), .A2(n1060), .ZN(n1080) );
NAND2_X1 U781 ( .A1(KEYINPUT57), .A2(n1086), .ZN(n1051) );
NAND4_X1 U782 ( .A1(n1054), .A2(n1058), .A3(n1067), .A4(n1087), .ZN(n1086) );
NOR3_X1 U783 ( .A1(n1072), .A2(n1088), .A3(n1071), .ZN(n1087) );
XNOR2_X1 U784 ( .A(KEYINPUT11), .B(n1089), .ZN(n1054) );
NAND4_X1 U785 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1047) );
NOR4_X1 U786 ( .A1(n1094), .A2(n1083), .A3(n1095), .A4(n1096), .ZN(n1093) );
XOR2_X1 U787 ( .A(n1097), .B(n1098), .Z(n1095) );
NOR2_X1 U788 ( .A1(KEYINPUT17), .A2(n1099), .ZN(n1098) );
XOR2_X1 U789 ( .A(n1100), .B(KEYINPUT62), .Z(n1099) );
NOR3_X1 U790 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1092) );
NOR2_X1 U791 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XOR2_X1 U792 ( .A(n1106), .B(KEYINPUT29), .Z(n1105) );
NOR2_X1 U793 ( .A1(n1107), .A2(n1106), .ZN(n1102) );
XNOR2_X1 U794 ( .A(G472), .B(n1108), .ZN(n1101) );
XNOR2_X1 U795 ( .A(n1109), .B(n1110), .ZN(n1091) );
NAND2_X1 U796 ( .A1(KEYINPUT38), .A2(n1111), .ZN(n1109) );
XOR2_X1 U797 ( .A(n1112), .B(n1113), .Z(n1090) );
XOR2_X1 U798 ( .A(KEYINPUT48), .B(G469), .Z(n1113) );
XOR2_X1 U799 ( .A(n1114), .B(n1115), .Z(G72) );
NOR2_X1 U800 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U801 ( .A(n1118), .B(KEYINPUT5), .Z(n1117) );
NAND3_X1 U802 ( .A1(n1119), .A2(n1048), .A3(n1120), .ZN(n1118) );
NOR2_X1 U803 ( .A1(n1121), .A2(n1120), .ZN(n1116) );
NAND2_X1 U804 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
NAND2_X1 U805 ( .A1(G953), .A2(n1124), .ZN(n1123) );
XOR2_X1 U806 ( .A(n1125), .B(n1126), .Z(n1122) );
NOR2_X1 U807 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
XOR2_X1 U808 ( .A(n1129), .B(KEYINPUT42), .Z(n1128) );
NAND2_X1 U809 ( .A1(G140), .A2(n1130), .ZN(n1129) );
NOR2_X1 U810 ( .A1(G140), .A2(n1130), .ZN(n1127) );
XNOR2_X1 U811 ( .A(KEYINPUT35), .B(n1131), .ZN(n1130) );
NOR2_X1 U812 ( .A1(G953), .A2(n1132), .ZN(n1121) );
NAND2_X1 U813 ( .A1(G953), .A2(n1133), .ZN(n1114) );
NAND2_X1 U814 ( .A1(G900), .A2(G227), .ZN(n1133) );
XOR2_X1 U815 ( .A(n1134), .B(n1135), .Z(G69) );
XOR2_X1 U816 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U817 ( .A1(G953), .A2(n1138), .ZN(n1137) );
NAND2_X1 U818 ( .A1(G898), .A2(G224), .ZN(n1138) );
NAND2_X1 U819 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
NAND2_X1 U820 ( .A1(G953), .A2(n1141), .ZN(n1140) );
XNOR2_X1 U821 ( .A(n1142), .B(n1143), .ZN(n1139) );
NOR2_X1 U822 ( .A1(KEYINPUT2), .A2(n1144), .ZN(n1142) );
NOR2_X1 U823 ( .A1(n1145), .A2(G953), .ZN(n1134) );
NOR2_X1 U824 ( .A1(n1146), .A2(n1147), .ZN(G66) );
NOR3_X1 U825 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1147) );
NOR2_X1 U826 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U827 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U828 ( .A(KEYINPUT50), .B(n1155), .Z(n1154) );
NOR3_X1 U829 ( .A1(n1156), .A2(n1155), .A3(n1153), .ZN(n1149) );
AND2_X1 U830 ( .A1(n1153), .A2(n1155), .ZN(n1148) );
NOR2_X1 U831 ( .A1(n1157), .A2(n1100), .ZN(n1155) );
INV_X1 U832 ( .A(KEYINPUT63), .ZN(n1153) );
NOR2_X1 U833 ( .A1(n1146), .A2(n1158), .ZN(G63) );
NOR3_X1 U834 ( .A1(n1111), .A2(n1159), .A3(n1160), .ZN(n1158) );
AND3_X1 U835 ( .A1(n1161), .A2(G478), .A3(n1162), .ZN(n1160) );
NOR2_X1 U836 ( .A1(n1163), .A2(n1161), .ZN(n1159) );
NOR2_X1 U837 ( .A1(n1053), .A2(n1110), .ZN(n1163) );
NOR2_X1 U838 ( .A1(n1146), .A2(n1164), .ZN(G60) );
XOR2_X1 U839 ( .A(n1165), .B(n1166), .Z(n1164) );
AND2_X1 U840 ( .A1(G475), .A2(n1162), .ZN(n1165) );
XOR2_X1 U841 ( .A(G104), .B(n1167), .Z(G6) );
NOR2_X1 U842 ( .A1(n1168), .A2(n1169), .ZN(G57) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U844 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NOR2_X1 U845 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NOR2_X1 U846 ( .A1(n1176), .A2(n1157), .ZN(n1175) );
NOR2_X1 U847 ( .A1(n1177), .A2(n1178), .ZN(n1174) );
AND2_X1 U848 ( .A1(n1179), .A2(KEYINPUT51), .ZN(n1177) );
NOR2_X1 U849 ( .A1(n1180), .A2(n1179), .ZN(n1172) );
XNOR2_X1 U850 ( .A(n1181), .B(n1182), .ZN(n1179) );
XNOR2_X1 U851 ( .A(KEYINPUT14), .B(n1183), .ZN(n1181) );
NOR2_X1 U852 ( .A1(KEYINPUT25), .A2(n1184), .ZN(n1183) );
XOR2_X1 U853 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U854 ( .A1(KEYINPUT26), .A2(n1187), .ZN(n1185) );
NOR2_X1 U855 ( .A1(n1188), .A2(n1189), .ZN(n1180) );
INV_X1 U856 ( .A(KEYINPUT51), .ZN(n1189) );
NOR3_X1 U857 ( .A1(n1178), .A2(n1176), .A3(n1157), .ZN(n1188) );
INV_X1 U858 ( .A(KEYINPUT32), .ZN(n1178) );
NAND2_X1 U859 ( .A1(n1190), .A2(KEYINPUT56), .ZN(n1170) );
XNOR2_X1 U860 ( .A(n1191), .B(G101), .ZN(n1190) );
NOR2_X1 U861 ( .A1(G952), .A2(n1192), .ZN(n1168) );
XNOR2_X1 U862 ( .A(G953), .B(KEYINPUT33), .ZN(n1192) );
NOR2_X1 U863 ( .A1(n1146), .A2(n1193), .ZN(G54) );
XOR2_X1 U864 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U865 ( .A(n1196), .B(n1197), .Z(n1195) );
XNOR2_X1 U866 ( .A(n1198), .B(G110), .ZN(n1197) );
NOR2_X1 U867 ( .A1(KEYINPUT53), .A2(n1199), .ZN(n1196) );
XNOR2_X1 U868 ( .A(n1200), .B(n1201), .ZN(n1199) );
NOR2_X1 U869 ( .A1(KEYINPUT6), .A2(n1187), .ZN(n1201) );
XOR2_X1 U870 ( .A(n1202), .B(n1186), .Z(n1194) );
XOR2_X1 U871 ( .A(n1203), .B(n1204), .Z(n1202) );
AND2_X1 U872 ( .A1(G469), .A2(n1162), .ZN(n1204) );
NOR2_X1 U873 ( .A1(n1146), .A2(n1205), .ZN(G51) );
XOR2_X1 U874 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U875 ( .A(n1208), .B(n1209), .Z(n1207) );
NOR2_X1 U876 ( .A1(n1106), .A2(n1157), .ZN(n1209) );
INV_X1 U877 ( .A(n1162), .ZN(n1157) );
NOR2_X1 U878 ( .A1(n1210), .A2(n1053), .ZN(n1162) );
AND2_X1 U879 ( .A1(n1145), .A2(n1132), .ZN(n1053) );
INV_X1 U880 ( .A(n1119), .ZN(n1132) );
NAND4_X1 U881 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1119) );
NOR4_X1 U882 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
INV_X1 U883 ( .A(n1219), .ZN(n1217) );
NOR2_X1 U884 ( .A1(n1220), .A2(n1221), .ZN(n1213) );
NAND3_X1 U885 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1212) );
NAND2_X1 U886 ( .A1(n1225), .A2(n1226), .ZN(n1223) );
NAND3_X1 U887 ( .A1(n1063), .A2(n1227), .A3(KEYINPUT19), .ZN(n1226) );
NAND3_X1 U888 ( .A1(n1228), .A2(n1229), .A3(n1063), .ZN(n1211) );
INV_X1 U889 ( .A(KEYINPUT19), .ZN(n1229) );
AND2_X1 U890 ( .A1(n1230), .A2(n1231), .ZN(n1145) );
NOR4_X1 U891 ( .A1(n1232), .A2(n1167), .A3(n1046), .A4(n1233), .ZN(n1231) );
AND3_X1 U892 ( .A1(n1222), .A2(n1234), .A3(n1067), .ZN(n1046) );
AND3_X1 U893 ( .A1(n1067), .A2(n1234), .A3(n1235), .ZN(n1167) );
NOR4_X1 U894 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1230) );
INV_X1 U895 ( .A(n1240), .ZN(n1238) );
INV_X1 U896 ( .A(n1241), .ZN(n1237) );
NOR2_X1 U897 ( .A1(KEYINPUT22), .A2(n1242), .ZN(n1208) );
NOR3_X1 U898 ( .A1(n1243), .A2(n1244), .A3(n1245), .ZN(n1242) );
NOR3_X1 U899 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1245) );
AND2_X1 U900 ( .A1(n1246), .A2(n1247), .ZN(n1244) );
AND2_X1 U901 ( .A1(n1187), .A2(n1249), .ZN(n1247) );
XNOR2_X1 U902 ( .A(KEYINPUT41), .B(n1131), .ZN(n1249) );
NOR2_X1 U903 ( .A1(n1048), .A2(G952), .ZN(n1146) );
XOR2_X1 U904 ( .A(G146), .B(n1216), .Z(G48) );
NOR3_X1 U905 ( .A1(n1250), .A2(n1077), .A3(n1225), .ZN(n1216) );
XOR2_X1 U906 ( .A(G143), .B(n1215), .Z(G45) );
AND4_X1 U907 ( .A1(n1251), .A2(n1096), .A3(n1252), .A4(n1253), .ZN(n1215) );
NOR2_X1 U908 ( .A1(n1065), .A2(n1250), .ZN(n1253) );
INV_X1 U909 ( .A(n1227), .ZN(n1065) );
XNOR2_X1 U910 ( .A(n1198), .B(n1221), .ZN(G42) );
AND2_X1 U911 ( .A1(n1254), .A2(n1255), .ZN(n1221) );
XOR2_X1 U912 ( .A(G137), .B(n1220), .Z(G39) );
AND4_X1 U913 ( .A1(n1063), .A2(n1224), .A3(n1256), .A4(n1058), .ZN(n1220) );
XNOR2_X1 U914 ( .A(G134), .B(n1257), .ZN(G36) );
NOR2_X1 U915 ( .A1(KEYINPUT49), .A2(n1258), .ZN(n1257) );
NOR2_X1 U916 ( .A1(n1259), .A2(n1228), .ZN(n1258) );
NAND3_X1 U917 ( .A1(n1227), .A2(n1222), .A3(n1224), .ZN(n1228) );
XNOR2_X1 U918 ( .A(n1260), .B(n1218), .ZN(G33) );
AND2_X1 U919 ( .A1(n1254), .A2(n1227), .ZN(n1218) );
NOR3_X1 U920 ( .A1(n1250), .A2(n1077), .A3(n1259), .ZN(n1254) );
INV_X1 U921 ( .A(n1063), .ZN(n1259) );
NOR2_X1 U922 ( .A1(n1071), .A2(n1094), .ZN(n1063) );
INV_X1 U923 ( .A(n1072), .ZN(n1094) );
XNOR2_X1 U924 ( .A(G128), .B(n1261), .ZN(G30) );
NAND4_X1 U925 ( .A1(n1262), .A2(n1222), .A3(n1263), .A4(n1264), .ZN(n1261) );
OR2_X1 U926 ( .A1(n1224), .A2(KEYINPUT61), .ZN(n1264) );
INV_X1 U927 ( .A(n1250), .ZN(n1224) );
NAND2_X1 U928 ( .A1(n1265), .A2(n1266), .ZN(n1250) );
NAND2_X1 U929 ( .A1(KEYINPUT61), .A2(n1267), .ZN(n1263) );
NAND2_X1 U930 ( .A1(n1265), .A2(n1082), .ZN(n1267) );
INV_X1 U931 ( .A(n1266), .ZN(n1082) );
INV_X1 U932 ( .A(n1225), .ZN(n1262) );
NAND2_X1 U933 ( .A1(n1256), .A2(n1252), .ZN(n1225) );
XOR2_X1 U934 ( .A(G101), .B(n1232), .Z(G3) );
AND3_X1 U935 ( .A1(n1234), .A2(n1058), .A3(n1227), .ZN(n1232) );
XNOR2_X1 U936 ( .A(G125), .B(n1219), .ZN(G27) );
NAND4_X1 U937 ( .A1(n1265), .A2(n1060), .A3(n1268), .A4(n1255), .ZN(n1219) );
NOR2_X1 U938 ( .A1(n1069), .A2(n1077), .ZN(n1268) );
INV_X1 U939 ( .A(n1235), .ZN(n1077) );
AND3_X1 U940 ( .A1(n1089), .A2(n1269), .A3(n1270), .ZN(n1265) );
NAND2_X1 U941 ( .A1(G953), .A2(n1271), .ZN(n1270) );
NAND2_X1 U942 ( .A1(G902), .A2(n1124), .ZN(n1271) );
INV_X1 U943 ( .A(G900), .ZN(n1124) );
XOR2_X1 U944 ( .A(n1239), .B(n1272), .Z(G24) );
NOR2_X1 U945 ( .A1(KEYINPUT31), .A2(n1273), .ZN(n1272) );
AND4_X1 U946 ( .A1(n1274), .A2(n1067), .A3(n1251), .A4(n1096), .ZN(n1239) );
NOR2_X1 U947 ( .A1(n1275), .A2(n1276), .ZN(n1067) );
XNOR2_X1 U948 ( .A(G119), .B(n1240), .ZN(G21) );
NAND3_X1 U949 ( .A1(n1274), .A2(n1058), .A3(n1256), .ZN(n1240) );
AND2_X1 U950 ( .A1(n1276), .A2(n1275), .ZN(n1256) );
INV_X1 U951 ( .A(n1277), .ZN(n1276) );
NAND2_X1 U952 ( .A1(n1278), .A2(n1279), .ZN(G18) );
NAND2_X1 U953 ( .A1(G116), .A2(n1241), .ZN(n1279) );
XOR2_X1 U954 ( .A(n1280), .B(KEYINPUT4), .Z(n1278) );
OR2_X1 U955 ( .A1(n1241), .A2(G116), .ZN(n1280) );
NAND3_X1 U956 ( .A1(n1227), .A2(n1222), .A3(n1274), .ZN(n1241) );
INV_X1 U957 ( .A(n1078), .ZN(n1222) );
NAND2_X1 U958 ( .A1(n1281), .A2(n1251), .ZN(n1078) );
XNOR2_X1 U959 ( .A(n1096), .B(KEYINPUT8), .ZN(n1281) );
XOR2_X1 U960 ( .A(G113), .B(n1236), .Z(G15) );
AND3_X1 U961 ( .A1(n1227), .A2(n1235), .A3(n1274), .ZN(n1236) );
AND2_X1 U962 ( .A1(n1060), .A2(n1282), .ZN(n1274) );
INV_X1 U963 ( .A(n1088), .ZN(n1060) );
NAND2_X1 U964 ( .A1(n1084), .A2(n1283), .ZN(n1088) );
NOR2_X1 U965 ( .A1(n1277), .A2(n1275), .ZN(n1227) );
XOR2_X1 U966 ( .A(G110), .B(n1233), .Z(G12) );
AND3_X1 U967 ( .A1(n1234), .A2(n1058), .A3(n1255), .ZN(n1233) );
INV_X1 U968 ( .A(n1066), .ZN(n1255) );
NAND2_X1 U969 ( .A1(n1277), .A2(n1275), .ZN(n1066) );
XOR2_X1 U970 ( .A(n1100), .B(n1097), .Z(n1275) );
NAND2_X1 U971 ( .A1(n1151), .A2(n1210), .ZN(n1097) );
INV_X1 U972 ( .A(n1156), .ZN(n1151) );
NAND2_X1 U973 ( .A1(n1284), .A2(n1285), .ZN(n1156) );
NAND3_X1 U974 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1285) );
XOR2_X1 U975 ( .A(KEYINPUT54), .B(n1289), .Z(n1286) );
NAND2_X1 U976 ( .A1(n1290), .A2(n1291), .ZN(n1284) );
NAND2_X1 U977 ( .A1(n1288), .A2(n1287), .ZN(n1291) );
NAND2_X1 U978 ( .A1(n1292), .A2(n1293), .ZN(n1287) );
XNOR2_X1 U979 ( .A(n1294), .B(n1295), .ZN(n1293) );
XNOR2_X1 U980 ( .A(n1296), .B(n1297), .ZN(n1292) );
XOR2_X1 U981 ( .A(n1298), .B(KEYINPUT10), .Z(n1288) );
NAND2_X1 U982 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XNOR2_X1 U983 ( .A(n1301), .B(n1296), .ZN(n1300) );
XNOR2_X1 U984 ( .A(n1302), .B(n1303), .ZN(n1296) );
NOR2_X1 U985 ( .A1(KEYINPUT34), .A2(n1304), .ZN(n1303) );
NOR2_X1 U986 ( .A1(G110), .A2(KEYINPUT21), .ZN(n1302) );
XNOR2_X1 U987 ( .A(n1294), .B(n1305), .ZN(n1299) );
NOR2_X1 U988 ( .A1(KEYINPUT30), .A2(G146), .ZN(n1294) );
XOR2_X1 U989 ( .A(KEYINPUT23), .B(n1289), .Z(n1290) );
XNOR2_X1 U990 ( .A(n1306), .B(G137), .ZN(n1289) );
NAND3_X1 U991 ( .A1(G234), .A2(n1048), .A3(G221), .ZN(n1306) );
NAND2_X1 U992 ( .A1(G217), .A2(n1307), .ZN(n1100) );
XOR2_X1 U993 ( .A(n1308), .B(n1176), .Z(n1277) );
INV_X1 U994 ( .A(G472), .ZN(n1176) );
NAND2_X1 U995 ( .A1(KEYINPUT40), .A2(n1309), .ZN(n1308) );
XNOR2_X1 U996 ( .A(KEYINPUT7), .B(n1108), .ZN(n1309) );
NAND2_X1 U997 ( .A1(n1310), .A2(n1210), .ZN(n1108) );
XOR2_X1 U998 ( .A(n1311), .B(n1312), .Z(n1310) );
XOR2_X1 U999 ( .A(G101), .B(n1313), .Z(n1312) );
NOR2_X1 U1000 ( .A1(KEYINPUT24), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1001 ( .A(n1315), .B(n1126), .Z(n1314) );
NOR2_X1 U1002 ( .A1(KEYINPUT3), .A2(n1316), .ZN(n1315) );
XOR2_X1 U1003 ( .A(KEYINPUT27), .B(n1182), .Z(n1316) );
NOR2_X1 U1004 ( .A1(n1317), .A2(n1318), .ZN(n1311) );
NOR2_X1 U1005 ( .A1(KEYINPUT9), .A2(n1191), .ZN(n1318) );
INV_X1 U1006 ( .A(n1319), .ZN(n1191) );
NOR2_X1 U1007 ( .A1(KEYINPUT0), .A2(n1319), .ZN(n1317) );
NAND3_X1 U1008 ( .A1(n1320), .A2(n1048), .A3(G210), .ZN(n1319) );
NAND2_X1 U1009 ( .A1(n1321), .A2(n1322), .ZN(n1058) );
OR3_X1 U1010 ( .A1(n1251), .A2(n1096), .A3(KEYINPUT8), .ZN(n1322) );
NAND2_X1 U1011 ( .A1(KEYINPUT8), .A2(n1235), .ZN(n1321) );
NOR2_X1 U1012 ( .A1(n1323), .A2(n1251), .ZN(n1235) );
XOR2_X1 U1013 ( .A(n1110), .B(n1324), .Z(n1251) );
NOR2_X1 U1014 ( .A1(n1111), .A2(KEYINPUT13), .ZN(n1324) );
NOR2_X1 U1015 ( .A1(n1161), .A2(G902), .ZN(n1111) );
XNOR2_X1 U1016 ( .A(n1325), .B(n1326), .ZN(n1161) );
XNOR2_X1 U1017 ( .A(n1327), .B(n1328), .ZN(n1326) );
NOR2_X1 U1018 ( .A1(G107), .A2(KEYINPUT15), .ZN(n1328) );
NAND2_X1 U1019 ( .A1(n1329), .A2(KEYINPUT16), .ZN(n1327) );
XOR2_X1 U1020 ( .A(n1330), .B(G134), .Z(n1329) );
NAND2_X1 U1021 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NAND2_X1 U1022 ( .A1(G143), .A2(n1297), .ZN(n1332) );
XOR2_X1 U1023 ( .A(KEYINPUT20), .B(n1333), .Z(n1331) );
NOR2_X1 U1024 ( .A1(G143), .A2(n1297), .ZN(n1333) );
XOR2_X1 U1025 ( .A(n1334), .B(n1335), .Z(n1325) );
AND4_X1 U1026 ( .A1(n1336), .A2(n1048), .A3(G234), .A4(G217), .ZN(n1335) );
INV_X1 U1027 ( .A(KEYINPUT60), .ZN(n1336) );
XNOR2_X1 U1028 ( .A(G116), .B(G122), .ZN(n1334) );
INV_X1 U1029 ( .A(G478), .ZN(n1110) );
INV_X1 U1030 ( .A(n1096), .ZN(n1323) );
XNOR2_X1 U1031 ( .A(n1337), .B(G475), .ZN(n1096) );
OR2_X1 U1032 ( .A1(n1166), .A2(G902), .ZN(n1337) );
XNOR2_X1 U1033 ( .A(n1338), .B(n1339), .ZN(n1166) );
XOR2_X1 U1034 ( .A(G104), .B(n1340), .Z(n1339) );
NOR2_X1 U1035 ( .A1(KEYINPUT1), .A2(n1341), .ZN(n1340) );
XOR2_X1 U1036 ( .A(n1342), .B(n1343), .Z(n1341) );
XOR2_X1 U1037 ( .A(n1344), .B(n1345), .Z(n1343) );
NAND2_X1 U1038 ( .A1(KEYINPUT45), .A2(n1260), .ZN(n1345) );
INV_X1 U1039 ( .A(G131), .ZN(n1260) );
NAND2_X1 U1040 ( .A1(KEYINPUT36), .A2(n1295), .ZN(n1344) );
INV_X1 U1041 ( .A(n1305), .ZN(n1295) );
XNOR2_X1 U1042 ( .A(G140), .B(n1131), .ZN(n1305) );
XNOR2_X1 U1043 ( .A(G146), .B(n1346), .ZN(n1342) );
NAND3_X1 U1044 ( .A1(n1347), .A2(n1348), .A3(n1349), .ZN(n1346) );
NAND2_X1 U1045 ( .A1(KEYINPUT37), .A2(n1350), .ZN(n1349) );
OR3_X1 U1046 ( .A1(n1350), .A2(KEYINPUT37), .A3(G143), .ZN(n1348) );
NAND2_X1 U1047 ( .A1(G143), .A2(n1351), .ZN(n1347) );
NAND2_X1 U1048 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
INV_X1 U1049 ( .A(KEYINPUT37), .ZN(n1353) );
XNOR2_X1 U1050 ( .A(n1350), .B(KEYINPUT58), .ZN(n1352) );
AND3_X1 U1051 ( .A1(n1320), .A2(n1048), .A3(G214), .ZN(n1350) );
XNOR2_X1 U1052 ( .A(G113), .B(G122), .ZN(n1338) );
AND2_X1 U1053 ( .A1(n1282), .A2(n1266), .ZN(n1234) );
NOR2_X1 U1054 ( .A1(n1084), .A2(n1354), .ZN(n1266) );
XNOR2_X1 U1055 ( .A(KEYINPUT44), .B(n1083), .ZN(n1354) );
INV_X1 U1056 ( .A(n1283), .ZN(n1083) );
NAND2_X1 U1057 ( .A1(n1355), .A2(n1307), .ZN(n1283) );
NAND2_X1 U1058 ( .A1(G234), .A2(n1210), .ZN(n1307) );
XNOR2_X1 U1059 ( .A(G221), .B(KEYINPUT52), .ZN(n1355) );
XNOR2_X1 U1060 ( .A(n1356), .B(G469), .ZN(n1084) );
NAND2_X1 U1061 ( .A1(KEYINPUT55), .A2(n1112), .ZN(n1356) );
NAND2_X1 U1062 ( .A1(n1357), .A2(n1210), .ZN(n1112) );
XOR2_X1 U1063 ( .A(n1126), .B(n1358), .Z(n1357) );
XNOR2_X1 U1064 ( .A(n1359), .B(n1360), .ZN(n1358) );
INV_X1 U1065 ( .A(n1200), .ZN(n1360) );
NOR2_X1 U1066 ( .A1(KEYINPUT12), .A2(n1361), .ZN(n1359) );
XOR2_X1 U1067 ( .A(n1362), .B(n1363), .Z(n1361) );
XNOR2_X1 U1068 ( .A(n1364), .B(n1365), .ZN(n1363) );
NOR2_X1 U1069 ( .A1(KEYINPUT18), .A2(n1203), .ZN(n1365) );
NAND2_X1 U1070 ( .A1(G227), .A2(n1048), .ZN(n1203) );
NAND2_X1 U1071 ( .A1(KEYINPUT28), .A2(n1198), .ZN(n1364) );
INV_X1 U1072 ( .A(G140), .ZN(n1198) );
XNOR2_X1 U1073 ( .A(G110), .B(KEYINPUT43), .ZN(n1362) );
XOR2_X1 U1074 ( .A(n1186), .B(n1366), .Z(n1126) );
XOR2_X1 U1075 ( .A(G131), .B(n1367), .Z(n1186) );
XOR2_X1 U1076 ( .A(G137), .B(G134), .Z(n1367) );
AND4_X1 U1077 ( .A1(n1252), .A2(n1368), .A3(n1089), .A4(n1269), .ZN(n1282) );
OR2_X1 U1078 ( .A1(G953), .A2(G952), .ZN(n1269) );
NAND2_X1 U1079 ( .A1(G237), .A2(G234), .ZN(n1089) );
NAND2_X1 U1080 ( .A1(G953), .A2(n1369), .ZN(n1368) );
NAND2_X1 U1081 ( .A1(G902), .A2(n1141), .ZN(n1369) );
INV_X1 U1082 ( .A(G898), .ZN(n1141) );
INV_X1 U1083 ( .A(n1069), .ZN(n1252) );
NAND2_X1 U1084 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NAND2_X1 U1085 ( .A1(G214), .A2(n1370), .ZN(n1072) );
XNOR2_X1 U1086 ( .A(n1107), .B(n1106), .ZN(n1071) );
NAND2_X1 U1087 ( .A1(G210), .A2(n1370), .ZN(n1106) );
NAND2_X1 U1088 ( .A1(n1320), .A2(n1210), .ZN(n1370) );
INV_X1 U1089 ( .A(G237), .ZN(n1320) );
INV_X1 U1090 ( .A(n1104), .ZN(n1107) );
NAND2_X1 U1091 ( .A1(n1371), .A2(n1210), .ZN(n1104) );
INV_X1 U1092 ( .A(G902), .ZN(n1210) );
XOR2_X1 U1093 ( .A(n1206), .B(n1372), .Z(n1371) );
NOR4_X1 U1094 ( .A1(n1373), .A2(n1374), .A3(KEYINPUT47), .A4(n1243), .ZN(n1372) );
AND2_X1 U1095 ( .A1(n1248), .A2(n1246), .ZN(n1243) );
NOR2_X1 U1096 ( .A1(n1187), .A2(G125), .ZN(n1248) );
INV_X1 U1097 ( .A(n1366), .ZN(n1187) );
NOR3_X1 U1098 ( .A1(G125), .A2(n1366), .A3(n1246), .ZN(n1374) );
NOR2_X1 U1099 ( .A1(n1375), .A2(n1131), .ZN(n1373) );
INV_X1 U1100 ( .A(G125), .ZN(n1131) );
XNOR2_X1 U1101 ( .A(n1246), .B(n1366), .ZN(n1375) );
XOR2_X1 U1102 ( .A(n1376), .B(n1297), .Z(n1366) );
INV_X1 U1103 ( .A(n1301), .ZN(n1297) );
XOR2_X1 U1104 ( .A(G128), .B(KEYINPUT59), .Z(n1301) );
XNOR2_X1 U1105 ( .A(G146), .B(G143), .ZN(n1376) );
NAND2_X1 U1106 ( .A1(G224), .A2(n1048), .ZN(n1246) );
INV_X1 U1107 ( .A(G953), .ZN(n1048) );
XNOR2_X1 U1108 ( .A(n1144), .B(n1377), .ZN(n1206) );
NOR2_X1 U1109 ( .A1(KEYINPUT46), .A2(n1143), .ZN(n1377) );
XNOR2_X1 U1110 ( .A(n1182), .B(n1200), .ZN(n1143) );
XOR2_X1 U1111 ( .A(G101), .B(n1378), .Z(n1200) );
XOR2_X1 U1112 ( .A(G107), .B(G104), .Z(n1378) );
XOR2_X1 U1113 ( .A(G113), .B(n1379), .Z(n1182) );
XNOR2_X1 U1114 ( .A(n1304), .B(G116), .ZN(n1379) );
INV_X1 U1115 ( .A(G119), .ZN(n1304) );
XNOR2_X1 U1116 ( .A(G110), .B(n1273), .ZN(n1144) );
INV_X1 U1117 ( .A(G122), .ZN(n1273) );
endmodule


