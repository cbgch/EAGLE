//Key = 1001100011001001111100001011110111010101000001000000011100001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366;

XNOR2_X1 U753 ( .A(n1044), .B(n1045), .ZN(G9) );
XNOR2_X1 U754 ( .A(G107), .B(KEYINPUT51), .ZN(n1045) );
NOR2_X1 U755 ( .A1(n1046), .A2(n1047), .ZN(G75) );
NOR4_X1 U756 ( .A1(n1048), .A2(n1049), .A3(G953), .A4(n1050), .ZN(n1047) );
NOR2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR3_X1 U759 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NOR3_X1 U760 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1056) );
NOR2_X1 U761 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U762 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U763 ( .A1(n1065), .A2(n1066), .ZN(n1059) );
XNOR2_X1 U764 ( .A(n1067), .B(KEYINPUT20), .ZN(n1065) );
AND2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1058) );
NOR3_X1 U766 ( .A1(n1062), .A2(n1069), .A3(n1070), .ZN(n1053) );
NOR2_X1 U767 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR2_X1 U768 ( .A1(n1073), .A2(n1055), .ZN(n1072) );
NOR2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U771 ( .A1(n1078), .A2(n1057), .ZN(n1071) );
NOR2_X1 U772 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U773 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
INV_X1 U774 ( .A(n1083), .ZN(n1062) );
INV_X1 U775 ( .A(n1084), .ZN(n1051) );
NAND2_X1 U776 ( .A1(n1085), .A2(G952), .ZN(n1048) );
NOR3_X1 U777 ( .A1(n1086), .A2(G953), .A3(n1050), .ZN(n1046) );
AND3_X1 U778 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1050) );
NOR3_X1 U779 ( .A1(n1090), .A2(n1091), .A3(n1070), .ZN(n1089) );
XNOR2_X1 U780 ( .A(n1092), .B(n1093), .ZN(n1091) );
NOR2_X1 U781 ( .A1(G475), .A2(KEYINPUT50), .ZN(n1093) );
XOR2_X1 U782 ( .A(KEYINPUT36), .B(G952), .Z(n1086) );
XOR2_X1 U783 ( .A(n1094), .B(n1095), .Z(G72) );
NOR2_X1 U784 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U785 ( .A(KEYINPUT1), .B(n1098), .Z(n1097) );
AND2_X1 U786 ( .A1(G227), .A2(G900), .ZN(n1098) );
NAND2_X1 U787 ( .A1(n1099), .A2(n1100), .ZN(n1094) );
NAND2_X1 U788 ( .A1(n1101), .A2(n1096), .ZN(n1100) );
XOR2_X1 U789 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND3_X1 U790 ( .A1(G900), .A2(n1103), .A3(G953), .ZN(n1099) );
XOR2_X1 U791 ( .A(n1104), .B(n1105), .Z(n1103) );
XNOR2_X1 U792 ( .A(n1106), .B(n1107), .ZN(n1104) );
NOR2_X1 U793 ( .A1(KEYINPUT7), .A2(n1108), .ZN(n1107) );
XOR2_X1 U794 ( .A(n1109), .B(n1110), .Z(n1108) );
XNOR2_X1 U795 ( .A(n1111), .B(G131), .ZN(n1110) );
NOR2_X1 U796 ( .A1(KEYINPUT41), .A2(n1112), .ZN(n1109) );
XOR2_X1 U797 ( .A(n1113), .B(n1114), .Z(G69) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U799 ( .A(n1117), .B(KEYINPUT0), .Z(n1116) );
OR3_X1 U800 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1117) );
INV_X1 U801 ( .A(n1121), .ZN(n1118) );
NOR2_X1 U802 ( .A1(n1122), .A2(n1121), .ZN(n1115) );
NAND2_X1 U803 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
NAND2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XNOR2_X1 U805 ( .A(KEYINPUT17), .B(n1127), .ZN(n1126) );
INV_X1 U806 ( .A(n1128), .ZN(n1125) );
XNOR2_X1 U807 ( .A(G953), .B(KEYINPUT34), .ZN(n1123) );
NOR2_X1 U808 ( .A1(n1119), .A2(n1120), .ZN(n1122) );
XNOR2_X1 U809 ( .A(n1129), .B(n1130), .ZN(n1120) );
NOR3_X1 U810 ( .A1(KEYINPUT47), .A2(n1131), .A3(n1132), .ZN(n1130) );
NOR3_X1 U811 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
INV_X1 U812 ( .A(KEYINPUT30), .ZN(n1133) );
NOR2_X1 U813 ( .A1(KEYINPUT30), .A2(n1136), .ZN(n1131) );
NAND2_X1 U814 ( .A1(G953), .A2(n1137), .ZN(n1113) );
NAND2_X1 U815 ( .A1(G898), .A2(G224), .ZN(n1137) );
NOR2_X1 U816 ( .A1(n1138), .A2(n1139), .ZN(G66) );
XOR2_X1 U817 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND3_X1 U818 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1140) );
XNOR2_X1 U819 ( .A(G217), .B(KEYINPUT15), .ZN(n1144) );
NOR2_X1 U820 ( .A1(n1138), .A2(n1145), .ZN(G63) );
NOR2_X1 U821 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U822 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U823 ( .A1(KEYINPUT33), .A2(n1150), .ZN(n1149) );
NAND2_X1 U824 ( .A1(n1142), .A2(G478), .ZN(n1148) );
NOR2_X1 U825 ( .A1(KEYINPUT33), .A2(n1150), .ZN(n1146) );
NOR2_X1 U826 ( .A1(n1138), .A2(n1151), .ZN(G60) );
NOR3_X1 U827 ( .A1(n1092), .A2(n1152), .A3(n1153), .ZN(n1151) );
AND3_X1 U828 ( .A1(n1154), .A2(G475), .A3(n1142), .ZN(n1153) );
NOR2_X1 U829 ( .A1(n1155), .A2(n1154), .ZN(n1152) );
NOR2_X1 U830 ( .A1(n1085), .A2(n1156), .ZN(n1155) );
NAND2_X1 U831 ( .A1(n1157), .A2(n1158), .ZN(G6) );
NAND2_X1 U832 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U833 ( .A(KEYINPUT39), .B(n1161), .Z(n1157) );
NOR2_X1 U834 ( .A1(n1159), .A2(n1160), .ZN(n1161) );
INV_X1 U835 ( .A(n1162), .ZN(n1159) );
NOR3_X1 U836 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(G57) );
AND3_X1 U837 ( .A1(KEYINPUT14), .A2(G953), .A3(G952), .ZN(n1165) );
NOR2_X1 U838 ( .A1(KEYINPUT14), .A2(n1166), .ZN(n1164) );
INV_X1 U839 ( .A(n1138), .ZN(n1166) );
NOR2_X1 U840 ( .A1(n1167), .A2(n1168), .ZN(n1163) );
XOR2_X1 U841 ( .A(KEYINPUT10), .B(n1169), .Z(n1168) );
NOR2_X1 U842 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XNOR2_X1 U843 ( .A(n1172), .B(n1173), .ZN(n1171) );
INV_X1 U844 ( .A(n1174), .ZN(n1170) );
NOR2_X1 U845 ( .A1(n1175), .A2(n1174), .ZN(n1167) );
XOR2_X1 U846 ( .A(n1176), .B(n1177), .Z(n1174) );
XNOR2_X1 U847 ( .A(n1173), .B(n1178), .ZN(n1175) );
INV_X1 U848 ( .A(n1172), .ZN(n1178) );
XOR2_X1 U849 ( .A(n1179), .B(n1180), .Z(n1173) );
NOR2_X1 U850 ( .A1(KEYINPUT56), .A2(n1181), .ZN(n1180) );
NAND2_X1 U851 ( .A1(n1142), .A2(G472), .ZN(n1179) );
NOR2_X1 U852 ( .A1(n1138), .A2(n1182), .ZN(G54) );
XNOR2_X1 U853 ( .A(n1183), .B(n1184), .ZN(n1182) );
XOR2_X1 U854 ( .A(n1185), .B(n1186), .Z(n1183) );
NOR2_X1 U855 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U856 ( .A(n1189), .B(KEYINPUT26), .Z(n1188) );
NAND2_X1 U857 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U858 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
NAND2_X1 U859 ( .A1(n1142), .A2(n1192), .ZN(n1185) );
XOR2_X1 U860 ( .A(KEYINPUT5), .B(G469), .Z(n1192) );
NOR2_X1 U861 ( .A1(n1138), .A2(n1193), .ZN(G51) );
XOR2_X1 U862 ( .A(n1194), .B(n1195), .Z(n1193) );
NAND2_X1 U863 ( .A1(n1142), .A2(n1196), .ZN(n1195) );
NOR2_X1 U864 ( .A1(n1197), .A2(n1085), .ZN(n1142) );
NOR3_X1 U865 ( .A1(n1128), .A2(n1044), .A3(n1102), .ZN(n1085) );
NAND4_X1 U866 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1102) );
NOR4_X1 U867 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
NAND2_X1 U868 ( .A1(n1075), .A2(n1206), .ZN(n1200) );
NAND2_X1 U869 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND3_X1 U870 ( .A1(n1090), .A2(n1209), .A3(n1210), .ZN(n1208) );
XNOR2_X1 U871 ( .A(n1211), .B(KEYINPUT57), .ZN(n1207) );
NAND4_X1 U872 ( .A1(n1212), .A2(n1064), .A3(n1213), .A4(n1088), .ZN(n1198) );
INV_X1 U873 ( .A(n1127), .ZN(n1044) );
NAND3_X1 U874 ( .A1(n1068), .A2(n1067), .A3(n1214), .ZN(n1127) );
NAND4_X1 U875 ( .A1(n1215), .A2(n1162), .A3(n1216), .A4(n1217), .ZN(n1128) );
AND4_X1 U876 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1217) );
OR2_X1 U877 ( .A1(n1222), .A2(n1223), .ZN(n1216) );
NAND3_X1 U878 ( .A1(n1214), .A2(n1067), .A3(n1213), .ZN(n1162) );
NAND3_X1 U879 ( .A1(n1063), .A2(n1213), .A3(n1224), .ZN(n1215) );
NAND2_X1 U880 ( .A1(n1225), .A2(n1226), .ZN(n1194) );
NAND2_X1 U881 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
XOR2_X1 U882 ( .A(KEYINPUT28), .B(n1229), .Z(n1225) );
NOR2_X1 U883 ( .A1(n1228), .A2(n1227), .ZN(n1229) );
XNOR2_X1 U884 ( .A(KEYINPUT48), .B(n1230), .ZN(n1227) );
NOR2_X1 U885 ( .A1(n1096), .A2(G952), .ZN(n1138) );
XNOR2_X1 U886 ( .A(G146), .B(n1231), .ZN(G48) );
NAND3_X1 U887 ( .A1(n1211), .A2(n1075), .A3(KEYINPUT29), .ZN(n1231) );
AND2_X1 U888 ( .A1(n1232), .A2(n1213), .ZN(n1211) );
XNOR2_X1 U889 ( .A(G143), .B(n1233), .ZN(G45) );
NAND4_X1 U890 ( .A1(n1210), .A2(n1234), .A3(n1090), .A4(n1209), .ZN(n1233) );
XNOR2_X1 U891 ( .A(KEYINPUT6), .B(n1223), .ZN(n1234) );
XOR2_X1 U892 ( .A(n1235), .B(n1236), .Z(G42) );
XNOR2_X1 U893 ( .A(G140), .B(KEYINPUT46), .ZN(n1236) );
NAND4_X1 U894 ( .A1(n1064), .A2(n1213), .A3(KEYINPUT53), .A4(n1237), .ZN(n1235) );
NOR3_X1 U895 ( .A1(n1057), .A2(n1238), .A3(n1239), .ZN(n1237) );
XNOR2_X1 U896 ( .A(n1080), .B(KEYINPUT2), .ZN(n1239) );
NAND2_X1 U897 ( .A1(n1240), .A2(n1241), .ZN(G39) );
NAND2_X1 U898 ( .A1(n1242), .A2(n1199), .ZN(n1241) );
NAND2_X1 U899 ( .A1(n1111), .A2(n1243), .ZN(n1242) );
NAND2_X1 U900 ( .A1(KEYINPUT63), .A2(n1244), .ZN(n1243) );
NAND3_X1 U901 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1240) );
INV_X1 U902 ( .A(KEYINPUT63), .ZN(n1247) );
NAND2_X1 U903 ( .A1(G137), .A2(n1244), .ZN(n1246) );
INV_X1 U904 ( .A(KEYINPUT21), .ZN(n1244) );
NAND2_X1 U905 ( .A1(n1248), .A2(n1111), .ZN(n1245) );
OR2_X1 U906 ( .A1(n1199), .A2(KEYINPUT21), .ZN(n1248) );
NAND3_X1 U907 ( .A1(n1232), .A2(n1088), .A3(n1083), .ZN(n1199) );
XOR2_X1 U908 ( .A(n1203), .B(n1249), .Z(G36) );
NOR2_X1 U909 ( .A1(KEYINPUT42), .A2(n1112), .ZN(n1249) );
INV_X1 U910 ( .A(G134), .ZN(n1112) );
AND3_X1 U911 ( .A1(n1088), .A2(n1068), .A3(n1210), .ZN(n1203) );
XNOR2_X1 U912 ( .A(n1250), .B(n1205), .ZN(G33) );
AND3_X1 U913 ( .A1(n1213), .A2(n1088), .A3(n1210), .ZN(n1205) );
AND2_X1 U914 ( .A1(n1212), .A2(n1063), .ZN(n1210) );
INV_X1 U915 ( .A(n1057), .ZN(n1088) );
NAND2_X1 U916 ( .A1(n1251), .A2(n1077), .ZN(n1057) );
INV_X1 U917 ( .A(n1076), .ZN(n1251) );
XNOR2_X1 U918 ( .A(n1252), .B(n1204), .ZN(G30) );
AND3_X1 U919 ( .A1(n1068), .A2(n1075), .A3(n1232), .ZN(n1204) );
AND3_X1 U920 ( .A1(n1253), .A2(n1254), .A3(n1212), .ZN(n1232) );
NOR2_X1 U921 ( .A1(n1255), .A2(n1238), .ZN(n1212) );
XNOR2_X1 U922 ( .A(G101), .B(n1221), .ZN(G3) );
NAND3_X1 U923 ( .A1(n1063), .A2(n1214), .A3(n1083), .ZN(n1221) );
XOR2_X1 U924 ( .A(n1202), .B(n1256), .Z(G27) );
NOR2_X1 U925 ( .A1(KEYINPUT11), .A2(n1257), .ZN(n1256) );
AND4_X1 U926 ( .A1(n1064), .A2(n1213), .A3(n1258), .A4(n1087), .ZN(n1202) );
NOR2_X1 U927 ( .A1(n1238), .A2(n1223), .ZN(n1258) );
AND2_X1 U928 ( .A1(n1259), .A2(n1260), .ZN(n1238) );
NAND4_X1 U929 ( .A1(n1261), .A2(G953), .A3(n1084), .A4(n1262), .ZN(n1260) );
INV_X1 U930 ( .A(G900), .ZN(n1262) );
NAND2_X1 U931 ( .A1(n1263), .A2(n1264), .ZN(G24) );
OR2_X1 U932 ( .A1(n1265), .A2(G122), .ZN(n1264) );
NAND2_X1 U933 ( .A1(n1266), .A2(G122), .ZN(n1263) );
NAND2_X1 U934 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
OR2_X1 U935 ( .A1(n1220), .A2(KEYINPUT31), .ZN(n1268) );
INV_X1 U936 ( .A(n1269), .ZN(n1220) );
NAND2_X1 U937 ( .A1(KEYINPUT31), .A2(n1265), .ZN(n1267) );
NAND2_X1 U938 ( .A1(KEYINPUT37), .A2(n1269), .ZN(n1265) );
NOR4_X1 U939 ( .A1(n1270), .A2(n1070), .A3(n1271), .A4(n1272), .ZN(n1269) );
INV_X1 U940 ( .A(n1067), .ZN(n1070) );
NOR2_X1 U941 ( .A1(n1254), .A2(n1253), .ZN(n1067) );
XNOR2_X1 U942 ( .A(G119), .B(n1219), .ZN(G21) );
NAND4_X1 U943 ( .A1(n1224), .A2(n1083), .A3(n1253), .A4(n1254), .ZN(n1219) );
INV_X1 U944 ( .A(n1270), .ZN(n1224) );
XNOR2_X1 U945 ( .A(G116), .B(n1273), .ZN(G18) );
NAND2_X1 U946 ( .A1(n1274), .A2(n1075), .ZN(n1273) );
XOR2_X1 U947 ( .A(n1222), .B(KEYINPUT16), .Z(n1274) );
NAND4_X1 U948 ( .A1(n1063), .A2(n1087), .A3(n1068), .A4(n1275), .ZN(n1222) );
NOR2_X1 U949 ( .A1(n1209), .A2(n1271), .ZN(n1068) );
INV_X1 U950 ( .A(n1090), .ZN(n1271) );
XOR2_X1 U951 ( .A(G113), .B(n1276), .Z(G15) );
NOR4_X1 U952 ( .A1(KEYINPUT58), .A2(n1066), .A3(n1277), .A4(n1270), .ZN(n1276) );
NAND3_X1 U953 ( .A1(n1075), .A2(n1275), .A3(n1087), .ZN(n1270) );
INV_X1 U954 ( .A(n1055), .ZN(n1087) );
NAND2_X1 U955 ( .A1(n1278), .A2(n1082), .ZN(n1055) );
INV_X1 U956 ( .A(n1081), .ZN(n1278) );
INV_X1 U957 ( .A(n1063), .ZN(n1277) );
NOR2_X1 U958 ( .A1(n1253), .A2(n1279), .ZN(n1063) );
INV_X1 U959 ( .A(n1213), .ZN(n1066) );
NOR2_X1 U960 ( .A1(n1090), .A2(n1272), .ZN(n1213) );
INV_X1 U961 ( .A(n1209), .ZN(n1272) );
XNOR2_X1 U962 ( .A(G110), .B(n1218), .ZN(G12) );
NAND3_X1 U963 ( .A1(n1064), .A2(n1214), .A3(n1083), .ZN(n1218) );
NOR2_X1 U964 ( .A1(n1090), .A2(n1209), .ZN(n1083) );
NAND3_X1 U965 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1209) );
OR2_X1 U966 ( .A1(n1156), .A2(KEYINPUT9), .ZN(n1282) );
NAND3_X1 U967 ( .A1(KEYINPUT9), .A2(n1156), .A3(n1092), .ZN(n1281) );
NAND2_X1 U968 ( .A1(n1283), .A2(n1284), .ZN(n1280) );
INV_X1 U969 ( .A(n1092), .ZN(n1284) );
NOR2_X1 U970 ( .A1(n1154), .A2(G902), .ZN(n1092) );
XOR2_X1 U971 ( .A(n1285), .B(n1286), .Z(n1154) );
XOR2_X1 U972 ( .A(n1287), .B(n1288), .Z(n1286) );
XNOR2_X1 U973 ( .A(G113), .B(n1160), .ZN(n1288) );
XNOR2_X1 U974 ( .A(G143), .B(n1289), .ZN(n1287) );
XNOR2_X1 U975 ( .A(n1290), .B(n1291), .ZN(n1285) );
INV_X1 U976 ( .A(n1106), .ZN(n1291) );
XOR2_X1 U977 ( .A(n1292), .B(n1293), .Z(n1290) );
AND3_X1 U978 ( .A1(G214), .A2(n1096), .A3(n1294), .ZN(n1293) );
NAND2_X1 U979 ( .A1(KEYINPUT8), .A2(n1250), .ZN(n1292) );
INV_X1 U980 ( .A(G131), .ZN(n1250) );
NAND2_X1 U981 ( .A1(KEYINPUT9), .A2(n1295), .ZN(n1283) );
XNOR2_X1 U982 ( .A(KEYINPUT19), .B(n1156), .ZN(n1295) );
INV_X1 U983 ( .A(G475), .ZN(n1156) );
XNOR2_X1 U984 ( .A(n1296), .B(G478), .ZN(n1090) );
NAND2_X1 U985 ( .A1(n1150), .A2(n1197), .ZN(n1296) );
XOR2_X1 U986 ( .A(n1297), .B(n1298), .Z(n1150) );
XNOR2_X1 U987 ( .A(G107), .B(n1299), .ZN(n1298) );
NAND2_X1 U988 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NAND2_X1 U989 ( .A1(G116), .A2(n1289), .ZN(n1301) );
XOR2_X1 U990 ( .A(KEYINPUT18), .B(n1302), .Z(n1300) );
NOR2_X1 U991 ( .A1(G116), .A2(n1289), .ZN(n1302) );
NAND2_X1 U992 ( .A1(n1303), .A2(n1304), .ZN(n1297) );
NAND2_X1 U993 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
INV_X1 U994 ( .A(n1307), .ZN(n1306) );
XOR2_X1 U995 ( .A(KEYINPUT24), .B(n1308), .Z(n1305) );
NAND2_X1 U996 ( .A1(n1309), .A2(n1307), .ZN(n1303) );
XOR2_X1 U997 ( .A(G128), .B(n1310), .Z(n1307) );
XOR2_X1 U998 ( .A(KEYINPUT44), .B(G143), .Z(n1310) );
XOR2_X1 U999 ( .A(KEYINPUT49), .B(n1308), .Z(n1309) );
XNOR2_X1 U1000 ( .A(n1311), .B(G134), .ZN(n1308) );
NAND3_X1 U1001 ( .A1(G234), .A2(n1096), .A3(G217), .ZN(n1311) );
AND3_X1 U1002 ( .A1(n1075), .A2(n1275), .A3(n1080), .ZN(n1214) );
INV_X1 U1003 ( .A(n1255), .ZN(n1080) );
NAND2_X1 U1004 ( .A1(n1081), .A2(n1082), .ZN(n1255) );
NAND2_X1 U1005 ( .A1(G221), .A2(n1143), .ZN(n1082) );
NAND2_X1 U1006 ( .A1(G234), .A2(n1312), .ZN(n1143) );
XNOR2_X1 U1007 ( .A(n1313), .B(G469), .ZN(n1081) );
NAND2_X1 U1008 ( .A1(n1314), .A2(n1197), .ZN(n1313) );
XOR2_X1 U1009 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1010 ( .A(n1317), .B(KEYINPUT62), .ZN(n1316) );
NAND2_X1 U1011 ( .A1(KEYINPUT61), .A2(n1184), .ZN(n1317) );
XOR2_X1 U1012 ( .A(n1318), .B(n1319), .Z(n1184) );
XOR2_X1 U1013 ( .A(n1320), .B(n1321), .Z(n1319) );
XNOR2_X1 U1014 ( .A(KEYINPUT40), .B(n1322), .ZN(n1321) );
NOR2_X1 U1015 ( .A1(KEYINPUT59), .A2(n1177), .ZN(n1322) );
XNOR2_X1 U1016 ( .A(n1323), .B(n1105), .ZN(n1318) );
XNOR2_X1 U1017 ( .A(n1324), .B(n1325), .ZN(n1105) );
NOR2_X1 U1018 ( .A1(G143), .A2(KEYINPUT22), .ZN(n1325) );
NAND2_X1 U1019 ( .A1(KEYINPUT4), .A2(n1252), .ZN(n1324) );
XNOR2_X1 U1020 ( .A(n1190), .B(n1191), .ZN(n1315) );
NAND2_X1 U1021 ( .A1(G227), .A2(n1096), .ZN(n1191) );
XNOR2_X1 U1022 ( .A(G110), .B(n1326), .ZN(n1190) );
NAND2_X1 U1023 ( .A1(n1259), .A2(n1327), .ZN(n1275) );
NAND3_X1 U1024 ( .A1(n1261), .A2(n1084), .A3(n1119), .ZN(n1327) );
NOR2_X1 U1025 ( .A1(n1096), .A2(G898), .ZN(n1119) );
XNOR2_X1 U1026 ( .A(G902), .B(KEYINPUT54), .ZN(n1261) );
NAND3_X1 U1027 ( .A1(n1084), .A2(n1096), .A3(G952), .ZN(n1259) );
NAND2_X1 U1028 ( .A1(n1328), .A2(G237), .ZN(n1084) );
XNOR2_X1 U1029 ( .A(G234), .B(KEYINPUT55), .ZN(n1328) );
INV_X1 U1030 ( .A(n1223), .ZN(n1075) );
NAND2_X1 U1031 ( .A1(n1076), .A2(n1077), .ZN(n1223) );
NAND2_X1 U1032 ( .A1(G214), .A2(n1329), .ZN(n1077) );
XNOR2_X1 U1033 ( .A(n1330), .B(n1196), .ZN(n1076) );
AND2_X1 U1034 ( .A1(G210), .A2(n1329), .ZN(n1196) );
NAND2_X1 U1035 ( .A1(n1312), .A2(n1294), .ZN(n1329) );
NAND2_X1 U1036 ( .A1(n1331), .A2(n1197), .ZN(n1330) );
XOR2_X1 U1037 ( .A(n1228), .B(n1230), .Z(n1331) );
XNOR2_X1 U1038 ( .A(n1129), .B(n1136), .ZN(n1230) );
XNOR2_X1 U1039 ( .A(n1135), .B(n1134), .ZN(n1136) );
XNOR2_X1 U1040 ( .A(n1332), .B(n1333), .ZN(n1134) );
NAND2_X1 U1041 ( .A1(KEYINPUT12), .A2(n1334), .ZN(n1332) );
XNOR2_X1 U1042 ( .A(G101), .B(n1323), .ZN(n1135) );
XNOR2_X1 U1043 ( .A(G107), .B(n1160), .ZN(n1323) );
INV_X1 U1044 ( .A(G104), .ZN(n1160) );
XNOR2_X1 U1045 ( .A(n1335), .B(n1289), .ZN(n1129) );
INV_X1 U1046 ( .A(G122), .ZN(n1289) );
NAND2_X1 U1047 ( .A1(KEYINPUT3), .A2(n1336), .ZN(n1335) );
INV_X1 U1048 ( .A(G110), .ZN(n1336) );
XOR2_X1 U1049 ( .A(n1337), .B(n1338), .Z(n1228) );
XOR2_X1 U1050 ( .A(n1339), .B(n1340), .Z(n1337) );
NAND2_X1 U1051 ( .A1(G224), .A2(n1096), .ZN(n1339) );
AND2_X1 U1052 ( .A1(n1279), .A2(n1253), .ZN(n1064) );
XNOR2_X1 U1053 ( .A(n1341), .B(n1342), .ZN(n1253) );
NOR2_X1 U1054 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
INV_X1 U1055 ( .A(G217), .ZN(n1344) );
AND2_X1 U1056 ( .A1(n1312), .A2(G234), .ZN(n1343) );
XOR2_X1 U1057 ( .A(G902), .B(KEYINPUT35), .Z(n1312) );
NAND2_X1 U1058 ( .A1(n1141), .A2(n1197), .ZN(n1341) );
XNOR2_X1 U1059 ( .A(n1345), .B(n1106), .ZN(n1141) );
XOR2_X1 U1060 ( .A(n1326), .B(n1340), .Z(n1106) );
XNOR2_X1 U1061 ( .A(n1257), .B(G146), .ZN(n1340) );
INV_X1 U1062 ( .A(G125), .ZN(n1257) );
XOR2_X1 U1063 ( .A(G140), .B(KEYINPUT60), .Z(n1326) );
XNOR2_X1 U1064 ( .A(n1346), .B(n1347), .ZN(n1345) );
NOR2_X1 U1065 ( .A1(KEYINPUT13), .A2(n1348), .ZN(n1347) );
XOR2_X1 U1066 ( .A(n1349), .B(n1350), .Z(n1348) );
XNOR2_X1 U1067 ( .A(G119), .B(G110), .ZN(n1350) );
NAND2_X1 U1068 ( .A1(KEYINPUT45), .A2(n1252), .ZN(n1349) );
NOR2_X1 U1069 ( .A1(KEYINPUT43), .A2(n1351), .ZN(n1346) );
XNOR2_X1 U1070 ( .A(n1111), .B(n1352), .ZN(n1351) );
AND3_X1 U1071 ( .A1(G221), .A2(n1096), .A3(G234), .ZN(n1352) );
INV_X1 U1072 ( .A(n1254), .ZN(n1279) );
XNOR2_X1 U1073 ( .A(n1353), .B(G472), .ZN(n1254) );
NAND2_X1 U1074 ( .A1(n1354), .A2(n1197), .ZN(n1353) );
INV_X1 U1075 ( .A(G902), .ZN(n1197) );
XNOR2_X1 U1076 ( .A(n1172), .B(n1355), .ZN(n1354) );
XOR2_X1 U1077 ( .A(n1356), .B(n1181), .Z(n1355) );
XNOR2_X1 U1078 ( .A(n1320), .B(n1338), .ZN(n1181) );
XNOR2_X1 U1079 ( .A(n1357), .B(G143), .ZN(n1338) );
NAND2_X1 U1080 ( .A1(KEYINPUT27), .A2(n1252), .ZN(n1357) );
INV_X1 U1081 ( .A(G128), .ZN(n1252) );
XOR2_X1 U1082 ( .A(n1358), .B(n1359), .Z(n1320) );
NOR2_X1 U1083 ( .A1(KEYINPUT25), .A2(n1360), .ZN(n1359) );
XNOR2_X1 U1084 ( .A(n1111), .B(G134), .ZN(n1360) );
INV_X1 U1085 ( .A(G137), .ZN(n1111) );
XNOR2_X1 U1086 ( .A(G146), .B(G131), .ZN(n1358) );
NAND3_X1 U1087 ( .A1(n1361), .A2(n1362), .A3(n1363), .ZN(n1356) );
NAND2_X1 U1088 ( .A1(KEYINPUT23), .A2(n1176), .ZN(n1363) );
NAND3_X1 U1089 ( .A1(n1364), .A2(n1365), .A3(n1177), .ZN(n1362) );
INV_X1 U1090 ( .A(KEYINPUT23), .ZN(n1365) );
OR2_X1 U1091 ( .A1(n1177), .A2(n1364), .ZN(n1361) );
NOR2_X1 U1092 ( .A1(KEYINPUT52), .A2(n1176), .ZN(n1364) );
NAND3_X1 U1093 ( .A1(n1294), .A2(n1096), .A3(G210), .ZN(n1176) );
INV_X1 U1094 ( .A(G953), .ZN(n1096) );
INV_X1 U1095 ( .A(G237), .ZN(n1294) );
INV_X1 U1096 ( .A(G101), .ZN(n1177) );
XOR2_X1 U1097 ( .A(n1334), .B(n1366), .Z(n1172) );
XOR2_X1 U1098 ( .A(KEYINPUT38), .B(n1333), .Z(n1366) );
XOR2_X1 U1099 ( .A(G113), .B(G119), .Z(n1333) );
XOR2_X1 U1100 ( .A(G116), .B(KEYINPUT32), .Z(n1334) );
endmodule


