//Key = 1011110010111100110000100111000100100000011111001001110110111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309;

XNOR2_X1 U723 ( .A(G107), .B(n999), .ZN(G9) );
NOR2_X1 U724 ( .A1(n1000), .A2(n1001), .ZN(G75) );
NOR4_X1 U725 ( .A1(G953), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n1001) );
NOR2_X1 U726 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
NOR2_X1 U727 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR3_X1 U728 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1008) );
NOR2_X1 U729 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR2_X1 U730 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NOR2_X1 U731 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR2_X1 U732 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NOR2_X1 U733 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR2_X1 U734 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U735 ( .A1(n1024), .A2(n1025), .ZN(n1016) );
NOR2_X1 U736 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U737 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NOR3_X1 U738 ( .A1(n1019), .A2(n1030), .A3(n1025), .ZN(n1012) );
NOR2_X1 U739 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR4_X1 U740 ( .A1(n1033), .A2(n1025), .A3(n1019), .A4(n1015), .ZN(n1007) );
INV_X1 U741 ( .A(n1034), .ZN(n1025) );
NOR2_X1 U742 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U743 ( .A1(n1009), .A2(n1037), .ZN(n1035) );
NOR3_X1 U744 ( .A1(n1002), .A2(G953), .A3(G952), .ZN(n1000) );
AND4_X1 U745 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1002) );
NOR3_X1 U746 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
XOR2_X1 U747 ( .A(KEYINPUT46), .B(n1045), .Z(n1044) );
XOR2_X1 U748 ( .A(G475), .B(n1046), .Z(n1043) );
NAND4_X1 U749 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1042) );
NAND3_X1 U750 ( .A1(G478), .A2(n1051), .A3(n1052), .ZN(n1050) );
OR2_X1 U751 ( .A1(n1052), .A2(G478), .ZN(n1049) );
INV_X1 U752 ( .A(KEYINPUT50), .ZN(n1052) );
OR2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(n1048) );
NAND2_X1 U754 ( .A1(n1055), .A2(n1053), .ZN(n1047) );
XOR2_X1 U755 ( .A(KEYINPUT32), .B(n1054), .Z(n1055) );
NOR3_X1 U756 ( .A1(n1010), .A2(n1056), .A3(n1057), .ZN(n1040) );
XNOR2_X1 U757 ( .A(n1058), .B(n1059), .ZN(n1039) );
NOR2_X1 U758 ( .A1(G472), .A2(KEYINPUT20), .ZN(n1059) );
XNOR2_X1 U759 ( .A(n1060), .B(n1061), .ZN(n1038) );
XOR2_X1 U760 ( .A(n1062), .B(n1063), .Z(G72) );
XOR2_X1 U761 ( .A(n1064), .B(n1065), .Z(n1063) );
NOR2_X1 U762 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
AND2_X1 U763 ( .A1(G227), .A2(G900), .ZN(n1066) );
NAND2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1064) );
NAND2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
XOR2_X1 U766 ( .A(n1072), .B(n1073), .Z(n1068) );
XNOR2_X1 U767 ( .A(n1074), .B(n1075), .ZN(n1073) );
NOR2_X1 U768 ( .A1(KEYINPUT14), .A2(n1076), .ZN(n1075) );
XNOR2_X1 U769 ( .A(n1077), .B(n1078), .ZN(n1072) );
NAND2_X1 U770 ( .A1(n1067), .A2(n1079), .ZN(n1062) );
XOR2_X1 U771 ( .A(n1080), .B(n1081), .Z(G69) );
XOR2_X1 U772 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XOR2_X1 U774 ( .A(n1086), .B(n1087), .Z(n1085) );
AND2_X1 U775 ( .A1(n1088), .A2(n1070), .ZN(n1084) );
NAND2_X1 U776 ( .A1(n1067), .A2(n1089), .ZN(n1082) );
NAND3_X1 U777 ( .A1(n1090), .A2(n999), .A3(n1091), .ZN(n1089) );
XOR2_X1 U778 ( .A(n1092), .B(KEYINPUT47), .Z(n1091) );
NAND2_X1 U779 ( .A1(G953), .A2(n1093), .ZN(n1080) );
NAND2_X1 U780 ( .A1(G898), .A2(G224), .ZN(n1093) );
NOR2_X1 U781 ( .A1(n1094), .A2(n1095), .ZN(G66) );
NOR2_X1 U782 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U783 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U784 ( .A1(n1053), .A2(n1100), .ZN(n1099) );
NOR2_X1 U785 ( .A1(KEYINPUT62), .A2(n1101), .ZN(n1098) );
XNOR2_X1 U786 ( .A(KEYINPUT59), .B(n1102), .ZN(n1101) );
NOR2_X1 U787 ( .A1(n1103), .A2(n1104), .ZN(n1096) );
INV_X1 U788 ( .A(KEYINPUT62), .ZN(n1104) );
XOR2_X1 U789 ( .A(n1102), .B(KEYINPUT59), .Z(n1103) );
NOR2_X1 U790 ( .A1(n1094), .A2(n1105), .ZN(G63) );
XOR2_X1 U791 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U792 ( .A1(n1100), .A2(n1108), .ZN(n1106) );
XOR2_X1 U793 ( .A(KEYINPUT48), .B(G478), .Z(n1108) );
NOR2_X1 U794 ( .A1(n1094), .A2(n1109), .ZN(G60) );
NOR3_X1 U795 ( .A1(n1046), .A2(n1110), .A3(n1111), .ZN(n1109) );
NOR3_X1 U796 ( .A1(n1112), .A2(n1113), .A3(n1100), .ZN(n1111) );
INV_X1 U797 ( .A(n1114), .ZN(n1112) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1114), .ZN(n1110) );
NOR2_X1 U799 ( .A1(n1116), .A2(n1113), .ZN(n1115) );
XNOR2_X1 U800 ( .A(G475), .B(KEYINPUT24), .ZN(n1113) );
INV_X1 U801 ( .A(n1004), .ZN(n1116) );
XNOR2_X1 U802 ( .A(G104), .B(n1117), .ZN(G6) );
NOR2_X1 U803 ( .A1(n1094), .A2(n1118), .ZN(G57) );
XOR2_X1 U804 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U805 ( .A(n1121), .B(n1122), .Z(n1120) );
XNOR2_X1 U806 ( .A(n1123), .B(n1124), .ZN(n1122) );
NOR2_X1 U807 ( .A1(KEYINPUT15), .A2(n1125), .ZN(n1124) );
NAND2_X1 U808 ( .A1(KEYINPUT2), .A2(n1126), .ZN(n1123) );
NOR2_X1 U809 ( .A1(n1127), .A2(n1100), .ZN(n1121) );
XOR2_X1 U810 ( .A(n1128), .B(n1129), .Z(n1119) );
NOR2_X1 U811 ( .A1(n1094), .A2(n1130), .ZN(G54) );
XOR2_X1 U812 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U813 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U814 ( .A1(n1135), .A2(n1100), .ZN(n1133) );
XOR2_X1 U815 ( .A(n1136), .B(n1137), .Z(n1131) );
XNOR2_X1 U816 ( .A(KEYINPUT19), .B(n1138), .ZN(n1137) );
NAND2_X1 U817 ( .A1(KEYINPUT26), .A2(n1139), .ZN(n1136) );
NOR2_X1 U818 ( .A1(n1094), .A2(n1140), .ZN(G51) );
XOR2_X1 U819 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U820 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR3_X1 U821 ( .A1(n1100), .A2(KEYINPUT49), .A3(n1145), .ZN(n1144) );
INV_X1 U822 ( .A(G210), .ZN(n1145) );
NAND2_X1 U823 ( .A1(G902), .A2(n1004), .ZN(n1100) );
NAND4_X1 U824 ( .A1(n1146), .A2(n1147), .A3(n1090), .A4(n1092), .ZN(n1004) );
AND4_X1 U825 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1090) );
AND3_X1 U826 ( .A1(n1117), .A2(n1152), .A3(n1153), .ZN(n1151) );
NAND3_X1 U827 ( .A1(n1154), .A2(n1034), .A3(n1032), .ZN(n1117) );
INV_X1 U828 ( .A(n1079), .ZN(n1147) );
NAND4_X1 U829 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1079) );
AND4_X1 U830 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1158) );
NAND2_X1 U831 ( .A1(n1032), .A2(n1163), .ZN(n1157) );
NAND2_X1 U832 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U833 ( .A1(n1166), .A2(n1021), .ZN(n1165) );
OR2_X1 U834 ( .A1(n1167), .A2(n1168), .ZN(n1164) );
NAND4_X1 U835 ( .A1(n1031), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1155) );
NAND2_X1 U836 ( .A1(KEYINPUT13), .A2(n1167), .ZN(n1171) );
NAND2_X1 U837 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
INV_X1 U838 ( .A(KEYINPUT13), .ZN(n1173) );
NAND2_X1 U839 ( .A1(n1174), .A2(n1175), .ZN(n1172) );
XOR2_X1 U840 ( .A(n999), .B(KEYINPUT40), .Z(n1146) );
NAND3_X1 U841 ( .A1(n1031), .A2(n1034), .A3(n1154), .ZN(n999) );
XOR2_X1 U842 ( .A(n1176), .B(n1177), .Z(n1141) );
NOR2_X1 U843 ( .A1(KEYINPUT33), .A2(n1178), .ZN(n1177) );
XOR2_X1 U844 ( .A(n1179), .B(KEYINPUT41), .Z(n1176) );
NOR2_X1 U845 ( .A1(n1067), .A2(G952), .ZN(n1094) );
XOR2_X1 U846 ( .A(G146), .B(n1180), .Z(G48) );
NOR3_X1 U847 ( .A1(n1167), .A2(n1181), .A3(n1182), .ZN(n1180) );
XNOR2_X1 U848 ( .A(n1168), .B(KEYINPUT10), .ZN(n1181) );
NAND2_X1 U849 ( .A1(n1183), .A2(n1184), .ZN(G45) );
OR2_X1 U850 ( .A1(n1156), .A2(G143), .ZN(n1184) );
XOR2_X1 U851 ( .A(n1185), .B(KEYINPUT9), .Z(n1183) );
NAND2_X1 U852 ( .A1(G143), .A2(n1156), .ZN(n1185) );
NAND4_X1 U853 ( .A1(n1021), .A2(n1036), .A3(n1186), .A4(n1187), .ZN(n1156) );
NOR3_X1 U854 ( .A1(n1175), .A2(n1188), .A3(n1168), .ZN(n1187) );
XOR2_X1 U855 ( .A(n1162), .B(n1189), .Z(G42) );
NAND2_X1 U856 ( .A1(KEYINPUT25), .A2(G140), .ZN(n1189) );
NAND2_X1 U857 ( .A1(n1166), .A2(n1190), .ZN(n1162) );
XNOR2_X1 U858 ( .A(G137), .B(n1161), .ZN(G39) );
NAND2_X1 U859 ( .A1(n1191), .A2(n1166), .ZN(n1161) );
NAND2_X1 U860 ( .A1(n1192), .A2(n1193), .ZN(G36) );
NAND2_X1 U861 ( .A1(G134), .A2(n1160), .ZN(n1193) );
XOR2_X1 U862 ( .A(KEYINPUT11), .B(n1194), .Z(n1192) );
NOR2_X1 U863 ( .A1(G134), .A2(n1160), .ZN(n1194) );
NAND3_X1 U864 ( .A1(n1021), .A2(n1031), .A3(n1166), .ZN(n1160) );
NOR4_X1 U865 ( .A1(n1009), .A2(n1175), .A3(n1168), .A4(n1010), .ZN(n1166) );
INV_X1 U866 ( .A(n1027), .ZN(n1175) );
XOR2_X1 U867 ( .A(n1195), .B(n1196), .Z(G33) );
NAND2_X1 U868 ( .A1(KEYINPUT45), .A2(G131), .ZN(n1196) );
NAND4_X1 U869 ( .A1(n1021), .A2(n1027), .A3(n1032), .A4(n1197), .ZN(n1195) );
NOR3_X1 U870 ( .A1(n1009), .A2(n1010), .A3(n1198), .ZN(n1197) );
XNOR2_X1 U871 ( .A(n1168), .B(KEYINPUT4), .ZN(n1198) );
INV_X1 U872 ( .A(n1037), .ZN(n1010) );
XOR2_X1 U873 ( .A(G128), .B(n1199), .Z(G30) );
NOR4_X1 U874 ( .A1(KEYINPUT29), .A2(n1168), .A3(n1200), .A4(n1167), .ZN(n1199) );
NAND2_X1 U875 ( .A1(n1174), .A2(n1027), .ZN(n1167) );
NOR3_X1 U876 ( .A1(n1201), .A2(n1022), .A3(n1202), .ZN(n1174) );
INV_X1 U877 ( .A(n1169), .ZN(n1168) );
XNOR2_X1 U878 ( .A(G101), .B(n1203), .ZN(G3) );
NAND2_X1 U879 ( .A1(KEYINPUT17), .A2(n1204), .ZN(n1203) );
INV_X1 U880 ( .A(n1153), .ZN(n1204) );
NAND3_X1 U881 ( .A1(n1021), .A2(n1154), .A3(n1205), .ZN(n1153) );
XNOR2_X1 U882 ( .A(G125), .B(n1159), .ZN(G27) );
NAND4_X1 U883 ( .A1(n1190), .A2(n1206), .A3(n1036), .A4(n1169), .ZN(n1159) );
NAND2_X1 U884 ( .A1(n1006), .A2(n1207), .ZN(n1169) );
NAND4_X1 U885 ( .A1(G902), .A2(n1070), .A3(n1208), .A4(n1071), .ZN(n1207) );
INV_X1 U886 ( .A(G900), .ZN(n1071) );
NOR3_X1 U887 ( .A1(n1023), .A2(n1022), .A3(n1182), .ZN(n1190) );
XNOR2_X1 U888 ( .A(G122), .B(n1152), .ZN(G24) );
NAND4_X1 U889 ( .A1(n1186), .A2(n1209), .A3(n1034), .A4(n1210), .ZN(n1152) );
NOR2_X1 U890 ( .A1(n1211), .A2(n1023), .ZN(n1034) );
XOR2_X1 U891 ( .A(G119), .B(n1212), .Z(G21) );
NOR3_X1 U892 ( .A1(KEYINPUT18), .A2(n1213), .A3(n1214), .ZN(n1212) );
NOR2_X1 U893 ( .A1(KEYINPUT8), .A2(n1215), .ZN(n1214) );
NOR4_X1 U894 ( .A1(n1202), .A2(n1019), .A3(n1216), .A4(n1217), .ZN(n1215) );
INV_X1 U895 ( .A(n1191), .ZN(n1216) );
INV_X1 U896 ( .A(n1206), .ZN(n1019) );
AND2_X1 U897 ( .A1(n1150), .A2(KEYINPUT8), .ZN(n1213) );
NAND2_X1 U898 ( .A1(n1191), .A2(n1209), .ZN(n1150) );
NOR3_X1 U899 ( .A1(n1201), .A2(n1022), .A3(n1015), .ZN(n1191) );
NAND2_X1 U900 ( .A1(n1218), .A2(n1219), .ZN(G18) );
NAND2_X1 U901 ( .A1(G116), .A2(n1092), .ZN(n1219) );
XOR2_X1 U902 ( .A(KEYINPUT27), .B(n1220), .Z(n1218) );
NOR2_X1 U903 ( .A1(G116), .A2(n1092), .ZN(n1220) );
NAND3_X1 U904 ( .A1(n1209), .A2(n1031), .A3(n1021), .ZN(n1092) );
INV_X1 U905 ( .A(n1200), .ZN(n1031) );
NAND2_X1 U906 ( .A1(n1221), .A2(n1210), .ZN(n1200) );
INV_X1 U907 ( .A(n1188), .ZN(n1210) );
XNOR2_X1 U908 ( .A(n1148), .B(n1222), .ZN(G15) );
NOR2_X1 U909 ( .A1(KEYINPUT6), .A2(n1223), .ZN(n1222) );
INV_X1 U910 ( .A(G113), .ZN(n1223) );
NAND3_X1 U911 ( .A1(n1021), .A2(n1209), .A3(n1032), .ZN(n1148) );
INV_X1 U912 ( .A(n1182), .ZN(n1032) );
NAND2_X1 U913 ( .A1(n1188), .A2(n1186), .ZN(n1182) );
XOR2_X1 U914 ( .A(n1224), .B(KEYINPUT35), .Z(n1186) );
AND3_X1 U915 ( .A1(n1036), .A2(n1217), .A3(n1206), .ZN(n1209) );
NOR2_X1 U916 ( .A1(n1028), .A2(n1056), .ZN(n1206) );
NOR2_X1 U917 ( .A1(n1211), .A2(n1201), .ZN(n1021) );
XNOR2_X1 U918 ( .A(G110), .B(n1149), .ZN(G12) );
NAND4_X1 U919 ( .A1(n1205), .A2(n1154), .A3(n1201), .A4(n1211), .ZN(n1149) );
INV_X1 U920 ( .A(n1022), .ZN(n1211) );
XOR2_X1 U921 ( .A(n1054), .B(n1053), .Z(n1022) );
NAND2_X1 U922 ( .A1(G217), .A2(n1225), .ZN(n1053) );
NOR2_X1 U923 ( .A1(n1102), .A2(G902), .ZN(n1054) );
XOR2_X1 U924 ( .A(n1226), .B(n1227), .Z(n1102) );
XNOR2_X1 U925 ( .A(KEYINPUT31), .B(n1074), .ZN(n1227) );
XOR2_X1 U926 ( .A(n1228), .B(n1229), .Z(n1226) );
NOR2_X1 U927 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
INV_X1 U928 ( .A(G221), .ZN(n1230) );
NAND2_X1 U929 ( .A1(n1232), .A2(n1233), .ZN(n1228) );
NAND2_X1 U930 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U931 ( .A(KEYINPUT60), .B(n1236), .Z(n1232) );
NOR2_X1 U932 ( .A1(n1235), .A2(n1234), .ZN(n1236) );
XOR2_X1 U933 ( .A(n1237), .B(G110), .Z(n1234) );
NAND2_X1 U934 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND2_X1 U935 ( .A1(G128), .A2(n1240), .ZN(n1239) );
XOR2_X1 U936 ( .A(n1241), .B(KEYINPUT61), .Z(n1238) );
OR2_X1 U937 ( .A1(n1240), .A2(G128), .ZN(n1241) );
INV_X1 U938 ( .A(n1023), .ZN(n1201) );
XOR2_X1 U939 ( .A(n1058), .B(n1127), .Z(n1023) );
INV_X1 U940 ( .A(G472), .ZN(n1127) );
NAND2_X1 U941 ( .A1(n1242), .A2(n1243), .ZN(n1058) );
XOR2_X1 U942 ( .A(n1244), .B(n1245), .Z(n1242) );
XOR2_X1 U943 ( .A(n1246), .B(n1125), .Z(n1245) );
NOR2_X1 U944 ( .A1(KEYINPUT57), .A2(n1129), .ZN(n1246) );
XNOR2_X1 U945 ( .A(n1128), .B(n1126), .ZN(n1244) );
XOR2_X1 U946 ( .A(n1247), .B(G101), .Z(n1128) );
NAND3_X1 U947 ( .A1(n1248), .A2(n1249), .A3(G210), .ZN(n1247) );
AND3_X1 U948 ( .A1(n1027), .A2(n1217), .A3(n1036), .ZN(n1154) );
INV_X1 U949 ( .A(n1202), .ZN(n1036) );
NAND2_X1 U950 ( .A1(n1250), .A2(n1037), .ZN(n1202) );
NAND2_X1 U951 ( .A1(G214), .A2(n1251), .ZN(n1037) );
XOR2_X1 U952 ( .A(KEYINPUT54), .B(n1009), .Z(n1250) );
XNOR2_X1 U953 ( .A(n1252), .B(n1061), .ZN(n1009) );
AND2_X1 U954 ( .A1(G210), .A2(n1251), .ZN(n1061) );
NAND2_X1 U955 ( .A1(n1249), .A2(n1243), .ZN(n1251) );
NAND2_X1 U956 ( .A1(KEYINPUT52), .A2(n1060), .ZN(n1252) );
AND2_X1 U957 ( .A1(n1253), .A2(n1243), .ZN(n1060) );
XOR2_X1 U958 ( .A(n1178), .B(n1254), .Z(n1253) );
XOR2_X1 U959 ( .A(n1255), .B(KEYINPUT5), .Z(n1254) );
NAND2_X1 U960 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND2_X1 U961 ( .A1(KEYINPUT30), .A2(n1143), .ZN(n1257) );
XNOR2_X1 U962 ( .A(n1258), .B(n1179), .ZN(n1256) );
NAND2_X1 U963 ( .A1(G224), .A2(n1248), .ZN(n1179) );
OR2_X1 U964 ( .A1(n1143), .A2(KEYINPUT30), .ZN(n1258) );
XNOR2_X1 U965 ( .A(n1125), .B(G125), .ZN(n1143) );
XOR2_X1 U966 ( .A(n1259), .B(n1260), .Z(n1125) );
NAND2_X1 U967 ( .A1(KEYINPUT43), .A2(n1261), .ZN(n1259) );
XOR2_X1 U968 ( .A(n1262), .B(n1087), .Z(n1178) );
XOR2_X1 U969 ( .A(G110), .B(G122), .Z(n1087) );
NAND2_X1 U970 ( .A1(KEYINPUT56), .A2(n1086), .ZN(n1262) );
XNOR2_X1 U971 ( .A(n1263), .B(n1126), .ZN(n1086) );
XOR2_X1 U972 ( .A(n1264), .B(n1240), .Z(n1126) );
XOR2_X1 U973 ( .A(G119), .B(KEYINPUT22), .Z(n1240) );
XNOR2_X1 U974 ( .A(G113), .B(G116), .ZN(n1264) );
NAND2_X1 U975 ( .A1(n1265), .A2(n1266), .ZN(n1217) );
NAND4_X1 U976 ( .A1(G902), .A2(n1070), .A3(n1208), .A4(n1088), .ZN(n1266) );
INV_X1 U977 ( .A(G898), .ZN(n1088) );
XOR2_X1 U978 ( .A(G953), .B(KEYINPUT37), .Z(n1070) );
XOR2_X1 U979 ( .A(n1006), .B(KEYINPUT36), .Z(n1265) );
NAND3_X1 U980 ( .A1(n1208), .A2(n1067), .A3(G952), .ZN(n1006) );
NAND2_X1 U981 ( .A1(G237), .A2(n1267), .ZN(n1208) );
NOR2_X1 U982 ( .A1(n1268), .A2(n1056), .ZN(n1027) );
INV_X1 U983 ( .A(n1029), .ZN(n1056) );
NAND2_X1 U984 ( .A1(G221), .A2(n1225), .ZN(n1029) );
NAND2_X1 U985 ( .A1(n1267), .A2(n1243), .ZN(n1225) );
XNOR2_X1 U986 ( .A(G234), .B(KEYINPUT12), .ZN(n1267) );
INV_X1 U987 ( .A(n1028), .ZN(n1268) );
XOR2_X1 U988 ( .A(n1045), .B(KEYINPUT7), .Z(n1028) );
XOR2_X1 U989 ( .A(n1269), .B(n1135), .Z(n1045) );
INV_X1 U990 ( .A(G469), .ZN(n1135) );
NAND2_X1 U991 ( .A1(n1270), .A2(n1243), .ZN(n1269) );
INV_X1 U992 ( .A(G902), .ZN(n1243) );
XOR2_X1 U993 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U994 ( .A(KEYINPUT53), .B(n1273), .Z(n1272) );
NOR2_X1 U995 ( .A1(KEYINPUT39), .A2(n1138), .ZN(n1273) );
NAND2_X1 U996 ( .A1(G227), .A2(n1248), .ZN(n1138) );
XNOR2_X1 U997 ( .A(n1139), .B(n1134), .ZN(n1271) );
XOR2_X1 U998 ( .A(n1129), .B(n1274), .Z(n1134) );
XOR2_X1 U999 ( .A(G140), .B(G110), .Z(n1274) );
XNOR2_X1 U1000 ( .A(n1275), .B(n1077), .ZN(n1129) );
XNOR2_X1 U1001 ( .A(G131), .B(n1276), .ZN(n1077) );
NAND2_X1 U1002 ( .A1(n1277), .A2(n1074), .ZN(n1275) );
INV_X1 U1003 ( .A(G137), .ZN(n1074) );
XNOR2_X1 U1004 ( .A(KEYINPUT55), .B(KEYINPUT3), .ZN(n1277) );
XNOR2_X1 U1005 ( .A(n1263), .B(n1078), .ZN(n1139) );
XOR2_X1 U1006 ( .A(n1260), .B(n1261), .Z(n1078) );
XNOR2_X1 U1007 ( .A(G128), .B(KEYINPUT44), .ZN(n1261) );
XNOR2_X1 U1008 ( .A(G146), .B(G143), .ZN(n1260) );
XNOR2_X1 U1009 ( .A(G101), .B(n1278), .ZN(n1263) );
XNOR2_X1 U1010 ( .A(G107), .B(n1279), .ZN(n1278) );
INV_X1 U1011 ( .A(n1015), .ZN(n1205) );
NAND2_X1 U1012 ( .A1(n1188), .A2(n1221), .ZN(n1015) );
XNOR2_X1 U1013 ( .A(n1224), .B(KEYINPUT21), .ZN(n1221) );
NAND2_X1 U1014 ( .A1(n1280), .A2(n1281), .ZN(n1224) );
NAND2_X1 U1015 ( .A1(G475), .A2(n1282), .ZN(n1281) );
XOR2_X1 U1016 ( .A(KEYINPUT0), .B(n1283), .Z(n1280) );
NOR2_X1 U1017 ( .A1(G475), .A2(n1282), .ZN(n1283) );
XOR2_X1 U1018 ( .A(KEYINPUT42), .B(n1046), .Z(n1282) );
NOR2_X1 U1019 ( .A1(n1114), .A2(G902), .ZN(n1046) );
XOR2_X1 U1020 ( .A(n1284), .B(n1235), .Z(n1114) );
XNOR2_X1 U1021 ( .A(G146), .B(n1076), .ZN(n1235) );
XOR2_X1 U1022 ( .A(G125), .B(G140), .Z(n1076) );
XOR2_X1 U1023 ( .A(n1285), .B(n1286), .Z(n1284) );
NOR2_X1 U1024 ( .A1(KEYINPUT28), .A2(n1287), .ZN(n1286) );
XNOR2_X1 U1025 ( .A(G131), .B(n1288), .ZN(n1287) );
NAND2_X1 U1026 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
NAND4_X1 U1027 ( .A1(G143), .A2(G214), .A3(n1248), .A4(n1249), .ZN(n1290) );
NAND2_X1 U1028 ( .A1(n1291), .A2(n1292), .ZN(n1289) );
NAND3_X1 U1029 ( .A1(n1248), .A2(n1249), .A3(G214), .ZN(n1292) );
INV_X1 U1030 ( .A(G237), .ZN(n1249) );
XOR2_X1 U1031 ( .A(KEYINPUT58), .B(G143), .Z(n1291) );
NAND2_X1 U1032 ( .A1(n1293), .A2(n1294), .ZN(n1285) );
NAND2_X1 U1033 ( .A1(n1295), .A2(n1279), .ZN(n1294) );
XOR2_X1 U1034 ( .A(n1296), .B(KEYINPUT1), .Z(n1293) );
OR2_X1 U1035 ( .A1(n1295), .A2(n1279), .ZN(n1296) );
INV_X1 U1036 ( .A(G104), .ZN(n1279) );
XOR2_X1 U1037 ( .A(G113), .B(n1297), .Z(n1295) );
XOR2_X1 U1038 ( .A(KEYINPUT16), .B(G122), .Z(n1297) );
NOR2_X1 U1039 ( .A1(n1057), .A2(n1298), .ZN(n1188) );
AND2_X1 U1040 ( .A1(G478), .A2(n1051), .ZN(n1298) );
NOR2_X1 U1041 ( .A1(n1051), .A2(G478), .ZN(n1057) );
OR2_X1 U1042 ( .A1(n1107), .A2(G902), .ZN(n1051) );
XNOR2_X1 U1043 ( .A(n1299), .B(n1300), .ZN(n1107) );
XOR2_X1 U1044 ( .A(n1301), .B(n1302), .Z(n1300) );
XNOR2_X1 U1045 ( .A(G116), .B(G122), .ZN(n1302) );
NAND2_X1 U1046 ( .A1(KEYINPUT34), .A2(n1303), .ZN(n1301) );
XOR2_X1 U1047 ( .A(n1304), .B(n1305), .Z(n1303) );
XNOR2_X1 U1048 ( .A(G128), .B(G143), .ZN(n1305) );
NAND2_X1 U1049 ( .A1(KEYINPUT63), .A2(n1276), .ZN(n1304) );
INV_X1 U1050 ( .A(G134), .ZN(n1276) );
XNOR2_X1 U1051 ( .A(n1306), .B(n1307), .ZN(n1299) );
NOR2_X1 U1052 ( .A1(n1308), .A2(KEYINPUT23), .ZN(n1307) );
NOR2_X1 U1053 ( .A1(n1231), .A2(n1309), .ZN(n1308) );
INV_X1 U1054 ( .A(G217), .ZN(n1309) );
NAND2_X1 U1055 ( .A1(G234), .A2(n1248), .ZN(n1231) );
XNOR2_X1 U1056 ( .A(n1067), .B(KEYINPUT51), .ZN(n1248) );
INV_X1 U1057 ( .A(G953), .ZN(n1067) );
NOR2_X1 U1058 ( .A1(G107), .A2(KEYINPUT38), .ZN(n1306) );
endmodule


