//Key = 0011101001011100011111100000011110010101101100011100110101001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347;

XNOR2_X1 U730 ( .A(n1013), .B(n1014), .ZN(G9) );
NOR2_X1 U731 ( .A1(n1015), .A2(n1016), .ZN(G75) );
NOR4_X1 U732 ( .A1(G953), .A2(n1017), .A3(n1018), .A4(n1019), .ZN(n1016) );
NOR2_X1 U733 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR2_X1 U734 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR3_X1 U735 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
NOR3_X1 U736 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1025) );
NOR3_X1 U737 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
XNOR2_X1 U738 ( .A(KEYINPUT20), .B(n1033), .ZN(n1030) );
NOR2_X1 U739 ( .A1(n1034), .A2(n1035), .ZN(n1027) );
NOR3_X1 U740 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1034) );
NOR3_X1 U741 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
INV_X1 U742 ( .A(KEYINPUT42), .ZN(n1039) );
NOR2_X1 U743 ( .A1(KEYINPUT42), .A2(n1033), .ZN(n1037) );
XNOR2_X1 U744 ( .A(KEYINPUT24), .B(n1042), .ZN(n1036) );
NOR3_X1 U745 ( .A1(n1035), .A2(n1043), .A3(n1033), .ZN(n1022) );
NOR3_X1 U746 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NOR2_X1 U747 ( .A1(n1047), .A2(n1026), .ZN(n1046) );
NOR2_X1 U748 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
INV_X1 U749 ( .A(n1050), .ZN(n1045) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1024), .ZN(n1044) );
INV_X1 U751 ( .A(n1052), .ZN(n1035) );
NOR3_X1 U752 ( .A1(n1017), .A2(G953), .A3(G952), .ZN(n1015) );
AND4_X1 U753 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1017) );
NOR4_X1 U754 ( .A1(n1057), .A2(n1058), .A3(n1033), .A4(n1059), .ZN(n1056) );
XOR2_X1 U755 ( .A(n1060), .B(n1061), .Z(n1059) );
NOR3_X1 U756 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1055) );
NOR2_X1 U757 ( .A1(n1065), .A2(n1066), .ZN(n1062) );
INV_X1 U758 ( .A(G478), .ZN(n1066) );
NOR2_X1 U759 ( .A1(G902), .A2(n1067), .ZN(n1065) );
NAND2_X1 U760 ( .A1(G472), .A2(n1068), .ZN(n1054) );
XOR2_X1 U761 ( .A(KEYINPUT32), .B(n1069), .Z(n1053) );
XOR2_X1 U762 ( .A(n1070), .B(n1071), .Z(G72) );
NOR2_X1 U763 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U764 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XOR2_X1 U765 ( .A(n1076), .B(KEYINPUT61), .Z(n1075) );
NAND2_X1 U766 ( .A1(G900), .A2(G227), .ZN(n1076) );
NOR3_X1 U767 ( .A1(G953), .A2(KEYINPUT50), .A3(n1077), .ZN(n1072) );
NOR2_X1 U768 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(n1070) );
NAND2_X1 U770 ( .A1(G953), .A2(n1082), .ZN(n1081) );
XOR2_X1 U771 ( .A(n1083), .B(KEYINPUT21), .Z(n1080) );
NAND2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U773 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U774 ( .A(n1088), .B(KEYINPUT48), .Z(n1087) );
XNOR2_X1 U775 ( .A(KEYINPUT56), .B(n1089), .ZN(n1086) );
NAND2_X1 U776 ( .A1(n1090), .A2(n1091), .ZN(n1084) );
XOR2_X1 U777 ( .A(n1088), .B(KEYINPUT58), .Z(n1091) );
XOR2_X1 U778 ( .A(n1092), .B(n1093), .Z(n1088) );
NOR2_X1 U779 ( .A1(KEYINPUT14), .A2(n1094), .ZN(n1093) );
XNOR2_X1 U780 ( .A(G131), .B(n1095), .ZN(n1094) );
NOR2_X1 U781 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U782 ( .A1(KEYINPUT13), .A2(n1098), .ZN(n1097) );
NOR2_X1 U783 ( .A1(KEYINPUT28), .A2(n1099), .ZN(n1096) );
INV_X1 U784 ( .A(n1098), .ZN(n1099) );
XOR2_X1 U785 ( .A(KEYINPUT56), .B(n1089), .Z(n1090) );
XOR2_X1 U786 ( .A(n1100), .B(n1101), .Z(G69) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U788 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XNOR2_X1 U789 ( .A(G953), .B(KEYINPUT54), .ZN(n1105) );
NOR2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NAND2_X1 U791 ( .A1(n1108), .A2(n1109), .ZN(n1102) );
NAND2_X1 U792 ( .A1(G953), .A2(n1107), .ZN(n1109) );
XOR2_X1 U793 ( .A(n1110), .B(n1111), .Z(n1108) );
NAND3_X1 U794 ( .A1(n1112), .A2(n1074), .A3(KEYINPUT55), .ZN(n1100) );
NOR2_X1 U795 ( .A1(n1113), .A2(n1114), .ZN(G66) );
XNOR2_X1 U796 ( .A(n1115), .B(n1116), .ZN(n1114) );
NOR2_X1 U797 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NOR2_X1 U798 ( .A1(n1119), .A2(n1120), .ZN(G63) );
XNOR2_X1 U799 ( .A(n1121), .B(n1067), .ZN(n1120) );
NAND3_X1 U800 ( .A1(n1122), .A2(n1123), .A3(G478), .ZN(n1121) );
NAND2_X1 U801 ( .A1(KEYINPUT30), .A2(n1118), .ZN(n1123) );
NAND2_X1 U802 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
INV_X1 U803 ( .A(KEYINPUT30), .ZN(n1125) );
NAND2_X1 U804 ( .A1(n1126), .A2(G902), .ZN(n1124) );
XOR2_X1 U805 ( .A(KEYINPUT10), .B(n1113), .Z(n1119) );
NOR2_X1 U806 ( .A1(n1113), .A2(n1127), .ZN(G60) );
XOR2_X1 U807 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U808 ( .A1(n1130), .A2(n1118), .ZN(n1128) );
XNOR2_X1 U809 ( .A(n1131), .B(n1132), .ZN(G6) );
NOR2_X1 U810 ( .A1(n1113), .A2(n1133), .ZN(G57) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U812 ( .A(n1136), .B(n1137), .Z(n1135) );
NOR2_X1 U813 ( .A1(n1138), .A2(n1118), .ZN(n1137) );
INV_X1 U814 ( .A(G472), .ZN(n1138) );
NOR2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
XOR2_X1 U816 ( .A(KEYINPUT5), .B(n1141), .Z(n1140) );
NOR2_X1 U817 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
AND2_X1 U818 ( .A1(n1143), .A2(n1142), .ZN(n1139) );
XNOR2_X1 U819 ( .A(n1144), .B(n1145), .ZN(n1134) );
NOR2_X1 U820 ( .A1(n1113), .A2(n1146), .ZN(G54) );
XOR2_X1 U821 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U822 ( .A(n1149), .B(n1150), .Z(n1148) );
NAND2_X1 U823 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
XOR2_X1 U824 ( .A(n1153), .B(KEYINPUT34), .Z(n1151) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1147) );
NOR2_X1 U826 ( .A1(KEYINPUT25), .A2(G140), .ZN(n1155) );
XNOR2_X1 U827 ( .A(G110), .B(n1156), .ZN(n1154) );
NOR2_X1 U828 ( .A1(n1157), .A2(n1118), .ZN(n1156) );
XNOR2_X1 U829 ( .A(G469), .B(KEYINPUT36), .ZN(n1157) );
NOR2_X1 U830 ( .A1(n1113), .A2(n1158), .ZN(G51) );
XOR2_X1 U831 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U832 ( .A(G125), .B(n1161), .Z(n1160) );
NOR2_X1 U833 ( .A1(n1162), .A2(KEYINPUT44), .ZN(n1161) );
NOR2_X1 U834 ( .A1(n1061), .A2(n1118), .ZN(n1162) );
NAND2_X1 U835 ( .A1(G902), .A2(n1019), .ZN(n1118) );
INV_X1 U836 ( .A(n1126), .ZN(n1019) );
NOR3_X1 U837 ( .A1(n1079), .A2(n1112), .A3(n1163), .ZN(n1126) );
XOR2_X1 U838 ( .A(KEYINPUT59), .B(n1078), .Z(n1163) );
NAND2_X1 U839 ( .A1(n1164), .A2(n1165), .ZN(n1078) );
NAND4_X1 U840 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
AND3_X1 U841 ( .A1(n1170), .A2(n1171), .A3(n1058), .ZN(n1168) );
NOR2_X1 U842 ( .A1(n1172), .A2(n1051), .ZN(n1166) );
OR2_X1 U843 ( .A1(n1173), .A2(n1169), .ZN(n1164) );
INV_X1 U844 ( .A(KEYINPUT18), .ZN(n1169) );
NAND4_X1 U845 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1112) );
NOR4_X1 U846 ( .A1(n1178), .A2(n1132), .A3(n1179), .A4(n1180), .ZN(n1177) );
NOR2_X1 U847 ( .A1(n1181), .A2(n1050), .ZN(n1180) );
NOR3_X1 U848 ( .A1(n1182), .A2(n1183), .A3(n1051), .ZN(n1179) );
NOR3_X1 U849 ( .A1(n1026), .A2(n1181), .A3(n1184), .ZN(n1132) );
NOR2_X1 U850 ( .A1(n1014), .A2(n1185), .ZN(n1176) );
NOR3_X1 U851 ( .A1(n1026), .A2(n1181), .A3(n1183), .ZN(n1014) );
NAND4_X1 U852 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1079) );
NOR4_X1 U853 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
NAND3_X1 U854 ( .A1(n1052), .A2(n1194), .A3(n1195), .ZN(n1188) );
NOR2_X1 U855 ( .A1(n1074), .A2(G952), .ZN(n1113) );
XNOR2_X1 U856 ( .A(G146), .B(n1186), .ZN(G48) );
NAND3_X1 U857 ( .A1(n1049), .A2(n1196), .A3(n1194), .ZN(n1186) );
INV_X1 U858 ( .A(n1197), .ZN(n1194) );
XOR2_X1 U859 ( .A(n1173), .B(n1198), .Z(G45) );
NOR2_X1 U860 ( .A1(G143), .A2(KEYINPUT23), .ZN(n1198) );
NAND4_X1 U861 ( .A1(n1199), .A2(n1196), .A3(n1058), .A4(n1171), .ZN(n1173) );
XNOR2_X1 U862 ( .A(G140), .B(n1187), .ZN(G42) );
NAND3_X1 U863 ( .A1(n1200), .A2(n1170), .A3(n1052), .ZN(n1187) );
XOR2_X1 U864 ( .A(G137), .B(n1201), .Z(G39) );
NOR3_X1 U865 ( .A1(n1024), .A2(n1202), .A3(n1197), .ZN(n1201) );
XNOR2_X1 U866 ( .A(n1052), .B(KEYINPUT51), .ZN(n1202) );
XNOR2_X1 U867 ( .A(n1203), .B(n1193), .ZN(G36) );
AND3_X1 U868 ( .A1(n1199), .A2(n1048), .A3(n1052), .ZN(n1193) );
XNOR2_X1 U869 ( .A(n1204), .B(n1192), .ZN(G33) );
AND3_X1 U870 ( .A1(n1199), .A2(n1049), .A3(n1052), .ZN(n1192) );
NOR2_X1 U871 ( .A1(n1031), .A2(n1064), .ZN(n1052) );
INV_X1 U872 ( .A(n1032), .ZN(n1064) );
NOR3_X1 U873 ( .A1(n1042), .A2(n1167), .A3(n1051), .ZN(n1199) );
INV_X1 U874 ( .A(n1205), .ZN(n1167) );
XOR2_X1 U875 ( .A(G128), .B(n1191), .Z(G30) );
NOR3_X1 U876 ( .A1(n1183), .A2(n1172), .A3(n1197), .ZN(n1191) );
NAND4_X1 U877 ( .A1(n1170), .A2(n1057), .A3(n1205), .A4(n1206), .ZN(n1197) );
XNOR2_X1 U878 ( .A(n1143), .B(n1178), .ZN(G3) );
NOR3_X1 U879 ( .A1(n1051), .A2(n1181), .A3(n1024), .ZN(n1178) );
INV_X1 U880 ( .A(n1195), .ZN(n1024) );
INV_X1 U881 ( .A(G101), .ZN(n1143) );
XOR2_X1 U882 ( .A(G125), .B(n1190), .Z(G27) );
AND2_X1 U883 ( .A1(n1200), .A2(n1028), .ZN(n1190) );
AND4_X1 U884 ( .A1(n1049), .A2(n1205), .A3(n1207), .A4(n1208), .ZN(n1200) );
OR2_X1 U885 ( .A1(n1209), .A2(KEYINPUT35), .ZN(n1208) );
NAND2_X1 U886 ( .A1(KEYINPUT35), .A2(n1210), .ZN(n1207) );
NAND2_X1 U887 ( .A1(n1211), .A2(n1057), .ZN(n1210) );
NAND2_X1 U888 ( .A1(n1021), .A2(n1212), .ZN(n1205) );
NAND4_X1 U889 ( .A1(G953), .A2(G902), .A3(n1213), .A4(n1082), .ZN(n1212) );
INV_X1 U890 ( .A(G900), .ZN(n1082) );
INV_X1 U891 ( .A(n1184), .ZN(n1049) );
XNOR2_X1 U892 ( .A(G122), .B(n1174), .ZN(G24) );
NAND4_X1 U893 ( .A1(n1214), .A2(n1209), .A3(n1058), .A4(n1171), .ZN(n1174) );
INV_X1 U894 ( .A(n1026), .ZN(n1209) );
NAND2_X1 U895 ( .A1(n1215), .A2(n1211), .ZN(n1026) );
XNOR2_X1 U896 ( .A(G119), .B(n1175), .ZN(G21) );
NAND4_X1 U897 ( .A1(n1214), .A2(n1195), .A3(n1057), .A4(n1206), .ZN(n1175) );
INV_X1 U898 ( .A(n1182), .ZN(n1214) );
XNOR2_X1 U899 ( .A(n1216), .B(n1217), .ZN(G18) );
NOR3_X1 U900 ( .A1(n1218), .A2(n1183), .A3(n1182), .ZN(n1217) );
INV_X1 U901 ( .A(n1048), .ZN(n1183) );
NOR2_X1 U902 ( .A1(n1058), .A2(n1219), .ZN(n1048) );
XNOR2_X1 U903 ( .A(KEYINPUT17), .B(n1051), .ZN(n1218) );
XNOR2_X1 U904 ( .A(n1220), .B(n1185), .ZN(G15) );
NOR3_X1 U905 ( .A1(n1051), .A2(n1184), .A3(n1182), .ZN(n1185) );
NAND2_X1 U906 ( .A1(n1028), .A2(n1221), .ZN(n1182) );
NOR2_X1 U907 ( .A1(n1033), .A2(n1172), .ZN(n1028) );
NAND2_X1 U908 ( .A1(n1222), .A2(n1041), .ZN(n1033) );
NAND2_X1 U909 ( .A1(n1219), .A2(n1058), .ZN(n1184) );
NAND2_X1 U910 ( .A1(n1215), .A2(n1206), .ZN(n1051) );
INV_X1 U911 ( .A(n1057), .ZN(n1215) );
XOR2_X1 U912 ( .A(n1223), .B(n1224), .Z(G12) );
NOR3_X1 U913 ( .A1(n1050), .A2(n1225), .A3(n1226), .ZN(n1224) );
NOR2_X1 U914 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
AND3_X1 U915 ( .A1(n1170), .A2(n1221), .A3(n1172), .ZN(n1227) );
AND2_X1 U916 ( .A1(n1228), .A2(n1181), .ZN(n1225) );
NAND3_X1 U917 ( .A1(n1170), .A2(n1221), .A3(n1196), .ZN(n1181) );
INV_X1 U918 ( .A(n1172), .ZN(n1196) );
NAND2_X1 U919 ( .A1(n1031), .A2(n1032), .ZN(n1172) );
NAND2_X1 U920 ( .A1(G214), .A2(n1229), .ZN(n1032) );
XNOR2_X1 U921 ( .A(n1230), .B(n1061), .ZN(n1031) );
NAND2_X1 U922 ( .A1(G210), .A2(n1229), .ZN(n1061) );
NAND2_X1 U923 ( .A1(n1231), .A2(n1232), .ZN(n1229) );
NAND2_X1 U924 ( .A1(n1233), .A2(KEYINPUT29), .ZN(n1230) );
XOR2_X1 U925 ( .A(n1060), .B(KEYINPUT46), .Z(n1233) );
NAND2_X1 U926 ( .A1(n1234), .A2(n1232), .ZN(n1060) );
XOR2_X1 U927 ( .A(n1235), .B(n1236), .Z(n1234) );
XOR2_X1 U928 ( .A(KEYINPUT45), .B(KEYINPUT15), .Z(n1236) );
XNOR2_X1 U929 ( .A(n1159), .B(n1237), .ZN(n1235) );
NOR2_X1 U930 ( .A1(G125), .A2(KEYINPUT41), .ZN(n1237) );
XNOR2_X1 U931 ( .A(n1238), .B(n1239), .ZN(n1159) );
XOR2_X1 U932 ( .A(n1110), .B(n1240), .Z(n1239) );
XOR2_X1 U933 ( .A(n1241), .B(n1242), .Z(n1110) );
XOR2_X1 U934 ( .A(n1243), .B(n1244), .Z(n1242) );
XNOR2_X1 U935 ( .A(KEYINPUT37), .B(n1013), .ZN(n1244) );
NOR2_X1 U936 ( .A1(KEYINPUT7), .A2(n1131), .ZN(n1243) );
INV_X1 U937 ( .A(G104), .ZN(n1131) );
XOR2_X1 U938 ( .A(n1245), .B(n1246), .Z(n1241) );
NAND2_X1 U939 ( .A1(n1247), .A2(n1248), .ZN(n1245) );
NAND2_X1 U940 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
INV_X1 U941 ( .A(KEYINPUT1), .ZN(n1250) );
NAND3_X1 U942 ( .A1(G113), .A2(n1251), .A3(KEYINPUT1), .ZN(n1247) );
XOR2_X1 U943 ( .A(n1252), .B(n1253), .Z(n1238) );
NOR2_X1 U944 ( .A1(G953), .A2(n1106), .ZN(n1253) );
INV_X1 U945 ( .A(G224), .ZN(n1106) );
NAND2_X1 U946 ( .A1(KEYINPUT40), .A2(n1111), .ZN(n1252) );
XNOR2_X1 U947 ( .A(n1254), .B(n1255), .ZN(n1111) );
NOR2_X1 U948 ( .A1(KEYINPUT26), .A2(n1256), .ZN(n1255) );
INV_X1 U949 ( .A(G122), .ZN(n1256) );
NAND2_X1 U950 ( .A1(n1257), .A2(n1021), .ZN(n1221) );
NAND3_X1 U951 ( .A1(n1213), .A2(n1074), .A3(G952), .ZN(n1021) );
NAND4_X1 U952 ( .A1(G953), .A2(G902), .A3(n1213), .A4(n1107), .ZN(n1257) );
INV_X1 U953 ( .A(G898), .ZN(n1107) );
NAND2_X1 U954 ( .A1(G237), .A2(G234), .ZN(n1213) );
INV_X1 U955 ( .A(n1042), .ZN(n1170) );
NAND2_X1 U956 ( .A1(n1040), .A2(n1041), .ZN(n1042) );
NAND2_X1 U957 ( .A1(G221), .A2(n1258), .ZN(n1041) );
INV_X1 U958 ( .A(n1222), .ZN(n1040) );
XOR2_X1 U959 ( .A(n1259), .B(G469), .Z(n1222) );
NAND3_X1 U960 ( .A1(n1260), .A2(n1261), .A3(n1232), .ZN(n1259) );
NAND2_X1 U961 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NAND2_X1 U962 ( .A1(n1152), .A2(n1153), .ZN(n1263) );
NAND2_X1 U963 ( .A1(n1264), .A2(n1145), .ZN(n1153) );
INV_X1 U964 ( .A(n1265), .ZN(n1264) );
NAND2_X1 U965 ( .A1(n1265), .A2(n1266), .ZN(n1152) );
NAND2_X1 U966 ( .A1(n1267), .A2(n1268), .ZN(n1260) );
INV_X1 U967 ( .A(n1262), .ZN(n1268) );
XNOR2_X1 U968 ( .A(n1269), .B(n1270), .ZN(n1262) );
NOR2_X1 U969 ( .A1(KEYINPUT63), .A2(n1150), .ZN(n1270) );
AND2_X1 U970 ( .A1(G227), .A2(n1074), .ZN(n1150) );
XNOR2_X1 U971 ( .A(G110), .B(G140), .ZN(n1269) );
XNOR2_X1 U972 ( .A(n1145), .B(n1265), .ZN(n1267) );
XNOR2_X1 U973 ( .A(n1092), .B(n1271), .ZN(n1265) );
XNOR2_X1 U974 ( .A(n1272), .B(n1246), .ZN(n1271) );
XOR2_X1 U975 ( .A(G101), .B(KEYINPUT27), .Z(n1246) );
NAND3_X1 U976 ( .A1(n1273), .A2(n1274), .A3(KEYINPUT19), .ZN(n1272) );
NAND2_X1 U977 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
INV_X1 U978 ( .A(KEYINPUT8), .ZN(n1276) );
XNOR2_X1 U979 ( .A(G104), .B(G107), .ZN(n1275) );
NAND3_X1 U980 ( .A1(G104), .A2(n1013), .A3(KEYINPUT8), .ZN(n1273) );
INV_X1 U981 ( .A(G107), .ZN(n1013) );
NAND2_X1 U982 ( .A1(n1277), .A2(n1278), .ZN(n1092) );
NAND2_X1 U983 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
INV_X1 U984 ( .A(G146), .ZN(n1280) );
NAND2_X1 U985 ( .A1(n1281), .A2(G146), .ZN(n1277) );
XOR2_X1 U986 ( .A(KEYINPUT9), .B(n1279), .Z(n1281) );
INV_X1 U987 ( .A(KEYINPUT16), .ZN(n1228) );
NAND3_X1 U988 ( .A1(n1211), .A2(n1195), .A3(n1282), .ZN(n1050) );
XNOR2_X1 U989 ( .A(n1057), .B(KEYINPUT35), .ZN(n1282) );
XOR2_X1 U990 ( .A(n1283), .B(n1117), .Z(n1057) );
NAND2_X1 U991 ( .A1(G217), .A2(n1258), .ZN(n1117) );
NAND2_X1 U992 ( .A1(G234), .A2(n1232), .ZN(n1258) );
NAND2_X1 U993 ( .A1(n1115), .A2(n1232), .ZN(n1283) );
XNOR2_X1 U994 ( .A(n1284), .B(n1285), .ZN(n1115) );
XOR2_X1 U995 ( .A(n1286), .B(n1287), .Z(n1285) );
NAND2_X1 U996 ( .A1(G221), .A2(n1288), .ZN(n1287) );
NAND2_X1 U997 ( .A1(KEYINPUT22), .A2(n1289), .ZN(n1286) );
XOR2_X1 U998 ( .A(n1290), .B(n1291), .Z(n1289) );
XNOR2_X1 U999 ( .A(n1292), .B(n1293), .ZN(n1291) );
NAND3_X1 U1000 ( .A1(n1294), .A2(n1295), .A3(n1296), .ZN(n1292) );
OR2_X1 U1001 ( .A1(n1297), .A2(G128), .ZN(n1296) );
NAND2_X1 U1002 ( .A1(n1298), .A2(n1299), .ZN(n1295) );
INV_X1 U1003 ( .A(KEYINPUT12), .ZN(n1299) );
NAND2_X1 U1004 ( .A1(n1300), .A2(n1297), .ZN(n1298) );
XNOR2_X1 U1005 ( .A(KEYINPUT2), .B(G128), .ZN(n1300) );
NAND2_X1 U1006 ( .A1(KEYINPUT12), .A2(n1301), .ZN(n1294) );
NAND2_X1 U1007 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
OR2_X1 U1008 ( .A1(G128), .A2(KEYINPUT2), .ZN(n1303) );
NAND3_X1 U1009 ( .A1(G128), .A2(n1297), .A3(KEYINPUT2), .ZN(n1302) );
INV_X1 U1010 ( .A(G119), .ZN(n1297) );
XNOR2_X1 U1011 ( .A(KEYINPUT53), .B(n1254), .ZN(n1290) );
XNOR2_X1 U1012 ( .A(G137), .B(KEYINPUT0), .ZN(n1284) );
NOR2_X1 U1013 ( .A1(n1171), .A2(n1058), .ZN(n1195) );
XOR2_X1 U1014 ( .A(n1304), .B(n1130), .Z(n1058) );
INV_X1 U1015 ( .A(G475), .ZN(n1130) );
OR2_X1 U1016 ( .A1(n1129), .A2(G902), .ZN(n1304) );
XNOR2_X1 U1017 ( .A(n1305), .B(n1306), .ZN(n1129) );
XOR2_X1 U1018 ( .A(n1293), .B(n1307), .Z(n1306) );
XOR2_X1 U1019 ( .A(n1308), .B(n1309), .Z(n1307) );
NAND2_X1 U1020 ( .A1(KEYINPUT6), .A2(n1220), .ZN(n1309) );
NAND2_X1 U1021 ( .A1(n1310), .A2(n1311), .ZN(n1308) );
NAND2_X1 U1022 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NAND2_X1 U1023 ( .A1(KEYINPUT57), .A2(n1314), .ZN(n1312) );
NAND4_X1 U1024 ( .A1(KEYINPUT60), .A2(G214), .A3(n1231), .A4(n1074), .ZN(n1314) );
NAND2_X1 U1025 ( .A1(n1315), .A2(n1316), .ZN(n1310) );
NAND3_X1 U1026 ( .A1(n1231), .A2(n1074), .A3(G214), .ZN(n1316) );
NAND2_X1 U1027 ( .A1(KEYINPUT60), .A2(n1317), .ZN(n1315) );
NAND2_X1 U1028 ( .A1(KEYINPUT57), .A2(G143), .ZN(n1317) );
XOR2_X1 U1029 ( .A(G146), .B(n1089), .Z(n1293) );
XOR2_X1 U1030 ( .A(G125), .B(G140), .Z(n1089) );
XOR2_X1 U1031 ( .A(n1318), .B(n1319), .Z(n1305) );
XNOR2_X1 U1032 ( .A(KEYINPUT11), .B(n1204), .ZN(n1319) );
XNOR2_X1 U1033 ( .A(G104), .B(G122), .ZN(n1318) );
INV_X1 U1034 ( .A(n1219), .ZN(n1171) );
NOR2_X1 U1035 ( .A1(n1320), .A2(n1069), .ZN(n1219) );
NOR3_X1 U1036 ( .A1(G478), .A2(G902), .A3(n1067), .ZN(n1069) );
AND2_X1 U1037 ( .A1(G478), .A2(n1321), .ZN(n1320) );
NAND2_X1 U1038 ( .A1(n1322), .A2(n1232), .ZN(n1321) );
INV_X1 U1039 ( .A(n1067), .ZN(n1322) );
XNOR2_X1 U1040 ( .A(n1323), .B(n1324), .ZN(n1067) );
XOR2_X1 U1041 ( .A(n1325), .B(n1326), .Z(n1324) );
XNOR2_X1 U1042 ( .A(n1327), .B(n1328), .ZN(n1326) );
NAND2_X1 U1043 ( .A1(KEYINPUT49), .A2(n1203), .ZN(n1328) );
INV_X1 U1044 ( .A(G134), .ZN(n1203) );
NAND2_X1 U1045 ( .A1(KEYINPUT52), .A2(G128), .ZN(n1327) );
NAND2_X1 U1046 ( .A1(G217), .A2(n1288), .ZN(n1325) );
AND2_X1 U1047 ( .A1(G234), .A2(n1074), .ZN(n1288) );
XOR2_X1 U1048 ( .A(n1329), .B(n1330), .Z(n1323) );
NOR2_X1 U1049 ( .A1(KEYINPUT38), .A2(n1331), .ZN(n1330) );
XNOR2_X1 U1050 ( .A(G116), .B(G122), .ZN(n1331) );
XNOR2_X1 U1051 ( .A(G107), .B(G143), .ZN(n1329) );
XOR2_X1 U1052 ( .A(n1206), .B(KEYINPUT43), .Z(n1211) );
NAND3_X1 U1053 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1206) );
INV_X1 U1054 ( .A(n1063), .ZN(n1334) );
NOR2_X1 U1055 ( .A1(n1068), .A2(G472), .ZN(n1063) );
OR2_X1 U1056 ( .A1(G472), .A2(KEYINPUT47), .ZN(n1333) );
NAND3_X1 U1057 ( .A1(G472), .A2(n1068), .A3(KEYINPUT47), .ZN(n1332) );
NAND2_X1 U1058 ( .A1(n1335), .A2(n1232), .ZN(n1068) );
INV_X1 U1059 ( .A(G902), .ZN(n1232) );
XOR2_X1 U1060 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1061 ( .A(KEYINPUT4), .B(n1338), .Z(n1337) );
NOR2_X1 U1062 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
XOR2_X1 U1063 ( .A(n1341), .B(KEYINPUT39), .Z(n1340) );
NAND2_X1 U1064 ( .A1(G101), .A2(n1342), .ZN(n1341) );
NOR2_X1 U1065 ( .A1(G101), .A2(n1342), .ZN(n1339) );
XNOR2_X1 U1066 ( .A(KEYINPUT62), .B(n1142), .ZN(n1342) );
NAND3_X1 U1067 ( .A1(n1231), .A2(n1074), .A3(G210), .ZN(n1142) );
INV_X1 U1068 ( .A(G953), .ZN(n1074) );
INV_X1 U1069 ( .A(G237), .ZN(n1231) );
NAND2_X1 U1070 ( .A1(n1343), .A2(n1344), .ZN(n1336) );
NAND2_X1 U1071 ( .A1(n1345), .A2(n1266), .ZN(n1344) );
INV_X1 U1072 ( .A(n1145), .ZN(n1266) );
NAND2_X1 U1073 ( .A1(n1346), .A2(n1145), .ZN(n1343) );
XOR2_X1 U1074 ( .A(n1347), .B(n1204), .Z(n1145) );
INV_X1 U1075 ( .A(G131), .ZN(n1204) );
NAND2_X1 U1076 ( .A1(KEYINPUT3), .A2(n1098), .ZN(n1347) );
XOR2_X1 U1077 ( .A(G134), .B(G137), .Z(n1098) );
XNOR2_X1 U1078 ( .A(KEYINPUT33), .B(n1345), .ZN(n1346) );
INV_X1 U1079 ( .A(n1144), .ZN(n1345) );
XNOR2_X1 U1080 ( .A(n1240), .B(n1249), .ZN(n1144) );
XNOR2_X1 U1081 ( .A(n1220), .B(n1251), .ZN(n1249) );
XNOR2_X1 U1082 ( .A(n1216), .B(G119), .ZN(n1251) );
INV_X1 U1083 ( .A(G116), .ZN(n1216) );
INV_X1 U1084 ( .A(G113), .ZN(n1220) );
XNOR2_X1 U1085 ( .A(G146), .B(n1279), .ZN(n1240) );
XNOR2_X1 U1086 ( .A(n1313), .B(G128), .ZN(n1279) );
INV_X1 U1087 ( .A(G143), .ZN(n1313) );
NAND2_X1 U1088 ( .A1(KEYINPUT31), .A2(n1254), .ZN(n1223) );
INV_X1 U1089 ( .A(G110), .ZN(n1254) );
endmodule


