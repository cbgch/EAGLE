//Key = 0110101100010001000111101101111001001100011001101100011011010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367;

XOR2_X1 U742 ( .A(n1028), .B(n1029), .Z(G9) );
NOR2_X1 U743 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U744 ( .A1(n1032), .A2(n1033), .A3(G953), .A4(n1034), .ZN(n1031) );
NOR2_X1 U745 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U746 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR3_X1 U747 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NOR2_X1 U748 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U749 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U750 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U751 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U752 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR2_X1 U753 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR3_X1 U754 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1046) );
NOR2_X1 U755 ( .A1(n1057), .A2(n1055), .ZN(n1042) );
NOR2_X1 U756 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
AND2_X1 U757 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR4_X1 U758 ( .A1(n1062), .A2(n1055), .A3(n1045), .A4(n1049), .ZN(n1037) );
NOR2_X1 U759 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U760 ( .A1(n1065), .A2(n1041), .ZN(n1063) );
NAND3_X1 U761 ( .A1(n1066), .A2(G952), .A3(n1067), .ZN(n1032) );
NOR3_X1 U762 ( .A1(n1034), .A2(n1068), .A3(n1069), .ZN(n1030) );
NOR2_X1 U763 ( .A1(KEYINPUT38), .A2(n1070), .ZN(n1069) );
NOR2_X1 U764 ( .A1(G953), .A2(G952), .ZN(n1070) );
NOR2_X1 U765 ( .A1(n1071), .A2(n1072), .ZN(n1068) );
INV_X1 U766 ( .A(KEYINPUT38), .ZN(n1072) );
AND4_X1 U767 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1034) );
NOR3_X1 U768 ( .A1(n1077), .A2(n1039), .A3(n1078), .ZN(n1076) );
NAND3_X1 U769 ( .A1(n1053), .A2(n1079), .A3(n1054), .ZN(n1077) );
NOR3_X1 U770 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1075) );
NOR3_X1 U771 ( .A1(n1083), .A2(KEYINPUT3), .A3(n1084), .ZN(n1082) );
NOR2_X1 U772 ( .A1(G902), .A2(n1085), .ZN(n1084) );
AND2_X1 U773 ( .A1(n1083), .A2(KEYINPUT3), .ZN(n1081) );
XOR2_X1 U774 ( .A(G472), .B(n1086), .Z(n1080) );
NOR2_X1 U775 ( .A1(KEYINPUT5), .A2(n1087), .ZN(n1086) );
XNOR2_X1 U776 ( .A(n1088), .B(n1089), .ZN(n1074) );
XOR2_X1 U777 ( .A(n1090), .B(G469), .Z(n1073) );
XOR2_X1 U778 ( .A(n1091), .B(n1092), .Z(G72) );
NOR2_X1 U779 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR2_X1 U780 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NAND2_X1 U781 ( .A1(n1097), .A2(n1098), .ZN(n1091) );
NAND2_X1 U782 ( .A1(n1099), .A2(n1094), .ZN(n1098) );
XOR2_X1 U783 ( .A(n1100), .B(n1067), .Z(n1099) );
OR3_X1 U784 ( .A1(n1100), .A2(n1096), .A3(n1094), .ZN(n1097) );
NAND2_X1 U785 ( .A1(KEYINPUT2), .A2(n1101), .ZN(n1100) );
XOR2_X1 U786 ( .A(KEYINPUT60), .B(n1102), .Z(n1101) );
NOR2_X1 U787 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XOR2_X1 U788 ( .A(n1105), .B(KEYINPUT19), .Z(n1104) );
NAND2_X1 U789 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1103) );
XNOR2_X1 U791 ( .A(n1108), .B(n1109), .ZN(n1107) );
XOR2_X1 U792 ( .A(G131), .B(n1110), .Z(n1109) );
XNOR2_X1 U793 ( .A(KEYINPUT1), .B(n1111), .ZN(n1106) );
NAND2_X1 U794 ( .A1(n1112), .A2(n1113), .ZN(G69) );
NAND3_X1 U795 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1113) );
XOR2_X1 U796 ( .A(KEYINPUT33), .B(n1117), .Z(n1112) );
NOR2_X1 U797 ( .A1(n1118), .A2(n1116), .ZN(n1117) );
AND2_X1 U798 ( .A1(n1119), .A2(n1120), .ZN(n1116) );
NAND2_X1 U799 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U800 ( .A1(n1123), .A2(n1094), .ZN(n1122) );
INV_X1 U801 ( .A(n1124), .ZN(n1121) );
NAND3_X1 U802 ( .A1(n1123), .A2(n1094), .A3(n1124), .ZN(n1119) );
NAND2_X1 U803 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U804 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U805 ( .A(KEYINPUT0), .B(G953), .Z(n1127) );
XNOR2_X1 U806 ( .A(n1129), .B(n1130), .ZN(n1125) );
XOR2_X1 U807 ( .A(G122), .B(n1131), .Z(n1130) );
NOR2_X1 U808 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XOR2_X1 U809 ( .A(KEYINPUT34), .B(n1134), .Z(n1133) );
NOR2_X1 U810 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NOR2_X1 U811 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
INV_X1 U812 ( .A(n1135), .ZN(n1138) );
XNOR2_X1 U813 ( .A(n1136), .B(KEYINPUT32), .ZN(n1137) );
XOR2_X1 U814 ( .A(G113), .B(n1139), .Z(n1136) );
AND2_X1 U815 ( .A1(n1115), .A2(n1114), .ZN(n1118) );
XNOR2_X1 U816 ( .A(G953), .B(KEYINPUT49), .ZN(n1114) );
NAND2_X1 U817 ( .A1(G898), .A2(G224), .ZN(n1115) );
NOR2_X1 U818 ( .A1(n1071), .A2(n1140), .ZN(G66) );
XOR2_X1 U819 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U820 ( .A(KEYINPUT20), .B(n1143), .Z(n1142) );
NOR2_X1 U821 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NOR2_X1 U822 ( .A1(n1071), .A2(n1146), .ZN(G63) );
XNOR2_X1 U823 ( .A(n1147), .B(n1148), .ZN(n1146) );
NOR2_X1 U824 ( .A1(n1149), .A2(n1145), .ZN(n1148) );
INV_X1 U825 ( .A(G478), .ZN(n1149) );
NOR2_X1 U826 ( .A1(n1071), .A2(n1150), .ZN(G60) );
XOR2_X1 U827 ( .A(n1085), .B(n1151), .Z(n1150) );
NOR2_X1 U828 ( .A1(n1083), .A2(n1145), .ZN(n1151) );
XNOR2_X1 U829 ( .A(G104), .B(n1152), .ZN(G6) );
NOR2_X1 U830 ( .A1(n1071), .A2(n1153), .ZN(G57) );
XOR2_X1 U831 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U832 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U833 ( .A(n1158), .B(n1159), .Z(n1154) );
NOR2_X1 U834 ( .A1(n1160), .A2(n1145), .ZN(n1159) );
INV_X1 U835 ( .A(G472), .ZN(n1160) );
XNOR2_X1 U836 ( .A(n1161), .B(n1162), .ZN(n1158) );
NOR2_X1 U837 ( .A1(KEYINPUT9), .A2(n1163), .ZN(n1162) );
XOR2_X1 U838 ( .A(n1164), .B(KEYINPUT39), .Z(n1163) );
NOR2_X1 U839 ( .A1(KEYINPUT12), .A2(n1165), .ZN(n1161) );
XOR2_X1 U840 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U841 ( .A1(n1071), .A2(n1168), .ZN(G54) );
XOR2_X1 U842 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U843 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U844 ( .A1(KEYINPUT35), .A2(n1173), .ZN(n1172) );
XOR2_X1 U845 ( .A(G140), .B(G110), .Z(n1173) );
NOR2_X1 U846 ( .A1(n1174), .A2(n1175), .ZN(n1171) );
INV_X1 U847 ( .A(KEYINPUT35), .ZN(n1175) );
NOR2_X1 U848 ( .A1(n1176), .A2(n1177), .ZN(n1174) );
XOR2_X1 U849 ( .A(n1178), .B(n1179), .Z(n1169) );
NOR2_X1 U850 ( .A1(n1180), .A2(n1145), .ZN(n1179) );
INV_X1 U851 ( .A(G469), .ZN(n1180) );
NOR2_X1 U852 ( .A1(n1071), .A2(n1181), .ZN(G51) );
XOR2_X1 U853 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U854 ( .A(KEYINPUT29), .B(n1184), .Z(n1183) );
NOR2_X1 U855 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U856 ( .A(n1187), .B(KEYINPUT46), .Z(n1186) );
NAND2_X1 U857 ( .A1(n1188), .A2(G125), .ZN(n1187) );
NOR2_X1 U858 ( .A1(G125), .A2(n1188), .ZN(n1185) );
XOR2_X1 U859 ( .A(n1189), .B(n1190), .Z(n1182) );
NOR2_X1 U860 ( .A1(n1089), .A2(n1145), .ZN(n1190) );
NAND2_X1 U861 ( .A1(G902), .A2(n1191), .ZN(n1145) );
NAND2_X1 U862 ( .A1(n1067), .A2(n1066), .ZN(n1191) );
INV_X1 U863 ( .A(n1123), .ZN(n1066) );
NAND4_X1 U864 ( .A1(n1192), .A2(n1029), .A3(n1193), .A4(n1194), .ZN(n1123) );
AND3_X1 U865 ( .A1(n1195), .A2(n1196), .A3(n1152), .ZN(n1194) );
NAND3_X1 U866 ( .A1(n1065), .A2(n1197), .A3(n1198), .ZN(n1152) );
OR2_X1 U867 ( .A1(n1199), .A2(n1200), .ZN(n1195) );
NOR2_X1 U868 ( .A1(n1201), .A2(n1202), .ZN(n1199) );
INV_X1 U869 ( .A(n1203), .ZN(n1202) );
AND2_X1 U870 ( .A1(n1059), .A2(n1064), .ZN(n1201) );
NAND2_X1 U871 ( .A1(n1204), .A2(n1205), .ZN(n1059) );
NAND2_X1 U872 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U873 ( .A1(n1198), .A2(n1061), .ZN(n1204) );
NAND3_X1 U874 ( .A1(n1065), .A2(n1197), .A3(n1060), .ZN(n1029) );
AND4_X1 U875 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1067) );
NOR4_X1 U876 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1211) );
INV_X1 U877 ( .A(n1216), .ZN(n1213) );
NOR3_X1 U878 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1210) );
NOR3_X1 U879 ( .A1(n1220), .A2(n1221), .A3(n1055), .ZN(n1219) );
INV_X1 U880 ( .A(n1222), .ZN(n1055) );
INV_X1 U881 ( .A(KEYINPUT23), .ZN(n1220) );
NOR2_X1 U882 ( .A1(KEYINPUT23), .A2(n1223), .ZN(n1218) );
NOR2_X1 U883 ( .A1(n1094), .A2(G952), .ZN(n1071) );
XOR2_X1 U884 ( .A(G146), .B(n1217), .Z(G48) );
AND3_X1 U885 ( .A1(n1224), .A2(n1051), .A3(n1198), .ZN(n1217) );
XNOR2_X1 U886 ( .A(G143), .B(n1208), .ZN(G45) );
NAND4_X1 U887 ( .A1(n1064), .A2(n1225), .A3(n1226), .A4(n1051), .ZN(n1208) );
NOR2_X1 U888 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NAND2_X1 U889 ( .A1(n1229), .A2(n1230), .ZN(G42) );
OR2_X1 U890 ( .A1(G140), .A2(KEYINPUT63), .ZN(n1230) );
XNOR2_X1 U891 ( .A(n1231), .B(n1223), .ZN(n1229) );
NAND2_X1 U892 ( .A1(n1221), .A2(n1222), .ZN(n1223) );
AND4_X1 U893 ( .A1(n1198), .A2(n1225), .A3(n1232), .A4(n1039), .ZN(n1221) );
NAND2_X1 U894 ( .A1(KEYINPUT63), .A2(G140), .ZN(n1231) );
XOR2_X1 U895 ( .A(n1233), .B(n1212), .Z(G39) );
AND3_X1 U896 ( .A1(n1224), .A2(n1222), .A3(n1206), .ZN(n1212) );
NAND2_X1 U897 ( .A1(KEYINPUT30), .A2(n1234), .ZN(n1233) );
INV_X1 U898 ( .A(G137), .ZN(n1234) );
XNOR2_X1 U899 ( .A(G134), .B(n1209), .ZN(G36) );
NAND2_X1 U900 ( .A1(n1235), .A2(n1060), .ZN(n1209) );
XOR2_X1 U901 ( .A(n1236), .B(n1215), .Z(G33) );
AND2_X1 U902 ( .A1(n1235), .A2(n1198), .ZN(n1215) );
AND3_X1 U903 ( .A1(n1222), .A2(n1225), .A3(n1064), .ZN(n1235) );
NOR2_X1 U904 ( .A1(n1052), .A2(n1237), .ZN(n1222) );
XNOR2_X1 U905 ( .A(n1238), .B(KEYINPUT47), .ZN(n1052) );
XNOR2_X1 U906 ( .A(G131), .B(KEYINPUT27), .ZN(n1236) );
XOR2_X1 U907 ( .A(G128), .B(n1214), .Z(G30) );
AND3_X1 U908 ( .A1(n1060), .A2(n1051), .A3(n1224), .ZN(n1214) );
AND3_X1 U909 ( .A1(n1239), .A2(n1240), .A3(n1225), .ZN(n1224) );
AND2_X1 U910 ( .A1(n1207), .A2(n1241), .ZN(n1225) );
INV_X1 U911 ( .A(n1242), .ZN(n1207) );
OR2_X1 U912 ( .A1(n1243), .A2(n1064), .ZN(n1240) );
NAND2_X1 U913 ( .A1(n1244), .A2(n1243), .ZN(n1239) );
NAND2_X1 U914 ( .A1(n1041), .A2(n1039), .ZN(n1244) );
XOR2_X1 U915 ( .A(n1245), .B(n1246), .Z(G3) );
NOR2_X1 U916 ( .A1(KEYINPUT50), .A2(n1166), .ZN(n1246) );
NOR3_X1 U917 ( .A1(n1247), .A2(n1242), .A3(n1045), .ZN(n1245) );
NAND3_X1 U918 ( .A1(n1248), .A2(n1249), .A3(n1064), .ZN(n1247) );
OR2_X1 U919 ( .A1(n1250), .A2(KEYINPUT52), .ZN(n1249) );
NAND2_X1 U920 ( .A1(KEYINPUT52), .A2(n1251), .ZN(n1248) );
NAND2_X1 U921 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
XOR2_X1 U922 ( .A(n1254), .B(n1216), .Z(G27) );
NAND4_X1 U923 ( .A1(n1039), .A2(n1241), .A3(n1051), .A4(n1255), .ZN(n1216) );
AND3_X1 U924 ( .A1(n1198), .A2(n1061), .A3(n1232), .ZN(n1255) );
NAND2_X1 U925 ( .A1(n1256), .A2(n1257), .ZN(n1241) );
NAND4_X1 U926 ( .A1(G953), .A2(G902), .A3(n1258), .A4(n1096), .ZN(n1257) );
INV_X1 U927 ( .A(G900), .ZN(n1096) );
XNOR2_X1 U928 ( .A(KEYINPUT28), .B(n1036), .ZN(n1256) );
XOR2_X1 U929 ( .A(n1259), .B(n1260), .Z(G24) );
NOR4_X1 U930 ( .A1(n1261), .A2(n1262), .A3(KEYINPUT40), .A4(n1203), .ZN(n1260) );
NAND3_X1 U931 ( .A1(n1065), .A2(n1061), .A3(n1263), .ZN(n1203) );
NOR3_X1 U932 ( .A1(n1041), .A2(n1227), .A3(n1228), .ZN(n1263) );
NOR2_X1 U933 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
INV_X1 U934 ( .A(KEYINPUT26), .ZN(n1265) );
NOR2_X1 U935 ( .A1(n1253), .A2(n1252), .ZN(n1264) );
NOR2_X1 U936 ( .A1(KEYINPUT26), .A2(n1250), .ZN(n1261) );
XNOR2_X1 U937 ( .A(G122), .B(KEYINPUT4), .ZN(n1259) );
XNOR2_X1 U938 ( .A(G119), .B(n1196), .ZN(G21) );
NAND4_X1 U939 ( .A1(n1061), .A2(n1206), .A3(n1266), .A4(n1250), .ZN(n1196) );
NOR2_X1 U940 ( .A1(n1232), .A2(n1267), .ZN(n1266) );
XOR2_X1 U941 ( .A(n1243), .B(n1039), .Z(n1267) );
INV_X1 U942 ( .A(KEYINPUT31), .ZN(n1243) );
XNOR2_X1 U943 ( .A(G116), .B(n1193), .ZN(G18) );
NAND4_X1 U944 ( .A1(n1064), .A2(n1061), .A3(n1060), .A4(n1250), .ZN(n1193) );
INV_X1 U945 ( .A(n1200), .ZN(n1250) );
NOR2_X1 U946 ( .A1(n1268), .A2(n1228), .ZN(n1060) );
XOR2_X1 U947 ( .A(n1269), .B(n1270), .Z(G15) );
XOR2_X1 U948 ( .A(KEYINPUT56), .B(G113), .Z(n1270) );
NAND3_X1 U949 ( .A1(n1271), .A2(n1064), .A3(n1272), .ZN(n1269) );
AND3_X1 U950 ( .A1(n1198), .A2(n1252), .A3(n1061), .ZN(n1272) );
INV_X1 U951 ( .A(n1049), .ZN(n1061) );
NAND2_X1 U952 ( .A1(n1273), .A2(n1054), .ZN(n1049) );
NOR2_X1 U953 ( .A1(n1078), .A2(n1227), .ZN(n1198) );
INV_X1 U954 ( .A(n1228), .ZN(n1078) );
NOR2_X1 U955 ( .A1(n1039), .A2(n1232), .ZN(n1064) );
XOR2_X1 U956 ( .A(n1253), .B(KEYINPUT48), .Z(n1271) );
INV_X1 U957 ( .A(n1051), .ZN(n1253) );
XOR2_X1 U958 ( .A(n1274), .B(n1192), .Z(G12) );
NAND3_X1 U959 ( .A1(n1197), .A2(n1039), .A3(n1206), .ZN(n1192) );
INV_X1 U960 ( .A(n1045), .ZN(n1206) );
NAND2_X1 U961 ( .A1(n1228), .A2(n1227), .ZN(n1045) );
INV_X1 U962 ( .A(n1268), .ZN(n1227) );
NAND2_X1 U963 ( .A1(n1079), .A2(n1275), .ZN(n1268) );
NAND2_X1 U964 ( .A1(G475), .A2(n1276), .ZN(n1275) );
NAND2_X1 U965 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND3_X1 U966 ( .A1(n1083), .A2(n1278), .A3(n1277), .ZN(n1079) );
INV_X1 U967 ( .A(n1085), .ZN(n1277) );
XOR2_X1 U968 ( .A(n1279), .B(n1280), .Z(n1085) );
XOR2_X1 U969 ( .A(n1281), .B(n1282), .Z(n1280) );
XOR2_X1 U970 ( .A(G104), .B(n1283), .Z(n1282) );
NOR2_X1 U971 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U972 ( .A(n1286), .B(KEYINPUT54), .Z(n1285) );
NAND4_X1 U973 ( .A1(G143), .A2(G214), .A3(n1287), .A4(n1094), .ZN(n1286) );
NOR2_X1 U974 ( .A1(n1288), .A2(n1289), .ZN(n1284) );
XOR2_X1 U975 ( .A(KEYINPUT61), .B(G143), .Z(n1289) );
AND3_X1 U976 ( .A1(G214), .A2(n1094), .A3(n1287), .ZN(n1288) );
XOR2_X1 U977 ( .A(KEYINPUT57), .B(G131), .Z(n1281) );
XNOR2_X1 U978 ( .A(n1290), .B(n1291), .ZN(n1279) );
XOR2_X1 U979 ( .A(n1292), .B(n1111), .Z(n1291) );
NOR2_X1 U980 ( .A1(G146), .A2(KEYINPUT44), .ZN(n1292) );
INV_X1 U981 ( .A(G475), .ZN(n1083) );
XOR2_X1 U982 ( .A(n1293), .B(G478), .Z(n1228) );
NAND2_X1 U983 ( .A1(n1147), .A2(n1278), .ZN(n1293) );
XNOR2_X1 U984 ( .A(n1294), .B(n1295), .ZN(n1147) );
XOR2_X1 U985 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U986 ( .A(G122), .B(G116), .Z(n1297) );
XOR2_X1 U987 ( .A(G143), .B(G134), .Z(n1296) );
XNOR2_X1 U988 ( .A(n1298), .B(n1299), .ZN(n1294) );
XOR2_X1 U989 ( .A(n1300), .B(G107), .Z(n1298) );
NAND2_X1 U990 ( .A1(G217), .A2(n1301), .ZN(n1300) );
INV_X1 U991 ( .A(n1065), .ZN(n1039) );
XNOR2_X1 U992 ( .A(n1302), .B(n1144), .ZN(n1065) );
NAND2_X1 U993 ( .A1(G217), .A2(n1303), .ZN(n1144) );
NAND2_X1 U994 ( .A1(n1304), .A2(n1278), .ZN(n1302) );
XOR2_X1 U995 ( .A(KEYINPUT8), .B(n1141), .Z(n1304) );
XNOR2_X1 U996 ( .A(n1305), .B(n1306), .ZN(n1141) );
XOR2_X1 U997 ( .A(n1307), .B(n1308), .Z(n1306) );
XOR2_X1 U998 ( .A(G119), .B(G110), .Z(n1308) );
XOR2_X1 U999 ( .A(KEYINPUT36), .B(G146), .Z(n1307) );
XOR2_X1 U1000 ( .A(n1309), .B(n1310), .Z(n1305) );
XNOR2_X1 U1001 ( .A(n1299), .B(n1111), .ZN(n1310) );
XOR2_X1 U1002 ( .A(G125), .B(G140), .Z(n1111) );
XOR2_X1 U1003 ( .A(n1311), .B(n1312), .Z(n1309) );
NOR2_X1 U1004 ( .A1(G137), .A2(KEYINPUT55), .ZN(n1312) );
NAND2_X1 U1005 ( .A1(n1313), .A2(n1301), .ZN(n1311) );
AND2_X1 U1006 ( .A1(G234), .A2(n1094), .ZN(n1301) );
XNOR2_X1 U1007 ( .A(G221), .B(KEYINPUT41), .ZN(n1313) );
NOR3_X1 U1008 ( .A1(n1041), .A2(n1242), .A3(n1200), .ZN(n1197) );
NAND2_X1 U1009 ( .A1(n1051), .A2(n1252), .ZN(n1200) );
NAND2_X1 U1010 ( .A1(n1036), .A2(n1314), .ZN(n1252) );
NAND4_X1 U1011 ( .A1(G953), .A2(G902), .A3(n1258), .A4(n1128), .ZN(n1314) );
INV_X1 U1012 ( .A(G898), .ZN(n1128) );
NAND3_X1 U1013 ( .A1(n1258), .A2(n1094), .A3(G952), .ZN(n1036) );
NAND2_X1 U1014 ( .A1(G237), .A2(G234), .ZN(n1258) );
NOR2_X1 U1015 ( .A1(n1238), .A2(n1237), .ZN(n1051) );
XOR2_X1 U1016 ( .A(n1053), .B(KEYINPUT6), .Z(n1237) );
NAND2_X1 U1017 ( .A1(G214), .A2(n1315), .ZN(n1053) );
XNOR2_X1 U1018 ( .A(n1088), .B(n1316), .ZN(n1238) );
NOR2_X1 U1019 ( .A1(KEYINPUT58), .A2(n1317), .ZN(n1316) );
XOR2_X1 U1020 ( .A(n1089), .B(KEYINPUT24), .Z(n1317) );
NAND2_X1 U1021 ( .A1(G210), .A2(n1315), .ZN(n1089) );
NAND2_X1 U1022 ( .A1(n1287), .A2(n1278), .ZN(n1315) );
NAND2_X1 U1023 ( .A1(n1318), .A2(n1278), .ZN(n1088) );
XOR2_X1 U1024 ( .A(n1319), .B(n1320), .Z(n1318) );
INV_X1 U1025 ( .A(n1189), .ZN(n1320) );
XOR2_X1 U1026 ( .A(n1321), .B(n1322), .Z(n1189) );
XOR2_X1 U1027 ( .A(n1139), .B(n1323), .Z(n1322) );
XOR2_X1 U1028 ( .A(n1129), .B(n1324), .Z(n1323) );
NAND2_X1 U1029 ( .A1(G224), .A2(n1094), .ZN(n1324) );
NAND2_X1 U1030 ( .A1(n1325), .A2(KEYINPUT53), .ZN(n1129) );
XOR2_X1 U1031 ( .A(n1274), .B(KEYINPUT18), .Z(n1325) );
XOR2_X1 U1032 ( .A(n1135), .B(n1290), .Z(n1321) );
XOR2_X1 U1033 ( .A(G113), .B(G122), .Z(n1290) );
XOR2_X1 U1034 ( .A(n1326), .B(KEYINPUT14), .Z(n1135) );
NAND3_X1 U1035 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1326) );
NAND2_X1 U1036 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
INV_X1 U1037 ( .A(KEYINPUT25), .ZN(n1331) );
NAND3_X1 U1038 ( .A1(KEYINPUT25), .A2(n1332), .A3(n1166), .ZN(n1328) );
OR2_X1 U1039 ( .A1(n1166), .A2(n1332), .ZN(n1327) );
NOR2_X1 U1040 ( .A1(n1333), .A2(n1330), .ZN(n1332) );
XNOR2_X1 U1041 ( .A(n1334), .B(G104), .ZN(n1330) );
NAND2_X1 U1042 ( .A1(KEYINPUT11), .A2(n1028), .ZN(n1334) );
INV_X1 U1043 ( .A(G107), .ZN(n1028) );
INV_X1 U1044 ( .A(KEYINPUT7), .ZN(n1333) );
NOR2_X1 U1045 ( .A1(KEYINPUT10), .A2(n1335), .ZN(n1319) );
NOR2_X1 U1046 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XOR2_X1 U1047 ( .A(n1338), .B(KEYINPUT37), .Z(n1337) );
NAND2_X1 U1048 ( .A1(n1157), .A2(n1254), .ZN(n1338) );
NOR2_X1 U1049 ( .A1(n1254), .A2(n1157), .ZN(n1336) );
INV_X1 U1050 ( .A(G125), .ZN(n1254) );
NAND2_X1 U1051 ( .A1(n1056), .A2(n1054), .ZN(n1242) );
NAND2_X1 U1052 ( .A1(G221), .A2(n1303), .ZN(n1054) );
NAND2_X1 U1053 ( .A1(G234), .A2(n1278), .ZN(n1303) );
INV_X1 U1054 ( .A(n1273), .ZN(n1056) );
XNOR2_X1 U1055 ( .A(n1339), .B(n1090), .ZN(n1273) );
NAND2_X1 U1056 ( .A1(n1340), .A2(n1278), .ZN(n1090) );
XOR2_X1 U1057 ( .A(n1178), .B(n1341), .Z(n1340) );
NOR2_X1 U1058 ( .A1(n1177), .A2(n1342), .ZN(n1341) );
XOR2_X1 U1059 ( .A(KEYINPUT13), .B(n1176), .Z(n1342) );
NOR2_X1 U1060 ( .A1(G140), .A2(n1274), .ZN(n1176) );
AND2_X1 U1061 ( .A1(G140), .A2(n1274), .ZN(n1177) );
XOR2_X1 U1062 ( .A(n1343), .B(n1344), .Z(n1178) );
XOR2_X1 U1063 ( .A(G101), .B(n1345), .Z(n1344) );
XOR2_X1 U1064 ( .A(G107), .B(G104), .Z(n1345) );
XOR2_X1 U1065 ( .A(n1108), .B(n1346), .Z(n1343) );
XOR2_X1 U1066 ( .A(n1347), .B(n1348), .Z(n1346) );
INV_X1 U1067 ( .A(n1156), .ZN(n1348) );
NOR2_X1 U1068 ( .A1(G953), .A2(n1095), .ZN(n1347) );
INV_X1 U1069 ( .A(G227), .ZN(n1095) );
XOR2_X1 U1070 ( .A(n1349), .B(n1350), .Z(n1108) );
NAND2_X1 U1071 ( .A1(KEYINPUT15), .A2(n1351), .ZN(n1349) );
NAND2_X1 U1072 ( .A1(KEYINPUT59), .A2(G469), .ZN(n1339) );
INV_X1 U1073 ( .A(n1232), .ZN(n1041) );
XOR2_X1 U1074 ( .A(n1087), .B(G472), .Z(n1232) );
NAND2_X1 U1075 ( .A1(n1352), .A2(n1278), .ZN(n1087) );
INV_X1 U1076 ( .A(G902), .ZN(n1278) );
XOR2_X1 U1077 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1078 ( .A(n1355), .B(n1356), .Z(n1354) );
NOR2_X1 U1079 ( .A1(KEYINPUT62), .A2(n1156), .ZN(n1356) );
XNOR2_X1 U1080 ( .A(n1110), .B(n1357), .ZN(n1156) );
NOR2_X1 U1081 ( .A1(G131), .A2(KEYINPUT16), .ZN(n1357) );
XOR2_X1 U1082 ( .A(G134), .B(G137), .Z(n1110) );
NOR3_X1 U1083 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1355) );
NOR3_X1 U1084 ( .A1(n1361), .A2(n1362), .A3(n1167), .ZN(n1360) );
AND2_X1 U1085 ( .A1(n1361), .A2(n1167), .ZN(n1359) );
INV_X1 U1086 ( .A(KEYINPUT42), .ZN(n1361) );
NOR2_X1 U1087 ( .A1(n1363), .A2(n1166), .ZN(n1358) );
INV_X1 U1088 ( .A(G101), .ZN(n1166) );
NOR2_X1 U1089 ( .A1(n1364), .A2(n1167), .ZN(n1363) );
NAND3_X1 U1090 ( .A1(n1287), .A2(n1094), .A3(G210), .ZN(n1167) );
INV_X1 U1091 ( .A(G953), .ZN(n1094) );
INV_X1 U1092 ( .A(G237), .ZN(n1287) );
INV_X1 U1093 ( .A(n1362), .ZN(n1364) );
XOR2_X1 U1094 ( .A(n1365), .B(G101), .Z(n1362) );
XNOR2_X1 U1095 ( .A(KEYINPUT43), .B(KEYINPUT21), .ZN(n1365) );
XOR2_X1 U1096 ( .A(n1164), .B(n1157), .Z(n1353) );
INV_X1 U1097 ( .A(n1188), .ZN(n1157) );
XOR2_X1 U1098 ( .A(n1366), .B(n1350), .Z(n1188) );
XNOR2_X1 U1099 ( .A(n1299), .B(KEYINPUT22), .ZN(n1350) );
XNOR2_X1 U1100 ( .A(G128), .B(KEYINPUT51), .ZN(n1299) );
XNOR2_X1 U1101 ( .A(n1351), .B(KEYINPUT45), .ZN(n1366) );
XOR2_X1 U1102 ( .A(G143), .B(G146), .Z(n1351) );
XNOR2_X1 U1103 ( .A(G113), .B(n1367), .ZN(n1164) );
NOR2_X1 U1104 ( .A1(KEYINPUT17), .A2(n1139), .ZN(n1367) );
XOR2_X1 U1105 ( .A(G116), .B(G119), .Z(n1139) );
INV_X1 U1106 ( .A(G110), .ZN(n1274) );
endmodule


