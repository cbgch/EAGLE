//Key = 0010100011001000010011000000100001100111100000110110000000010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330;

XNOR2_X1 U729 ( .A(G107), .B(n1014), .ZN(G9) );
NAND2_X1 U730 ( .A1(n1015), .A2(n1016), .ZN(G75) );
NAND2_X1 U731 ( .A1(G952), .A2(n1017), .ZN(n1016) );
NAND4_X1 U732 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
AND3_X1 U733 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1021) );
NAND3_X1 U734 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1019) );
NAND2_X1 U735 ( .A1(n1028), .A2(n1029), .ZN(n1025) );
NAND3_X1 U736 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NAND2_X1 U737 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NAND2_X1 U738 ( .A1(KEYINPUT29), .A2(n1035), .ZN(n1033) );
NAND4_X1 U739 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1030) );
NAND2_X1 U740 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NAND2_X1 U741 ( .A1(n1042), .A2(n1043), .ZN(n1037) );
OR2_X1 U742 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U743 ( .A1(n1035), .A2(n1046), .ZN(n1036) );
INV_X1 U744 ( .A(KEYINPUT29), .ZN(n1046) );
NAND2_X1 U745 ( .A1(n1047), .A2(n1048), .ZN(n1028) );
NAND2_X1 U746 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U747 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
INV_X1 U748 ( .A(n1053), .ZN(n1049) );
NAND3_X1 U749 ( .A1(n1032), .A2(n1054), .A3(n1047), .ZN(n1018) );
AND3_X1 U750 ( .A1(n1041), .A2(n1042), .A3(n1039), .ZN(n1047) );
INV_X1 U751 ( .A(n1034), .ZN(n1039) );
NAND2_X1 U752 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U753 ( .A1(n1057), .A2(n1027), .ZN(n1056) );
INV_X1 U754 ( .A(n1058), .ZN(n1055) );
NAND2_X1 U755 ( .A1(n1059), .A2(n1060), .ZN(n1015) );
INV_X1 U756 ( .A(G952), .ZN(n1060) );
NAND2_X1 U757 ( .A1(n1061), .A2(n1023), .ZN(n1059) );
NAND4_X1 U758 ( .A1(n1062), .A2(n1051), .A3(n1063), .A4(n1064), .ZN(n1023) );
NOR4_X1 U759 ( .A1(n1052), .A2(n1057), .A3(n1065), .A4(n1066), .ZN(n1064) );
XNOR2_X1 U760 ( .A(n1067), .B(n1068), .ZN(n1066) );
NAND2_X1 U761 ( .A1(KEYINPUT47), .A2(n1069), .ZN(n1067) );
XOR2_X1 U762 ( .A(n1070), .B(n1071), .Z(n1065) );
NOR2_X1 U763 ( .A1(G469), .A2(KEYINPUT58), .ZN(n1071) );
NOR2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(n1063) );
XNOR2_X1 U765 ( .A(n1074), .B(n1075), .ZN(n1072) );
XNOR2_X1 U766 ( .A(n1076), .B(KEYINPUT59), .ZN(n1074) );
XOR2_X1 U767 ( .A(n1024), .B(KEYINPUT35), .Z(n1061) );
XOR2_X1 U768 ( .A(n1077), .B(n1078), .Z(G72) );
NOR2_X1 U769 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U770 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NAND2_X1 U771 ( .A1(n1083), .A2(n1084), .ZN(n1077) );
NAND2_X1 U772 ( .A1(n1085), .A2(n1080), .ZN(n1084) );
XOR2_X1 U773 ( .A(n1086), .B(n1087), .Z(n1085) );
OR3_X1 U774 ( .A1(n1082), .A2(n1087), .A3(n1080), .ZN(n1083) );
XNOR2_X1 U775 ( .A(n1088), .B(n1089), .ZN(n1087) );
XOR2_X1 U776 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U777 ( .A1(KEYINPUT63), .A2(n1092), .ZN(n1090) );
XNOR2_X1 U778 ( .A(n1093), .B(n1094), .ZN(n1088) );
NAND2_X1 U779 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NAND2_X1 U780 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U781 ( .A1(KEYINPUT62), .A2(n1099), .ZN(n1098) );
NAND2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
INV_X1 U783 ( .A(n1102), .ZN(n1097) );
NAND2_X1 U784 ( .A1(G131), .A2(n1103), .ZN(n1095) );
NAND2_X1 U785 ( .A1(n1101), .A2(n1104), .ZN(n1103) );
NAND2_X1 U786 ( .A1(KEYINPUT62), .A2(n1102), .ZN(n1104) );
INV_X1 U787 ( .A(KEYINPUT30), .ZN(n1101) );
NAND2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(G69) );
NAND2_X1 U789 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U790 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U791 ( .A1(G953), .A2(G224), .ZN(n1110) );
INV_X1 U792 ( .A(n1111), .ZN(n1107) );
NAND3_X1 U793 ( .A1(n1112), .A2(n1109), .A3(n1111), .ZN(n1105) );
NAND3_X1 U794 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1111) );
XOR2_X1 U795 ( .A(n1116), .B(KEYINPUT10), .Z(n1115) );
OR2_X1 U796 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U797 ( .A1(n1118), .A2(n1117), .ZN(n1114) );
XNOR2_X1 U798 ( .A(n1119), .B(KEYINPUT49), .ZN(n1117) );
NAND2_X1 U799 ( .A1(G953), .A2(n1120), .ZN(n1113) );
NAND4_X1 U800 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1109) );
AND3_X1 U801 ( .A1(n1020), .A2(n1080), .A3(n1014), .ZN(n1124) );
XNOR2_X1 U802 ( .A(n1125), .B(KEYINPUT12), .ZN(n1123) );
NAND3_X1 U803 ( .A1(G953), .A2(G224), .A3(G898), .ZN(n1112) );
NOR2_X1 U804 ( .A1(n1126), .A2(n1127), .ZN(G66) );
XOR2_X1 U805 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND2_X1 U806 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
INV_X1 U807 ( .A(n1075), .ZN(n1131) );
NOR2_X1 U808 ( .A1(n1126), .A2(n1132), .ZN(G63) );
XOR2_X1 U809 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U810 ( .A(n1135), .B(KEYINPUT36), .Z(n1133) );
NAND2_X1 U811 ( .A1(n1130), .A2(G478), .ZN(n1135) );
NOR2_X1 U812 ( .A1(n1126), .A2(n1136), .ZN(G60) );
XOR2_X1 U813 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U814 ( .A1(n1130), .A2(G475), .ZN(n1137) );
XNOR2_X1 U815 ( .A(G104), .B(n1121), .ZN(G6) );
NOR2_X1 U816 ( .A1(n1126), .A2(n1139), .ZN(G57) );
XOR2_X1 U817 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U818 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NOR2_X1 U819 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XNOR2_X1 U820 ( .A(n1146), .B(KEYINPUT52), .ZN(n1145) );
NOR2_X1 U821 ( .A1(n1147), .A2(n1148), .ZN(n1142) );
XNOR2_X1 U822 ( .A(n1146), .B(KEYINPUT38), .ZN(n1148) );
XOR2_X1 U823 ( .A(n1149), .B(n1150), .Z(n1140) );
NAND2_X1 U824 ( .A1(n1130), .A2(G472), .ZN(n1149) );
NOR2_X1 U825 ( .A1(n1126), .A2(n1151), .ZN(G54) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1151) );
XNOR2_X1 U827 ( .A(n1154), .B(n1155), .ZN(n1153) );
NAND2_X1 U828 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U829 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U830 ( .A1(n1160), .A2(n1161), .ZN(n1156) );
XNOR2_X1 U831 ( .A(n1158), .B(KEYINPUT25), .ZN(n1160) );
XOR2_X1 U832 ( .A(n1162), .B(n1163), .Z(n1152) );
NAND2_X1 U833 ( .A1(n1130), .A2(G469), .ZN(n1162) );
NOR2_X1 U834 ( .A1(n1126), .A2(n1164), .ZN(G51) );
XOR2_X1 U835 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U836 ( .A(n1167), .B(n1168), .Z(n1166) );
XNOR2_X1 U837 ( .A(n1169), .B(n1170), .ZN(n1165) );
XOR2_X1 U838 ( .A(n1171), .B(KEYINPUT17), .Z(n1169) );
NAND2_X1 U839 ( .A1(n1130), .A2(n1172), .ZN(n1171) );
AND2_X1 U840 ( .A1(n1173), .A2(n1174), .ZN(n1130) );
NAND2_X1 U841 ( .A1(n1022), .A2(n1020), .ZN(n1174) );
OR2_X1 U842 ( .A1(n1175), .A2(n1176), .ZN(n1020) );
INV_X1 U843 ( .A(n1177), .ZN(n1176) );
AND3_X1 U844 ( .A1(n1086), .A2(n1125), .A3(n1178), .ZN(n1022) );
AND3_X1 U845 ( .A1(n1121), .A2(n1014), .A3(n1122), .ZN(n1178) );
NAND3_X1 U846 ( .A1(n1042), .A2(n1179), .A3(n1045), .ZN(n1014) );
NAND3_X1 U847 ( .A1(n1042), .A2(n1179), .A3(n1044), .ZN(n1121) );
AND4_X1 U848 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1125) );
AND4_X1 U849 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1086) );
AND4_X1 U850 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187) );
NOR2_X1 U851 ( .A1(n1192), .A2(n1193), .ZN(n1186) );
NOR2_X1 U852 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
XOR2_X1 U853 ( .A(n1196), .B(KEYINPUT11), .Z(n1194) );
INV_X1 U854 ( .A(n1197), .ZN(n1192) );
XNOR2_X1 U855 ( .A(KEYINPUT56), .B(n1198), .ZN(n1173) );
NOR2_X1 U856 ( .A1(n1080), .A2(G952), .ZN(n1126) );
XNOR2_X1 U857 ( .A(G146), .B(n1197), .ZN(G48) );
NAND4_X1 U858 ( .A1(n1199), .A2(n1044), .A3(n1058), .A4(n1053), .ZN(n1197) );
XNOR2_X1 U859 ( .A(G143), .B(n1184), .ZN(G45) );
NAND4_X1 U860 ( .A1(n1200), .A2(n1053), .A3(n1201), .A4(n1073), .ZN(n1184) );
XNOR2_X1 U861 ( .A(G140), .B(n1185), .ZN(G42) );
NAND3_X1 U862 ( .A1(n1032), .A2(n1058), .A3(n1202), .ZN(n1185) );
XNOR2_X1 U863 ( .A(G137), .B(n1191), .ZN(G39) );
NAND4_X1 U864 ( .A1(n1199), .A2(n1032), .A3(n1041), .A4(n1058), .ZN(n1191) );
XNOR2_X1 U865 ( .A(G134), .B(n1190), .ZN(G36) );
NAND3_X1 U866 ( .A1(n1032), .A2(n1045), .A3(n1200), .ZN(n1190) );
INV_X1 U867 ( .A(n1195), .ZN(n1032) );
NAND2_X1 U868 ( .A1(n1203), .A2(n1204), .ZN(G33) );
NAND2_X1 U869 ( .A1(n1205), .A2(n1100), .ZN(n1204) );
XNOR2_X1 U870 ( .A(n1206), .B(KEYINPUT33), .ZN(n1205) );
NAND2_X1 U871 ( .A1(n1207), .A2(G131), .ZN(n1203) );
XOR2_X1 U872 ( .A(KEYINPUT21), .B(n1206), .Z(n1207) );
NOR2_X1 U873 ( .A1(n1196), .A2(n1195), .ZN(n1206) );
NAND2_X1 U874 ( .A1(n1051), .A2(n1208), .ZN(n1195) );
XOR2_X1 U875 ( .A(KEYINPUT40), .B(n1052), .Z(n1208) );
NAND2_X1 U876 ( .A1(n1200), .A2(n1044), .ZN(n1196) );
AND3_X1 U877 ( .A1(n1058), .A2(n1209), .A3(n1040), .ZN(n1200) );
XNOR2_X1 U878 ( .A(G128), .B(n1189), .ZN(G30) );
NAND4_X1 U879 ( .A1(n1199), .A2(n1045), .A3(n1053), .A4(n1177), .ZN(n1189) );
AND3_X1 U880 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1199) );
XNOR2_X1 U881 ( .A(G101), .B(n1212), .ZN(G3) );
NOR2_X1 U882 ( .A1(KEYINPUT41), .A2(n1213), .ZN(n1212) );
NOR2_X1 U883 ( .A1(n1214), .A2(n1175), .ZN(n1213) );
NAND3_X1 U884 ( .A1(n1041), .A2(n1215), .A3(n1040), .ZN(n1175) );
XNOR2_X1 U885 ( .A(n1177), .B(KEYINPUT53), .ZN(n1214) );
XNOR2_X1 U886 ( .A(G125), .B(n1188), .ZN(G27) );
NAND4_X1 U887 ( .A1(n1027), .A2(n1202), .A3(n1053), .A4(n1026), .ZN(n1188) );
AND3_X1 U888 ( .A1(n1216), .A2(n1209), .A3(n1044), .ZN(n1202) );
NAND2_X1 U889 ( .A1(n1034), .A2(n1217), .ZN(n1209) );
NAND4_X1 U890 ( .A1(G953), .A2(G902), .A3(n1218), .A4(n1082), .ZN(n1217) );
INV_X1 U891 ( .A(G900), .ZN(n1082) );
XNOR2_X1 U892 ( .A(G122), .B(n1180), .ZN(G24) );
NAND4_X1 U893 ( .A1(n1219), .A2(n1042), .A3(n1201), .A4(n1073), .ZN(n1180) );
AND2_X1 U894 ( .A1(n1062), .A2(n1220), .ZN(n1042) );
XNOR2_X1 U895 ( .A(G119), .B(n1181), .ZN(G21) );
NAND4_X1 U896 ( .A1(n1211), .A2(n1219), .A3(n1041), .A4(n1210), .ZN(n1181) );
XNOR2_X1 U897 ( .A(G116), .B(n1182), .ZN(G18) );
NAND3_X1 U898 ( .A1(n1040), .A2(n1045), .A3(n1219), .ZN(n1182) );
NOR2_X1 U899 ( .A1(n1073), .A2(n1221), .ZN(n1045) );
XNOR2_X1 U900 ( .A(G113), .B(n1183), .ZN(G15) );
NAND3_X1 U901 ( .A1(n1044), .A2(n1040), .A3(n1219), .ZN(n1183) );
AND3_X1 U902 ( .A1(n1215), .A2(n1026), .A3(n1027), .ZN(n1219) );
AND2_X1 U903 ( .A1(n1211), .A2(n1220), .ZN(n1040) );
XNOR2_X1 U904 ( .A(KEYINPUT31), .B(n1210), .ZN(n1220) );
XOR2_X1 U905 ( .A(n1062), .B(KEYINPUT8), .Z(n1211) );
AND2_X1 U906 ( .A1(n1221), .A2(n1073), .ZN(n1044) );
INV_X1 U907 ( .A(n1201), .ZN(n1221) );
XNOR2_X1 U908 ( .A(G110), .B(n1122), .ZN(G12) );
NAND2_X1 U909 ( .A1(n1035), .A2(n1179), .ZN(n1122) );
AND2_X1 U910 ( .A1(n1215), .A2(n1177), .ZN(n1179) );
XOR2_X1 U911 ( .A(n1058), .B(KEYINPUT15), .Z(n1177) );
NOR2_X1 U912 ( .A1(n1027), .A2(n1057), .ZN(n1058) );
INV_X1 U913 ( .A(n1026), .ZN(n1057) );
NAND2_X1 U914 ( .A1(G221), .A2(n1222), .ZN(n1026) );
XOR2_X1 U915 ( .A(n1070), .B(G469), .Z(n1027) );
NAND2_X1 U916 ( .A1(n1223), .A2(n1198), .ZN(n1070) );
XOR2_X1 U917 ( .A(n1224), .B(n1225), .Z(n1223) );
XNOR2_X1 U918 ( .A(n1163), .B(n1159), .ZN(n1225) );
INV_X1 U919 ( .A(n1161), .ZN(n1159) );
XNOR2_X1 U920 ( .A(n1226), .B(n1227), .ZN(n1161) );
XNOR2_X1 U921 ( .A(n1228), .B(n1229), .ZN(n1227) );
NOR2_X1 U922 ( .A1(G107), .A2(KEYINPUT14), .ZN(n1229) );
NOR2_X1 U923 ( .A1(n1081), .A2(G953), .ZN(n1163) );
INV_X1 U924 ( .A(G227), .ZN(n1081) );
XNOR2_X1 U925 ( .A(n1158), .B(n1230), .ZN(n1224) );
NOR2_X1 U926 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NOR3_X1 U927 ( .A1(KEYINPUT34), .A2(G110), .A3(n1094), .ZN(n1232) );
NOR2_X1 U928 ( .A1(n1154), .A2(n1233), .ZN(n1231) );
INV_X1 U929 ( .A(KEYINPUT34), .ZN(n1233) );
XNOR2_X1 U930 ( .A(G110), .B(n1094), .ZN(n1154) );
INV_X1 U931 ( .A(G140), .ZN(n1094) );
XOR2_X1 U932 ( .A(n1091), .B(n1234), .Z(n1158) );
XNOR2_X1 U933 ( .A(n1235), .B(n1236), .ZN(n1091) );
XNOR2_X1 U934 ( .A(KEYINPUT20), .B(n1237), .ZN(n1235) );
NOR2_X1 U935 ( .A1(G128), .A2(KEYINPUT55), .ZN(n1237) );
AND2_X1 U936 ( .A1(n1053), .A2(n1238), .ZN(n1215) );
NAND2_X1 U937 ( .A1(n1034), .A2(n1239), .ZN(n1238) );
NAND4_X1 U938 ( .A1(G953), .A2(G902), .A3(n1218), .A4(n1120), .ZN(n1239) );
INV_X1 U939 ( .A(G898), .ZN(n1120) );
NAND3_X1 U940 ( .A1(n1024), .A2(n1218), .A3(G952), .ZN(n1034) );
NAND2_X1 U941 ( .A1(G237), .A2(G234), .ZN(n1218) );
XNOR2_X1 U942 ( .A(G953), .B(KEYINPUT60), .ZN(n1024) );
NOR2_X1 U943 ( .A1(n1240), .A2(n1051), .ZN(n1053) );
XOR2_X1 U944 ( .A(n1241), .B(n1172), .Z(n1051) );
AND2_X1 U945 ( .A1(G210), .A2(n1242), .ZN(n1172) );
NAND2_X1 U946 ( .A1(n1243), .A2(n1198), .ZN(n1241) );
XOR2_X1 U947 ( .A(n1244), .B(n1167), .Z(n1243) );
XNOR2_X1 U948 ( .A(n1119), .B(n1118), .ZN(n1167) );
XNOR2_X1 U949 ( .A(G110), .B(G122), .ZN(n1118) );
XNOR2_X1 U950 ( .A(n1147), .B(n1245), .ZN(n1119) );
XNOR2_X1 U951 ( .A(G101), .B(n1246), .ZN(n1245) );
NAND2_X1 U952 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND2_X1 U953 ( .A1(G107), .A2(n1226), .ZN(n1248) );
XOR2_X1 U954 ( .A(n1249), .B(KEYINPUT24), .Z(n1247) );
OR2_X1 U955 ( .A1(n1226), .A2(G107), .ZN(n1249) );
NAND3_X1 U956 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1244) );
NAND2_X1 U957 ( .A1(KEYINPUT7), .A2(n1253), .ZN(n1252) );
OR3_X1 U958 ( .A1(n1253), .A2(KEYINPUT7), .A3(n1254), .ZN(n1251) );
NAND2_X1 U959 ( .A1(n1254), .A2(n1255), .ZN(n1250) );
NAND2_X1 U960 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
INV_X1 U961 ( .A(KEYINPUT7), .ZN(n1257) );
XNOR2_X1 U962 ( .A(n1253), .B(KEYINPUT42), .ZN(n1256) );
XNOR2_X1 U963 ( .A(n1168), .B(KEYINPUT4), .ZN(n1253) );
XOR2_X1 U964 ( .A(n1258), .B(n1092), .Z(n1168) );
XNOR2_X1 U965 ( .A(n1170), .B(KEYINPUT23), .ZN(n1254) );
NAND2_X1 U966 ( .A1(G224), .A2(n1080), .ZN(n1170) );
XNOR2_X1 U967 ( .A(KEYINPUT40), .B(n1052), .ZN(n1240) );
AND2_X1 U968 ( .A1(n1259), .A2(n1242), .ZN(n1052) );
NAND2_X1 U969 ( .A1(n1260), .A2(n1198), .ZN(n1242) );
XOR2_X1 U970 ( .A(KEYINPUT26), .B(G214), .Z(n1259) );
AND2_X1 U971 ( .A1(n1041), .A2(n1216), .ZN(n1035) );
AND2_X1 U972 ( .A1(n1261), .A2(n1210), .ZN(n1216) );
NAND2_X1 U973 ( .A1(n1262), .A2(n1263), .ZN(n1210) );
NAND2_X1 U974 ( .A1(n1076), .A2(n1075), .ZN(n1263) );
XOR2_X1 U975 ( .A(KEYINPUT46), .B(n1264), .Z(n1262) );
NOR2_X1 U976 ( .A1(n1076), .A2(n1075), .ZN(n1264) );
NAND2_X1 U977 ( .A1(G217), .A2(n1222), .ZN(n1075) );
NAND2_X1 U978 ( .A1(G234), .A2(n1198), .ZN(n1222) );
AND2_X1 U979 ( .A1(n1129), .A2(n1198), .ZN(n1076) );
XOR2_X1 U980 ( .A(n1265), .B(n1266), .Z(n1129) );
XOR2_X1 U981 ( .A(n1267), .B(n1268), .Z(n1266) );
NAND2_X1 U982 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
NAND2_X1 U983 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND2_X1 U984 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
OR2_X1 U985 ( .A1(n1275), .A2(KEYINPUT48), .ZN(n1274) );
INV_X1 U986 ( .A(KEYINPUT16), .ZN(n1273) );
NAND2_X1 U987 ( .A1(n1275), .A2(n1276), .ZN(n1269) );
NAND2_X1 U988 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
OR2_X1 U989 ( .A1(n1271), .A2(KEYINPUT16), .ZN(n1278) );
XOR2_X1 U990 ( .A(n1279), .B(n1280), .Z(n1271) );
INV_X1 U991 ( .A(KEYINPUT48), .ZN(n1277) );
XOR2_X1 U992 ( .A(n1281), .B(n1282), .Z(n1275) );
NOR2_X1 U993 ( .A1(KEYINPUT5), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U994 ( .A(G119), .B(G128), .ZN(n1283) );
XNOR2_X1 U995 ( .A(G110), .B(KEYINPUT2), .ZN(n1281) );
NAND2_X1 U996 ( .A1(G221), .A2(n1284), .ZN(n1267) );
NAND2_X1 U997 ( .A1(KEYINPUT37), .A2(n1285), .ZN(n1265) );
INV_X1 U998 ( .A(G137), .ZN(n1285) );
XOR2_X1 U999 ( .A(n1062), .B(KEYINPUT18), .Z(n1261) );
XOR2_X1 U1000 ( .A(n1286), .B(G472), .Z(n1062) );
NAND2_X1 U1001 ( .A1(n1287), .A2(n1198), .ZN(n1286) );
XOR2_X1 U1002 ( .A(n1288), .B(n1289), .Z(n1287) );
XNOR2_X1 U1003 ( .A(n1150), .B(n1146), .ZN(n1289) );
XNOR2_X1 U1004 ( .A(n1290), .B(n1234), .ZN(n1146) );
XNOR2_X1 U1005 ( .A(n1291), .B(n1292), .ZN(n1234) );
XNOR2_X1 U1006 ( .A(KEYINPUT43), .B(n1100), .ZN(n1292) );
NAND2_X1 U1007 ( .A1(n1293), .A2(n1294), .ZN(n1291) );
NAND2_X1 U1008 ( .A1(n1102), .A2(n1295), .ZN(n1294) );
XOR2_X1 U1009 ( .A(G137), .B(n1296), .Z(n1102) );
OR3_X1 U1010 ( .A1(n1296), .A2(G137), .A3(n1295), .ZN(n1293) );
INV_X1 U1011 ( .A(KEYINPUT0), .ZN(n1295) );
XOR2_X1 U1012 ( .A(n1258), .B(KEYINPUT61), .Z(n1290) );
NAND2_X1 U1013 ( .A1(n1297), .A2(n1298), .ZN(n1258) );
NAND2_X1 U1014 ( .A1(G128), .A2(n1236), .ZN(n1298) );
XOR2_X1 U1015 ( .A(n1299), .B(KEYINPUT19), .Z(n1297) );
OR2_X1 U1016 ( .A1(n1236), .A2(G128), .ZN(n1299) );
XNOR2_X1 U1017 ( .A(G143), .B(n1280), .ZN(n1236) );
INV_X1 U1018 ( .A(G146), .ZN(n1280) );
XOR2_X1 U1019 ( .A(n1300), .B(n1228), .Z(n1150) );
INV_X1 U1020 ( .A(G101), .ZN(n1228) );
NAND3_X1 U1021 ( .A1(n1260), .A2(n1080), .A3(G210), .ZN(n1300) );
XNOR2_X1 U1022 ( .A(KEYINPUT44), .B(n1301), .ZN(n1288) );
NOR2_X1 U1023 ( .A1(KEYINPUT27), .A2(n1144), .ZN(n1301) );
INV_X1 U1024 ( .A(n1147), .ZN(n1144) );
XOR2_X1 U1025 ( .A(G113), .B(n1302), .Z(n1147) );
XOR2_X1 U1026 ( .A(G119), .B(G116), .Z(n1302) );
NOR2_X1 U1027 ( .A1(n1201), .A2(n1073), .ZN(n1041) );
XNOR2_X1 U1028 ( .A(n1303), .B(G475), .ZN(n1073) );
NAND2_X1 U1029 ( .A1(n1138), .A2(n1198), .ZN(n1303) );
XOR2_X1 U1030 ( .A(n1304), .B(n1305), .Z(n1138) );
XOR2_X1 U1031 ( .A(n1279), .B(n1306), .Z(n1305) );
XOR2_X1 U1032 ( .A(n1307), .B(n1226), .Z(n1306) );
XNOR2_X1 U1033 ( .A(G104), .B(KEYINPUT57), .ZN(n1226) );
NAND2_X1 U1034 ( .A1(n1308), .A2(KEYINPUT28), .ZN(n1307) );
XNOR2_X1 U1035 ( .A(G122), .B(n1309), .ZN(n1308) );
NOR2_X1 U1036 ( .A1(KEYINPUT13), .A2(n1310), .ZN(n1309) );
XOR2_X1 U1037 ( .A(KEYINPUT9), .B(G113), .Z(n1310) );
XOR2_X1 U1038 ( .A(G140), .B(n1092), .Z(n1279) );
XOR2_X1 U1039 ( .A(G125), .B(KEYINPUT3), .Z(n1092) );
XOR2_X1 U1040 ( .A(n1311), .B(n1312), .Z(n1304) );
XNOR2_X1 U1041 ( .A(KEYINPUT51), .B(n1100), .ZN(n1312) );
INV_X1 U1042 ( .A(G131), .ZN(n1100) );
XNOR2_X1 U1043 ( .A(n1313), .B(n1314), .ZN(n1311) );
NOR2_X1 U1044 ( .A1(G146), .A2(KEYINPUT22), .ZN(n1314) );
NOR2_X1 U1045 ( .A1(KEYINPUT6), .A2(n1315), .ZN(n1313) );
NOR2_X1 U1046 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XOR2_X1 U1047 ( .A(n1318), .B(KEYINPUT39), .Z(n1317) );
NAND2_X1 U1048 ( .A1(G143), .A2(n1319), .ZN(n1318) );
NOR2_X1 U1049 ( .A1(G143), .A2(n1319), .ZN(n1316) );
AND3_X1 U1050 ( .A1(n1260), .A2(n1080), .A3(G214), .ZN(n1319) );
INV_X1 U1051 ( .A(G237), .ZN(n1260) );
XOR2_X1 U1052 ( .A(n1068), .B(n1069), .Z(n1201) );
INV_X1 U1053 ( .A(G478), .ZN(n1069) );
NAND2_X1 U1054 ( .A1(n1134), .A2(n1198), .ZN(n1068) );
INV_X1 U1055 ( .A(G902), .ZN(n1198) );
XNOR2_X1 U1056 ( .A(n1320), .B(n1321), .ZN(n1134) );
NOR2_X1 U1057 ( .A1(KEYINPUT54), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1058 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1059 ( .A(n1325), .B(n1296), .Z(n1324) );
XOR2_X1 U1060 ( .A(G134), .B(KEYINPUT50), .Z(n1296) );
XNOR2_X1 U1061 ( .A(G107), .B(n1326), .ZN(n1325) );
NOR2_X1 U1062 ( .A1(KEYINPUT45), .A2(n1327), .ZN(n1326) );
XNOR2_X1 U1063 ( .A(G122), .B(KEYINPUT1), .ZN(n1327) );
XOR2_X1 U1064 ( .A(n1328), .B(n1329), .Z(n1323) );
XNOR2_X1 U1065 ( .A(KEYINPUT32), .B(n1330), .ZN(n1329) );
INV_X1 U1066 ( .A(G143), .ZN(n1330) );
XNOR2_X1 U1067 ( .A(G116), .B(G128), .ZN(n1328) );
NAND2_X1 U1068 ( .A1(G217), .A2(n1284), .ZN(n1320) );
AND2_X1 U1069 ( .A1(G234), .A2(n1080), .ZN(n1284) );
INV_X1 U1070 ( .A(G953), .ZN(n1080) );
endmodule


