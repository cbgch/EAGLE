//Key = 0011000101011101100001111011000001101011001011101100001111000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
n1408;

XOR2_X1 U769 ( .A(G107), .B(n1068), .Z(G9) );
NOR2_X1 U770 ( .A1(n1069), .A2(n1070), .ZN(G75) );
NOR3_X1 U771 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1070) );
NOR2_X1 U772 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR2_X1 U776 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR3_X1 U777 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1082) );
NOR2_X1 U778 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR3_X1 U780 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1085) );
NOR2_X1 U781 ( .A1(n1094), .A2(n1095), .ZN(n1084) );
NOR2_X1 U782 ( .A1(n1094), .A2(n1096), .ZN(n1080) );
NOR2_X1 U783 ( .A1(n1097), .A2(n1093), .ZN(n1096) );
NOR3_X1 U784 ( .A1(n1088), .A2(n1098), .A3(n1099), .ZN(n1097) );
NOR2_X1 U785 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U786 ( .A1(KEYINPUT35), .A2(n1102), .ZN(n1100) );
AND2_X1 U787 ( .A1(n1103), .A2(n1093), .ZN(n1094) );
NAND4_X1 U788 ( .A1(KEYINPUT35), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1103) );
INV_X1 U789 ( .A(n1101), .ZN(n1104) );
NOR4_X1 U790 ( .A1(n1107), .A2(n1088), .A3(n1083), .A4(n1093), .ZN(n1076) );
INV_X1 U791 ( .A(n1106), .ZN(n1088) );
NOR2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U793 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
XOR2_X1 U794 ( .A(n1112), .B(KEYINPUT17), .Z(n1111) );
NAND3_X1 U795 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1071) );
NAND3_X1 U796 ( .A1(n1116), .A2(n1091), .A3(n1117), .ZN(n1115) );
INV_X1 U797 ( .A(n1079), .ZN(n1117) );
INV_X1 U798 ( .A(KEYINPUT12), .ZN(n1091) );
OR4_X1 U799 ( .A1(n1075), .A2(n1093), .A3(n1083), .A4(n1092), .ZN(n1116) );
XNOR2_X1 U800 ( .A(n1118), .B(KEYINPUT31), .ZN(n1092) );
INV_X1 U801 ( .A(n1119), .ZN(n1093) );
NOR3_X1 U802 ( .A1(n1120), .A2(G953), .A3(G952), .ZN(n1069) );
INV_X1 U803 ( .A(n1113), .ZN(n1120) );
NAND4_X1 U804 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1113) );
NOR4_X1 U805 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1124) );
XOR2_X1 U806 ( .A(n1112), .B(KEYINPUT9), .Z(n1128) );
XOR2_X1 U807 ( .A(n1129), .B(n1130), .Z(n1127) );
XOR2_X1 U808 ( .A(KEYINPUT62), .B(KEYINPUT13), .Z(n1130) );
XOR2_X1 U809 ( .A(n1131), .B(G478), .Z(n1129) );
NOR2_X1 U810 ( .A1(n1132), .A2(n1133), .ZN(n1126) );
NOR2_X1 U811 ( .A1(G902), .A2(n1134), .ZN(n1132) );
NOR2_X1 U812 ( .A1(n1083), .A2(n1135), .ZN(n1123) );
XOR2_X1 U813 ( .A(n1136), .B(KEYINPUT10), .Z(n1122) );
XNOR2_X1 U814 ( .A(n1137), .B(n1138), .ZN(n1121) );
XOR2_X1 U815 ( .A(n1139), .B(n1140), .Z(G72) );
XOR2_X1 U816 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U817 ( .A1(n1143), .A2(n1114), .ZN(n1142) );
AND2_X1 U818 ( .A1(G227), .A2(G900), .ZN(n1143) );
NOR2_X1 U819 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
XOR2_X1 U820 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U821 ( .A(G140), .B(G125), .Z(n1147) );
NOR2_X1 U822 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
XOR2_X1 U823 ( .A(n1150), .B(KEYINPUT39), .Z(n1149) );
NAND3_X1 U824 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
NOR2_X1 U825 ( .A1(n1154), .A2(n1153), .ZN(n1148) );
XOR2_X1 U826 ( .A(n1155), .B(KEYINPUT16), .Z(n1153) );
AND2_X1 U827 ( .A1(n1152), .A2(n1151), .ZN(n1154) );
NOR2_X1 U828 ( .A1(G900), .A2(n1114), .ZN(n1144) );
NOR2_X1 U829 ( .A1(n1156), .A2(G953), .ZN(n1139) );
XOR2_X1 U830 ( .A(n1157), .B(n1158), .Z(G69) );
NOR2_X1 U831 ( .A1(n1159), .A2(n1114), .ZN(n1158) );
AND2_X1 U832 ( .A1(G224), .A2(G898), .ZN(n1159) );
NOR2_X1 U833 ( .A1(KEYINPUT50), .A2(n1160), .ZN(n1157) );
XOR2_X1 U834 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U835 ( .A1(n1163), .A2(G953), .ZN(n1162) );
NAND3_X1 U836 ( .A1(n1164), .A2(n1165), .A3(KEYINPUT23), .ZN(n1161) );
NAND2_X1 U837 ( .A1(G953), .A2(n1166), .ZN(n1165) );
XOR2_X1 U838 ( .A(n1167), .B(KEYINPUT30), .Z(n1164) );
NAND2_X1 U839 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U840 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NAND2_X1 U841 ( .A1(n1172), .A2(n1173), .ZN(n1168) );
INV_X1 U842 ( .A(n1171), .ZN(n1173) );
XNOR2_X1 U843 ( .A(G122), .B(n1174), .ZN(n1171) );
XOR2_X1 U844 ( .A(n1170), .B(n1175), .Z(n1172) );
XNOR2_X1 U845 ( .A(KEYINPUT61), .B(KEYINPUT0), .ZN(n1175) );
XOR2_X1 U846 ( .A(n1176), .B(n1177), .Z(n1170) );
NOR2_X1 U847 ( .A1(KEYINPUT60), .A2(n1178), .ZN(n1177) );
NOR2_X1 U848 ( .A1(n1179), .A2(n1180), .ZN(G66) );
XNOR2_X1 U849 ( .A(n1181), .B(n1182), .ZN(n1180) );
XNOR2_X1 U850 ( .A(KEYINPUT2), .B(n1183), .ZN(n1182) );
NOR3_X1 U851 ( .A1(n1184), .A2(KEYINPUT19), .A3(n1185), .ZN(n1183) );
NOR2_X1 U852 ( .A1(n1179), .A2(n1186), .ZN(G63) );
NOR3_X1 U853 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1186) );
NOR3_X1 U854 ( .A1(n1190), .A2(n1191), .A3(n1184), .ZN(n1189) );
NOR2_X1 U855 ( .A1(n1192), .A2(n1193), .ZN(n1188) );
INV_X1 U856 ( .A(n1190), .ZN(n1193) );
AND2_X1 U857 ( .A1(n1073), .A2(G478), .ZN(n1192) );
NOR2_X1 U858 ( .A1(n1179), .A2(n1194), .ZN(G60) );
XOR2_X1 U859 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U860 ( .A(KEYINPUT49), .B(n1197), .Z(n1196) );
NOR2_X1 U861 ( .A1(n1133), .A2(n1184), .ZN(n1197) );
XOR2_X1 U862 ( .A(G104), .B(n1198), .Z(G6) );
NOR2_X1 U863 ( .A1(n1179), .A2(n1199), .ZN(G57) );
XOR2_X1 U864 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U865 ( .A(n1202), .B(n1203), .Z(n1201) );
NOR2_X1 U866 ( .A1(KEYINPUT51), .A2(n1204), .ZN(n1202) );
XOR2_X1 U867 ( .A(n1205), .B(n1206), .Z(n1200) );
NOR2_X1 U868 ( .A1(n1207), .A2(n1184), .ZN(n1206) );
INV_X1 U869 ( .A(G472), .ZN(n1207) );
NOR2_X1 U870 ( .A1(n1179), .A2(n1208), .ZN(G54) );
XOR2_X1 U871 ( .A(n1209), .B(n1210), .Z(n1208) );
XOR2_X1 U872 ( .A(n1211), .B(n1212), .Z(n1210) );
NOR2_X1 U873 ( .A1(n1213), .A2(n1184), .ZN(n1212) );
INV_X1 U874 ( .A(G469), .ZN(n1213) );
NAND2_X1 U875 ( .A1(KEYINPUT27), .A2(n1214), .ZN(n1211) );
XOR2_X1 U876 ( .A(n1155), .B(n1215), .Z(n1214) );
NOR2_X1 U877 ( .A1(n1179), .A2(n1216), .ZN(G51) );
XOR2_X1 U878 ( .A(n1217), .B(n1218), .Z(n1216) );
XOR2_X1 U879 ( .A(n1219), .B(n1220), .Z(n1218) );
XOR2_X1 U880 ( .A(KEYINPUT55), .B(KEYINPUT21), .Z(n1220) );
NOR2_X1 U881 ( .A1(n1138), .A2(n1184), .ZN(n1219) );
NAND2_X1 U882 ( .A1(G902), .A2(n1073), .ZN(n1184) );
NAND2_X1 U883 ( .A1(n1163), .A2(n1156), .ZN(n1073) );
AND4_X1 U884 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1156) );
AND4_X1 U885 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1224) );
NAND2_X1 U886 ( .A1(n1229), .A2(n1230), .ZN(n1223) );
NAND2_X1 U887 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND2_X1 U888 ( .A1(n1233), .A2(n1090), .ZN(n1232) );
XOR2_X1 U889 ( .A(n1234), .B(KEYINPUT11), .Z(n1233) );
NAND2_X1 U890 ( .A1(n1235), .A2(n1089), .ZN(n1231) );
AND4_X1 U891 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1163) );
NOR4_X1 U892 ( .A1(n1240), .A2(n1068), .A3(n1241), .A4(n1242), .ZN(n1239) );
INV_X1 U893 ( .A(n1243), .ZN(n1242) );
AND3_X1 U894 ( .A1(n1106), .A2(n1089), .A3(n1244), .ZN(n1068) );
INV_X1 U895 ( .A(n1245), .ZN(n1240) );
NOR2_X1 U896 ( .A1(n1246), .A2(n1198), .ZN(n1238) );
AND3_X1 U897 ( .A1(n1244), .A2(n1106), .A3(n1090), .ZN(n1198) );
XOR2_X1 U898 ( .A(n1247), .B(n1248), .Z(n1217) );
NAND2_X1 U899 ( .A1(KEYINPUT15), .A2(n1204), .ZN(n1247) );
NOR2_X1 U900 ( .A1(n1114), .A2(G952), .ZN(n1179) );
NAND2_X1 U901 ( .A1(n1249), .A2(n1250), .ZN(G48) );
OR2_X1 U902 ( .A1(n1251), .A2(G146), .ZN(n1250) );
XOR2_X1 U903 ( .A(n1252), .B(KEYINPUT25), .Z(n1249) );
NAND2_X1 U904 ( .A1(G146), .A2(n1251), .ZN(n1252) );
NAND3_X1 U905 ( .A1(n1235), .A2(n1090), .A3(n1229), .ZN(n1251) );
XOR2_X1 U906 ( .A(n1253), .B(n1221), .Z(G45) );
NAND4_X1 U907 ( .A1(n1229), .A2(n1118), .A3(n1254), .A4(n1255), .ZN(n1221) );
XOR2_X1 U908 ( .A(n1256), .B(n1222), .Z(G42) );
NAND3_X1 U909 ( .A1(n1090), .A2(n1257), .A3(n1258), .ZN(n1222) );
XOR2_X1 U910 ( .A(n1259), .B(n1228), .Z(G39) );
NAND3_X1 U911 ( .A1(n1235), .A2(n1119), .A3(n1258), .ZN(n1228) );
XOR2_X1 U912 ( .A(n1260), .B(n1227), .Z(G36) );
NAND3_X1 U913 ( .A1(n1118), .A2(n1089), .A3(n1258), .ZN(n1227) );
XNOR2_X1 U914 ( .A(G131), .B(n1226), .ZN(G33) );
NAND3_X1 U915 ( .A1(n1090), .A2(n1118), .A3(n1258), .ZN(n1226) );
NOR2_X1 U916 ( .A1(n1261), .A2(n1079), .ZN(n1258) );
NAND2_X1 U917 ( .A1(n1262), .A2(n1112), .ZN(n1079) );
INV_X1 U918 ( .A(n1110), .ZN(n1262) );
XOR2_X1 U919 ( .A(n1263), .B(KEYINPUT29), .Z(n1110) );
NAND3_X1 U920 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(G30) );
NAND4_X1 U921 ( .A1(n1267), .A2(n1268), .A3(n1089), .A4(n1269), .ZN(n1266) );
NOR2_X1 U922 ( .A1(n1234), .A2(n1261), .ZN(n1269) );
NAND2_X1 U923 ( .A1(n1270), .A2(n1271), .ZN(n1268) );
XOR2_X1 U924 ( .A(KEYINPUT4), .B(G128), .Z(n1270) );
XOR2_X1 U925 ( .A(KEYINPUT52), .B(n1109), .Z(n1267) );
NAND2_X1 U926 ( .A1(KEYINPUT20), .A2(n1272), .ZN(n1265) );
NAND3_X1 U927 ( .A1(n1273), .A2(n1271), .A3(G128), .ZN(n1264) );
INV_X1 U928 ( .A(KEYINPUT20), .ZN(n1271) );
NAND4_X1 U929 ( .A1(n1235), .A2(n1089), .A3(n1274), .A4(n1275), .ZN(n1273) );
OR2_X1 U930 ( .A1(n1229), .A2(KEYINPUT52), .ZN(n1275) );
NOR2_X1 U931 ( .A1(n1261), .A2(n1276), .ZN(n1229) );
NAND2_X1 U932 ( .A1(KEYINPUT52), .A2(n1277), .ZN(n1274) );
OR2_X1 U933 ( .A1(n1261), .A2(n1109), .ZN(n1277) );
NAND3_X1 U934 ( .A1(n1278), .A2(n1101), .A3(n1102), .ZN(n1261) );
XOR2_X1 U935 ( .A(G101), .B(n1246), .Z(G3) );
AND3_X1 U936 ( .A1(n1118), .A2(n1244), .A3(n1119), .ZN(n1246) );
XOR2_X1 U937 ( .A(n1279), .B(n1225), .Z(G27) );
NAND4_X1 U938 ( .A1(n1109), .A2(n1278), .A3(n1098), .A4(n1280), .ZN(n1225) );
AND2_X1 U939 ( .A1(n1257), .A2(n1090), .ZN(n1280) );
NAND2_X1 U940 ( .A1(n1075), .A2(n1281), .ZN(n1278) );
NAND4_X1 U941 ( .A1(G953), .A2(G902), .A3(n1282), .A4(n1283), .ZN(n1281) );
INV_X1 U942 ( .A(G900), .ZN(n1283) );
XNOR2_X1 U943 ( .A(G122), .B(n1236), .ZN(G24) );
NAND4_X1 U944 ( .A1(n1284), .A2(n1106), .A3(n1254), .A4(n1255), .ZN(n1236) );
NOR2_X1 U945 ( .A1(n1135), .A2(n1285), .ZN(n1106) );
XOR2_X1 U946 ( .A(n1286), .B(n1237), .Z(G21) );
NAND3_X1 U947 ( .A1(n1119), .A2(n1284), .A3(n1235), .ZN(n1237) );
INV_X1 U948 ( .A(n1234), .ZN(n1235) );
NAND2_X1 U949 ( .A1(n1285), .A2(n1135), .ZN(n1234) );
XOR2_X1 U950 ( .A(n1287), .B(n1245), .Z(G18) );
NAND3_X1 U951 ( .A1(n1284), .A2(n1089), .A3(n1118), .ZN(n1245) );
AND2_X1 U952 ( .A1(n1288), .A2(n1254), .ZN(n1089) );
XNOR2_X1 U953 ( .A(n1289), .B(KEYINPUT57), .ZN(n1254) );
XOR2_X1 U954 ( .A(n1290), .B(n1243), .Z(G15) );
NAND3_X1 U955 ( .A1(n1118), .A2(n1284), .A3(n1090), .ZN(n1243) );
NOR2_X1 U956 ( .A1(n1289), .A2(n1288), .ZN(n1090) );
AND2_X1 U957 ( .A1(n1098), .A2(n1291), .ZN(n1284) );
INV_X1 U958 ( .A(n1083), .ZN(n1098) );
NAND2_X1 U959 ( .A1(n1105), .A2(n1101), .ZN(n1083) );
NOR2_X1 U960 ( .A1(n1292), .A2(n1135), .ZN(n1118) );
XOR2_X1 U961 ( .A(n1241), .B(n1293), .Z(G12) );
NOR2_X1 U962 ( .A1(KEYINPUT63), .A2(n1294), .ZN(n1293) );
AND3_X1 U963 ( .A1(n1257), .A2(n1244), .A3(n1119), .ZN(n1241) );
NOR2_X1 U964 ( .A1(n1255), .A2(n1289), .ZN(n1119) );
NAND2_X1 U965 ( .A1(n1295), .A2(n1296), .ZN(n1289) );
NAND2_X1 U966 ( .A1(G478), .A2(n1131), .ZN(n1296) );
XOR2_X1 U967 ( .A(n1297), .B(KEYINPUT14), .Z(n1295) );
NAND2_X1 U968 ( .A1(n1187), .A2(n1191), .ZN(n1297) );
INV_X1 U969 ( .A(G478), .ZN(n1191) );
INV_X1 U970 ( .A(n1131), .ZN(n1187) );
NAND2_X1 U971 ( .A1(n1190), .A2(n1298), .ZN(n1131) );
XOR2_X1 U972 ( .A(n1299), .B(n1300), .Z(n1190) );
XOR2_X1 U973 ( .A(G128), .B(n1301), .Z(n1300) );
XOR2_X1 U974 ( .A(G143), .B(G134), .Z(n1301) );
XOR2_X1 U975 ( .A(n1302), .B(n1303), .Z(n1299) );
NOR2_X1 U976 ( .A1(KEYINPUT47), .A2(n1304), .ZN(n1303) );
XOR2_X1 U977 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U978 ( .A(G122), .B(n1287), .Z(n1306) );
NAND2_X1 U979 ( .A1(KEYINPUT34), .A2(G107), .ZN(n1305) );
NAND2_X1 U980 ( .A1(n1307), .A2(G217), .ZN(n1302) );
INV_X1 U981 ( .A(n1288), .ZN(n1255) );
NOR2_X1 U982 ( .A1(n1308), .A2(n1125), .ZN(n1288) );
NOR3_X1 U983 ( .A1(G475), .A2(G902), .A3(n1134), .ZN(n1125) );
INV_X1 U984 ( .A(n1195), .ZN(n1134) );
AND2_X1 U985 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
NAND2_X1 U986 ( .A1(n1195), .A2(n1298), .ZN(n1310) );
XOR2_X1 U987 ( .A(n1311), .B(n1312), .Z(n1195) );
XNOR2_X1 U988 ( .A(n1313), .B(n1314), .ZN(n1312) );
XOR2_X1 U989 ( .A(n1315), .B(n1316), .Z(n1314) );
NAND2_X1 U990 ( .A1(KEYINPUT44), .A2(n1317), .ZN(n1315) );
XOR2_X1 U991 ( .A(n1318), .B(n1319), .Z(n1311) );
NOR2_X1 U992 ( .A1(G140), .A2(KEYINPUT37), .ZN(n1319) );
XOR2_X1 U993 ( .A(n1320), .B(G113), .Z(n1318) );
NAND2_X1 U994 ( .A1(KEYINPUT33), .A2(n1321), .ZN(n1320) );
XOR2_X1 U995 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U996 ( .A(G131), .B(n1253), .Z(n1323) );
NAND2_X1 U997 ( .A1(n1324), .A2(G214), .ZN(n1322) );
XOR2_X1 U998 ( .A(n1133), .B(KEYINPUT36), .Z(n1309) );
INV_X1 U999 ( .A(G475), .ZN(n1133) );
AND3_X1 U1000 ( .A1(n1102), .A2(n1101), .A3(n1291), .ZN(n1244) );
AND2_X1 U1001 ( .A1(n1109), .A2(n1325), .ZN(n1291) );
NAND2_X1 U1002 ( .A1(n1075), .A2(n1326), .ZN(n1325) );
NAND4_X1 U1003 ( .A1(G953), .A2(G902), .A3(n1282), .A4(n1166), .ZN(n1326) );
INV_X1 U1004 ( .A(G898), .ZN(n1166) );
NAND3_X1 U1005 ( .A1(n1282), .A2(n1114), .A3(G952), .ZN(n1075) );
NAND2_X1 U1006 ( .A1(G237), .A2(G234), .ZN(n1282) );
INV_X1 U1007 ( .A(n1276), .ZN(n1109) );
NAND2_X1 U1008 ( .A1(n1263), .A2(n1112), .ZN(n1276) );
NAND2_X1 U1009 ( .A1(G214), .A2(n1327), .ZN(n1112) );
XNOR2_X1 U1010 ( .A(n1328), .B(n1137), .ZN(n1263) );
NAND2_X1 U1011 ( .A1(n1329), .A2(n1298), .ZN(n1137) );
XOR2_X1 U1012 ( .A(n1204), .B(n1248), .Z(n1329) );
XNOR2_X1 U1013 ( .A(n1330), .B(n1331), .ZN(n1248) );
XOR2_X1 U1014 ( .A(n1313), .B(n1174), .Z(n1331) );
XOR2_X1 U1015 ( .A(G110), .B(KEYINPUT45), .Z(n1174) );
XOR2_X1 U1016 ( .A(G122), .B(G125), .Z(n1313) );
XOR2_X1 U1017 ( .A(n1332), .B(n1333), .Z(n1330) );
NOR2_X1 U1018 ( .A1(KEYINPUT58), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1019 ( .A(n1335), .B(n1178), .Z(n1334) );
XOR2_X1 U1020 ( .A(n1336), .B(n1337), .Z(n1178) );
XOR2_X1 U1021 ( .A(KEYINPUT38), .B(G107), .Z(n1337) );
XOR2_X1 U1022 ( .A(n1338), .B(n1316), .Z(n1336) );
NAND2_X1 U1023 ( .A1(KEYINPUT22), .A2(n1176), .ZN(n1335) );
XOR2_X1 U1024 ( .A(n1290), .B(n1339), .Z(n1176) );
NOR2_X1 U1025 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
XOR2_X1 U1026 ( .A(KEYINPUT41), .B(n1342), .Z(n1341) );
NOR2_X1 U1027 ( .A1(G116), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1028 ( .A(KEYINPUT42), .B(G119), .Z(n1343) );
NAND2_X1 U1029 ( .A1(G224), .A2(n1114), .ZN(n1332) );
NAND2_X1 U1030 ( .A1(KEYINPUT3), .A2(n1138), .ZN(n1328) );
NAND2_X1 U1031 ( .A1(G210), .A2(n1327), .ZN(n1138) );
NAND2_X1 U1032 ( .A1(n1344), .A2(n1298), .ZN(n1327) );
INV_X1 U1033 ( .A(G237), .ZN(n1344) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1345), .ZN(n1101) );
INV_X1 U1035 ( .A(n1105), .ZN(n1102) );
XOR2_X1 U1036 ( .A(n1346), .B(G469), .Z(n1105) );
NAND2_X1 U1037 ( .A1(n1347), .A2(n1298), .ZN(n1346) );
XOR2_X1 U1038 ( .A(n1348), .B(n1209), .Z(n1347) );
XOR2_X1 U1039 ( .A(n1349), .B(n1350), .Z(n1209) );
XOR2_X1 U1040 ( .A(n1205), .B(n1351), .Z(n1350) );
NAND2_X1 U1041 ( .A1(G227), .A2(n1114), .ZN(n1351) );
XOR2_X1 U1042 ( .A(n1294), .B(G140), .Z(n1349) );
INV_X1 U1043 ( .A(G110), .ZN(n1294) );
NAND3_X1 U1044 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1348) );
NAND2_X1 U1045 ( .A1(KEYINPUT28), .A2(n1155), .ZN(n1354) );
NAND3_X1 U1046 ( .A1(n1355), .A2(n1356), .A3(n1215), .ZN(n1353) );
INV_X1 U1047 ( .A(n1155), .ZN(n1355) );
NAND2_X1 U1048 ( .A1(n1357), .A2(n1358), .ZN(n1352) );
NAND2_X1 U1049 ( .A1(n1359), .A2(n1356), .ZN(n1358) );
INV_X1 U1050 ( .A(KEYINPUT28), .ZN(n1356) );
XOR2_X1 U1051 ( .A(n1155), .B(KEYINPUT24), .Z(n1359) );
XNOR2_X1 U1052 ( .A(n1360), .B(n1361), .ZN(n1155) );
XOR2_X1 U1053 ( .A(KEYINPUT8), .B(n1362), .Z(n1361) );
INV_X1 U1054 ( .A(n1215), .ZN(n1357) );
XOR2_X1 U1055 ( .A(n1363), .B(G101), .Z(n1215) );
NAND3_X1 U1056 ( .A1(n1364), .A2(n1365), .A3(n1366), .ZN(n1363) );
NAND2_X1 U1057 ( .A1(KEYINPUT6), .A2(n1367), .ZN(n1366) );
NAND3_X1 U1058 ( .A1(n1316), .A2(n1368), .A3(G107), .ZN(n1365) );
NAND2_X1 U1059 ( .A1(n1369), .A2(n1370), .ZN(n1364) );
INV_X1 U1060 ( .A(G107), .ZN(n1370) );
NAND2_X1 U1061 ( .A1(n1371), .A2(n1368), .ZN(n1369) );
INV_X1 U1062 ( .A(KEYINPUT6), .ZN(n1368) );
XOR2_X1 U1063 ( .A(KEYINPUT18), .B(n1316), .Z(n1371) );
INV_X1 U1064 ( .A(n1367), .ZN(n1316) );
XNOR2_X1 U1065 ( .A(G104), .B(KEYINPUT7), .ZN(n1367) );
INV_X1 U1066 ( .A(n1095), .ZN(n1257) );
NAND2_X1 U1067 ( .A1(n1292), .A2(n1135), .ZN(n1095) );
XNOR2_X1 U1068 ( .A(n1372), .B(n1373), .ZN(n1135) );
NOR2_X1 U1069 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
XOR2_X1 U1070 ( .A(n1185), .B(KEYINPUT40), .Z(n1375) );
INV_X1 U1071 ( .A(G217), .ZN(n1185) );
INV_X1 U1072 ( .A(n1345), .ZN(n1374) );
NAND2_X1 U1073 ( .A1(G234), .A2(n1298), .ZN(n1345) );
NAND2_X1 U1074 ( .A1(n1181), .A2(n1298), .ZN(n1372) );
XNOR2_X1 U1075 ( .A(n1376), .B(n1377), .ZN(n1181) );
XOR2_X1 U1076 ( .A(n1378), .B(n1379), .Z(n1377) );
XOR2_X1 U1077 ( .A(G137), .B(G110), .Z(n1379) );
NOR3_X1 U1078 ( .A1(KEYINPUT53), .A2(n1380), .A3(n1381), .ZN(n1378) );
NOR3_X1 U1079 ( .A1(KEYINPUT54), .A2(G119), .A3(n1272), .ZN(n1381) );
INV_X1 U1080 ( .A(G128), .ZN(n1272) );
NOR2_X1 U1081 ( .A1(n1382), .A2(n1383), .ZN(n1380) );
INV_X1 U1082 ( .A(KEYINPUT54), .ZN(n1383) );
XOR2_X1 U1083 ( .A(G128), .B(G119), .Z(n1382) );
XOR2_X1 U1084 ( .A(n1384), .B(n1385), .Z(n1376) );
AND2_X1 U1085 ( .A1(G221), .A2(n1307), .ZN(n1385) );
AND2_X1 U1086 ( .A1(G234), .A2(n1114), .ZN(n1307) );
INV_X1 U1087 ( .A(G953), .ZN(n1114) );
NAND2_X1 U1088 ( .A1(n1386), .A2(n1387), .ZN(n1384) );
NAND2_X1 U1089 ( .A1(n1388), .A2(n1317), .ZN(n1387) );
XOR2_X1 U1090 ( .A(KEYINPUT26), .B(n1389), .Z(n1386) );
NOR2_X1 U1091 ( .A1(n1317), .A2(n1388), .ZN(n1389) );
XNOR2_X1 U1092 ( .A(n1390), .B(n1391), .ZN(n1388) );
NOR2_X1 U1093 ( .A1(KEYINPUT59), .A2(n1279), .ZN(n1391) );
INV_X1 U1094 ( .A(G125), .ZN(n1279) );
XOR2_X1 U1095 ( .A(n1256), .B(KEYINPUT46), .Z(n1390) );
INV_X1 U1096 ( .A(G140), .ZN(n1256) );
INV_X1 U1097 ( .A(n1285), .ZN(n1292) );
XOR2_X1 U1098 ( .A(n1136), .B(KEYINPUT56), .Z(n1285) );
XOR2_X1 U1099 ( .A(n1392), .B(G472), .Z(n1136) );
NAND2_X1 U1100 ( .A1(n1393), .A2(n1298), .ZN(n1392) );
INV_X1 U1101 ( .A(G902), .ZN(n1298) );
XOR2_X1 U1102 ( .A(n1394), .B(n1395), .Z(n1393) );
XOR2_X1 U1103 ( .A(n1396), .B(n1203), .Z(n1395) );
XNOR2_X1 U1104 ( .A(n1397), .B(n1398), .ZN(n1203) );
XOR2_X1 U1105 ( .A(n1338), .B(n1399), .Z(n1398) );
NAND3_X1 U1106 ( .A1(n1400), .A2(n1401), .A3(n1402), .ZN(n1399) );
NAND2_X1 U1107 ( .A1(n1340), .A2(n1290), .ZN(n1402) );
NOR2_X1 U1108 ( .A1(n1287), .A2(G119), .ZN(n1340) );
NAND3_X1 U1109 ( .A1(G113), .A2(n1287), .A3(n1286), .ZN(n1401) );
INV_X1 U1110 ( .A(G119), .ZN(n1286) );
INV_X1 U1111 ( .A(G116), .ZN(n1287) );
NAND2_X1 U1112 ( .A1(G119), .A2(n1403), .ZN(n1400) );
XOR2_X1 U1113 ( .A(n1290), .B(G116), .Z(n1403) );
INV_X1 U1114 ( .A(G113), .ZN(n1290) );
INV_X1 U1115 ( .A(G101), .ZN(n1338) );
NAND2_X1 U1116 ( .A1(n1324), .A2(G210), .ZN(n1397) );
NOR2_X1 U1117 ( .A1(G953), .A2(G237), .ZN(n1324) );
NOR2_X1 U1118 ( .A1(KEYINPUT43), .A2(n1204), .ZN(n1396) );
XNOR2_X1 U1119 ( .A(n1404), .B(n1362), .ZN(n1204) );
XOR2_X1 U1120 ( .A(G128), .B(KEYINPUT32), .Z(n1362) );
NAND2_X1 U1121 ( .A1(KEYINPUT48), .A2(n1360), .ZN(n1404) );
XOR2_X1 U1122 ( .A(n1253), .B(n1317), .Z(n1360) );
INV_X1 U1123 ( .A(G146), .ZN(n1317) );
INV_X1 U1124 ( .A(G143), .ZN(n1253) );
XNOR2_X1 U1125 ( .A(KEYINPUT5), .B(n1205), .ZN(n1394) );
NAND3_X1 U1126 ( .A1(n1405), .A2(n1406), .A3(n1151), .ZN(n1205) );
NAND2_X1 U1127 ( .A1(G137), .A2(n1407), .ZN(n1151) );
OR2_X1 U1128 ( .A1(n1152), .A2(KEYINPUT1), .ZN(n1406) );
NAND2_X1 U1129 ( .A1(n1408), .A2(n1259), .ZN(n1152) );
INV_X1 U1130 ( .A(G137), .ZN(n1259) );
XOR2_X1 U1131 ( .A(G131), .B(n1260), .Z(n1408) );
INV_X1 U1132 ( .A(G134), .ZN(n1260) );
NAND2_X1 U1133 ( .A1(n1407), .A2(KEYINPUT1), .ZN(n1405) );
XOR2_X1 U1134 ( .A(G134), .B(G131), .Z(n1407) );
endmodule


