//Key = 1111001011011111100000101011011101001111100010001100101001010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290;

XOR2_X1 U707 ( .A(n992), .B(n993), .Z(G9) );
XOR2_X1 U708 ( .A(KEYINPUT10), .B(G107), .Z(n993) );
NOR2_X1 U709 ( .A1(n994), .A2(n995), .ZN(G75) );
NOR4_X1 U710 ( .A1(G953), .A2(n996), .A3(n997), .A4(n998), .ZN(n995) );
NOR2_X1 U711 ( .A1(n999), .A2(n1000), .ZN(n997) );
NOR2_X1 U712 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NOR3_X1 U713 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1002) );
NOR2_X1 U714 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NOR2_X1 U715 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NOR3_X1 U716 ( .A1(n1010), .A2(n1011), .A3(n1012), .ZN(n1006) );
NOR3_X1 U717 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NOR2_X1 U718 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR2_X1 U719 ( .A1(n1018), .A2(n1019), .ZN(n1011) );
NOR4_X1 U720 ( .A1(n1013), .A2(n1020), .A3(n1010), .A4(n1009), .ZN(n1001) );
NOR2_X1 U721 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U722 ( .A1(n1023), .A2(n1003), .ZN(n1022) );
NOR2_X1 U723 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
XNOR2_X1 U724 ( .A(KEYINPUT41), .B(n1026), .ZN(n1025) );
NOR2_X1 U725 ( .A1(n1027), .A2(n1028), .ZN(n1024) );
NOR2_X1 U726 ( .A1(n1029), .A2(n1005), .ZN(n1021) );
NOR2_X1 U727 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR3_X1 U728 ( .A1(n996), .A2(G953), .A3(G952), .ZN(n994) );
AND4_X1 U729 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n996) );
NOR4_X1 U730 ( .A1(n1013), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1035) );
XNOR2_X1 U731 ( .A(n1039), .B(n1040), .ZN(n1038) );
XNOR2_X1 U732 ( .A(KEYINPUT4), .B(KEYINPUT0), .ZN(n1039) );
XOR2_X1 U733 ( .A(n1041), .B(n1042), .Z(n1037) );
NAND2_X1 U734 ( .A1(KEYINPUT31), .A2(n1043), .ZN(n1041) );
AND2_X1 U735 ( .A1(n1044), .A2(n1045), .ZN(n1036) );
NOR2_X1 U736 ( .A1(n1046), .A2(n1047), .ZN(n1034) );
XNOR2_X1 U737 ( .A(G469), .B(n1048), .ZN(n1047) );
XOR2_X1 U738 ( .A(KEYINPUT43), .B(n1049), .Z(n1046) );
NOR2_X1 U739 ( .A1(n1045), .A2(n1044), .ZN(n1049) );
NAND2_X1 U740 ( .A1(n1050), .A2(n1051), .ZN(G72) );
NAND2_X1 U741 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XNOR2_X1 U742 ( .A(n1054), .B(n1055), .ZN(n1052) );
NOR2_X1 U743 ( .A1(KEYINPUT20), .A2(n1056), .ZN(n1054) );
NAND2_X1 U744 ( .A1(n1057), .A2(G953), .ZN(n1050) );
XOR2_X1 U745 ( .A(n1055), .B(n1058), .Z(n1057) );
AND2_X1 U746 ( .A1(G227), .A2(G900), .ZN(n1058) );
NAND2_X1 U747 ( .A1(n1059), .A2(n1060), .ZN(n1055) );
NAND2_X1 U748 ( .A1(G953), .A2(n1061), .ZN(n1060) );
XOR2_X1 U749 ( .A(n1062), .B(n1063), .Z(n1059) );
XOR2_X1 U750 ( .A(n1064), .B(n1065), .Z(n1063) );
XOR2_X1 U751 ( .A(n1066), .B(KEYINPUT47), .Z(n1062) );
NAND2_X1 U752 ( .A1(n1067), .A2(n1068), .ZN(G69) );
NAND2_X1 U753 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XOR2_X1 U754 ( .A(KEYINPUT11), .B(n1071), .Z(n1067) );
NOR2_X1 U755 ( .A1(n1069), .A2(n1070), .ZN(n1071) );
NAND2_X1 U756 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NAND3_X1 U757 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
NAND2_X1 U758 ( .A1(G953), .A2(n1077), .ZN(n1074) );
XOR2_X1 U759 ( .A(KEYINPUT30), .B(n1078), .Z(n1072) );
NOR3_X1 U760 ( .A1(n1075), .A2(G953), .A3(n1076), .ZN(n1078) );
XNOR2_X1 U761 ( .A(n1079), .B(KEYINPUT51), .ZN(n1075) );
NAND2_X1 U762 ( .A1(G953), .A2(n1080), .ZN(n1069) );
NAND2_X1 U763 ( .A1(G898), .A2(G224), .ZN(n1080) );
NOR2_X1 U764 ( .A1(n1081), .A2(n1082), .ZN(G66) );
NOR3_X1 U765 ( .A1(n1045), .A2(n1083), .A3(n1084), .ZN(n1082) );
NOR3_X1 U766 ( .A1(n1085), .A2(n1044), .A3(n1086), .ZN(n1084) );
INV_X1 U767 ( .A(n1087), .ZN(n1086) );
NOR2_X1 U768 ( .A1(n1088), .A2(n1089), .ZN(n1083) );
NOR2_X1 U769 ( .A1(n1090), .A2(n1044), .ZN(n1088) );
NOR2_X1 U770 ( .A1(n1081), .A2(n1091), .ZN(G63) );
XOR2_X1 U771 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND2_X1 U772 ( .A1(n1087), .A2(G478), .ZN(n1092) );
NOR2_X1 U773 ( .A1(n1081), .A2(n1094), .ZN(G60) );
NOR3_X1 U774 ( .A1(n1042), .A2(n1095), .A3(n1096), .ZN(n1094) );
AND3_X1 U775 ( .A1(n1097), .A2(G475), .A3(n1087), .ZN(n1096) );
NOR2_X1 U776 ( .A1(n1098), .A2(n1097), .ZN(n1095) );
NOR2_X1 U777 ( .A1(n1090), .A2(n1043), .ZN(n1098) );
XNOR2_X1 U778 ( .A(G104), .B(n1099), .ZN(G6) );
NAND4_X1 U779 ( .A1(n1100), .A2(n1101), .A3(n1018), .A4(n1102), .ZN(n1099) );
NOR2_X1 U780 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U781 ( .A(KEYINPUT58), .B(n1105), .ZN(n1104) );
NOR2_X1 U782 ( .A1(n1081), .A2(n1106), .ZN(G57) );
XOR2_X1 U783 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND2_X1 U784 ( .A1(n1087), .A2(G472), .ZN(n1107) );
NOR3_X1 U785 ( .A1(n1109), .A2(n1081), .A3(n1110), .ZN(G54) );
NOR3_X1 U786 ( .A1(n1111), .A2(KEYINPUT32), .A3(n1112), .ZN(n1110) );
XOR2_X1 U787 ( .A(n1113), .B(n1114), .Z(n1111) );
NAND2_X1 U788 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U789 ( .A1(n1117), .A2(n1118), .ZN(n1109) );
XOR2_X1 U790 ( .A(n1113), .B(n1119), .Z(n1118) );
NAND2_X1 U791 ( .A1(n1120), .A2(n1116), .ZN(n1119) );
INV_X1 U792 ( .A(KEYINPUT46), .ZN(n1116) );
NAND2_X1 U793 ( .A1(n1087), .A2(G469), .ZN(n1113) );
NOR2_X1 U794 ( .A1(KEYINPUT32), .A2(n1112), .ZN(n1117) );
XOR2_X1 U795 ( .A(n1121), .B(n1122), .Z(n1112) );
XNOR2_X1 U796 ( .A(n1123), .B(n1065), .ZN(n1121) );
NOR2_X1 U797 ( .A1(n1081), .A2(n1124), .ZN(G51) );
XOR2_X1 U798 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U799 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND2_X1 U800 ( .A1(KEYINPUT36), .A2(n1129), .ZN(n1128) );
XOR2_X1 U801 ( .A(KEYINPUT9), .B(n1130), .Z(n1129) );
NAND2_X1 U802 ( .A1(n1087), .A2(n1131), .ZN(n1127) );
XOR2_X1 U803 ( .A(KEYINPUT17), .B(G210), .Z(n1131) );
NOR2_X1 U804 ( .A1(n1132), .A2(n1090), .ZN(n1087) );
INV_X1 U805 ( .A(n998), .ZN(n1090) );
NAND2_X1 U806 ( .A1(n1076), .A2(n1056), .ZN(n998) );
AND2_X1 U807 ( .A1(n1133), .A2(n1134), .ZN(n1056) );
NOR4_X1 U808 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1134) );
NOR4_X1 U809 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1133) );
NOR3_X1 U810 ( .A1(n1143), .A2(n1026), .A3(n1103), .ZN(n1142) );
NOR3_X1 U811 ( .A1(n1144), .A2(n1008), .A3(n1005), .ZN(n1141) );
INV_X1 U812 ( .A(n1145), .ZN(n1140) );
AND2_X1 U813 ( .A1(n1146), .A2(n1147), .ZN(n1076) );
NOR4_X1 U814 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1147) );
NOR4_X1 U815 ( .A1(n1152), .A2(n992), .A3(n1153), .A4(n1154), .ZN(n1146) );
NOR3_X1 U816 ( .A1(n1103), .A2(n1009), .A3(n1155), .ZN(n1154) );
NOR3_X1 U817 ( .A1(n1155), .A2(n1009), .A3(n1156), .ZN(n992) );
NOR2_X1 U818 ( .A1(n1026), .A2(n1157), .ZN(n1152) );
NOR2_X1 U819 ( .A1(n1158), .A2(G952), .ZN(n1081) );
XNOR2_X1 U820 ( .A(KEYINPUT21), .B(G953), .ZN(n1158) );
XNOR2_X1 U821 ( .A(G146), .B(n1159), .ZN(G48) );
NAND2_X1 U822 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U823 ( .A(KEYINPUT56), .B(n1162), .Z(n1161) );
NOR2_X1 U824 ( .A1(n1103), .A2(n1143), .ZN(n1162) );
INV_X1 U825 ( .A(n1031), .ZN(n1103) );
NAND2_X1 U826 ( .A1(n1163), .A2(n1164), .ZN(G45) );
NAND2_X1 U827 ( .A1(n1165), .A2(n1145), .ZN(n1164) );
XOR2_X1 U828 ( .A(KEYINPUT26), .B(n1166), .Z(n1163) );
NOR2_X1 U829 ( .A1(n1145), .A2(n1165), .ZN(n1166) );
XNOR2_X1 U830 ( .A(KEYINPUT61), .B(n1167), .ZN(n1165) );
NAND4_X1 U831 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1145) );
NOR3_X1 U832 ( .A1(n1172), .A2(n1026), .A3(n1008), .ZN(n1171) );
XNOR2_X1 U833 ( .A(G140), .B(n1173), .ZN(G42) );
NAND3_X1 U834 ( .A1(n1101), .A2(n1174), .A3(n1175), .ZN(n1173) );
INV_X1 U835 ( .A(n1144), .ZN(n1175) );
XNOR2_X1 U836 ( .A(KEYINPUT53), .B(n1005), .ZN(n1174) );
XNOR2_X1 U837 ( .A(n1176), .B(n1139), .ZN(G39) );
NOR3_X1 U838 ( .A1(n1003), .A2(n1005), .A3(n1143), .ZN(n1139) );
XOR2_X1 U839 ( .A(G134), .B(n1138), .Z(G36) );
AND3_X1 U840 ( .A1(n1030), .A2(n1169), .A3(n1177), .ZN(n1138) );
XOR2_X1 U841 ( .A(n1137), .B(n1178), .Z(G33) );
XOR2_X1 U842 ( .A(KEYINPUT23), .B(G131), .Z(n1178) );
AND3_X1 U843 ( .A1(n1031), .A2(n1169), .A3(n1177), .ZN(n1137) );
NOR3_X1 U844 ( .A1(n1005), .A2(n1008), .A3(n1172), .ZN(n1177) );
INV_X1 U845 ( .A(n1033), .ZN(n1005) );
NOR2_X1 U846 ( .A1(n1027), .A2(n1179), .ZN(n1033) );
INV_X1 U847 ( .A(n1028), .ZN(n1179) );
XNOR2_X1 U848 ( .A(G128), .B(n1180), .ZN(G30) );
NAND2_X1 U849 ( .A1(KEYINPUT48), .A2(n1136), .ZN(n1180) );
NOR3_X1 U850 ( .A1(n1156), .A2(n1026), .A3(n1143), .ZN(n1136) );
NAND4_X1 U851 ( .A1(n1181), .A2(n1101), .A3(n1017), .A4(n1169), .ZN(n1143) );
INV_X1 U852 ( .A(n1030), .ZN(n1156) );
XOR2_X1 U853 ( .A(n1151), .B(n1182), .Z(G3) );
NOR2_X1 U854 ( .A1(KEYINPUT19), .A2(n1183), .ZN(n1182) );
INV_X1 U855 ( .A(G101), .ZN(n1183) );
NOR3_X1 U856 ( .A1(n1172), .A2(n1155), .A3(n1003), .ZN(n1151) );
XNOR2_X1 U857 ( .A(n1135), .B(n1184), .ZN(G27) );
NOR2_X1 U858 ( .A1(G125), .A2(KEYINPUT42), .ZN(n1184) );
NOR4_X1 U859 ( .A1(n1144), .A2(n1026), .A3(n1010), .A4(n1013), .ZN(n1135) );
NAND4_X1 U860 ( .A1(n1040), .A2(n1031), .A3(n1181), .A4(n1169), .ZN(n1144) );
NAND2_X1 U861 ( .A1(n1185), .A2(n1186), .ZN(n1169) );
NAND4_X1 U862 ( .A1(G953), .A2(G902), .A3(n1187), .A4(n1061), .ZN(n1186) );
INV_X1 U863 ( .A(G900), .ZN(n1061) );
XNOR2_X1 U864 ( .A(KEYINPUT6), .B(n1000), .ZN(n1185) );
XNOR2_X1 U865 ( .A(n1150), .B(n1188), .ZN(G24) );
XNOR2_X1 U866 ( .A(KEYINPUT33), .B(n1189), .ZN(n1188) );
AND3_X1 U867 ( .A1(n1190), .A2(n1018), .A3(n1191), .ZN(n1150) );
NOR3_X1 U868 ( .A1(n1026), .A2(n1032), .A3(n1192), .ZN(n1191) );
INV_X1 U869 ( .A(n1009), .ZN(n1018) );
NAND2_X1 U870 ( .A1(n1193), .A2(n1040), .ZN(n1009) );
XOR2_X1 U871 ( .A(G119), .B(n1149), .Z(G21) );
AND4_X1 U872 ( .A1(n1194), .A2(n1190), .A3(n1195), .A4(n1181), .ZN(n1149) );
INV_X1 U873 ( .A(n1016), .ZN(n1181) );
NOR2_X1 U874 ( .A1(n1040), .A2(n1026), .ZN(n1195) );
INV_X1 U875 ( .A(n1017), .ZN(n1040) );
XNOR2_X1 U876 ( .A(G116), .B(n1196), .ZN(G18) );
NAND3_X1 U877 ( .A1(n1160), .A2(n1197), .A3(KEYINPUT8), .ZN(n1196) );
XNOR2_X1 U878 ( .A(KEYINPUT50), .B(n1157), .ZN(n1197) );
NAND3_X1 U879 ( .A1(n1014), .A2(n1030), .A3(n1190), .ZN(n1157) );
NOR2_X1 U880 ( .A1(n1170), .A2(n1032), .ZN(n1030) );
INV_X1 U881 ( .A(n1168), .ZN(n1032) );
NAND2_X1 U882 ( .A1(n1198), .A2(n1199), .ZN(G15) );
NAND2_X1 U883 ( .A1(n1148), .A2(n1200), .ZN(n1199) );
XOR2_X1 U884 ( .A(KEYINPUT52), .B(n1201), .Z(n1198) );
NOR2_X1 U885 ( .A1(n1148), .A2(n1200), .ZN(n1201) );
AND4_X1 U886 ( .A1(n1190), .A2(n1031), .A3(n1100), .A4(n1014), .ZN(n1148) );
INV_X1 U887 ( .A(n1172), .ZN(n1014) );
NAND2_X1 U888 ( .A1(n1193), .A2(n1017), .ZN(n1172) );
XNOR2_X1 U889 ( .A(n1016), .B(KEYINPUT57), .ZN(n1193) );
NOR2_X1 U890 ( .A1(n1168), .A2(n1192), .ZN(n1031) );
NOR3_X1 U891 ( .A1(n1013), .A2(n1202), .A3(n1010), .ZN(n1190) );
INV_X1 U892 ( .A(n1105), .ZN(n1202) );
INV_X1 U893 ( .A(n1019), .ZN(n1013) );
XOR2_X1 U894 ( .A(n1153), .B(n1203), .Z(G12) );
XOR2_X1 U895 ( .A(KEYINPUT35), .B(G110), .Z(n1203) );
NOR4_X1 U896 ( .A1(n1003), .A2(n1155), .A3(n1016), .A4(n1017), .ZN(n1153) );
XNOR2_X1 U897 ( .A(n1204), .B(G472), .ZN(n1017) );
NAND2_X1 U898 ( .A1(n1205), .A2(n1132), .ZN(n1204) );
XOR2_X1 U899 ( .A(n1108), .B(KEYINPUT25), .Z(n1205) );
XOR2_X1 U900 ( .A(n1206), .B(n1207), .Z(n1108) );
XOR2_X1 U901 ( .A(n1208), .B(n1209), .Z(n1207) );
XNOR2_X1 U902 ( .A(G119), .B(n1210), .ZN(n1209) );
NAND2_X1 U903 ( .A1(G210), .A2(n1211), .ZN(n1210) );
NOR2_X1 U904 ( .A1(G116), .A2(KEYINPUT28), .ZN(n1208) );
XOR2_X1 U905 ( .A(n1212), .B(n1130), .Z(n1206) );
XOR2_X1 U906 ( .A(n1123), .B(n1213), .Z(n1212) );
XNOR2_X1 U907 ( .A(n1044), .B(n1214), .ZN(n1016) );
NOR2_X1 U908 ( .A1(KEYINPUT18), .A2(n1215), .ZN(n1214) );
XNOR2_X1 U909 ( .A(n1045), .B(KEYINPUT44), .ZN(n1215) );
NOR2_X1 U910 ( .A1(n1089), .A2(G902), .ZN(n1045) );
INV_X1 U911 ( .A(n1085), .ZN(n1089) );
XNOR2_X1 U912 ( .A(n1216), .B(n1217), .ZN(n1085) );
XOR2_X1 U913 ( .A(G110), .B(n1218), .Z(n1217) );
XNOR2_X1 U914 ( .A(n1219), .B(G119), .ZN(n1218) );
INV_X1 U915 ( .A(G128), .ZN(n1219) );
XOR2_X1 U916 ( .A(n1220), .B(n1221), .Z(n1216) );
NOR2_X1 U917 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NOR2_X1 U918 ( .A1(n1224), .A2(G137), .ZN(n1223) );
NOR3_X1 U919 ( .A1(n1225), .A2(G953), .A3(n1226), .ZN(n1224) );
NOR4_X1 U920 ( .A1(G953), .A2(n1227), .A3(n1226), .A4(n1225), .ZN(n1222) );
INV_X1 U921 ( .A(G221), .ZN(n1225) );
INV_X1 U922 ( .A(G234), .ZN(n1226) );
XNOR2_X1 U923 ( .A(G137), .B(KEYINPUT5), .ZN(n1227) );
NAND2_X1 U924 ( .A1(KEYINPUT22), .A2(n1228), .ZN(n1220) );
XOR2_X1 U925 ( .A(G146), .B(n1229), .Z(n1228) );
NOR2_X1 U926 ( .A1(KEYINPUT55), .A2(n1064), .ZN(n1229) );
NAND2_X1 U927 ( .A1(G217), .A2(n1230), .ZN(n1044) );
NAND3_X1 U928 ( .A1(n1100), .A2(n1105), .A3(n1101), .ZN(n1155) );
INV_X1 U929 ( .A(n1008), .ZN(n1101) );
NAND2_X1 U930 ( .A1(n1010), .A2(n1019), .ZN(n1008) );
NAND2_X1 U931 ( .A1(G221), .A2(n1230), .ZN(n1019) );
NAND2_X1 U932 ( .A1(G234), .A2(n1132), .ZN(n1230) );
XNOR2_X1 U933 ( .A(n1231), .B(n1048), .ZN(n1010) );
NAND2_X1 U934 ( .A1(n1232), .A2(n1132), .ZN(n1048) );
XOR2_X1 U935 ( .A(n1233), .B(n1234), .Z(n1232) );
XNOR2_X1 U936 ( .A(n1123), .B(n1120), .ZN(n1234) );
INV_X1 U937 ( .A(n1115), .ZN(n1120) );
XNOR2_X1 U938 ( .A(n1235), .B(n1236), .ZN(n1115) );
XOR2_X1 U939 ( .A(G140), .B(G110), .Z(n1236) );
NAND2_X1 U940 ( .A1(G227), .A2(n1053), .ZN(n1235) );
XOR2_X1 U941 ( .A(n1066), .B(KEYINPUT45), .Z(n1123) );
XOR2_X1 U942 ( .A(n1237), .B(n1238), .Z(n1066) );
XNOR2_X1 U943 ( .A(KEYINPUT14), .B(n1176), .ZN(n1238) );
INV_X1 U944 ( .A(G137), .ZN(n1176) );
XNOR2_X1 U945 ( .A(G134), .B(n1239), .ZN(n1237) );
XOR2_X1 U946 ( .A(n1240), .B(KEYINPUT7), .Z(n1233) );
NAND2_X1 U947 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
NAND2_X1 U948 ( .A1(n1122), .A2(n1065), .ZN(n1242) );
XOR2_X1 U949 ( .A(KEYINPUT24), .B(n1243), .Z(n1241) );
NOR2_X1 U950 ( .A1(n1122), .A2(n1065), .ZN(n1243) );
XNOR2_X1 U951 ( .A(G128), .B(n1244), .ZN(n1065) );
XOR2_X1 U952 ( .A(n1245), .B(n1246), .Z(n1122) );
XNOR2_X1 U953 ( .A(G101), .B(KEYINPUT62), .ZN(n1245) );
NAND2_X1 U954 ( .A1(KEYINPUT40), .A2(n1247), .ZN(n1231) );
INV_X1 U955 ( .A(G469), .ZN(n1247) );
NAND2_X1 U956 ( .A1(n1000), .A2(n1248), .ZN(n1105) );
NAND4_X1 U957 ( .A1(G953), .A2(G902), .A3(n1187), .A4(n1077), .ZN(n1248) );
INV_X1 U958 ( .A(G898), .ZN(n1077) );
NAND3_X1 U959 ( .A1(n1187), .A2(n1053), .A3(G952), .ZN(n1000) );
NAND2_X1 U960 ( .A1(G237), .A2(G234), .ZN(n1187) );
XNOR2_X1 U961 ( .A(n1160), .B(KEYINPUT63), .ZN(n1100) );
INV_X1 U962 ( .A(n1026), .ZN(n1160) );
NAND2_X1 U963 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U964 ( .A1(G214), .A2(n1249), .ZN(n1028) );
XOR2_X1 U965 ( .A(KEYINPUT2), .B(n1250), .Z(n1249) );
NOR2_X1 U966 ( .A1(G237), .A2(G902), .ZN(n1250) );
NAND3_X1 U967 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1027) );
NAND2_X1 U968 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
OR3_X1 U969 ( .A1(n1255), .A2(n1254), .A3(G902), .ZN(n1252) );
AND2_X1 U970 ( .A1(G210), .A2(G237), .ZN(n1254) );
XNOR2_X1 U971 ( .A(n1256), .B(n1257), .ZN(n1255) );
XOR2_X1 U972 ( .A(KEYINPUT49), .B(KEYINPUT27), .Z(n1257) );
XOR2_X1 U973 ( .A(n1125), .B(n1130), .Z(n1256) );
XNOR2_X1 U974 ( .A(n1258), .B(n1259), .ZN(n1130) );
XNOR2_X1 U975 ( .A(n1167), .B(G128), .ZN(n1259) );
NAND2_X1 U976 ( .A1(KEYINPUT59), .A2(G146), .ZN(n1258) );
XOR2_X1 U977 ( .A(n1260), .B(n1261), .Z(n1125) );
XNOR2_X1 U978 ( .A(G125), .B(n1262), .ZN(n1261) );
XNOR2_X1 U979 ( .A(KEYINPUT3), .B(KEYINPUT29), .ZN(n1262) );
XOR2_X1 U980 ( .A(n1079), .B(n1263), .Z(n1260) );
AND2_X1 U981 ( .A1(n1053), .A2(G224), .ZN(n1263) );
XOR2_X1 U982 ( .A(n1264), .B(n1265), .Z(n1079) );
XNOR2_X1 U983 ( .A(n1213), .B(n1266), .ZN(n1265) );
XNOR2_X1 U984 ( .A(n1267), .B(n1268), .ZN(n1266) );
NAND2_X1 U985 ( .A1(KEYINPUT38), .A2(n1189), .ZN(n1268) );
NAND2_X1 U986 ( .A1(KEYINPUT54), .A2(G119), .ZN(n1267) );
XNOR2_X1 U987 ( .A(G101), .B(n1200), .ZN(n1213) );
XOR2_X1 U988 ( .A(n1269), .B(n1270), .Z(n1264) );
XOR2_X1 U989 ( .A(KEYINPUT37), .B(G116), .Z(n1270) );
XOR2_X1 U990 ( .A(n1271), .B(G110), .Z(n1269) );
NAND2_X1 U991 ( .A1(n1272), .A2(KEYINPUT12), .ZN(n1271) );
XNOR2_X1 U992 ( .A(n1246), .B(KEYINPUT15), .ZN(n1272) );
XNOR2_X1 U993 ( .A(n1273), .B(n1274), .ZN(n1246) );
XNOR2_X1 U994 ( .A(G107), .B(KEYINPUT16), .ZN(n1273) );
NAND2_X1 U995 ( .A1(G210), .A2(G902), .ZN(n1251) );
INV_X1 U996 ( .A(n1194), .ZN(n1003) );
NOR2_X1 U997 ( .A1(n1168), .A2(n1170), .ZN(n1194) );
INV_X1 U998 ( .A(n1192), .ZN(n1170) );
XOR2_X1 U999 ( .A(n1042), .B(n1043), .Z(n1192) );
INV_X1 U1000 ( .A(G475), .ZN(n1043) );
NOR2_X1 U1001 ( .A1(n1097), .A2(G902), .ZN(n1042) );
XOR2_X1 U1002 ( .A(n1275), .B(n1276), .Z(n1097) );
XOR2_X1 U1003 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U1004 ( .A(n1274), .B(n1244), .Z(n1278) );
XNOR2_X1 U1005 ( .A(n1167), .B(G146), .ZN(n1244) );
INV_X1 U1006 ( .A(G143), .ZN(n1167) );
XOR2_X1 U1007 ( .A(G104), .B(KEYINPUT60), .Z(n1274) );
XNOR2_X1 U1008 ( .A(n1239), .B(n1064), .ZN(n1277) );
XNOR2_X1 U1009 ( .A(G125), .B(G140), .ZN(n1064) );
XOR2_X1 U1010 ( .A(G131), .B(KEYINPUT13), .Z(n1239) );
XOR2_X1 U1011 ( .A(n1279), .B(n1280), .Z(n1275) );
XNOR2_X1 U1012 ( .A(KEYINPUT39), .B(n1189), .ZN(n1280) );
XNOR2_X1 U1013 ( .A(n1281), .B(n1200), .ZN(n1279) );
INV_X1 U1014 ( .A(G113), .ZN(n1200) );
NAND2_X1 U1015 ( .A1(G214), .A2(n1211), .ZN(n1281) );
NOR2_X1 U1016 ( .A1(G953), .A2(G237), .ZN(n1211) );
XNOR2_X1 U1017 ( .A(n1282), .B(G478), .ZN(n1168) );
NAND2_X1 U1018 ( .A1(n1093), .A2(n1132), .ZN(n1282) );
INV_X1 U1019 ( .A(G902), .ZN(n1132) );
XNOR2_X1 U1020 ( .A(n1283), .B(n1284), .ZN(n1093) );
XOR2_X1 U1021 ( .A(n1285), .B(n1286), .Z(n1284) );
NAND3_X1 U1022 ( .A1(G217), .A2(n1053), .A3(G234), .ZN(n1286) );
INV_X1 U1023 ( .A(G953), .ZN(n1053) );
NAND2_X1 U1024 ( .A1(n1287), .A2(KEYINPUT1), .ZN(n1285) );
XNOR2_X1 U1025 ( .A(G107), .B(n1288), .ZN(n1287) );
XNOR2_X1 U1026 ( .A(n1189), .B(G116), .ZN(n1288) );
INV_X1 U1027 ( .A(G122), .ZN(n1189) );
XOR2_X1 U1028 ( .A(n1289), .B(n1290), .Z(n1283) );
NOR2_X1 U1029 ( .A1(KEYINPUT34), .A2(G128), .ZN(n1290) );
XNOR2_X1 U1030 ( .A(G134), .B(G143), .ZN(n1289) );
endmodule


