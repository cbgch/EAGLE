//Key = 0010101111101100011011100000100010101010100110010010010101100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300;

XOR2_X1 U716 ( .A(G107), .B(n994), .Z(G9) );
NOR2_X1 U717 ( .A1(n995), .A2(n996), .ZN(G75) );
NOR4_X1 U718 ( .A1(n997), .A2(n998), .A3(G953), .A4(n999), .ZN(n996) );
NOR2_X1 U719 ( .A1(n1000), .A2(n1001), .ZN(n998) );
NOR2_X1 U720 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NOR2_X1 U721 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NOR2_X1 U722 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NOR2_X1 U723 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NOR2_X1 U724 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NOR2_X1 U725 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR2_X1 U726 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
XOR2_X1 U727 ( .A(KEYINPUT41), .B(n1016), .Z(n1015) );
NOR2_X1 U728 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
XNOR2_X1 U729 ( .A(n1019), .B(KEYINPUT53), .ZN(n1014) );
NOR2_X1 U730 ( .A1(n1020), .A2(n1021), .ZN(n1010) );
NOR2_X1 U731 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U732 ( .A1(n1024), .A2(n1025), .ZN(n1006) );
XNOR2_X1 U733 ( .A(n1026), .B(n1027), .ZN(n1025) );
NOR3_X1 U734 ( .A1(n1009), .A2(n1028), .A3(n1024), .ZN(n1002) );
INV_X1 U735 ( .A(n1029), .ZN(n1024) );
NOR2_X1 U736 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NAND3_X1 U737 ( .A1(n1032), .A2(n1033), .A3(KEYINPUT32), .ZN(n997) );
NOR3_X1 U738 ( .A1(n999), .A2(G953), .A3(G952), .ZN(n995) );
AND3_X1 U739 ( .A1(n1034), .A2(n1029), .A3(n1035), .ZN(n999) );
NOR3_X1 U740 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
XOR2_X1 U741 ( .A(n1039), .B(n1040), .Z(n1038) );
NAND2_X1 U742 ( .A1(KEYINPUT43), .A2(n1041), .ZN(n1039) );
NOR2_X1 U743 ( .A1(n1021), .A2(n1013), .ZN(n1029) );
XNOR2_X1 U744 ( .A(n1042), .B(n1043), .ZN(n1034) );
XOR2_X1 U745 ( .A(n1044), .B(n1045), .Z(G72) );
XOR2_X1 U746 ( .A(n1046), .B(n1047), .Z(n1045) );
NAND2_X1 U747 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U748 ( .A1(G953), .A2(n1050), .ZN(n1049) );
XOR2_X1 U749 ( .A(n1051), .B(n1052), .Z(n1048) );
XNOR2_X1 U750 ( .A(G125), .B(n1053), .ZN(n1052) );
XNOR2_X1 U751 ( .A(KEYINPUT59), .B(KEYINPUT5), .ZN(n1053) );
XOR2_X1 U752 ( .A(n1054), .B(n1055), .Z(n1051) );
XOR2_X1 U753 ( .A(n1056), .B(n1057), .Z(n1055) );
NOR2_X1 U754 ( .A1(G140), .A2(KEYINPUT30), .ZN(n1056) );
NAND2_X1 U755 ( .A1(n1058), .A2(n1059), .ZN(n1046) );
NAND2_X1 U756 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
XNOR2_X1 U757 ( .A(KEYINPUT58), .B(n1062), .ZN(n1058) );
NOR2_X1 U758 ( .A1(n1063), .A2(n1062), .ZN(n1044) );
AND2_X1 U759 ( .A1(G227), .A2(G900), .ZN(n1063) );
NAND2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(G69) );
NAND2_X1 U761 ( .A1(G953), .A2(n1066), .ZN(n1065) );
XOR2_X1 U762 ( .A(n1067), .B(n1068), .Z(n1064) );
NOR2_X1 U763 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NOR2_X1 U764 ( .A1(G953), .A2(n1032), .ZN(n1070) );
NOR2_X1 U765 ( .A1(G224), .A2(n1062), .ZN(n1069) );
NOR2_X1 U766 ( .A1(KEYINPUT51), .A2(n1071), .ZN(n1067) );
XOR2_X1 U767 ( .A(n1072), .B(n1073), .Z(n1071) );
XOR2_X1 U768 ( .A(KEYINPUT48), .B(n1074), .Z(n1073) );
NOR2_X1 U769 ( .A1(KEYINPUT61), .A2(n1075), .ZN(n1074) );
NOR2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(G66) );
XOR2_X1 U771 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U772 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR2_X1 U773 ( .A1(n1076), .A2(n1082), .ZN(G63) );
NOR3_X1 U774 ( .A1(n1040), .A2(n1083), .A3(n1084), .ZN(n1082) );
AND3_X1 U775 ( .A1(n1085), .A2(G478), .A3(n1086), .ZN(n1084) );
NOR2_X1 U776 ( .A1(n1087), .A2(n1085), .ZN(n1083) );
NOR2_X1 U777 ( .A1(n1088), .A2(n1041), .ZN(n1087) );
INV_X1 U778 ( .A(G478), .ZN(n1041) );
NOR2_X1 U779 ( .A1(n1076), .A2(n1089), .ZN(G60) );
XNOR2_X1 U780 ( .A(n1090), .B(n1091), .ZN(n1089) );
AND2_X1 U781 ( .A1(G475), .A2(n1086), .ZN(n1091) );
XNOR2_X1 U782 ( .A(G104), .B(n1092), .ZN(G6) );
NOR2_X1 U783 ( .A1(KEYINPUT1), .A2(n1093), .ZN(n1092) );
NOR3_X1 U784 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
XNOR2_X1 U785 ( .A(n1097), .B(KEYINPUT16), .ZN(n1095) );
NOR2_X1 U786 ( .A1(n1076), .A2(n1098), .ZN(G57) );
XOR2_X1 U787 ( .A(n1099), .B(n1100), .Z(n1098) );
XOR2_X1 U788 ( .A(n1101), .B(n1102), .Z(n1100) );
AND2_X1 U789 ( .A1(G472), .A2(n1086), .ZN(n1102) );
XNOR2_X1 U790 ( .A(n1103), .B(KEYINPUT2), .ZN(n1099) );
NOR2_X1 U791 ( .A1(n1076), .A2(n1104), .ZN(G54) );
XOR2_X1 U792 ( .A(n1105), .B(n1106), .Z(n1104) );
XOR2_X1 U793 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U794 ( .A1(n1043), .A2(n1081), .ZN(n1108) );
INV_X1 U795 ( .A(n1086), .ZN(n1081) );
NOR2_X1 U796 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
XOR2_X1 U797 ( .A(n1111), .B(n1112), .Z(n1105) );
NOR2_X1 U798 ( .A1(KEYINPUT35), .A2(n1113), .ZN(n1112) );
NOR2_X1 U799 ( .A1(n1076), .A2(n1114), .ZN(G51) );
XNOR2_X1 U800 ( .A(n1115), .B(n1116), .ZN(n1114) );
XOR2_X1 U801 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U802 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XOR2_X1 U803 ( .A(n1121), .B(KEYINPUT22), .Z(n1120) );
NAND2_X1 U804 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U805 ( .A1(n1122), .A2(n1124), .ZN(n1119) );
XNOR2_X1 U806 ( .A(KEYINPUT63), .B(n1123), .ZN(n1124) );
XOR2_X1 U807 ( .A(n1125), .B(KEYINPUT14), .Z(n1123) );
XNOR2_X1 U808 ( .A(n1126), .B(n1127), .ZN(n1122) );
NAND2_X1 U809 ( .A1(KEYINPUT50), .A2(n1128), .ZN(n1126) );
NAND3_X1 U810 ( .A1(n1086), .A2(n1129), .A3(KEYINPUT57), .ZN(n1117) );
NOR2_X1 U811 ( .A1(n1130), .A2(n1088), .ZN(n1086) );
AND2_X1 U812 ( .A1(n1131), .A2(n1033), .ZN(n1088) );
AND2_X1 U813 ( .A1(n1132), .A2(n1060), .ZN(n1033) );
AND4_X1 U814 ( .A1(n1133), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n1060) );
AND4_X1 U815 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1136) );
NAND2_X1 U816 ( .A1(n1141), .A2(n1142), .ZN(n1135) );
INV_X1 U817 ( .A(n1143), .ZN(n1142) );
XNOR2_X1 U818 ( .A(n1144), .B(KEYINPUT36), .ZN(n1141) );
NAND3_X1 U819 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(n1133) );
XNOR2_X1 U820 ( .A(n1144), .B(KEYINPUT9), .ZN(n1147) );
XOR2_X1 U821 ( .A(n1061), .B(KEYINPUT25), .Z(n1132) );
XNOR2_X1 U822 ( .A(n1032), .B(KEYINPUT10), .ZN(n1131) );
AND2_X1 U823 ( .A1(n1148), .A2(n1149), .ZN(n1032) );
NOR4_X1 U824 ( .A1(n1150), .A2(n1151), .A3(n994), .A4(n1152), .ZN(n1149) );
INV_X1 U825 ( .A(n1153), .ZN(n1152) );
AND3_X1 U826 ( .A1(n1154), .A2(n1030), .A3(n1097), .ZN(n994) );
NOR4_X1 U827 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1148) );
NOR2_X1 U828 ( .A1(n1159), .A2(n1096), .ZN(n1158) );
INV_X1 U829 ( .A(n1154), .ZN(n1096) );
NOR2_X1 U830 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR2_X1 U831 ( .A1(n1013), .A2(n1094), .ZN(n1161) );
INV_X1 U832 ( .A(n1097), .ZN(n1013) );
NOR2_X1 U833 ( .A1(n1162), .A2(n1163), .ZN(n1160) );
XNOR2_X1 U834 ( .A(KEYINPUT55), .B(n1005), .ZN(n1163) );
INV_X1 U835 ( .A(n1164), .ZN(n1157) );
NOR2_X1 U836 ( .A1(n1165), .A2(n1166), .ZN(n1156) );
INV_X1 U837 ( .A(KEYINPUT21), .ZN(n1165) );
NOR3_X1 U838 ( .A1(KEYINPUT21), .A2(n1167), .A3(n1168), .ZN(n1155) );
NOR2_X1 U839 ( .A1(n1062), .A2(G952), .ZN(n1076) );
XNOR2_X1 U840 ( .A(G146), .B(n1134), .ZN(G48) );
NAND2_X1 U841 ( .A1(n1145), .A2(n1169), .ZN(n1134) );
XNOR2_X1 U842 ( .A(G143), .B(n1140), .ZN(G45) );
NAND3_X1 U843 ( .A1(n1170), .A2(n1023), .A3(n1171), .ZN(n1140) );
XNOR2_X1 U844 ( .A(G140), .B(n1061), .ZN(G42) );
NAND4_X1 U845 ( .A1(n1171), .A2(n1031), .A3(n1022), .A4(n1144), .ZN(n1061) );
XOR2_X1 U846 ( .A(G137), .B(n1172), .Z(G39) );
NOR3_X1 U847 ( .A1(n1173), .A2(n1021), .A3(n1005), .ZN(n1172) );
XOR2_X1 U848 ( .A(G134), .B(n1174), .Z(G36) );
NOR2_X1 U849 ( .A1(n1021), .A2(n1143), .ZN(n1174) );
NAND3_X1 U850 ( .A1(n1023), .A2(n1030), .A3(n1171), .ZN(n1143) );
XNOR2_X1 U851 ( .A(G131), .B(n1137), .ZN(G33) );
NAND4_X1 U852 ( .A1(n1171), .A2(n1031), .A3(n1023), .A4(n1144), .ZN(n1137) );
INV_X1 U853 ( .A(n1021), .ZN(n1144) );
NAND2_X1 U854 ( .A1(n1175), .A2(n1018), .ZN(n1021) );
INV_X1 U855 ( .A(n1017), .ZN(n1175) );
INV_X1 U856 ( .A(n1094), .ZN(n1031) );
XNOR2_X1 U857 ( .A(G128), .B(n1139), .ZN(G30) );
NAND3_X1 U858 ( .A1(n1030), .A2(n1019), .A3(n1145), .ZN(n1139) );
INV_X1 U859 ( .A(n1173), .ZN(n1145) );
NAND3_X1 U860 ( .A1(n1176), .A2(n1177), .A3(n1171), .ZN(n1173) );
AND3_X1 U861 ( .A1(n1178), .A2(n1026), .A3(n1179), .ZN(n1171) );
XNOR2_X1 U862 ( .A(G101), .B(n1180), .ZN(G3) );
NAND4_X1 U863 ( .A1(KEYINPUT38), .A2(n1023), .A3(n1146), .A4(n1154), .ZN(n1180) );
NAND2_X1 U864 ( .A1(n1181), .A2(n1182), .ZN(G27) );
NAND2_X1 U865 ( .A1(n1183), .A2(n1138), .ZN(n1182) );
XOR2_X1 U866 ( .A(KEYINPUT20), .B(n1184), .Z(n1181) );
NOR2_X1 U867 ( .A1(n1138), .A2(n1183), .ZN(n1184) );
XNOR2_X1 U868 ( .A(KEYINPUT27), .B(n1127), .ZN(n1183) );
NAND4_X1 U869 ( .A1(n1169), .A2(n1185), .A3(n1022), .A4(n1178), .ZN(n1138) );
NAND2_X1 U870 ( .A1(n1001), .A2(n1186), .ZN(n1178) );
NAND4_X1 U871 ( .A1(G953), .A2(G902), .A3(n1187), .A4(n1050), .ZN(n1186) );
INV_X1 U872 ( .A(G900), .ZN(n1050) );
XNOR2_X1 U873 ( .A(G122), .B(n1164), .ZN(G24) );
NAND4_X1 U874 ( .A1(n1170), .A2(n1185), .A3(n1097), .A4(n1188), .ZN(n1164) );
NOR2_X1 U875 ( .A1(n1189), .A2(n1177), .ZN(n1097) );
NOR3_X1 U876 ( .A1(n1190), .A2(n1191), .A3(n1168), .ZN(n1170) );
XNOR2_X1 U877 ( .A(n1151), .B(n1192), .ZN(G21) );
NOR2_X1 U878 ( .A1(G119), .A2(KEYINPUT31), .ZN(n1192) );
AND4_X1 U879 ( .A1(n1176), .A2(n1146), .A3(n1185), .A4(n1193), .ZN(n1151) );
NOR3_X1 U880 ( .A1(n1168), .A2(n1194), .A3(n1195), .ZN(n1193) );
NAND2_X1 U881 ( .A1(n1196), .A2(n1197), .ZN(G18) );
NAND2_X1 U882 ( .A1(KEYINPUT49), .A2(n1198), .ZN(n1197) );
XOR2_X1 U883 ( .A(n1166), .B(n1199), .Z(n1196) );
NOR2_X1 U884 ( .A1(KEYINPUT49), .A2(n1198), .ZN(n1199) );
NAND2_X1 U885 ( .A1(n1167), .A2(n1019), .ZN(n1166) );
INV_X1 U886 ( .A(n1168), .ZN(n1019) );
AND2_X1 U887 ( .A1(n1200), .A2(n1030), .ZN(n1167) );
NOR2_X1 U888 ( .A1(n1036), .A2(n1190), .ZN(n1030) );
XOR2_X1 U889 ( .A(G113), .B(n1201), .Z(G15) );
NOR2_X1 U890 ( .A1(KEYINPUT3), .A2(n1153), .ZN(n1201) );
NAND2_X1 U891 ( .A1(n1200), .A2(n1169), .ZN(n1153) );
NOR2_X1 U892 ( .A1(n1094), .A2(n1168), .ZN(n1169) );
NAND2_X1 U893 ( .A1(n1190), .A2(n1036), .ZN(n1094) );
NOR3_X1 U894 ( .A1(n1009), .A2(n1194), .A3(n1162), .ZN(n1200) );
INV_X1 U895 ( .A(n1023), .ZN(n1162) );
NOR2_X1 U896 ( .A1(n1189), .A2(n1195), .ZN(n1023) );
INV_X1 U897 ( .A(n1185), .ZN(n1009) );
NOR2_X1 U898 ( .A1(n1179), .A2(n1037), .ZN(n1185) );
INV_X1 U899 ( .A(n1027), .ZN(n1179) );
XNOR2_X1 U900 ( .A(n1202), .B(n1150), .ZN(G12) );
AND3_X1 U901 ( .A1(n1022), .A2(n1154), .A3(n1146), .ZN(n1150) );
INV_X1 U902 ( .A(n1005), .ZN(n1146) );
NAND2_X1 U903 ( .A1(n1190), .A2(n1191), .ZN(n1005) );
INV_X1 U904 ( .A(n1036), .ZN(n1191) );
XNOR2_X1 U905 ( .A(n1203), .B(G475), .ZN(n1036) );
NAND2_X1 U906 ( .A1(n1090), .A2(n1130), .ZN(n1203) );
XNOR2_X1 U907 ( .A(n1204), .B(n1205), .ZN(n1090) );
XOR2_X1 U908 ( .A(n1206), .B(n1207), .Z(n1205) );
XNOR2_X1 U909 ( .A(KEYINPUT19), .B(n1208), .ZN(n1207) );
NOR2_X1 U910 ( .A1(KEYINPUT37), .A2(n1209), .ZN(n1206) );
XNOR2_X1 U911 ( .A(n1210), .B(KEYINPUT54), .ZN(n1209) );
XOR2_X1 U912 ( .A(n1211), .B(n1212), .Z(n1204) );
NOR2_X1 U913 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
AND4_X1 U914 ( .A1(n1215), .A2(G214), .A3(n1216), .A4(n1217), .ZN(n1214) );
NOR2_X1 U915 ( .A1(n1218), .A2(n1215), .ZN(n1213) );
XOR2_X1 U916 ( .A(n1219), .B(KEYINPUT28), .Z(n1215) );
AND3_X1 U917 ( .A1(G214), .A2(n1216), .A3(n1217), .ZN(n1218) );
XOR2_X1 U918 ( .A(n1220), .B(n1221), .Z(n1211) );
NOR2_X1 U919 ( .A1(KEYINPUT11), .A2(n1222), .ZN(n1221) );
INV_X1 U920 ( .A(G131), .ZN(n1222) );
NAND2_X1 U921 ( .A1(n1223), .A2(n1224), .ZN(n1220) );
NAND2_X1 U922 ( .A1(G104), .A2(n1225), .ZN(n1224) );
XOR2_X1 U923 ( .A(KEYINPUT4), .B(n1226), .Z(n1223) );
NOR2_X1 U924 ( .A1(G104), .A2(n1225), .ZN(n1226) );
XNOR2_X1 U925 ( .A(n1227), .B(G113), .ZN(n1225) );
XNOR2_X1 U926 ( .A(n1040), .B(G478), .ZN(n1190) );
NOR2_X1 U927 ( .A1(n1085), .A2(G902), .ZN(n1040) );
XNOR2_X1 U928 ( .A(n1228), .B(n1229), .ZN(n1085) );
XNOR2_X1 U929 ( .A(n1227), .B(G107), .ZN(n1229) );
XOR2_X1 U930 ( .A(n1230), .B(n1231), .Z(n1228) );
AND3_X1 U931 ( .A1(G234), .A2(n1217), .A3(G217), .ZN(n1231) );
XOR2_X1 U932 ( .A(n1232), .B(n1233), .Z(n1230) );
XNOR2_X1 U933 ( .A(n1234), .B(n1235), .ZN(n1233) );
XOR2_X1 U934 ( .A(G128), .B(n1236), .Z(n1235) );
NOR2_X1 U935 ( .A1(G116), .A2(KEYINPUT29), .ZN(n1236) );
XOR2_X1 U936 ( .A(n1237), .B(G134), .Z(n1232) );
XNOR2_X1 U937 ( .A(KEYINPUT26), .B(KEYINPUT18), .ZN(n1237) );
NOR4_X1 U938 ( .A1(n1027), .A2(n1168), .A3(n1037), .A4(n1194), .ZN(n1154) );
INV_X1 U939 ( .A(n1188), .ZN(n1194) );
NAND2_X1 U940 ( .A1(n1001), .A2(n1238), .ZN(n1188) );
NAND4_X1 U941 ( .A1(G953), .A2(G902), .A3(n1187), .A4(n1066), .ZN(n1238) );
INV_X1 U942 ( .A(G898), .ZN(n1066) );
NAND3_X1 U943 ( .A1(n1187), .A2(n1062), .A3(G952), .ZN(n1001) );
NAND2_X1 U944 ( .A1(G237), .A2(G234), .ZN(n1187) );
INV_X1 U945 ( .A(n1026), .ZN(n1037) );
NAND2_X1 U946 ( .A1(G221), .A2(n1239), .ZN(n1026) );
NAND2_X1 U947 ( .A1(G234), .A2(n1130), .ZN(n1239) );
NAND2_X1 U948 ( .A1(n1017), .A2(n1018), .ZN(n1168) );
NAND2_X1 U949 ( .A1(G214), .A2(n1240), .ZN(n1018) );
XNOR2_X1 U950 ( .A(n1241), .B(n1129), .ZN(n1017) );
AND2_X1 U951 ( .A1(G210), .A2(n1240), .ZN(n1129) );
NAND2_X1 U952 ( .A1(n1242), .A2(n1130), .ZN(n1240) );
XNOR2_X1 U953 ( .A(G237), .B(KEYINPUT0), .ZN(n1242) );
NAND2_X1 U954 ( .A1(n1243), .A2(n1130), .ZN(n1241) );
XOR2_X1 U955 ( .A(n1244), .B(n1245), .Z(n1243) );
XNOR2_X1 U956 ( .A(n1103), .B(n1246), .ZN(n1245) );
NAND2_X1 U957 ( .A1(KEYINPUT40), .A2(n1127), .ZN(n1246) );
XNOR2_X1 U958 ( .A(n1125), .B(n1247), .ZN(n1244) );
INV_X1 U959 ( .A(n1115), .ZN(n1247) );
XNOR2_X1 U960 ( .A(n1072), .B(n1075), .ZN(n1115) );
XNOR2_X1 U961 ( .A(n1248), .B(n1249), .ZN(n1075) );
XNOR2_X1 U962 ( .A(G113), .B(KEYINPUT45), .ZN(n1248) );
XOR2_X1 U963 ( .A(n1250), .B(n1251), .Z(n1072) );
NOR2_X1 U964 ( .A1(KEYINPUT23), .A2(n1252), .ZN(n1251) );
XOR2_X1 U965 ( .A(n1253), .B(G101), .Z(n1250) );
NAND3_X1 U966 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1253) );
NAND2_X1 U967 ( .A1(n1257), .A2(n1227), .ZN(n1256) );
INV_X1 U968 ( .A(G122), .ZN(n1227) );
NAND2_X1 U969 ( .A1(KEYINPUT12), .A2(n1258), .ZN(n1257) );
XNOR2_X1 U970 ( .A(KEYINPUT17), .B(n1202), .ZN(n1258) );
NAND3_X1 U971 ( .A1(KEYINPUT12), .A2(G122), .A3(n1202), .ZN(n1255) );
OR2_X1 U972 ( .A1(n1202), .A2(KEYINPUT12), .ZN(n1254) );
NAND2_X1 U973 ( .A1(G224), .A2(n1259), .ZN(n1125) );
XOR2_X1 U974 ( .A(KEYINPUT46), .B(n1217), .Z(n1259) );
XOR2_X1 U975 ( .A(n1260), .B(n1042), .Z(n1027) );
NAND2_X1 U976 ( .A1(n1261), .A2(n1130), .ZN(n1042) );
XOR2_X1 U977 ( .A(n1262), .B(n1263), .Z(n1261) );
NOR2_X1 U978 ( .A1(n1110), .A2(n1264), .ZN(n1263) );
XOR2_X1 U979 ( .A(KEYINPUT60), .B(n1109), .Z(n1264) );
AND2_X1 U980 ( .A1(n1265), .A2(n1266), .ZN(n1109) );
NOR2_X1 U981 ( .A1(n1266), .A2(n1265), .ZN(n1110) );
XNOR2_X1 U982 ( .A(G140), .B(n1202), .ZN(n1265) );
NAND2_X1 U983 ( .A1(G227), .A2(n1217), .ZN(n1266) );
NAND2_X1 U984 ( .A1(n1267), .A2(KEYINPUT6), .ZN(n1262) );
XOR2_X1 U985 ( .A(n1113), .B(n1268), .Z(n1267) );
NOR2_X1 U986 ( .A1(KEYINPUT42), .A2(n1111), .ZN(n1268) );
XOR2_X1 U987 ( .A(n1269), .B(n1270), .Z(n1111) );
XOR2_X1 U988 ( .A(KEYINPUT15), .B(G101), .Z(n1270) );
XOR2_X1 U989 ( .A(n1054), .B(n1252), .Z(n1269) );
XOR2_X1 U990 ( .A(G107), .B(G104), .Z(n1252) );
XOR2_X1 U991 ( .A(n1271), .B(n1272), .Z(n1054) );
XNOR2_X1 U992 ( .A(n1273), .B(n1234), .ZN(n1272) );
INV_X1 U993 ( .A(n1219), .ZN(n1234) );
NOR2_X1 U994 ( .A1(KEYINPUT39), .A2(n1208), .ZN(n1273) );
NAND2_X1 U995 ( .A1(KEYINPUT13), .A2(n1043), .ZN(n1260) );
INV_X1 U996 ( .A(G469), .ZN(n1043) );
AND2_X1 U997 ( .A1(n1176), .A2(n1195), .ZN(n1022) );
INV_X1 U998 ( .A(n1177), .ZN(n1195) );
XNOR2_X1 U999 ( .A(n1274), .B(G472), .ZN(n1177) );
NAND2_X1 U1000 ( .A1(n1275), .A2(n1130), .ZN(n1274) );
INV_X1 U1001 ( .A(G902), .ZN(n1130) );
XOR2_X1 U1002 ( .A(n1101), .B(n1276), .Z(n1275) );
NOR2_X1 U1003 ( .A1(n1103), .A2(KEYINPUT56), .ZN(n1276) );
INV_X1 U1004 ( .A(n1128), .ZN(n1103) );
NAND2_X1 U1005 ( .A1(n1277), .A2(n1278), .ZN(n1128) );
NAND2_X1 U1006 ( .A1(n1271), .A2(n1279), .ZN(n1278) );
XOR2_X1 U1007 ( .A(KEYINPUT34), .B(n1280), .Z(n1277) );
NOR2_X1 U1008 ( .A1(n1271), .A2(n1279), .ZN(n1280) );
XNOR2_X1 U1009 ( .A(n1208), .B(n1219), .ZN(n1279) );
XOR2_X1 U1010 ( .A(G143), .B(KEYINPUT44), .Z(n1219) );
XNOR2_X1 U1011 ( .A(G128), .B(KEYINPUT33), .ZN(n1271) );
XOR2_X1 U1012 ( .A(n1281), .B(n1282), .Z(n1101) );
XNOR2_X1 U1013 ( .A(G101), .B(n1283), .ZN(n1282) );
NAND3_X1 U1014 ( .A1(n1217), .A2(n1216), .A3(G210), .ZN(n1283) );
INV_X1 U1015 ( .A(G237), .ZN(n1216) );
XOR2_X1 U1016 ( .A(n1113), .B(n1284), .Z(n1281) );
NOR2_X1 U1017 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
XOR2_X1 U1018 ( .A(KEYINPUT62), .B(n1287), .Z(n1286) );
NOR2_X1 U1019 ( .A1(G113), .A2(n1249), .ZN(n1287) );
AND2_X1 U1020 ( .A1(n1249), .A2(G113), .ZN(n1285) );
XNOR2_X1 U1021 ( .A(G119), .B(n1198), .ZN(n1249) );
INV_X1 U1022 ( .A(G116), .ZN(n1198) );
XOR2_X1 U1023 ( .A(n1288), .B(n1057), .Z(n1113) );
XNOR2_X1 U1024 ( .A(n1289), .B(n1290), .ZN(n1057) );
XOR2_X1 U1025 ( .A(KEYINPUT24), .B(G137), .Z(n1290) );
XNOR2_X1 U1026 ( .A(G131), .B(G134), .ZN(n1289) );
XNOR2_X1 U1027 ( .A(KEYINPUT8), .B(KEYINPUT47), .ZN(n1288) );
XOR2_X1 U1028 ( .A(n1189), .B(KEYINPUT52), .Z(n1176) );
NAND3_X1 U1029 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n1189) );
NAND2_X1 U1030 ( .A1(n1294), .A2(n1078), .ZN(n1293) );
OR3_X1 U1031 ( .A1(n1078), .A2(n1294), .A3(G902), .ZN(n1292) );
NOR2_X1 U1032 ( .A1(n1080), .A2(G234), .ZN(n1294) );
INV_X1 U1033 ( .A(G217), .ZN(n1080) );
XOR2_X1 U1034 ( .A(n1295), .B(n1296), .Z(n1078) );
XOR2_X1 U1035 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U1036 ( .A(G128), .B(G119), .Z(n1298) );
XNOR2_X1 U1037 ( .A(n1208), .B(G137), .ZN(n1297) );
INV_X1 U1038 ( .A(G146), .ZN(n1208) );
XOR2_X1 U1039 ( .A(n1299), .B(n1210), .Z(n1295) );
XNOR2_X1 U1040 ( .A(G140), .B(n1127), .ZN(n1210) );
INV_X1 U1041 ( .A(G125), .ZN(n1127) );
XNOR2_X1 U1042 ( .A(n1300), .B(n1202), .ZN(n1299) );
NAND3_X1 U1043 ( .A1(G221), .A2(n1217), .A3(G234), .ZN(n1300) );
XNOR2_X1 U1044 ( .A(n1062), .B(KEYINPUT7), .ZN(n1217) );
INV_X1 U1045 ( .A(G953), .ZN(n1062) );
NAND2_X1 U1046 ( .A1(G902), .A2(G217), .ZN(n1291) );
INV_X1 U1047 ( .A(G110), .ZN(n1202) );
endmodule


