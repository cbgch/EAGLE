//Key = 1111110010011011001101011110111011011101101001111101011111100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301;

NAND3_X1 U711 ( .A1(n996), .A2(n997), .A3(n998), .ZN(G9) );
NAND2_X1 U712 ( .A1(G107), .A2(n999), .ZN(n998) );
NAND2_X1 U713 ( .A1(KEYINPUT7), .A2(n1000), .ZN(n997) );
NAND2_X1 U714 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
INV_X1 U715 ( .A(n999), .ZN(n1002) );
XNOR2_X1 U716 ( .A(KEYINPUT10), .B(G107), .ZN(n1001) );
NAND2_X1 U717 ( .A1(n1003), .A2(n1004), .ZN(n996) );
INV_X1 U718 ( .A(KEYINPUT7), .ZN(n1004) );
NAND2_X1 U719 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
OR3_X1 U720 ( .A1(n999), .A2(G107), .A3(KEYINPUT10), .ZN(n1006) );
NAND2_X1 U721 ( .A1(KEYINPUT10), .A2(G107), .ZN(n1005) );
NOR2_X1 U722 ( .A1(n1007), .A2(n1008), .ZN(G75) );
NOR4_X1 U723 ( .A1(G953), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1008) );
NOR2_X1 U724 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NOR2_X1 U725 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR3_X1 U726 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1015) );
NOR3_X1 U727 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1017) );
NOR3_X1 U728 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1021) );
NOR2_X1 U729 ( .A1(n1025), .A2(n1026), .ZN(n1019) );
NOR2_X1 U730 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR2_X1 U731 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR3_X1 U732 ( .A1(n1023), .A2(n1031), .A3(n1032), .ZN(n1014) );
NOR4_X1 U733 ( .A1(n1026), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1032) );
AND2_X1 U734 ( .A1(n1036), .A2(KEYINPUT0), .ZN(n1035) );
NOR2_X1 U735 ( .A1(n1037), .A2(n1018), .ZN(n1034) );
NOR2_X1 U736 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR2_X1 U737 ( .A1(n1040), .A2(n1016), .ZN(n1033) );
NOR2_X1 U738 ( .A1(n1041), .A2(n1042), .ZN(n1031) );
NOR2_X1 U739 ( .A1(KEYINPUT0), .A2(n1043), .ZN(n1042) );
NOR3_X1 U740 ( .A1(n1009), .A2(G953), .A3(G952), .ZN(n1007) );
AND4_X1 U741 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1009) );
XOR2_X1 U742 ( .A(KEYINPUT62), .B(n1048), .Z(n1047) );
NOR3_X1 U743 ( .A1(n1026), .A2(n1049), .A3(n1050), .ZN(n1048) );
XNOR2_X1 U744 ( .A(G469), .B(n1051), .ZN(n1050) );
NOR2_X1 U745 ( .A1(n1052), .A2(KEYINPUT52), .ZN(n1051) );
NOR2_X1 U746 ( .A1(n1053), .A2(n1054), .ZN(n1046) );
XOR2_X1 U747 ( .A(n1055), .B(n1056), .Z(n1054) );
NAND2_X1 U748 ( .A1(KEYINPUT4), .A2(n1057), .ZN(n1055) );
XOR2_X1 U749 ( .A(n1058), .B(KEYINPUT46), .Z(n1045) );
NAND2_X1 U750 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XOR2_X1 U751 ( .A(n1061), .B(KEYINPUT43), .Z(n1059) );
XOR2_X1 U752 ( .A(n1062), .B(n1063), .Z(n1044) );
XOR2_X1 U753 ( .A(n1064), .B(n1065), .Z(G72) );
NOR2_X1 U754 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U755 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NAND2_X1 U756 ( .A1(n1070), .A2(n1071), .ZN(n1064) );
NAND2_X1 U757 ( .A1(n1072), .A2(n1067), .ZN(n1071) );
XNOR2_X1 U758 ( .A(n1073), .B(n1074), .ZN(n1072) );
NAND3_X1 U759 ( .A1(G900), .A2(n1073), .A3(G953), .ZN(n1070) );
XNOR2_X1 U760 ( .A(n1075), .B(n1076), .ZN(n1073) );
NAND2_X1 U761 ( .A1(n1077), .A2(KEYINPUT57), .ZN(n1075) );
XOR2_X1 U762 ( .A(n1078), .B(n1079), .Z(n1077) );
XOR2_X1 U763 ( .A(KEYINPUT16), .B(G140), .Z(n1079) );
XOR2_X1 U764 ( .A(n1080), .B(n1081), .Z(G69) );
XOR2_X1 U765 ( .A(n1082), .B(n1083), .Z(n1081) );
OR2_X1 U766 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U767 ( .A1(n1086), .A2(G953), .ZN(n1082) );
XOR2_X1 U768 ( .A(n1087), .B(KEYINPUT38), .Z(n1086) );
NAND2_X1 U769 ( .A1(G898), .A2(G224), .ZN(n1087) );
NOR2_X1 U770 ( .A1(n1088), .A2(G953), .ZN(n1080) );
NOR2_X1 U771 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR2_X1 U772 ( .A1(n1091), .A2(n1092), .ZN(G66) );
XOR2_X1 U773 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND2_X1 U774 ( .A1(n1095), .A2(G217), .ZN(n1094) );
NOR2_X1 U775 ( .A1(n1091), .A2(n1096), .ZN(G63) );
NOR3_X1 U776 ( .A1(n1056), .A2(n1097), .A3(n1098), .ZN(n1096) );
AND3_X1 U777 ( .A1(n1099), .A2(G478), .A3(n1095), .ZN(n1098) );
NOR2_X1 U778 ( .A1(n1100), .A2(n1099), .ZN(n1097) );
NOR2_X1 U779 ( .A1(n1101), .A2(n1057), .ZN(n1100) );
INV_X1 U780 ( .A(G478), .ZN(n1057) );
NOR2_X1 U781 ( .A1(n1091), .A2(n1102), .ZN(G60) );
NOR3_X1 U782 ( .A1(n1062), .A2(n1103), .A3(n1104), .ZN(n1102) );
AND3_X1 U783 ( .A1(n1105), .A2(G475), .A3(n1095), .ZN(n1104) );
NOR2_X1 U784 ( .A1(n1106), .A2(n1105), .ZN(n1103) );
NOR2_X1 U785 ( .A1(n1101), .A2(n1063), .ZN(n1106) );
XOR2_X1 U786 ( .A(G104), .B(n1107), .Z(G6) );
NOR2_X1 U787 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U788 ( .A1(n1091), .A2(n1110), .ZN(G57) );
XOR2_X1 U789 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U790 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U791 ( .A(n1115), .B(n1116), .Z(n1111) );
NAND2_X1 U792 ( .A1(n1095), .A2(n1117), .ZN(n1115) );
XOR2_X1 U793 ( .A(KEYINPUT34), .B(G472), .Z(n1117) );
NOR2_X1 U794 ( .A1(n1091), .A2(n1118), .ZN(G54) );
XOR2_X1 U795 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U796 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U797 ( .A(n1123), .B(n1124), .Z(n1119) );
NAND2_X1 U798 ( .A1(n1095), .A2(G469), .ZN(n1124) );
NOR2_X1 U799 ( .A1(n1125), .A2(n1101), .ZN(n1095) );
NAND2_X1 U800 ( .A1(KEYINPUT11), .A2(n1126), .ZN(n1123) );
NOR2_X1 U801 ( .A1(n1091), .A2(n1127), .ZN(G51) );
XOR2_X1 U802 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U803 ( .A(n1130), .B(n1084), .Z(n1129) );
XOR2_X1 U804 ( .A(n1131), .B(n1132), .Z(n1128) );
XNOR2_X1 U805 ( .A(KEYINPUT17), .B(n1133), .ZN(n1132) );
NAND3_X1 U806 ( .A1(n1134), .A2(n1135), .A3(G902), .ZN(n1131) );
XOR2_X1 U807 ( .A(KEYINPUT23), .B(n1101), .Z(n1135) );
INV_X1 U808 ( .A(n1011), .ZN(n1101) );
NAND3_X1 U809 ( .A1(n1074), .A2(n1136), .A3(n1137), .ZN(n1011) );
XOR2_X1 U810 ( .A(n1089), .B(KEYINPUT12), .Z(n1137) );
NAND4_X1 U811 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1089) );
NAND3_X1 U812 ( .A1(n1142), .A2(n1020), .A3(n1143), .ZN(n1139) );
XOR2_X1 U813 ( .A(n1144), .B(KEYINPUT9), .Z(n1143) );
NAND3_X1 U814 ( .A1(n1145), .A2(n1038), .A3(n1146), .ZN(n1138) );
INV_X1 U815 ( .A(n1090), .ZN(n1136) );
NAND4_X1 U816 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n999), .ZN(n1090) );
NAND3_X1 U817 ( .A1(n1150), .A2(n1151), .A3(n1038), .ZN(n999) );
NAND2_X1 U818 ( .A1(n1152), .A2(n1153), .ZN(n1147) );
XOR2_X1 U819 ( .A(n1109), .B(KEYINPUT35), .Z(n1152) );
NAND4_X1 U820 ( .A1(n1039), .A2(n1150), .A3(n1028), .A4(n1144), .ZN(n1109) );
AND2_X1 U821 ( .A1(n1154), .A2(n1155), .ZN(n1074) );
AND4_X1 U822 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
NOR4_X1 U823 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1154) );
NOR3_X1 U824 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1162) );
INV_X1 U825 ( .A(n1167), .ZN(n1161) );
NOR2_X1 U826 ( .A1(n1067), .A2(G952), .ZN(n1091) );
XNOR2_X1 U827 ( .A(G146), .B(n1158), .ZN(G48) );
NAND3_X1 U828 ( .A1(n1168), .A2(n1039), .A3(n1169), .ZN(n1158) );
XOR2_X1 U829 ( .A(n1157), .B(n1170), .Z(G45) );
NAND2_X1 U830 ( .A1(KEYINPUT30), .A2(G143), .ZN(n1170) );
NAND4_X1 U831 ( .A1(n1145), .A2(n1168), .A3(n1171), .A4(n1172), .ZN(n1157) );
XOR2_X1 U832 ( .A(n1173), .B(n1156), .Z(G42) );
NAND4_X1 U833 ( .A1(n1174), .A2(n1039), .A3(n1175), .A4(n1041), .ZN(n1156) );
XOR2_X1 U834 ( .A(n1176), .B(n1167), .Z(G39) );
NAND3_X1 U835 ( .A1(n1175), .A2(n1041), .A3(n1142), .ZN(n1167) );
XOR2_X1 U836 ( .A(G134), .B(n1160), .Z(G36) );
AND4_X1 U837 ( .A1(n1145), .A2(n1175), .A3(n1041), .A4(n1038), .ZN(n1160) );
XOR2_X1 U838 ( .A(n1177), .B(n1178), .Z(G33) );
NAND2_X1 U839 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NAND3_X1 U840 ( .A1(n1041), .A2(n1181), .A3(n1182), .ZN(n1180) );
INV_X1 U841 ( .A(KEYINPUT39), .ZN(n1182) );
INV_X1 U842 ( .A(n1026), .ZN(n1041) );
NAND2_X1 U843 ( .A1(n1163), .A2(KEYINPUT39), .ZN(n1179) );
NOR2_X1 U844 ( .A1(n1181), .A2(n1026), .ZN(n1163) );
NAND2_X1 U845 ( .A1(n1183), .A2(n1022), .ZN(n1026) );
NAND3_X1 U846 ( .A1(n1039), .A2(n1175), .A3(n1145), .ZN(n1181) );
NAND2_X1 U847 ( .A1(KEYINPUT54), .A2(n1184), .ZN(n1177) );
INV_X1 U848 ( .A(G131), .ZN(n1184) );
XOR2_X1 U849 ( .A(n1185), .B(n1186), .Z(G30) );
NAND3_X1 U850 ( .A1(n1038), .A2(n1187), .A3(n1168), .ZN(n1186) );
INV_X1 U851 ( .A(n1166), .ZN(n1168) );
NAND2_X1 U852 ( .A1(n1175), .A2(n1153), .ZN(n1166) );
AND2_X1 U853 ( .A1(n1028), .A2(n1188), .ZN(n1175) );
XOR2_X1 U854 ( .A(KEYINPUT63), .B(n1169), .Z(n1187) );
INV_X1 U855 ( .A(n1164), .ZN(n1169) );
XNOR2_X1 U856 ( .A(G101), .B(n1148), .ZN(G3) );
NAND3_X1 U857 ( .A1(n1145), .A2(n1151), .A3(n1189), .ZN(n1148) );
XOR2_X1 U858 ( .A(n1159), .B(n1190), .Z(G27) );
NAND2_X1 U859 ( .A1(KEYINPUT55), .A2(G125), .ZN(n1190) );
NAND4_X1 U860 ( .A1(n1020), .A2(n1174), .A3(n1039), .A4(n1188), .ZN(n1159) );
NAND2_X1 U861 ( .A1(n1013), .A2(n1191), .ZN(n1188) );
NAND4_X1 U862 ( .A1(G902), .A2(G953), .A3(n1192), .A4(n1069), .ZN(n1191) );
INV_X1 U863 ( .A(G900), .ZN(n1069) );
XOR2_X1 U864 ( .A(n1140), .B(n1193), .Z(G24) );
NOR2_X1 U865 ( .A1(G122), .A2(KEYINPUT31), .ZN(n1193) );
NAND4_X1 U866 ( .A1(n1146), .A2(n1150), .A3(n1171), .A4(n1172), .ZN(n1140) );
INV_X1 U867 ( .A(n1018), .ZN(n1150) );
NAND2_X1 U868 ( .A1(n1194), .A2(n1195), .ZN(n1018) );
INV_X1 U869 ( .A(n1053), .ZN(n1195) );
XOR2_X1 U870 ( .A(G119), .B(n1196), .Z(G21) );
AND2_X1 U871 ( .A1(n1142), .A2(n1146), .ZN(n1196) );
NOR2_X1 U872 ( .A1(n1016), .A2(n1164), .ZN(n1142) );
NAND2_X1 U873 ( .A1(n1053), .A2(n1197), .ZN(n1164) );
NAND2_X1 U874 ( .A1(n1198), .A2(n1199), .ZN(G18) );
NAND2_X1 U875 ( .A1(G116), .A2(n1200), .ZN(n1199) );
XOR2_X1 U876 ( .A(n1201), .B(KEYINPUT60), .Z(n1198) );
OR2_X1 U877 ( .A1(n1200), .A2(G116), .ZN(n1201) );
NAND4_X1 U878 ( .A1(n1020), .A2(n1145), .A3(n1038), .A4(n1202), .ZN(n1200) );
XNOR2_X1 U879 ( .A(KEYINPUT28), .B(n1144), .ZN(n1202) );
INV_X1 U880 ( .A(n1165), .ZN(n1038) );
NAND2_X1 U881 ( .A1(n1203), .A2(n1171), .ZN(n1165) );
XOR2_X1 U882 ( .A(n1141), .B(n1204), .Z(G15) );
XNOR2_X1 U883 ( .A(G113), .B(KEYINPUT59), .ZN(n1204) );
NAND3_X1 U884 ( .A1(n1145), .A2(n1039), .A3(n1146), .ZN(n1141) );
AND2_X1 U885 ( .A1(n1020), .A2(n1144), .ZN(n1146) );
NOR2_X1 U886 ( .A1(n1023), .A2(n1108), .ZN(n1020) );
OR2_X1 U887 ( .A1(n1029), .A2(n1049), .ZN(n1023) );
INV_X1 U888 ( .A(n1030), .ZN(n1049) );
NOR2_X1 U889 ( .A1(n1171), .A2(n1205), .ZN(n1039) );
INV_X1 U890 ( .A(n1172), .ZN(n1205) );
INV_X1 U891 ( .A(n1040), .ZN(n1145) );
NAND2_X1 U892 ( .A1(n1053), .A2(n1194), .ZN(n1040) );
XOR2_X1 U893 ( .A(n1197), .B(KEYINPUT2), .Z(n1194) );
XNOR2_X1 U894 ( .A(n1206), .B(n1149), .ZN(G12) );
NAND2_X1 U895 ( .A1(n1036), .A2(n1151), .ZN(n1149) );
AND3_X1 U896 ( .A1(n1153), .A2(n1144), .A3(n1028), .ZN(n1151) );
AND2_X1 U897 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND2_X1 U898 ( .A1(G221), .A2(n1207), .ZN(n1030) );
NAND2_X1 U899 ( .A1(G234), .A2(n1125), .ZN(n1207) );
XOR2_X1 U900 ( .A(n1052), .B(G469), .Z(n1029) );
AND2_X1 U901 ( .A1(n1208), .A2(n1125), .ZN(n1052) );
XOR2_X1 U902 ( .A(n1209), .B(n1121), .Z(n1208) );
XNOR2_X1 U903 ( .A(n1210), .B(n1211), .ZN(n1121) );
XOR2_X1 U904 ( .A(G107), .B(G101), .Z(n1211) );
XOR2_X1 U905 ( .A(n1212), .B(n1076), .Z(n1210) );
INV_X1 U906 ( .A(n1116), .ZN(n1076) );
NAND2_X1 U907 ( .A1(KEYINPUT56), .A2(G104), .ZN(n1212) );
NOR2_X1 U908 ( .A1(KEYINPUT6), .A2(n1213), .ZN(n1209) );
XOR2_X1 U909 ( .A(n1126), .B(n1122), .Z(n1213) );
XOR2_X1 U910 ( .A(G140), .B(n1214), .Z(n1122) );
NOR2_X1 U911 ( .A1(G953), .A2(n1068), .ZN(n1214) );
INV_X1 U912 ( .A(G227), .ZN(n1068) );
NAND2_X1 U913 ( .A1(n1013), .A2(n1215), .ZN(n1144) );
NAND3_X1 U914 ( .A1(n1085), .A2(n1192), .A3(G902), .ZN(n1215) );
NOR2_X1 U915 ( .A1(n1067), .A2(G898), .ZN(n1085) );
NAND3_X1 U916 ( .A1(n1192), .A2(n1067), .A3(G952), .ZN(n1013) );
NAND2_X1 U917 ( .A1(G237), .A2(G234), .ZN(n1192) );
INV_X1 U918 ( .A(n1108), .ZN(n1153) );
NAND2_X1 U919 ( .A1(n1024), .A2(n1022), .ZN(n1108) );
NAND2_X1 U920 ( .A1(G214), .A2(n1216), .ZN(n1022) );
INV_X1 U921 ( .A(n1183), .ZN(n1024) );
XOR2_X1 U922 ( .A(n1217), .B(n1134), .Z(n1183) );
AND2_X1 U923 ( .A1(G210), .A2(n1216), .ZN(n1134) );
NAND2_X1 U924 ( .A1(n1218), .A2(n1125), .ZN(n1216) );
INV_X1 U925 ( .A(G237), .ZN(n1218) );
NAND2_X1 U926 ( .A1(n1219), .A2(n1125), .ZN(n1217) );
XOR2_X1 U927 ( .A(n1220), .B(n1221), .Z(n1219) );
XNOR2_X1 U928 ( .A(n1222), .B(n1130), .ZN(n1221) );
XNOR2_X1 U929 ( .A(n1223), .B(G125), .ZN(n1130) );
NAND2_X1 U930 ( .A1(KEYINPUT40), .A2(n1084), .ZN(n1222) );
XNOR2_X1 U931 ( .A(n1224), .B(n1225), .ZN(n1084) );
XOR2_X1 U932 ( .A(n1226), .B(n1227), .Z(n1225) );
XNOR2_X1 U933 ( .A(n1228), .B(n1229), .ZN(n1227) );
NOR2_X1 U934 ( .A1(KEYINPUT41), .A2(n1230), .ZN(n1229) );
NAND2_X1 U935 ( .A1(n1231), .A2(KEYINPUT18), .ZN(n1228) );
XOR2_X1 U936 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U937 ( .A(KEYINPUT20), .B(G107), .Z(n1233) );
XNOR2_X1 U938 ( .A(G101), .B(n1234), .ZN(n1224) );
XOR2_X1 U939 ( .A(KEYINPUT25), .B(G110), .Z(n1234) );
XNOR2_X1 U940 ( .A(n1235), .B(KEYINPUT58), .ZN(n1220) );
NAND2_X1 U941 ( .A1(KEYINPUT26), .A2(n1133), .ZN(n1235) );
NAND2_X1 U942 ( .A1(G224), .A2(n1067), .ZN(n1133) );
INV_X1 U943 ( .A(n1043), .ZN(n1036) );
NAND2_X1 U944 ( .A1(n1189), .A2(n1174), .ZN(n1043) );
AND2_X1 U945 ( .A1(n1236), .A2(n1197), .ZN(n1174) );
NAND2_X1 U946 ( .A1(n1061), .A2(n1060), .ZN(n1197) );
NAND3_X1 U947 ( .A1(n1093), .A2(n1125), .A3(n1237), .ZN(n1060) );
NAND2_X1 U948 ( .A1(G217), .A2(n1238), .ZN(n1237) );
NAND2_X1 U949 ( .A1(G217), .A2(n1239), .ZN(n1061) );
NAND2_X1 U950 ( .A1(n1240), .A2(n1125), .ZN(n1239) );
OR2_X1 U951 ( .A1(n1093), .A2(G234), .ZN(n1240) );
NAND2_X1 U952 ( .A1(n1241), .A2(n1242), .ZN(n1093) );
NAND3_X1 U953 ( .A1(n1243), .A2(n1244), .A3(n1245), .ZN(n1242) );
NAND2_X1 U954 ( .A1(n1246), .A2(n1247), .ZN(n1241) );
NAND2_X1 U955 ( .A1(n1243), .A2(n1244), .ZN(n1247) );
NAND2_X1 U956 ( .A1(n1248), .A2(n1249), .ZN(n1244) );
XOR2_X1 U957 ( .A(KEYINPUT50), .B(n1250), .Z(n1249) );
XNOR2_X1 U958 ( .A(n1251), .B(KEYINPUT37), .ZN(n1243) );
OR2_X1 U959 ( .A1(n1250), .A2(n1248), .ZN(n1251) );
XNOR2_X1 U960 ( .A(n1252), .B(G146), .ZN(n1248) );
NAND2_X1 U961 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NAND2_X1 U962 ( .A1(n1255), .A2(G125), .ZN(n1254) );
NAND2_X1 U963 ( .A1(n1256), .A2(n1078), .ZN(n1253) );
XOR2_X1 U964 ( .A(n1255), .B(KEYINPUT47), .Z(n1256) );
XNOR2_X1 U965 ( .A(n1257), .B(n1258), .ZN(n1250) );
XOR2_X1 U966 ( .A(n1126), .B(G128), .Z(n1257) );
XOR2_X1 U967 ( .A(KEYINPUT29), .B(n1245), .Z(n1246) );
XOR2_X1 U968 ( .A(n1259), .B(n1176), .Z(n1245) );
INV_X1 U969 ( .A(G137), .ZN(n1176) );
NAND3_X1 U970 ( .A1(G234), .A2(n1067), .A3(G221), .ZN(n1259) );
XOR2_X1 U971 ( .A(n1053), .B(KEYINPUT19), .Z(n1236) );
XOR2_X1 U972 ( .A(n1260), .B(n1261), .Z(n1053) );
XOR2_X1 U973 ( .A(KEYINPUT49), .B(G472), .Z(n1261) );
NAND2_X1 U974 ( .A1(n1262), .A2(n1125), .ZN(n1260) );
INV_X1 U975 ( .A(G902), .ZN(n1125) );
XOR2_X1 U976 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U977 ( .A(n1265), .B(KEYINPUT5), .ZN(n1264) );
NAND2_X1 U978 ( .A1(KEYINPUT14), .A2(n1116), .ZN(n1265) );
XOR2_X1 U979 ( .A(n1266), .B(n1267), .Z(n1116) );
XOR2_X1 U980 ( .A(G137), .B(G134), .Z(n1267) );
XOR2_X1 U981 ( .A(n1223), .B(G131), .Z(n1266) );
XOR2_X1 U982 ( .A(n1185), .B(n1268), .Z(n1223) );
XNOR2_X1 U983 ( .A(n1114), .B(n1113), .ZN(n1263) );
XOR2_X1 U984 ( .A(n1226), .B(KEYINPUT13), .Z(n1113) );
XNOR2_X1 U985 ( .A(n1269), .B(n1258), .ZN(n1226) );
XOR2_X1 U986 ( .A(G119), .B(KEYINPUT8), .Z(n1258) );
XNOR2_X1 U987 ( .A(G113), .B(G116), .ZN(n1269) );
XNOR2_X1 U988 ( .A(n1270), .B(G101), .ZN(n1114) );
NAND2_X1 U989 ( .A1(G210), .A2(n1271), .ZN(n1270) );
INV_X1 U990 ( .A(n1016), .ZN(n1189) );
NAND2_X1 U991 ( .A1(n1203), .A2(n1272), .ZN(n1016) );
XOR2_X1 U992 ( .A(KEYINPUT48), .B(n1171), .Z(n1272) );
XOR2_X1 U993 ( .A(n1056), .B(G478), .Z(n1171) );
NOR2_X1 U994 ( .A1(n1099), .A2(G902), .ZN(n1056) );
XOR2_X1 U995 ( .A(n1273), .B(n1274), .Z(n1099) );
NOR3_X1 U996 ( .A1(n1238), .A2(n1275), .A3(n1276), .ZN(n1274) );
INV_X1 U997 ( .A(G217), .ZN(n1276) );
XOR2_X1 U998 ( .A(n1067), .B(KEYINPUT36), .Z(n1275) );
INV_X1 U999 ( .A(G953), .ZN(n1067) );
INV_X1 U1000 ( .A(G234), .ZN(n1238) );
NAND3_X1 U1001 ( .A1(n1277), .A2(n1278), .A3(KEYINPUT3), .ZN(n1273) );
OR3_X1 U1002 ( .A1(n1279), .A2(n1280), .A3(KEYINPUT15), .ZN(n1278) );
NAND2_X1 U1003 ( .A1(n1281), .A2(KEYINPUT15), .ZN(n1277) );
XNOR2_X1 U1004 ( .A(n1282), .B(n1280), .ZN(n1281) );
XNOR2_X1 U1005 ( .A(n1283), .B(n1284), .ZN(n1280) );
XOR2_X1 U1006 ( .A(KEYINPUT21), .B(G134), .Z(n1284) );
NAND2_X1 U1007 ( .A1(KEYINPUT45), .A2(n1285), .ZN(n1283) );
XNOR2_X1 U1008 ( .A(G143), .B(n1286), .ZN(n1285) );
NAND2_X1 U1009 ( .A1(KEYINPUT1), .A2(n1185), .ZN(n1286) );
INV_X1 U1010 ( .A(G128), .ZN(n1185) );
NAND2_X1 U1011 ( .A1(n1279), .A2(n1287), .ZN(n1282) );
XOR2_X1 U1012 ( .A(KEYINPUT61), .B(KEYINPUT53), .Z(n1287) );
XOR2_X1 U1013 ( .A(n1288), .B(n1230), .Z(n1279) );
XNOR2_X1 U1014 ( .A(G116), .B(G107), .ZN(n1288) );
XNOR2_X1 U1015 ( .A(n1172), .B(KEYINPUT44), .ZN(n1203) );
XNOR2_X1 U1016 ( .A(n1289), .B(n1290), .ZN(n1172) );
XOR2_X1 U1017 ( .A(KEYINPUT42), .B(n1062), .Z(n1290) );
NOR2_X1 U1018 ( .A1(n1105), .A2(G902), .ZN(n1062) );
XNOR2_X1 U1019 ( .A(n1291), .B(n1292), .ZN(n1105) );
XOR2_X1 U1020 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U1021 ( .A(G131), .B(n1295), .Z(n1294) );
NOR2_X1 U1022 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
XOR2_X1 U1023 ( .A(n1298), .B(KEYINPUT24), .Z(n1297) );
NAND2_X1 U1024 ( .A1(n1299), .A2(n1232), .ZN(n1298) );
NOR2_X1 U1025 ( .A1(n1299), .A2(n1232), .ZN(n1296) );
INV_X1 U1026 ( .A(G104), .ZN(n1232) );
XNOR2_X1 U1027 ( .A(G113), .B(n1230), .ZN(n1299) );
XOR2_X1 U1028 ( .A(G122), .B(KEYINPUT27), .Z(n1230) );
AND2_X1 U1029 ( .A1(n1271), .A2(G214), .ZN(n1293) );
NOR2_X1 U1030 ( .A1(G953), .A2(G237), .ZN(n1271) );
XOR2_X1 U1031 ( .A(n1255), .B(n1300), .Z(n1291) );
XOR2_X1 U1032 ( .A(n1301), .B(n1268), .Z(n1300) );
XOR2_X1 U1033 ( .A(G143), .B(G146), .Z(n1268) );
NOR2_X1 U1034 ( .A1(KEYINPUT22), .A2(n1078), .ZN(n1301) );
INV_X1 U1035 ( .A(G125), .ZN(n1078) );
XOR2_X1 U1036 ( .A(n1173), .B(KEYINPUT33), .Z(n1255) );
INV_X1 U1037 ( .A(G140), .ZN(n1173) );
NAND2_X1 U1038 ( .A1(KEYINPUT32), .A2(n1063), .ZN(n1289) );
INV_X1 U1039 ( .A(G475), .ZN(n1063) );
NAND2_X1 U1040 ( .A1(KEYINPUT51), .A2(n1126), .ZN(n1206) );
INV_X1 U1041 ( .A(G110), .ZN(n1126) );
endmodule


