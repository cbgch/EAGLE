//Key = 1000101001100011011011110100110011010010000010011010010001101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385;

XNOR2_X1 U753 ( .A(G107), .B(n1046), .ZN(G9) );
NOR2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(G75) );
NOR4_X1 U755 ( .A1(n1049), .A2(n1050), .A3(KEYINPUT19), .A4(G953), .ZN(n1048) );
NAND2_X1 U756 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NAND3_X1 U757 ( .A1(n1053), .A2(n1054), .A3(KEYINPUT63), .ZN(n1052) );
NAND2_X1 U758 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NAND3_X1 U759 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
XNOR2_X1 U760 ( .A(n1060), .B(n1061), .ZN(n1059) );
NAND4_X1 U761 ( .A1(n1062), .A2(n1063), .A3(n1061), .A4(n1064), .ZN(n1055) );
NOR3_X1 U762 ( .A1(n1065), .A2(n1060), .A3(n1066), .ZN(n1064) );
NOR2_X1 U763 ( .A1(n1067), .A2(n1058), .ZN(n1066) );
NOR2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
INV_X1 U765 ( .A(n1057), .ZN(n1069) );
NOR2_X1 U766 ( .A1(n1070), .A2(n1071), .ZN(n1057) );
NOR2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1068) );
NOR2_X1 U768 ( .A1(n1074), .A2(n1075), .ZN(n1065) );
NOR2_X1 U769 ( .A1(n1076), .A2(n1071), .ZN(n1075) );
NOR2_X1 U770 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
OR2_X1 U771 ( .A1(n1079), .A2(n1080), .ZN(n1063) );
NAND3_X1 U772 ( .A1(n1081), .A2(n1079), .A3(n1080), .ZN(n1062) );
NAND2_X1 U773 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND4_X1 U774 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1083) );
NOR3_X1 U775 ( .A1(n1050), .A2(G953), .A3(G952), .ZN(n1047) );
AND4_X1 U776 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1050) );
NOR4_X1 U777 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1091) );
XNOR2_X1 U778 ( .A(n1096), .B(n1097), .ZN(n1095) );
NOR2_X1 U779 ( .A1(KEYINPUT41), .A2(n1098), .ZN(n1097) );
XNOR2_X1 U780 ( .A(n1099), .B(n1100), .ZN(n1092) );
NOR2_X1 U781 ( .A1(G475), .A2(KEYINPUT24), .ZN(n1100) );
AND3_X1 U782 ( .A1(n1101), .A2(n1079), .A3(n1102), .ZN(n1090) );
INV_X1 U783 ( .A(n1103), .ZN(n1079) );
XNOR2_X1 U784 ( .A(n1104), .B(n1105), .ZN(n1088) );
NAND2_X1 U785 ( .A1(KEYINPUT17), .A2(n1106), .ZN(n1105) );
XOR2_X1 U786 ( .A(n1107), .B(n1108), .Z(G72) );
NOR2_X1 U787 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U788 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
INV_X1 U789 ( .A(n1113), .ZN(n1112) );
NOR2_X1 U790 ( .A1(G227), .A2(n1114), .ZN(n1111) );
NOR2_X1 U791 ( .A1(n1115), .A2(n1114), .ZN(n1109) );
NOR2_X1 U792 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
INV_X1 U793 ( .A(G900), .ZN(n1117) );
NOR2_X1 U794 ( .A1(G227), .A2(n1113), .ZN(n1116) );
XNOR2_X1 U795 ( .A(n1118), .B(n1119), .ZN(n1113) );
XNOR2_X1 U796 ( .A(n1120), .B(n1121), .ZN(n1119) );
NAND2_X1 U797 ( .A1(KEYINPUT47), .A2(n1122), .ZN(n1120) );
XNOR2_X1 U798 ( .A(n1123), .B(n1124), .ZN(n1118) );
NOR2_X1 U799 ( .A1(G134), .A2(KEYINPUT8), .ZN(n1124) );
NOR2_X1 U800 ( .A1(KEYINPUT49), .A2(n1125), .ZN(n1123) );
NAND2_X1 U801 ( .A1(n1114), .A2(n1126), .ZN(n1107) );
XOR2_X1 U802 ( .A(n1127), .B(n1128), .Z(G69) );
XOR2_X1 U803 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U804 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XNOR2_X1 U805 ( .A(n1133), .B(n1134), .ZN(n1132) );
XOR2_X1 U806 ( .A(n1135), .B(n1136), .Z(n1133) );
NAND2_X1 U807 ( .A1(KEYINPUT10), .A2(n1137), .ZN(n1135) );
NOR2_X1 U808 ( .A1(G898), .A2(n1114), .ZN(n1131) );
NAND2_X1 U809 ( .A1(n1138), .A2(n1114), .ZN(n1129) );
NAND2_X1 U810 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XNOR2_X1 U811 ( .A(KEYINPUT0), .B(n1141), .ZN(n1140) );
INV_X1 U812 ( .A(n1142), .ZN(n1139) );
NAND2_X1 U813 ( .A1(G953), .A2(n1143), .ZN(n1127) );
NAND2_X1 U814 ( .A1(G898), .A2(G224), .ZN(n1143) );
NOR2_X1 U815 ( .A1(n1144), .A2(n1145), .ZN(G66) );
XNOR2_X1 U816 ( .A(n1146), .B(n1147), .ZN(n1145) );
NOR2_X1 U817 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NOR2_X1 U818 ( .A1(n1144), .A2(n1150), .ZN(G63) );
NOR3_X1 U819 ( .A1(n1104), .A2(n1151), .A3(n1152), .ZN(n1150) );
NOR3_X1 U820 ( .A1(n1153), .A2(n1106), .A3(n1149), .ZN(n1152) );
NOR2_X1 U821 ( .A1(n1154), .A2(n1155), .ZN(n1151) );
NOR2_X1 U822 ( .A1(n1051), .A2(n1106), .ZN(n1154) );
NOR2_X1 U823 ( .A1(n1144), .A2(n1156), .ZN(G60) );
NOR3_X1 U824 ( .A1(n1099), .A2(n1157), .A3(n1158), .ZN(n1156) );
NOR4_X1 U825 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1149), .ZN(n1158) );
INV_X1 U826 ( .A(n1162), .ZN(n1159) );
NOR2_X1 U827 ( .A1(n1163), .A2(n1162), .ZN(n1157) );
NOR3_X1 U828 ( .A1(n1160), .A2(n1051), .A3(n1161), .ZN(n1163) );
INV_X1 U829 ( .A(KEYINPUT23), .ZN(n1160) );
XNOR2_X1 U830 ( .A(G104), .B(n1141), .ZN(G6) );
NOR2_X1 U831 ( .A1(n1144), .A2(n1164), .ZN(G57) );
XOR2_X1 U832 ( .A(n1165), .B(n1166), .Z(n1164) );
XNOR2_X1 U833 ( .A(n1167), .B(n1168), .ZN(n1166) );
NAND3_X1 U834 ( .A1(n1169), .A2(n1170), .A3(KEYINPUT14), .ZN(n1168) );
NAND2_X1 U835 ( .A1(KEYINPUT33), .A2(n1171), .ZN(n1170) );
XOR2_X1 U836 ( .A(n1172), .B(n1173), .Z(n1171) );
OR3_X1 U837 ( .A1(n1172), .A2(n1173), .A3(KEYINPUT33), .ZN(n1169) );
NAND3_X1 U838 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1172) );
NAND2_X1 U839 ( .A1(KEYINPUT3), .A2(n1177), .ZN(n1176) );
NAND3_X1 U840 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1175) );
NAND2_X1 U841 ( .A1(n1181), .A2(n1182), .ZN(n1174) );
NAND2_X1 U842 ( .A1(n1183), .A2(n1179), .ZN(n1182) );
INV_X1 U843 ( .A(KEYINPUT3), .ZN(n1179) );
XNOR2_X1 U844 ( .A(KEYINPUT27), .B(n1177), .ZN(n1183) );
XOR2_X1 U845 ( .A(n1184), .B(n1185), .Z(n1165) );
NOR2_X1 U846 ( .A1(n1186), .A2(n1149), .ZN(n1185) );
NAND2_X1 U847 ( .A1(KEYINPUT28), .A2(n1187), .ZN(n1184) );
NOR2_X1 U848 ( .A1(n1144), .A2(n1188), .ZN(G54) );
XOR2_X1 U849 ( .A(n1189), .B(n1190), .Z(n1188) );
XNOR2_X1 U850 ( .A(n1177), .B(n1191), .ZN(n1190) );
XOR2_X1 U851 ( .A(n1192), .B(n1193), .Z(n1189) );
NOR2_X1 U852 ( .A1(n1096), .A2(n1149), .ZN(n1193) );
NOR2_X1 U853 ( .A1(n1194), .A2(n1195), .ZN(n1192) );
XOR2_X1 U854 ( .A(n1196), .B(n1197), .Z(n1195) );
XOR2_X1 U855 ( .A(n1198), .B(n1199), .Z(n1197) );
NAND2_X1 U856 ( .A1(KEYINPUT15), .A2(n1200), .ZN(n1199) );
NAND2_X1 U857 ( .A1(n1201), .A2(n1202), .ZN(n1198) );
NOR2_X1 U858 ( .A1(n1201), .A2(n1202), .ZN(n1194) );
INV_X1 U859 ( .A(KEYINPUT37), .ZN(n1202) );
NOR2_X1 U860 ( .A1(n1144), .A2(n1203), .ZN(G51) );
XOR2_X1 U861 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U862 ( .A(n1206), .B(n1207), .Z(n1205) );
NOR2_X1 U863 ( .A1(KEYINPUT40), .A2(n1208), .ZN(n1206) );
INV_X1 U864 ( .A(n1209), .ZN(n1208) );
XOR2_X1 U865 ( .A(n1210), .B(n1211), .Z(n1204) );
NOR2_X1 U866 ( .A1(n1212), .A2(n1149), .ZN(n1211) );
OR2_X1 U867 ( .A1(n1213), .A2(n1051), .ZN(n1149) );
NOR3_X1 U868 ( .A1(n1142), .A2(n1214), .A3(n1126), .ZN(n1051) );
NAND4_X1 U869 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1126) );
NOR4_X1 U870 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1218) );
NOR2_X1 U871 ( .A1(n1223), .A2(n1224), .ZN(n1217) );
NOR3_X1 U872 ( .A1(n1225), .A2(n1226), .A3(n1227), .ZN(n1224) );
XNOR2_X1 U873 ( .A(KEYINPUT50), .B(n1070), .ZN(n1225) );
INV_X1 U874 ( .A(n1141), .ZN(n1214) );
NAND3_X1 U875 ( .A1(n1228), .A2(n1058), .A3(n1078), .ZN(n1141) );
NAND4_X1 U876 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1142) );
AND4_X1 U877 ( .A1(n1233), .A2(n1046), .A3(n1234), .A4(n1235), .ZN(n1232) );
NAND3_X1 U878 ( .A1(n1077), .A2(n1058), .A3(n1228), .ZN(n1046) );
NAND4_X1 U879 ( .A1(n1236), .A2(n1078), .A3(n1072), .A4(n1237), .ZN(n1231) );
XNOR2_X1 U880 ( .A(KEYINPUT53), .B(n1238), .ZN(n1237) );
NOR2_X1 U881 ( .A1(n1239), .A2(G952), .ZN(n1144) );
XNOR2_X1 U882 ( .A(n1114), .B(KEYINPUT48), .ZN(n1239) );
NAND3_X1 U883 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(G48) );
NAND2_X1 U884 ( .A1(KEYINPUT16), .A2(n1223), .ZN(n1242) );
NAND3_X1 U885 ( .A1(n1243), .A2(n1244), .A3(G146), .ZN(n1241) );
NAND2_X1 U886 ( .A1(n1245), .A2(n1246), .ZN(n1240) );
NAND2_X1 U887 ( .A1(n1247), .A2(n1244), .ZN(n1245) );
INV_X1 U888 ( .A(KEYINPUT16), .ZN(n1244) );
XNOR2_X1 U889 ( .A(n1223), .B(KEYINPUT43), .ZN(n1247) );
INV_X1 U890 ( .A(n1243), .ZN(n1223) );
NAND3_X1 U891 ( .A1(n1248), .A2(n1078), .A3(n1249), .ZN(n1243) );
XOR2_X1 U892 ( .A(n1216), .B(n1250), .Z(G45) );
NAND2_X1 U893 ( .A1(KEYINPUT25), .A2(G143), .ZN(n1250) );
NAND4_X1 U894 ( .A1(n1251), .A2(n1249), .A3(n1072), .A4(n1252), .ZN(n1216) );
NAND3_X1 U895 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(G42) );
OR2_X1 U896 ( .A1(n1256), .A2(KEYINPUT29), .ZN(n1255) );
NAND3_X1 U897 ( .A1(KEYINPUT29), .A2(n1256), .A3(n1222), .ZN(n1254) );
NAND2_X1 U898 ( .A1(n1257), .A2(n1258), .ZN(n1253) );
INV_X1 U899 ( .A(n1222), .ZN(n1258) );
NOR3_X1 U900 ( .A1(n1085), .A2(n1084), .A3(n1227), .ZN(n1222) );
INV_X1 U901 ( .A(n1073), .ZN(n1084) );
NAND2_X1 U902 ( .A1(KEYINPUT29), .A2(n1259), .ZN(n1257) );
XNOR2_X1 U903 ( .A(KEYINPUT35), .B(n1256), .ZN(n1259) );
XOR2_X1 U904 ( .A(G137), .B(n1260), .Z(G39) );
NOR4_X1 U905 ( .A1(KEYINPUT2), .A2(n1226), .A3(n1227), .A4(n1070), .ZN(n1260) );
INV_X1 U906 ( .A(n1074), .ZN(n1070) );
INV_X1 U907 ( .A(n1248), .ZN(n1226) );
XOR2_X1 U908 ( .A(G134), .B(n1221), .Z(G36) );
NOR3_X1 U909 ( .A1(n1086), .A2(n1087), .A3(n1227), .ZN(n1221) );
INV_X1 U910 ( .A(n1077), .ZN(n1086) );
XNOR2_X1 U911 ( .A(n1122), .B(n1220), .ZN(G33) );
NOR3_X1 U912 ( .A1(n1085), .A2(n1087), .A3(n1227), .ZN(n1220) );
NAND4_X1 U913 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1102), .ZN(n1227) );
INV_X1 U914 ( .A(n1071), .ZN(n1262) );
NAND2_X1 U915 ( .A1(n1082), .A2(n1080), .ZN(n1071) );
XNOR2_X1 U916 ( .A(n1103), .B(KEYINPUT42), .ZN(n1082) );
INV_X1 U917 ( .A(n1072), .ZN(n1087) );
XOR2_X1 U918 ( .A(G128), .B(n1219), .Z(G30) );
AND3_X1 U919 ( .A1(n1248), .A2(n1077), .A3(n1249), .ZN(n1219) );
AND3_X1 U920 ( .A1(n1261), .A2(n1263), .A3(n1264), .ZN(n1249) );
XNOR2_X1 U921 ( .A(G101), .B(n1229), .ZN(G3) );
NAND3_X1 U922 ( .A1(n1228), .A2(n1072), .A3(n1074), .ZN(n1229) );
NAND2_X1 U923 ( .A1(n1265), .A2(n1266), .ZN(G27) );
NAND2_X1 U924 ( .A1(G125), .A2(n1215), .ZN(n1266) );
XOR2_X1 U925 ( .A(n1267), .B(KEYINPUT52), .Z(n1265) );
OR2_X1 U926 ( .A1(n1215), .A2(G125), .ZN(n1267) );
NAND4_X1 U927 ( .A1(n1236), .A2(n1078), .A3(n1073), .A4(n1263), .ZN(n1215) );
NAND2_X1 U928 ( .A1(n1268), .A2(n1269), .ZN(n1263) );
NAND4_X1 U929 ( .A1(n1270), .A2(G953), .A3(G902), .A4(n1054), .ZN(n1269) );
XNOR2_X1 U930 ( .A(G900), .B(KEYINPUT36), .ZN(n1270) );
XNOR2_X1 U931 ( .A(n1230), .B(n1271), .ZN(G24) );
NOR2_X1 U932 ( .A1(KEYINPUT59), .A2(n1272), .ZN(n1271) );
NAND4_X1 U933 ( .A1(n1251), .A2(n1273), .A3(n1058), .A4(n1252), .ZN(n1230) );
NAND2_X1 U934 ( .A1(n1274), .A2(n1275), .ZN(n1058) );
NAND2_X1 U935 ( .A1(n1072), .A2(n1276), .ZN(n1275) );
NAND3_X1 U936 ( .A1(n1277), .A2(n1278), .A3(KEYINPUT9), .ZN(n1274) );
XNOR2_X1 U937 ( .A(G119), .B(n1235), .ZN(G21) );
NAND3_X1 U938 ( .A1(n1074), .A2(n1248), .A3(n1273), .ZN(n1235) );
XNOR2_X1 U939 ( .A(G116), .B(n1234), .ZN(G18) );
NAND2_X1 U940 ( .A1(n1279), .A2(n1077), .ZN(n1234) );
NOR2_X1 U941 ( .A1(n1251), .A2(n1280), .ZN(n1077) );
INV_X1 U942 ( .A(n1252), .ZN(n1280) );
XOR2_X1 U943 ( .A(n1281), .B(n1282), .Z(G15) );
NAND2_X1 U944 ( .A1(n1279), .A2(n1078), .ZN(n1282) );
INV_X1 U945 ( .A(n1085), .ZN(n1078) );
NAND2_X1 U946 ( .A1(n1283), .A2(n1251), .ZN(n1085) );
XNOR2_X1 U947 ( .A(n1252), .B(KEYINPUT61), .ZN(n1283) );
AND2_X1 U948 ( .A1(n1273), .A2(n1072), .ZN(n1279) );
NOR2_X1 U949 ( .A1(n1094), .A2(n1277), .ZN(n1072) );
AND2_X1 U950 ( .A1(n1236), .A2(n1238), .ZN(n1273) );
AND2_X1 U951 ( .A1(n1264), .A2(n1061), .ZN(n1236) );
NAND2_X1 U952 ( .A1(KEYINPUT6), .A2(G113), .ZN(n1281) );
XNOR2_X1 U953 ( .A(G110), .B(n1233), .ZN(G12) );
NAND3_X1 U954 ( .A1(n1228), .A2(n1073), .A3(n1074), .ZN(n1233) );
NOR2_X1 U955 ( .A1(n1252), .A2(n1251), .ZN(n1074) );
XOR2_X1 U956 ( .A(n1161), .B(n1284), .Z(n1251) );
NOR2_X1 U957 ( .A1(KEYINPUT46), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U958 ( .A(n1099), .B(KEYINPUT60), .ZN(n1285) );
NOR2_X1 U959 ( .A1(n1162), .A2(G902), .ZN(n1099) );
XNOR2_X1 U960 ( .A(n1286), .B(n1287), .ZN(n1162) );
XOR2_X1 U961 ( .A(n1288), .B(n1289), .Z(n1287) );
XNOR2_X1 U962 ( .A(n1122), .B(n1290), .ZN(n1289) );
NOR2_X1 U963 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XOR2_X1 U964 ( .A(n1293), .B(KEYINPUT62), .Z(n1292) );
OR3_X1 U965 ( .A1(n1294), .A2(G104), .A3(n1295), .ZN(n1293) );
NOR2_X1 U966 ( .A1(n1296), .A2(n1297), .ZN(n1291) );
NOR2_X1 U967 ( .A1(n1294), .A2(n1295), .ZN(n1296) );
XNOR2_X1 U968 ( .A(n1298), .B(KEYINPUT31), .ZN(n1295) );
NAND2_X1 U969 ( .A1(G122), .A2(n1299), .ZN(n1298) );
NOR2_X1 U970 ( .A1(n1299), .A2(G122), .ZN(n1294) );
INV_X1 U971 ( .A(G131), .ZN(n1122) );
NOR2_X1 U972 ( .A1(n1300), .A2(n1301), .ZN(n1288) );
XOR2_X1 U973 ( .A(KEYINPUT1), .B(n1302), .Z(n1301) );
NOR2_X1 U974 ( .A1(n1303), .A2(G143), .ZN(n1302) );
NOR3_X1 U975 ( .A1(n1304), .A2(G953), .A3(G237), .ZN(n1303) );
NOR4_X1 U976 ( .A1(G953), .A2(G237), .A3(n1304), .A4(n1305), .ZN(n1300) );
XNOR2_X1 U977 ( .A(n1306), .B(n1307), .ZN(n1286) );
INV_X1 U978 ( .A(G475), .ZN(n1161) );
XOR2_X1 U979 ( .A(n1104), .B(n1308), .Z(n1252) );
NOR2_X1 U980 ( .A1(KEYINPUT5), .A2(n1106), .ZN(n1308) );
INV_X1 U981 ( .A(G478), .ZN(n1106) );
NOR2_X1 U982 ( .A1(n1155), .A2(G902), .ZN(n1104) );
INV_X1 U983 ( .A(n1153), .ZN(n1155) );
XNOR2_X1 U984 ( .A(n1309), .B(n1310), .ZN(n1153) );
XNOR2_X1 U985 ( .A(n1311), .B(n1312), .ZN(n1310) );
XNOR2_X1 U986 ( .A(G134), .B(n1272), .ZN(n1312) );
INV_X1 U987 ( .A(G122), .ZN(n1272) );
XOR2_X1 U988 ( .A(n1313), .B(n1314), .Z(n1309) );
AND2_X1 U989 ( .A1(n1315), .A2(G217), .ZN(n1314) );
XNOR2_X1 U990 ( .A(G107), .B(n1316), .ZN(n1313) );
NOR2_X1 U991 ( .A1(KEYINPUT55), .A2(n1317), .ZN(n1316) );
NAND2_X1 U992 ( .A1(n1318), .A2(n1319), .ZN(n1073) );
NAND2_X1 U993 ( .A1(n1248), .A2(n1276), .ZN(n1319) );
INV_X1 U994 ( .A(KEYINPUT9), .ZN(n1276) );
NOR2_X1 U995 ( .A1(n1278), .A2(n1277), .ZN(n1248) );
INV_X1 U996 ( .A(n1094), .ZN(n1278) );
NAND3_X1 U997 ( .A1(n1277), .A2(n1094), .A3(KEYINPUT9), .ZN(n1318) );
XOR2_X1 U998 ( .A(n1320), .B(n1148), .Z(n1094) );
NAND2_X1 U999 ( .A1(G217), .A2(n1321), .ZN(n1148) );
NAND2_X1 U1000 ( .A1(n1146), .A2(n1213), .ZN(n1320) );
XNOR2_X1 U1001 ( .A(n1322), .B(n1323), .ZN(n1146) );
XNOR2_X1 U1002 ( .A(n1324), .B(n1325), .ZN(n1323) );
XOR2_X1 U1003 ( .A(n1326), .B(n1327), .Z(n1325) );
NAND2_X1 U1004 ( .A1(n1315), .A2(G221), .ZN(n1327) );
AND2_X1 U1005 ( .A1(G234), .A2(n1114), .ZN(n1315) );
NAND2_X1 U1006 ( .A1(KEYINPUT58), .A2(n1328), .ZN(n1326) );
INV_X1 U1007 ( .A(n1121), .ZN(n1324) );
XOR2_X1 U1008 ( .A(n1329), .B(n1306), .Z(n1121) );
XNOR2_X1 U1009 ( .A(G125), .B(n1256), .ZN(n1306) );
INV_X1 U1010 ( .A(G140), .ZN(n1256) );
XOR2_X1 U1011 ( .A(n1330), .B(n1331), .Z(n1322) );
NOR2_X1 U1012 ( .A1(KEYINPUT54), .A2(n1307), .ZN(n1331) );
XNOR2_X1 U1013 ( .A(G110), .B(G128), .ZN(n1330) );
AND3_X1 U1014 ( .A1(n1332), .A2(n1333), .A3(n1101), .ZN(n1277) );
NAND2_X1 U1015 ( .A1(n1334), .A2(n1186), .ZN(n1101) );
INV_X1 U1016 ( .A(G472), .ZN(n1186) );
OR2_X1 U1017 ( .A1(n1089), .A2(KEYINPUT11), .ZN(n1333) );
NAND2_X1 U1018 ( .A1(G472), .A2(n1335), .ZN(n1089) );
NAND2_X1 U1019 ( .A1(KEYINPUT11), .A2(n1334), .ZN(n1332) );
INV_X1 U1020 ( .A(n1335), .ZN(n1334) );
NAND2_X1 U1021 ( .A1(n1336), .A2(n1213), .ZN(n1335) );
XOR2_X1 U1022 ( .A(n1337), .B(n1338), .Z(n1336) );
XNOR2_X1 U1023 ( .A(n1177), .B(n1180), .ZN(n1338) );
XNOR2_X1 U1024 ( .A(n1173), .B(n1339), .ZN(n1337) );
XNOR2_X1 U1025 ( .A(n1187), .B(n1167), .ZN(n1339) );
NOR3_X1 U1026 ( .A1(G237), .A2(G953), .A3(n1212), .ZN(n1167) );
INV_X1 U1027 ( .A(G101), .ZN(n1187) );
XNOR2_X1 U1028 ( .A(n1340), .B(n1341), .ZN(n1173) );
XNOR2_X1 U1029 ( .A(KEYINPUT56), .B(n1311), .ZN(n1341) );
XNOR2_X1 U1030 ( .A(n1342), .B(n1299), .ZN(n1340) );
INV_X1 U1031 ( .A(G113), .ZN(n1299) );
NAND2_X1 U1032 ( .A1(KEYINPUT57), .A2(n1328), .ZN(n1342) );
AND3_X1 U1033 ( .A1(n1261), .A2(n1238), .A3(n1264), .ZN(n1228) );
NOR3_X1 U1034 ( .A1(n1060), .A2(n1103), .A3(n1080), .ZN(n1264) );
XOR2_X1 U1035 ( .A(n1093), .B(KEYINPUT44), .Z(n1080) );
XNOR2_X1 U1036 ( .A(n1343), .B(n1344), .ZN(n1093) );
NOR2_X1 U1037 ( .A1(n1212), .A2(n1345), .ZN(n1344) );
XOR2_X1 U1038 ( .A(KEYINPUT30), .B(n1346), .Z(n1345) );
INV_X1 U1039 ( .A(G210), .ZN(n1212) );
NAND2_X1 U1040 ( .A1(n1347), .A2(n1213), .ZN(n1343) );
XOR2_X1 U1041 ( .A(n1348), .B(n1349), .Z(n1347) );
NAND2_X1 U1042 ( .A1(KEYINPUT18), .A2(n1207), .ZN(n1349) );
XNOR2_X1 U1043 ( .A(n1350), .B(n1136), .ZN(n1207) );
XNOR2_X1 U1044 ( .A(n1200), .B(G122), .ZN(n1136) );
NAND2_X1 U1045 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
NAND2_X1 U1046 ( .A1(n1134), .A2(n1137), .ZN(n1352) );
XOR2_X1 U1047 ( .A(n1353), .B(KEYINPUT7), .Z(n1351) );
OR2_X1 U1048 ( .A1(n1137), .A2(n1134), .ZN(n1353) );
XOR2_X1 U1049 ( .A(n1354), .B(G113), .Z(n1134) );
NAND3_X1 U1050 ( .A1(n1355), .A2(n1356), .A3(n1357), .ZN(n1354) );
NAND2_X1 U1051 ( .A1(G116), .A2(n1328), .ZN(n1357) );
NAND2_X1 U1052 ( .A1(KEYINPUT51), .A2(n1358), .ZN(n1356) );
NAND2_X1 U1053 ( .A1(n1359), .A2(n1311), .ZN(n1358) );
INV_X1 U1054 ( .A(G116), .ZN(n1311) );
XNOR2_X1 U1055 ( .A(KEYINPUT12), .B(n1328), .ZN(n1359) );
NAND2_X1 U1056 ( .A1(n1360), .A2(n1361), .ZN(n1355) );
INV_X1 U1057 ( .A(KEYINPUT51), .ZN(n1361) );
NAND2_X1 U1058 ( .A1(n1362), .A2(n1363), .ZN(n1360) );
NAND2_X1 U1059 ( .A1(KEYINPUT12), .A2(n1328), .ZN(n1363) );
OR3_X1 U1060 ( .A1(G116), .A2(KEYINPUT12), .A3(n1328), .ZN(n1362) );
INV_X1 U1061 ( .A(G119), .ZN(n1328) );
XOR2_X1 U1062 ( .A(G101), .B(n1364), .Z(n1137) );
NAND3_X1 U1063 ( .A1(n1365), .A2(n1366), .A3(n1367), .ZN(n1348) );
NAND2_X1 U1064 ( .A1(n1210), .A2(n1368), .ZN(n1367) );
INV_X1 U1065 ( .A(KEYINPUT22), .ZN(n1368) );
NAND3_X1 U1066 ( .A1(KEYINPUT22), .A2(n1369), .A3(n1209), .ZN(n1366) );
OR2_X1 U1067 ( .A1(n1209), .A2(n1369), .ZN(n1365) );
NOR2_X1 U1068 ( .A1(KEYINPUT34), .A2(n1210), .ZN(n1369) );
NAND2_X1 U1069 ( .A1(G224), .A2(n1114), .ZN(n1210) );
XOR2_X1 U1070 ( .A(G125), .B(n1181), .Z(n1209) );
INV_X1 U1071 ( .A(n1180), .ZN(n1181) );
XNOR2_X1 U1072 ( .A(n1317), .B(n1307), .ZN(n1180) );
XOR2_X1 U1073 ( .A(G128), .B(n1305), .Z(n1317) );
NOR2_X1 U1074 ( .A1(n1304), .A2(n1346), .ZN(n1103) );
NOR2_X1 U1075 ( .A1(G902), .A2(G237), .ZN(n1346) );
INV_X1 U1076 ( .A(G214), .ZN(n1304) );
INV_X1 U1077 ( .A(n1102), .ZN(n1060) );
NAND2_X1 U1078 ( .A1(G221), .A2(n1321), .ZN(n1102) );
NAND2_X1 U1079 ( .A1(G234), .A2(n1213), .ZN(n1321) );
NAND2_X1 U1080 ( .A1(n1268), .A2(n1370), .ZN(n1238) );
NAND4_X1 U1081 ( .A1(G953), .A2(G902), .A3(n1054), .A4(n1371), .ZN(n1370) );
INV_X1 U1082 ( .A(G898), .ZN(n1371) );
NAND3_X1 U1083 ( .A1(n1054), .A2(n1114), .A3(G952), .ZN(n1268) );
NAND2_X1 U1084 ( .A1(G237), .A2(G234), .ZN(n1054) );
INV_X1 U1085 ( .A(n1061), .ZN(n1261) );
XNOR2_X1 U1086 ( .A(n1098), .B(n1372), .ZN(n1061) );
XNOR2_X1 U1087 ( .A(KEYINPUT38), .B(n1096), .ZN(n1372) );
INV_X1 U1088 ( .A(G469), .ZN(n1096) );
NAND2_X1 U1089 ( .A1(n1373), .A2(n1213), .ZN(n1098) );
INV_X1 U1090 ( .A(G902), .ZN(n1213) );
XOR2_X1 U1091 ( .A(n1374), .B(n1375), .Z(n1373) );
XNOR2_X1 U1092 ( .A(n1196), .B(n1177), .ZN(n1375) );
INV_X1 U1093 ( .A(n1178), .ZN(n1177) );
XOR2_X1 U1094 ( .A(n1376), .B(n1377), .Z(n1178) );
INV_X1 U1095 ( .A(n1329), .ZN(n1377) );
XOR2_X1 U1096 ( .A(G137), .B(KEYINPUT20), .Z(n1329) );
XNOR2_X1 U1097 ( .A(G131), .B(G134), .ZN(n1376) );
XNOR2_X1 U1098 ( .A(G140), .B(KEYINPUT39), .ZN(n1196) );
XOR2_X1 U1099 ( .A(n1378), .B(n1201), .Z(n1374) );
AND2_X1 U1100 ( .A1(G227), .A2(n1114), .ZN(n1201) );
INV_X1 U1101 ( .A(G953), .ZN(n1114) );
XNOR2_X1 U1102 ( .A(n1379), .B(n1200), .ZN(n1378) );
INV_X1 U1103 ( .A(G110), .ZN(n1200) );
NAND2_X1 U1104 ( .A1(KEYINPUT32), .A2(n1191), .ZN(n1379) );
XOR2_X1 U1105 ( .A(n1364), .B(n1380), .Z(n1191) );
XOR2_X1 U1106 ( .A(n1381), .B(n1125), .Z(n1380) );
XNOR2_X1 U1107 ( .A(G128), .B(n1382), .ZN(n1125) );
NOR2_X1 U1108 ( .A1(KEYINPUT13), .A2(n1383), .ZN(n1382) );
XOR2_X1 U1109 ( .A(n1307), .B(n1384), .Z(n1383) );
XNOR2_X1 U1110 ( .A(KEYINPUT45), .B(n1305), .ZN(n1384) );
INV_X1 U1111 ( .A(G143), .ZN(n1305) );
XNOR2_X1 U1112 ( .A(n1246), .B(KEYINPUT4), .ZN(n1307) );
INV_X1 U1113 ( .A(G146), .ZN(n1246) );
NAND2_X1 U1114 ( .A1(n1385), .A2(KEYINPUT21), .ZN(n1381) );
XNOR2_X1 U1115 ( .A(G101), .B(KEYINPUT26), .ZN(n1385) );
XNOR2_X1 U1116 ( .A(G107), .B(n1297), .ZN(n1364) );
INV_X1 U1117 ( .A(G104), .ZN(n1297) );
endmodule


