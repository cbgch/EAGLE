//Key = 1001110001010101011100100110001101100110010100111011011100010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;

XNOR2_X1 U745 ( .A(G107), .B(n1025), .ZN(G9) );
NOR2_X1 U746 ( .A1(n1026), .A2(n1027), .ZN(G75) );
AND3_X1 U747 ( .A1(n1028), .A2(G952), .A3(n1029), .ZN(n1027) );
AND3_X1 U748 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1028) );
NAND2_X1 U749 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U750 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND4_X1 U751 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1036) );
NAND2_X1 U752 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U753 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
XNOR2_X1 U754 ( .A(KEYINPUT26), .B(n1045), .ZN(n1043) );
NAND3_X1 U755 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1041) );
OR2_X1 U756 ( .A1(n1049), .A2(n1045), .ZN(n1047) );
OR3_X1 U757 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1046) );
NAND3_X1 U758 ( .A1(n1045), .A2(n1053), .A3(n1054), .ZN(n1035) );
NAND2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NAND2_X1 U760 ( .A1(n1038), .A2(n1057), .ZN(n1056) );
NAND2_X1 U761 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U762 ( .A1(n1037), .A2(n1060), .ZN(n1059) );
OR2_X1 U763 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U764 ( .A1(n1063), .A2(n1039), .ZN(n1058) );
NAND2_X1 U765 ( .A1(n1039), .A2(n1064), .ZN(n1055) );
INV_X1 U766 ( .A(n1065), .ZN(n1033) );
NOR3_X1 U767 ( .A1(n1066), .A2(G953), .A3(n1067), .ZN(n1026) );
INV_X1 U768 ( .A(n1030), .ZN(n1067) );
NAND4_X1 U769 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1030) );
NOR4_X1 U770 ( .A1(n1063), .A2(n1052), .A3(n1072), .A4(n1073), .ZN(n1071) );
XOR2_X1 U771 ( .A(n1074), .B(n1075), .Z(n1073) );
NOR2_X1 U772 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XNOR2_X1 U773 ( .A(KEYINPUT52), .B(KEYINPUT19), .ZN(n1077) );
XOR2_X1 U774 ( .A(n1078), .B(n1079), .Z(n1072) );
NAND2_X1 U775 ( .A1(KEYINPUT15), .A2(n1080), .ZN(n1078) );
NOR2_X1 U776 ( .A1(n1081), .A2(n1082), .ZN(n1070) );
XOR2_X1 U777 ( .A(n1083), .B(n1084), .Z(n1082) );
NAND2_X1 U778 ( .A1(KEYINPUT53), .A2(G475), .ZN(n1084) );
XOR2_X1 U779 ( .A(n1038), .B(KEYINPUT57), .Z(n1069) );
XOR2_X1 U780 ( .A(n1085), .B(G469), .Z(n1068) );
XOR2_X1 U781 ( .A(KEYINPUT62), .B(G952), .Z(n1066) );
XOR2_X1 U782 ( .A(n1086), .B(n1087), .Z(G72) );
XOR2_X1 U783 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U784 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NAND2_X1 U786 ( .A1(n1094), .A2(n1095), .ZN(n1088) );
NAND2_X1 U787 ( .A1(G953), .A2(n1093), .ZN(n1095) );
XOR2_X1 U788 ( .A(n1096), .B(n1097), .Z(n1094) );
XNOR2_X1 U789 ( .A(n1098), .B(KEYINPUT32), .ZN(n1097) );
NAND2_X1 U790 ( .A1(n1099), .A2(KEYINPUT25), .ZN(n1098) );
XNOR2_X1 U791 ( .A(G128), .B(n1100), .ZN(n1099) );
XNOR2_X1 U792 ( .A(n1101), .B(n1102), .ZN(n1096) );
NAND2_X1 U793 ( .A1(n1031), .A2(n1103), .ZN(n1086) );
NAND2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(G69) );
NAND3_X1 U795 ( .A1(n1106), .A2(n1107), .A3(KEYINPUT18), .ZN(n1105) );
NAND2_X1 U796 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND3_X1 U797 ( .A1(n1109), .A2(n1110), .A3(n1108), .ZN(n1104) );
INV_X1 U798 ( .A(n1091), .ZN(n1108) );
XOR2_X1 U799 ( .A(G953), .B(KEYINPUT5), .Z(n1091) );
NAND2_X1 U800 ( .A1(KEYINPUT18), .A2(n1106), .ZN(n1110) );
XOR2_X1 U801 ( .A(n1111), .B(n1112), .Z(n1106) );
NAND4_X1 U802 ( .A1(n1113), .A2(KEYINPUT9), .A3(n1114), .A4(n1115), .ZN(n1112) );
NAND2_X1 U803 ( .A1(G953), .A2(n1116), .ZN(n1114) );
NAND2_X1 U804 ( .A1(n1117), .A2(n1031), .ZN(n1111) );
NAND2_X1 U805 ( .A1(G898), .A2(G224), .ZN(n1109) );
NOR3_X1 U806 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(G66) );
NOR3_X1 U807 ( .A1(n1121), .A2(G953), .A3(G952), .ZN(n1120) );
AND2_X1 U808 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
INV_X1 U809 ( .A(KEYINPUT21), .ZN(n1121) );
XOR2_X1 U810 ( .A(n1123), .B(n1124), .Z(n1118) );
NAND2_X1 U811 ( .A1(n1125), .A2(n1076), .ZN(n1123) );
INV_X1 U812 ( .A(n1126), .ZN(n1076) );
NOR2_X1 U813 ( .A1(n1122), .A2(n1127), .ZN(G63) );
XOR2_X1 U814 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND2_X1 U815 ( .A1(KEYINPUT33), .A2(n1130), .ZN(n1129) );
NAND2_X1 U816 ( .A1(n1125), .A2(G478), .ZN(n1128) );
NOR2_X1 U817 ( .A1(n1122), .A2(n1131), .ZN(G60) );
XOR2_X1 U818 ( .A(n1132), .B(n1133), .Z(n1131) );
AND2_X1 U819 ( .A1(G475), .A2(n1125), .ZN(n1133) );
NAND2_X1 U820 ( .A1(KEYINPUT31), .A2(n1134), .ZN(n1132) );
XOR2_X1 U821 ( .A(G104), .B(n1135), .Z(G6) );
NOR2_X1 U822 ( .A1(n1122), .A2(n1136), .ZN(G57) );
XOR2_X1 U823 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U824 ( .A1(KEYINPUT43), .A2(n1139), .ZN(n1137) );
XOR2_X1 U825 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U826 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND4_X1 U827 ( .A1(KEYINPUT17), .A2(G472), .A3(n1144), .A4(n1145), .ZN(n1142) );
OR2_X1 U828 ( .A1(n1125), .A2(KEYINPUT23), .ZN(n1145) );
NAND2_X1 U829 ( .A1(KEYINPUT23), .A2(n1146), .ZN(n1144) );
NAND2_X1 U830 ( .A1(n1029), .A2(G902), .ZN(n1146) );
XNOR2_X1 U831 ( .A(n1147), .B(KEYINPUT46), .ZN(n1140) );
NAND2_X1 U832 ( .A1(KEYINPUT11), .A2(n1101), .ZN(n1147) );
NOR2_X1 U833 ( .A1(n1122), .A2(n1148), .ZN(G54) );
XOR2_X1 U834 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U835 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U836 ( .A1(n1125), .A2(G469), .ZN(n1151) );
XOR2_X1 U837 ( .A(n1153), .B(n1154), .Z(n1149) );
NOR2_X1 U838 ( .A1(KEYINPUT28), .A2(n1155), .ZN(n1154) );
NOR2_X1 U839 ( .A1(n1156), .A2(n1157), .ZN(n1153) );
XOR2_X1 U840 ( .A(n1158), .B(KEYINPUT41), .Z(n1157) );
NAND2_X1 U841 ( .A1(G110), .A2(n1159), .ZN(n1158) );
NOR2_X1 U842 ( .A1(G110), .A2(n1159), .ZN(n1156) );
NOR2_X1 U843 ( .A1(n1122), .A2(n1160), .ZN(G51) );
XOR2_X1 U844 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U845 ( .A(n1163), .B(n1164), .Z(n1162) );
NAND2_X1 U846 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
OR2_X1 U847 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND3_X1 U848 ( .A1(n1125), .A2(n1169), .A3(KEYINPUT63), .ZN(n1161) );
NOR2_X1 U849 ( .A1(n1170), .A2(n1029), .ZN(n1125) );
NOR2_X1 U850 ( .A1(n1103), .A2(n1117), .ZN(n1029) );
NAND4_X1 U851 ( .A1(n1171), .A2(n1025), .A3(n1172), .A4(n1173), .ZN(n1117) );
NOR4_X1 U852 ( .A1(n1174), .A2(n1175), .A3(n1135), .A4(n1176), .ZN(n1173) );
NOR2_X1 U853 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR3_X1 U854 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1177) );
NOR2_X1 U855 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
XNOR2_X1 U856 ( .A(n1061), .B(KEYINPUT42), .ZN(n1182) );
INV_X1 U857 ( .A(n1184), .ZN(n1180) );
NOR2_X1 U858 ( .A1(KEYINPUT6), .A2(n1185), .ZN(n1179) );
AND3_X1 U859 ( .A1(n1039), .A2(n1186), .A3(n1051), .ZN(n1135) );
NOR2_X1 U860 ( .A1(n1187), .A2(n1188), .ZN(n1175) );
XOR2_X1 U861 ( .A(n1189), .B(KEYINPUT49), .Z(n1188) );
NOR4_X1 U862 ( .A1(n1064), .A2(n1190), .A3(n1191), .A4(n1185), .ZN(n1174) );
INV_X1 U863 ( .A(KEYINPUT6), .ZN(n1190) );
NAND3_X1 U864 ( .A1(n1050), .A2(n1186), .A3(n1039), .ZN(n1025) );
NAND4_X1 U865 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1103) );
NOR4_X1 U866 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1195) );
NAND2_X1 U867 ( .A1(n1200), .A2(n1201), .ZN(n1194) );
NAND2_X1 U868 ( .A1(n1185), .A2(n1184), .ZN(n1201) );
NOR2_X1 U869 ( .A1(n1031), .A2(G952), .ZN(n1122) );
XNOR2_X1 U870 ( .A(G146), .B(n1192), .ZN(G48) );
NAND3_X1 U871 ( .A1(n1051), .A2(n1044), .A3(n1202), .ZN(n1192) );
XNOR2_X1 U872 ( .A(G143), .B(n1193), .ZN(G45) );
NAND4_X1 U873 ( .A1(n1064), .A2(n1203), .A3(n1061), .A4(n1204), .ZN(n1193) );
AND3_X1 U874 ( .A1(n1044), .A2(n1205), .A3(n1206), .ZN(n1204) );
NAND2_X1 U875 ( .A1(n1207), .A2(n1208), .ZN(G42) );
NAND2_X1 U876 ( .A1(n1199), .A2(n1159), .ZN(n1208) );
XOR2_X1 U877 ( .A(KEYINPUT54), .B(n1209), .Z(n1207) );
NOR2_X1 U878 ( .A1(n1199), .A2(n1159), .ZN(n1209) );
AND3_X1 U879 ( .A1(n1051), .A2(n1062), .A3(n1200), .ZN(n1199) );
INV_X1 U880 ( .A(n1210), .ZN(n1200) );
XNOR2_X1 U881 ( .A(n1211), .B(n1212), .ZN(G39) );
NOR2_X1 U882 ( .A1(n1210), .A2(n1184), .ZN(n1212) );
XOR2_X1 U883 ( .A(G134), .B(n1213), .Z(G36) );
NOR2_X1 U884 ( .A1(n1210), .A2(n1185), .ZN(n1213) );
XNOR2_X1 U885 ( .A(n1214), .B(n1198), .ZN(G33) );
NOR3_X1 U886 ( .A1(n1210), .A2(n1183), .A3(n1215), .ZN(n1198) );
NAND4_X1 U887 ( .A1(n1037), .A2(n1038), .A3(n1044), .A4(n1205), .ZN(n1210) );
XNOR2_X1 U888 ( .A(n1063), .B(KEYINPUT45), .ZN(n1037) );
XNOR2_X1 U889 ( .A(n1216), .B(n1197), .ZN(G30) );
AND3_X1 U890 ( .A1(n1217), .A2(n1050), .A3(n1202), .ZN(n1197) );
AND4_X1 U891 ( .A1(n1064), .A2(n1205), .A3(n1218), .A4(n1219), .ZN(n1202) );
NAND2_X1 U892 ( .A1(KEYINPUT29), .A2(n1215), .ZN(n1219) );
NAND2_X1 U893 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
INV_X1 U894 ( .A(KEYINPUT29), .ZN(n1221) );
NAND2_X1 U895 ( .A1(n1222), .A2(n1081), .ZN(n1220) );
XOR2_X1 U896 ( .A(G101), .B(n1223), .Z(G3) );
NOR2_X1 U897 ( .A1(n1187), .A2(n1189), .ZN(n1223) );
NAND4_X1 U898 ( .A1(n1217), .A2(n1061), .A3(n1045), .A4(n1224), .ZN(n1189) );
XOR2_X1 U899 ( .A(n1196), .B(n1225), .Z(G27) );
NOR2_X1 U900 ( .A1(KEYINPUT36), .A2(n1226), .ZN(n1225) );
XOR2_X1 U901 ( .A(KEYINPUT47), .B(G125), .Z(n1226) );
AND4_X1 U902 ( .A1(n1051), .A2(n1062), .A3(n1227), .A4(n1064), .ZN(n1196) );
AND2_X1 U903 ( .A1(n1205), .A2(n1054), .ZN(n1227) );
NAND2_X1 U904 ( .A1(n1065), .A2(n1228), .ZN(n1205) );
NAND4_X1 U905 ( .A1(G953), .A2(G902), .A3(n1229), .A4(n1093), .ZN(n1228) );
INV_X1 U906 ( .A(G900), .ZN(n1093) );
XNOR2_X1 U907 ( .A(G122), .B(n1172), .ZN(G24) );
NAND4_X1 U908 ( .A1(n1230), .A2(n1039), .A3(n1203), .A4(n1206), .ZN(n1172) );
NOR2_X1 U909 ( .A1(n1081), .A2(n1222), .ZN(n1039) );
INV_X1 U910 ( .A(n1231), .ZN(n1222) );
XOR2_X1 U911 ( .A(n1232), .B(n1233), .Z(G21) );
NOR2_X1 U912 ( .A1(KEYINPUT2), .A2(n1234), .ZN(n1233) );
NOR3_X1 U913 ( .A1(n1184), .A2(n1235), .A3(n1236), .ZN(n1232) );
NOR2_X1 U914 ( .A1(KEYINPUT30), .A2(n1237), .ZN(n1236) );
NOR2_X1 U915 ( .A1(n1064), .A2(n1191), .ZN(n1237) );
AND2_X1 U916 ( .A1(n1178), .A2(KEYINPUT30), .ZN(n1235) );
NAND3_X1 U917 ( .A1(n1045), .A2(n1081), .A3(n1238), .ZN(n1184) );
XNOR2_X1 U918 ( .A(KEYINPUT29), .B(n1231), .ZN(n1238) );
NAND2_X1 U919 ( .A1(n1239), .A2(n1240), .ZN(G18) );
NAND2_X1 U920 ( .A1(KEYINPUT40), .A2(n1241), .ZN(n1240) );
XOR2_X1 U921 ( .A(n1242), .B(n1243), .Z(n1239) );
NOR2_X1 U922 ( .A1(n1178), .A2(n1185), .ZN(n1243) );
NAND2_X1 U923 ( .A1(n1061), .A2(n1050), .ZN(n1185) );
NOR2_X1 U924 ( .A1(n1244), .A2(n1206), .ZN(n1050) );
INV_X1 U925 ( .A(n1215), .ZN(n1061) );
OR2_X1 U926 ( .A1(n1241), .A2(KEYINPUT40), .ZN(n1242) );
XNOR2_X1 U927 ( .A(n1245), .B(n1246), .ZN(G15) );
NOR3_X1 U928 ( .A1(n1178), .A2(n1183), .A3(n1215), .ZN(n1246) );
NAND2_X1 U929 ( .A1(n1231), .A2(n1081), .ZN(n1215) );
INV_X1 U930 ( .A(n1230), .ZN(n1178) );
NOR2_X1 U931 ( .A1(n1191), .A2(n1187), .ZN(n1230) );
INV_X1 U932 ( .A(n1064), .ZN(n1187) );
NAND2_X1 U933 ( .A1(n1054), .A2(n1224), .ZN(n1191) );
XNOR2_X1 U934 ( .A(G110), .B(n1247), .ZN(G12) );
NOR2_X1 U935 ( .A1(n1248), .A2(KEYINPUT12), .ZN(n1247) );
INV_X1 U936 ( .A(n1171), .ZN(n1248) );
NAND3_X1 U937 ( .A1(n1186), .A2(n1045), .A3(n1062), .ZN(n1171) );
NOR2_X1 U938 ( .A1(n1231), .A2(n1081), .ZN(n1062) );
XNOR2_X1 U939 ( .A(n1249), .B(G472), .ZN(n1081) );
NAND2_X1 U940 ( .A1(n1250), .A2(n1170), .ZN(n1249) );
XOR2_X1 U941 ( .A(n1143), .B(n1251), .Z(n1250) );
XOR2_X1 U942 ( .A(n1252), .B(n1138), .Z(n1251) );
XOR2_X1 U943 ( .A(n1253), .B(n1254), .Z(n1138) );
NAND2_X1 U944 ( .A1(G210), .A2(n1255), .ZN(n1253) );
NAND2_X1 U945 ( .A1(KEYINPUT22), .A2(n1256), .ZN(n1252) );
XOR2_X1 U946 ( .A(n1257), .B(n1258), .Z(n1143) );
XNOR2_X1 U947 ( .A(n1259), .B(n1245), .ZN(n1257) );
XOR2_X1 U948 ( .A(n1260), .B(n1074), .Z(n1231) );
NAND2_X1 U949 ( .A1(n1124), .A2(n1170), .ZN(n1074) );
XNOR2_X1 U950 ( .A(n1261), .B(n1262), .ZN(n1124) );
XOR2_X1 U951 ( .A(n1263), .B(n1264), .Z(n1262) );
NAND2_X1 U952 ( .A1(G221), .A2(n1265), .ZN(n1264) );
NAND2_X1 U953 ( .A1(n1266), .A2(n1267), .ZN(n1263) );
NAND2_X1 U954 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XOR2_X1 U955 ( .A(n1270), .B(KEYINPUT24), .Z(n1266) );
OR2_X1 U956 ( .A1(n1268), .A2(n1269), .ZN(n1270) );
INV_X1 U957 ( .A(G146), .ZN(n1269) );
XOR2_X1 U958 ( .A(n1102), .B(KEYINPUT38), .Z(n1268) );
XNOR2_X1 U959 ( .A(G137), .B(n1271), .ZN(n1261) );
NOR2_X1 U960 ( .A1(KEYINPUT16), .A2(n1272), .ZN(n1271) );
XOR2_X1 U961 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U962 ( .A(n1234), .B(G110), .ZN(n1274) );
XNOR2_X1 U963 ( .A(KEYINPUT51), .B(n1216), .ZN(n1273) );
NAND2_X1 U964 ( .A1(KEYINPUT50), .A2(n1126), .ZN(n1260) );
NAND2_X1 U965 ( .A1(G217), .A2(n1275), .ZN(n1126) );
NAND2_X1 U966 ( .A1(n1276), .A2(n1277), .ZN(n1045) );
OR3_X1 U967 ( .A1(n1206), .A2(n1203), .A3(KEYINPUT56), .ZN(n1277) );
INV_X1 U968 ( .A(n1244), .ZN(n1203) );
NAND2_X1 U969 ( .A1(KEYINPUT56), .A2(n1051), .ZN(n1276) );
INV_X1 U970 ( .A(n1183), .ZN(n1051) );
NAND2_X1 U971 ( .A1(n1206), .A2(n1244), .ZN(n1183) );
NAND3_X1 U972 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1244) );
NAND2_X1 U973 ( .A1(n1079), .A2(n1281), .ZN(n1280) );
OR3_X1 U974 ( .A1(n1281), .A2(n1079), .A3(n1282), .ZN(n1279) );
NOR2_X1 U975 ( .A1(n1130), .A2(G902), .ZN(n1079) );
XOR2_X1 U976 ( .A(n1283), .B(n1284), .Z(n1130) );
XOR2_X1 U977 ( .A(n1285), .B(n1286), .Z(n1284) );
XOR2_X1 U978 ( .A(G143), .B(G134), .Z(n1286) );
XOR2_X1 U979 ( .A(KEYINPUT39), .B(KEYINPUT13), .Z(n1285) );
XOR2_X1 U980 ( .A(n1287), .B(n1288), .Z(n1283) );
XOR2_X1 U981 ( .A(n1289), .B(n1290), .Z(n1288) );
NOR2_X1 U982 ( .A1(G122), .A2(KEYINPUT44), .ZN(n1289) );
XNOR2_X1 U983 ( .A(n1291), .B(n1241), .ZN(n1287) );
INV_X1 U984 ( .A(G116), .ZN(n1241) );
NAND2_X1 U985 ( .A1(G217), .A2(n1265), .ZN(n1291) );
AND2_X1 U986 ( .A1(G234), .A2(n1031), .ZN(n1265) );
NAND2_X1 U987 ( .A1(KEYINPUT4), .A2(n1080), .ZN(n1281) );
INV_X1 U988 ( .A(G478), .ZN(n1080) );
NAND2_X1 U989 ( .A1(G478), .A2(n1282), .ZN(n1278) );
INV_X1 U990 ( .A(KEYINPUT0), .ZN(n1282) );
XNOR2_X1 U991 ( .A(n1083), .B(G475), .ZN(n1206) );
NAND2_X1 U992 ( .A1(n1134), .A2(n1170), .ZN(n1083) );
XNOR2_X1 U993 ( .A(n1292), .B(n1293), .ZN(n1134) );
XOR2_X1 U994 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U995 ( .A(n1245), .B(G104), .ZN(n1295) );
INV_X1 U996 ( .A(G113), .ZN(n1245) );
XNOR2_X1 U997 ( .A(n1214), .B(G122), .ZN(n1294) );
INV_X1 U998 ( .A(G131), .ZN(n1214) );
XOR2_X1 U999 ( .A(n1296), .B(n1102), .Z(n1292) );
XNOR2_X1 U1000 ( .A(G125), .B(n1159), .ZN(n1102) );
XNOR2_X1 U1001 ( .A(n1297), .B(n1298), .ZN(n1296) );
NAND2_X1 U1002 ( .A1(G214), .A2(n1255), .ZN(n1297) );
NOR2_X1 U1003 ( .A1(G953), .A2(G237), .ZN(n1255) );
AND3_X1 U1004 ( .A1(n1217), .A2(n1224), .A3(n1064), .ZN(n1186) );
NOR2_X1 U1005 ( .A1(n1038), .A2(n1063), .ZN(n1064) );
AND2_X1 U1006 ( .A1(G214), .A2(n1299), .ZN(n1063) );
XNOR2_X1 U1007 ( .A(n1169), .B(n1300), .ZN(n1038) );
NOR3_X1 U1008 ( .A1(n1301), .A2(G902), .A3(n1302), .ZN(n1300) );
NOR2_X1 U1009 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
XOR2_X1 U1010 ( .A(n1305), .B(KEYINPUT10), .Z(n1303) );
XOR2_X1 U1011 ( .A(n1306), .B(KEYINPUT55), .Z(n1301) );
NAND2_X1 U1012 ( .A1(n1305), .A2(n1304), .ZN(n1306) );
NAND3_X1 U1013 ( .A1(n1307), .A2(n1308), .A3(n1165), .ZN(n1304) );
NAND2_X1 U1014 ( .A1(n1168), .A2(n1167), .ZN(n1165) );
OR3_X1 U1015 ( .A1(n1167), .A2(n1168), .A3(KEYINPUT7), .ZN(n1308) );
AND2_X1 U1016 ( .A1(G224), .A2(n1031), .ZN(n1168) );
NAND2_X1 U1017 ( .A1(KEYINPUT7), .A2(n1167), .ZN(n1307) );
XNOR2_X1 U1018 ( .A(G125), .B(n1258), .ZN(n1167) );
XNOR2_X1 U1019 ( .A(n1216), .B(n1309), .ZN(n1258) );
NOR2_X1 U1020 ( .A1(KEYINPUT35), .A2(n1298), .ZN(n1309) );
XOR2_X1 U1021 ( .A(n1163), .B(KEYINPUT58), .Z(n1305) );
NAND3_X1 U1022 ( .A1(n1310), .A2(n1311), .A3(n1115), .ZN(n1163) );
NAND2_X1 U1023 ( .A1(n1312), .A2(n1313), .ZN(n1115) );
NAND2_X1 U1024 ( .A1(KEYINPUT61), .A2(n1314), .ZN(n1311) );
NAND3_X1 U1025 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n1314) );
INV_X1 U1026 ( .A(n1312), .ZN(n1317) );
NOR2_X1 U1027 ( .A1(n1318), .A2(n1319), .ZN(n1312) );
NAND2_X1 U1028 ( .A1(n1313), .A2(n1320), .ZN(n1316) );
NAND3_X1 U1029 ( .A1(n1321), .A2(n1318), .A3(n1319), .ZN(n1315) );
OR2_X1 U1030 ( .A1(n1113), .A2(KEYINPUT61), .ZN(n1310) );
AND2_X1 U1031 ( .A1(n1322), .A2(n1323), .ZN(n1113) );
NAND2_X1 U1032 ( .A1(n1324), .A2(n1319), .ZN(n1323) );
XNOR2_X1 U1033 ( .A(n1313), .B(n1318), .ZN(n1324) );
INV_X1 U1034 ( .A(n1321), .ZN(n1313) );
NAND3_X1 U1035 ( .A1(n1321), .A2(n1318), .A3(n1320), .ZN(n1322) );
INV_X1 U1036 ( .A(n1319), .ZN(n1320) );
XNOR2_X1 U1037 ( .A(G122), .B(G110), .ZN(n1319) );
XNOR2_X1 U1038 ( .A(G113), .B(n1325), .ZN(n1318) );
NOR2_X1 U1039 ( .A1(KEYINPUT27), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1040 ( .A(n1259), .B(KEYINPUT48), .Z(n1326) );
XNOR2_X1 U1041 ( .A(G116), .B(n1327), .ZN(n1259) );
XNOR2_X1 U1042 ( .A(KEYINPUT60), .B(n1234), .ZN(n1327) );
INV_X1 U1043 ( .A(G119), .ZN(n1234) );
XOR2_X1 U1044 ( .A(G107), .B(n1328), .Z(n1321) );
AND2_X1 U1045 ( .A1(G210), .A2(n1299), .ZN(n1169) );
OR2_X1 U1046 ( .A1(G902), .A2(G237), .ZN(n1299) );
NAND2_X1 U1047 ( .A1(n1065), .A2(n1329), .ZN(n1224) );
NAND4_X1 U1048 ( .A1(G953), .A2(G902), .A3(n1229), .A4(n1116), .ZN(n1329) );
INV_X1 U1049 ( .A(G898), .ZN(n1116) );
NAND3_X1 U1050 ( .A1(n1229), .A2(n1031), .A3(G952), .ZN(n1065) );
INV_X1 U1051 ( .A(G953), .ZN(n1031) );
NAND2_X1 U1052 ( .A1(G237), .A2(G234), .ZN(n1229) );
XNOR2_X1 U1053 ( .A(n1044), .B(KEYINPUT34), .ZN(n1217) );
NAND2_X1 U1054 ( .A1(n1330), .A2(n1331), .ZN(n1044) );
NAND2_X1 U1055 ( .A1(n1054), .A2(n1332), .ZN(n1331) );
AND2_X1 U1056 ( .A1(n1048), .A2(n1049), .ZN(n1054) );
OR3_X1 U1057 ( .A1(n1048), .A2(n1052), .A3(n1332), .ZN(n1330) );
INV_X1 U1058 ( .A(KEYINPUT59), .ZN(n1332) );
INV_X1 U1059 ( .A(n1049), .ZN(n1052) );
NAND2_X1 U1060 ( .A1(G221), .A2(n1275), .ZN(n1049) );
NAND2_X1 U1061 ( .A1(n1333), .A2(G234), .ZN(n1275) );
XNOR2_X1 U1062 ( .A(G902), .B(KEYINPUT14), .ZN(n1333) );
XNOR2_X1 U1063 ( .A(n1334), .B(G469), .ZN(n1048) );
NAND2_X1 U1064 ( .A1(KEYINPUT37), .A2(n1085), .ZN(n1334) );
NAND2_X1 U1065 ( .A1(n1335), .A2(n1170), .ZN(n1085) );
INV_X1 U1066 ( .A(G902), .ZN(n1170) );
XOR2_X1 U1067 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1068 ( .A(G110), .B(n1338), .Z(n1337) );
NOR2_X1 U1069 ( .A1(KEYINPUT8), .A2(n1159), .ZN(n1338) );
INV_X1 U1070 ( .A(G140), .ZN(n1159) );
XOR2_X1 U1071 ( .A(n1152), .B(n1155), .Z(n1336) );
XNOR2_X1 U1072 ( .A(n1256), .B(KEYINPUT20), .ZN(n1155) );
INV_X1 U1073 ( .A(n1101), .ZN(n1256) );
XOR2_X1 U1074 ( .A(G131), .B(n1339), .Z(n1101) );
XNOR2_X1 U1075 ( .A(n1211), .B(G134), .ZN(n1339) );
INV_X1 U1076 ( .A(G137), .ZN(n1211) );
XOR2_X1 U1077 ( .A(n1340), .B(n1341), .Z(n1152) );
XOR2_X1 U1078 ( .A(n1342), .B(n1290), .Z(n1341) );
XNOR2_X1 U1079 ( .A(G107), .B(n1216), .ZN(n1290) );
INV_X1 U1080 ( .A(G128), .ZN(n1216) );
NOR2_X1 U1081 ( .A1(G953), .A2(n1092), .ZN(n1342) );
INV_X1 U1082 ( .A(G227), .ZN(n1092) );
XNOR2_X1 U1083 ( .A(n1328), .B(n1100), .ZN(n1340) );
XNOR2_X1 U1084 ( .A(n1298), .B(KEYINPUT3), .ZN(n1100) );
XNOR2_X1 U1085 ( .A(G143), .B(G146), .ZN(n1298) );
XOR2_X1 U1086 ( .A(G104), .B(n1254), .Z(n1328) );
XOR2_X1 U1087 ( .A(G101), .B(KEYINPUT1), .Z(n1254) );
endmodule


