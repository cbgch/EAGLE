//Key = 1000110011011101110101111001100100011000010110000010001011010110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345;

XNOR2_X1 U736 ( .A(G107), .B(n1024), .ZN(G9) );
NOR2_X1 U737 ( .A1(n1025), .A2(n1026), .ZN(G75) );
NOR4_X1 U738 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
NAND3_X1 U739 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1027) );
NAND2_X1 U740 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U741 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U742 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NAND2_X1 U743 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NAND2_X1 U744 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
OR2_X1 U745 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U746 ( .A1(n1047), .A2(n1048), .ZN(n1041) );
OR2_X1 U747 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND3_X1 U748 ( .A1(n1047), .A2(n1051), .A3(n1043), .ZN(n1036) );
NAND3_X1 U749 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1051) );
NAND2_X1 U750 ( .A1(n1040), .A2(n1055), .ZN(n1054) );
NAND2_X1 U751 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U752 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
INV_X1 U753 ( .A(n1060), .ZN(n1056) );
NAND3_X1 U754 ( .A1(n1061), .A2(n1062), .A3(n1038), .ZN(n1052) );
NOR3_X1 U755 ( .A1(n1030), .A2(G952), .A3(n1063), .ZN(n1025) );
INV_X1 U756 ( .A(n1032), .ZN(n1063) );
NAND4_X1 U757 ( .A1(n1064), .A2(n1038), .A3(n1065), .A4(n1066), .ZN(n1032) );
NOR4_X1 U758 ( .A1(n1062), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1066) );
XNOR2_X1 U759 ( .A(n1070), .B(KEYINPUT17), .ZN(n1068) );
XOR2_X1 U760 ( .A(n1071), .B(n1072), .Z(n1067) );
NOR2_X1 U761 ( .A1(G475), .A2(KEYINPUT40), .ZN(n1072) );
XNOR2_X1 U762 ( .A(G478), .B(n1073), .ZN(n1065) );
NOR2_X1 U763 ( .A1(KEYINPUT10), .A2(n1074), .ZN(n1073) );
XNOR2_X1 U764 ( .A(n1075), .B(n1076), .ZN(n1064) );
NOR2_X1 U765 ( .A1(KEYINPUT14), .A2(n1077), .ZN(n1076) );
XOR2_X1 U766 ( .A(n1078), .B(n1079), .Z(G72) );
NOR2_X1 U767 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
AND2_X1 U768 ( .A1(G227), .A2(G900), .ZN(n1080) );
NAND2_X1 U769 ( .A1(n1082), .A2(n1083), .ZN(n1078) );
NAND2_X1 U770 ( .A1(n1084), .A2(n1081), .ZN(n1083) );
XOR2_X1 U771 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U772 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
XNOR2_X1 U773 ( .A(KEYINPUT41), .B(n1031), .ZN(n1088) );
INV_X1 U774 ( .A(n1089), .ZN(n1031) );
INV_X1 U775 ( .A(n1028), .ZN(n1087) );
NAND3_X1 U776 ( .A1(n1086), .A2(G900), .A3(G953), .ZN(n1082) );
XNOR2_X1 U777 ( .A(n1090), .B(n1091), .ZN(n1086) );
NOR2_X1 U778 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR2_X1 U779 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
INV_X1 U780 ( .A(n1096), .ZN(n1095) );
XOR2_X1 U781 ( .A(KEYINPUT32), .B(n1097), .Z(n1094) );
NOR2_X1 U782 ( .A1(n1096), .A2(n1098), .ZN(n1092) );
XOR2_X1 U783 ( .A(KEYINPUT13), .B(n1097), .Z(n1098) );
NOR2_X1 U784 ( .A1(KEYINPUT53), .A2(n1099), .ZN(n1097) );
XNOR2_X1 U785 ( .A(G131), .B(n1100), .ZN(n1099) );
NAND3_X1 U786 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1100) );
NAND2_X1 U787 ( .A1(KEYINPUT51), .A2(G134), .ZN(n1103) );
NAND3_X1 U788 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1102) );
INV_X1 U789 ( .A(KEYINPUT51), .ZN(n1105) );
OR2_X1 U790 ( .A1(n1106), .A2(n1104), .ZN(n1101) );
NOR2_X1 U791 ( .A1(G134), .A2(KEYINPUT7), .ZN(n1104) );
NAND2_X1 U792 ( .A1(n1107), .A2(n1108), .ZN(G69) );
NAND2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
INV_X1 U794 ( .A(n1111), .ZN(n1110) );
NAND2_X1 U795 ( .A1(n1112), .A2(n1113), .ZN(n1109) );
NAND2_X1 U796 ( .A1(G953), .A2(n1114), .ZN(n1113) );
NAND2_X1 U797 ( .A1(n1111), .A2(n1112), .ZN(n1107) );
AND2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1112) );
OR2_X1 U799 ( .A1(n1081), .A2(G224), .ZN(n1116) );
NAND2_X1 U800 ( .A1(n1029), .A2(n1081), .ZN(n1115) );
NOR3_X1 U801 ( .A1(KEYINPUT46), .A2(n1117), .A3(n1118), .ZN(n1111) );
XOR2_X1 U802 ( .A(n1119), .B(n1120), .Z(n1118) );
NOR2_X1 U803 ( .A1(KEYINPUT48), .A2(n1121), .ZN(n1120) );
XNOR2_X1 U804 ( .A(G122), .B(n1122), .ZN(n1121) );
INV_X1 U805 ( .A(G110), .ZN(n1122) );
NOR2_X1 U806 ( .A1(G898), .A2(n1081), .ZN(n1117) );
NOR2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(G66) );
XOR2_X1 U808 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND3_X1 U809 ( .A1(n1127), .A2(n1128), .A3(KEYINPUT31), .ZN(n1125) );
NOR2_X1 U810 ( .A1(n1123), .A2(n1129), .ZN(G63) );
XOR2_X1 U811 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U812 ( .A1(n1132), .A2(KEYINPUT25), .ZN(n1130) );
NOR2_X1 U813 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U814 ( .A1(n1123), .A2(n1135), .ZN(G60) );
XNOR2_X1 U815 ( .A(n1136), .B(n1137), .ZN(n1135) );
NOR3_X1 U816 ( .A1(n1134), .A2(KEYINPUT58), .A3(n1138), .ZN(n1137) );
XNOR2_X1 U817 ( .A(G104), .B(n1139), .ZN(G6) );
NOR2_X1 U818 ( .A1(n1123), .A2(n1140), .ZN(G57) );
XNOR2_X1 U819 ( .A(n1141), .B(n1142), .ZN(n1140) );
XNOR2_X1 U820 ( .A(n1143), .B(n1144), .ZN(n1142) );
NOR2_X1 U821 ( .A1(n1077), .A2(n1134), .ZN(n1143) );
INV_X1 U822 ( .A(G472), .ZN(n1077) );
NOR3_X1 U823 ( .A1(n1123), .A2(n1145), .A3(n1146), .ZN(G54) );
NOR2_X1 U824 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
INV_X1 U825 ( .A(n1149), .ZN(n1148) );
NOR2_X1 U826 ( .A1(n1150), .A2(n1151), .ZN(n1147) );
NOR3_X1 U827 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
AND2_X1 U828 ( .A1(n1152), .A2(n1153), .ZN(n1150) );
INV_X1 U829 ( .A(KEYINPUT62), .ZN(n1152) );
NOR2_X1 U830 ( .A1(n1155), .A2(n1149), .ZN(n1145) );
XNOR2_X1 U831 ( .A(n1156), .B(n1157), .ZN(n1149) );
XNOR2_X1 U832 ( .A(n1158), .B(n1159), .ZN(n1157) );
NOR2_X1 U833 ( .A1(KEYINPUT33), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U834 ( .A(n1090), .B(n1161), .ZN(n1156) );
NOR2_X1 U835 ( .A1(n1153), .A2(n1154), .ZN(n1155) );
INV_X1 U836 ( .A(KEYINPUT44), .ZN(n1154) );
NAND2_X1 U837 ( .A1(n1127), .A2(G469), .ZN(n1153) );
INV_X1 U838 ( .A(n1134), .ZN(n1127) );
NOR2_X1 U839 ( .A1(n1123), .A2(n1162), .ZN(G51) );
XOR2_X1 U840 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U841 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U842 ( .A1(n1167), .A2(n1134), .ZN(n1165) );
NAND2_X1 U843 ( .A1(G902), .A2(n1168), .ZN(n1134) );
OR3_X1 U844 ( .A1(n1029), .A2(n1089), .A3(n1028), .ZN(n1168) );
NAND4_X1 U845 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1028) );
NOR3_X1 U846 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1172) );
NAND2_X1 U847 ( .A1(n1176), .A2(n1040), .ZN(n1171) );
NAND3_X1 U848 ( .A1(n1177), .A2(n1178), .A3(n1045), .ZN(n1169) );
NAND2_X1 U849 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NAND2_X1 U850 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XNOR2_X1 U851 ( .A(KEYINPUT38), .B(n1183), .ZN(n1182) );
NAND2_X1 U852 ( .A1(n1040), .A2(n1050), .ZN(n1179) );
NAND4_X1 U853 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1029) );
AND4_X1 U854 ( .A1(n1024), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1187) );
NAND3_X1 U855 ( .A1(n1047), .A2(n1191), .A3(n1050), .ZN(n1024) );
AND2_X1 U856 ( .A1(n1192), .A2(n1139), .ZN(n1186) );
NAND3_X1 U857 ( .A1(n1191), .A2(n1049), .A3(n1047), .ZN(n1139) );
NAND4_X1 U858 ( .A1(n1193), .A2(n1181), .A3(n1194), .A4(n1047), .ZN(n1185) );
XNOR2_X1 U859 ( .A(n1195), .B(KEYINPUT45), .ZN(n1193) );
NAND2_X1 U860 ( .A1(n1196), .A2(n1197), .ZN(n1184) );
XNOR2_X1 U861 ( .A(KEYINPUT52), .B(n1198), .ZN(n1197) );
NOR2_X1 U862 ( .A1(n1199), .A2(n1200), .ZN(n1163) );
AND2_X1 U863 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NOR2_X1 U864 ( .A1(n1202), .A2(n1203), .ZN(n1199) );
XOR2_X1 U865 ( .A(n1201), .B(KEYINPUT37), .Z(n1203) );
XNOR2_X1 U866 ( .A(n1204), .B(n1205), .ZN(n1202) );
NOR2_X1 U867 ( .A1(G125), .A2(n1206), .ZN(n1205) );
XNOR2_X1 U868 ( .A(KEYINPUT9), .B(KEYINPUT39), .ZN(n1206) );
NOR2_X1 U869 ( .A1(n1081), .A2(G952), .ZN(n1123) );
XOR2_X1 U870 ( .A(G146), .B(n1173), .Z(G48) );
AND4_X1 U871 ( .A1(n1177), .A2(n1207), .A3(n1196), .A4(n1049), .ZN(n1173) );
XNOR2_X1 U872 ( .A(G143), .B(n1208), .ZN(G45) );
NAND4_X1 U873 ( .A1(n1181), .A2(n1045), .A3(n1177), .A4(n1196), .ZN(n1208) );
XNOR2_X1 U874 ( .A(G140), .B(n1209), .ZN(G42) );
NAND2_X1 U875 ( .A1(n1210), .A2(n1040), .ZN(n1209) );
XNOR2_X1 U876 ( .A(n1176), .B(KEYINPUT57), .ZN(n1210) );
AND3_X1 U877 ( .A1(n1177), .A2(n1049), .A3(n1046), .ZN(n1176) );
XOR2_X1 U878 ( .A(n1175), .B(n1211), .Z(G39) );
NOR2_X1 U879 ( .A1(KEYINPUT29), .A2(n1106), .ZN(n1211) );
AND4_X1 U880 ( .A1(n1040), .A2(n1177), .A3(n1043), .A4(n1207), .ZN(n1175) );
XNOR2_X1 U881 ( .A(G134), .B(n1212), .ZN(G36) );
NAND4_X1 U882 ( .A1(n1213), .A2(n1040), .A3(n1177), .A4(n1050), .ZN(n1212) );
XNOR2_X1 U883 ( .A(n1045), .B(KEYINPUT61), .ZN(n1213) );
XNOR2_X1 U884 ( .A(G131), .B(n1214), .ZN(G33) );
NAND2_X1 U885 ( .A1(KEYINPUT15), .A2(n1174), .ZN(n1214) );
AND4_X1 U886 ( .A1(n1040), .A2(n1045), .A3(n1177), .A4(n1049), .ZN(n1174) );
AND2_X1 U887 ( .A1(n1060), .A2(n1215), .ZN(n1177) );
AND2_X1 U888 ( .A1(n1061), .A2(n1216), .ZN(n1040) );
INV_X1 U889 ( .A(n1069), .ZN(n1061) );
XNOR2_X1 U890 ( .A(n1217), .B(n1218), .ZN(G30) );
NAND2_X1 U891 ( .A1(n1219), .A2(n1220), .ZN(n1217) );
OR3_X1 U892 ( .A1(n1221), .A2(n1222), .A3(KEYINPUT24), .ZN(n1220) );
NAND2_X1 U893 ( .A1(n1089), .A2(KEYINPUT24), .ZN(n1219) );
NOR2_X1 U894 ( .A1(n1221), .A2(n1223), .ZN(n1089) );
NAND4_X1 U895 ( .A1(n1207), .A2(n1050), .A3(n1196), .A4(n1215), .ZN(n1221) );
XNOR2_X1 U896 ( .A(G101), .B(n1192), .ZN(G3) );
NAND3_X1 U897 ( .A1(n1043), .A2(n1191), .A3(n1045), .ZN(n1192) );
XNOR2_X1 U898 ( .A(G125), .B(n1170), .ZN(G27) );
NAND4_X1 U899 ( .A1(n1194), .A2(n1046), .A3(n1049), .A4(n1215), .ZN(n1170) );
NAND2_X1 U900 ( .A1(n1224), .A2(n1225), .ZN(n1215) );
NAND2_X1 U901 ( .A1(n1226), .A2(n1227), .ZN(n1224) );
INV_X1 U902 ( .A(G900), .ZN(n1227) );
XOR2_X1 U903 ( .A(n1228), .B(n1229), .Z(G24) );
NOR2_X1 U904 ( .A1(G122), .A2(KEYINPUT55), .ZN(n1229) );
NAND4_X1 U905 ( .A1(n1181), .A2(n1194), .A3(n1047), .A4(n1230), .ZN(n1228) );
XNOR2_X1 U906 ( .A(KEYINPUT16), .B(n1231), .ZN(n1230) );
NOR2_X1 U907 ( .A1(n1232), .A2(n1070), .ZN(n1047) );
AND2_X1 U908 ( .A1(n1233), .A2(n1234), .ZN(n1181) );
XNOR2_X1 U909 ( .A(KEYINPUT8), .B(n1235), .ZN(n1233) );
XNOR2_X1 U910 ( .A(G119), .B(n1190), .ZN(G21) );
NAND4_X1 U911 ( .A1(n1194), .A2(n1043), .A3(n1207), .A4(n1231), .ZN(n1190) );
NOR2_X1 U912 ( .A1(n1236), .A2(n1237), .ZN(n1207) );
XNOR2_X1 U913 ( .A(G116), .B(n1189), .ZN(G18) );
NAND4_X1 U914 ( .A1(n1194), .A2(n1045), .A3(n1050), .A4(n1231), .ZN(n1189) );
NOR2_X1 U915 ( .A1(n1235), .A2(n1238), .ZN(n1050) );
INV_X1 U916 ( .A(n1053), .ZN(n1194) );
NAND2_X1 U917 ( .A1(n1038), .A2(n1196), .ZN(n1053) );
INV_X1 U918 ( .A(n1183), .ZN(n1196) );
XOR2_X1 U919 ( .A(G113), .B(n1239), .Z(G15) );
NOR2_X1 U920 ( .A1(n1183), .A2(n1198), .ZN(n1239) );
NAND4_X1 U921 ( .A1(n1045), .A2(n1038), .A3(n1049), .A4(n1231), .ZN(n1198) );
NAND2_X1 U922 ( .A1(n1240), .A2(n1241), .ZN(n1049) );
NAND2_X1 U923 ( .A1(n1043), .A2(n1242), .ZN(n1241) );
INV_X1 U924 ( .A(KEYINPUT8), .ZN(n1242) );
NAND3_X1 U925 ( .A1(n1238), .A2(n1235), .A3(KEYINPUT8), .ZN(n1240) );
NOR2_X1 U926 ( .A1(n1243), .A2(n1058), .ZN(n1038) );
NOR2_X1 U927 ( .A1(n1070), .A2(n1237), .ZN(n1045) );
INV_X1 U928 ( .A(n1232), .ZN(n1237) );
XOR2_X1 U929 ( .A(n1188), .B(n1244), .Z(G12) );
XNOR2_X1 U930 ( .A(G110), .B(KEYINPUT2), .ZN(n1244) );
NAND3_X1 U931 ( .A1(n1043), .A2(n1191), .A3(n1046), .ZN(n1188) );
NOR2_X1 U932 ( .A1(n1232), .A2(n1236), .ZN(n1046) );
INV_X1 U933 ( .A(n1070), .ZN(n1236) );
XNOR2_X1 U934 ( .A(n1245), .B(n1128), .ZN(n1070) );
AND2_X1 U935 ( .A1(G217), .A2(n1246), .ZN(n1128) );
NAND2_X1 U936 ( .A1(n1126), .A2(n1247), .ZN(n1245) );
XOR2_X1 U937 ( .A(n1248), .B(n1249), .Z(n1126) );
XOR2_X1 U938 ( .A(n1250), .B(n1251), .Z(n1249) );
XNOR2_X1 U939 ( .A(n1252), .B(n1253), .ZN(n1251) );
NAND2_X1 U940 ( .A1(KEYINPUT50), .A2(n1218), .ZN(n1253) );
NAND2_X1 U941 ( .A1(n1254), .A2(KEYINPUT56), .ZN(n1252) );
XOR2_X1 U942 ( .A(n1255), .B(n1256), .Z(n1254) );
NAND2_X1 U943 ( .A1(G221), .A2(n1257), .ZN(n1250) );
XNOR2_X1 U944 ( .A(G110), .B(n1258), .ZN(n1248) );
XNOR2_X1 U945 ( .A(n1106), .B(G119), .ZN(n1258) );
NAND2_X1 U946 ( .A1(n1259), .A2(n1260), .ZN(n1232) );
NAND2_X1 U947 ( .A1(n1075), .A2(n1261), .ZN(n1260) );
XOR2_X1 U948 ( .A(n1262), .B(KEYINPUT20), .Z(n1259) );
OR2_X1 U949 ( .A1(n1261), .A2(n1075), .ZN(n1262) );
AND2_X1 U950 ( .A1(n1247), .A2(n1263), .ZN(n1075) );
NAND2_X1 U951 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NAND2_X1 U952 ( .A1(n1141), .A2(n1144), .ZN(n1265) );
XOR2_X1 U953 ( .A(KEYINPUT5), .B(n1266), .Z(n1264) );
NOR2_X1 U954 ( .A1(n1141), .A2(n1144), .ZN(n1266) );
XOR2_X1 U955 ( .A(n1204), .B(n1267), .Z(n1144) );
XOR2_X1 U956 ( .A(n1160), .B(n1268), .Z(n1267) );
XOR2_X1 U957 ( .A(n1269), .B(G101), .Z(n1141) );
NAND3_X1 U958 ( .A1(n1270), .A2(n1271), .A3(G210), .ZN(n1269) );
XOR2_X1 U959 ( .A(G472), .B(KEYINPUT22), .Z(n1261) );
NOR3_X1 U960 ( .A1(n1223), .A2(n1195), .A3(n1183), .ZN(n1191) );
NAND2_X1 U961 ( .A1(n1216), .A2(n1069), .ZN(n1183) );
XOR2_X1 U962 ( .A(n1272), .B(n1167), .Z(n1069) );
NAND2_X1 U963 ( .A1(G210), .A2(n1273), .ZN(n1167) );
NAND2_X1 U964 ( .A1(n1274), .A2(n1247), .ZN(n1272) );
XOR2_X1 U965 ( .A(n1275), .B(n1276), .Z(n1274) );
XNOR2_X1 U966 ( .A(G125), .B(n1201), .ZN(n1276) );
NAND2_X1 U967 ( .A1(G224), .A2(n1270), .ZN(n1201) );
XOR2_X1 U968 ( .A(n1204), .B(n1166), .Z(n1275) );
XNOR2_X1 U969 ( .A(n1277), .B(n1278), .ZN(n1166) );
NOR2_X1 U970 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NOR2_X1 U971 ( .A1(n1281), .A2(n1119), .ZN(n1280) );
XNOR2_X1 U972 ( .A(n1282), .B(n1268), .ZN(n1119) );
INV_X1 U973 ( .A(KEYINPUT0), .ZN(n1281) );
NOR3_X1 U974 ( .A1(KEYINPUT0), .A2(n1268), .A3(n1282), .ZN(n1279) );
XNOR2_X1 U975 ( .A(G101), .B(n1283), .ZN(n1282) );
XNOR2_X1 U976 ( .A(n1284), .B(G104), .ZN(n1283) );
XNOR2_X1 U977 ( .A(G113), .B(n1285), .ZN(n1268) );
XOR2_X1 U978 ( .A(G119), .B(G116), .Z(n1285) );
NAND2_X1 U979 ( .A1(n1286), .A2(KEYINPUT19), .ZN(n1277) );
XNOR2_X1 U980 ( .A(G110), .B(G122), .ZN(n1286) );
NAND2_X1 U981 ( .A1(n1287), .A2(n1288), .ZN(n1204) );
NAND2_X1 U982 ( .A1(n1289), .A2(n1218), .ZN(n1288) );
XOR2_X1 U983 ( .A(KEYINPUT60), .B(n1290), .Z(n1289) );
NAND2_X1 U984 ( .A1(G128), .A2(n1291), .ZN(n1287) );
XNOR2_X1 U985 ( .A(n1290), .B(KEYINPUT3), .ZN(n1291) );
XNOR2_X1 U986 ( .A(G143), .B(n1255), .ZN(n1290) );
XOR2_X1 U987 ( .A(n1062), .B(KEYINPUT43), .Z(n1216) );
AND2_X1 U988 ( .A1(G214), .A2(n1273), .ZN(n1062) );
NAND2_X1 U989 ( .A1(n1292), .A2(n1271), .ZN(n1273) );
INV_X1 U990 ( .A(n1231), .ZN(n1195) );
NAND2_X1 U991 ( .A1(n1293), .A2(n1225), .ZN(n1231) );
NAND2_X1 U992 ( .A1(n1034), .A2(n1294), .ZN(n1225) );
INV_X1 U993 ( .A(n1030), .ZN(n1294) );
XOR2_X1 U994 ( .A(G953), .B(KEYINPUT6), .Z(n1030) );
AND2_X1 U995 ( .A1(G952), .A2(n1295), .ZN(n1034) );
NAND2_X1 U996 ( .A1(n1226), .A2(n1114), .ZN(n1293) );
INV_X1 U997 ( .A(G898), .ZN(n1114) );
AND3_X1 U998 ( .A1(G902), .A2(n1295), .A3(G953), .ZN(n1226) );
NAND2_X1 U999 ( .A1(G237), .A2(n1296), .ZN(n1295) );
INV_X1 U1000 ( .A(n1222), .ZN(n1223) );
XOR2_X1 U1001 ( .A(n1060), .B(KEYINPUT63), .Z(n1222) );
NOR2_X1 U1002 ( .A1(n1059), .A2(n1058), .ZN(n1060) );
AND2_X1 U1003 ( .A1(G221), .A2(n1246), .ZN(n1058) );
NAND2_X1 U1004 ( .A1(n1296), .A2(n1292), .ZN(n1246) );
XOR2_X1 U1005 ( .A(G234), .B(KEYINPUT18), .Z(n1296) );
INV_X1 U1006 ( .A(n1243), .ZN(n1059) );
XNOR2_X1 U1007 ( .A(n1297), .B(G469), .ZN(n1243) );
NAND3_X1 U1008 ( .A1(n1298), .A2(n1299), .A3(n1247), .ZN(n1297) );
NAND2_X1 U1009 ( .A1(KEYINPUT59), .A2(n1300), .ZN(n1299) );
XOR2_X1 U1010 ( .A(n1301), .B(n1161), .Z(n1300) );
NAND3_X1 U1011 ( .A1(n1301), .A2(n1161), .A3(n1302), .ZN(n1298) );
INV_X1 U1012 ( .A(KEYINPUT59), .ZN(n1302) );
XOR2_X1 U1013 ( .A(n1303), .B(n1304), .Z(n1161) );
XNOR2_X1 U1014 ( .A(n1305), .B(G110), .ZN(n1304) );
INV_X1 U1015 ( .A(G140), .ZN(n1305) );
NAND2_X1 U1016 ( .A1(G227), .A2(n1270), .ZN(n1303) );
NAND2_X1 U1017 ( .A1(n1306), .A2(n1307), .ZN(n1301) );
NAND2_X1 U1018 ( .A1(n1308), .A2(n1159), .ZN(n1307) );
INV_X1 U1019 ( .A(n1309), .ZN(n1159) );
NAND2_X1 U1020 ( .A1(n1309), .A2(n1310), .ZN(n1306) );
XNOR2_X1 U1021 ( .A(n1308), .B(KEYINPUT42), .ZN(n1310) );
XOR2_X1 U1022 ( .A(n1090), .B(n1160), .Z(n1308) );
XNOR2_X1 U1023 ( .A(G131), .B(n1311), .ZN(n1160) );
XNOR2_X1 U1024 ( .A(n1106), .B(G134), .ZN(n1311) );
INV_X1 U1025 ( .A(G137), .ZN(n1106) );
XNOR2_X1 U1026 ( .A(n1312), .B(n1255), .ZN(n1090) );
XNOR2_X1 U1027 ( .A(n1313), .B(n1218), .ZN(n1312) );
NAND2_X1 U1028 ( .A1(n1314), .A2(KEYINPUT27), .ZN(n1313) );
XNOR2_X1 U1029 ( .A(G143), .B(KEYINPUT30), .ZN(n1314) );
XNOR2_X1 U1030 ( .A(n1315), .B(n1316), .ZN(n1309) );
NOR2_X1 U1031 ( .A1(G101), .A2(KEYINPUT49), .ZN(n1316) );
NAND2_X1 U1032 ( .A1(n1317), .A2(n1318), .ZN(n1315) );
NAND2_X1 U1033 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
XNOR2_X1 U1034 ( .A(KEYINPUT36), .B(n1321), .ZN(n1320) );
INV_X1 U1035 ( .A(G104), .ZN(n1321) );
XNOR2_X1 U1036 ( .A(KEYINPUT54), .B(n1284), .ZN(n1319) );
INV_X1 U1037 ( .A(G107), .ZN(n1284) );
NAND2_X1 U1038 ( .A1(n1322), .A2(n1323), .ZN(n1317) );
XNOR2_X1 U1039 ( .A(KEYINPUT36), .B(G104), .ZN(n1323) );
XNOR2_X1 U1040 ( .A(G107), .B(KEYINPUT28), .ZN(n1322) );
NOR2_X1 U1041 ( .A1(n1235), .A2(n1234), .ZN(n1043) );
INV_X1 U1042 ( .A(n1238), .ZN(n1234) );
XOR2_X1 U1043 ( .A(n1324), .B(n1133), .Z(n1238) );
INV_X1 U1044 ( .A(G478), .ZN(n1133) );
NAND2_X1 U1045 ( .A1(KEYINPUT11), .A2(n1074), .ZN(n1324) );
NAND2_X1 U1046 ( .A1(n1131), .A2(n1247), .ZN(n1074) );
XNOR2_X1 U1047 ( .A(n1325), .B(n1326), .ZN(n1131) );
XOR2_X1 U1048 ( .A(n1327), .B(n1328), .Z(n1326) );
NAND2_X1 U1049 ( .A1(KEYINPUT4), .A2(n1329), .ZN(n1328) );
XOR2_X1 U1050 ( .A(G122), .B(G116), .Z(n1329) );
NAND2_X1 U1051 ( .A1(n1330), .A2(n1331), .ZN(n1327) );
OR2_X1 U1052 ( .A1(n1332), .A2(G134), .ZN(n1331) );
XOR2_X1 U1053 ( .A(n1333), .B(KEYINPUT47), .Z(n1330) );
NAND2_X1 U1054 ( .A1(G134), .A2(n1332), .ZN(n1333) );
XNOR2_X1 U1055 ( .A(G143), .B(n1218), .ZN(n1332) );
INV_X1 U1056 ( .A(G128), .ZN(n1218) );
XNOR2_X1 U1057 ( .A(G107), .B(n1334), .ZN(n1325) );
AND2_X1 U1058 ( .A1(n1257), .A2(G217), .ZN(n1334) );
AND2_X1 U1059 ( .A1(G234), .A2(n1270), .ZN(n1257) );
XOR2_X1 U1060 ( .A(n1071), .B(n1138), .Z(n1235) );
INV_X1 U1061 ( .A(G475), .ZN(n1138) );
NAND2_X1 U1062 ( .A1(n1136), .A2(n1247), .ZN(n1071) );
XNOR2_X1 U1063 ( .A(n1292), .B(KEYINPUT23), .ZN(n1247) );
INV_X1 U1064 ( .A(G902), .ZN(n1292) );
XNOR2_X1 U1065 ( .A(n1335), .B(n1336), .ZN(n1136) );
XOR2_X1 U1066 ( .A(n1337), .B(n1338), .Z(n1336) );
XNOR2_X1 U1067 ( .A(n1339), .B(G131), .ZN(n1338) );
INV_X1 U1068 ( .A(G143), .ZN(n1339) );
NOR2_X1 U1069 ( .A1(KEYINPUT34), .A2(n1340), .ZN(n1337) );
XOR2_X1 U1070 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1071 ( .A(KEYINPUT1), .B(G122), .Z(n1342) );
XNOR2_X1 U1072 ( .A(G113), .B(G104), .ZN(n1341) );
XNOR2_X1 U1073 ( .A(n1256), .B(n1343), .ZN(n1335) );
XOR2_X1 U1074 ( .A(n1344), .B(n1345), .Z(n1343) );
NAND2_X1 U1075 ( .A1(KEYINPUT35), .A2(n1255), .ZN(n1345) );
XNOR2_X1 U1076 ( .A(G146), .B(KEYINPUT26), .ZN(n1255) );
NAND3_X1 U1077 ( .A1(n1270), .A2(n1271), .A3(G214), .ZN(n1344) );
INV_X1 U1078 ( .A(G237), .ZN(n1271) );
XNOR2_X1 U1079 ( .A(n1081), .B(KEYINPUT21), .ZN(n1270) );
INV_X1 U1080 ( .A(G953), .ZN(n1081) );
XOR2_X1 U1081 ( .A(n1096), .B(KEYINPUT12), .Z(n1256) );
XOR2_X1 U1082 ( .A(G140), .B(G125), .Z(n1096) );
endmodule


