//Key = 0110101001011111000100110000001010110111101000000110001111101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267;

XNOR2_X1 U704 ( .A(n966), .B(n967), .ZN(G9) );
NOR2_X1 U705 ( .A1(n968), .A2(n969), .ZN(n967) );
NOR2_X1 U706 ( .A1(n970), .A2(n971), .ZN(G75) );
NOR3_X1 U707 ( .A1(n972), .A2(n973), .A3(n974), .ZN(n971) );
NOR2_X1 U708 ( .A1(n975), .A2(n976), .ZN(n973) );
INV_X1 U709 ( .A(n977), .ZN(n976) );
NOR2_X1 U710 ( .A1(n978), .A2(n979), .ZN(n975) );
NOR2_X1 U711 ( .A1(KEYINPUT49), .A2(n980), .ZN(n979) );
AND4_X1 U712 ( .A1(n981), .A2(n982), .A3(n983), .A4(n984), .ZN(n980) );
NOR2_X1 U713 ( .A1(n985), .A2(n986), .ZN(n978) );
NOR2_X1 U714 ( .A1(n987), .A2(n988), .ZN(n985) );
NOR2_X1 U715 ( .A1(n989), .A2(n990), .ZN(n988) );
NOR2_X1 U716 ( .A1(n991), .A2(n992), .ZN(n989) );
AND2_X1 U717 ( .A1(n981), .A2(n993), .ZN(n992) );
NOR2_X1 U718 ( .A1(n994), .A2(n995), .ZN(n991) );
NOR2_X1 U719 ( .A1(n996), .A2(n997), .ZN(n994) );
XOR2_X1 U720 ( .A(KEYINPUT17), .B(n998), .Z(n997) );
AND4_X1 U721 ( .A1(n981), .A2(n982), .A3(n983), .A4(KEYINPUT49), .ZN(n987) );
NAND3_X1 U722 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n972) );
NAND3_X1 U723 ( .A1(n981), .A2(n1002), .A3(n984), .ZN(n1001) );
INV_X1 U724 ( .A(n986), .ZN(n984) );
NAND2_X1 U725 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND3_X1 U726 ( .A1(n982), .A2(n1005), .A3(n977), .ZN(n1004) );
NAND2_X1 U727 ( .A1(n1006), .A2(n1007), .ZN(n1003) );
NAND3_X1 U728 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1007) );
NAND3_X1 U729 ( .A1(n1011), .A2(n982), .A3(n1012), .ZN(n1010) );
INV_X1 U730 ( .A(n995), .ZN(n982) );
INV_X1 U731 ( .A(n1013), .ZN(n1009) );
NAND3_X1 U732 ( .A1(n1014), .A2(n977), .A3(n1015), .ZN(n1008) );
NOR3_X1 U733 ( .A1(n1016), .A2(G953), .A3(G952), .ZN(n970) );
INV_X1 U734 ( .A(n999), .ZN(n1016) );
NAND4_X1 U735 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n999) );
NOR4_X1 U736 ( .A1(n1012), .A2(n1021), .A3(n995), .A4(n1022), .ZN(n1020) );
XNOR2_X1 U737 ( .A(n1023), .B(n1011), .ZN(n1019) );
XNOR2_X1 U738 ( .A(KEYINPUT10), .B(KEYINPUT0), .ZN(n1023) );
XOR2_X1 U739 ( .A(n1024), .B(n1025), .Z(n1018) );
XOR2_X1 U740 ( .A(KEYINPUT27), .B(G478), .Z(n1025) );
XNOR2_X1 U741 ( .A(n1026), .B(n1027), .ZN(n1017) );
NAND2_X1 U742 ( .A1(KEYINPUT34), .A2(n1028), .ZN(n1026) );
XOR2_X1 U743 ( .A(n1029), .B(n1030), .Z(G72) );
NOR2_X1 U744 ( .A1(n1031), .A2(n1000), .ZN(n1030) );
NOR2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U746 ( .A1(n1034), .A2(n1035), .ZN(n1029) );
NAND2_X1 U747 ( .A1(n1036), .A2(n1000), .ZN(n1035) );
XNOR2_X1 U748 ( .A(n1037), .B(n1038), .ZN(n1036) );
NAND3_X1 U749 ( .A1(n1037), .A2(G900), .A3(G953), .ZN(n1034) );
NOR2_X1 U750 ( .A1(KEYINPUT44), .A2(n1039), .ZN(n1037) );
XOR2_X1 U751 ( .A(n1040), .B(n1041), .Z(n1039) );
XNOR2_X1 U752 ( .A(n1042), .B(n1043), .ZN(n1041) );
NOR2_X1 U753 ( .A1(G125), .A2(KEYINPUT31), .ZN(n1043) );
INV_X1 U754 ( .A(G131), .ZN(n1042) );
XOR2_X1 U755 ( .A(n1044), .B(n1045), .Z(n1040) );
NOR3_X1 U756 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
NOR2_X1 U757 ( .A1(KEYINPUT14), .A2(n1049), .ZN(n1048) );
NOR3_X1 U758 ( .A1(G134), .A2(n1050), .A3(n1051), .ZN(n1047) );
NOR2_X1 U759 ( .A1(G137), .A2(n1052), .ZN(n1046) );
NOR2_X1 U760 ( .A1(n1051), .A2(n1053), .ZN(n1052) );
XNOR2_X1 U761 ( .A(KEYINPUT3), .B(n1049), .ZN(n1053) );
INV_X1 U762 ( .A(G134), .ZN(n1049) );
INV_X1 U763 ( .A(KEYINPUT14), .ZN(n1051) );
XOR2_X1 U764 ( .A(n1054), .B(n1055), .Z(G69) );
NAND2_X1 U765 ( .A1(G953), .A2(n1056), .ZN(n1055) );
NAND2_X1 U766 ( .A1(G898), .A2(G224), .ZN(n1056) );
NAND4_X1 U767 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1054) );
NAND4_X1 U768 ( .A1(KEYINPUT2), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1060) );
INV_X1 U769 ( .A(n1064), .ZN(n1063) );
NAND2_X1 U770 ( .A1(n1064), .A2(n1065), .ZN(n1059) );
NAND3_X1 U771 ( .A1(n1066), .A2(n1000), .A3(KEYINPUT2), .ZN(n1065) );
XNOR2_X1 U772 ( .A(n1067), .B(n1068), .ZN(n1064) );
NAND2_X1 U773 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NAND2_X1 U774 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XOR2_X1 U775 ( .A(n1073), .B(KEYINPUT36), .Z(n1069) );
OR2_X1 U776 ( .A1(n1072), .A2(n1071), .ZN(n1073) );
NAND2_X1 U777 ( .A1(G953), .A2(n1074), .ZN(n1058) );
OR2_X1 U778 ( .A1(n1061), .A2(n1062), .ZN(n1057) );
NOR2_X1 U779 ( .A1(G953), .A2(n1075), .ZN(n1062) );
INV_X1 U780 ( .A(KEYINPUT25), .ZN(n1061) );
NOR2_X1 U781 ( .A1(n1076), .A2(n1077), .ZN(G66) );
XOR2_X1 U782 ( .A(n1078), .B(n1079), .Z(n1077) );
NAND2_X1 U783 ( .A1(n1080), .A2(n1028), .ZN(n1078) );
NOR2_X1 U784 ( .A1(n1081), .A2(n1082), .ZN(G63) );
XNOR2_X1 U785 ( .A(n1083), .B(n1084), .ZN(n1082) );
XOR2_X1 U786 ( .A(n1085), .B(KEYINPUT54), .Z(n1083) );
NAND2_X1 U787 ( .A1(n1080), .A2(G478), .ZN(n1085) );
NOR2_X1 U788 ( .A1(G952), .A2(n1086), .ZN(n1081) );
XNOR2_X1 U789 ( .A(KEYINPUT1), .B(n1000), .ZN(n1086) );
NOR2_X1 U790 ( .A1(n1076), .A2(n1087), .ZN(G60) );
XOR2_X1 U791 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U792 ( .A1(n1090), .A2(n1080), .ZN(n1088) );
XNOR2_X1 U793 ( .A(G475), .B(KEYINPUT56), .ZN(n1090) );
XOR2_X1 U794 ( .A(n1091), .B(n1092), .Z(G6) );
NAND2_X1 U795 ( .A1(KEYINPUT4), .A2(G104), .ZN(n1092) );
NOR2_X1 U796 ( .A1(n1076), .A2(n1093), .ZN(G57) );
XOR2_X1 U797 ( .A(n1094), .B(n1095), .Z(n1093) );
XNOR2_X1 U798 ( .A(n1096), .B(n1097), .ZN(n1095) );
NAND2_X1 U799 ( .A1(KEYINPUT12), .A2(n1098), .ZN(n1097) );
XNOR2_X1 U800 ( .A(n1099), .B(n1100), .ZN(n1098) );
NAND2_X1 U801 ( .A1(KEYINPUT40), .A2(n1101), .ZN(n1100) );
NAND2_X1 U802 ( .A1(n1102), .A2(KEYINPUT37), .ZN(n1096) );
XOR2_X1 U803 ( .A(n1103), .B(n1104), .Z(n1102) );
XNOR2_X1 U804 ( .A(n1105), .B(n1106), .ZN(n1104) );
NAND2_X1 U805 ( .A1(n1080), .A2(G472), .ZN(n1094) );
NOR2_X1 U806 ( .A1(n1076), .A2(n1107), .ZN(G54) );
XOR2_X1 U807 ( .A(n1108), .B(n1109), .Z(n1107) );
AND2_X1 U808 ( .A1(G469), .A2(n1080), .ZN(n1109) );
NOR2_X1 U809 ( .A1(KEYINPUT41), .A2(n1110), .ZN(n1108) );
XOR2_X1 U810 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U811 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U812 ( .A(n1115), .B(KEYINPUT15), .Z(n1114) );
NAND2_X1 U813 ( .A1(n1116), .A2(KEYINPUT32), .ZN(n1113) );
XOR2_X1 U814 ( .A(n1117), .B(G110), .Z(n1116) );
NAND2_X1 U815 ( .A1(KEYINPUT30), .A2(n1118), .ZN(n1117) );
XOR2_X1 U816 ( .A(n1119), .B(n1120), .Z(n1111) );
XNOR2_X1 U817 ( .A(n1121), .B(n1122), .ZN(n1119) );
NOR2_X1 U818 ( .A1(n1076), .A2(n1123), .ZN(G51) );
XNOR2_X1 U819 ( .A(n1124), .B(n1125), .ZN(n1123) );
XOR2_X1 U820 ( .A(n1126), .B(KEYINPUT6), .Z(n1125) );
NAND2_X1 U821 ( .A1(n1080), .A2(n1127), .ZN(n1126) );
AND2_X1 U822 ( .A1(G902), .A2(n974), .ZN(n1080) );
NAND2_X1 U823 ( .A1(n1038), .A2(n1075), .ZN(n974) );
INV_X1 U824 ( .A(n1066), .ZN(n1075) );
NAND4_X1 U825 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1066) );
AND4_X1 U826 ( .A1(n1091), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1131) );
NAND4_X1 U827 ( .A1(n981), .A2(n1135), .A3(n993), .A4(n1136), .ZN(n1091) );
NOR2_X1 U828 ( .A1(n969), .A2(n1137), .ZN(n1136) );
NOR2_X1 U829 ( .A1(n1138), .A2(n1139), .ZN(n1130) );
NOR2_X1 U830 ( .A1(n1140), .A2(n969), .ZN(n1139) );
XOR2_X1 U831 ( .A(n968), .B(KEYINPUT21), .Z(n1140) );
NAND4_X1 U832 ( .A1(n993), .A2(n1005), .A3(n981), .A4(n1135), .ZN(n968) );
INV_X1 U833 ( .A(n1141), .ZN(n1138) );
AND4_X1 U834 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1038) );
NOR4_X1 U835 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1145) );
INV_X1 U836 ( .A(n1150), .ZN(n1148) );
INV_X1 U837 ( .A(n1151), .ZN(n1147) );
NOR2_X1 U838 ( .A1(n1152), .A2(n1153), .ZN(n1144) );
NOR2_X1 U839 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XNOR2_X1 U840 ( .A(KEYINPUT13), .B(n1137), .ZN(n1155) );
NOR2_X1 U841 ( .A1(n1000), .A2(G952), .ZN(n1076) );
XNOR2_X1 U842 ( .A(n1156), .B(n1152), .ZN(G48) );
AND3_X1 U843 ( .A1(n1157), .A2(n1158), .A3(n983), .ZN(n1152) );
XOR2_X1 U844 ( .A(n1142), .B(n1159), .Z(G45) );
NAND2_X1 U845 ( .A1(KEYINPUT55), .A2(G143), .ZN(n1159) );
NAND4_X1 U846 ( .A1(n1158), .A2(n993), .A3(n996), .A4(n1160), .ZN(n1142) );
AND3_X1 U847 ( .A1(n1161), .A2(n1162), .A3(n1021), .ZN(n1160) );
XNOR2_X1 U848 ( .A(G140), .B(n1163), .ZN(G42) );
NOR2_X1 U849 ( .A1(n1164), .A2(KEYINPUT43), .ZN(n1163) );
INV_X1 U850 ( .A(n1143), .ZN(n1164) );
NAND3_X1 U851 ( .A1(n983), .A2(n1165), .A3(n998), .ZN(n1143) );
XOR2_X1 U852 ( .A(n1166), .B(n1167), .Z(G39) );
XNOR2_X1 U853 ( .A(KEYINPUT60), .B(n1050), .ZN(n1167) );
NAND2_X1 U854 ( .A1(KEYINPUT23), .A2(n1149), .ZN(n1166) );
AND3_X1 U855 ( .A1(n977), .A2(n1157), .A3(n1006), .ZN(n1149) );
XNOR2_X1 U856 ( .A(G134), .B(n1150), .ZN(G36) );
NAND3_X1 U857 ( .A1(n1165), .A2(n1005), .A3(n996), .ZN(n1150) );
XNOR2_X1 U858 ( .A(G131), .B(n1151), .ZN(G33) );
NAND3_X1 U859 ( .A1(n983), .A2(n1165), .A3(n996), .ZN(n1151) );
AND3_X1 U860 ( .A1(n993), .A2(n1162), .A3(n977), .ZN(n1165) );
NOR2_X1 U861 ( .A1(n1168), .A2(n1012), .ZN(n977) );
XOR2_X1 U862 ( .A(G128), .B(n1146), .Z(G30) );
AND3_X1 U863 ( .A1(n1158), .A2(n1005), .A3(n1157), .ZN(n1146) );
AND4_X1 U864 ( .A1(n993), .A2(n1169), .A3(n1022), .A4(n1162), .ZN(n1157) );
NAND2_X1 U865 ( .A1(n1170), .A2(n1171), .ZN(G3) );
NAND2_X1 U866 ( .A1(n1172), .A2(n1141), .ZN(n1171) );
XOR2_X1 U867 ( .A(KEYINPUT19), .B(n1173), .Z(n1170) );
NOR2_X1 U868 ( .A1(n1141), .A2(n1172), .ZN(n1173) );
XNOR2_X1 U869 ( .A(KEYINPUT45), .B(n1101), .ZN(n1172) );
NAND2_X1 U870 ( .A1(n1174), .A2(n996), .ZN(n1141) );
XOR2_X1 U871 ( .A(G125), .B(n1175), .Z(G27) );
NOR3_X1 U872 ( .A1(n1154), .A2(KEYINPUT16), .A3(n1137), .ZN(n1175) );
NAND3_X1 U873 ( .A1(n998), .A2(n1162), .A3(n1013), .ZN(n1154) );
NAND2_X1 U874 ( .A1(n986), .A2(n1176), .ZN(n1162) );
NAND4_X1 U875 ( .A1(G953), .A2(G902), .A3(n1177), .A4(n1033), .ZN(n1176) );
INV_X1 U876 ( .A(G900), .ZN(n1033) );
XNOR2_X1 U877 ( .A(G122), .B(n1128), .ZN(G24) );
NAND4_X1 U878 ( .A1(n1178), .A2(n981), .A3(n1161), .A4(n1021), .ZN(n1128) );
NOR2_X1 U879 ( .A1(n1022), .A2(n1169), .ZN(n981) );
XNOR2_X1 U880 ( .A(G119), .B(n1129), .ZN(G21) );
NAND4_X1 U881 ( .A1(n1178), .A2(n1006), .A3(n1169), .A4(n1022), .ZN(n1129) );
XNOR2_X1 U882 ( .A(G116), .B(n1134), .ZN(G18) );
NAND3_X1 U883 ( .A1(n996), .A2(n1005), .A3(n1178), .ZN(n1134) );
AND2_X1 U884 ( .A1(n1179), .A2(n1161), .ZN(n1005) );
XNOR2_X1 U885 ( .A(n1180), .B(KEYINPUT51), .ZN(n1161) );
XOR2_X1 U886 ( .A(n1133), .B(n1181), .Z(G15) );
NOR2_X1 U887 ( .A1(KEYINPUT61), .A2(n1182), .ZN(n1181) );
XOR2_X1 U888 ( .A(KEYINPUT29), .B(G113), .Z(n1182) );
NAND3_X1 U889 ( .A1(n996), .A2(n983), .A3(n1178), .ZN(n1133) );
AND2_X1 U890 ( .A1(n1013), .A2(n1135), .ZN(n1178) );
NOR2_X1 U891 ( .A1(n995), .A2(n969), .ZN(n1013) );
INV_X1 U892 ( .A(n1158), .ZN(n969) );
NAND2_X1 U893 ( .A1(n1014), .A2(n1183), .ZN(n995) );
INV_X1 U894 ( .A(n1137), .ZN(n983) );
NAND2_X1 U895 ( .A1(n1180), .A2(n1021), .ZN(n1137) );
NOR2_X1 U896 ( .A1(n1169), .A2(n1184), .ZN(n996) );
XNOR2_X1 U897 ( .A(G110), .B(n1132), .ZN(G12) );
NAND2_X1 U898 ( .A1(n1174), .A2(n998), .ZN(n1132) );
AND2_X1 U899 ( .A1(n1184), .A2(n1169), .ZN(n998) );
XNOR2_X1 U900 ( .A(n1027), .B(n1028), .ZN(n1169) );
AND2_X1 U901 ( .A1(G217), .A2(n1185), .ZN(n1028) );
NAND2_X1 U902 ( .A1(n1186), .A2(n1187), .ZN(n1027) );
XOR2_X1 U903 ( .A(KEYINPUT18), .B(n1079), .Z(n1187) );
XNOR2_X1 U904 ( .A(n1188), .B(n1189), .ZN(n1079) );
XOR2_X1 U905 ( .A(n1190), .B(n1191), .Z(n1189) );
AND2_X1 U906 ( .A1(G221), .A2(n1192), .ZN(n1190) );
XNOR2_X1 U907 ( .A(n1193), .B(n1050), .ZN(n1188) );
NAND2_X1 U908 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
OR2_X1 U909 ( .A1(n1196), .A2(G110), .ZN(n1195) );
XOR2_X1 U910 ( .A(n1197), .B(KEYINPUT8), .Z(n1194) );
NAND2_X1 U911 ( .A1(G110), .A2(n1196), .ZN(n1197) );
XOR2_X1 U912 ( .A(G119), .B(G128), .Z(n1196) );
INV_X1 U913 ( .A(n1022), .ZN(n1184) );
XNOR2_X1 U914 ( .A(n1198), .B(G472), .ZN(n1022) );
NAND3_X1 U915 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1198) );
XNOR2_X1 U916 ( .A(KEYINPUT35), .B(n1186), .ZN(n1201) );
NAND2_X1 U917 ( .A1(n1202), .A2(n1203), .ZN(n1200) );
NAND2_X1 U918 ( .A1(KEYINPUT9), .A2(n1101), .ZN(n1203) );
XOR2_X1 U919 ( .A(n1204), .B(n1205), .Z(n1202) );
NOR2_X1 U920 ( .A1(n1099), .A2(KEYINPUT47), .ZN(n1204) );
INV_X1 U921 ( .A(n1206), .ZN(n1099) );
NAND3_X1 U922 ( .A1(KEYINPUT9), .A2(n1101), .A3(n1207), .ZN(n1199) );
XOR2_X1 U923 ( .A(n1208), .B(n1205), .Z(n1207) );
XNOR2_X1 U924 ( .A(n1209), .B(n1210), .ZN(n1205) );
XNOR2_X1 U925 ( .A(n1211), .B(n1106), .ZN(n1210) );
XOR2_X1 U926 ( .A(G146), .B(n1212), .Z(n1106) );
NAND2_X1 U927 ( .A1(KEYINPUT39), .A2(n1103), .ZN(n1211) );
NAND2_X1 U928 ( .A1(n1213), .A2(n1214), .ZN(n1209) );
OR2_X1 U929 ( .A1(KEYINPUT26), .A2(n1105), .ZN(n1214) );
NAND2_X1 U930 ( .A1(KEYINPUT7), .A2(n1105), .ZN(n1213) );
XNOR2_X1 U931 ( .A(G113), .B(n1215), .ZN(n1105) );
NOR2_X1 U932 ( .A1(KEYINPUT46), .A2(n1216), .ZN(n1215) );
XNOR2_X1 U933 ( .A(G116), .B(G119), .ZN(n1216) );
NOR2_X1 U934 ( .A1(KEYINPUT47), .A2(n1206), .ZN(n1208) );
NAND2_X1 U935 ( .A1(n1217), .A2(G210), .ZN(n1206) );
INV_X1 U936 ( .A(G101), .ZN(n1101) );
AND4_X1 U937 ( .A1(n1006), .A2(n1158), .A3(n993), .A4(n1135), .ZN(n1174) );
NAND2_X1 U938 ( .A1(n986), .A2(n1218), .ZN(n1135) );
NAND4_X1 U939 ( .A1(G953), .A2(G902), .A3(n1177), .A4(n1074), .ZN(n1218) );
INV_X1 U940 ( .A(G898), .ZN(n1074) );
NAND3_X1 U941 ( .A1(n1177), .A2(n1000), .A3(G952), .ZN(n986) );
NAND2_X1 U942 ( .A1(G237), .A2(G234), .ZN(n1177) );
NOR2_X1 U943 ( .A1(n1014), .A2(n1015), .ZN(n993) );
INV_X1 U944 ( .A(n1183), .ZN(n1015) );
NAND2_X1 U945 ( .A1(G221), .A2(n1185), .ZN(n1183) );
NAND2_X1 U946 ( .A1(G234), .A2(n1219), .ZN(n1185) );
XOR2_X1 U947 ( .A(n1220), .B(G469), .Z(n1014) );
NAND2_X1 U948 ( .A1(n1221), .A2(n1186), .ZN(n1220) );
XOR2_X1 U949 ( .A(n1222), .B(n1223), .Z(n1221) );
XNOR2_X1 U950 ( .A(n1120), .B(n1044), .ZN(n1223) );
XOR2_X1 U951 ( .A(n1224), .B(n1225), .Z(n1044) );
XNOR2_X1 U952 ( .A(n1115), .B(n1118), .ZN(n1224) );
INV_X1 U953 ( .A(G140), .ZN(n1118) );
NAND2_X1 U954 ( .A1(KEYINPUT57), .A2(n1156), .ZN(n1115) );
INV_X1 U955 ( .A(G146), .ZN(n1156) );
XNOR2_X1 U956 ( .A(n1226), .B(n1227), .ZN(n1120) );
NOR2_X1 U957 ( .A1(G953), .A2(n1032), .ZN(n1227) );
INV_X1 U958 ( .A(G227), .ZN(n1032) );
XOR2_X1 U959 ( .A(n1228), .B(n1229), .Z(n1222) );
NOR2_X1 U960 ( .A1(KEYINPUT20), .A2(n1103), .ZN(n1229) );
XNOR2_X1 U961 ( .A(n1122), .B(G134), .ZN(n1103) );
XOR2_X1 U962 ( .A(G131), .B(n1230), .Z(n1122) );
XNOR2_X1 U963 ( .A(KEYINPUT38), .B(n1050), .ZN(n1230) );
INV_X1 U964 ( .A(G137), .ZN(n1050) );
XNOR2_X1 U965 ( .A(G110), .B(KEYINPUT11), .ZN(n1228) );
NOR2_X1 U966 ( .A1(n1011), .A2(n1012), .ZN(n1158) );
AND2_X1 U967 ( .A1(G214), .A2(n1231), .ZN(n1012) );
INV_X1 U968 ( .A(n1168), .ZN(n1011) );
XNOR2_X1 U969 ( .A(n1232), .B(n1127), .ZN(n1168) );
AND2_X1 U970 ( .A1(G210), .A2(n1231), .ZN(n1127) );
NAND2_X1 U971 ( .A1(n1233), .A2(n1219), .ZN(n1231) );
INV_X1 U972 ( .A(G902), .ZN(n1219) );
INV_X1 U973 ( .A(G237), .ZN(n1233) );
NAND2_X1 U974 ( .A1(n1186), .A2(n1124), .ZN(n1232) );
XNOR2_X1 U975 ( .A(n1234), .B(n1235), .ZN(n1124) );
XOR2_X1 U976 ( .A(n1071), .B(n1236), .Z(n1235) );
XNOR2_X1 U977 ( .A(n1068), .B(n1212), .ZN(n1236) );
XNOR2_X1 U978 ( .A(n1237), .B(n1238), .ZN(n1212) );
NOR2_X1 U979 ( .A1(G128), .A2(KEYINPUT59), .ZN(n1238) );
NAND2_X1 U980 ( .A1(KEYINPUT42), .A2(n1239), .ZN(n1237) );
XOR2_X1 U981 ( .A(G122), .B(G110), .Z(n1068) );
XOR2_X1 U982 ( .A(n1226), .B(KEYINPUT53), .Z(n1071) );
XNOR2_X1 U983 ( .A(G101), .B(n1240), .ZN(n1226) );
XNOR2_X1 U984 ( .A(n966), .B(G104), .ZN(n1240) );
XOR2_X1 U985 ( .A(n1241), .B(n1242), .Z(n1234) );
XOR2_X1 U986 ( .A(KEYINPUT22), .B(n1243), .Z(n1242) );
AND2_X1 U987 ( .A1(n1000), .A2(G224), .ZN(n1243) );
XOR2_X1 U988 ( .A(n1244), .B(n1245), .Z(n1241) );
NAND2_X1 U989 ( .A1(KEYINPUT58), .A2(n1072), .ZN(n1244) );
XNOR2_X1 U990 ( .A(n1246), .B(n1247), .ZN(n1072) );
XOR2_X1 U991 ( .A(G113), .B(n1248), .Z(n1247) );
NOR2_X1 U992 ( .A1(G119), .A2(KEYINPUT52), .ZN(n1248) );
XNOR2_X1 U993 ( .A(G116), .B(KEYINPUT48), .ZN(n1246) );
INV_X1 U994 ( .A(n990), .ZN(n1006) );
NAND2_X1 U995 ( .A1(n1179), .A2(n1180), .ZN(n990) );
XNOR2_X1 U996 ( .A(n1249), .B(G478), .ZN(n1180) );
NAND2_X1 U997 ( .A1(n1250), .A2(KEYINPUT50), .ZN(n1249) );
XOR2_X1 U998 ( .A(n1024), .B(KEYINPUT33), .Z(n1250) );
NAND2_X1 U999 ( .A1(n1084), .A2(n1186), .ZN(n1024) );
XOR2_X1 U1000 ( .A(n1251), .B(n1252), .Z(n1084) );
XOR2_X1 U1001 ( .A(n1253), .B(n1254), .Z(n1252) );
XNOR2_X1 U1002 ( .A(G122), .B(KEYINPUT62), .ZN(n1254) );
NAND2_X1 U1003 ( .A1(n1255), .A2(n1256), .ZN(n1253) );
INV_X1 U1004 ( .A(G116), .ZN(n1256) );
XNOR2_X1 U1005 ( .A(KEYINPUT5), .B(KEYINPUT24), .ZN(n1255) );
XNOR2_X1 U1006 ( .A(n1257), .B(n1258), .ZN(n1251) );
INV_X1 U1007 ( .A(n1121), .ZN(n1258) );
XOR2_X1 U1008 ( .A(G134), .B(n1225), .Z(n1121) );
XOR2_X1 U1009 ( .A(G128), .B(G143), .Z(n1225) );
XOR2_X1 U1010 ( .A(n1259), .B(n1260), .Z(n1257) );
NOR2_X1 U1011 ( .A1(KEYINPUT63), .A2(n966), .ZN(n1260) );
INV_X1 U1012 ( .A(G107), .ZN(n966) );
NAND2_X1 U1013 ( .A1(G217), .A2(n1192), .ZN(n1259) );
AND2_X1 U1014 ( .A1(G234), .A2(n1000), .ZN(n1192) );
INV_X1 U1015 ( .A(G953), .ZN(n1000) );
INV_X1 U1016 ( .A(n1021), .ZN(n1179) );
XNOR2_X1 U1017 ( .A(n1261), .B(G475), .ZN(n1021) );
NAND2_X1 U1018 ( .A1(n1186), .A2(n1089), .ZN(n1261) );
XNOR2_X1 U1019 ( .A(n1262), .B(n1263), .ZN(n1089) );
XOR2_X1 U1020 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U1021 ( .A(G122), .B(G113), .Z(n1265) );
XNOR2_X1 U1022 ( .A(n1239), .B(G131), .ZN(n1264) );
INV_X1 U1023 ( .A(G143), .ZN(n1239) );
XNOR2_X1 U1024 ( .A(n1191), .B(n1266), .ZN(n1262) );
XNOR2_X1 U1025 ( .A(G104), .B(n1267), .ZN(n1266) );
NAND2_X1 U1026 ( .A1(n1217), .A2(G214), .ZN(n1267) );
NOR2_X1 U1027 ( .A1(G953), .A2(G237), .ZN(n1217) );
XOR2_X1 U1028 ( .A(G140), .B(n1245), .Z(n1191) );
XOR2_X1 U1029 ( .A(G125), .B(G146), .Z(n1245) );
XNOR2_X1 U1030 ( .A(G902), .B(KEYINPUT28), .ZN(n1186) );
endmodule


