//Key = 0111000110110001010001101110000101000100001100011001100001000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404;

XNOR2_X1 U778 ( .A(n1075), .B(n1076), .ZN(G9) );
NOR2_X1 U779 ( .A1(n1077), .A2(n1078), .ZN(G75) );
NOR3_X1 U780 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NAND3_X1 U781 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1079) );
NAND2_X1 U782 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U783 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND4_X1 U784 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1088) );
NAND3_X1 U785 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1090) );
NAND2_X1 U786 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
OR2_X1 U787 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U788 ( .A1(n1100), .A2(n1101), .ZN(n1094) );
NAND2_X1 U789 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND2_X1 U790 ( .A1(KEYINPUT42), .A2(n1104), .ZN(n1103) );
NAND2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1102) );
OR3_X1 U792 ( .A1(n1107), .A2(KEYINPUT42), .A3(n1100), .ZN(n1093) );
NAND3_X1 U793 ( .A1(n1096), .A2(n1108), .A3(n1100), .ZN(n1087) );
NAND2_X1 U794 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND3_X1 U795 ( .A1(n1111), .A2(n1112), .A3(n1092), .ZN(n1110) );
NAND2_X1 U796 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
OR3_X1 U797 ( .A1(n1115), .A2(n1116), .A3(n1113), .ZN(n1111) );
NAND2_X1 U798 ( .A1(n1089), .A2(n1117), .ZN(n1109) );
INV_X1 U799 ( .A(n1118), .ZN(n1085) );
NOR3_X1 U800 ( .A1(n1119), .A2(G953), .A3(n1120), .ZN(n1077) );
INV_X1 U801 ( .A(n1082), .ZN(n1120) );
NAND4_X1 U802 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1082) );
NOR4_X1 U803 ( .A1(n1105), .A2(n1113), .A3(n1125), .A4(n1126), .ZN(n1124) );
XNOR2_X1 U804 ( .A(n1127), .B(n1128), .ZN(n1126) );
XNOR2_X1 U805 ( .A(n1129), .B(KEYINPUT2), .ZN(n1127) );
XNOR2_X1 U806 ( .A(G475), .B(n1130), .ZN(n1125) );
NOR2_X1 U807 ( .A1(n1131), .A2(KEYINPUT49), .ZN(n1130) );
NOR3_X1 U808 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1123) );
NOR2_X1 U809 ( .A1(KEYINPUT6), .A2(n1135), .ZN(n1134) );
NOR2_X1 U810 ( .A1(n1136), .A2(n1137), .ZN(n1133) );
INV_X1 U811 ( .A(KEYINPUT6), .ZN(n1137) );
NOR2_X1 U812 ( .A1(n1138), .A2(n1139), .ZN(n1136) );
NOR2_X1 U813 ( .A1(G902), .A2(n1140), .ZN(n1138) );
XNOR2_X1 U814 ( .A(n1141), .B(n1142), .ZN(n1132) );
XNOR2_X1 U815 ( .A(KEYINPUT15), .B(n1143), .ZN(n1122) );
XNOR2_X1 U816 ( .A(KEYINPUT30), .B(n1080), .ZN(n1119) );
INV_X1 U817 ( .A(G952), .ZN(n1080) );
XOR2_X1 U818 ( .A(n1144), .B(n1145), .Z(G72) );
NOR2_X1 U819 ( .A1(n1146), .A2(KEYINPUT44), .ZN(n1145) );
NOR2_X1 U820 ( .A1(G953), .A2(n1147), .ZN(n1146) );
XOR2_X1 U821 ( .A(n1148), .B(n1149), .Z(n1144) );
NOR2_X1 U822 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XOR2_X1 U823 ( .A(n1152), .B(n1153), .Z(n1151) );
XNOR2_X1 U824 ( .A(n1154), .B(n1155), .ZN(n1153) );
XNOR2_X1 U825 ( .A(G140), .B(n1156), .ZN(n1152) );
NOR2_X1 U826 ( .A1(G125), .A2(n1157), .ZN(n1156) );
XNOR2_X1 U827 ( .A(KEYINPUT55), .B(KEYINPUT22), .ZN(n1157) );
NAND2_X1 U828 ( .A1(n1158), .A2(n1159), .ZN(n1148) );
NAND2_X1 U829 ( .A1(G900), .A2(G227), .ZN(n1159) );
XNOR2_X1 U830 ( .A(KEYINPUT45), .B(n1083), .ZN(n1158) );
XOR2_X1 U831 ( .A(n1160), .B(n1161), .Z(G69) );
XOR2_X1 U832 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U833 ( .A1(G953), .A2(n1164), .ZN(n1163) );
NAND2_X1 U834 ( .A1(G898), .A2(G224), .ZN(n1164) );
NAND2_X1 U835 ( .A1(n1165), .A2(n1166), .ZN(n1162) );
NAND2_X1 U836 ( .A1(G953), .A2(n1167), .ZN(n1166) );
XNOR2_X1 U837 ( .A(n1168), .B(n1169), .ZN(n1165) );
NOR2_X1 U838 ( .A1(n1170), .A2(G953), .ZN(n1160) );
NOR2_X1 U839 ( .A1(n1171), .A2(n1172), .ZN(G66) );
XOR2_X1 U840 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U841 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND2_X1 U842 ( .A1(KEYINPUT21), .A2(n1177), .ZN(n1173) );
NOR2_X1 U843 ( .A1(n1171), .A2(n1178), .ZN(G63) );
XOR2_X1 U844 ( .A(n1179), .B(n1180), .Z(n1178) );
NAND2_X1 U845 ( .A1(n1181), .A2(G478), .ZN(n1179) );
NOR2_X1 U846 ( .A1(n1171), .A2(n1182), .ZN(G60) );
NOR3_X1 U847 ( .A1(n1131), .A2(n1183), .A3(n1184), .ZN(n1182) );
AND3_X1 U848 ( .A1(n1185), .A2(G475), .A3(n1181), .ZN(n1184) );
NOR2_X1 U849 ( .A1(n1186), .A2(n1185), .ZN(n1183) );
AND2_X1 U850 ( .A1(n1081), .A2(G475), .ZN(n1186) );
NAND2_X1 U851 ( .A1(n1187), .A2(n1188), .ZN(G6) );
NAND2_X1 U852 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U853 ( .A1(n1191), .A2(n1192), .ZN(n1189) );
NAND2_X1 U854 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
INV_X1 U855 ( .A(KEYINPUT3), .ZN(n1194) );
NAND2_X1 U856 ( .A1(KEYINPUT3), .A2(n1195), .ZN(n1191) );
OR2_X1 U857 ( .A1(n1195), .A2(n1190), .ZN(n1187) );
NAND2_X1 U858 ( .A1(KEYINPUT26), .A2(n1193), .ZN(n1195) );
NAND4_X1 U859 ( .A1(n1098), .A2(n1089), .A3(n1196), .A4(n1197), .ZN(n1193) );
NAND2_X1 U860 ( .A1(KEYINPUT47), .A2(n1198), .ZN(n1197) );
NAND2_X1 U861 ( .A1(n1199), .A2(n1200), .ZN(n1196) );
INV_X1 U862 ( .A(KEYINPUT47), .ZN(n1200) );
NAND2_X1 U863 ( .A1(n1201), .A2(n1107), .ZN(n1199) );
NOR2_X1 U864 ( .A1(n1171), .A2(n1202), .ZN(G57) );
XOR2_X1 U865 ( .A(n1203), .B(n1204), .Z(n1202) );
XNOR2_X1 U866 ( .A(n1205), .B(n1206), .ZN(n1204) );
NAND2_X1 U867 ( .A1(KEYINPUT51), .A2(n1207), .ZN(n1205) );
NAND2_X1 U868 ( .A1(n1208), .A2(n1209), .ZN(n1203) );
NAND2_X1 U869 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND2_X1 U870 ( .A1(n1212), .A2(n1213), .ZN(n1208) );
INV_X1 U871 ( .A(n1211), .ZN(n1213) );
XNOR2_X1 U872 ( .A(n1214), .B(n1215), .ZN(n1211) );
NAND2_X1 U873 ( .A1(KEYINPUT1), .A2(n1216), .ZN(n1214) );
XNOR2_X1 U874 ( .A(n1210), .B(KEYINPUT58), .ZN(n1212) );
NOR2_X1 U875 ( .A1(n1176), .A2(n1139), .ZN(n1210) );
NOR2_X1 U876 ( .A1(n1217), .A2(n1218), .ZN(G54) );
XOR2_X1 U877 ( .A(KEYINPUT32), .B(n1219), .Z(n1218) );
NOR2_X1 U878 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
XNOR2_X1 U879 ( .A(G953), .B(KEYINPUT39), .ZN(n1220) );
XOR2_X1 U880 ( .A(n1222), .B(n1223), .Z(n1217) );
XNOR2_X1 U881 ( .A(n1224), .B(n1155), .ZN(n1223) );
XOR2_X1 U882 ( .A(n1225), .B(n1226), .Z(n1222) );
NOR2_X1 U883 ( .A1(KEYINPUT53), .A2(n1154), .ZN(n1226) );
XOR2_X1 U884 ( .A(n1227), .B(n1228), .Z(n1225) );
NOR2_X1 U885 ( .A1(KEYINPUT60), .A2(n1229), .ZN(n1228) );
NAND3_X1 U886 ( .A1(n1230), .A2(n1081), .A3(G469), .ZN(n1227) );
XNOR2_X1 U887 ( .A(KEYINPUT9), .B(n1231), .ZN(n1230) );
NOR2_X1 U888 ( .A1(n1171), .A2(n1232), .ZN(G51) );
XOR2_X1 U889 ( .A(n1233), .B(n1234), .Z(n1232) );
XOR2_X1 U890 ( .A(n1235), .B(n1236), .Z(n1234) );
NOR2_X1 U891 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XOR2_X1 U892 ( .A(n1239), .B(KEYINPUT57), .Z(n1238) );
NAND2_X1 U893 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NOR2_X1 U894 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
XOR2_X1 U895 ( .A(KEYINPUT10), .B(n1242), .Z(n1240) );
NAND2_X1 U896 ( .A1(n1181), .A2(n1243), .ZN(n1235) );
INV_X1 U897 ( .A(n1176), .ZN(n1181) );
NAND2_X1 U898 ( .A1(G902), .A2(n1081), .ZN(n1176) );
NAND2_X1 U899 ( .A1(n1170), .A2(n1147), .ZN(n1081) );
AND2_X1 U900 ( .A1(n1244), .A2(n1245), .ZN(n1147) );
NOR4_X1 U901 ( .A1(n1246), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1245) );
NOR4_X1 U902 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1244) );
INV_X1 U903 ( .A(n1254), .ZN(n1252) );
AND4_X1 U904 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1170) );
NOR4_X1 U905 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1076), .ZN(n1258) );
NOR3_X1 U906 ( .A1(n1198), .A2(n1262), .A3(n1114), .ZN(n1076) );
INV_X1 U907 ( .A(n1263), .ZN(n1260) );
NOR2_X1 U908 ( .A1(n1264), .A2(n1265), .ZN(n1257) );
NOR4_X1 U909 ( .A1(n1266), .A2(n1267), .A3(n1268), .A4(n1114), .ZN(n1265) );
INV_X1 U910 ( .A(KEYINPUT46), .ZN(n1266) );
NOR2_X1 U911 ( .A1(KEYINPUT46), .A2(n1269), .ZN(n1264) );
NAND2_X1 U912 ( .A1(n1098), .A2(n1270), .ZN(n1256) );
NAND2_X1 U913 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND3_X1 U914 ( .A1(n1273), .A2(n1274), .A3(n1089), .ZN(n1272) );
OR2_X1 U915 ( .A1(n1275), .A2(KEYINPUT14), .ZN(n1274) );
NAND2_X1 U916 ( .A1(KEYINPUT14), .A2(n1276), .ZN(n1273) );
NAND3_X1 U917 ( .A1(n1277), .A2(n1278), .A3(n1104), .ZN(n1276) );
NAND2_X1 U918 ( .A1(n1116), .A2(n1279), .ZN(n1271) );
NAND3_X1 U919 ( .A1(n1100), .A2(n1275), .A3(n1115), .ZN(n1255) );
NOR2_X1 U920 ( .A1(n1221), .A2(n1083), .ZN(n1171) );
XOR2_X1 U921 ( .A(G952), .B(KEYINPUT0), .Z(n1221) );
XOR2_X1 U922 ( .A(G146), .B(n1253), .Z(G48) );
AND3_X1 U923 ( .A1(n1098), .A2(n1280), .A3(n1281), .ZN(n1253) );
XNOR2_X1 U924 ( .A(G143), .B(n1254), .ZN(G45) );
NAND3_X1 U925 ( .A1(n1268), .A2(n1116), .A3(n1281), .ZN(n1254) );
XNOR2_X1 U926 ( .A(n1282), .B(n1250), .ZN(G42) );
AND3_X1 U927 ( .A1(n1115), .A2(n1098), .A3(n1283), .ZN(n1250) );
XOR2_X1 U928 ( .A(n1251), .B(n1284), .Z(G39) );
XOR2_X1 U929 ( .A(KEYINPUT56), .B(G137), .Z(n1284) );
AND3_X1 U930 ( .A1(n1100), .A2(n1280), .A3(n1283), .ZN(n1251) );
XOR2_X1 U931 ( .A(G134), .B(n1249), .Z(G36) );
AND3_X1 U932 ( .A1(n1116), .A2(n1099), .A3(n1283), .ZN(n1249) );
XOR2_X1 U933 ( .A(G131), .B(n1248), .Z(G33) );
AND3_X1 U934 ( .A1(n1098), .A2(n1116), .A3(n1283), .ZN(n1248) );
AND4_X1 U935 ( .A1(n1104), .A2(n1285), .A3(n1091), .A4(n1092), .ZN(n1283) );
XOR2_X1 U936 ( .A(G128), .B(n1247), .Z(G30) );
AND3_X1 U937 ( .A1(n1280), .A2(n1099), .A3(n1281), .ZN(n1247) );
NOR3_X1 U938 ( .A1(n1278), .A2(n1286), .A3(n1107), .ZN(n1281) );
INV_X1 U939 ( .A(n1104), .ZN(n1107) );
NAND2_X1 U940 ( .A1(n1287), .A2(n1288), .ZN(G3) );
NAND2_X1 U941 ( .A1(n1261), .A2(n1207), .ZN(n1288) );
XOR2_X1 U942 ( .A(KEYINPUT17), .B(n1289), .Z(n1287) );
NOR2_X1 U943 ( .A1(n1261), .A2(n1207), .ZN(n1289) );
AND3_X1 U944 ( .A1(n1116), .A2(n1275), .A3(n1100), .ZN(n1261) );
XOR2_X1 U945 ( .A(G125), .B(n1246), .Z(G27) );
AND4_X1 U946 ( .A1(n1115), .A2(n1098), .A3(n1290), .A4(n1096), .ZN(n1246) );
NOR2_X1 U947 ( .A1(n1286), .A2(n1278), .ZN(n1290) );
INV_X1 U948 ( .A(n1117), .ZN(n1278) );
INV_X1 U949 ( .A(n1285), .ZN(n1286) );
NAND2_X1 U950 ( .A1(n1118), .A2(n1291), .ZN(n1285) );
NAND3_X1 U951 ( .A1(G902), .A2(n1292), .A3(n1150), .ZN(n1291) );
NOR2_X1 U952 ( .A1(n1083), .A2(G900), .ZN(n1150) );
XNOR2_X1 U953 ( .A(G122), .B(n1269), .ZN(G24) );
NAND3_X1 U954 ( .A1(n1279), .A2(n1089), .A3(n1268), .ZN(n1269) );
NOR2_X1 U955 ( .A1(n1293), .A2(n1143), .ZN(n1268) );
INV_X1 U956 ( .A(n1114), .ZN(n1089) );
NAND2_X1 U957 ( .A1(n1135), .A2(n1121), .ZN(n1114) );
XNOR2_X1 U958 ( .A(G119), .B(n1263), .ZN(G21) );
NAND3_X1 U959 ( .A1(n1280), .A2(n1279), .A3(n1100), .ZN(n1263) );
NOR2_X1 U960 ( .A1(n1121), .A2(n1135), .ZN(n1280) );
INV_X1 U961 ( .A(n1294), .ZN(n1121) );
XOR2_X1 U962 ( .A(G116), .B(n1259), .Z(G18) );
AND3_X1 U963 ( .A1(n1279), .A2(n1099), .A3(n1116), .ZN(n1259) );
INV_X1 U964 ( .A(n1262), .ZN(n1099) );
NAND2_X1 U965 ( .A1(n1293), .A2(n1295), .ZN(n1262) );
NAND3_X1 U966 ( .A1(n1296), .A2(n1297), .A3(n1298), .ZN(G15) );
NAND2_X1 U967 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
NAND2_X1 U968 ( .A1(n1301), .A2(n1302), .ZN(n1297) );
INV_X1 U969 ( .A(KEYINPUT33), .ZN(n1302) );
NAND2_X1 U970 ( .A1(n1303), .A2(G113), .ZN(n1301) );
XNOR2_X1 U971 ( .A(n1299), .B(KEYINPUT16), .ZN(n1303) );
NAND2_X1 U972 ( .A1(KEYINPUT33), .A2(n1304), .ZN(n1296) );
NAND2_X1 U973 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
OR3_X1 U974 ( .A1(n1300), .A2(n1299), .A3(KEYINPUT16), .ZN(n1306) );
INV_X1 U975 ( .A(G113), .ZN(n1300) );
NAND2_X1 U976 ( .A1(KEYINPUT16), .A2(n1299), .ZN(n1305) );
AND3_X1 U977 ( .A1(n1279), .A2(n1307), .A3(n1098), .ZN(n1299) );
NOR2_X1 U978 ( .A1(n1293), .A2(n1295), .ZN(n1098) );
XOR2_X1 U979 ( .A(KEYINPUT20), .B(n1116), .Z(n1307) );
NOR2_X1 U980 ( .A1(n1294), .A2(n1135), .ZN(n1116) );
INV_X1 U981 ( .A(n1267), .ZN(n1279) );
NAND2_X1 U982 ( .A1(n1096), .A2(n1201), .ZN(n1267) );
NOR2_X1 U983 ( .A1(n1308), .A2(n1105), .ZN(n1096) );
XNOR2_X1 U984 ( .A(G110), .B(n1309), .ZN(G12) );
NAND3_X1 U985 ( .A1(n1275), .A2(n1310), .A3(n1115), .ZN(n1309) );
AND2_X1 U986 ( .A1(n1135), .A2(n1294), .ZN(n1115) );
XOR2_X1 U987 ( .A(n1311), .B(n1175), .Z(n1294) );
NAND2_X1 U988 ( .A1(G217), .A2(n1312), .ZN(n1175) );
NAND2_X1 U989 ( .A1(n1177), .A2(n1231), .ZN(n1311) );
XOR2_X1 U990 ( .A(n1313), .B(n1314), .Z(n1177) );
XOR2_X1 U991 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U992 ( .A(G125), .B(n1317), .ZN(n1316) );
XNOR2_X1 U993 ( .A(n1282), .B(G137), .ZN(n1315) );
XOR2_X1 U994 ( .A(n1318), .B(n1319), .Z(n1313) );
XOR2_X1 U995 ( .A(n1320), .B(n1321), .Z(n1318) );
NOR2_X1 U996 ( .A1(G110), .A2(n1322), .ZN(n1321) );
XNOR2_X1 U997 ( .A(KEYINPUT40), .B(KEYINPUT24), .ZN(n1322) );
NAND2_X1 U998 ( .A1(G221), .A2(n1323), .ZN(n1320) );
XNOR2_X1 U999 ( .A(n1324), .B(n1139), .ZN(n1135) );
INV_X1 U1000 ( .A(G472), .ZN(n1139) );
OR2_X1 U1001 ( .A1(n1140), .A2(G902), .ZN(n1324) );
XNOR2_X1 U1002 ( .A(n1325), .B(n1326), .ZN(n1140) );
XOR2_X1 U1003 ( .A(n1206), .B(n1327), .Z(n1326) );
XNOR2_X1 U1004 ( .A(G101), .B(KEYINPUT29), .ZN(n1327) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1328), .ZN(n1206) );
XOR2_X1 U1006 ( .A(n1215), .B(n1216), .Z(n1325) );
XOR2_X1 U1007 ( .A(n1329), .B(n1330), .Z(n1216) );
XNOR2_X1 U1008 ( .A(KEYINPUT38), .B(n1317), .ZN(n1330) );
XNOR2_X1 U1009 ( .A(G116), .B(G113), .ZN(n1329) );
XOR2_X1 U1010 ( .A(n1331), .B(n1154), .Z(n1215) );
XOR2_X1 U1011 ( .A(KEYINPUT5), .B(n1100), .Z(n1310) );
AND2_X1 U1012 ( .A1(n1143), .A2(n1293), .ZN(n1100) );
NAND2_X1 U1013 ( .A1(n1332), .A2(n1333), .ZN(n1293) );
NAND2_X1 U1014 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
INV_X1 U1015 ( .A(G475), .ZN(n1335) );
XNOR2_X1 U1016 ( .A(n1131), .B(KEYINPUT34), .ZN(n1334) );
NAND2_X1 U1017 ( .A1(n1336), .A2(G475), .ZN(n1332) );
XOR2_X1 U1018 ( .A(KEYINPUT59), .B(n1131), .Z(n1336) );
NOR2_X1 U1019 ( .A1(n1185), .A2(G902), .ZN(n1131) );
XNOR2_X1 U1020 ( .A(n1337), .B(n1338), .ZN(n1185) );
XNOR2_X1 U1021 ( .A(G113), .B(n1339), .ZN(n1338) );
XNOR2_X1 U1022 ( .A(KEYINPUT48), .B(KEYINPUT13), .ZN(n1339) );
XOR2_X1 U1023 ( .A(n1340), .B(n1341), .Z(n1337) );
XNOR2_X1 U1024 ( .A(n1342), .B(n1190), .ZN(n1340) );
NAND2_X1 U1025 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
NAND2_X1 U1026 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
XOR2_X1 U1027 ( .A(KEYINPUT43), .B(n1347), .Z(n1343) );
NOR2_X1 U1028 ( .A1(n1345), .A2(n1346), .ZN(n1347) );
XOR2_X1 U1029 ( .A(n1348), .B(n1349), .Z(n1346) );
XNOR2_X1 U1030 ( .A(n1350), .B(G131), .ZN(n1349) );
NAND2_X1 U1031 ( .A1(G214), .A2(n1328), .ZN(n1348) );
NOR2_X1 U1032 ( .A1(G953), .A2(G237), .ZN(n1328) );
XNOR2_X1 U1033 ( .A(n1351), .B(n1352), .ZN(n1345) );
XNOR2_X1 U1034 ( .A(n1353), .B(KEYINPUT28), .ZN(n1352) );
NAND2_X1 U1035 ( .A1(n1354), .A2(KEYINPUT11), .ZN(n1353) );
XOR2_X1 U1036 ( .A(n1355), .B(G125), .Z(n1354) );
NAND2_X1 U1037 ( .A1(KEYINPUT52), .A2(n1282), .ZN(n1355) );
INV_X1 U1038 ( .A(n1295), .ZN(n1143) );
XNOR2_X1 U1039 ( .A(n1356), .B(G478), .ZN(n1295) );
NAND2_X1 U1040 ( .A1(n1180), .A2(n1231), .ZN(n1356) );
XOR2_X1 U1041 ( .A(n1357), .B(n1358), .Z(n1180) );
XOR2_X1 U1042 ( .A(n1359), .B(n1360), .Z(n1358) );
AND2_X1 U1043 ( .A1(G217), .A2(n1323), .ZN(n1360) );
AND2_X1 U1044 ( .A1(G234), .A2(n1083), .ZN(n1323) );
NOR2_X1 U1045 ( .A1(KEYINPUT54), .A2(G134), .ZN(n1359) );
XOR2_X1 U1046 ( .A(n1361), .B(n1362), .Z(n1357) );
NOR2_X1 U1047 ( .A1(KEYINPUT63), .A2(n1363), .ZN(n1362) );
XOR2_X1 U1048 ( .A(n1364), .B(n1341), .Z(n1363) );
XNOR2_X1 U1049 ( .A(G107), .B(G116), .ZN(n1364) );
XNOR2_X1 U1050 ( .A(G128), .B(G143), .ZN(n1361) );
INV_X1 U1051 ( .A(n1198), .ZN(n1275) );
NAND2_X1 U1052 ( .A1(n1104), .A2(n1201), .ZN(n1198) );
AND2_X1 U1053 ( .A1(n1117), .A2(n1277), .ZN(n1201) );
NAND2_X1 U1054 ( .A1(n1118), .A2(n1365), .ZN(n1277) );
NAND4_X1 U1055 ( .A1(G953), .A2(G902), .A3(n1292), .A4(n1167), .ZN(n1365) );
INV_X1 U1056 ( .A(G898), .ZN(n1167) );
NAND3_X1 U1057 ( .A1(n1292), .A2(n1083), .A3(G952), .ZN(n1118) );
NAND2_X1 U1058 ( .A1(G237), .A2(G234), .ZN(n1292) );
NOR2_X1 U1059 ( .A1(n1092), .A2(n1113), .ZN(n1117) );
INV_X1 U1060 ( .A(n1091), .ZN(n1113) );
NAND2_X1 U1061 ( .A1(G214), .A2(n1366), .ZN(n1091) );
NAND3_X1 U1062 ( .A1(n1367), .A2(n1368), .A3(n1369), .ZN(n1092) );
NAND2_X1 U1063 ( .A1(n1129), .A2(n1370), .ZN(n1369) );
OR3_X1 U1064 ( .A1(n1370), .A2(n1129), .A3(KEYINPUT18), .ZN(n1368) );
AND2_X1 U1065 ( .A1(n1371), .A2(n1231), .ZN(n1129) );
XOR2_X1 U1066 ( .A(n1233), .B(n1372), .Z(n1371) );
XNOR2_X1 U1067 ( .A(n1242), .B(n1241), .ZN(n1372) );
XNOR2_X1 U1068 ( .A(n1331), .B(G125), .ZN(n1241) );
XOR2_X1 U1069 ( .A(n1373), .B(n1319), .Z(n1331) );
XOR2_X1 U1070 ( .A(G128), .B(n1351), .Z(n1319) );
NAND2_X1 U1071 ( .A1(KEYINPUT37), .A2(n1350), .ZN(n1373) );
INV_X1 U1072 ( .A(G143), .ZN(n1350) );
NAND2_X1 U1073 ( .A1(G224), .A2(n1083), .ZN(n1242) );
XOR2_X1 U1074 ( .A(n1168), .B(n1374), .Z(n1233) );
NOR2_X1 U1075 ( .A1(KEYINPUT50), .A2(n1169), .ZN(n1374) );
XNOR2_X1 U1076 ( .A(n1375), .B(n1376), .ZN(n1169) );
XNOR2_X1 U1077 ( .A(n1207), .B(n1377), .ZN(n1376) );
NOR2_X1 U1078 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
XOR2_X1 U1079 ( .A(n1380), .B(KEYINPUT62), .Z(n1379) );
NAND2_X1 U1080 ( .A1(n1381), .A2(G113), .ZN(n1380) );
NOR2_X1 U1081 ( .A1(G113), .A2(n1381), .ZN(n1378) );
XOR2_X1 U1082 ( .A(n1382), .B(G116), .Z(n1381) );
NAND2_X1 U1083 ( .A1(KEYINPUT7), .A2(n1317), .ZN(n1382) );
INV_X1 U1084 ( .A(G119), .ZN(n1317) );
INV_X1 U1085 ( .A(G101), .ZN(n1207) );
NAND2_X1 U1086 ( .A1(n1383), .A2(n1384), .ZN(n1375) );
NAND2_X1 U1087 ( .A1(KEYINPUT25), .A2(n1385), .ZN(n1384) );
OR3_X1 U1088 ( .A1(n1190), .A2(G107), .A3(KEYINPUT25), .ZN(n1383) );
XOR2_X1 U1089 ( .A(n1386), .B(n1341), .Z(n1168) );
XOR2_X1 U1090 ( .A(G122), .B(KEYINPUT23), .Z(n1341) );
NAND2_X1 U1091 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
INV_X1 U1092 ( .A(G110), .ZN(n1388) );
XNOR2_X1 U1093 ( .A(KEYINPUT41), .B(KEYINPUT19), .ZN(n1387) );
NAND2_X1 U1094 ( .A1(KEYINPUT31), .A2(n1128), .ZN(n1370) );
NAND2_X1 U1095 ( .A1(KEYINPUT18), .A2(n1243), .ZN(n1367) );
INV_X1 U1096 ( .A(n1128), .ZN(n1243) );
NAND2_X1 U1097 ( .A1(G210), .A2(n1366), .ZN(n1128) );
NAND2_X1 U1098 ( .A1(n1389), .A2(n1231), .ZN(n1366) );
INV_X1 U1099 ( .A(G237), .ZN(n1389) );
NOR2_X1 U1100 ( .A1(n1106), .A2(n1105), .ZN(n1104) );
AND2_X1 U1101 ( .A1(G221), .A2(n1312), .ZN(n1105) );
NAND2_X1 U1102 ( .A1(G234), .A2(n1231), .ZN(n1312) );
INV_X1 U1103 ( .A(n1308), .ZN(n1106) );
XOR2_X1 U1104 ( .A(n1142), .B(n1390), .Z(n1308) );
NOR2_X1 U1105 ( .A1(KEYINPUT4), .A2(n1141), .ZN(n1390) );
INV_X1 U1106 ( .A(G469), .ZN(n1141) );
AND2_X1 U1107 ( .A1(n1391), .A2(n1231), .ZN(n1142) );
INV_X1 U1108 ( .A(G902), .ZN(n1231) );
XNOR2_X1 U1109 ( .A(n1392), .B(n1393), .ZN(n1391) );
INV_X1 U1110 ( .A(n1224), .ZN(n1393) );
XNOR2_X1 U1111 ( .A(n1394), .B(n1395), .ZN(n1224) );
XNOR2_X1 U1112 ( .A(n1282), .B(G110), .ZN(n1395) );
INV_X1 U1113 ( .A(G140), .ZN(n1282) );
NAND2_X1 U1114 ( .A1(G227), .A2(n1083), .ZN(n1394) );
INV_X1 U1115 ( .A(G953), .ZN(n1083) );
NOR3_X1 U1116 ( .A1(n1396), .A2(KEYINPUT12), .A3(n1397), .ZN(n1392) );
NOR2_X1 U1117 ( .A1(n1154), .A2(n1398), .ZN(n1397) );
XOR2_X1 U1118 ( .A(n1399), .B(KEYINPUT8), .Z(n1396) );
NAND2_X1 U1119 ( .A1(n1398), .A2(n1154), .ZN(n1399) );
XNOR2_X1 U1120 ( .A(G131), .B(n1400), .ZN(n1154) );
XOR2_X1 U1121 ( .A(G137), .B(G134), .Z(n1400) );
XNOR2_X1 U1122 ( .A(n1229), .B(n1155), .ZN(n1398) );
XOR2_X1 U1123 ( .A(G128), .B(n1401), .Z(n1155) );
NOR2_X1 U1124 ( .A1(KEYINPUT35), .A2(n1402), .ZN(n1401) );
XOR2_X1 U1125 ( .A(n1403), .B(n1404), .Z(n1402) );
XOR2_X1 U1126 ( .A(KEYINPUT61), .B(KEYINPUT36), .Z(n1404) );
XNOR2_X1 U1127 ( .A(G143), .B(n1351), .ZN(n1403) );
XOR2_X1 U1128 ( .A(G146), .B(KEYINPUT27), .Z(n1351) );
XNOR2_X1 U1129 ( .A(G101), .B(n1385), .ZN(n1229) );
XNOR2_X1 U1130 ( .A(n1190), .B(n1075), .ZN(n1385) );
INV_X1 U1131 ( .A(G107), .ZN(n1075) );
INV_X1 U1132 ( .A(G104), .ZN(n1190) );
endmodule


