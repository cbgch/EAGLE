//Key = 0100011001110010010010010111110011110101100001000110010110001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327;

XOR2_X1 U725 ( .A(G107), .B(n1004), .Z(G9) );
NOR2_X1 U726 ( .A1(n1005), .A2(n1006), .ZN(G75) );
NOR3_X1 U727 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1006) );
NAND3_X1 U728 ( .A1(n1010), .A2(n1011), .A3(n1012), .ZN(n1007) );
NAND2_X1 U729 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U730 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NAND4_X1 U731 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
NAND2_X1 U732 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U733 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND3_X1 U734 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1019) );
NAND2_X1 U735 ( .A1(n1023), .A2(n1028), .ZN(n1026) );
NAND2_X1 U736 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND2_X1 U737 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
INV_X1 U738 ( .A(n1033), .ZN(n1029) );
NAND2_X1 U739 ( .A1(n1024), .A2(n1034), .ZN(n1025) );
NAND2_X1 U740 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND3_X1 U741 ( .A1(G214), .A2(n1037), .A3(n1038), .ZN(n1036) );
NAND4_X1 U742 ( .A1(n1039), .A2(n1027), .A3(n1024), .A4(n1040), .ZN(n1015) );
NAND2_X1 U743 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR2_X1 U744 ( .A1(n1043), .A2(n1044), .ZN(n1039) );
NOR2_X1 U745 ( .A1(n1045), .A2(n1018), .ZN(n1044) );
NOR2_X1 U746 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U747 ( .A1(n1041), .A2(n1042), .ZN(n1046) );
INV_X1 U748 ( .A(KEYINPUT48), .ZN(n1042) );
NOR2_X1 U749 ( .A1(n1048), .A2(n1049), .ZN(n1043) );
NOR2_X1 U750 ( .A1(n1050), .A2(n1041), .ZN(n1049) );
NOR2_X1 U751 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U752 ( .A1(n1053), .A2(G953), .A3(G952), .ZN(n1005) );
INV_X1 U753 ( .A(n1010), .ZN(n1053) );
NAND3_X1 U754 ( .A1(n1054), .A2(n1031), .A3(n1055), .ZN(n1010) );
NOR3_X1 U755 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
XNOR2_X1 U756 ( .A(G478), .B(n1059), .ZN(n1058) );
NOR2_X1 U757 ( .A1(KEYINPUT46), .A2(n1060), .ZN(n1059) );
XOR2_X1 U758 ( .A(KEYINPUT12), .B(n1061), .Z(n1060) );
NOR3_X1 U759 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1057) );
NOR2_X1 U760 ( .A1(KEYINPUT55), .A2(n1065), .ZN(n1064) );
XNOR2_X1 U761 ( .A(KEYINPUT30), .B(G475), .ZN(n1065) );
NOR3_X1 U762 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1063) );
INV_X1 U763 ( .A(KEYINPUT55), .ZN(n1066) );
AND2_X1 U764 ( .A1(n1068), .A2(n1067), .ZN(n1062) );
OR2_X1 U765 ( .A1(KEYINPUT62), .A2(n1069), .ZN(n1068) );
XNOR2_X1 U766 ( .A(KEYINPUT30), .B(n1070), .ZN(n1069) );
XNOR2_X1 U767 ( .A(n1032), .B(KEYINPUT26), .ZN(n1056) );
XOR2_X1 U768 ( .A(n1071), .B(KEYINPUT17), .Z(n1054) );
NAND3_X1 U769 ( .A1(n1072), .A2(n1018), .A3(n1023), .ZN(n1071) );
XNOR2_X1 U770 ( .A(KEYINPUT20), .B(n1027), .ZN(n1072) );
NAND3_X1 U771 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(G72) );
INV_X1 U772 ( .A(n1076), .ZN(n1075) );
NAND2_X1 U773 ( .A1(n1077), .A2(n1011), .ZN(n1074) );
NAND2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1080), .A2(n1008), .ZN(n1079) );
NAND2_X1 U776 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
INV_X1 U778 ( .A(KEYINPUT33), .ZN(n1084) );
NAND3_X1 U779 ( .A1(n1085), .A2(n1086), .A3(KEYINPUT33), .ZN(n1081) );
INV_X1 U780 ( .A(KEYINPUT36), .ZN(n1086) );
NAND2_X1 U781 ( .A1(n1083), .A2(n1087), .ZN(n1078) );
NAND2_X1 U782 ( .A1(n1088), .A2(G953), .ZN(n1073) );
XNOR2_X1 U783 ( .A(n1083), .B(G227), .ZN(n1088) );
NOR2_X1 U784 ( .A1(n1085), .A2(KEYINPUT36), .ZN(n1083) );
XOR2_X1 U785 ( .A(n1089), .B(n1090), .Z(n1085) );
XOR2_X1 U786 ( .A(n1091), .B(n1092), .Z(n1090) );
XNOR2_X1 U787 ( .A(G125), .B(KEYINPUT1), .ZN(n1092) );
NAND2_X1 U788 ( .A1(KEYINPUT5), .A2(n1093), .ZN(n1091) );
XOR2_X1 U789 ( .A(n1094), .B(n1095), .Z(n1089) );
NAND2_X1 U790 ( .A1(n1096), .A2(n1097), .ZN(G69) );
NAND2_X1 U791 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U792 ( .A1(G953), .A2(n1100), .ZN(n1099) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1100) );
NAND2_X1 U794 ( .A1(n1101), .A2(n1102), .ZN(n1096) );
NAND2_X1 U795 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND2_X1 U796 ( .A1(G953), .A2(n1105), .ZN(n1104) );
INV_X1 U797 ( .A(n1098), .ZN(n1101) );
XNOR2_X1 U798 ( .A(n1106), .B(n1107), .ZN(n1098) );
NOR2_X1 U799 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XNOR2_X1 U800 ( .A(G953), .B(KEYINPUT53), .ZN(n1109) );
NAND2_X1 U801 ( .A1(n1110), .A2(n1103), .ZN(n1106) );
INV_X1 U802 ( .A(n1111), .ZN(n1103) );
XOR2_X1 U803 ( .A(n1112), .B(n1113), .Z(n1110) );
NOR2_X1 U804 ( .A1(KEYINPUT13), .A2(n1114), .ZN(n1112) );
NOR2_X1 U805 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U806 ( .A(n1117), .B(KEYINPUT60), .Z(n1116) );
NAND2_X1 U807 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U808 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
XNOR2_X1 U809 ( .A(n1120), .B(KEYINPUT24), .ZN(n1119) );
NOR2_X1 U810 ( .A1(n1121), .A2(n1122), .ZN(G66) );
XOR2_X1 U811 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U812 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR2_X1 U813 ( .A1(n1121), .A2(n1127), .ZN(G63) );
XOR2_X1 U814 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U815 ( .A1(n1130), .A2(n1126), .ZN(n1128) );
INV_X1 U816 ( .A(G478), .ZN(n1130) );
NOR2_X1 U817 ( .A1(n1121), .A2(n1131), .ZN(G60) );
XOR2_X1 U818 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U819 ( .A1(n1070), .A2(n1126), .ZN(n1132) );
XOR2_X1 U820 ( .A(G104), .B(n1134), .Z(G6) );
NOR2_X1 U821 ( .A1(n1121), .A2(n1135), .ZN(G57) );
XOR2_X1 U822 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U823 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U824 ( .A1(n1140), .A2(n1126), .ZN(n1138) );
XNOR2_X1 U825 ( .A(G101), .B(n1141), .ZN(n1136) );
NOR2_X1 U826 ( .A1(n1121), .A2(n1142), .ZN(G54) );
XOR2_X1 U827 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U828 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR3_X1 U829 ( .A1(n1126), .A2(KEYINPUT58), .A3(n1147), .ZN(n1146) );
XOR2_X1 U830 ( .A(n1148), .B(n1149), .Z(n1143) );
XNOR2_X1 U831 ( .A(n1093), .B(G110), .ZN(n1149) );
NOR2_X1 U832 ( .A1(n1121), .A2(n1150), .ZN(G51) );
XOR2_X1 U833 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U834 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U835 ( .A(KEYINPUT61), .B(n1155), .Z(n1154) );
NOR2_X1 U836 ( .A1(KEYINPUT3), .A2(n1156), .ZN(n1155) );
NOR2_X1 U837 ( .A1(n1157), .A2(n1126), .ZN(n1153) );
NAND2_X1 U838 ( .A1(n1158), .A2(n1159), .ZN(n1126) );
NAND2_X1 U839 ( .A1(n1108), .A2(n1087), .ZN(n1159) );
INV_X1 U840 ( .A(n1008), .ZN(n1087) );
NAND4_X1 U841 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1008) );
NOR4_X1 U842 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1163) );
INV_X1 U843 ( .A(n1168), .ZN(n1167) );
AND2_X1 U844 ( .A1(n1169), .A2(n1170), .ZN(n1162) );
NAND2_X1 U845 ( .A1(n1023), .A2(n1171), .ZN(n1161) );
NAND2_X1 U846 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NAND2_X1 U847 ( .A1(KEYINPUT0), .A2(n1174), .ZN(n1173) );
NAND2_X1 U848 ( .A1(n1175), .A2(n1017), .ZN(n1172) );
NAND2_X1 U849 ( .A1(n1176), .A2(n1177), .ZN(n1160) );
INV_X1 U850 ( .A(KEYINPUT0), .ZN(n1177) );
INV_X1 U851 ( .A(n1009), .ZN(n1108) );
NAND2_X1 U852 ( .A1(n1178), .A2(n1179), .ZN(n1009) );
NOR4_X1 U853 ( .A1(n1180), .A2(n1181), .A3(n1004), .A4(n1182), .ZN(n1179) );
INV_X1 U854 ( .A(n1183), .ZN(n1182) );
AND3_X1 U855 ( .A1(n1052), .A2(n1024), .A3(n1184), .ZN(n1004) );
INV_X1 U856 ( .A(n1185), .ZN(n1181) );
NOR4_X1 U857 ( .A1(n1186), .A2(n1187), .A3(n1134), .A4(n1188), .ZN(n1178) );
NOR2_X1 U858 ( .A1(n1189), .A2(n1035), .ZN(n1188) );
XOR2_X1 U859 ( .A(n1190), .B(KEYINPUT42), .Z(n1189) );
AND3_X1 U860 ( .A1(n1184), .A2(n1024), .A3(n1051), .ZN(n1134) );
INV_X1 U861 ( .A(n1191), .ZN(n1187) );
INV_X1 U862 ( .A(n1192), .ZN(n1186) );
XNOR2_X1 U863 ( .A(KEYINPUT4), .B(n1193), .ZN(n1158) );
XNOR2_X1 U864 ( .A(n1194), .B(n1195), .ZN(n1151) );
NOR2_X1 U865 ( .A1(KEYINPUT7), .A2(n1196), .ZN(n1195) );
NOR2_X1 U866 ( .A1(n1011), .A2(G952), .ZN(n1121) );
XOR2_X1 U867 ( .A(n1170), .B(n1197), .Z(G48) );
NAND2_X1 U868 ( .A1(KEYINPUT14), .A2(G146), .ZN(n1197) );
NAND3_X1 U869 ( .A1(n1051), .A2(n1198), .A3(n1175), .ZN(n1170) );
XNOR2_X1 U870 ( .A(G143), .B(n1169), .ZN(G45) );
NAND3_X1 U871 ( .A1(n1199), .A2(n1033), .A3(n1200), .ZN(n1169) );
NOR3_X1 U872 ( .A1(n1035), .A2(n1201), .A3(n1202), .ZN(n1200) );
XNOR2_X1 U873 ( .A(G140), .B(n1168), .ZN(G42) );
NAND3_X1 U874 ( .A1(n1199), .A2(n1023), .A3(n1203), .ZN(n1168) );
XNOR2_X1 U875 ( .A(n1204), .B(n1205), .ZN(G39) );
NOR4_X1 U876 ( .A1(KEYINPUT52), .A2(n1041), .A3(n1047), .A4(n1206), .ZN(n1205) );
XNOR2_X1 U877 ( .A(G134), .B(n1207), .ZN(G36) );
NAND2_X1 U878 ( .A1(KEYINPUT11), .A2(n1165), .ZN(n1207) );
AND4_X1 U879 ( .A1(n1199), .A2(n1033), .A3(n1023), .A4(n1052), .ZN(n1165) );
INV_X1 U880 ( .A(n1041), .ZN(n1023) );
XOR2_X1 U881 ( .A(n1208), .B(n1176), .Z(G33) );
NOR2_X1 U882 ( .A1(n1174), .A2(n1041), .ZN(n1176) );
NAND2_X1 U883 ( .A1(n1038), .A2(n1209), .ZN(n1041) );
NAND2_X1 U884 ( .A1(G214), .A2(n1037), .ZN(n1209) );
NAND3_X1 U885 ( .A1(n1051), .A2(n1033), .A3(n1199), .ZN(n1174) );
XNOR2_X1 U886 ( .A(G131), .B(KEYINPUT28), .ZN(n1208) );
XOR2_X1 U887 ( .A(n1164), .B(n1210), .Z(G30) );
NOR2_X1 U888 ( .A1(KEYINPUT38), .A2(n1211), .ZN(n1210) );
AND3_X1 U889 ( .A1(n1052), .A2(n1198), .A3(n1175), .ZN(n1164) );
INV_X1 U890 ( .A(n1206), .ZN(n1175) );
NAND3_X1 U891 ( .A1(n1032), .A2(n1212), .A3(n1199), .ZN(n1206) );
AND3_X1 U892 ( .A1(n1213), .A2(n1018), .A3(n1021), .ZN(n1199) );
XNOR2_X1 U893 ( .A(n1214), .B(n1215), .ZN(G3) );
NOR2_X1 U894 ( .A1(n1035), .A2(n1190), .ZN(n1215) );
NAND3_X1 U895 ( .A1(n1033), .A2(n1017), .A3(n1216), .ZN(n1190) );
NOR3_X1 U896 ( .A1(n1027), .A2(n1048), .A3(n1217), .ZN(n1216) );
XOR2_X1 U897 ( .A(G125), .B(n1166), .Z(G27) );
AND3_X1 U898 ( .A1(n1218), .A2(n1213), .A3(n1203), .ZN(n1166) );
AND3_X1 U899 ( .A1(n1031), .A2(n1032), .A3(n1051), .ZN(n1203) );
NAND2_X1 U900 ( .A1(n1219), .A2(n1220), .ZN(n1213) );
NAND3_X1 U901 ( .A1(G902), .A2(n1014), .A3(n1076), .ZN(n1220) );
NOR2_X1 U902 ( .A1(G900), .A2(n1011), .ZN(n1076) );
XNOR2_X1 U903 ( .A(G122), .B(n1191), .ZN(G24) );
NAND4_X1 U904 ( .A1(n1221), .A2(n1024), .A3(n1222), .A4(n1223), .ZN(n1191) );
NOR2_X1 U905 ( .A1(n1212), .A2(n1032), .ZN(n1024) );
XNOR2_X1 U906 ( .A(n1224), .B(n1225), .ZN(G21) );
NOR2_X1 U907 ( .A1(KEYINPUT51), .A2(n1183), .ZN(n1225) );
NAND4_X1 U908 ( .A1(n1221), .A2(n1017), .A3(n1032), .A4(n1212), .ZN(n1183) );
XNOR2_X1 U909 ( .A(G116), .B(n1185), .ZN(G18) );
NAND3_X1 U910 ( .A1(n1221), .A2(n1052), .A3(n1033), .ZN(n1185) );
NOR2_X1 U911 ( .A1(n1223), .A2(n1202), .ZN(n1052) );
INV_X1 U912 ( .A(n1222), .ZN(n1202) );
XNOR2_X1 U913 ( .A(n1226), .B(KEYINPUT43), .ZN(n1222) );
XOR2_X1 U914 ( .A(n1227), .B(G113), .Z(G15) );
NAND2_X1 U915 ( .A1(KEYINPUT35), .A2(n1192), .ZN(n1227) );
NAND3_X1 U916 ( .A1(n1033), .A2(n1221), .A3(n1051), .ZN(n1192) );
AND2_X1 U917 ( .A1(n1226), .A2(n1223), .ZN(n1051) );
AND2_X1 U918 ( .A1(n1218), .A2(n1228), .ZN(n1221) );
NOR3_X1 U919 ( .A1(n1035), .A2(n1048), .A3(n1021), .ZN(n1218) );
NOR2_X1 U920 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
XNOR2_X1 U921 ( .A(G110), .B(n1229), .ZN(G12) );
NAND2_X1 U922 ( .A1(KEYINPUT9), .A2(n1180), .ZN(n1229) );
AND4_X1 U923 ( .A1(n1017), .A2(n1184), .A3(n1031), .A4(n1032), .ZN(n1180) );
XOR2_X1 U924 ( .A(n1230), .B(n1125), .Z(n1032) );
NAND2_X1 U925 ( .A1(G217), .A2(n1231), .ZN(n1125) );
NAND2_X1 U926 ( .A1(n1232), .A2(n1193), .ZN(n1230) );
XOR2_X1 U927 ( .A(n1123), .B(KEYINPUT32), .Z(n1232) );
XOR2_X1 U928 ( .A(n1233), .B(n1234), .Z(n1123) );
XOR2_X1 U929 ( .A(n1235), .B(n1236), .Z(n1234) );
NAND2_X1 U930 ( .A1(KEYINPUT34), .A2(n1237), .ZN(n1236) );
NAND2_X1 U931 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
OR2_X1 U932 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
XOR2_X1 U933 ( .A(n1242), .B(KEYINPUT21), .Z(n1238) );
NAND2_X1 U934 ( .A1(n1241), .A2(n1240), .ZN(n1242) );
XNOR2_X1 U935 ( .A(n1243), .B(n1244), .ZN(n1240) );
XNOR2_X1 U936 ( .A(KEYINPUT31), .B(n1211), .ZN(n1244) );
INV_X1 U937 ( .A(G128), .ZN(n1211) );
XNOR2_X1 U938 ( .A(G110), .B(G119), .ZN(n1243) );
XNOR2_X1 U939 ( .A(n1245), .B(n1246), .ZN(n1241) );
NOR2_X1 U940 ( .A1(KEYINPUT57), .A2(G125), .ZN(n1246) );
XNOR2_X1 U941 ( .A(G140), .B(G146), .ZN(n1245) );
NAND2_X1 U942 ( .A1(n1247), .A2(G221), .ZN(n1235) );
XNOR2_X1 U943 ( .A(G137), .B(KEYINPUT44), .ZN(n1233) );
INV_X1 U944 ( .A(n1212), .ZN(n1031) );
XOR2_X1 U945 ( .A(n1248), .B(n1140), .Z(n1212) );
INV_X1 U946 ( .A(G472), .ZN(n1140) );
NAND2_X1 U947 ( .A1(n1193), .A2(n1249), .ZN(n1248) );
NAND2_X1 U948 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NAND2_X1 U949 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
XOR2_X1 U950 ( .A(KEYINPUT23), .B(n1139), .Z(n1253) );
XNOR2_X1 U951 ( .A(n1254), .B(n1214), .ZN(n1252) );
XOR2_X1 U952 ( .A(n1255), .B(KEYINPUT8), .Z(n1250) );
NAND2_X1 U953 ( .A1(n1256), .A2(n1139), .ZN(n1255) );
XNOR2_X1 U954 ( .A(n1257), .B(n1258), .ZN(n1139) );
XNOR2_X1 U955 ( .A(n1156), .B(n1259), .ZN(n1258) );
XOR2_X1 U956 ( .A(n1260), .B(n1261), .Z(n1257) );
NAND2_X1 U957 ( .A1(n1262), .A2(n1263), .ZN(n1260) );
NAND2_X1 U958 ( .A1(G116), .A2(n1224), .ZN(n1263) );
XOR2_X1 U959 ( .A(KEYINPUT56), .B(n1264), .Z(n1262) );
NOR2_X1 U960 ( .A1(G116), .A2(n1224), .ZN(n1264) );
INV_X1 U961 ( .A(G119), .ZN(n1224) );
XNOR2_X1 U962 ( .A(G101), .B(n1254), .ZN(n1256) );
NAND2_X1 U963 ( .A1(KEYINPUT10), .A2(n1265), .ZN(n1254) );
INV_X1 U964 ( .A(n1141), .ZN(n1265) );
NAND3_X1 U965 ( .A1(n1266), .A2(n1011), .A3(G210), .ZN(n1141) );
NOR4_X1 U966 ( .A1(n1035), .A2(n1027), .A3(n1217), .A4(n1048), .ZN(n1184) );
INV_X1 U967 ( .A(n1018), .ZN(n1048) );
NAND2_X1 U968 ( .A1(G221), .A2(n1231), .ZN(n1018) );
NAND2_X1 U969 ( .A1(G234), .A2(n1267), .ZN(n1231) );
INV_X1 U970 ( .A(n1228), .ZN(n1217) );
NAND2_X1 U971 ( .A1(n1219), .A2(n1268), .ZN(n1228) );
NAND3_X1 U972 ( .A1(G902), .A2(n1014), .A3(n1111), .ZN(n1268) );
NOR2_X1 U973 ( .A1(n1011), .A2(G898), .ZN(n1111) );
NAND3_X1 U974 ( .A1(n1014), .A2(n1011), .A3(G952), .ZN(n1219) );
NAND2_X1 U975 ( .A1(G234), .A2(n1269), .ZN(n1014) );
XNOR2_X1 U976 ( .A(KEYINPUT54), .B(n1266), .ZN(n1269) );
INV_X1 U977 ( .A(n1021), .ZN(n1027) );
XOR2_X1 U978 ( .A(n1270), .B(n1147), .Z(n1021) );
INV_X1 U979 ( .A(G469), .ZN(n1147) );
NAND2_X1 U980 ( .A1(n1271), .A2(n1193), .ZN(n1270) );
XOR2_X1 U981 ( .A(n1145), .B(n1272), .Z(n1271) );
NOR2_X1 U982 ( .A1(KEYINPUT16), .A2(n1273), .ZN(n1272) );
XOR2_X1 U983 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U984 ( .A(n1148), .B(n1276), .ZN(n1275) );
NOR2_X1 U985 ( .A1(G140), .A2(KEYINPUT15), .ZN(n1276) );
NAND2_X1 U986 ( .A1(G227), .A2(n1011), .ZN(n1148) );
XNOR2_X1 U987 ( .A(G110), .B(KEYINPUT6), .ZN(n1274) );
XNOR2_X1 U988 ( .A(n1277), .B(n1120), .ZN(n1145) );
XNOR2_X1 U989 ( .A(n1261), .B(n1095), .ZN(n1277) );
XNOR2_X1 U990 ( .A(n1278), .B(n1279), .ZN(n1095) );
XNOR2_X1 U991 ( .A(G146), .B(n1280), .ZN(n1279) );
XNOR2_X1 U992 ( .A(KEYINPUT50), .B(KEYINPUT41), .ZN(n1280) );
XOR2_X1 U993 ( .A(n1281), .B(n1282), .Z(n1278) );
NOR2_X1 U994 ( .A1(G128), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U995 ( .A(KEYINPUT27), .B(KEYINPUT22), .ZN(n1283) );
XNOR2_X1 U996 ( .A(G131), .B(G143), .ZN(n1281) );
NOR2_X1 U997 ( .A1(KEYINPUT59), .A2(n1094), .ZN(n1261) );
XNOR2_X1 U998 ( .A(G134), .B(n1284), .ZN(n1094) );
XNOR2_X1 U999 ( .A(KEYINPUT40), .B(n1204), .ZN(n1284) );
INV_X1 U1000 ( .A(G137), .ZN(n1204) );
INV_X1 U1001 ( .A(n1198), .ZN(n1035) );
NOR2_X1 U1002 ( .A1(n1038), .A2(n1285), .ZN(n1198) );
AND2_X1 U1003 ( .A1(G214), .A2(n1037), .ZN(n1285) );
XNOR2_X1 U1004 ( .A(n1286), .B(n1157), .ZN(n1038) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1037), .ZN(n1157) );
NAND2_X1 U1006 ( .A1(n1267), .A2(n1266), .ZN(n1037) );
XNOR2_X1 U1007 ( .A(n1193), .B(KEYINPUT45), .ZN(n1267) );
NAND2_X1 U1008 ( .A1(n1287), .A2(n1193), .ZN(n1286) );
INV_X1 U1009 ( .A(G902), .ZN(n1193) );
XNOR2_X1 U1010 ( .A(n1288), .B(n1196), .ZN(n1287) );
XOR2_X1 U1011 ( .A(n1289), .B(n1290), .Z(n1196) );
XNOR2_X1 U1012 ( .A(KEYINPUT25), .B(n1120), .ZN(n1290) );
XOR2_X1 U1013 ( .A(n1214), .B(n1291), .Z(n1120) );
XOR2_X1 U1014 ( .A(G107), .B(G104), .Z(n1291) );
INV_X1 U1015 ( .A(G101), .ZN(n1214) );
XOR2_X1 U1016 ( .A(n1118), .B(n1113), .Z(n1289) );
XNOR2_X1 U1017 ( .A(n1292), .B(n1293), .ZN(n1113) );
NOR2_X1 U1018 ( .A1(KEYINPUT19), .A2(n1294), .ZN(n1293) );
INV_X1 U1019 ( .A(G110), .ZN(n1292) );
XOR2_X1 U1020 ( .A(n1295), .B(G113), .Z(n1118) );
NAND2_X1 U1021 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
NAND2_X1 U1022 ( .A1(G119), .A2(n1298), .ZN(n1297) );
XOR2_X1 U1023 ( .A(KEYINPUT29), .B(n1299), .Z(n1296) );
NOR2_X1 U1024 ( .A1(G119), .A2(n1298), .ZN(n1299) );
INV_X1 U1025 ( .A(G116), .ZN(n1298) );
NOR2_X1 U1026 ( .A1(KEYINPUT2), .A2(n1300), .ZN(n1288) );
XNOR2_X1 U1027 ( .A(n1156), .B(n1194), .ZN(n1300) );
XOR2_X1 U1028 ( .A(G125), .B(n1301), .Z(n1194) );
NOR2_X1 U1029 ( .A1(G953), .A2(n1105), .ZN(n1301) );
INV_X1 U1030 ( .A(G224), .ZN(n1105) );
XOR2_X1 U1031 ( .A(n1302), .B(n1303), .Z(n1156) );
XNOR2_X1 U1032 ( .A(KEYINPUT37), .B(n1304), .ZN(n1303) );
XNOR2_X1 U1033 ( .A(G128), .B(G143), .ZN(n1302) );
INV_X1 U1034 ( .A(n1047), .ZN(n1017) );
NAND2_X1 U1035 ( .A1(n1201), .A2(n1226), .ZN(n1047) );
XNOR2_X1 U1036 ( .A(n1061), .B(G478), .ZN(n1226) );
NOR2_X1 U1037 ( .A1(n1129), .A2(G902), .ZN(n1061) );
XNOR2_X1 U1038 ( .A(n1305), .B(n1306), .ZN(n1129) );
XOR2_X1 U1039 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U1040 ( .A(G107), .B(n1309), .ZN(n1308) );
NOR2_X1 U1041 ( .A1(G143), .A2(KEYINPUT18), .ZN(n1309) );
NAND2_X1 U1042 ( .A1(G217), .A2(n1247), .ZN(n1307) );
AND2_X1 U1043 ( .A1(G234), .A2(n1011), .ZN(n1247) );
XOR2_X1 U1044 ( .A(n1310), .B(n1311), .Z(n1305) );
XNOR2_X1 U1045 ( .A(n1294), .B(G116), .ZN(n1311) );
XNOR2_X1 U1046 ( .A(G134), .B(G128), .ZN(n1310) );
INV_X1 U1047 ( .A(n1223), .ZN(n1201) );
XOR2_X1 U1048 ( .A(n1067), .B(n1312), .Z(n1223) );
XNOR2_X1 U1049 ( .A(KEYINPUT47), .B(n1070), .ZN(n1312) );
INV_X1 U1050 ( .A(G475), .ZN(n1070) );
NOR2_X1 U1051 ( .A1(n1133), .A2(G902), .ZN(n1067) );
XNOR2_X1 U1052 ( .A(n1313), .B(n1314), .ZN(n1133) );
XOR2_X1 U1053 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1054 ( .A(n1294), .B(G104), .ZN(n1316) );
INV_X1 U1055 ( .A(G122), .ZN(n1294) );
AND3_X1 U1056 ( .A1(G214), .A2(n1011), .A3(n1266), .ZN(n1315) );
INV_X1 U1057 ( .A(G237), .ZN(n1266) );
INV_X1 U1058 ( .A(G953), .ZN(n1011) );
XNOR2_X1 U1059 ( .A(n1259), .B(n1317), .ZN(n1313) );
XOR2_X1 U1060 ( .A(n1318), .B(n1319), .Z(n1317) );
NAND2_X1 U1061 ( .A1(KEYINPUT39), .A2(G143), .ZN(n1319) );
NAND2_X1 U1062 ( .A1(n1320), .A2(n1321), .ZN(n1318) );
NAND2_X1 U1063 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NAND2_X1 U1064 ( .A1(KEYINPUT49), .A2(n1324), .ZN(n1323) );
NAND2_X1 U1065 ( .A1(KEYINPUT63), .A2(G146), .ZN(n1324) );
NAND2_X1 U1066 ( .A1(n1325), .A2(n1304), .ZN(n1320) );
INV_X1 U1067 ( .A(G146), .ZN(n1304) );
NAND2_X1 U1068 ( .A1(KEYINPUT63), .A2(n1326), .ZN(n1325) );
NAND2_X1 U1069 ( .A1(KEYINPUT49), .A2(n1327), .ZN(n1326) );
INV_X1 U1070 ( .A(n1322), .ZN(n1327) );
XOR2_X1 U1071 ( .A(G125), .B(n1093), .Z(n1322) );
INV_X1 U1072 ( .A(G140), .ZN(n1093) );
XOR2_X1 U1073 ( .A(G113), .B(G131), .Z(n1259) );
endmodule


