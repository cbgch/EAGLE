//Key = 1110011110111000110000010010011011110101100011100011001011101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409;

XNOR2_X1 U770 ( .A(G107), .B(n1070), .ZN(G9) );
NOR2_X1 U771 ( .A1(n1071), .A2(n1072), .ZN(G75) );
NOR4_X1 U772 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1072) );
NAND4_X1 U773 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1073) );
NAND4_X1 U774 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1078) );
NAND2_X1 U775 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NAND3_X1 U776 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NAND3_X1 U777 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1088) );
INV_X1 U778 ( .A(n1093), .ZN(n1091) );
NAND2_X1 U779 ( .A1(n1094), .A2(n1095), .ZN(n1090) );
INV_X1 U780 ( .A(KEYINPUT51), .ZN(n1095) );
NAND2_X1 U781 ( .A1(n1094), .A2(n1096), .ZN(n1085) );
NAND3_X1 U782 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
NAND2_X1 U783 ( .A1(n1087), .A2(n1100), .ZN(n1099) );
NAND2_X1 U784 ( .A1(KEYINPUT34), .A2(n1089), .ZN(n1100) );
NAND4_X1 U785 ( .A1(KEYINPUT51), .A2(n1101), .A3(n1102), .A4(n1089), .ZN(n1097) );
NAND2_X1 U786 ( .A1(n1089), .A2(n1103), .ZN(n1077) );
NAND2_X1 U787 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND3_X1 U788 ( .A1(n1087), .A2(n1094), .A3(n1106), .ZN(n1105) );
NOR3_X1 U789 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1106) );
NOR2_X1 U790 ( .A1(n1110), .A2(n1084), .ZN(n1109) );
AND2_X1 U791 ( .A1(n1082), .A2(KEYINPUT34), .ZN(n1110) );
NOR2_X1 U792 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
NAND2_X1 U793 ( .A1(n1113), .A2(n1084), .ZN(n1104) );
XOR2_X1 U794 ( .A(n1114), .B(KEYINPUT63), .Z(n1113) );
NAND4_X1 U795 ( .A1(n1081), .A2(n1087), .A3(n1115), .A4(n1094), .ZN(n1114) );
INV_X1 U796 ( .A(n1107), .ZN(n1081) );
AND3_X1 U797 ( .A1(n1079), .A2(n1080), .A3(n1116), .ZN(n1071) );
NAND4_X1 U798 ( .A1(n1117), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1079) );
NOR4_X1 U799 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1120) );
NOR2_X1 U800 ( .A1(G478), .A2(n1125), .ZN(n1124) );
AND3_X1 U801 ( .A1(n1125), .A2(n1126), .A3(G478), .ZN(n1123) );
INV_X1 U802 ( .A(KEYINPUT41), .ZN(n1125) );
NAND3_X1 U803 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1121) );
XOR2_X1 U804 ( .A(KEYINPUT56), .B(n1130), .Z(n1128) );
NOR3_X1 U805 ( .A1(n1112), .A2(n1131), .A3(n1132), .ZN(n1119) );
INV_X1 U806 ( .A(n1133), .ZN(n1132) );
NAND2_X1 U807 ( .A1(G475), .A2(n1134), .ZN(n1118) );
XNOR2_X1 U808 ( .A(KEYINPUT5), .B(n1135), .ZN(n1117) );
XOR2_X1 U809 ( .A(n1136), .B(n1137), .Z(G72) );
XOR2_X1 U810 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U811 ( .A1(G953), .A2(n1140), .ZN(n1139) );
NAND2_X1 U812 ( .A1(G900), .A2(G227), .ZN(n1140) );
NAND2_X1 U813 ( .A1(n1141), .A2(n1142), .ZN(n1138) );
NAND2_X1 U814 ( .A1(G953), .A2(n1143), .ZN(n1142) );
XOR2_X1 U815 ( .A(n1144), .B(n1145), .Z(n1141) );
XNOR2_X1 U816 ( .A(n1146), .B(n1147), .ZN(n1145) );
NOR2_X1 U817 ( .A1(KEYINPUT31), .A2(n1148), .ZN(n1147) );
XOR2_X1 U818 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U819 ( .A(n1151), .B(G137), .Z(n1150) );
INV_X1 U820 ( .A(G131), .ZN(n1151) );
NAND2_X1 U821 ( .A1(KEYINPUT32), .A2(n1152), .ZN(n1149) );
NAND2_X1 U822 ( .A1(n1153), .A2(n1154), .ZN(n1144) );
NAND2_X1 U823 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND2_X1 U824 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
NAND2_X1 U825 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NAND2_X1 U826 ( .A1(n1161), .A2(G146), .ZN(n1153) );
XOR2_X1 U827 ( .A(G140), .B(G125), .Z(n1161) );
AND2_X1 U828 ( .A1(n1075), .A2(n1080), .ZN(n1136) );
XOR2_X1 U829 ( .A(n1162), .B(n1163), .Z(G69) );
NOR2_X1 U830 ( .A1(n1080), .A2(n1164), .ZN(n1163) );
XOR2_X1 U831 ( .A(KEYINPUT59), .B(n1165), .Z(n1164) );
NOR2_X1 U832 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XNOR2_X1 U833 ( .A(G224), .B(KEYINPUT27), .ZN(n1166) );
NAND3_X1 U834 ( .A1(n1168), .A2(n1169), .A3(KEYINPUT58), .ZN(n1162) );
NAND3_X1 U835 ( .A1(n1170), .A2(n1080), .A3(n1171), .ZN(n1169) );
INV_X1 U836 ( .A(n1172), .ZN(n1171) );
XOR2_X1 U837 ( .A(KEYINPUT26), .B(n1173), .Z(n1168) );
NOR2_X1 U838 ( .A1(n1174), .A2(n1170), .ZN(n1173) );
NAND2_X1 U839 ( .A1(n1175), .A2(n1176), .ZN(n1170) );
NAND2_X1 U840 ( .A1(n1177), .A2(G953), .ZN(n1176) );
XOR2_X1 U841 ( .A(n1167), .B(KEYINPUT25), .Z(n1177) );
XOR2_X1 U842 ( .A(n1178), .B(n1179), .Z(n1175) );
NOR2_X1 U843 ( .A1(KEYINPUT52), .A2(n1180), .ZN(n1179) );
XNOR2_X1 U844 ( .A(n1181), .B(n1182), .ZN(n1180) );
XOR2_X1 U845 ( .A(G113), .B(n1183), .Z(n1182) );
NOR2_X1 U846 ( .A1(KEYINPUT53), .A2(n1184), .ZN(n1183) );
XNOR2_X1 U847 ( .A(G101), .B(n1185), .ZN(n1184) );
XNOR2_X1 U848 ( .A(G122), .B(G110), .ZN(n1178) );
NOR2_X1 U849 ( .A1(n1172), .A2(G953), .ZN(n1174) );
NOR2_X1 U850 ( .A1(n1074), .A2(n1186), .ZN(n1172) );
NOR2_X1 U851 ( .A1(n1187), .A2(n1188), .ZN(G66) );
XOR2_X1 U852 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U853 ( .A1(n1191), .A2(n1192), .ZN(n1189) );
NOR2_X1 U854 ( .A1(n1187), .A2(n1193), .ZN(G63) );
XOR2_X1 U855 ( .A(n1194), .B(n1195), .Z(n1193) );
NAND3_X1 U856 ( .A1(n1196), .A2(G478), .A3(KEYINPUT35), .ZN(n1194) );
NOR2_X1 U857 ( .A1(n1187), .A2(n1197), .ZN(G60) );
XOR2_X1 U858 ( .A(n1198), .B(n1199), .Z(n1197) );
XOR2_X1 U859 ( .A(KEYINPUT28), .B(n1200), .Z(n1199) );
AND2_X1 U860 ( .A1(G475), .A2(n1196), .ZN(n1200) );
XNOR2_X1 U861 ( .A(G104), .B(n1201), .ZN(G6) );
NOR2_X1 U862 ( .A1(n1187), .A2(n1202), .ZN(G57) );
XOR2_X1 U863 ( .A(n1203), .B(n1204), .Z(n1202) );
XNOR2_X1 U864 ( .A(n1205), .B(n1206), .ZN(n1204) );
NOR3_X1 U865 ( .A1(n1192), .A2(KEYINPUT36), .A3(n1207), .ZN(n1206) );
INV_X1 U866 ( .A(G472), .ZN(n1207) );
NAND2_X1 U867 ( .A1(KEYINPUT44), .A2(G101), .ZN(n1205) );
XOR2_X1 U868 ( .A(n1208), .B(n1209), .Z(n1203) );
NAND2_X1 U869 ( .A1(n1210), .A2(n1211), .ZN(n1208) );
NAND3_X1 U870 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1211) );
XOR2_X1 U871 ( .A(KEYINPUT46), .B(n1215), .Z(n1210) );
NOR2_X1 U872 ( .A1(n1216), .A2(n1214), .ZN(n1215) );
XNOR2_X1 U873 ( .A(n1181), .B(n1217), .ZN(n1214) );
AND2_X1 U874 ( .A1(n1212), .A2(n1213), .ZN(n1216) );
NAND2_X1 U875 ( .A1(n1218), .A2(n1219), .ZN(n1213) );
XOR2_X1 U876 ( .A(KEYINPUT42), .B(n1220), .Z(n1218) );
OR2_X1 U877 ( .A1(n1220), .A2(n1219), .ZN(n1212) );
NOR2_X1 U878 ( .A1(n1187), .A2(n1221), .ZN(G54) );
XOR2_X1 U879 ( .A(n1222), .B(n1223), .Z(n1221) );
XOR2_X1 U880 ( .A(n1224), .B(n1225), .Z(n1223) );
NAND2_X1 U881 ( .A1(n1226), .A2(n1227), .ZN(n1224) );
XOR2_X1 U882 ( .A(KEYINPUT40), .B(n1228), .Z(n1226) );
XOR2_X1 U883 ( .A(n1229), .B(n1230), .Z(n1222) );
XNOR2_X1 U884 ( .A(n1231), .B(n1232), .ZN(n1230) );
AND2_X1 U885 ( .A1(G469), .A2(n1196), .ZN(n1232) );
NAND2_X1 U886 ( .A1(KEYINPUT2), .A2(n1233), .ZN(n1229) );
NOR4_X1 U887 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(G51) );
NOR2_X1 U888 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
XOR2_X1 U889 ( .A(KEYINPUT12), .B(n1240), .Z(n1238) );
NOR2_X1 U890 ( .A1(n1240), .A2(n1241), .ZN(n1236) );
INV_X1 U891 ( .A(n1239), .ZN(n1241) );
XOR2_X1 U892 ( .A(n1242), .B(n1243), .Z(n1239) );
NAND3_X1 U893 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1242) );
NAND2_X1 U894 ( .A1(n1247), .A2(n1248), .ZN(n1245) );
INV_X1 U895 ( .A(KEYINPUT0), .ZN(n1248) );
XOR2_X1 U896 ( .A(n1249), .B(n1250), .Z(n1247) );
NOR2_X1 U897 ( .A1(G125), .A2(n1219), .ZN(n1250) );
NAND2_X1 U898 ( .A1(KEYINPUT0), .A2(n1251), .ZN(n1244) );
AND2_X1 U899 ( .A1(n1196), .A2(G210), .ZN(n1240) );
INV_X1 U900 ( .A(n1192), .ZN(n1196) );
NAND2_X1 U901 ( .A1(G902), .A2(n1252), .ZN(n1192) );
OR3_X1 U902 ( .A1(n1076), .A2(n1075), .A3(n1074), .ZN(n1252) );
NAND4_X1 U903 ( .A1(n1201), .A2(n1253), .A3(n1254), .A4(n1070), .ZN(n1074) );
NAND3_X1 U904 ( .A1(n1094), .A2(n1255), .A3(n1115), .ZN(n1070) );
NAND3_X1 U905 ( .A1(n1255), .A2(n1256), .A3(n1082), .ZN(n1253) );
NAND3_X1 U906 ( .A1(n1094), .A2(n1255), .A3(n1111), .ZN(n1201) );
NAND4_X1 U907 ( .A1(n1257), .A2(n1258), .A3(n1259), .A4(n1260), .ZN(n1075) );
AND4_X1 U908 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1260) );
NOR2_X1 U909 ( .A1(n1265), .A2(n1266), .ZN(n1259) );
INV_X1 U910 ( .A(n1267), .ZN(n1265) );
XNOR2_X1 U911 ( .A(n1186), .B(KEYINPUT54), .ZN(n1076) );
NAND4_X1 U912 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1186) );
NOR3_X1 U913 ( .A1(n1272), .A2(n1080), .A3(n1116), .ZN(n1235) );
INV_X1 U914 ( .A(G952), .ZN(n1116) );
AND2_X1 U915 ( .A1(n1272), .A2(n1187), .ZN(n1234) );
NOR2_X1 U916 ( .A1(n1080), .A2(G952), .ZN(n1187) );
INV_X1 U917 ( .A(KEYINPUT18), .ZN(n1272) );
XOR2_X1 U918 ( .A(n1156), .B(n1261), .Z(G48) );
NAND3_X1 U919 ( .A1(n1111), .A2(n1273), .A3(n1274), .ZN(n1261) );
XOR2_X1 U920 ( .A(n1275), .B(n1257), .Z(G45) );
NAND4_X1 U921 ( .A1(n1274), .A2(n1093), .A3(n1276), .A4(n1277), .ZN(n1257) );
XOR2_X1 U922 ( .A(n1160), .B(n1264), .Z(G42) );
NAND3_X1 U923 ( .A1(n1111), .A2(n1256), .A3(n1278), .ZN(n1264) );
XOR2_X1 U924 ( .A(n1258), .B(n1279), .Z(G39) );
NOR2_X1 U925 ( .A1(G137), .A2(KEYINPUT47), .ZN(n1279) );
NAND3_X1 U926 ( .A1(n1273), .A2(n1082), .A3(n1278), .ZN(n1258) );
NAND2_X1 U927 ( .A1(n1280), .A2(n1281), .ZN(G36) );
OR2_X1 U928 ( .A1(n1263), .A2(G134), .ZN(n1281) );
XOR2_X1 U929 ( .A(n1282), .B(KEYINPUT4), .Z(n1280) );
NAND2_X1 U930 ( .A1(G134), .A2(n1263), .ZN(n1282) );
NAND3_X1 U931 ( .A1(n1093), .A2(n1115), .A3(n1278), .ZN(n1263) );
XOR2_X1 U932 ( .A(G131), .B(n1266), .Z(G33) );
AND3_X1 U933 ( .A1(n1111), .A2(n1093), .A3(n1278), .ZN(n1266) );
NOR3_X1 U934 ( .A1(n1283), .A2(n1112), .A3(n1098), .ZN(n1278) );
OR3_X1 U935 ( .A1(n1102), .A2(n1101), .A3(n1284), .ZN(n1098) );
XOR2_X1 U936 ( .A(n1285), .B(n1267), .Z(G30) );
NAND3_X1 U937 ( .A1(n1273), .A2(n1115), .A3(n1274), .ZN(n1267) );
AND2_X1 U938 ( .A1(n1286), .A2(n1287), .ZN(n1274) );
XNOR2_X1 U939 ( .A(G101), .B(n1288), .ZN(G3) );
NAND2_X1 U940 ( .A1(KEYINPUT62), .A2(n1289), .ZN(n1288) );
INV_X1 U941 ( .A(n1254), .ZN(n1289) );
NAND3_X1 U942 ( .A1(n1093), .A2(n1255), .A3(n1082), .ZN(n1254) );
AND2_X1 U943 ( .A1(n1286), .A2(n1290), .ZN(n1255) );
XOR2_X1 U944 ( .A(n1159), .B(n1262), .Z(G27) );
NAND4_X1 U945 ( .A1(n1087), .A2(n1256), .A3(n1111), .A4(n1291), .ZN(n1262) );
NOR3_X1 U946 ( .A1(n1283), .A2(n1089), .A3(n1112), .ZN(n1291) );
INV_X1 U947 ( .A(n1287), .ZN(n1283) );
NAND2_X1 U948 ( .A1(n1107), .A2(n1292), .ZN(n1287) );
NAND4_X1 U949 ( .A1(G953), .A2(G902), .A3(n1293), .A4(n1143), .ZN(n1292) );
INV_X1 U950 ( .A(G900), .ZN(n1143) );
XNOR2_X1 U951 ( .A(G122), .B(n1268), .ZN(G24) );
NAND4_X1 U952 ( .A1(n1294), .A2(n1094), .A3(n1276), .A4(n1277), .ZN(n1268) );
AND2_X1 U953 ( .A1(n1129), .A2(n1295), .ZN(n1094) );
XOR2_X1 U954 ( .A(n1296), .B(n1127), .Z(n1295) );
XOR2_X1 U955 ( .A(n1269), .B(n1297), .Z(G21) );
NAND2_X1 U956 ( .A1(KEYINPUT23), .A2(G119), .ZN(n1297) );
NAND3_X1 U957 ( .A1(n1273), .A2(n1082), .A3(n1294), .ZN(n1269) );
XNOR2_X1 U958 ( .A(G116), .B(n1270), .ZN(G18) );
NAND3_X1 U959 ( .A1(n1093), .A2(n1115), .A3(n1294), .ZN(n1270) );
NOR2_X1 U960 ( .A1(n1277), .A2(n1298), .ZN(n1115) );
NAND2_X1 U961 ( .A1(n1299), .A2(n1300), .ZN(G15) );
OR2_X1 U962 ( .A1(n1271), .A2(G113), .ZN(n1300) );
XOR2_X1 U963 ( .A(n1301), .B(KEYINPUT22), .Z(n1299) );
NAND2_X1 U964 ( .A1(G113), .A2(n1271), .ZN(n1301) );
NAND3_X1 U965 ( .A1(n1111), .A2(n1093), .A3(n1294), .ZN(n1271) );
AND4_X1 U966 ( .A1(n1087), .A2(n1290), .A3(n1084), .A4(n1284), .ZN(n1294) );
INV_X1 U967 ( .A(n1122), .ZN(n1087) );
NAND2_X1 U968 ( .A1(n1102), .A2(n1302), .ZN(n1122) );
NOR2_X1 U969 ( .A1(n1303), .A2(n1127), .ZN(n1093) );
NOR2_X1 U970 ( .A1(n1276), .A2(n1304), .ZN(n1111) );
XNOR2_X1 U971 ( .A(G110), .B(n1305), .ZN(G12) );
NAND3_X1 U972 ( .A1(n1082), .A2(n1286), .A3(n1306), .ZN(n1305) );
NOR3_X1 U973 ( .A1(n1307), .A2(KEYINPUT61), .A3(n1092), .ZN(n1306) );
INV_X1 U974 ( .A(n1256), .ZN(n1092) );
NAND2_X1 U975 ( .A1(n1308), .A2(n1309), .ZN(n1256) );
NAND2_X1 U976 ( .A1(n1273), .A2(n1296), .ZN(n1309) );
INV_X1 U977 ( .A(KEYINPUT37), .ZN(n1296) );
NOR2_X1 U978 ( .A1(n1127), .A2(n1129), .ZN(n1273) );
NAND3_X1 U979 ( .A1(n1303), .A2(n1127), .A3(KEYINPUT37), .ZN(n1308) );
XOR2_X1 U980 ( .A(n1310), .B(G472), .Z(n1127) );
NAND2_X1 U981 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U982 ( .A(n1313), .B(n1314), .Z(n1311) );
XNOR2_X1 U983 ( .A(n1217), .B(n1315), .ZN(n1314) );
XOR2_X1 U984 ( .A(n1316), .B(n1220), .Z(n1315) );
INV_X1 U985 ( .A(n1317), .ZN(n1316) );
XNOR2_X1 U986 ( .A(n1318), .B(KEYINPUT16), .ZN(n1217) );
NAND2_X1 U987 ( .A1(KEYINPUT45), .A2(n1319), .ZN(n1318) );
INV_X1 U988 ( .A(G113), .ZN(n1319) );
XOR2_X1 U989 ( .A(n1320), .B(n1321), .Z(n1313) );
XOR2_X1 U990 ( .A(KEYINPUT7), .B(KEYINPUT49), .Z(n1321) );
XOR2_X1 U991 ( .A(n1219), .B(n1209), .Z(n1320) );
AND3_X1 U992 ( .A1(n1322), .A2(n1080), .A3(G210), .ZN(n1209) );
INV_X1 U993 ( .A(n1129), .ZN(n1303) );
XNOR2_X1 U994 ( .A(n1323), .B(n1191), .ZN(n1129) );
NAND2_X1 U995 ( .A1(G217), .A2(n1324), .ZN(n1191) );
OR2_X1 U996 ( .A1(n1190), .A2(G902), .ZN(n1323) );
XNOR2_X1 U997 ( .A(n1325), .B(n1326), .ZN(n1190) );
XOR2_X1 U998 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U999 ( .A(n1329), .B(n1330), .ZN(n1328) );
NOR2_X1 U1000 ( .A1(KEYINPUT14), .A2(n1331), .ZN(n1330) );
XNOR2_X1 U1001 ( .A(G110), .B(KEYINPUT21), .ZN(n1331) );
NAND2_X1 U1002 ( .A1(n1332), .A2(KEYINPUT1), .ZN(n1329) );
XOR2_X1 U1003 ( .A(n1156), .B(n1333), .Z(n1332) );
NOR2_X1 U1004 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NOR2_X1 U1005 ( .A1(G140), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1006 ( .A(KEYINPUT24), .B(G125), .Z(n1336) );
NOR2_X1 U1007 ( .A1(n1337), .A2(n1338), .ZN(n1327) );
INV_X1 U1008 ( .A(G221), .ZN(n1338) );
XOR2_X1 U1009 ( .A(n1339), .B(n1340), .Z(n1325) );
XOR2_X1 U1010 ( .A(KEYINPUT48), .B(G137), .Z(n1340) );
XOR2_X1 U1011 ( .A(G119), .B(n1285), .Z(n1339) );
XOR2_X1 U1012 ( .A(n1290), .B(KEYINPUT50), .Z(n1307) );
NAND2_X1 U1013 ( .A1(n1107), .A2(n1341), .ZN(n1290) );
NAND4_X1 U1014 ( .A1(G953), .A2(G902), .A3(n1293), .A4(n1167), .ZN(n1341) );
INV_X1 U1015 ( .A(G898), .ZN(n1167) );
NAND3_X1 U1016 ( .A1(n1293), .A2(n1080), .A3(G952), .ZN(n1107) );
NAND2_X1 U1017 ( .A1(G237), .A2(G234), .ZN(n1293) );
NOR4_X1 U1018 ( .A1(n1102), .A2(n1101), .A3(n1112), .A4(n1089), .ZN(n1286) );
INV_X1 U1019 ( .A(n1284), .ZN(n1089) );
NAND2_X1 U1020 ( .A1(n1133), .A2(n1135), .ZN(n1284) );
NAND3_X1 U1021 ( .A1(G210), .A2(n1342), .A3(n1343), .ZN(n1135) );
NAND2_X1 U1022 ( .A1(n1344), .A2(n1312), .ZN(n1342) );
NAND3_X1 U1023 ( .A1(n1345), .A2(n1312), .A3(n1344), .ZN(n1133) );
XNOR2_X1 U1024 ( .A(n1346), .B(n1243), .ZN(n1344) );
XNOR2_X1 U1025 ( .A(n1347), .B(n1348), .ZN(n1243) );
XOR2_X1 U1026 ( .A(n1185), .B(n1349), .Z(n1348) );
XNOR2_X1 U1027 ( .A(G110), .B(KEYINPUT6), .ZN(n1349) );
NAND2_X1 U1028 ( .A1(KEYINPUT60), .A2(n1350), .ZN(n1185) );
XNOR2_X1 U1029 ( .A(G107), .B(n1351), .ZN(n1350) );
NAND2_X1 U1030 ( .A1(KEYINPUT33), .A2(G104), .ZN(n1351) );
XOR2_X1 U1031 ( .A(n1317), .B(n1352), .Z(n1347) );
XOR2_X1 U1032 ( .A(G101), .B(n1181), .Z(n1317) );
XNOR2_X1 U1033 ( .A(G116), .B(G119), .ZN(n1181) );
NAND2_X1 U1034 ( .A1(n1353), .A2(n1246), .ZN(n1346) );
NAND3_X1 U1035 ( .A1(n1249), .A2(n1219), .A3(G125), .ZN(n1246) );
INV_X1 U1036 ( .A(n1251), .ZN(n1353) );
NAND2_X1 U1037 ( .A1(n1354), .A2(n1355), .ZN(n1251) );
NAND2_X1 U1038 ( .A1(n1356), .A2(n1159), .ZN(n1355) );
XOR2_X1 U1039 ( .A(n1219), .B(n1249), .Z(n1356) );
OR3_X1 U1040 ( .A1(n1249), .A2(n1219), .A3(n1159), .ZN(n1354) );
NAND2_X1 U1041 ( .A1(n1357), .A2(n1358), .ZN(n1219) );
NAND2_X1 U1042 ( .A1(n1359), .A2(n1285), .ZN(n1358) );
XOR2_X1 U1043 ( .A(n1360), .B(KEYINPUT13), .Z(n1357) );
OR2_X1 U1044 ( .A1(n1359), .A2(n1285), .ZN(n1360) );
XNOR2_X1 U1045 ( .A(n1361), .B(G143), .ZN(n1359) );
NAND2_X1 U1046 ( .A1(KEYINPUT57), .A2(n1156), .ZN(n1361) );
INV_X1 U1047 ( .A(G146), .ZN(n1156) );
NAND2_X1 U1048 ( .A1(G224), .A2(n1080), .ZN(n1249) );
NAND2_X1 U1049 ( .A1(n1343), .A2(G210), .ZN(n1345) );
XOR2_X1 U1050 ( .A(n1362), .B(KEYINPUT38), .Z(n1343) );
INV_X1 U1051 ( .A(n1084), .ZN(n1112) );
NAND2_X1 U1052 ( .A1(G214), .A2(n1362), .ZN(n1084) );
NAND2_X1 U1053 ( .A1(n1312), .A2(n1322), .ZN(n1362) );
INV_X1 U1054 ( .A(n1302), .ZN(n1101) );
NAND2_X1 U1055 ( .A1(G221), .A2(n1324), .ZN(n1302) );
NAND2_X1 U1056 ( .A1(G234), .A2(n1312), .ZN(n1324) );
XOR2_X1 U1057 ( .A(n1363), .B(G469), .Z(n1102) );
NAND2_X1 U1058 ( .A1(n1364), .A2(n1312), .ZN(n1363) );
XOR2_X1 U1059 ( .A(n1365), .B(n1366), .Z(n1364) );
XOR2_X1 U1060 ( .A(n1231), .B(n1367), .Z(n1366) );
XNOR2_X1 U1061 ( .A(KEYINPUT20), .B(n1368), .ZN(n1367) );
NOR2_X1 U1062 ( .A1(KEYINPUT3), .A2(n1369), .ZN(n1368) );
NOR2_X1 U1063 ( .A1(n1228), .A2(n1370), .ZN(n1369) );
XNOR2_X1 U1064 ( .A(KEYINPUT9), .B(n1227), .ZN(n1370) );
NAND2_X1 U1065 ( .A1(G110), .A2(n1160), .ZN(n1227) );
NOR2_X1 U1066 ( .A1(G110), .A2(n1160), .ZN(n1228) );
INV_X1 U1067 ( .A(G140), .ZN(n1160) );
NAND2_X1 U1068 ( .A1(G227), .A2(n1080), .ZN(n1231) );
XOR2_X1 U1069 ( .A(n1225), .B(n1371), .Z(n1365) );
NOR2_X1 U1070 ( .A1(n1220), .A2(n1372), .ZN(n1371) );
XOR2_X1 U1071 ( .A(KEYINPUT43), .B(KEYINPUT15), .Z(n1372) );
INV_X1 U1072 ( .A(n1233), .ZN(n1220) );
XOR2_X1 U1073 ( .A(n1373), .B(G131), .Z(n1233) );
NAND2_X1 U1074 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
NAND2_X1 U1075 ( .A1(G137), .A2(n1152), .ZN(n1375) );
XOR2_X1 U1076 ( .A(n1376), .B(KEYINPUT55), .Z(n1374) );
OR2_X1 U1077 ( .A1(n1152), .A2(G137), .ZN(n1376) );
XOR2_X1 U1078 ( .A(n1377), .B(n1378), .Z(n1225) );
XOR2_X1 U1079 ( .A(G107), .B(G101), .Z(n1378) );
XNOR2_X1 U1080 ( .A(n1379), .B(n1146), .ZN(n1377) );
XOR2_X1 U1081 ( .A(n1380), .B(KEYINPUT29), .Z(n1146) );
NOR2_X1 U1082 ( .A1(n1276), .A2(n1277), .ZN(n1082) );
INV_X1 U1083 ( .A(n1304), .ZN(n1277) );
NOR2_X1 U1084 ( .A1(n1381), .A2(n1130), .ZN(n1304) );
NOR3_X1 U1085 ( .A1(G475), .A2(G902), .A3(n1198), .ZN(n1130) );
INV_X1 U1086 ( .A(n1382), .ZN(n1198) );
AND2_X1 U1087 ( .A1(G475), .A2(n1134), .ZN(n1381) );
NAND2_X1 U1088 ( .A1(n1382), .A2(n1312), .ZN(n1134) );
XOR2_X1 U1089 ( .A(n1383), .B(n1384), .Z(n1382) );
XOR2_X1 U1090 ( .A(n1385), .B(n1386), .Z(n1384) );
XOR2_X1 U1091 ( .A(KEYINPUT11), .B(G131), .Z(n1386) );
NOR2_X1 U1092 ( .A1(n1387), .A2(n1388), .ZN(n1385) );
XOR2_X1 U1093 ( .A(n1389), .B(KEYINPUT17), .Z(n1388) );
NAND2_X1 U1094 ( .A1(n1275), .A2(n1390), .ZN(n1389) );
NOR2_X1 U1095 ( .A1(n1390), .A2(n1275), .ZN(n1387) );
NAND3_X1 U1096 ( .A1(n1322), .A2(n1080), .A3(G214), .ZN(n1390) );
INV_X1 U1097 ( .A(G237), .ZN(n1322) );
XOR2_X1 U1098 ( .A(n1391), .B(n1379), .Z(n1383) );
XOR2_X1 U1099 ( .A(G104), .B(G146), .Z(n1379) );
XOR2_X1 U1100 ( .A(n1392), .B(n1352), .Z(n1391) );
XOR2_X1 U1101 ( .A(G113), .B(G122), .Z(n1352) );
NAND2_X1 U1102 ( .A1(n1393), .A2(n1394), .ZN(n1392) );
NAND2_X1 U1103 ( .A1(n1395), .A2(n1159), .ZN(n1394) );
INV_X1 U1104 ( .A(G125), .ZN(n1159) );
NAND2_X1 U1105 ( .A1(KEYINPUT39), .A2(G140), .ZN(n1395) );
NAND2_X1 U1106 ( .A1(n1334), .A2(KEYINPUT39), .ZN(n1393) );
INV_X1 U1107 ( .A(n1157), .ZN(n1334) );
NAND2_X1 U1108 ( .A1(G125), .A2(G140), .ZN(n1157) );
INV_X1 U1109 ( .A(n1298), .ZN(n1276) );
NOR2_X1 U1110 ( .A1(n1131), .A2(n1396), .ZN(n1298) );
AND2_X1 U1111 ( .A1(G478), .A2(n1126), .ZN(n1396) );
NOR2_X1 U1112 ( .A1(n1126), .A2(G478), .ZN(n1131) );
NAND2_X1 U1113 ( .A1(n1195), .A2(n1312), .ZN(n1126) );
INV_X1 U1114 ( .A(G902), .ZN(n1312) );
XNOR2_X1 U1115 ( .A(n1397), .B(n1398), .ZN(n1195) );
XOR2_X1 U1116 ( .A(n1399), .B(n1400), .Z(n1398) );
XOR2_X1 U1117 ( .A(G122), .B(G116), .Z(n1400) );
NOR2_X1 U1118 ( .A1(G107), .A2(n1401), .ZN(n1399) );
XNOR2_X1 U1119 ( .A(KEYINPUT30), .B(KEYINPUT19), .ZN(n1401) );
XOR2_X1 U1120 ( .A(n1402), .B(n1403), .Z(n1397) );
NOR2_X1 U1121 ( .A1(n1337), .A2(n1404), .ZN(n1403) );
INV_X1 U1122 ( .A(G217), .ZN(n1404) );
NAND2_X1 U1123 ( .A1(G234), .A2(n1080), .ZN(n1337) );
INV_X1 U1124 ( .A(G953), .ZN(n1080) );
NAND3_X1 U1125 ( .A1(n1405), .A2(n1406), .A3(n1407), .ZN(n1402) );
NAND2_X1 U1126 ( .A1(G134), .A2(n1408), .ZN(n1407) );
NAND3_X1 U1127 ( .A1(n1409), .A2(n1152), .A3(KEYINPUT10), .ZN(n1406) );
INV_X1 U1128 ( .A(G134), .ZN(n1152) );
INV_X1 U1129 ( .A(n1408), .ZN(n1409) );
NAND2_X1 U1130 ( .A1(KEYINPUT8), .A2(n1380), .ZN(n1408) );
OR2_X1 U1131 ( .A1(n1380), .A2(KEYINPUT10), .ZN(n1405) );
XOR2_X1 U1132 ( .A(n1285), .B(n1275), .Z(n1380) );
INV_X1 U1133 ( .A(G143), .ZN(n1275) );
INV_X1 U1134 ( .A(G128), .ZN(n1285) );
endmodule


