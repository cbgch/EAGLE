//Key = 0001000110001111000101000011011010011010110010011010000001101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320;

XNOR2_X1 U738 ( .A(G107), .B(n1012), .ZN(G9) );
NAND4_X1 U739 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(G75) );
NAND3_X1 U740 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1015) );
NOR3_X1 U741 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1019) );
XOR2_X1 U742 ( .A(n1023), .B(KEYINPUT45), .Z(n1020) );
NAND4_X1 U743 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1023) );
XNOR2_X1 U744 ( .A(n1028), .B(n1029), .ZN(n1025) );
XOR2_X1 U745 ( .A(n1030), .B(KEYINPUT60), .Z(n1024) );
NAND3_X1 U746 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
OR2_X1 U747 ( .A1(G478), .A2(KEYINPUT14), .ZN(n1032) );
NAND3_X1 U748 ( .A1(G478), .A2(n1034), .A3(KEYINPUT14), .ZN(n1031) );
XNOR2_X1 U749 ( .A(n1035), .B(n1036), .ZN(n1018) );
XNOR2_X1 U750 ( .A(n1037), .B(n1038), .ZN(n1017) );
NAND2_X1 U751 ( .A1(n1039), .A2(n1040), .ZN(n1014) );
NAND2_X1 U752 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND4_X1 U753 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
NAND2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U756 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U757 ( .A1(n1053), .A2(n1054), .ZN(n1047) );
NAND2_X1 U758 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U759 ( .A1(n1021), .A2(n1057), .ZN(n1056) );
NAND3_X1 U760 ( .A1(n1053), .A2(n1058), .A3(n1049), .ZN(n1041) );
NAND2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND3_X1 U762 ( .A1(n1061), .A2(n1062), .A3(n1044), .ZN(n1060) );
OR2_X1 U763 ( .A1(n1046), .A2(n1043), .ZN(n1062) );
OR3_X1 U764 ( .A1(n1063), .A2(n1064), .A3(n1022), .ZN(n1061) );
NAND2_X1 U765 ( .A1(n1043), .A2(n1065), .ZN(n1059) );
INV_X1 U766 ( .A(n1066), .ZN(n1039) );
INV_X1 U767 ( .A(n1067), .ZN(n1013) );
XOR2_X1 U768 ( .A(n1068), .B(n1069), .Z(G72) );
XOR2_X1 U769 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U771 ( .A1(G953), .A2(n1074), .ZN(n1073) );
XOR2_X1 U772 ( .A(n1075), .B(n1076), .Z(n1072) );
XNOR2_X1 U773 ( .A(n1077), .B(n1078), .ZN(n1076) );
XOR2_X1 U774 ( .A(n1079), .B(n1080), .Z(n1075) );
XOR2_X1 U775 ( .A(KEYINPUT2), .B(G125), .Z(n1080) );
NOR2_X1 U776 ( .A1(G140), .A2(KEYINPUT55), .ZN(n1079) );
NAND2_X1 U777 ( .A1(G953), .A2(n1081), .ZN(n1070) );
NAND2_X1 U778 ( .A1(n1082), .A2(G900), .ZN(n1081) );
XNOR2_X1 U779 ( .A(G227), .B(KEYINPUT58), .ZN(n1082) );
NOR2_X1 U780 ( .A1(n1083), .A2(G953), .ZN(n1068) );
XOR2_X1 U781 ( .A(n1084), .B(n1085), .Z(G69) );
XOR2_X1 U782 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U783 ( .A1(n1088), .A2(n1016), .ZN(n1087) );
NOR2_X1 U784 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U785 ( .A1(n1091), .A2(n1092), .ZN(n1086) );
NAND2_X1 U786 ( .A1(G953), .A2(n1090), .ZN(n1092) );
XOR2_X1 U787 ( .A(n1093), .B(n1094), .Z(n1091) );
XNOR2_X1 U788 ( .A(n1095), .B(n1096), .ZN(n1094) );
NOR2_X1 U789 ( .A1(KEYINPUT17), .A2(n1097), .ZN(n1096) );
XNOR2_X1 U790 ( .A(n1098), .B(n1099), .ZN(n1097) );
NAND2_X1 U791 ( .A1(n1016), .A2(n1100), .ZN(n1084) );
NAND2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XNOR2_X1 U793 ( .A(KEYINPUT7), .B(n1103), .ZN(n1102) );
NOR2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(G66) );
XOR2_X1 U795 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U796 ( .A1(n1029), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U797 ( .A(n1109), .B(KEYINPUT30), .ZN(n1104) );
NOR2_X1 U798 ( .A1(n1109), .A2(n1110), .ZN(G63) );
XOR2_X1 U799 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U800 ( .A1(n1113), .A2(n1108), .ZN(n1111) );
NOR2_X1 U801 ( .A1(n1109), .A2(n1114), .ZN(G60) );
XOR2_X1 U802 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U803 ( .A1(n1117), .A2(n1108), .ZN(n1115) );
XNOR2_X1 U804 ( .A(G104), .B(n1103), .ZN(G6) );
NOR2_X1 U805 ( .A1(n1109), .A2(n1118), .ZN(G57) );
XOR2_X1 U806 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U807 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U808 ( .A1(KEYINPUT49), .A2(n1123), .ZN(n1121) );
XOR2_X1 U809 ( .A(KEYINPUT46), .B(n1124), .Z(n1119) );
NOR2_X1 U810 ( .A1(n1125), .A2(n1108), .ZN(n1124) );
XNOR2_X1 U811 ( .A(G472), .B(KEYINPUT25), .ZN(n1125) );
NOR2_X1 U812 ( .A1(n1126), .A2(n1127), .ZN(G54) );
XOR2_X1 U813 ( .A(KEYINPUT51), .B(n1109), .Z(n1127) );
XOR2_X1 U814 ( .A(n1128), .B(n1129), .Z(n1126) );
XOR2_X1 U815 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U816 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U817 ( .A1(KEYINPUT9), .A2(n1134), .ZN(n1133) );
NOR2_X1 U818 ( .A1(n1036), .A2(n1108), .ZN(n1132) );
INV_X1 U819 ( .A(G469), .ZN(n1036) );
XNOR2_X1 U820 ( .A(G140), .B(n1135), .ZN(n1130) );
XNOR2_X1 U821 ( .A(n1136), .B(n1137), .ZN(n1128) );
XNOR2_X1 U822 ( .A(n1138), .B(n1139), .ZN(n1136) );
NOR2_X1 U823 ( .A1(n1109), .A2(n1140), .ZN(G51) );
XOR2_X1 U824 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U825 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U826 ( .A1(n1038), .A2(n1108), .ZN(n1144) );
NAND2_X1 U827 ( .A1(G902), .A2(n1067), .ZN(n1108) );
NAND3_X1 U828 ( .A1(n1101), .A2(n1103), .A3(n1083), .ZN(n1067) );
AND4_X1 U829 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1083) );
NOR4_X1 U830 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1148) );
NOR2_X1 U831 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
XNOR2_X1 U832 ( .A(KEYINPUT40), .B(n1051), .ZN(n1154) );
AND2_X1 U833 ( .A1(n1155), .A2(n1156), .ZN(n1147) );
NAND3_X1 U834 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1145) );
XOR2_X1 U835 ( .A(KEYINPUT56), .B(n1049), .Z(n1158) );
NAND3_X1 U836 ( .A1(n1160), .A2(n1053), .A3(n1064), .ZN(n1103) );
AND4_X1 U837 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1101) );
NOR4_X1 U838 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
INV_X1 U839 ( .A(n1012), .ZN(n1168) );
NAND3_X1 U840 ( .A1(n1063), .A2(n1053), .A3(n1160), .ZN(n1012) );
NAND3_X1 U841 ( .A1(n1160), .A2(n1169), .A3(n1043), .ZN(n1163) );
NOR2_X1 U842 ( .A1(KEYINPUT43), .A2(n1170), .ZN(n1143) );
XOR2_X1 U843 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U844 ( .A(G125), .B(n1173), .Z(n1172) );
NOR2_X1 U845 ( .A1(KEYINPUT0), .A2(n1174), .ZN(n1171) );
INV_X1 U846 ( .A(n1175), .ZN(n1174) );
NOR2_X1 U847 ( .A1(n1016), .A2(G952), .ZN(n1109) );
XNOR2_X1 U848 ( .A(G146), .B(n1146), .ZN(G48) );
NAND3_X1 U849 ( .A1(n1176), .A2(n1177), .A3(n1159), .ZN(n1146) );
XNOR2_X1 U850 ( .A(G143), .B(n1156), .ZN(G45) );
NAND3_X1 U851 ( .A1(n1157), .A2(n1178), .A3(n1179), .ZN(n1156) );
NOR3_X1 U852 ( .A1(n1055), .A2(n1180), .A3(n1026), .ZN(n1179) );
XNOR2_X1 U853 ( .A(G140), .B(n1181), .ZN(G42) );
OR2_X1 U854 ( .A1(n1153), .A2(n1051), .ZN(n1181) );
NAND2_X1 U855 ( .A1(n1182), .A2(n1183), .ZN(G39) );
OR2_X1 U856 ( .A1(n1155), .A2(G137), .ZN(n1183) );
XOR2_X1 U857 ( .A(n1184), .B(KEYINPUT10), .Z(n1182) );
NAND2_X1 U858 ( .A1(G137), .A2(n1155), .ZN(n1184) );
NAND4_X1 U859 ( .A1(n1043), .A2(n1049), .A3(n1178), .A4(n1176), .ZN(n1155) );
XOR2_X1 U860 ( .A(G134), .B(n1150), .Z(G36) );
AND4_X1 U861 ( .A1(n1157), .A2(n1049), .A3(n1178), .A4(n1063), .ZN(n1150) );
XOR2_X1 U862 ( .A(n1185), .B(n1186), .Z(G33) );
NOR2_X1 U863 ( .A1(KEYINPUT39), .A2(n1187), .ZN(n1186) );
NOR2_X1 U864 ( .A1(n1052), .A2(n1153), .ZN(n1185) );
NAND2_X1 U865 ( .A1(n1159), .A2(n1049), .ZN(n1153) );
AND2_X1 U866 ( .A1(n1057), .A2(n1188), .ZN(n1049) );
XNOR2_X1 U867 ( .A(n1189), .B(KEYINPUT42), .ZN(n1057) );
AND2_X1 U868 ( .A1(n1064), .A2(n1178), .ZN(n1159) );
AND2_X1 U869 ( .A1(n1065), .A2(n1190), .ZN(n1178) );
XNOR2_X1 U870 ( .A(n1191), .B(KEYINPUT26), .ZN(n1065) );
XNOR2_X1 U871 ( .A(G128), .B(n1192), .ZN(G30) );
NAND2_X1 U872 ( .A1(KEYINPUT41), .A2(n1149), .ZN(n1192) );
AND4_X1 U873 ( .A1(n1176), .A2(n1063), .A3(n1193), .A4(n1191), .ZN(n1149) );
NOR2_X1 U874 ( .A1(n1194), .A2(n1055), .ZN(n1193) );
XNOR2_X1 U875 ( .A(G101), .B(n1161), .ZN(G3) );
NAND3_X1 U876 ( .A1(n1157), .A2(n1160), .A3(n1043), .ZN(n1161) );
NOR3_X1 U877 ( .A1(n1055), .A2(n1195), .A3(n1196), .ZN(n1160) );
INV_X1 U878 ( .A(n1191), .ZN(n1196) );
XOR2_X1 U879 ( .A(G125), .B(n1152), .Z(G27) );
AND4_X1 U880 ( .A1(n1169), .A2(n1177), .A3(n1064), .A4(n1197), .ZN(n1152) );
NOR3_X1 U881 ( .A1(n1198), .A2(n1022), .A3(n1194), .ZN(n1197) );
INV_X1 U882 ( .A(n1190), .ZN(n1194) );
NAND2_X1 U883 ( .A1(n1066), .A2(n1199), .ZN(n1190) );
NAND4_X1 U884 ( .A1(G953), .A2(G902), .A3(n1200), .A4(n1074), .ZN(n1199) );
INV_X1 U885 ( .A(G900), .ZN(n1074) );
XOR2_X1 U886 ( .A(n1162), .B(n1201), .Z(G24) );
NAND2_X1 U887 ( .A1(KEYINPUT32), .A2(G122), .ZN(n1201) );
NAND4_X1 U888 ( .A1(n1202), .A2(n1053), .A3(n1203), .A4(n1204), .ZN(n1162) );
NAND2_X1 U889 ( .A1(n1205), .A2(n1206), .ZN(n1053) );
OR2_X1 U890 ( .A1(n1051), .A2(KEYINPUT35), .ZN(n1206) );
INV_X1 U891 ( .A(n1169), .ZN(n1051) );
NAND3_X1 U892 ( .A1(n1207), .A2(n1027), .A3(KEYINPUT35), .ZN(n1205) );
XOR2_X1 U893 ( .A(G119), .B(n1167), .Z(G21) );
AND3_X1 U894 ( .A1(n1043), .A2(n1176), .A3(n1202), .ZN(n1167) );
NOR2_X1 U895 ( .A1(n1207), .A2(n1027), .ZN(n1176) );
INV_X1 U896 ( .A(n1208), .ZN(n1027) );
XOR2_X1 U897 ( .A(G116), .B(n1166), .Z(G18) );
AND3_X1 U898 ( .A1(n1157), .A2(n1063), .A3(n1202), .ZN(n1166) );
NOR2_X1 U899 ( .A1(n1203), .A2(n1180), .ZN(n1063) );
INV_X1 U900 ( .A(n1204), .ZN(n1180) );
XOR2_X1 U901 ( .A(n1209), .B(n1165), .Z(G15) );
AND3_X1 U902 ( .A1(n1064), .A2(n1157), .A3(n1202), .ZN(n1165) );
NOR4_X1 U903 ( .A1(n1055), .A2(n1198), .A3(n1022), .A4(n1195), .ZN(n1202) );
INV_X1 U904 ( .A(n1044), .ZN(n1198) );
INV_X1 U905 ( .A(n1052), .ZN(n1157) );
NAND2_X1 U906 ( .A1(n1210), .A2(n1208), .ZN(n1052) );
XNOR2_X1 U907 ( .A(KEYINPUT35), .B(n1207), .ZN(n1210) );
NOR2_X1 U908 ( .A1(n1204), .A2(n1026), .ZN(n1064) );
INV_X1 U909 ( .A(n1203), .ZN(n1026) );
NAND2_X1 U910 ( .A1(KEYINPUT21), .A2(n1098), .ZN(n1209) );
XNOR2_X1 U911 ( .A(G110), .B(n1211), .ZN(G12) );
NAND4_X1 U912 ( .A1(n1043), .A2(n1169), .A3(n1212), .A4(n1191), .ZN(n1211) );
NOR2_X1 U913 ( .A1(n1044), .A2(n1022), .ZN(n1191) );
INV_X1 U914 ( .A(n1046), .ZN(n1022) );
NAND2_X1 U915 ( .A1(G221), .A2(n1213), .ZN(n1046) );
XNOR2_X1 U916 ( .A(n1035), .B(n1214), .ZN(n1044) );
NOR2_X1 U917 ( .A1(G469), .A2(KEYINPUT5), .ZN(n1214) );
NAND2_X1 U918 ( .A1(n1215), .A2(n1216), .ZN(n1035) );
XOR2_X1 U919 ( .A(n1217), .B(n1218), .Z(n1215) );
XNOR2_X1 U920 ( .A(n1219), .B(n1077), .ZN(n1218) );
INV_X1 U921 ( .A(n1138), .ZN(n1077) );
NOR2_X1 U922 ( .A1(KEYINPUT1), .A2(n1220), .ZN(n1219) );
XNOR2_X1 U923 ( .A(n1137), .B(n1078), .ZN(n1220) );
XOR2_X1 U924 ( .A(n1135), .B(n1221), .Z(n1078) );
NAND2_X1 U925 ( .A1(KEYINPUT44), .A2(n1222), .ZN(n1135) );
XNOR2_X1 U926 ( .A(n1223), .B(G143), .ZN(n1222) );
INV_X1 U927 ( .A(G146), .ZN(n1223) );
NAND2_X1 U928 ( .A1(n1224), .A2(n1225), .ZN(n1137) );
NAND2_X1 U929 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
INV_X1 U930 ( .A(G107), .ZN(n1227) );
XOR2_X1 U931 ( .A(KEYINPUT50), .B(n1228), .Z(n1226) );
NAND2_X1 U932 ( .A1(n1228), .A2(G107), .ZN(n1224) );
NAND2_X1 U933 ( .A1(n1229), .A2(n1230), .ZN(n1217) );
NAND2_X1 U934 ( .A1(KEYINPUT13), .A2(n1231), .ZN(n1230) );
INV_X1 U935 ( .A(n1232), .ZN(n1231) );
NAND2_X1 U936 ( .A1(KEYINPUT28), .A2(n1232), .ZN(n1229) );
XNOR2_X1 U937 ( .A(n1134), .B(n1233), .ZN(n1232) );
NOR2_X1 U938 ( .A1(KEYINPUT16), .A2(n1234), .ZN(n1233) );
XNOR2_X1 U939 ( .A(G140), .B(n1235), .ZN(n1234) );
NOR2_X1 U940 ( .A1(KEYINPUT24), .A2(n1236), .ZN(n1235) );
NAND2_X1 U941 ( .A1(G227), .A2(n1016), .ZN(n1134) );
NOR2_X1 U942 ( .A1(n1195), .A2(n1237), .ZN(n1212) );
XNOR2_X1 U943 ( .A(n1177), .B(KEYINPUT37), .ZN(n1237) );
INV_X1 U944 ( .A(n1055), .ZN(n1177) );
NAND2_X1 U945 ( .A1(n1238), .A2(n1189), .ZN(n1055) );
XOR2_X1 U946 ( .A(n1239), .B(n1240), .Z(n1189) );
NOR2_X1 U947 ( .A1(n1241), .A2(KEYINPUT18), .ZN(n1240) );
INV_X1 U948 ( .A(n1038), .ZN(n1241) );
NAND2_X1 U949 ( .A1(G210), .A2(n1242), .ZN(n1038) );
XOR2_X1 U950 ( .A(n1037), .B(KEYINPUT33), .Z(n1239) );
NAND2_X1 U951 ( .A1(n1243), .A2(n1216), .ZN(n1037) );
XOR2_X1 U952 ( .A(n1244), .B(n1245), .Z(n1243) );
NOR2_X1 U953 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XOR2_X1 U954 ( .A(n1248), .B(KEYINPUT48), .Z(n1247) );
NAND2_X1 U955 ( .A1(G125), .A2(n1175), .ZN(n1248) );
NOR2_X1 U956 ( .A1(G125), .A2(n1175), .ZN(n1246) );
XNOR2_X1 U957 ( .A(n1249), .B(n1250), .ZN(n1244) );
NOR2_X1 U958 ( .A1(KEYINPUT11), .A2(n1141), .ZN(n1250) );
XNOR2_X1 U959 ( .A(n1093), .B(n1251), .ZN(n1141) );
XOR2_X1 U960 ( .A(n1099), .B(n1252), .Z(n1251) );
XNOR2_X1 U961 ( .A(n1253), .B(n1228), .ZN(n1093) );
XNOR2_X1 U962 ( .A(G104), .B(n1254), .ZN(n1228) );
XNOR2_X1 U963 ( .A(G107), .B(G110), .ZN(n1253) );
NOR2_X1 U964 ( .A1(KEYINPUT4), .A2(n1255), .ZN(n1249) );
XNOR2_X1 U965 ( .A(n1173), .B(KEYINPUT23), .ZN(n1255) );
NOR2_X1 U966 ( .A1(n1089), .A2(G953), .ZN(n1173) );
INV_X1 U967 ( .A(G224), .ZN(n1089) );
XNOR2_X1 U968 ( .A(n1021), .B(KEYINPUT22), .ZN(n1238) );
INV_X1 U969 ( .A(n1188), .ZN(n1021) );
NAND2_X1 U970 ( .A1(G214), .A2(n1242), .ZN(n1188) );
NAND2_X1 U971 ( .A1(n1256), .A2(n1216), .ZN(n1242) );
INV_X1 U972 ( .A(G237), .ZN(n1256) );
AND2_X1 U973 ( .A1(n1257), .A2(n1066), .ZN(n1195) );
NAND3_X1 U974 ( .A1(n1200), .A2(n1016), .A3(G952), .ZN(n1066) );
NAND4_X1 U975 ( .A1(G953), .A2(G902), .A3(n1200), .A4(n1090), .ZN(n1257) );
INV_X1 U976 ( .A(G898), .ZN(n1090) );
NAND2_X1 U977 ( .A1(G237), .A2(G234), .ZN(n1200) );
NOR2_X1 U978 ( .A1(n1207), .A2(n1208), .ZN(n1169) );
XNOR2_X1 U979 ( .A(n1258), .B(G472), .ZN(n1208) );
NAND2_X1 U980 ( .A1(n1259), .A2(n1216), .ZN(n1258) );
XOR2_X1 U981 ( .A(n1123), .B(n1122), .Z(n1259) );
XNOR2_X1 U982 ( .A(n1260), .B(n1261), .ZN(n1122) );
XNOR2_X1 U983 ( .A(n1138), .B(n1175), .ZN(n1261) );
NAND2_X1 U984 ( .A1(n1262), .A2(n1263), .ZN(n1175) );
NAND2_X1 U985 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
XOR2_X1 U986 ( .A(KEYINPUT6), .B(n1266), .Z(n1264) );
NAND2_X1 U987 ( .A1(n1267), .A2(G143), .ZN(n1262) );
XOR2_X1 U988 ( .A(KEYINPUT36), .B(n1266), .Z(n1267) );
XNOR2_X1 U989 ( .A(n1268), .B(G146), .ZN(n1266) );
NAND2_X1 U990 ( .A1(KEYINPUT29), .A2(n1221), .ZN(n1268) );
INV_X1 U991 ( .A(G128), .ZN(n1221) );
XOR2_X1 U992 ( .A(G131), .B(n1269), .Z(n1138) );
XOR2_X1 U993 ( .A(G137), .B(G134), .Z(n1269) );
XOR2_X1 U994 ( .A(n1270), .B(KEYINPUT15), .Z(n1260) );
NAND3_X1 U995 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1270) );
NAND2_X1 U996 ( .A1(G113), .A2(n1274), .ZN(n1273) );
OR3_X1 U997 ( .A1(n1274), .A2(G113), .A3(KEYINPUT20), .ZN(n1272) );
NAND2_X1 U998 ( .A1(KEYINPUT47), .A2(n1099), .ZN(n1274) );
INV_X1 U999 ( .A(n1275), .ZN(n1099) );
NAND2_X1 U1000 ( .A1(KEYINPUT20), .A2(n1275), .ZN(n1271) );
XNOR2_X1 U1001 ( .A(G116), .B(n1276), .ZN(n1275) );
AND2_X1 U1002 ( .A1(n1277), .A2(n1278), .ZN(n1123) );
NAND2_X1 U1003 ( .A1(n1279), .A2(n1254), .ZN(n1278) );
INV_X1 U1004 ( .A(G101), .ZN(n1254) );
NAND2_X1 U1005 ( .A1(n1280), .A2(G210), .ZN(n1279) );
NAND3_X1 U1006 ( .A1(n1280), .A2(G210), .A3(G101), .ZN(n1277) );
XOR2_X1 U1007 ( .A(n1281), .B(n1029), .Z(n1207) );
NAND2_X1 U1008 ( .A1(G217), .A2(n1213), .ZN(n1029) );
NAND2_X1 U1009 ( .A1(G234), .A2(n1216), .ZN(n1213) );
INV_X1 U1010 ( .A(G902), .ZN(n1216) );
NAND2_X1 U1011 ( .A1(KEYINPUT8), .A2(n1028), .ZN(n1281) );
OR2_X1 U1012 ( .A1(n1107), .A2(G902), .ZN(n1028) );
XNOR2_X1 U1013 ( .A(n1282), .B(n1283), .ZN(n1107) );
XOR2_X1 U1014 ( .A(G137), .B(n1284), .Z(n1283) );
NOR2_X1 U1015 ( .A1(KEYINPUT52), .A2(n1285), .ZN(n1284) );
XOR2_X1 U1016 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U1017 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U1018 ( .A(KEYINPUT61), .B(KEYINPUT38), .Z(n1289) );
NOR2_X1 U1019 ( .A1(KEYINPUT31), .A2(n1290), .ZN(n1288) );
XNOR2_X1 U1020 ( .A(n1291), .B(n1292), .ZN(n1290) );
NOR2_X1 U1021 ( .A1(KEYINPUT54), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U1022 ( .A(n1276), .B(n1139), .ZN(n1286) );
XNOR2_X1 U1023 ( .A(n1236), .B(G128), .ZN(n1139) );
INV_X1 U1024 ( .A(G110), .ZN(n1236) );
XOR2_X1 U1025 ( .A(G119), .B(KEYINPUT34), .Z(n1276) );
NAND2_X1 U1026 ( .A1(n1294), .A2(G221), .ZN(n1282) );
NOR2_X1 U1027 ( .A1(n1204), .A2(n1203), .ZN(n1043) );
XOR2_X1 U1028 ( .A(n1295), .B(n1117), .Z(n1203) );
INV_X1 U1029 ( .A(G475), .ZN(n1117) );
OR2_X1 U1030 ( .A1(n1116), .A2(G902), .ZN(n1295) );
XNOR2_X1 U1031 ( .A(n1296), .B(n1297), .ZN(n1116) );
XOR2_X1 U1032 ( .A(G104), .B(n1298), .Z(n1297) );
NOR2_X1 U1033 ( .A1(KEYINPUT59), .A2(n1299), .ZN(n1298) );
XOR2_X1 U1034 ( .A(n1300), .B(n1301), .Z(n1299) );
XNOR2_X1 U1035 ( .A(n1302), .B(n1265), .ZN(n1301) );
NAND2_X1 U1036 ( .A1(n1280), .A2(G214), .ZN(n1302) );
NOR2_X1 U1037 ( .A1(G953), .A2(G237), .ZN(n1280) );
NAND2_X1 U1038 ( .A1(KEYINPUT63), .A2(n1187), .ZN(n1300) );
INV_X1 U1039 ( .A(G131), .ZN(n1187) );
XOR2_X1 U1040 ( .A(n1303), .B(n1252), .Z(n1296) );
XNOR2_X1 U1041 ( .A(n1098), .B(G122), .ZN(n1252) );
INV_X1 U1042 ( .A(G113), .ZN(n1098) );
NAND3_X1 U1043 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n1303) );
NAND2_X1 U1044 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
INV_X1 U1045 ( .A(n1291), .ZN(n1307) );
NAND3_X1 U1046 ( .A1(n1309), .A2(n1291), .A3(KEYINPUT57), .ZN(n1305) );
XOR2_X1 U1047 ( .A(G146), .B(KEYINPUT62), .Z(n1291) );
INV_X1 U1048 ( .A(n1308), .ZN(n1309) );
NAND2_X1 U1049 ( .A1(KEYINPUT12), .A2(n1293), .ZN(n1308) );
OR2_X1 U1050 ( .A1(n1293), .A2(KEYINPUT57), .ZN(n1304) );
XOR2_X1 U1051 ( .A(G140), .B(G125), .Z(n1293) );
NAND2_X1 U1052 ( .A1(n1033), .A2(n1310), .ZN(n1204) );
NAND2_X1 U1053 ( .A1(G478), .A2(n1034), .ZN(n1310) );
INV_X1 U1054 ( .A(n1311), .ZN(n1034) );
NAND2_X1 U1055 ( .A1(n1311), .A2(n1113), .ZN(n1033) );
INV_X1 U1056 ( .A(G478), .ZN(n1113) );
NOR2_X1 U1057 ( .A1(n1112), .A2(G902), .ZN(n1311) );
XNOR2_X1 U1058 ( .A(n1312), .B(n1313), .ZN(n1112) );
XNOR2_X1 U1059 ( .A(n1314), .B(n1315), .ZN(n1313) );
NOR2_X1 U1060 ( .A1(G107), .A2(KEYINPUT53), .ZN(n1315) );
NAND2_X1 U1061 ( .A1(KEYINPUT3), .A2(n1095), .ZN(n1314) );
INV_X1 U1062 ( .A(G122), .ZN(n1095) );
XOR2_X1 U1063 ( .A(n1316), .B(n1317), .Z(n1312) );
XNOR2_X1 U1064 ( .A(G116), .B(n1318), .ZN(n1317) );
NAND2_X1 U1065 ( .A1(n1319), .A2(KEYINPUT19), .ZN(n1318) );
XNOR2_X1 U1066 ( .A(G128), .B(n1320), .ZN(n1319) );
XNOR2_X1 U1067 ( .A(n1265), .B(G134), .ZN(n1320) );
INV_X1 U1068 ( .A(G143), .ZN(n1265) );
NAND3_X1 U1069 ( .A1(G217), .A2(n1294), .A3(KEYINPUT27), .ZN(n1316) );
AND2_X1 U1070 ( .A1(G234), .A2(n1016), .ZN(n1294) );
INV_X1 U1071 ( .A(G953), .ZN(n1016) );
endmodule


