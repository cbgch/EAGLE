//Key = 1100011000010111100000111001111111101101000101000000010100110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381;

XOR2_X1 U738 ( .A(G107), .B(n1040), .Z(G9) );
NOR2_X1 U739 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR2_X1 U740 ( .A1(n1043), .A2(n1044), .ZN(G75) );
NOR3_X1 U741 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NOR2_X1 U742 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR3_X1 U743 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1048) );
NOR2_X1 U744 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
INV_X1 U745 ( .A(n1055), .ZN(n1054) );
NOR2_X1 U746 ( .A1(n1056), .A2(n1057), .ZN(n1053) );
NOR2_X1 U747 ( .A1(KEYINPUT51), .A2(n1058), .ZN(n1056) );
NOR3_X1 U748 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1051) );
NOR2_X1 U749 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U750 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U751 ( .A1(n1066), .A2(n1067), .ZN(n1062) );
NOR2_X1 U752 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
XOR2_X1 U753 ( .A(n1070), .B(KEYINPUT36), .Z(n1050) );
NAND4_X1 U754 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1070) );
NOR2_X1 U755 ( .A1(n1059), .A2(n1075), .ZN(n1074) );
INV_X1 U756 ( .A(n1076), .ZN(n1071) );
NAND3_X1 U757 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1045) );
NAND2_X1 U758 ( .A1(n1055), .A2(n1080), .ZN(n1079) );
NAND2_X1 U759 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND3_X1 U760 ( .A1(n1083), .A2(n1049), .A3(KEYINPUT51), .ZN(n1082) );
NAND2_X1 U761 ( .A1(n1072), .A2(n1084), .ZN(n1081) );
NAND2_X1 U762 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U763 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR3_X1 U764 ( .A1(n1065), .A2(n1067), .A3(n1059), .ZN(n1055) );
NOR3_X1 U765 ( .A1(n1089), .A2(G953), .A3(G952), .ZN(n1043) );
INV_X1 U766 ( .A(n1077), .ZN(n1089) );
NAND4_X1 U767 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1077) );
NOR4_X1 U768 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1093) );
XNOR2_X1 U769 ( .A(G472), .B(n1098), .ZN(n1097) );
XOR2_X1 U770 ( .A(n1099), .B(n1100), .Z(n1095) );
XOR2_X1 U771 ( .A(KEYINPUT38), .B(n1101), .Z(n1100) );
NOR2_X1 U772 ( .A1(KEYINPUT21), .A2(G469), .ZN(n1101) );
XOR2_X1 U773 ( .A(n1102), .B(n1103), .Z(n1094) );
NOR2_X1 U774 ( .A1(KEYINPUT49), .A2(n1104), .ZN(n1103) );
XNOR2_X1 U775 ( .A(G478), .B(KEYINPUT2), .ZN(n1102) );
NOR3_X1 U776 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1092) );
XOR2_X1 U777 ( .A(n1108), .B(n1109), .Z(n1090) );
NOR2_X1 U778 ( .A1(n1110), .A2(KEYINPUT9), .ZN(n1109) );
INV_X1 U779 ( .A(n1111), .ZN(n1110) );
XOR2_X1 U780 ( .A(n1112), .B(n1113), .Z(G72) );
XOR2_X1 U781 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U782 ( .A1(G953), .A2(n1116), .ZN(n1115) );
NAND2_X1 U783 ( .A1(G900), .A2(G227), .ZN(n1116) );
NAND2_X1 U784 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
NAND2_X1 U785 ( .A1(G953), .A2(n1119), .ZN(n1118) );
XOR2_X1 U786 ( .A(n1120), .B(n1121), .Z(n1117) );
XOR2_X1 U787 ( .A(n1122), .B(n1123), .Z(n1121) );
XNOR2_X1 U788 ( .A(KEYINPUT17), .B(n1124), .ZN(n1123) );
XOR2_X1 U789 ( .A(KEYINPUT44), .B(KEYINPUT37), .Z(n1122) );
XOR2_X1 U790 ( .A(n1125), .B(n1126), .Z(n1120) );
XOR2_X1 U791 ( .A(n1127), .B(n1128), .Z(n1125) );
NOR2_X1 U792 ( .A1(G137), .A2(KEYINPUT56), .ZN(n1128) );
NOR2_X1 U793 ( .A1(n1129), .A2(G953), .ZN(n1112) );
NOR2_X1 U794 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U795 ( .A(KEYINPUT54), .B(n1132), .Z(n1131) );
NAND2_X1 U796 ( .A1(n1133), .A2(n1134), .ZN(G69) );
NAND2_X1 U797 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U798 ( .A1(G953), .A2(n1137), .ZN(n1135) );
NAND2_X1 U799 ( .A1(G898), .A2(G224), .ZN(n1137) );
NAND2_X1 U800 ( .A1(n1138), .A2(n1139), .ZN(n1133) );
NAND2_X1 U801 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U802 ( .A1(G953), .A2(n1142), .ZN(n1141) );
INV_X1 U803 ( .A(n1136), .ZN(n1138) );
NAND2_X1 U804 ( .A1(n1143), .A2(n1144), .ZN(n1136) );
NAND2_X1 U805 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U806 ( .A(KEYINPUT22), .B(n1147), .Z(n1143) );
NOR2_X1 U807 ( .A1(n1145), .A2(n1146), .ZN(n1147) );
NAND2_X1 U808 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
XNOR2_X1 U809 ( .A(G953), .B(KEYINPUT7), .ZN(n1148) );
AND3_X1 U810 ( .A1(n1150), .A2(n1151), .A3(n1140), .ZN(n1145) );
INV_X1 U811 ( .A(n1152), .ZN(n1140) );
OR2_X1 U812 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
NAND2_X1 U813 ( .A1(n1155), .A2(n1154), .ZN(n1150) );
XOR2_X1 U814 ( .A(KEYINPUT61), .B(n1153), .Z(n1155) );
NOR2_X1 U815 ( .A1(n1156), .A2(n1157), .ZN(G66) );
NOR3_X1 U816 ( .A1(n1108), .A2(n1158), .A3(n1159), .ZN(n1157) );
NOR3_X1 U817 ( .A1(n1160), .A2(n1111), .A3(n1161), .ZN(n1159) );
INV_X1 U818 ( .A(n1162), .ZN(n1160) );
NOR2_X1 U819 ( .A1(n1163), .A2(n1162), .ZN(n1158) );
NOR2_X1 U820 ( .A1(n1164), .A2(n1111), .ZN(n1163) );
NOR2_X1 U821 ( .A1(n1156), .A2(n1165), .ZN(G63) );
XOR2_X1 U822 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U823 ( .A(n1168), .B(KEYINPUT42), .Z(n1167) );
NAND3_X1 U824 ( .A1(n1169), .A2(n1170), .A3(G478), .ZN(n1168) );
NAND2_X1 U825 ( .A1(KEYINPUT43), .A2(n1161), .ZN(n1170) );
NAND2_X1 U826 ( .A1(n1171), .A2(n1172), .ZN(n1169) );
INV_X1 U827 ( .A(KEYINPUT43), .ZN(n1172) );
NAND2_X1 U828 ( .A1(n1164), .A2(G902), .ZN(n1171) );
NOR2_X1 U829 ( .A1(n1156), .A2(n1173), .ZN(G60) );
XNOR2_X1 U830 ( .A(n1174), .B(n1175), .ZN(n1173) );
NOR2_X1 U831 ( .A1(n1176), .A2(n1161), .ZN(n1175) );
XNOR2_X1 U832 ( .A(G104), .B(n1177), .ZN(G6) );
NOR2_X1 U833 ( .A1(n1178), .A2(KEYINPUT26), .ZN(n1177) );
NOR3_X1 U834 ( .A1(n1156), .A2(n1179), .A3(n1180), .ZN(G57) );
NOR2_X1 U835 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U836 ( .A(n1183), .B(n1184), .Z(n1182) );
OR2_X1 U837 ( .A1(n1185), .A2(KEYINPUT3), .ZN(n1183) );
INV_X1 U838 ( .A(n1186), .ZN(n1181) );
NOR2_X1 U839 ( .A1(n1186), .A2(n1187), .ZN(n1179) );
XOR2_X1 U840 ( .A(n1188), .B(n1184), .Z(n1187) );
XOR2_X1 U841 ( .A(n1189), .B(n1190), .Z(n1184) );
NOR2_X1 U842 ( .A1(n1191), .A2(n1161), .ZN(n1190) );
INV_X1 U843 ( .A(G472), .ZN(n1191) );
NAND2_X1 U844 ( .A1(n1185), .A2(n1192), .ZN(n1188) );
INV_X1 U845 ( .A(KEYINPUT3), .ZN(n1192) );
NOR2_X1 U846 ( .A1(n1156), .A2(n1193), .ZN(G54) );
XOR2_X1 U847 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U848 ( .A(n1196), .B(n1197), .Z(n1195) );
XNOR2_X1 U849 ( .A(G110), .B(n1198), .ZN(n1197) );
NOR2_X1 U850 ( .A1(n1199), .A2(n1161), .ZN(n1196) );
XOR2_X1 U851 ( .A(n1200), .B(n1201), .Z(n1194) );
XNOR2_X1 U852 ( .A(n1202), .B(n1203), .ZN(n1200) );
NOR2_X1 U853 ( .A1(KEYINPUT60), .A2(n1204), .ZN(n1203) );
NOR2_X1 U854 ( .A1(n1156), .A2(n1205), .ZN(G51) );
XOR2_X1 U855 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U856 ( .A(n1208), .B(n1209), .Z(n1207) );
NOR2_X1 U857 ( .A1(G125), .A2(KEYINPUT47), .ZN(n1209) );
NOR2_X1 U858 ( .A1(n1210), .A2(n1161), .ZN(n1208) );
NAND2_X1 U859 ( .A1(G902), .A2(n1047), .ZN(n1161) );
INV_X1 U860 ( .A(n1164), .ZN(n1047) );
NOR3_X1 U861 ( .A1(n1130), .A2(n1132), .A3(n1149), .ZN(n1164) );
NAND4_X1 U862 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1149) );
NOR3_X1 U863 ( .A1(n1215), .A2(n1216), .A3(n1178), .ZN(n1214) );
NOR2_X1 U864 ( .A1(n1217), .A2(n1041), .ZN(n1178) );
NAND2_X1 U865 ( .A1(n1072), .A2(n1218), .ZN(n1041) );
NOR2_X1 U866 ( .A1(n1219), .A2(n1220), .ZN(n1215) );
NOR3_X1 U867 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1219) );
NOR3_X1 U868 ( .A1(n1065), .A2(n1064), .A3(n1224), .ZN(n1223) );
NOR3_X1 U869 ( .A1(n1225), .A2(n1061), .A3(n1042), .ZN(n1222) );
INV_X1 U870 ( .A(n1072), .ZN(n1061) );
XNOR2_X1 U871 ( .A(KEYINPUT13), .B(n1064), .ZN(n1225) );
NOR2_X1 U872 ( .A1(n1067), .A2(n1226), .ZN(n1221) );
AND2_X1 U873 ( .A1(n1227), .A2(n1228), .ZN(n1132) );
XNOR2_X1 U874 ( .A(n1229), .B(KEYINPUT6), .ZN(n1227) );
NAND4_X1 U875 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1130) );
NOR4_X1 U876 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1233) );
NAND3_X1 U877 ( .A1(n1073), .A2(n1238), .A3(n1239), .ZN(n1232) );
AND2_X1 U878 ( .A1(n1240), .A2(G953), .ZN(n1156) );
XNOR2_X1 U879 ( .A(G952), .B(KEYINPUT20), .ZN(n1240) );
XNOR2_X1 U880 ( .A(G146), .B(n1241), .ZN(G48) );
NAND2_X1 U881 ( .A1(KEYINPUT29), .A2(n1242), .ZN(n1241) );
INV_X1 U882 ( .A(n1230), .ZN(n1242) );
NAND3_X1 U883 ( .A1(n1069), .A2(n1238), .A3(n1243), .ZN(n1230) );
XNOR2_X1 U884 ( .A(G143), .B(n1231), .ZN(G45) );
NAND4_X1 U885 ( .A1(n1243), .A2(n1083), .A3(n1096), .A4(n1244), .ZN(n1231) );
XNOR2_X1 U886 ( .A(n1245), .B(n1237), .ZN(G42) );
NOR3_X1 U887 ( .A1(n1217), .A2(n1224), .A3(n1246), .ZN(n1237) );
XOR2_X1 U888 ( .A(G137), .B(n1247), .Z(G39) );
NOR3_X1 U889 ( .A1(n1246), .A2(n1065), .A3(n1248), .ZN(n1247) );
XNOR2_X1 U890 ( .A(KEYINPUT40), .B(n1238), .ZN(n1248) );
INV_X1 U891 ( .A(n1073), .ZN(n1065) );
XOR2_X1 U892 ( .A(n1249), .B(n1236), .Z(G36) );
NOR3_X1 U893 ( .A1(n1042), .A2(n1058), .A3(n1246), .ZN(n1236) );
INV_X1 U894 ( .A(n1083), .ZN(n1058) );
INV_X1 U895 ( .A(n1068), .ZN(n1042) );
NAND2_X1 U896 ( .A1(KEYINPUT45), .A2(n1124), .ZN(n1249) );
XNOR2_X1 U897 ( .A(n1250), .B(n1235), .ZN(G33) );
NOR2_X1 U898 ( .A1(n1246), .A2(n1226), .ZN(n1235) );
INV_X1 U899 ( .A(n1239), .ZN(n1246) );
NOR3_X1 U900 ( .A1(n1064), .A2(n1251), .A3(n1049), .ZN(n1239) );
NAND2_X1 U901 ( .A1(n1088), .A2(n1091), .ZN(n1049) );
XOR2_X1 U902 ( .A(G128), .B(n1234), .Z(G30) );
AND3_X1 U903 ( .A1(n1068), .A2(n1238), .A3(n1243), .ZN(n1234) );
NOR3_X1 U904 ( .A1(n1085), .A2(n1251), .A3(n1064), .ZN(n1243) );
XOR2_X1 U905 ( .A(G101), .B(n1216), .Z(G3) );
AND3_X1 U906 ( .A1(n1218), .A2(n1083), .A3(n1073), .ZN(n1216) );
XNOR2_X1 U907 ( .A(G125), .B(n1252), .ZN(G27) );
NAND3_X1 U908 ( .A1(n1228), .A2(n1229), .A3(KEYINPUT5), .ZN(n1252) );
NOR4_X1 U909 ( .A1(n1217), .A2(n1224), .A3(n1085), .A4(n1251), .ZN(n1228) );
AND2_X1 U910 ( .A1(n1059), .A2(n1253), .ZN(n1251) );
NAND4_X1 U911 ( .A1(n1254), .A2(G902), .A3(G953), .A4(n1119), .ZN(n1253) );
INV_X1 U912 ( .A(G900), .ZN(n1119) );
XOR2_X1 U913 ( .A(n1255), .B(KEYINPUT35), .Z(n1254) );
INV_X1 U914 ( .A(n1256), .ZN(n1085) );
INV_X1 U915 ( .A(n1057), .ZN(n1224) );
XNOR2_X1 U916 ( .A(G122), .B(n1213), .ZN(G24) );
NAND4_X1 U917 ( .A1(n1257), .A2(n1072), .A3(n1096), .A4(n1244), .ZN(n1213) );
XOR2_X1 U918 ( .A(n1211), .B(n1258), .Z(G21) );
NAND2_X1 U919 ( .A1(KEYINPUT28), .A2(G119), .ZN(n1258) );
NAND3_X1 U920 ( .A1(n1257), .A2(n1238), .A3(n1073), .ZN(n1211) );
NAND2_X1 U921 ( .A1(n1259), .A2(n1260), .ZN(n1238) );
NAND2_X1 U922 ( .A1(n1057), .A2(n1261), .ZN(n1260) );
NAND3_X1 U923 ( .A1(n1262), .A2(n1263), .A3(KEYINPUT14), .ZN(n1259) );
XNOR2_X1 U924 ( .A(G116), .B(n1212), .ZN(G18) );
NAND3_X1 U925 ( .A1(n1068), .A2(n1083), .A3(n1257), .ZN(n1212) );
NOR2_X1 U926 ( .A1(n1096), .A2(n1264), .ZN(n1068) );
XNOR2_X1 U927 ( .A(n1265), .B(n1266), .ZN(G15) );
NOR3_X1 U928 ( .A1(n1226), .A2(KEYINPUT18), .A3(n1267), .ZN(n1266) );
INV_X1 U929 ( .A(n1257), .ZN(n1267) );
NOR2_X1 U930 ( .A1(n1067), .A2(n1220), .ZN(n1257) );
INV_X1 U931 ( .A(n1229), .ZN(n1067) );
NOR2_X1 U932 ( .A1(n1076), .A2(n1107), .ZN(n1229) );
INV_X1 U933 ( .A(n1075), .ZN(n1107) );
NAND2_X1 U934 ( .A1(n1069), .A2(n1083), .ZN(n1226) );
NAND2_X1 U935 ( .A1(n1268), .A2(n1269), .ZN(n1083) );
NAND2_X1 U936 ( .A1(n1072), .A2(n1261), .ZN(n1269) );
INV_X1 U937 ( .A(KEYINPUT14), .ZN(n1261) );
NOR2_X1 U938 ( .A1(n1263), .A2(n1262), .ZN(n1072) );
INV_X1 U939 ( .A(n1270), .ZN(n1262) );
NAND3_X1 U940 ( .A1(n1270), .A2(n1263), .A3(KEYINPUT14), .ZN(n1268) );
INV_X1 U941 ( .A(n1217), .ZN(n1069) );
NAND2_X1 U942 ( .A1(n1264), .A2(n1096), .ZN(n1217) );
XNOR2_X1 U943 ( .A(G110), .B(n1271), .ZN(G12) );
NAND4_X1 U944 ( .A1(n1272), .A2(KEYINPUT63), .A3(n1073), .A4(n1218), .ZN(n1271) );
NOR2_X1 U945 ( .A1(n1064), .A2(n1220), .ZN(n1218) );
NAND2_X1 U946 ( .A1(n1256), .A2(n1273), .ZN(n1220) );
NAND2_X1 U947 ( .A1(n1059), .A2(n1274), .ZN(n1273) );
NAND3_X1 U948 ( .A1(n1152), .A2(n1255), .A3(G902), .ZN(n1274) );
NOR2_X1 U949 ( .A1(n1078), .A2(G898), .ZN(n1152) );
NAND3_X1 U950 ( .A1(n1255), .A2(n1078), .A3(G952), .ZN(n1059) );
NAND2_X1 U951 ( .A1(G237), .A2(G234), .ZN(n1255) );
NOR2_X1 U952 ( .A1(n1087), .A2(n1088), .ZN(n1256) );
NOR2_X1 U953 ( .A1(n1275), .A2(n1105), .ZN(n1088) );
NOR3_X1 U954 ( .A1(n1276), .A2(G902), .A3(n1277), .ZN(n1105) );
AND2_X1 U955 ( .A1(G237), .A2(n1278), .ZN(n1276) );
XNOR2_X1 U956 ( .A(KEYINPUT32), .B(n1106), .ZN(n1275) );
AND2_X1 U957 ( .A1(n1278), .A2(n1279), .ZN(n1106) );
NAND2_X1 U958 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U959 ( .A1(n1277), .A2(G237), .ZN(n1281) );
XNOR2_X1 U960 ( .A(n1206), .B(n1282), .ZN(n1277) );
XNOR2_X1 U961 ( .A(n1283), .B(KEYINPUT50), .ZN(n1282) );
NAND2_X1 U962 ( .A1(KEYINPUT53), .A2(G125), .ZN(n1283) );
XNOR2_X1 U963 ( .A(n1284), .B(n1285), .ZN(n1206) );
XOR2_X1 U964 ( .A(n1154), .B(n1153), .Z(n1285) );
XOR2_X1 U965 ( .A(G122), .B(G110), .Z(n1153) );
XNOR2_X1 U966 ( .A(n1286), .B(n1287), .ZN(n1154) );
XOR2_X1 U967 ( .A(n1288), .B(n1289), .Z(n1286) );
NOR2_X1 U968 ( .A1(G113), .A2(KEYINPUT8), .ZN(n1289) );
NAND2_X1 U969 ( .A1(n1290), .A2(n1291), .ZN(n1288) );
NAND2_X1 U970 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND2_X1 U971 ( .A1(G101), .A2(n1294), .ZN(n1293) );
OR2_X1 U972 ( .A1(KEYINPUT4), .A2(KEYINPUT58), .ZN(n1294) );
NAND3_X1 U973 ( .A1(n1295), .A2(n1296), .A3(KEYINPUT58), .ZN(n1290) );
OR2_X1 U974 ( .A1(G101), .A2(KEYINPUT4), .ZN(n1296) );
NAND2_X1 U975 ( .A1(G101), .A2(n1297), .ZN(n1295) );
OR2_X1 U976 ( .A1(n1292), .A2(KEYINPUT4), .ZN(n1297) );
XOR2_X1 U977 ( .A(n1298), .B(n1299), .Z(n1284) );
NOR2_X1 U978 ( .A1(G953), .A2(n1142), .ZN(n1299) );
INV_X1 U979 ( .A(G224), .ZN(n1142) );
XNOR2_X1 U980 ( .A(n1210), .B(KEYINPUT10), .ZN(n1278) );
INV_X1 U981 ( .A(G210), .ZN(n1210) );
INV_X1 U982 ( .A(n1091), .ZN(n1087) );
NAND2_X1 U983 ( .A1(G214), .A2(n1300), .ZN(n1091) );
OR2_X1 U984 ( .A1(G237), .A2(G902), .ZN(n1300) );
NAND2_X1 U985 ( .A1(n1076), .A2(n1075), .ZN(n1064) );
NAND2_X1 U986 ( .A1(G221), .A2(n1301), .ZN(n1075) );
XOR2_X1 U987 ( .A(n1099), .B(n1199), .Z(n1076) );
INV_X1 U988 ( .A(G469), .ZN(n1199) );
NAND2_X1 U989 ( .A1(n1302), .A2(n1280), .ZN(n1099) );
XOR2_X1 U990 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U991 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U992 ( .A(KEYINPUT46), .B(KEYINPUT1), .ZN(n1306) );
NAND4_X1 U993 ( .A1(n1307), .A2(n1308), .A3(n1309), .A4(n1310), .ZN(n1305) );
NAND2_X1 U994 ( .A1(KEYINPUT41), .A2(n1311), .ZN(n1310) );
NAND3_X1 U995 ( .A1(n1312), .A2(n1313), .A3(G110), .ZN(n1309) );
INV_X1 U996 ( .A(KEYINPUT41), .ZN(n1313) );
XNOR2_X1 U997 ( .A(KEYINPUT55), .B(G140), .ZN(n1312) );
NAND3_X1 U998 ( .A1(KEYINPUT62), .A2(n1314), .A3(n1245), .ZN(n1308) );
NAND2_X1 U999 ( .A1(G110), .A2(KEYINPUT55), .ZN(n1314) );
NAND3_X1 U1000 ( .A1(n1315), .A2(n1316), .A3(G140), .ZN(n1307) );
INV_X1 U1001 ( .A(KEYINPUT62), .ZN(n1316) );
OR2_X1 U1002 ( .A1(n1311), .A2(KEYINPUT55), .ZN(n1315) );
XNOR2_X1 U1003 ( .A(n1317), .B(n1204), .ZN(n1303) );
XOR2_X1 U1004 ( .A(n1127), .B(G146), .Z(n1204) );
XOR2_X1 U1005 ( .A(n1318), .B(n1319), .Z(n1127) );
XNOR2_X1 U1006 ( .A(KEYINPUT59), .B(KEYINPUT11), .ZN(n1318) );
XNOR2_X1 U1007 ( .A(n1320), .B(n1202), .ZN(n1317) );
XNOR2_X1 U1008 ( .A(n1292), .B(n1321), .ZN(n1202) );
XOR2_X1 U1009 ( .A(G101), .B(n1322), .Z(n1321) );
AND2_X1 U1010 ( .A1(n1078), .A2(G227), .ZN(n1322) );
INV_X1 U1011 ( .A(G953), .ZN(n1078) );
XNOR2_X1 U1012 ( .A(G104), .B(G107), .ZN(n1292) );
NOR2_X1 U1013 ( .A1(n1244), .A2(n1096), .ZN(n1073) );
XOR2_X1 U1014 ( .A(n1323), .B(n1176), .Z(n1096) );
INV_X1 U1015 ( .A(G475), .ZN(n1176) );
NAND2_X1 U1016 ( .A1(n1174), .A2(n1280), .ZN(n1323) );
XNOR2_X1 U1017 ( .A(n1324), .B(n1325), .ZN(n1174) );
XNOR2_X1 U1018 ( .A(n1326), .B(n1126), .ZN(n1325) );
XOR2_X1 U1019 ( .A(n1201), .B(n1327), .Z(n1126) );
XNOR2_X1 U1020 ( .A(G131), .B(n1245), .ZN(n1201) );
NAND2_X1 U1021 ( .A1(KEYINPUT33), .A2(n1328), .ZN(n1326) );
XNOR2_X1 U1022 ( .A(G143), .B(n1329), .ZN(n1328) );
NAND2_X1 U1023 ( .A1(G214), .A2(n1330), .ZN(n1329) );
XNOR2_X1 U1024 ( .A(G104), .B(n1331), .ZN(n1324) );
XNOR2_X1 U1025 ( .A(n1332), .B(G113), .ZN(n1331) );
INV_X1 U1026 ( .A(n1264), .ZN(n1244) );
XNOR2_X1 U1027 ( .A(n1104), .B(G478), .ZN(n1264) );
AND2_X1 U1028 ( .A1(n1166), .A2(n1280), .ZN(n1104) );
XOR2_X1 U1029 ( .A(n1333), .B(n1334), .Z(n1166) );
NOR3_X1 U1030 ( .A1(n1335), .A2(G953), .A3(n1336), .ZN(n1334) );
INV_X1 U1031 ( .A(G217), .ZN(n1335) );
NAND2_X1 U1032 ( .A1(n1337), .A2(n1338), .ZN(n1333) );
OR2_X1 U1033 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
XOR2_X1 U1034 ( .A(n1341), .B(KEYINPUT57), .Z(n1337) );
NAND2_X1 U1035 ( .A1(n1340), .A2(n1339), .ZN(n1341) );
NAND2_X1 U1036 ( .A1(n1342), .A2(n1343), .ZN(n1339) );
NAND2_X1 U1037 ( .A1(G107), .A2(n1344), .ZN(n1343) );
XOR2_X1 U1038 ( .A(n1345), .B(KEYINPUT12), .Z(n1342) );
OR2_X1 U1039 ( .A1(n1344), .A2(G107), .ZN(n1345) );
XNOR2_X1 U1040 ( .A(G116), .B(n1332), .ZN(n1344) );
INV_X1 U1041 ( .A(G122), .ZN(n1332) );
XOR2_X1 U1042 ( .A(G134), .B(n1319), .Z(n1340) );
XNOR2_X1 U1043 ( .A(G128), .B(n1346), .ZN(n1319) );
XNOR2_X1 U1044 ( .A(n1057), .B(KEYINPUT24), .ZN(n1272) );
NOR2_X1 U1045 ( .A1(n1270), .A2(n1263), .ZN(n1057) );
NAND2_X1 U1046 ( .A1(n1347), .A2(n1348), .ZN(n1263) );
NAND2_X1 U1047 ( .A1(G472), .A2(n1098), .ZN(n1348) );
XOR2_X1 U1048 ( .A(n1349), .B(KEYINPUT48), .Z(n1347) );
OR2_X1 U1049 ( .A1(n1098), .A2(G472), .ZN(n1349) );
NAND2_X1 U1050 ( .A1(n1350), .A2(n1280), .ZN(n1098) );
XOR2_X1 U1051 ( .A(n1351), .B(n1352), .Z(n1350) );
XNOR2_X1 U1052 ( .A(n1186), .B(n1189), .ZN(n1352) );
XNOR2_X1 U1053 ( .A(n1353), .B(G101), .ZN(n1189) );
NAND2_X1 U1054 ( .A1(G210), .A2(n1330), .ZN(n1353) );
NOR2_X1 U1055 ( .A1(G953), .A2(G237), .ZN(n1330) );
XOR2_X1 U1056 ( .A(n1298), .B(n1354), .Z(n1186) );
INV_X1 U1057 ( .A(n1320), .ZN(n1354) );
XOR2_X1 U1058 ( .A(n1198), .B(n1250), .Z(n1320) );
INV_X1 U1059 ( .A(G131), .ZN(n1250) );
NAND4_X1 U1060 ( .A1(n1355), .A2(n1356), .A3(n1357), .A4(n1358), .ZN(n1198) );
NAND3_X1 U1061 ( .A1(n1359), .A2(n1124), .A3(n1360), .ZN(n1358) );
INV_X1 U1062 ( .A(KEYINPUT19), .ZN(n1360) );
XOR2_X1 U1063 ( .A(KEYINPUT16), .B(G137), .Z(n1359) );
NAND2_X1 U1064 ( .A1(G134), .A2(KEYINPUT19), .ZN(n1357) );
OR3_X1 U1065 ( .A1(n1361), .A2(G137), .A3(KEYINPUT27), .ZN(n1356) );
NOR2_X1 U1066 ( .A1(KEYINPUT16), .A2(G134), .ZN(n1361) );
NAND3_X1 U1067 ( .A1(G137), .A2(n1362), .A3(KEYINPUT27), .ZN(n1355) );
NAND2_X1 U1068 ( .A1(KEYINPUT16), .A2(n1124), .ZN(n1362) );
INV_X1 U1069 ( .A(G134), .ZN(n1124) );
XOR2_X1 U1070 ( .A(n1363), .B(G128), .Z(n1298) );
NAND3_X1 U1071 ( .A1(n1364), .A2(n1365), .A3(n1366), .ZN(n1363) );
OR2_X1 U1072 ( .A1(n1346), .A2(KEYINPUT15), .ZN(n1366) );
NAND3_X1 U1073 ( .A1(KEYINPUT15), .A2(n1346), .A3(G146), .ZN(n1365) );
INV_X1 U1074 ( .A(G143), .ZN(n1346) );
NAND2_X1 U1075 ( .A1(n1367), .A2(n1368), .ZN(n1364) );
NAND2_X1 U1076 ( .A1(n1369), .A2(KEYINPUT15), .ZN(n1367) );
XNOR2_X1 U1077 ( .A(G143), .B(KEYINPUT25), .ZN(n1369) );
XOR2_X1 U1078 ( .A(n1370), .B(KEYINPUT23), .Z(n1351) );
NAND2_X1 U1079 ( .A1(KEYINPUT39), .A2(n1185), .ZN(n1370) );
XOR2_X1 U1080 ( .A(n1371), .B(n1287), .Z(n1185) );
XOR2_X1 U1081 ( .A(G116), .B(G119), .Z(n1287) );
NAND2_X1 U1082 ( .A1(KEYINPUT30), .A2(n1265), .ZN(n1371) );
INV_X1 U1083 ( .A(G113), .ZN(n1265) );
XOR2_X1 U1084 ( .A(n1372), .B(n1111), .Z(n1270) );
NAND2_X1 U1085 ( .A1(G217), .A2(n1301), .ZN(n1111) );
NAND2_X1 U1086 ( .A1(G234), .A2(n1280), .ZN(n1301) );
INV_X1 U1087 ( .A(G902), .ZN(n1280) );
XNOR2_X1 U1088 ( .A(n1108), .B(KEYINPUT31), .ZN(n1372) );
NOR2_X1 U1089 ( .A1(n1162), .A2(G902), .ZN(n1108) );
XNOR2_X1 U1090 ( .A(n1373), .B(n1374), .ZN(n1162) );
XOR2_X1 U1091 ( .A(n1375), .B(n1376), .Z(n1374) );
XOR2_X1 U1092 ( .A(n1377), .B(n1378), .Z(n1376) );
NOR3_X1 U1093 ( .A1(n1379), .A2(G953), .A3(n1336), .ZN(n1378) );
XNOR2_X1 U1094 ( .A(G234), .B(KEYINPUT52), .ZN(n1336) );
INV_X1 U1095 ( .A(G221), .ZN(n1379) );
NAND2_X1 U1096 ( .A1(KEYINPUT0), .A2(n1380), .ZN(n1377) );
XNOR2_X1 U1097 ( .A(n1245), .B(n1327), .ZN(n1380) );
XNOR2_X1 U1098 ( .A(G125), .B(n1368), .ZN(n1327) );
INV_X1 U1099 ( .A(G146), .ZN(n1368) );
INV_X1 U1100 ( .A(G140), .ZN(n1245) );
NAND2_X1 U1101 ( .A1(KEYINPUT34), .A2(n1311), .ZN(n1375) );
INV_X1 U1102 ( .A(G110), .ZN(n1311) );
XNOR2_X1 U1103 ( .A(G119), .B(n1381), .ZN(n1373) );
XOR2_X1 U1104 ( .A(G137), .B(G128), .Z(n1381) );
endmodule


