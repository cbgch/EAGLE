//Key = 0010011100100101000001110100000011111001000000001110001001110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337;

XOR2_X1 U732 ( .A(G107), .B(n1018), .Z(G9) );
NOR2_X1 U733 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR2_X1 U734 ( .A1(n1021), .A2(n1022), .ZN(G75) );
NOR3_X1 U735 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NOR3_X1 U736 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1024) );
NOR2_X1 U737 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NOR3_X1 U738 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
NOR2_X1 U739 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
AND2_X1 U740 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR3_X1 U741 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1034) );
NOR3_X1 U742 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NOR2_X1 U743 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U744 ( .A1(n1046), .A2(n1047), .ZN(n1039) );
XNOR2_X1 U745 ( .A(KEYINPUT16), .B(n1048), .ZN(n1046) );
NOR3_X1 U746 ( .A1(n1049), .A2(n1050), .A3(n1048), .ZN(n1029) );
NOR2_X1 U747 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U748 ( .A1(n1053), .A2(n1033), .ZN(n1052) );
NOR2_X1 U749 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U750 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U751 ( .A1(KEYINPUT53), .A2(n1020), .ZN(n1054) );
NOR2_X1 U752 ( .A1(n1058), .A2(n1031), .ZN(n1051) );
NOR2_X1 U753 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
INV_X1 U754 ( .A(n1061), .ZN(n1027) );
NAND3_X1 U755 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1023) );
NAND3_X1 U756 ( .A1(n1065), .A2(n1066), .A3(KEYINPUT53), .ZN(n1064) );
NAND4_X1 U757 ( .A1(n1067), .A2(n1061), .A3(n1036), .A4(n1068), .ZN(n1066) );
NOR2_X1 U758 ( .A1(n1049), .A2(n1026), .ZN(n1068) );
INV_X1 U759 ( .A(KEYINPUT5), .ZN(n1026) );
INV_X1 U760 ( .A(n1069), .ZN(n1049) );
AND3_X1 U761 ( .A1(n1062), .A2(n1063), .A3(n1070), .ZN(n1021) );
NAND4_X1 U762 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1062) );
NOR4_X1 U763 ( .A1(n1075), .A2(n1041), .A3(n1076), .A4(n1045), .ZN(n1074) );
XNOR2_X1 U764 ( .A(n1077), .B(KEYINPUT49), .ZN(n1076) );
NOR2_X1 U765 ( .A1(n1078), .A2(n1079), .ZN(n1073) );
XNOR2_X1 U766 ( .A(n1080), .B(n1081), .ZN(n1079) );
NOR2_X1 U767 ( .A1(KEYINPUT26), .A2(n1082), .ZN(n1081) );
XOR2_X1 U768 ( .A(n1083), .B(G475), .Z(n1072) );
XNOR2_X1 U769 ( .A(n1038), .B(KEYINPUT14), .ZN(n1071) );
XOR2_X1 U770 ( .A(n1084), .B(n1085), .Z(G72) );
XOR2_X1 U771 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U772 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NOR2_X1 U773 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND3_X1 U774 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1086) );
INV_X1 U775 ( .A(n1094), .ZN(n1093) );
NAND2_X1 U776 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
NAND2_X1 U777 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
NAND2_X1 U778 ( .A1(KEYINPUT39), .A2(n1099), .ZN(n1098) );
NAND2_X1 U779 ( .A1(n1100), .A2(n1101), .ZN(n1097) );
INV_X1 U780 ( .A(KEYINPUT39), .ZN(n1101) );
OR2_X1 U781 ( .A1(n1096), .A2(n1099), .ZN(n1091) );
NAND2_X1 U782 ( .A1(KEYINPUT48), .A2(n1100), .ZN(n1099) );
XOR2_X1 U783 ( .A(G140), .B(n1102), .Z(n1100) );
NOR2_X1 U784 ( .A1(G125), .A2(KEYINPUT41), .ZN(n1102) );
XOR2_X1 U785 ( .A(n1103), .B(n1104), .Z(n1096) );
XNOR2_X1 U786 ( .A(n1105), .B(G131), .ZN(n1104) );
INV_X1 U787 ( .A(G134), .ZN(n1105) );
XOR2_X1 U788 ( .A(n1106), .B(n1107), .Z(n1103) );
NAND2_X1 U789 ( .A1(G953), .A2(n1108), .ZN(n1084) );
NAND2_X1 U790 ( .A1(G900), .A2(G227), .ZN(n1108) );
NAND2_X1 U791 ( .A1(n1109), .A2(n1110), .ZN(G69) );
NAND2_X1 U792 ( .A1(G953), .A2(n1111), .ZN(n1110) );
XOR2_X1 U793 ( .A(n1112), .B(n1113), .Z(n1109) );
NOR2_X1 U794 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U795 ( .A1(G953), .A2(n1116), .ZN(n1115) );
NOR2_X1 U796 ( .A1(G224), .A2(n1063), .ZN(n1114) );
NOR2_X1 U797 ( .A1(KEYINPUT63), .A2(n1117), .ZN(n1112) );
XOR2_X1 U798 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U799 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
XOR2_X1 U800 ( .A(n1122), .B(KEYINPUT34), .Z(n1121) );
NAND2_X1 U801 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U802 ( .A1(n1124), .A2(n1123), .ZN(n1120) );
XOR2_X1 U803 ( .A(n1125), .B(KEYINPUT40), .Z(n1123) );
NOR2_X1 U804 ( .A1(n1126), .A2(n1127), .ZN(G66) );
XOR2_X1 U805 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U806 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
NOR3_X1 U807 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(G63) );
AND2_X1 U808 ( .A1(KEYINPUT10), .A2(n1126), .ZN(n1134) );
NOR3_X1 U809 ( .A1(KEYINPUT10), .A2(n1063), .A3(n1070), .ZN(n1133) );
INV_X1 U810 ( .A(G952), .ZN(n1070) );
XOR2_X1 U811 ( .A(n1135), .B(n1136), .Z(n1132) );
AND2_X1 U812 ( .A1(G478), .A2(n1137), .ZN(n1136) );
NAND2_X1 U813 ( .A1(KEYINPUT57), .A2(n1138), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(G60) );
XOR2_X1 U815 ( .A(KEYINPUT46), .B(n1126), .Z(n1140) );
NOR2_X1 U816 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
XOR2_X1 U817 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND3_X1 U818 ( .A1(n1145), .A2(n1025), .A3(G475), .ZN(n1144) );
XNOR2_X1 U819 ( .A(KEYINPUT52), .B(n1146), .ZN(n1145) );
NAND2_X1 U820 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
NOR2_X1 U821 ( .A1(n1147), .A2(n1148), .ZN(n1141) );
INV_X1 U822 ( .A(KEYINPUT9), .ZN(n1148) );
XOR2_X1 U823 ( .A(n1149), .B(KEYINPUT17), .Z(n1147) );
XOR2_X1 U824 ( .A(G104), .B(n1150), .Z(G6) );
NOR2_X1 U825 ( .A1(n1126), .A2(n1151), .ZN(G57) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U827 ( .A(n1154), .B(n1155), .Z(n1153) );
XNOR2_X1 U828 ( .A(n1156), .B(n1157), .ZN(n1155) );
XOR2_X1 U829 ( .A(n1158), .B(n1159), .Z(n1152) );
XOR2_X1 U830 ( .A(n1160), .B(n1161), .Z(n1159) );
AND2_X1 U831 ( .A1(G472), .A2(n1137), .ZN(n1160) );
NOR2_X1 U832 ( .A1(n1126), .A2(n1162), .ZN(G54) );
XOR2_X1 U833 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U834 ( .A(n1165), .B(n1166), .Z(n1164) );
AND2_X1 U835 ( .A1(G469), .A2(n1137), .ZN(n1165) );
XOR2_X1 U836 ( .A(n1167), .B(n1168), .Z(n1163) );
XNOR2_X1 U837 ( .A(KEYINPUT19), .B(n1169), .ZN(n1168) );
NOR2_X1 U838 ( .A1(KEYINPUT28), .A2(n1170), .ZN(n1167) );
XOR2_X1 U839 ( .A(n1171), .B(KEYINPUT36), .Z(n1170) );
NOR2_X1 U840 ( .A1(n1126), .A2(n1172), .ZN(G51) );
XOR2_X1 U841 ( .A(n1173), .B(n1174), .Z(n1172) );
NAND3_X1 U842 ( .A1(KEYINPUT25), .A2(n1137), .A3(n1175), .ZN(n1174) );
XNOR2_X1 U843 ( .A(G210), .B(KEYINPUT58), .ZN(n1175) );
INV_X1 U844 ( .A(n1131), .ZN(n1137) );
NAND2_X1 U845 ( .A1(G902), .A2(n1025), .ZN(n1131) );
NAND3_X1 U846 ( .A1(n1176), .A2(n1116), .A3(n1177), .ZN(n1025) );
XOR2_X1 U847 ( .A(n1089), .B(KEYINPUT50), .Z(n1177) );
NAND4_X1 U848 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1089) );
NAND2_X1 U849 ( .A1(n1182), .A2(n1183), .ZN(n1178) );
XNOR2_X1 U850 ( .A(n1059), .B(KEYINPUT13), .ZN(n1182) );
AND4_X1 U851 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1116) );
NOR4_X1 U852 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1150), .ZN(n1187) );
AND4_X1 U853 ( .A1(n1036), .A2(n1191), .A3(n1037), .A4(n1192), .ZN(n1150) );
NOR2_X1 U854 ( .A1(n1020), .A2(n1193), .ZN(n1192) );
INV_X1 U855 ( .A(n1194), .ZN(n1189) );
NOR2_X1 U856 ( .A1(n1195), .A2(n1196), .ZN(n1186) );
NOR2_X1 U857 ( .A1(n1197), .A2(n1020), .ZN(n1196) );
XOR2_X1 U858 ( .A(n1019), .B(KEYINPUT56), .Z(n1197) );
NAND4_X1 U859 ( .A1(n1037), .A2(n1036), .A3(n1059), .A4(n1191), .ZN(n1019) );
INV_X1 U860 ( .A(n1090), .ZN(n1176) );
NAND3_X1 U861 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1090) );
NAND2_X1 U862 ( .A1(n1183), .A2(n1060), .ZN(n1200) );
INV_X1 U863 ( .A(n1201), .ZN(n1183) );
OR2_X1 U864 ( .A1(n1202), .A2(n1203), .ZN(n1199) );
NAND2_X1 U865 ( .A1(n1204), .A2(n1205), .ZN(n1198) );
NAND2_X1 U866 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U867 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XOR2_X1 U868 ( .A(n1210), .B(KEYINPUT20), .Z(n1206) );
NAND2_X1 U869 ( .A1(n1211), .A2(n1212), .ZN(n1173) );
NAND2_X1 U870 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XOR2_X1 U871 ( .A(KEYINPUT61), .B(n1215), .Z(n1211) );
NOR2_X1 U872 ( .A1(n1213), .A2(n1214), .ZN(n1215) );
XOR2_X1 U873 ( .A(n1216), .B(n1217), .Z(n1213) );
XNOR2_X1 U874 ( .A(n1218), .B(KEYINPUT24), .ZN(n1217) );
NAND2_X1 U875 ( .A1(KEYINPUT35), .A2(n1156), .ZN(n1218) );
NOR2_X1 U876 ( .A1(n1063), .A2(G952), .ZN(n1126) );
XNOR2_X1 U877 ( .A(n1219), .B(n1220), .ZN(G48) );
NOR2_X1 U878 ( .A1(n1193), .A2(n1201), .ZN(n1220) );
XNOR2_X1 U879 ( .A(n1221), .B(n1222), .ZN(G45) );
NOR2_X1 U880 ( .A1(n1223), .A2(n1202), .ZN(n1222) );
NAND4_X1 U881 ( .A1(n1209), .A2(n1065), .A3(n1224), .A4(n1078), .ZN(n1202) );
XNOR2_X1 U882 ( .A(n1042), .B(KEYINPUT18), .ZN(n1223) );
XOR2_X1 U883 ( .A(G140), .B(n1225), .Z(G42) );
NOR2_X1 U884 ( .A1(n1210), .A2(n1031), .ZN(n1225) );
INV_X1 U885 ( .A(n1204), .ZN(n1031) );
NAND2_X1 U886 ( .A1(n1226), .A2(n1209), .ZN(n1210) );
XNOR2_X1 U887 ( .A(G137), .B(n1227), .ZN(G39) );
NAND4_X1 U888 ( .A1(n1228), .A2(n1204), .A3(n1208), .A4(n1037), .ZN(n1227) );
XOR2_X1 U889 ( .A(n1229), .B(KEYINPUT4), .Z(n1228) );
XNOR2_X1 U890 ( .A(G134), .B(n1179), .ZN(G36) );
NAND2_X1 U891 ( .A1(n1230), .A2(n1059), .ZN(n1179) );
XNOR2_X1 U892 ( .A(G131), .B(n1180), .ZN(G33) );
NAND2_X1 U893 ( .A1(n1230), .A2(n1060), .ZN(n1180) );
AND3_X1 U894 ( .A1(n1042), .A2(n1209), .A3(n1204), .ZN(n1230) );
NOR2_X1 U895 ( .A1(n1056), .A2(n1075), .ZN(n1204) );
INV_X1 U896 ( .A(n1057), .ZN(n1075) );
XOR2_X1 U897 ( .A(G128), .B(n1231), .Z(G30) );
NOR2_X1 U898 ( .A1(n1232), .A2(n1201), .ZN(n1231) );
NAND4_X1 U899 ( .A1(n1209), .A2(n1065), .A3(n1077), .A4(n1045), .ZN(n1201) );
AND2_X1 U900 ( .A1(n1037), .A2(n1229), .ZN(n1209) );
XNOR2_X1 U901 ( .A(n1157), .B(n1195), .ZN(G3) );
AND2_X1 U902 ( .A1(n1233), .A2(n1042), .ZN(n1195) );
XNOR2_X1 U903 ( .A(G125), .B(n1181), .ZN(G27) );
NAND4_X1 U904 ( .A1(n1069), .A2(n1226), .A3(n1065), .A4(n1229), .ZN(n1181) );
NAND2_X1 U905 ( .A1(n1234), .A2(n1235), .ZN(n1229) );
NAND3_X1 U906 ( .A1(G902), .A2(n1061), .A3(n1094), .ZN(n1235) );
NOR2_X1 U907 ( .A1(n1063), .A2(G900), .ZN(n1094) );
NOR3_X1 U908 ( .A1(n1045), .A2(n1044), .A3(n1193), .ZN(n1226) );
XNOR2_X1 U909 ( .A(G122), .B(n1184), .ZN(G24) );
NAND4_X1 U910 ( .A1(n1236), .A2(n1036), .A3(n1224), .A4(n1078), .ZN(n1184) );
INV_X1 U911 ( .A(n1237), .ZN(n1224) );
INV_X1 U912 ( .A(n1048), .ZN(n1036) );
NAND2_X1 U913 ( .A1(n1238), .A2(n1239), .ZN(n1048) );
XOR2_X1 U914 ( .A(n1190), .B(n1240), .Z(G21) );
NOR2_X1 U915 ( .A1(KEYINPUT1), .A2(n1241), .ZN(n1240) );
INV_X1 U916 ( .A(G119), .ZN(n1241) );
AND2_X1 U917 ( .A1(n1236), .A2(n1208), .ZN(n1190) );
NOR3_X1 U918 ( .A1(n1044), .A2(n1238), .A3(n1033), .ZN(n1208) );
INV_X1 U919 ( .A(n1067), .ZN(n1033) );
XNOR2_X1 U920 ( .A(G116), .B(n1194), .ZN(G18) );
NAND3_X1 U921 ( .A1(n1042), .A2(n1059), .A3(n1236), .ZN(n1194) );
INV_X1 U922 ( .A(n1232), .ZN(n1059) );
NAND2_X1 U923 ( .A1(n1242), .A2(n1078), .ZN(n1232) );
XNOR2_X1 U924 ( .A(KEYINPUT54), .B(n1237), .ZN(n1242) );
XOR2_X1 U925 ( .A(G113), .B(n1188), .Z(G15) );
AND3_X1 U926 ( .A1(n1060), .A2(n1042), .A3(n1236), .ZN(n1188) );
AND3_X1 U927 ( .A1(n1065), .A2(n1191), .A3(n1069), .ZN(n1236) );
NOR2_X1 U928 ( .A1(n1038), .A2(n1041), .ZN(n1069) );
INV_X1 U929 ( .A(n1203), .ZN(n1042) );
NAND2_X1 U930 ( .A1(n1239), .A2(n1045), .ZN(n1203) );
XNOR2_X1 U931 ( .A(KEYINPUT21), .B(n1044), .ZN(n1239) );
INV_X1 U932 ( .A(n1077), .ZN(n1044) );
XNOR2_X1 U933 ( .A(G110), .B(n1185), .ZN(G12) );
NAND3_X1 U934 ( .A1(n1238), .A2(n1077), .A3(n1233), .ZN(n1185) );
AND4_X1 U935 ( .A1(n1065), .A2(n1037), .A3(n1067), .A4(n1191), .ZN(n1233) );
NAND2_X1 U936 ( .A1(n1234), .A2(n1243), .ZN(n1191) );
NAND4_X1 U937 ( .A1(G953), .A2(G902), .A3(n1061), .A4(n1111), .ZN(n1243) );
INV_X1 U938 ( .A(G898), .ZN(n1111) );
NAND3_X1 U939 ( .A1(n1061), .A2(n1063), .A3(G952), .ZN(n1234) );
NAND2_X1 U940 ( .A1(G237), .A2(G234), .ZN(n1061) );
NAND2_X1 U941 ( .A1(n1244), .A2(n1245), .ZN(n1067) );
OR2_X1 U942 ( .A1(n1193), .A2(KEYINPUT54), .ZN(n1245) );
INV_X1 U943 ( .A(n1060), .ZN(n1193) );
NOR2_X1 U944 ( .A1(n1078), .A2(n1237), .ZN(n1060) );
NAND3_X1 U945 ( .A1(n1237), .A2(n1246), .A3(KEYINPUT54), .ZN(n1244) );
INV_X1 U946 ( .A(n1078), .ZN(n1246) );
XNOR2_X1 U947 ( .A(n1247), .B(G478), .ZN(n1078) );
NAND2_X1 U948 ( .A1(n1248), .A2(n1146), .ZN(n1247) );
XOR2_X1 U949 ( .A(n1138), .B(KEYINPUT30), .Z(n1248) );
XOR2_X1 U950 ( .A(n1249), .B(n1250), .Z(n1138) );
XOR2_X1 U951 ( .A(n1251), .B(n1252), .Z(n1250) );
NOR2_X1 U952 ( .A1(n1253), .A2(n1254), .ZN(n1251) );
INV_X1 U953 ( .A(G217), .ZN(n1253) );
XOR2_X1 U954 ( .A(n1255), .B(n1256), .Z(n1249) );
XNOR2_X1 U955 ( .A(n1221), .B(G134), .ZN(n1256) );
NAND2_X1 U956 ( .A1(n1257), .A2(n1258), .ZN(n1255) );
NAND2_X1 U957 ( .A1(G122), .A2(n1259), .ZN(n1258) );
XOR2_X1 U958 ( .A(KEYINPUT22), .B(n1260), .Z(n1257) );
NOR2_X1 U959 ( .A1(G122), .A2(n1259), .ZN(n1260) );
INV_X1 U960 ( .A(G116), .ZN(n1259) );
XNOR2_X1 U961 ( .A(n1261), .B(G475), .ZN(n1237) );
NAND2_X1 U962 ( .A1(n1262), .A2(n1083), .ZN(n1261) );
NAND2_X1 U963 ( .A1(n1149), .A2(n1146), .ZN(n1083) );
XOR2_X1 U964 ( .A(n1263), .B(n1264), .Z(n1149) );
XNOR2_X1 U965 ( .A(n1265), .B(n1266), .ZN(n1264) );
XOR2_X1 U966 ( .A(n1267), .B(n1268), .Z(n1266) );
NOR2_X1 U967 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
XOR2_X1 U968 ( .A(n1271), .B(KEYINPUT6), .Z(n1270) );
NAND2_X1 U969 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NOR2_X1 U970 ( .A1(n1273), .A2(n1272), .ZN(n1269) );
XNOR2_X1 U971 ( .A(n1274), .B(G143), .ZN(n1272) );
NAND2_X1 U972 ( .A1(n1275), .A2(G214), .ZN(n1274) );
INV_X1 U973 ( .A(G131), .ZN(n1273) );
NAND2_X1 U974 ( .A1(n1276), .A2(KEYINPUT23), .ZN(n1267) );
XNOR2_X1 U975 ( .A(G146), .B(n1277), .ZN(n1276) );
XNOR2_X1 U976 ( .A(G113), .B(n1278), .ZN(n1263) );
XOR2_X1 U977 ( .A(KEYINPUT59), .B(G122), .Z(n1278) );
XNOR2_X1 U978 ( .A(KEYINPUT37), .B(KEYINPUT12), .ZN(n1262) );
NOR2_X1 U979 ( .A1(n1279), .A2(n1041), .ZN(n1037) );
INV_X1 U980 ( .A(n1047), .ZN(n1041) );
NAND2_X1 U981 ( .A1(G221), .A2(n1280), .ZN(n1047) );
XNOR2_X1 U982 ( .A(KEYINPUT15), .B(n1281), .ZN(n1280) );
INV_X1 U983 ( .A(n1038), .ZN(n1279) );
XNOR2_X1 U984 ( .A(n1282), .B(G469), .ZN(n1038) );
NAND2_X1 U985 ( .A1(n1283), .A2(n1146), .ZN(n1282) );
XNOR2_X1 U986 ( .A(n1166), .B(n1284), .ZN(n1283) );
XOR2_X1 U987 ( .A(n1171), .B(n1285), .Z(n1284) );
NOR2_X1 U988 ( .A1(KEYINPUT29), .A2(n1169), .ZN(n1285) );
XOR2_X1 U989 ( .A(n1286), .B(n1287), .Z(n1171) );
XOR2_X1 U990 ( .A(n1106), .B(n1252), .Z(n1286) );
XOR2_X1 U991 ( .A(G107), .B(G128), .Z(n1252) );
XOR2_X1 U992 ( .A(n1288), .B(KEYINPUT44), .Z(n1106) );
NAND2_X1 U993 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
NAND2_X1 U994 ( .A1(G143), .A2(n1219), .ZN(n1290) );
XOR2_X1 U995 ( .A(KEYINPUT62), .B(n1291), .Z(n1289) );
NOR2_X1 U996 ( .A1(G143), .A2(n1219), .ZN(n1291) );
XNOR2_X1 U997 ( .A(n1158), .B(n1292), .ZN(n1166) );
XNOR2_X1 U998 ( .A(G140), .B(n1293), .ZN(n1292) );
NAND2_X1 U999 ( .A1(n1294), .A2(n1063), .ZN(n1293) );
XOR2_X1 U1000 ( .A(KEYINPUT38), .B(G227), .Z(n1294) );
INV_X1 U1001 ( .A(n1020), .ZN(n1065) );
NAND2_X1 U1002 ( .A1(n1056), .A2(n1057), .ZN(n1020) );
NAND2_X1 U1003 ( .A1(G214), .A2(n1295), .ZN(n1057) );
XOR2_X1 U1004 ( .A(n1080), .B(n1082), .Z(n1056) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1295), .ZN(n1082) );
NAND2_X1 U1006 ( .A1(n1296), .A2(n1146), .ZN(n1295) );
INV_X1 U1007 ( .A(G237), .ZN(n1296) );
NAND2_X1 U1008 ( .A1(n1297), .A2(n1146), .ZN(n1080) );
XOR2_X1 U1009 ( .A(n1216), .B(n1298), .Z(n1297) );
XNOR2_X1 U1010 ( .A(n1156), .B(n1299), .ZN(n1298) );
NOR2_X1 U1011 ( .A1(KEYINPUT8), .A2(n1300), .ZN(n1299) );
INV_X1 U1012 ( .A(n1214), .ZN(n1300) );
XOR2_X1 U1013 ( .A(n1119), .B(n1301), .Z(n1214) );
XOR2_X1 U1014 ( .A(n1124), .B(n1125), .Z(n1301) );
XNOR2_X1 U1015 ( .A(n1287), .B(G107), .ZN(n1125) );
XOR2_X1 U1016 ( .A(G101), .B(n1265), .Z(n1287) );
XOR2_X1 U1017 ( .A(G104), .B(KEYINPUT0), .Z(n1265) );
XOR2_X1 U1018 ( .A(n1302), .B(n1303), .Z(n1124) );
NOR2_X1 U1019 ( .A1(KEYINPUT31), .A2(n1304), .ZN(n1303) );
XNOR2_X1 U1020 ( .A(n1305), .B(KEYINPUT60), .ZN(n1304) );
XNOR2_X1 U1021 ( .A(n1169), .B(G122), .ZN(n1119) );
INV_X1 U1022 ( .A(G110), .ZN(n1169) );
XNOR2_X1 U1023 ( .A(G125), .B(n1306), .ZN(n1216) );
AND2_X1 U1024 ( .A1(n1063), .A2(G224), .ZN(n1306) );
XOR2_X1 U1025 ( .A(n1307), .B(n1130), .Z(n1077) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1281), .ZN(n1130) );
NAND2_X1 U1027 ( .A1(n1308), .A2(n1146), .ZN(n1281) );
XOR2_X1 U1028 ( .A(KEYINPUT27), .B(G234), .Z(n1308) );
OR2_X1 U1029 ( .A1(n1129), .A2(G902), .ZN(n1307) );
XNOR2_X1 U1030 ( .A(n1309), .B(n1310), .ZN(n1129) );
XNOR2_X1 U1031 ( .A(n1107), .B(n1311), .ZN(n1310) );
XOR2_X1 U1032 ( .A(n1312), .B(n1313), .Z(n1311) );
NOR2_X1 U1033 ( .A1(n1314), .A2(n1254), .ZN(n1313) );
NAND2_X1 U1034 ( .A1(n1315), .A2(n1063), .ZN(n1254) );
INV_X1 U1035 ( .A(G953), .ZN(n1063) );
XOR2_X1 U1036 ( .A(KEYINPUT45), .B(G234), .Z(n1315) );
INV_X1 U1037 ( .A(G221), .ZN(n1314) );
NAND2_X1 U1038 ( .A1(KEYINPUT2), .A2(n1277), .ZN(n1312) );
XOR2_X1 U1039 ( .A(G125), .B(G140), .Z(n1277) );
XOR2_X1 U1040 ( .A(G128), .B(n1316), .Z(n1107) );
XOR2_X1 U1041 ( .A(n1317), .B(n1318), .Z(n1309) );
XNOR2_X1 U1042 ( .A(KEYINPUT47), .B(n1219), .ZN(n1318) );
INV_X1 U1043 ( .A(G146), .ZN(n1219) );
XNOR2_X1 U1044 ( .A(G119), .B(G110), .ZN(n1317) );
INV_X1 U1045 ( .A(n1045), .ZN(n1238) );
XNOR2_X1 U1046 ( .A(n1319), .B(G472), .ZN(n1045) );
NAND2_X1 U1047 ( .A1(n1320), .A2(n1146), .ZN(n1319) );
INV_X1 U1048 ( .A(G902), .ZN(n1146) );
XOR2_X1 U1049 ( .A(n1321), .B(n1322), .Z(n1320) );
XNOR2_X1 U1050 ( .A(n1161), .B(n1158), .ZN(n1322) );
XOR2_X1 U1051 ( .A(n1323), .B(n1324), .Z(n1158) );
NOR2_X1 U1052 ( .A1(KEYINPUT3), .A2(n1325), .ZN(n1324) );
XNOR2_X1 U1053 ( .A(G134), .B(n1316), .ZN(n1325) );
XOR2_X1 U1054 ( .A(G137), .B(KEYINPUT32), .Z(n1316) );
XNOR2_X1 U1055 ( .A(G131), .B(KEYINPUT51), .ZN(n1323) );
XOR2_X1 U1056 ( .A(n1302), .B(n1326), .Z(n1161) );
INV_X1 U1057 ( .A(n1305), .ZN(n1326) );
XOR2_X1 U1058 ( .A(G116), .B(KEYINPUT55), .Z(n1305) );
XNOR2_X1 U1059 ( .A(G113), .B(G119), .ZN(n1302) );
XOR2_X1 U1060 ( .A(n1327), .B(n1328), .Z(n1321) );
XNOR2_X1 U1061 ( .A(n1154), .B(n1329), .ZN(n1328) );
NOR2_X1 U1062 ( .A1(KEYINPUT42), .A2(n1156), .ZN(n1329) );
NAND2_X1 U1063 ( .A1(n1330), .A2(n1331), .ZN(n1156) );
NAND2_X1 U1064 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
XOR2_X1 U1065 ( .A(KEYINPUT7), .B(n1334), .Z(n1333) );
XNOR2_X1 U1066 ( .A(KEYINPUT44), .B(G128), .ZN(n1332) );
NAND2_X1 U1067 ( .A1(n1335), .A2(n1336), .ZN(n1330) );
XOR2_X1 U1068 ( .A(KEYINPUT11), .B(n1334), .Z(n1336) );
XNOR2_X1 U1069 ( .A(n1337), .B(G146), .ZN(n1334) );
NAND2_X1 U1070 ( .A1(KEYINPUT33), .A2(n1221), .ZN(n1337) );
INV_X1 U1071 ( .A(G143), .ZN(n1221) );
XOR2_X1 U1072 ( .A(KEYINPUT44), .B(G128), .Z(n1335) );
NAND2_X1 U1073 ( .A1(n1275), .A2(G210), .ZN(n1154) );
NOR2_X1 U1074 ( .A1(G953), .A2(G237), .ZN(n1275) );
NOR2_X1 U1075 ( .A1(KEYINPUT43), .A2(n1157), .ZN(n1327) );
INV_X1 U1076 ( .A(G101), .ZN(n1157) );
endmodule


