//Key = 0111111000010001101000111001111001010101100010001100100101110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373;

XNOR2_X1 U752 ( .A(G107), .B(n1039), .ZN(G9) );
NAND2_X1 U753 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
XOR2_X1 U754 ( .A(n1042), .B(KEYINPUT2), .Z(n1040) );
NAND4_X1 U755 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
XNOR2_X1 U756 ( .A(n1047), .B(KEYINPUT28), .ZN(n1043) );
NAND4_X1 U757 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(G75) );
NAND2_X1 U758 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U759 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND3_X1 U760 ( .A1(n1056), .A2(n1057), .A3(n1047), .ZN(n1055) );
NAND3_X1 U761 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1056) );
NAND2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NAND2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U764 ( .A1(KEYINPUT58), .A2(n1045), .ZN(n1064) );
NAND2_X1 U765 ( .A1(n1065), .A2(n1066), .ZN(n1058) );
INV_X1 U766 ( .A(KEYINPUT26), .ZN(n1066) );
NAND3_X1 U767 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1054) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NAND4_X1 U769 ( .A1(n1072), .A2(n1073), .A3(n1047), .A4(n1057), .ZN(n1071) );
NAND3_X1 U770 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1057) );
NAND2_X1 U771 ( .A1(KEYINPUT26), .A2(n1065), .ZN(n1076) );
OR3_X1 U772 ( .A1(n1077), .A2(KEYINPUT58), .A3(n1078), .ZN(n1074) );
NAND2_X1 U773 ( .A1(n1061), .A2(n1079), .ZN(n1070) );
NAND2_X1 U774 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U775 ( .A1(n1060), .A2(n1082), .ZN(n1081) );
NAND2_X1 U776 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U777 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U778 ( .A1(n1047), .A2(n1087), .ZN(n1080) );
NAND2_X1 U779 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
OR2_X1 U780 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
INV_X1 U781 ( .A(n1092), .ZN(n1052) );
NOR2_X1 U782 ( .A1(G953), .A2(n1093), .ZN(n1050) );
NOR4_X1 U783 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1093) );
NAND3_X1 U784 ( .A1(n1090), .A2(n1098), .A3(n1099), .ZN(n1095) );
NAND2_X1 U785 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
XOR2_X1 U786 ( .A(KEYINPUT38), .B(G478), .Z(n1100) );
NAND4_X1 U787 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1094) );
XOR2_X1 U788 ( .A(n1106), .B(G469), .Z(n1105) );
NAND2_X1 U789 ( .A1(KEYINPUT11), .A2(n1107), .ZN(n1106) );
XNOR2_X1 U790 ( .A(n1108), .B(n1109), .ZN(n1104) );
XOR2_X1 U791 ( .A(n1110), .B(KEYINPUT14), .Z(n1103) );
XOR2_X1 U792 ( .A(n1111), .B(G472), .Z(n1102) );
XOR2_X1 U793 ( .A(n1112), .B(n1113), .Z(G72) );
NOR2_X1 U794 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U795 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NAND2_X1 U796 ( .A1(n1118), .A2(n1119), .ZN(n1112) );
NAND2_X1 U797 ( .A1(n1120), .A2(n1115), .ZN(n1119) );
XOR2_X1 U798 ( .A(n1048), .B(n1121), .Z(n1120) );
OR3_X1 U799 ( .A1(n1117), .A2(n1121), .A3(n1115), .ZN(n1118) );
XNOR2_X1 U800 ( .A(n1122), .B(n1123), .ZN(n1121) );
XOR2_X1 U801 ( .A(n1124), .B(n1125), .Z(n1123) );
XNOR2_X1 U802 ( .A(n1126), .B(n1127), .ZN(n1122) );
XNOR2_X1 U803 ( .A(n1128), .B(KEYINPUT17), .ZN(n1127) );
NAND2_X1 U804 ( .A1(KEYINPUT59), .A2(n1129), .ZN(n1128) );
XOR2_X1 U805 ( .A(n1130), .B(n1131), .Z(G69) );
XOR2_X1 U806 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U807 ( .A1(G953), .A2(n1134), .ZN(n1133) );
NAND2_X1 U808 ( .A1(G898), .A2(G224), .ZN(n1134) );
NAND2_X1 U809 ( .A1(n1135), .A2(n1136), .ZN(n1132) );
XOR2_X1 U810 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U811 ( .A(n1139), .B(KEYINPUT20), .Z(n1135) );
NAND2_X1 U812 ( .A1(G953), .A2(n1140), .ZN(n1139) );
NOR2_X1 U813 ( .A1(n1049), .A2(G953), .ZN(n1130) );
NOR2_X1 U814 ( .A1(n1141), .A2(n1142), .ZN(G66) );
XOR2_X1 U815 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U816 ( .A1(KEYINPUT45), .A2(n1145), .ZN(n1144) );
NOR2_X1 U817 ( .A1(n1146), .A2(n1147), .ZN(n1143) );
NOR2_X1 U818 ( .A1(n1141), .A2(n1148), .ZN(G63) );
XOR2_X1 U819 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U820 ( .A(KEYINPUT61), .B(n1151), .Z(n1150) );
NOR2_X1 U821 ( .A1(n1152), .A2(n1147), .ZN(n1151) );
INV_X1 U822 ( .A(G478), .ZN(n1152) );
NOR2_X1 U823 ( .A1(n1141), .A2(n1153), .ZN(G60) );
XOR2_X1 U824 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U825 ( .A1(n1156), .A2(n1147), .ZN(n1155) );
XOR2_X1 U826 ( .A(n1157), .B(n1158), .Z(G6) );
NOR2_X1 U827 ( .A1(n1141), .A2(n1159), .ZN(G57) );
XOR2_X1 U828 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U829 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U830 ( .A1(n1164), .A2(n1147), .ZN(n1163) );
INV_X1 U831 ( .A(G472), .ZN(n1164) );
NOR2_X1 U832 ( .A1(KEYINPUT53), .A2(n1165), .ZN(n1162) );
XOR2_X1 U833 ( .A(KEYINPUT31), .B(G101), .Z(n1165) );
XOR2_X1 U834 ( .A(n1166), .B(n1167), .Z(n1160) );
NOR2_X1 U835 ( .A1(n1141), .A2(n1168), .ZN(G54) );
XOR2_X1 U836 ( .A(n1169), .B(n1170), .Z(n1168) );
XNOR2_X1 U837 ( .A(n1171), .B(n1172), .ZN(n1170) );
NAND2_X1 U838 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NAND3_X1 U839 ( .A1(n1125), .A2(n1175), .A3(n1176), .ZN(n1174) );
INV_X1 U840 ( .A(KEYINPUT29), .ZN(n1176) );
NAND2_X1 U841 ( .A1(n1177), .A2(KEYINPUT29), .ZN(n1173) );
XOR2_X1 U842 ( .A(n1178), .B(n1179), .Z(n1169) );
XOR2_X1 U843 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U844 ( .A1(G140), .A2(KEYINPUT42), .ZN(n1181) );
NOR3_X1 U845 ( .A1(n1116), .A2(KEYINPUT46), .A3(G953), .ZN(n1180) );
NOR3_X1 U846 ( .A1(n1147), .A2(KEYINPUT10), .A3(n1182), .ZN(n1178) );
INV_X1 U847 ( .A(G469), .ZN(n1182) );
NOR2_X1 U848 ( .A1(n1141), .A2(n1183), .ZN(G51) );
XOR2_X1 U849 ( .A(n1184), .B(n1185), .Z(n1183) );
XOR2_X1 U850 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U851 ( .A(n1188), .B(n1189), .Z(n1187) );
NOR2_X1 U852 ( .A1(n1109), .A2(n1147), .ZN(n1186) );
NAND2_X1 U853 ( .A1(G902), .A2(n1190), .ZN(n1147) );
NAND2_X1 U854 ( .A1(n1049), .A2(n1191), .ZN(n1190) );
XOR2_X1 U855 ( .A(KEYINPUT36), .B(n1048), .Z(n1191) );
AND4_X1 U856 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1048) );
NOR4_X1 U857 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1195) );
NAND2_X1 U858 ( .A1(n1200), .A2(n1201), .ZN(n1194) );
NAND2_X1 U859 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NAND2_X1 U860 ( .A1(n1060), .A2(n1204), .ZN(n1203) );
XOR2_X1 U861 ( .A(KEYINPUT8), .B(n1044), .Z(n1204) );
NAND2_X1 U862 ( .A1(n1061), .A2(n1041), .ZN(n1202) );
OR3_X1 U863 ( .A1(n1205), .A2(n1206), .A3(n1063), .ZN(n1192) );
AND4_X1 U864 ( .A1(n1158), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1049) );
AND4_X1 U865 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1209) );
NAND2_X1 U866 ( .A1(n1045), .A2(n1214), .ZN(n1208) );
NAND2_X1 U867 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND3_X1 U868 ( .A1(n1044), .A2(n1047), .A3(n1217), .ZN(n1216) );
NAND2_X1 U869 ( .A1(n1218), .A2(n1219), .ZN(n1215) );
NAND4_X1 U870 ( .A1(n1217), .A2(n1220), .A3(n1044), .A4(n1047), .ZN(n1158) );
XOR2_X1 U871 ( .A(n1221), .B(n1222), .Z(n1184) );
NAND2_X1 U872 ( .A1(KEYINPUT1), .A2(n1223), .ZN(n1221) );
NOR2_X1 U873 ( .A1(n1115), .A2(G952), .ZN(n1141) );
XOR2_X1 U874 ( .A(G146), .B(n1224), .Z(G48) );
NOR3_X1 U875 ( .A1(n1063), .A2(n1225), .A3(n1205), .ZN(n1224) );
XOR2_X1 U876 ( .A(n1206), .B(KEYINPUT41), .Z(n1225) );
XOR2_X1 U877 ( .A(G143), .B(n1199), .Z(G45) );
NOR4_X1 U878 ( .A1(n1226), .A2(n1088), .A3(n1067), .A4(n1069), .ZN(n1199) );
INV_X1 U879 ( .A(n1041), .ZN(n1088) );
NAND3_X1 U880 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(G42) );
NAND2_X1 U881 ( .A1(KEYINPUT63), .A2(n1230), .ZN(n1229) );
OR3_X1 U882 ( .A1(n1230), .A2(KEYINPUT63), .A3(G140), .ZN(n1228) );
NAND2_X1 U883 ( .A1(G140), .A2(n1231), .ZN(n1227) );
NAND2_X1 U884 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
INV_X1 U885 ( .A(KEYINPUT63), .ZN(n1233) );
XOR2_X1 U886 ( .A(n1230), .B(KEYINPUT3), .Z(n1232) );
NAND2_X1 U887 ( .A1(n1234), .A2(n1060), .ZN(n1230) );
XOR2_X1 U888 ( .A(n1235), .B(KEYINPUT27), .Z(n1234) );
NAND2_X1 U889 ( .A1(n1200), .A2(n1044), .ZN(n1235) );
INV_X1 U890 ( .A(n1236), .ZN(n1200) );
XOR2_X1 U891 ( .A(G137), .B(n1198), .Z(G39) );
AND4_X1 U892 ( .A1(n1237), .A2(n1238), .A3(n1086), .A4(n1239), .ZN(n1198) );
AND2_X1 U893 ( .A1(n1060), .A2(n1065), .ZN(n1239) );
XNOR2_X1 U894 ( .A(G134), .B(n1240), .ZN(G36) );
NOR2_X1 U895 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
NOR2_X1 U896 ( .A1(n1243), .A2(n1193), .ZN(n1242) );
OR3_X1 U897 ( .A1(n1226), .A2(n1077), .A3(n1075), .ZN(n1193) );
INV_X1 U898 ( .A(KEYINPUT35), .ZN(n1243) );
NOR4_X1 U899 ( .A1(KEYINPUT35), .A2(n1226), .A3(n1060), .A4(n1077), .ZN(n1241) );
XOR2_X1 U900 ( .A(G131), .B(n1197), .Z(G33) );
NOR3_X1 U901 ( .A1(n1075), .A2(n1226), .A3(n1063), .ZN(n1197) );
NAND3_X1 U902 ( .A1(n1044), .A2(n1237), .A3(n1219), .ZN(n1226) );
INV_X1 U903 ( .A(n1060), .ZN(n1075) );
NOR2_X1 U904 ( .A1(n1244), .A2(n1091), .ZN(n1060) );
XOR2_X1 U905 ( .A(G128), .B(n1196), .Z(G30) );
NOR3_X1 U906 ( .A1(n1206), .A2(n1077), .A3(n1205), .ZN(n1196) );
NAND4_X1 U907 ( .A1(n1041), .A2(n1086), .A3(n1237), .A4(n1238), .ZN(n1205) );
XOR2_X1 U908 ( .A(n1207), .B(n1245), .Z(G3) );
XOR2_X1 U909 ( .A(KEYINPUT44), .B(G101), .Z(n1245) );
NAND3_X1 U910 ( .A1(n1065), .A2(n1219), .A3(n1217), .ZN(n1207) );
NAND2_X1 U911 ( .A1(n1246), .A2(n1247), .ZN(G27) );
NAND2_X1 U912 ( .A1(G125), .A2(n1248), .ZN(n1247) );
XOR2_X1 U913 ( .A(n1249), .B(KEYINPUT19), .Z(n1246) );
OR2_X1 U914 ( .A1(n1248), .A2(G125), .ZN(n1249) );
NAND2_X1 U915 ( .A1(n1041), .A2(n1250), .ZN(n1248) );
XOR2_X1 U916 ( .A(KEYINPUT50), .B(n1251), .Z(n1250) );
NOR2_X1 U917 ( .A1(n1078), .A2(n1236), .ZN(n1251) );
NAND4_X1 U918 ( .A1(n1220), .A2(n1085), .A3(n1086), .A4(n1237), .ZN(n1236) );
NAND2_X1 U919 ( .A1(n1092), .A2(n1252), .ZN(n1237) );
NAND4_X1 U920 ( .A1(G953), .A2(n1253), .A3(n1254), .A4(n1117), .ZN(n1252) );
INV_X1 U921 ( .A(G900), .ZN(n1117) );
XOR2_X1 U922 ( .A(KEYINPUT34), .B(G902), .Z(n1253) );
XNOR2_X1 U923 ( .A(G122), .B(n1213), .ZN(G24) );
NAND4_X1 U924 ( .A1(n1218), .A2(n1047), .A3(n1097), .A4(n1255), .ZN(n1213) );
NOR2_X1 U925 ( .A1(n1238), .A2(n1086), .ZN(n1047) );
XOR2_X1 U926 ( .A(n1212), .B(n1256), .Z(G21) );
NAND2_X1 U927 ( .A1(KEYINPUT62), .A2(G119), .ZN(n1256) );
NAND4_X1 U928 ( .A1(n1218), .A2(n1069), .A3(n1257), .A4(n1067), .ZN(n1212) );
NOR2_X1 U929 ( .A1(n1085), .A2(n1110), .ZN(n1257) );
XOR2_X1 U930 ( .A(G116), .B(n1258), .Z(G18) );
NOR3_X1 U931 ( .A1(n1259), .A2(n1083), .A3(n1078), .ZN(n1258) );
NAND3_X1 U932 ( .A1(n1260), .A2(n1046), .A3(n1045), .ZN(n1259) );
INV_X1 U933 ( .A(n1077), .ZN(n1045) );
NAND2_X1 U934 ( .A1(n1067), .A2(n1255), .ZN(n1077) );
XOR2_X1 U935 ( .A(KEYINPUT13), .B(n1041), .Z(n1260) );
XNOR2_X1 U936 ( .A(G113), .B(n1211), .ZN(G15) );
NAND3_X1 U937 ( .A1(n1220), .A2(n1219), .A3(n1218), .ZN(n1211) );
AND2_X1 U938 ( .A1(n1217), .A2(n1061), .ZN(n1218) );
INV_X1 U939 ( .A(n1078), .ZN(n1061) );
NAND2_X1 U940 ( .A1(n1072), .A2(n1099), .ZN(n1078) );
INV_X1 U941 ( .A(n1083), .ZN(n1219) );
NAND2_X1 U942 ( .A1(n1110), .A2(n1238), .ZN(n1083) );
INV_X1 U943 ( .A(n1063), .ZN(n1220) );
NAND2_X1 U944 ( .A1(n1069), .A2(n1097), .ZN(n1063) );
INV_X1 U945 ( .A(n1255), .ZN(n1069) );
XOR2_X1 U946 ( .A(n1261), .B(n1210), .Z(G12) );
NAND4_X1 U947 ( .A1(n1217), .A2(n1065), .A3(n1085), .A4(n1086), .ZN(n1210) );
INV_X1 U948 ( .A(n1110), .ZN(n1086) );
XNOR2_X1 U949 ( .A(n1262), .B(n1146), .ZN(n1110) );
NAND2_X1 U950 ( .A1(G217), .A2(n1263), .ZN(n1146) );
NAND2_X1 U951 ( .A1(n1264), .A2(n1145), .ZN(n1262) );
NAND3_X1 U952 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1145) );
NAND2_X1 U953 ( .A1(KEYINPUT21), .A2(n1268), .ZN(n1267) );
OR3_X1 U954 ( .A1(n1268), .A2(KEYINPUT21), .A3(n1269), .ZN(n1266) );
NAND2_X1 U955 ( .A1(n1269), .A2(n1270), .ZN(n1265) );
NAND2_X1 U956 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
INV_X1 U957 ( .A(KEYINPUT21), .ZN(n1272) );
XNOR2_X1 U958 ( .A(KEYINPUT0), .B(n1268), .ZN(n1271) );
XOR2_X1 U959 ( .A(n1273), .B(n1274), .Z(n1268) );
XOR2_X1 U960 ( .A(n1275), .B(n1276), .Z(n1274) );
NAND2_X1 U961 ( .A1(KEYINPUT5), .A2(n1277), .ZN(n1276) );
INV_X1 U962 ( .A(G140), .ZN(n1277) );
NAND2_X1 U963 ( .A1(n1278), .A2(n1279), .ZN(n1275) );
NAND2_X1 U964 ( .A1(n1280), .A2(n1261), .ZN(n1279) );
XOR2_X1 U965 ( .A(KEYINPUT18), .B(n1281), .Z(n1278) );
NOR2_X1 U966 ( .A1(n1261), .A2(n1280), .ZN(n1281) );
XNOR2_X1 U967 ( .A(n1282), .B(n1283), .ZN(n1280) );
XOR2_X1 U968 ( .A(n1284), .B(KEYINPUT43), .Z(n1282) );
INV_X1 U969 ( .A(G119), .ZN(n1284) );
XOR2_X1 U970 ( .A(G146), .B(n1188), .Z(n1273) );
XNOR2_X1 U971 ( .A(G137), .B(n1285), .ZN(n1269) );
NOR3_X1 U972 ( .A1(n1286), .A2(KEYINPUT51), .A3(n1287), .ZN(n1285) );
INV_X1 U973 ( .A(G221), .ZN(n1287) );
INV_X1 U974 ( .A(n1238), .ZN(n1085) );
NAND2_X1 U975 ( .A1(n1288), .A2(n1289), .ZN(n1238) );
NAND2_X1 U976 ( .A1(G472), .A2(n1111), .ZN(n1289) );
XOR2_X1 U977 ( .A(KEYINPUT55), .B(n1290), .Z(n1288) );
NOR2_X1 U978 ( .A1(G472), .A2(n1111), .ZN(n1290) );
NAND2_X1 U979 ( .A1(n1291), .A2(n1264), .ZN(n1111) );
XOR2_X1 U980 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U981 ( .A(n1294), .B(n1166), .Z(n1293) );
XOR2_X1 U982 ( .A(n1295), .B(n1296), .Z(n1166) );
XOR2_X1 U983 ( .A(n1189), .B(n1297), .Z(n1295) );
AND2_X1 U984 ( .A1(G210), .A2(n1298), .ZN(n1297) );
NAND2_X1 U985 ( .A1(KEYINPUT33), .A2(n1299), .ZN(n1294) );
INV_X1 U986 ( .A(G101), .ZN(n1299) );
XNOR2_X1 U987 ( .A(n1300), .B(KEYINPUT32), .ZN(n1292) );
NAND2_X1 U988 ( .A1(KEYINPUT39), .A2(n1167), .ZN(n1300) );
XNOR2_X1 U989 ( .A(n1301), .B(n1302), .ZN(n1167) );
XOR2_X1 U990 ( .A(G119), .B(G116), .Z(n1302) );
NAND2_X1 U991 ( .A1(KEYINPUT30), .A2(G113), .ZN(n1301) );
NOR3_X1 U992 ( .A1(n1097), .A2(n1206), .A3(n1255), .ZN(n1065) );
NAND2_X1 U993 ( .A1(n1303), .A2(n1304), .ZN(n1255) );
NAND2_X1 U994 ( .A1(G478), .A2(n1101), .ZN(n1304) );
XOR2_X1 U995 ( .A(KEYINPUT22), .B(n1096), .Z(n1303) );
NOR2_X1 U996 ( .A1(n1101), .A2(G478), .ZN(n1096) );
OR2_X1 U997 ( .A1(n1149), .A2(G902), .ZN(n1101) );
XNOR2_X1 U998 ( .A(n1305), .B(n1306), .ZN(n1149) );
XOR2_X1 U999 ( .A(n1307), .B(n1308), .Z(n1306) );
XOR2_X1 U1000 ( .A(G116), .B(G107), .Z(n1308) );
XOR2_X1 U1001 ( .A(G143), .B(G134), .Z(n1307) );
XOR2_X1 U1002 ( .A(n1309), .B(n1310), .Z(n1305) );
XOR2_X1 U1003 ( .A(n1311), .B(n1283), .Z(n1309) );
NAND2_X1 U1004 ( .A1(G217), .A2(n1312), .ZN(n1311) );
INV_X1 U1005 ( .A(n1286), .ZN(n1312) );
NAND2_X1 U1006 ( .A1(G234), .A2(n1115), .ZN(n1286) );
INV_X1 U1007 ( .A(n1044), .ZN(n1206) );
NOR2_X1 U1008 ( .A1(n1072), .A2(n1073), .ZN(n1044) );
INV_X1 U1009 ( .A(n1099), .ZN(n1073) );
NAND2_X1 U1010 ( .A1(G221), .A2(n1263), .ZN(n1099) );
NAND2_X1 U1011 ( .A1(n1313), .A2(G234), .ZN(n1263) );
XOR2_X1 U1012 ( .A(n1264), .B(KEYINPUT12), .Z(n1313) );
XNOR2_X1 U1013 ( .A(n1107), .B(G469), .ZN(n1072) );
AND2_X1 U1014 ( .A1(n1314), .A2(n1264), .ZN(n1107) );
XOR2_X1 U1015 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1016 ( .A(G140), .B(n1317), .Z(n1316) );
NOR2_X1 U1017 ( .A1(G953), .A2(n1116), .ZN(n1317) );
INV_X1 U1018 ( .A(G227), .ZN(n1116) );
XNOR2_X1 U1019 ( .A(n1177), .B(n1171), .ZN(n1315) );
XNOR2_X1 U1020 ( .A(n1261), .B(n1296), .ZN(n1171) );
XNOR2_X1 U1021 ( .A(n1318), .B(n1126), .ZN(n1296) );
XOR2_X1 U1022 ( .A(G134), .B(G137), .Z(n1126) );
XOR2_X1 U1023 ( .A(n1129), .B(KEYINPUT40), .Z(n1318) );
XOR2_X1 U1024 ( .A(n1175), .B(n1125), .Z(n1177) );
XNOR2_X1 U1025 ( .A(n1319), .B(n1283), .ZN(n1125) );
XNOR2_X1 U1026 ( .A(n1320), .B(G101), .ZN(n1175) );
NAND2_X1 U1027 ( .A1(n1321), .A2(KEYINPUT15), .ZN(n1320) );
XOR2_X1 U1028 ( .A(n1157), .B(G107), .Z(n1321) );
INV_X1 U1029 ( .A(n1067), .ZN(n1097) );
XOR2_X1 U1030 ( .A(n1156), .B(n1322), .Z(n1067) );
NOR2_X1 U1031 ( .A1(n1154), .A2(G902), .ZN(n1322) );
AND2_X1 U1032 ( .A1(n1323), .A2(n1324), .ZN(n1154) );
NAND2_X1 U1033 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1034 ( .A(KEYINPUT16), .B(n1327), .Z(n1323) );
NOR2_X1 U1035 ( .A1(n1325), .A2(n1326), .ZN(n1327) );
XOR2_X1 U1036 ( .A(n1328), .B(n1124), .Z(n1326) );
XOR2_X1 U1037 ( .A(G125), .B(G140), .Z(n1124) );
XOR2_X1 U1038 ( .A(n1329), .B(G146), .Z(n1328) );
NAND4_X1 U1039 ( .A1(KEYINPUT6), .A2(n1330), .A3(n1331), .A4(n1332), .ZN(n1329) );
NAND2_X1 U1040 ( .A1(KEYINPUT25), .A2(n1333), .ZN(n1332) );
NAND2_X1 U1041 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
XOR2_X1 U1042 ( .A(KEYINPUT52), .B(n1129), .Z(n1334) );
INV_X1 U1043 ( .A(G131), .ZN(n1129) );
NAND2_X1 U1044 ( .A1(n1336), .A2(n1337), .ZN(n1331) );
INV_X1 U1045 ( .A(KEYINPUT25), .ZN(n1337) );
NAND2_X1 U1046 ( .A1(n1338), .A2(n1339), .ZN(n1336) );
OR2_X1 U1047 ( .A1(G131), .A2(KEYINPUT52), .ZN(n1339) );
NAND3_X1 U1048 ( .A1(G131), .A2(n1335), .A3(KEYINPUT52), .ZN(n1338) );
OR2_X1 U1049 ( .A1(n1335), .A2(G131), .ZN(n1330) );
XOR2_X1 U1050 ( .A(n1340), .B(G143), .Z(n1335) );
NAND2_X1 U1051 ( .A1(n1298), .A2(G214), .ZN(n1340) );
NOR2_X1 U1052 ( .A1(G953), .A2(G237), .ZN(n1298) );
XOR2_X1 U1053 ( .A(n1157), .B(n1341), .Z(n1325) );
NOR2_X1 U1054 ( .A1(KEYINPUT56), .A2(n1342), .ZN(n1341) );
XOR2_X1 U1055 ( .A(G113), .B(n1343), .Z(n1342) );
INV_X1 U1056 ( .A(G104), .ZN(n1157) );
INV_X1 U1057 ( .A(G475), .ZN(n1156) );
AND2_X1 U1058 ( .A1(n1041), .A2(n1046), .ZN(n1217) );
NAND2_X1 U1059 ( .A1(n1092), .A2(n1344), .ZN(n1046) );
NAND4_X1 U1060 ( .A1(G953), .A2(G902), .A3(n1254), .A4(n1140), .ZN(n1344) );
INV_X1 U1061 ( .A(G898), .ZN(n1140) );
NAND3_X1 U1062 ( .A1(n1254), .A2(n1115), .A3(G952), .ZN(n1092) );
NAND2_X1 U1063 ( .A1(G237), .A2(G234), .ZN(n1254) );
NOR2_X1 U1064 ( .A1(n1345), .A2(n1244), .ZN(n1041) );
XOR2_X1 U1065 ( .A(n1090), .B(KEYINPUT37), .Z(n1244) );
NAND2_X1 U1066 ( .A1(n1346), .A2(n1347), .ZN(n1090) );
XOR2_X1 U1067 ( .A(KEYINPUT54), .B(G214), .Z(n1346) );
INV_X1 U1068 ( .A(n1091), .ZN(n1345) );
XNOR2_X1 U1069 ( .A(n1348), .B(n1108), .ZN(n1091) );
NAND2_X1 U1070 ( .A1(n1349), .A2(n1264), .ZN(n1108) );
XOR2_X1 U1071 ( .A(n1350), .B(n1351), .Z(n1349) );
XNOR2_X1 U1072 ( .A(n1352), .B(n1222), .ZN(n1351) );
XNOR2_X1 U1073 ( .A(n1138), .B(n1353), .ZN(n1222) );
NOR2_X1 U1074 ( .A1(KEYINPUT47), .A2(n1137), .ZN(n1353) );
NAND2_X1 U1075 ( .A1(n1354), .A2(n1355), .ZN(n1137) );
NAND2_X1 U1076 ( .A1(G110), .A2(n1343), .ZN(n1355) );
XOR2_X1 U1077 ( .A(n1356), .B(KEYINPUT9), .Z(n1354) );
NAND2_X1 U1078 ( .A1(n1310), .A2(n1261), .ZN(n1356) );
INV_X1 U1079 ( .A(n1343), .ZN(n1310) );
XNOR2_X1 U1080 ( .A(G122), .B(KEYINPUT60), .ZN(n1343) );
XOR2_X1 U1081 ( .A(n1357), .B(n1358), .Z(n1138) );
XOR2_X1 U1082 ( .A(G104), .B(n1359), .Z(n1358) );
XOR2_X1 U1083 ( .A(G119), .B(G113), .Z(n1359) );
XOR2_X1 U1084 ( .A(n1360), .B(n1361), .Z(n1357) );
NOR2_X1 U1085 ( .A1(G107), .A2(KEYINPUT7), .ZN(n1361) );
XOR2_X1 U1086 ( .A(n1362), .B(G101), .Z(n1360) );
NAND2_X1 U1087 ( .A1(KEYINPUT24), .A2(n1363), .ZN(n1362) );
INV_X1 U1088 ( .A(G116), .ZN(n1363) );
NAND2_X1 U1089 ( .A1(KEYINPUT49), .A2(n1188), .ZN(n1352) );
INV_X1 U1090 ( .A(G125), .ZN(n1188) );
XOR2_X1 U1091 ( .A(n1189), .B(n1223), .Z(n1350) );
NAND2_X1 U1092 ( .A1(G224), .A2(n1115), .ZN(n1223) );
INV_X1 U1093 ( .A(G953), .ZN(n1115) );
NAND3_X1 U1094 ( .A1(n1364), .A2(n1365), .A3(n1366), .ZN(n1189) );
OR2_X1 U1095 ( .A1(n1283), .A2(n1319), .ZN(n1366) );
NAND2_X1 U1096 ( .A1(n1367), .A2(n1368), .ZN(n1365) );
INV_X1 U1097 ( .A(KEYINPUT57), .ZN(n1368) );
NAND2_X1 U1098 ( .A1(n1369), .A2(n1283), .ZN(n1367) );
XNOR2_X1 U1099 ( .A(KEYINPUT4), .B(n1319), .ZN(n1369) );
NAND2_X1 U1100 ( .A1(KEYINPUT57), .A2(n1370), .ZN(n1364) );
NAND2_X1 U1101 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
OR2_X1 U1102 ( .A1(n1319), .A2(KEYINPUT4), .ZN(n1372) );
NAND3_X1 U1103 ( .A1(n1283), .A2(n1319), .A3(KEYINPUT4), .ZN(n1371) );
XNOR2_X1 U1104 ( .A(G143), .B(G146), .ZN(n1319) );
XOR2_X1 U1105 ( .A(G128), .B(KEYINPUT23), .Z(n1283) );
NAND2_X1 U1106 ( .A1(KEYINPUT48), .A2(n1109), .ZN(n1348) );
NAND2_X1 U1107 ( .A1(G210), .A2(n1347), .ZN(n1109) );
NAND2_X1 U1108 ( .A1(n1373), .A2(n1264), .ZN(n1347) );
INV_X1 U1109 ( .A(G902), .ZN(n1264) );
INV_X1 U1110 ( .A(G237), .ZN(n1373) );
INV_X1 U1111 ( .A(G110), .ZN(n1261) );
endmodule


