//Key = 1000000011111001111111001111010110110011010011110000101111111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359;

XOR2_X1 U734 ( .A(n1024), .B(n1025), .Z(G9) );
NOR2_X1 U735 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR3_X1 U736 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
NAND3_X1 U737 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1028) );
NAND2_X1 U738 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U739 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U740 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U741 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND4_X1 U742 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1041) );
NAND3_X1 U743 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1040) );
NAND2_X1 U744 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NAND2_X1 U745 ( .A1(n1042), .A2(n1044), .ZN(n1050) );
NAND2_X1 U746 ( .A1(n1051), .A2(n1045), .ZN(n1046) );
NAND2_X1 U747 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U748 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U749 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
INV_X1 U750 ( .A(KEYINPUT19), .ZN(n1057) );
NAND3_X1 U751 ( .A1(n1058), .A2(n1059), .A3(n1042), .ZN(n1052) );
NAND2_X1 U752 ( .A1(KEYINPUT19), .A2(n1056), .ZN(n1059) );
XOR2_X1 U753 ( .A(KEYINPUT8), .B(n1060), .Z(n1058) );
NAND2_X1 U754 ( .A1(n1044), .A2(n1061), .ZN(n1036) );
NAND2_X1 U755 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND3_X1 U756 ( .A1(n1048), .A2(n1064), .A3(n1042), .ZN(n1063) );
NAND2_X1 U757 ( .A1(n1065), .A2(n1066), .ZN(n1062) );
NAND2_X1 U758 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U759 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XOR2_X1 U760 ( .A(n1055), .B(KEYINPUT26), .Z(n1069) );
NAND2_X1 U761 ( .A1(n1048), .A2(n1071), .ZN(n1067) );
NAND2_X1 U762 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
OR2_X1 U763 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
INV_X1 U764 ( .A(n1076), .ZN(n1034) );
NOR3_X1 U765 ( .A1(n1077), .A2(G953), .A3(G952), .ZN(n1026) );
INV_X1 U766 ( .A(n1031), .ZN(n1077) );
NAND2_X1 U767 ( .A1(n1078), .A2(n1079), .ZN(n1031) );
NOR4_X1 U768 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1049), .ZN(n1079) );
NOR2_X1 U769 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NAND3_X1 U770 ( .A1(n1085), .A2(n1086), .A3(n1074), .ZN(n1080) );
NOR4_X1 U771 ( .A1(n1087), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1078) );
XOR2_X1 U772 ( .A(n1091), .B(KEYINPUT10), .Z(n1090) );
NAND2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(n1091) );
XOR2_X1 U774 ( .A(G475), .B(KEYINPUT39), .Z(n1084) );
AND2_X1 U775 ( .A1(n1092), .A2(G478), .ZN(n1089) );
XNOR2_X1 U776 ( .A(n1093), .B(n1094), .ZN(n1088) );
NOR2_X1 U777 ( .A1(KEYINPUT1), .A2(n1095), .ZN(n1094) );
NAND4_X1 U778 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1087) );
OR2_X1 U779 ( .A1(n1100), .A2(KEYINPUT60), .ZN(n1099) );
NAND3_X1 U780 ( .A1(n1100), .A2(n1101), .A3(KEYINPUT60), .ZN(n1098) );
XOR2_X1 U781 ( .A(n1102), .B(KEYINPUT30), .Z(n1097) );
XOR2_X1 U782 ( .A(n1103), .B(KEYINPUT6), .Z(n1096) );
XOR2_X1 U783 ( .A(n1104), .B(n1105), .Z(G72) );
XOR2_X1 U784 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U785 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XOR2_X1 U786 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U787 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U788 ( .A(n1114), .B(n1115), .Z(n1110) );
XOR2_X1 U789 ( .A(KEYINPUT53), .B(n1116), .Z(n1115) );
NOR2_X1 U790 ( .A1(G900), .A2(n1117), .ZN(n1108) );
NAND2_X1 U791 ( .A1(n1032), .A2(n1029), .ZN(n1106) );
NAND2_X1 U792 ( .A1(G953), .A2(n1118), .ZN(n1104) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1118) );
XOR2_X1 U794 ( .A(n1119), .B(n1120), .Z(G69) );
NOR2_X1 U795 ( .A1(n1121), .A2(n1032), .ZN(n1120) );
AND2_X1 U796 ( .A1(G224), .A2(G898), .ZN(n1121) );
NAND2_X1 U797 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
NAND2_X1 U798 ( .A1(KEYINPUT36), .A2(n1124), .ZN(n1123) );
NAND2_X1 U799 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XOR2_X1 U800 ( .A(n1127), .B(n1128), .Z(n1122) );
AND2_X1 U801 ( .A1(n1032), .A2(n1030), .ZN(n1128) );
NAND3_X1 U802 ( .A1(n1126), .A2(n1129), .A3(n1125), .ZN(n1127) );
INV_X1 U803 ( .A(KEYINPUT36), .ZN(n1129) );
INV_X1 U804 ( .A(n1130), .ZN(n1126) );
NOR2_X1 U805 ( .A1(n1131), .A2(n1132), .ZN(G66) );
XOR2_X1 U806 ( .A(n1133), .B(n1134), .Z(n1132) );
XNOR2_X1 U807 ( .A(KEYINPUT29), .B(n1135), .ZN(n1133) );
NOR2_X1 U808 ( .A1(n1136), .A2(KEYINPUT40), .ZN(n1135) );
NOR2_X1 U809 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U810 ( .A1(n1131), .A2(n1139), .ZN(G63) );
XOR2_X1 U811 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U812 ( .A1(n1142), .A2(G478), .ZN(n1140) );
NOR2_X1 U813 ( .A1(n1131), .A2(n1143), .ZN(G60) );
NOR3_X1 U814 ( .A1(n1083), .A2(n1144), .A3(n1145), .ZN(n1143) );
AND3_X1 U815 ( .A1(n1146), .A2(G475), .A3(n1142), .ZN(n1145) );
NOR2_X1 U816 ( .A1(n1147), .A2(n1146), .ZN(n1144) );
NOR2_X1 U817 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
INV_X1 U818 ( .A(G475), .ZN(n1149) );
NOR2_X1 U819 ( .A1(n1029), .A2(n1030), .ZN(n1148) );
XNOR2_X1 U820 ( .A(G104), .B(n1150), .ZN(G6) );
NOR3_X1 U821 ( .A1(n1131), .A2(n1151), .A3(n1152), .ZN(G57) );
NOR2_X1 U822 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U823 ( .A1(n1155), .A2(n1156), .ZN(n1153) );
NOR2_X1 U824 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
INV_X1 U825 ( .A(KEYINPUT59), .ZN(n1158) );
NOR2_X1 U826 ( .A1(KEYINPUT59), .A2(n1159), .ZN(n1155) );
NOR2_X1 U827 ( .A1(G101), .A2(n1160), .ZN(n1151) );
NOR2_X1 U828 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U829 ( .A1(n1159), .A2(n1163), .ZN(n1162) );
INV_X1 U830 ( .A(KEYINPUT18), .ZN(n1163) );
AND2_X1 U831 ( .A1(n1164), .A2(n1165), .ZN(n1159) );
NAND2_X1 U832 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NAND2_X1 U833 ( .A1(n1168), .A2(n1169), .ZN(n1164) );
NOR2_X1 U834 ( .A1(KEYINPUT18), .A2(n1157), .ZN(n1161) );
AND2_X1 U835 ( .A1(n1170), .A2(n1171), .ZN(n1157) );
NAND2_X1 U836 ( .A1(n1169), .A2(n1167), .ZN(n1171) );
XOR2_X1 U837 ( .A(n1166), .B(KEYINPUT61), .Z(n1169) );
NAND2_X1 U838 ( .A1(n1166), .A2(n1168), .ZN(n1170) );
XOR2_X1 U839 ( .A(n1172), .B(n1173), .Z(n1166) );
XOR2_X1 U840 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND2_X1 U841 ( .A1(KEYINPUT57), .A2(n1176), .ZN(n1175) );
NAND2_X1 U842 ( .A1(n1142), .A2(G472), .ZN(n1174) );
XOR2_X1 U843 ( .A(n1177), .B(n1178), .Z(n1172) );
NOR2_X1 U844 ( .A1(n1131), .A2(n1179), .ZN(G54) );
XOR2_X1 U845 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U846 ( .A(n1182), .B(n1183), .Z(n1180) );
NAND2_X1 U847 ( .A1(n1142), .A2(G469), .ZN(n1182) );
INV_X1 U848 ( .A(n1138), .ZN(n1142) );
NOR2_X1 U849 ( .A1(n1131), .A2(n1184), .ZN(G51) );
XOR2_X1 U850 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U851 ( .A(n1187), .B(G125), .Z(n1185) );
OR2_X1 U852 ( .A1(n1138), .A2(n1095), .ZN(n1187) );
NAND2_X1 U853 ( .A1(G902), .A2(n1188), .ZN(n1138) );
OR2_X1 U854 ( .A1(n1030), .A2(n1029), .ZN(n1188) );
NAND4_X1 U855 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1029) );
AND4_X1 U856 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
OR2_X1 U857 ( .A1(n1197), .A2(n1072), .ZN(n1191) );
NAND3_X1 U858 ( .A1(n1048), .A2(n1198), .A3(n1199), .ZN(n1190) );
NAND2_X1 U859 ( .A1(n1070), .A2(n1200), .ZN(n1189) );
NAND2_X1 U860 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NAND3_X1 U861 ( .A1(n1203), .A2(n1204), .A3(n1056), .ZN(n1202) );
NAND2_X1 U862 ( .A1(KEYINPUT63), .A2(n1205), .ZN(n1204) );
NAND2_X1 U863 ( .A1(n1206), .A2(n1207), .ZN(n1203) );
INV_X1 U864 ( .A(KEYINPUT63), .ZN(n1207) );
NAND2_X1 U865 ( .A1(n1208), .A2(n1055), .ZN(n1206) );
INV_X1 U866 ( .A(n1042), .ZN(n1055) );
NAND3_X1 U867 ( .A1(n1209), .A2(n1210), .A3(n1060), .ZN(n1201) );
OR2_X1 U868 ( .A1(n1199), .A2(KEYINPUT7), .ZN(n1210) );
NAND2_X1 U869 ( .A1(KEYINPUT7), .A2(n1211), .ZN(n1209) );
NAND3_X1 U870 ( .A1(n1212), .A2(n1213), .A3(n1042), .ZN(n1211) );
NAND4_X1 U871 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1030) );
AND4_X1 U872 ( .A1(n1218), .A2(n1150), .A3(n1025), .A4(n1219), .ZN(n1217) );
NAND3_X1 U873 ( .A1(n1044), .A2(n1220), .A3(n1043), .ZN(n1025) );
NAND3_X1 U874 ( .A1(n1044), .A2(n1220), .A3(n1070), .ZN(n1150) );
NAND2_X1 U875 ( .A1(n1221), .A2(n1222), .ZN(n1216) );
NAND2_X1 U876 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XOR2_X1 U877 ( .A(KEYINPUT45), .B(n1056), .Z(n1223) );
NAND4_X1 U878 ( .A1(n1048), .A2(n1198), .A3(n1225), .A4(n1226), .ZN(n1214) );
NAND2_X1 U879 ( .A1(KEYINPUT34), .A2(n1227), .ZN(n1226) );
NAND2_X1 U880 ( .A1(n1228), .A2(n1229), .ZN(n1225) );
INV_X1 U881 ( .A(KEYINPUT34), .ZN(n1229) );
NAND3_X1 U882 ( .A1(n1065), .A2(n1230), .A3(n1231), .ZN(n1228) );
NOR2_X1 U883 ( .A1(n1032), .A2(G952), .ZN(n1131) );
NAND2_X1 U884 ( .A1(n1232), .A2(n1233), .ZN(G48) );
NAND2_X1 U885 ( .A1(G146), .A2(n1196), .ZN(n1233) );
XOR2_X1 U886 ( .A(KEYINPUT0), .B(n1234), .Z(n1232) );
NOR2_X1 U887 ( .A1(G146), .A2(n1196), .ZN(n1234) );
NAND2_X1 U888 ( .A1(n1235), .A2(n1070), .ZN(n1196) );
XOR2_X1 U889 ( .A(G143), .B(n1236), .Z(G45) );
NOR2_X1 U890 ( .A1(n1237), .A2(n1072), .ZN(n1236) );
XOR2_X1 U891 ( .A(n1197), .B(KEYINPUT48), .Z(n1237) );
NAND4_X1 U892 ( .A1(n1208), .A2(n1056), .A3(n1238), .A4(n1239), .ZN(n1197) );
XNOR2_X1 U893 ( .A(G140), .B(n1240), .ZN(G42) );
NAND3_X1 U894 ( .A1(n1241), .A2(n1060), .A3(KEYINPUT41), .ZN(n1240) );
XNOR2_X1 U895 ( .A(G137), .B(n1242), .ZN(G39) );
NAND3_X1 U896 ( .A1(n1199), .A2(n1048), .A3(n1243), .ZN(n1242) );
XOR2_X1 U897 ( .A(n1244), .B(KEYINPUT11), .Z(n1243) );
XNOR2_X1 U898 ( .A(G134), .B(n1195), .ZN(G36) );
NAND3_X1 U899 ( .A1(n1056), .A2(n1043), .A3(n1199), .ZN(n1195) );
XOR2_X1 U900 ( .A(n1245), .B(n1246), .Z(G33) );
NAND2_X1 U901 ( .A1(n1241), .A2(n1056), .ZN(n1246) );
AND2_X1 U902 ( .A1(n1199), .A2(n1070), .ZN(n1241) );
INV_X1 U903 ( .A(n1205), .ZN(n1199) );
NAND2_X1 U904 ( .A1(n1042), .A2(n1208), .ZN(n1205) );
NOR2_X1 U905 ( .A1(n1075), .A2(n1247), .ZN(n1042) );
INV_X1 U906 ( .A(n1074), .ZN(n1247) );
XOR2_X1 U907 ( .A(n1194), .B(n1248), .Z(G30) );
NAND2_X1 U908 ( .A1(KEYINPUT9), .A2(G128), .ZN(n1248) );
NAND2_X1 U909 ( .A1(n1235), .A2(n1043), .ZN(n1194) );
AND3_X1 U910 ( .A1(n1198), .A2(n1230), .A3(n1208), .ZN(n1235) );
NOR2_X1 U911 ( .A1(n1213), .A2(n1249), .ZN(n1208) );
INV_X1 U912 ( .A(n1244), .ZN(n1198) );
XOR2_X1 U913 ( .A(n1154), .B(n1250), .Z(G3) );
NAND2_X1 U914 ( .A1(n1221), .A2(n1056), .ZN(n1250) );
INV_X1 U915 ( .A(n1251), .ZN(n1221) );
XOR2_X1 U916 ( .A(n1252), .B(n1253), .Z(G27) );
XOR2_X1 U917 ( .A(n1254), .B(KEYINPUT56), .Z(n1253) );
NAND2_X1 U918 ( .A1(KEYINPUT35), .A2(n1193), .ZN(n1252) );
NAND4_X1 U919 ( .A1(n1060), .A2(n1070), .A3(n1255), .A4(n1065), .ZN(n1193) );
NOR2_X1 U920 ( .A1(n1249), .A2(n1072), .ZN(n1255) );
INV_X1 U921 ( .A(n1212), .ZN(n1249) );
NAND2_X1 U922 ( .A1(n1256), .A2(n1076), .ZN(n1212) );
NAND4_X1 U923 ( .A1(n1257), .A2(n1258), .A3(n1259), .A4(n1260), .ZN(n1256) );
INV_X1 U924 ( .A(G900), .ZN(n1260) );
XOR2_X1 U925 ( .A(KEYINPUT37), .B(G902), .Z(n1258) );
XOR2_X1 U926 ( .A(n1218), .B(n1261), .Z(G24) );
XNOR2_X1 U927 ( .A(G122), .B(KEYINPUT23), .ZN(n1261) );
NAND4_X1 U928 ( .A1(n1262), .A2(n1044), .A3(n1238), .A4(n1239), .ZN(n1218) );
NOR2_X1 U929 ( .A1(n1263), .A2(n1264), .ZN(n1044) );
XOR2_X1 U930 ( .A(G119), .B(n1265), .Z(G21) );
NOR4_X1 U931 ( .A1(KEYINPUT22), .A2(n1227), .A3(n1244), .A4(n1266), .ZN(n1265) );
NAND2_X1 U932 ( .A1(n1264), .A2(n1263), .ZN(n1244) );
XNOR2_X1 U933 ( .A(n1267), .B(n1215), .ZN(G18) );
NAND3_X1 U934 ( .A1(n1262), .A2(n1043), .A3(n1056), .ZN(n1215) );
AND2_X1 U935 ( .A1(n1268), .A2(n1239), .ZN(n1043) );
NAND2_X1 U936 ( .A1(KEYINPUT25), .A2(n1269), .ZN(n1267) );
NAND3_X1 U937 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(G15) );
NAND2_X1 U938 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U939 ( .A1(KEYINPUT58), .A2(n1275), .ZN(n1274) );
XOR2_X1 U940 ( .A(KEYINPUT33), .B(n1276), .Z(n1275) );
INV_X1 U941 ( .A(n1219), .ZN(n1273) );
NAND3_X1 U942 ( .A1(KEYINPUT58), .A2(n1219), .A3(n1276), .ZN(n1271) );
NAND3_X1 U943 ( .A1(n1070), .A2(n1262), .A3(n1056), .ZN(n1219) );
AND2_X1 U944 ( .A1(n1277), .A2(n1263), .ZN(n1056) );
INV_X1 U945 ( .A(n1227), .ZN(n1262) );
NAND3_X1 U946 ( .A1(n1230), .A2(n1278), .A3(n1065), .ZN(n1227) );
AND2_X1 U947 ( .A1(n1038), .A2(n1045), .ZN(n1065) );
INV_X1 U948 ( .A(n1072), .ZN(n1230) );
AND2_X1 U949 ( .A1(n1279), .A2(n1238), .ZN(n1070) );
OR2_X1 U950 ( .A1(n1276), .A2(KEYINPUT58), .ZN(n1270) );
XOR2_X1 U951 ( .A(G113), .B(KEYINPUT43), .Z(n1276) );
XOR2_X1 U952 ( .A(G110), .B(n1280), .Z(G12) );
NOR3_X1 U953 ( .A1(n1224), .A2(KEYINPUT13), .A3(n1251), .ZN(n1280) );
NAND2_X1 U954 ( .A1(n1048), .A2(n1220), .ZN(n1251) );
NOR3_X1 U955 ( .A1(n1072), .A2(n1231), .A3(n1213), .ZN(n1220) );
INV_X1 U956 ( .A(n1064), .ZN(n1213) );
NOR2_X1 U957 ( .A1(n1038), .A2(n1049), .ZN(n1064) );
INV_X1 U958 ( .A(n1045), .ZN(n1049) );
NAND2_X1 U959 ( .A1(G221), .A2(n1281), .ZN(n1045) );
XNOR2_X1 U960 ( .A(n1103), .B(KEYINPUT54), .ZN(n1038) );
XOR2_X1 U961 ( .A(n1282), .B(G469), .Z(n1103) );
NAND2_X1 U962 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
XOR2_X1 U963 ( .A(n1285), .B(n1286), .Z(n1283) );
XOR2_X1 U964 ( .A(KEYINPUT3), .B(G146), .Z(n1286) );
XOR2_X1 U965 ( .A(n1287), .B(n1183), .Z(n1285) );
XNOR2_X1 U966 ( .A(n1288), .B(n1289), .ZN(n1183) );
XOR2_X1 U967 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U968 ( .A(n1292), .B(n1293), .Z(n1291) );
AND2_X1 U969 ( .A1(n1032), .A2(G227), .ZN(n1293) );
NAND2_X1 U970 ( .A1(KEYINPUT20), .A2(n1294), .ZN(n1292) );
XOR2_X1 U971 ( .A(G104), .B(n1295), .Z(n1294) );
XOR2_X1 U972 ( .A(KEYINPUT42), .B(G107), .Z(n1295) );
XOR2_X1 U973 ( .A(n1177), .B(n1113), .Z(n1288) );
XOR2_X1 U974 ( .A(G143), .B(KEYINPUT50), .Z(n1113) );
XNOR2_X1 U975 ( .A(n1116), .B(n1296), .ZN(n1177) );
NAND2_X1 U976 ( .A1(n1297), .A2(KEYINPUT52), .ZN(n1287) );
XNOR2_X1 U977 ( .A(G140), .B(KEYINPUT62), .ZN(n1297) );
INV_X1 U978 ( .A(n1278), .ZN(n1231) );
NAND2_X1 U979 ( .A1(n1076), .A2(n1298), .ZN(n1278) );
NAND3_X1 U980 ( .A1(G902), .A2(n1259), .A3(n1130), .ZN(n1298) );
NOR2_X1 U981 ( .A1(n1117), .A2(G898), .ZN(n1130) );
INV_X1 U982 ( .A(n1257), .ZN(n1117) );
XOR2_X1 U983 ( .A(n1032), .B(KEYINPUT31), .Z(n1257) );
NAND3_X1 U984 ( .A1(n1259), .A2(n1032), .A3(G952), .ZN(n1076) );
NAND2_X1 U985 ( .A1(G237), .A2(G234), .ZN(n1259) );
NAND2_X1 U986 ( .A1(n1075), .A2(n1074), .ZN(n1072) );
NAND2_X1 U987 ( .A1(G214), .A2(n1299), .ZN(n1074) );
XOR2_X1 U988 ( .A(n1093), .B(n1095), .Z(n1075) );
NAND2_X1 U989 ( .A1(G210), .A2(n1299), .ZN(n1095) );
NAND2_X1 U990 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
XOR2_X1 U991 ( .A(KEYINPUT15), .B(G237), .Z(n1300) );
NAND2_X1 U992 ( .A1(n1302), .A2(n1284), .ZN(n1093) );
XNOR2_X1 U993 ( .A(n1186), .B(n1303), .ZN(n1302) );
XOR2_X1 U994 ( .A(n1304), .B(KEYINPUT44), .Z(n1303) );
NAND2_X1 U995 ( .A1(KEYINPUT46), .A2(n1254), .ZN(n1304) );
XNOR2_X1 U996 ( .A(n1305), .B(n1306), .ZN(n1186) );
XOR2_X1 U997 ( .A(n1125), .B(n1307), .Z(n1305) );
AND2_X1 U998 ( .A1(n1032), .A2(G224), .ZN(n1307) );
XOR2_X1 U999 ( .A(n1308), .B(n1309), .Z(n1125) );
XOR2_X1 U1000 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1001 ( .A(n1290), .B(n1312), .Z(n1308) );
NOR2_X1 U1002 ( .A1(KEYINPUT2), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1003 ( .A(n1314), .B(G119), .Z(n1313) );
NAND2_X1 U1004 ( .A1(KEYINPUT27), .A2(G116), .ZN(n1314) );
XOR2_X1 U1005 ( .A(n1154), .B(n1315), .Z(n1290) );
XOR2_X1 U1006 ( .A(KEYINPUT4), .B(G110), .Z(n1315) );
INV_X1 U1007 ( .A(G101), .ZN(n1154) );
INV_X1 U1008 ( .A(n1266), .ZN(n1048) );
NAND2_X1 U1009 ( .A1(n1279), .A2(n1268), .ZN(n1266) );
INV_X1 U1010 ( .A(n1238), .ZN(n1268) );
XOR2_X1 U1011 ( .A(n1083), .B(G475), .Z(n1238) );
NOR2_X1 U1012 ( .A1(n1146), .A2(G902), .ZN(n1083) );
XOR2_X1 U1013 ( .A(n1316), .B(n1317), .Z(n1146) );
XOR2_X1 U1014 ( .A(n1318), .B(n1112), .Z(n1317) );
NAND2_X1 U1015 ( .A1(KEYINPUT16), .A2(n1319), .ZN(n1318) );
XOR2_X1 U1016 ( .A(G122), .B(n1310), .Z(n1319) );
XOR2_X1 U1017 ( .A(G104), .B(G113), .Z(n1310) );
XOR2_X1 U1018 ( .A(n1320), .B(G131), .Z(n1316) );
NAND2_X1 U1019 ( .A1(KEYINPUT47), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1020 ( .A(n1322), .B(n1323), .Z(n1321) );
NAND2_X1 U1021 ( .A1(KEYINPUT38), .A2(G143), .ZN(n1323) );
NAND3_X1 U1022 ( .A1(n1324), .A2(n1032), .A3(G214), .ZN(n1322) );
XOR2_X1 U1023 ( .A(n1239), .B(KEYINPUT17), .Z(n1279) );
NAND2_X1 U1024 ( .A1(n1325), .A2(n1326), .ZN(n1239) );
NAND2_X1 U1025 ( .A1(G478), .A2(n1092), .ZN(n1326) );
XOR2_X1 U1026 ( .A(KEYINPUT24), .B(n1082), .Z(n1325) );
NOR2_X1 U1027 ( .A1(n1092), .A2(G478), .ZN(n1082) );
NAND2_X1 U1028 ( .A1(n1141), .A2(n1284), .ZN(n1092) );
XNOR2_X1 U1029 ( .A(n1327), .B(n1328), .ZN(n1141) );
XNOR2_X1 U1030 ( .A(n1329), .B(n1311), .ZN(n1328) );
XNOR2_X1 U1031 ( .A(n1024), .B(G122), .ZN(n1311) );
INV_X1 U1032 ( .A(G107), .ZN(n1024) );
NAND2_X1 U1033 ( .A1(KEYINPUT32), .A2(n1330), .ZN(n1329) );
XOR2_X1 U1034 ( .A(G143), .B(n1116), .Z(n1330) );
XOR2_X1 U1035 ( .A(G134), .B(G128), .Z(n1116) );
XOR2_X1 U1036 ( .A(n1331), .B(G116), .Z(n1327) );
NAND2_X1 U1037 ( .A1(G217), .A2(n1332), .ZN(n1331) );
INV_X1 U1038 ( .A(n1060), .ZN(n1224) );
NOR2_X1 U1039 ( .A1(n1263), .A2(n1277), .ZN(n1060) );
INV_X1 U1040 ( .A(n1264), .ZN(n1277) );
NAND2_X1 U1041 ( .A1(n1085), .A2(n1333), .ZN(n1264) );
NAND2_X1 U1042 ( .A1(n1100), .A2(n1101), .ZN(n1333) );
OR2_X1 U1043 ( .A1(n1101), .A2(n1100), .ZN(n1085) );
INV_X1 U1044 ( .A(n1137), .ZN(n1100) );
NAND2_X1 U1045 ( .A1(G217), .A2(n1281), .ZN(n1137) );
NAND2_X1 U1046 ( .A1(G234), .A2(n1301), .ZN(n1281) );
XOR2_X1 U1047 ( .A(G902), .B(KEYINPUT55), .Z(n1301) );
NAND2_X1 U1048 ( .A1(n1134), .A2(n1284), .ZN(n1101) );
XNOR2_X1 U1049 ( .A(n1334), .B(n1335), .ZN(n1134) );
XOR2_X1 U1050 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1051 ( .A(G119), .B(G110), .Z(n1337) );
XOR2_X1 U1052 ( .A(KEYINPUT49), .B(G137), .Z(n1336) );
XOR2_X1 U1053 ( .A(n1112), .B(n1338), .Z(n1334) );
XOR2_X1 U1054 ( .A(n1339), .B(n1340), .Z(n1338) );
NAND2_X1 U1055 ( .A1(KEYINPUT21), .A2(G128), .ZN(n1340) );
NAND2_X1 U1056 ( .A1(G221), .A2(n1332), .ZN(n1339) );
AND2_X1 U1057 ( .A1(G234), .A2(n1032), .ZN(n1332) );
XOR2_X1 U1058 ( .A(n1254), .B(n1181), .Z(n1112) );
XOR2_X1 U1059 ( .A(G140), .B(G146), .Z(n1181) );
INV_X1 U1060 ( .A(G125), .ZN(n1254) );
NAND2_X1 U1061 ( .A1(n1086), .A2(n1102), .ZN(n1263) );
NAND2_X1 U1062 ( .A1(n1341), .A2(n1342), .ZN(n1102) );
XOR2_X1 U1063 ( .A(KEYINPUT12), .B(G472), .Z(n1342) );
INV_X1 U1064 ( .A(n1343), .ZN(n1341) );
NAND2_X1 U1065 ( .A1(n1344), .A2(n1343), .ZN(n1086) );
NAND2_X1 U1066 ( .A1(n1345), .A2(n1284), .ZN(n1343) );
INV_X1 U1067 ( .A(G902), .ZN(n1284) );
XOR2_X1 U1068 ( .A(n1346), .B(n1347), .Z(n1345) );
XNOR2_X1 U1069 ( .A(n1306), .B(n1176), .ZN(n1347) );
XOR2_X1 U1070 ( .A(n1348), .B(G113), .Z(n1176) );
NAND2_X1 U1071 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
OR2_X1 U1072 ( .A1(n1269), .A2(G119), .ZN(n1350) );
XOR2_X1 U1073 ( .A(n1351), .B(KEYINPUT28), .Z(n1349) );
NAND2_X1 U1074 ( .A1(G119), .A2(n1269), .ZN(n1351) );
INV_X1 U1075 ( .A(G116), .ZN(n1269) );
XOR2_X1 U1076 ( .A(G128), .B(n1178), .Z(n1306) );
AND2_X1 U1077 ( .A1(n1352), .A2(n1353), .ZN(n1178) );
NAND2_X1 U1078 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
XOR2_X1 U1079 ( .A(n1356), .B(G146), .Z(n1354) );
OR3_X1 U1080 ( .A1(n1356), .A2(G146), .A3(n1355), .ZN(n1352) );
INV_X1 U1081 ( .A(KEYINPUT51), .ZN(n1355) );
INV_X1 U1082 ( .A(G143), .ZN(n1356) );
XOR2_X1 U1083 ( .A(n1168), .B(n1357), .Z(n1346) );
XOR2_X1 U1084 ( .A(G101), .B(n1358), .Z(n1357) );
NOR2_X1 U1085 ( .A1(KEYINPUT14), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1086 ( .A(G134), .B(n1296), .Z(n1359) );
XNOR2_X1 U1087 ( .A(n1114), .B(KEYINPUT5), .ZN(n1296) );
XOR2_X1 U1088 ( .A(n1245), .B(G137), .Z(n1114) );
INV_X1 U1089 ( .A(G131), .ZN(n1245) );
INV_X1 U1090 ( .A(n1167), .ZN(n1168) );
NAND3_X1 U1091 ( .A1(n1324), .A2(n1032), .A3(G210), .ZN(n1167) );
INV_X1 U1092 ( .A(G953), .ZN(n1032) );
INV_X1 U1093 ( .A(G237), .ZN(n1324) );
XNOR2_X1 U1094 ( .A(G472), .B(KEYINPUT12), .ZN(n1344) );
endmodule


