//Key = 1101110101010000110011000111111010010000110100001100111100101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386;

NAND2_X1 U751 ( .A1(n1053), .A2(n1054), .ZN(G9) );
NAND2_X1 U752 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XOR2_X1 U753 ( .A(KEYINPUT58), .B(n1057), .Z(n1055) );
NAND2_X1 U754 ( .A1(n1058), .A2(n1059), .ZN(n1053) );
XNOR2_X1 U755 ( .A(n1057), .B(KEYINPUT0), .ZN(n1059) );
XNOR2_X1 U756 ( .A(n1060), .B(KEYINPUT48), .ZN(n1057) );
NOR2_X1 U757 ( .A1(n1061), .A2(n1062), .ZN(G75) );
NOR4_X1 U758 ( .A1(G953), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1062) );
NOR2_X1 U759 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U760 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR3_X1 U761 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
NOR2_X1 U762 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U763 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U764 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NOR2_X1 U765 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U766 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NOR2_X1 U767 ( .A1(n1083), .A2(n1084), .ZN(n1077) );
NOR2_X1 U768 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NOR2_X1 U769 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR3_X1 U770 ( .A1(n1080), .A2(n1089), .A3(n1084), .ZN(n1073) );
NOR2_X1 U771 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR4_X1 U772 ( .A1(n1092), .A2(n1084), .A3(n1080), .A4(n1076), .ZN(n1068) );
NOR2_X1 U773 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR2_X1 U774 ( .A1(n1070), .A2(n1095), .ZN(n1093) );
NOR3_X1 U775 ( .A1(n1063), .A2(G953), .A3(G952), .ZN(n1061) );
AND4_X1 U776 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1063) );
NOR4_X1 U777 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1099) );
XOR2_X1 U778 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U779 ( .A(n1106), .B(n1107), .Z(n1102) );
XOR2_X1 U780 ( .A(n1108), .B(KEYINPUT47), .Z(n1107) );
XNOR2_X1 U781 ( .A(G469), .B(n1109), .ZN(n1101) );
NOR3_X1 U782 ( .A1(n1110), .A2(n1071), .A3(n1111), .ZN(n1098) );
INV_X1 U783 ( .A(n1112), .ZN(n1111) );
XOR2_X1 U784 ( .A(KEYINPUT21), .B(n1113), .Z(n1097) );
XOR2_X1 U785 ( .A(KEYINPUT40), .B(n1114), .Z(n1096) );
INV_X1 U786 ( .A(n1087), .ZN(n1114) );
XOR2_X1 U787 ( .A(n1115), .B(n1116), .Z(G72) );
NAND2_X1 U788 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U789 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U790 ( .A1(n1121), .A2(n1122), .ZN(n1115) );
NAND3_X1 U791 ( .A1(n1123), .A2(n1124), .A3(G900), .ZN(n1122) );
NAND2_X1 U792 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U793 ( .A1(n1127), .A2(G953), .ZN(n1125) );
NAND2_X1 U794 ( .A1(n1127), .A2(G227), .ZN(n1123) );
OR2_X1 U795 ( .A1(n1127), .A2(G953), .ZN(n1121) );
XOR2_X1 U796 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U797 ( .A1(KEYINPUT31), .A2(G125), .ZN(n1129) );
XOR2_X1 U798 ( .A(n1130), .B(n1131), .Z(n1128) );
NOR2_X1 U799 ( .A1(KEYINPUT19), .A2(n1132), .ZN(n1131) );
XOR2_X1 U800 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U801 ( .A(KEYINPUT53), .B(KEYINPUT34), .Z(n1134) );
NAND2_X1 U802 ( .A1(n1135), .A2(n1136), .ZN(G69) );
NAND2_X1 U803 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U804 ( .A1(G953), .A2(n1139), .ZN(n1138) );
NAND3_X1 U805 ( .A1(G953), .A2(n1140), .A3(n1141), .ZN(n1135) );
XNOR2_X1 U806 ( .A(n1137), .B(KEYINPUT8), .ZN(n1141) );
XNOR2_X1 U807 ( .A(n1142), .B(n1143), .ZN(n1137) );
NOR2_X1 U808 ( .A1(G953), .A2(n1144), .ZN(n1143) );
AND2_X1 U809 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U810 ( .A1(n1147), .A2(n1148), .ZN(n1142) );
NAND2_X1 U811 ( .A1(G953), .A2(n1149), .ZN(n1148) );
XOR2_X1 U812 ( .A(n1150), .B(n1151), .Z(n1147) );
XOR2_X1 U813 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U814 ( .A1(KEYINPUT1), .A2(n1154), .ZN(n1152) );
XOR2_X1 U815 ( .A(KEYINPUT61), .B(n1155), .Z(n1154) );
NAND2_X1 U816 ( .A1(G898), .A2(G224), .ZN(n1140) );
NOR2_X1 U817 ( .A1(n1156), .A2(n1157), .ZN(G66) );
XNOR2_X1 U818 ( .A(n1158), .B(n1159), .ZN(n1157) );
NOR2_X1 U819 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR2_X1 U820 ( .A1(n1156), .A2(n1162), .ZN(G63) );
NOR3_X1 U821 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1162) );
NOR3_X1 U822 ( .A1(n1166), .A2(n1108), .A3(n1161), .ZN(n1165) );
NOR2_X1 U823 ( .A1(n1167), .A2(n1168), .ZN(n1164) );
AND2_X1 U824 ( .A1(n1065), .A2(G478), .ZN(n1167) );
NOR2_X1 U825 ( .A1(n1156), .A2(n1169), .ZN(G60) );
XNOR2_X1 U826 ( .A(n1170), .B(n1171), .ZN(n1169) );
AND2_X1 U827 ( .A1(G475), .A2(n1172), .ZN(n1171) );
XNOR2_X1 U828 ( .A(n1145), .B(n1173), .ZN(G6) );
NOR2_X1 U829 ( .A1(KEYINPUT50), .A2(n1174), .ZN(n1173) );
NOR2_X1 U830 ( .A1(n1156), .A2(n1175), .ZN(G57) );
XOR2_X1 U831 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U832 ( .A1(n1178), .A2(n1179), .ZN(n1176) );
NOR2_X1 U833 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NOR2_X1 U834 ( .A1(n1182), .A2(n1183), .ZN(n1180) );
INV_X1 U835 ( .A(KEYINPUT60), .ZN(n1183) );
NOR2_X1 U836 ( .A1(KEYINPUT45), .A2(n1184), .ZN(n1182) );
INV_X1 U837 ( .A(n1185), .ZN(n1184) );
NOR2_X1 U838 ( .A1(n1186), .A2(n1185), .ZN(n1178) );
XOR2_X1 U839 ( .A(n1187), .B(n1188), .Z(n1185) );
XOR2_X1 U840 ( .A(n1189), .B(n1190), .Z(n1187) );
NOR2_X1 U841 ( .A1(n1191), .A2(KEYINPUT45), .ZN(n1186) );
AND2_X1 U842 ( .A1(n1181), .A2(KEYINPUT60), .ZN(n1191) );
NAND2_X1 U843 ( .A1(n1172), .A2(G472), .ZN(n1181) );
NOR3_X1 U844 ( .A1(n1192), .A2(n1156), .A3(n1193), .ZN(G54) );
NOR3_X1 U845 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1193) );
XOR2_X1 U846 ( .A(n1197), .B(n1198), .Z(n1194) );
NOR2_X1 U847 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
INV_X1 U848 ( .A(KEYINPUT35), .ZN(n1200) );
NOR2_X1 U849 ( .A1(n1201), .A2(n1202), .ZN(n1192) );
XOR2_X1 U850 ( .A(n1197), .B(n1203), .Z(n1202) );
AND2_X1 U851 ( .A1(n1199), .A2(KEYINPUT35), .ZN(n1203) );
AND2_X1 U852 ( .A1(n1172), .A2(G469), .ZN(n1197) );
INV_X1 U853 ( .A(n1161), .ZN(n1172) );
NOR2_X1 U854 ( .A1(n1195), .A2(n1196), .ZN(n1201) );
INV_X1 U855 ( .A(KEYINPUT27), .ZN(n1196) );
XOR2_X1 U856 ( .A(n1204), .B(n1205), .Z(n1195) );
XOR2_X1 U857 ( .A(KEYINPUT49), .B(G110), .Z(n1205) );
XOR2_X1 U858 ( .A(n1206), .B(n1207), .Z(n1204) );
NOR2_X1 U859 ( .A1(n1156), .A2(n1208), .ZN(G51) );
XOR2_X1 U860 ( .A(n1209), .B(n1210), .Z(n1208) );
XOR2_X1 U861 ( .A(n1211), .B(n1212), .Z(n1210) );
NAND2_X1 U862 ( .A1(n1213), .A2(KEYINPUT3), .ZN(n1211) );
XNOR2_X1 U863 ( .A(n1214), .B(KEYINPUT5), .ZN(n1213) );
XOR2_X1 U864 ( .A(n1215), .B(n1216), .Z(n1209) );
NOR2_X1 U865 ( .A1(n1105), .A2(n1161), .ZN(n1216) );
NAND2_X1 U866 ( .A1(G902), .A2(n1065), .ZN(n1161) );
NAND4_X1 U867 ( .A1(n1217), .A2(n1119), .A3(n1146), .A4(n1218), .ZN(n1065) );
XNOR2_X1 U868 ( .A(KEYINPUT26), .B(n1120), .ZN(n1218) );
NAND3_X1 U869 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1120) );
XOR2_X1 U870 ( .A(n1222), .B(KEYINPUT6), .Z(n1221) );
AND4_X1 U871 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1146) );
NOR3_X1 U872 ( .A1(n1227), .A2(n1058), .A3(n1228), .ZN(n1226) );
INV_X1 U873 ( .A(n1229), .ZN(n1228) );
INV_X1 U874 ( .A(n1056), .ZN(n1058) );
NAND3_X1 U875 ( .A1(n1090), .A2(n1230), .A3(n1231), .ZN(n1056) );
NAND2_X1 U876 ( .A1(n1082), .A2(n1232), .ZN(n1225) );
NAND2_X1 U877 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND2_X1 U878 ( .A1(n1235), .A2(n1091), .ZN(n1234) );
NAND2_X1 U879 ( .A1(n1236), .A2(n1231), .ZN(n1233) );
NAND4_X1 U880 ( .A1(n1237), .A2(n1094), .A3(n1238), .A4(n1239), .ZN(n1223) );
XOR2_X1 U881 ( .A(KEYINPUT22), .B(n1240), .Z(n1238) );
INV_X1 U882 ( .A(n1241), .ZN(n1237) );
AND4_X1 U883 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1119) );
NOR4_X1 U884 ( .A1(n1246), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1245) );
NAND3_X1 U885 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1244) );
XOR2_X1 U886 ( .A(n1076), .B(KEYINPUT25), .Z(n1252) );
XOR2_X1 U887 ( .A(n1145), .B(KEYINPUT24), .Z(n1217) );
NAND3_X1 U888 ( .A1(n1231), .A2(n1230), .A3(n1091), .ZN(n1145) );
NOR2_X1 U889 ( .A1(n1117), .A2(G952), .ZN(n1156) );
XOR2_X1 U890 ( .A(n1253), .B(n1242), .Z(G48) );
NAND4_X1 U891 ( .A1(n1251), .A2(n1091), .A3(n1254), .A4(n1086), .ZN(n1242) );
XNOR2_X1 U892 ( .A(G143), .B(n1255), .ZN(G45) );
NAND2_X1 U893 ( .A1(KEYINPUT30), .A2(n1249), .ZN(n1255) );
AND3_X1 U894 ( .A1(n1082), .A2(n1254), .A3(n1256), .ZN(n1249) );
NOR3_X1 U895 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1256) );
XOR2_X1 U896 ( .A(n1248), .B(n1260), .Z(G42) );
NOR2_X1 U897 ( .A1(KEYINPUT10), .A2(n1130), .ZN(n1260) );
AND3_X1 U898 ( .A1(n1091), .A2(n1081), .A3(n1250), .ZN(n1248) );
XOR2_X1 U899 ( .A(G137), .B(n1261), .Z(G39) );
NOR2_X1 U900 ( .A1(n1262), .A2(n1241), .ZN(n1261) );
XNOR2_X1 U901 ( .A(G134), .B(n1263), .ZN(G36) );
NAND3_X1 U902 ( .A1(n1219), .A2(n1250), .A3(KEYINPUT7), .ZN(n1263) );
XNOR2_X1 U903 ( .A(G131), .B(n1243), .ZN(G33) );
NAND3_X1 U904 ( .A1(n1250), .A2(n1091), .A3(n1082), .ZN(n1243) );
INV_X1 U905 ( .A(n1262), .ZN(n1250) );
NAND2_X1 U906 ( .A1(n1220), .A2(n1222), .ZN(n1262) );
NOR3_X1 U907 ( .A1(n1070), .A2(n1071), .A3(n1257), .ZN(n1220) );
INV_X1 U908 ( .A(n1095), .ZN(n1071) );
XOR2_X1 U909 ( .A(G128), .B(n1247), .Z(G30) );
AND4_X1 U910 ( .A1(n1251), .A2(n1254), .A3(n1090), .A4(n1264), .ZN(n1247) );
XOR2_X1 U911 ( .A(n1265), .B(n1266), .Z(G3) );
NAND2_X1 U912 ( .A1(KEYINPUT9), .A2(G101), .ZN(n1266) );
NAND4_X1 U913 ( .A1(n1264), .A2(n1239), .A3(n1267), .A4(n1268), .ZN(n1265) );
NOR2_X1 U914 ( .A1(n1269), .A2(n1076), .ZN(n1268) );
XOR2_X1 U915 ( .A(KEYINPUT42), .B(n1094), .Z(n1267) );
XNOR2_X1 U916 ( .A(n1246), .B(n1270), .ZN(G27) );
NAND2_X1 U917 ( .A1(KEYINPUT20), .A2(G125), .ZN(n1270) );
AND4_X1 U918 ( .A1(n1091), .A2(n1254), .A3(n1081), .A4(n1240), .ZN(n1246) );
AND2_X1 U919 ( .A1(n1094), .A2(n1222), .ZN(n1254) );
NAND2_X1 U920 ( .A1(n1067), .A2(n1271), .ZN(n1222) );
NAND4_X1 U921 ( .A1(G953), .A2(G902), .A3(n1272), .A4(n1273), .ZN(n1271) );
INV_X1 U922 ( .A(G900), .ZN(n1273) );
XOR2_X1 U923 ( .A(n1274), .B(G122), .Z(G24) );
NAND2_X1 U924 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
OR2_X1 U925 ( .A1(n1224), .A2(KEYINPUT46), .ZN(n1276) );
NAND2_X1 U926 ( .A1(n1277), .A2(n1235), .ZN(n1224) );
NAND4_X1 U927 ( .A1(n1278), .A2(n1277), .A3(n1279), .A4(KEYINPUT46), .ZN(n1275) );
NOR2_X1 U928 ( .A1(n1280), .A2(n1080), .ZN(n1279) );
NOR3_X1 U929 ( .A1(n1259), .A2(n1258), .A3(n1084), .ZN(n1277) );
INV_X1 U930 ( .A(n1230), .ZN(n1084) );
NOR2_X1 U931 ( .A1(n1281), .A2(n1100), .ZN(n1230) );
INV_X1 U932 ( .A(n1239), .ZN(n1278) );
XOR2_X1 U933 ( .A(G119), .B(n1282), .Z(G21) );
NOR2_X1 U934 ( .A1(n1283), .A2(n1241), .ZN(n1282) );
NAND2_X1 U935 ( .A1(n1236), .A2(n1251), .ZN(n1241) );
AND2_X1 U936 ( .A1(n1100), .A2(n1281), .ZN(n1251) );
XOR2_X1 U937 ( .A(G116), .B(n1227), .Z(G18) );
AND2_X1 U938 ( .A1(n1235), .A2(n1219), .ZN(n1227) );
AND2_X1 U939 ( .A1(n1082), .A2(n1090), .ZN(n1219) );
NOR2_X1 U940 ( .A1(n1113), .A2(n1258), .ZN(n1090) );
INV_X1 U941 ( .A(n1269), .ZN(n1082) );
INV_X1 U942 ( .A(n1283), .ZN(n1235) );
XOR2_X1 U943 ( .A(G113), .B(n1284), .Z(G15) );
NOR3_X1 U944 ( .A1(n1283), .A2(n1285), .A3(n1269), .ZN(n1284) );
NAND2_X1 U945 ( .A1(n1286), .A2(n1100), .ZN(n1269) );
XOR2_X1 U946 ( .A(n1281), .B(KEYINPUT4), .Z(n1286) );
XNOR2_X1 U947 ( .A(n1091), .B(KEYINPUT12), .ZN(n1285) );
AND2_X1 U948 ( .A1(n1258), .A2(n1113), .ZN(n1091) );
INV_X1 U949 ( .A(n1259), .ZN(n1113) );
NAND3_X1 U950 ( .A1(n1094), .A2(n1239), .A3(n1240), .ZN(n1283) );
INV_X1 U951 ( .A(n1080), .ZN(n1240) );
NAND2_X1 U952 ( .A1(n1287), .A2(n1087), .ZN(n1080) );
XOR2_X1 U953 ( .A(n1288), .B(n1229), .Z(G12) );
NAND3_X1 U954 ( .A1(n1081), .A2(n1231), .A3(n1236), .ZN(n1229) );
INV_X1 U955 ( .A(n1076), .ZN(n1236) );
NAND2_X1 U956 ( .A1(n1258), .A2(n1259), .ZN(n1076) );
XOR2_X1 U957 ( .A(n1289), .B(G475), .Z(n1259) );
NAND2_X1 U958 ( .A1(n1170), .A2(n1290), .ZN(n1289) );
XNOR2_X1 U959 ( .A(n1291), .B(n1292), .ZN(n1170) );
NOR2_X1 U960 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
AND3_X1 U961 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1294) );
XOR2_X1 U962 ( .A(n1298), .B(KEYINPUT28), .Z(n1297) );
NOR2_X1 U963 ( .A1(n1295), .A2(n1299), .ZN(n1293) );
NOR2_X1 U964 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
AND2_X1 U965 ( .A1(n1302), .A2(KEYINPUT28), .ZN(n1301) );
NOR2_X1 U966 ( .A1(KEYINPUT28), .A2(n1298), .ZN(n1300) );
INV_X1 U967 ( .A(n1303), .ZN(n1298) );
XNOR2_X1 U968 ( .A(n1304), .B(n1305), .ZN(n1295) );
XOR2_X1 U969 ( .A(G143), .B(G131), .Z(n1305) );
NAND2_X1 U970 ( .A1(n1306), .A2(G214), .ZN(n1304) );
NAND2_X1 U971 ( .A1(n1307), .A2(n1308), .ZN(n1291) );
NAND2_X1 U972 ( .A1(n1309), .A2(n1174), .ZN(n1308) );
XOR2_X1 U973 ( .A(n1310), .B(KEYINPUT18), .Z(n1307) );
OR2_X1 U974 ( .A1(n1309), .A2(n1174), .ZN(n1310) );
INV_X1 U975 ( .A(G104), .ZN(n1174) );
XOR2_X1 U976 ( .A(G122), .B(n1311), .Z(n1309) );
AND2_X1 U977 ( .A1(n1312), .A2(n1313), .ZN(n1258) );
NAND2_X1 U978 ( .A1(G478), .A2(n1106), .ZN(n1313) );
XOR2_X1 U979 ( .A(n1314), .B(KEYINPUT38), .Z(n1312) );
NAND2_X1 U980 ( .A1(n1163), .A2(n1108), .ZN(n1314) );
INV_X1 U981 ( .A(G478), .ZN(n1108) );
INV_X1 U982 ( .A(n1106), .ZN(n1163) );
NAND2_X1 U983 ( .A1(n1166), .A2(n1290), .ZN(n1106) );
INV_X1 U984 ( .A(n1168), .ZN(n1166) );
XOR2_X1 U985 ( .A(n1315), .B(n1316), .Z(n1168) );
AND2_X1 U986 ( .A1(n1317), .A2(G217), .ZN(n1316) );
NAND2_X1 U987 ( .A1(KEYINPUT52), .A2(n1318), .ZN(n1315) );
XOR2_X1 U988 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U989 ( .A(n1321), .B(n1322), .ZN(n1320) );
NAND2_X1 U990 ( .A1(KEYINPUT62), .A2(n1060), .ZN(n1322) );
NAND2_X1 U991 ( .A1(n1323), .A2(KEYINPUT55), .ZN(n1321) );
XNOR2_X1 U992 ( .A(G128), .B(n1324), .ZN(n1323) );
XOR2_X1 U993 ( .A(G143), .B(G134), .Z(n1324) );
XNOR2_X1 U994 ( .A(G116), .B(G122), .ZN(n1319) );
AND3_X1 U995 ( .A1(n1264), .A2(n1239), .A3(n1094), .ZN(n1231) );
INV_X1 U996 ( .A(n1280), .ZN(n1094) );
NAND2_X1 U997 ( .A1(n1070), .A2(n1095), .ZN(n1280) );
NAND2_X1 U998 ( .A1(G214), .A2(n1325), .ZN(n1095) );
XOR2_X1 U999 ( .A(n1104), .B(n1326), .Z(n1070) );
NOR2_X1 U1000 ( .A1(n1327), .A2(KEYINPUT57), .ZN(n1326) );
INV_X1 U1001 ( .A(n1105), .ZN(n1327) );
NAND2_X1 U1002 ( .A1(G210), .A2(n1325), .ZN(n1105) );
NAND2_X1 U1003 ( .A1(n1328), .A2(n1290), .ZN(n1325) );
INV_X1 U1004 ( .A(G237), .ZN(n1328) );
NAND3_X1 U1005 ( .A1(n1329), .A2(n1290), .A3(n1330), .ZN(n1104) );
XOR2_X1 U1006 ( .A(n1331), .B(KEYINPUT23), .Z(n1330) );
NAND2_X1 U1007 ( .A1(n1212), .A2(n1332), .ZN(n1331) );
OR2_X1 U1008 ( .A1(n1332), .A2(n1212), .ZN(n1329) );
XOR2_X1 U1009 ( .A(n1153), .B(n1333), .Z(n1212) );
NOR2_X1 U1010 ( .A1(KEYINPUT39), .A2(n1334), .ZN(n1333) );
XNOR2_X1 U1011 ( .A(n1155), .B(n1150), .ZN(n1334) );
XOR2_X1 U1012 ( .A(n1335), .B(n1336), .Z(n1150) );
NOR2_X1 U1013 ( .A1(G116), .A2(KEYINPUT44), .ZN(n1336) );
XOR2_X1 U1014 ( .A(n1337), .B(n1338), .Z(n1155) );
NOR2_X1 U1015 ( .A1(KEYINPUT13), .A2(n1060), .ZN(n1338) );
INV_X1 U1016 ( .A(G107), .ZN(n1060) );
XOR2_X1 U1017 ( .A(G122), .B(n1288), .Z(n1153) );
XNOR2_X1 U1018 ( .A(n1339), .B(n1214), .ZN(n1332) );
XOR2_X1 U1019 ( .A(G125), .B(n1340), .Z(n1214) );
NAND2_X1 U1020 ( .A1(KEYINPUT43), .A2(n1215), .ZN(n1339) );
NOR2_X1 U1021 ( .A1(n1139), .A2(G953), .ZN(n1215) );
INV_X1 U1022 ( .A(G224), .ZN(n1139) );
NAND2_X1 U1023 ( .A1(n1067), .A2(n1341), .ZN(n1239) );
NAND4_X1 U1024 ( .A1(G953), .A2(G902), .A3(n1272), .A4(n1149), .ZN(n1341) );
INV_X1 U1025 ( .A(G898), .ZN(n1149) );
NAND3_X1 U1026 ( .A1(n1272), .A2(n1117), .A3(G952), .ZN(n1067) );
NAND2_X1 U1027 ( .A1(G237), .A2(G234), .ZN(n1272) );
XOR2_X1 U1028 ( .A(n1086), .B(KEYINPUT36), .Z(n1264) );
INV_X1 U1029 ( .A(n1257), .ZN(n1086) );
NAND2_X1 U1030 ( .A1(n1088), .A2(n1087), .ZN(n1257) );
NAND2_X1 U1031 ( .A1(G221), .A2(n1342), .ZN(n1087) );
INV_X1 U1032 ( .A(n1287), .ZN(n1088) );
XNOR2_X1 U1033 ( .A(n1343), .B(n1109), .ZN(n1287) );
NAND2_X1 U1034 ( .A1(n1344), .A2(n1290), .ZN(n1109) );
XNOR2_X1 U1035 ( .A(n1345), .B(n1199), .ZN(n1344) );
XOR2_X1 U1036 ( .A(n1133), .B(n1346), .Z(n1199) );
XOR2_X1 U1037 ( .A(G107), .B(n1337), .Z(n1346) );
XOR2_X1 U1038 ( .A(G101), .B(G104), .Z(n1337) );
XNOR2_X1 U1039 ( .A(n1347), .B(n1348), .ZN(n1133) );
XOR2_X1 U1040 ( .A(n1349), .B(n1350), .Z(n1348) );
NOR2_X1 U1041 ( .A1(G128), .A2(KEYINPUT37), .ZN(n1349) );
NAND2_X1 U1042 ( .A1(n1351), .A2(n1352), .ZN(n1345) );
NAND2_X1 U1043 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
XOR2_X1 U1044 ( .A(n1288), .B(n1355), .Z(n1354) );
XNOR2_X1 U1045 ( .A(KEYINPUT11), .B(n1206), .ZN(n1353) );
XOR2_X1 U1046 ( .A(n1356), .B(KEYINPUT59), .Z(n1351) );
NAND2_X1 U1047 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
XOR2_X1 U1048 ( .A(G110), .B(n1355), .Z(n1358) );
NOR2_X1 U1049 ( .A1(KEYINPUT15), .A2(n1207), .ZN(n1355) );
XOR2_X1 U1050 ( .A(n1130), .B(KEYINPUT33), .Z(n1207) );
XOR2_X1 U1051 ( .A(KEYINPUT11), .B(n1206), .Z(n1357) );
NOR2_X1 U1052 ( .A1(n1126), .A2(G953), .ZN(n1206) );
INV_X1 U1053 ( .A(G227), .ZN(n1126) );
NAND2_X1 U1054 ( .A1(KEYINPUT17), .A2(G469), .ZN(n1343) );
NOR2_X1 U1055 ( .A1(n1100), .A2(n1359), .ZN(n1081) );
INV_X1 U1056 ( .A(n1281), .ZN(n1359) );
NAND3_X1 U1057 ( .A1(n1360), .A2(n1361), .A3(n1112), .ZN(n1281) );
NAND3_X1 U1058 ( .A1(n1160), .A2(n1290), .A3(n1158), .ZN(n1112) );
NAND2_X1 U1059 ( .A1(n1160), .A2(n1362), .ZN(n1361) );
INV_X1 U1060 ( .A(KEYINPUT54), .ZN(n1362) );
NAND2_X1 U1061 ( .A1(n1110), .A2(KEYINPUT54), .ZN(n1360) );
NOR2_X1 U1062 ( .A1(n1160), .A2(n1363), .ZN(n1110) );
AND2_X1 U1063 ( .A1(n1158), .A2(n1290), .ZN(n1363) );
XNOR2_X1 U1064 ( .A(n1364), .B(n1365), .ZN(n1158) );
XOR2_X1 U1065 ( .A(n1366), .B(n1367), .Z(n1365) );
XOR2_X1 U1066 ( .A(n1302), .B(n1368), .Z(n1367) );
NOR2_X1 U1067 ( .A1(KEYINPUT63), .A2(n1288), .ZN(n1368) );
NAND2_X1 U1068 ( .A1(n1303), .A2(n1296), .ZN(n1302) );
NAND2_X1 U1069 ( .A1(n1369), .A2(n1253), .ZN(n1296) );
INV_X1 U1070 ( .A(G146), .ZN(n1253) );
XOR2_X1 U1071 ( .A(G125), .B(n1130), .Z(n1369) );
INV_X1 U1072 ( .A(G140), .ZN(n1130) );
NAND2_X1 U1073 ( .A1(G146), .A2(n1370), .ZN(n1303) );
XOR2_X1 U1074 ( .A(G140), .B(G125), .Z(n1370) );
NAND2_X1 U1075 ( .A1(n1317), .A2(G221), .ZN(n1366) );
AND2_X1 U1076 ( .A1(G234), .A2(n1117), .ZN(n1317) );
INV_X1 U1077 ( .A(G953), .ZN(n1117) );
XOR2_X1 U1078 ( .A(n1371), .B(n1372), .Z(n1364) );
XOR2_X1 U1079 ( .A(KEYINPUT2), .B(G137), .Z(n1372) );
XNOR2_X1 U1080 ( .A(G119), .B(G128), .ZN(n1371) );
NAND2_X1 U1081 ( .A1(G217), .A2(n1342), .ZN(n1160) );
NAND2_X1 U1082 ( .A1(n1373), .A2(G234), .ZN(n1342) );
XOR2_X1 U1083 ( .A(n1290), .B(KEYINPUT56), .Z(n1373) );
INV_X1 U1084 ( .A(G902), .ZN(n1290) );
XNOR2_X1 U1085 ( .A(n1374), .B(G472), .ZN(n1100) );
NAND2_X1 U1086 ( .A1(n1375), .A2(n1376), .ZN(n1374) );
XOR2_X1 U1087 ( .A(n1377), .B(n1378), .Z(n1376) );
XNOR2_X1 U1088 ( .A(n1188), .B(n1177), .ZN(n1378) );
XNOR2_X1 U1089 ( .A(n1379), .B(G101), .ZN(n1177) );
NAND2_X1 U1090 ( .A1(n1306), .A2(G210), .ZN(n1379) );
NOR2_X1 U1091 ( .A1(G953), .A2(G237), .ZN(n1306) );
XNOR2_X1 U1092 ( .A(n1335), .B(n1380), .ZN(n1188) );
XOR2_X1 U1093 ( .A(KEYINPUT16), .B(G116), .Z(n1380) );
XNOR2_X1 U1094 ( .A(G119), .B(n1311), .ZN(n1335) );
XOR2_X1 U1095 ( .A(G113), .B(KEYINPUT41), .Z(n1311) );
XOR2_X1 U1096 ( .A(n1381), .B(KEYINPUT14), .Z(n1377) );
NAND2_X1 U1097 ( .A1(n1382), .A2(n1383), .ZN(n1381) );
NAND2_X1 U1098 ( .A1(n1190), .A2(n1340), .ZN(n1383) );
INV_X1 U1099 ( .A(n1189), .ZN(n1340) );
XOR2_X1 U1100 ( .A(n1384), .B(KEYINPUT51), .Z(n1382) );
NAND2_X1 U1101 ( .A1(n1189), .A2(n1385), .ZN(n1384) );
XOR2_X1 U1102 ( .A(KEYINPUT32), .B(n1190), .Z(n1385) );
INV_X1 U1103 ( .A(n1347), .ZN(n1190) );
XNOR2_X1 U1104 ( .A(G131), .B(n1386), .ZN(n1347) );
XOR2_X1 U1105 ( .A(G137), .B(G134), .Z(n1386) );
XNOR2_X1 U1106 ( .A(G128), .B(n1350), .ZN(n1189) );
XOR2_X1 U1107 ( .A(G143), .B(G146), .Z(n1350) );
XOR2_X1 U1108 ( .A(KEYINPUT29), .B(G902), .Z(n1375) );
INV_X1 U1109 ( .A(G110), .ZN(n1288) );
endmodule


