//Key = 1010101101110110010010001001100000101111011000010011110011000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355;

XOR2_X1 U740 ( .A(n1033), .B(n1034), .Z(G9) );
NAND2_X1 U741 ( .A1(KEYINPUT20), .A2(G107), .ZN(n1034) );
NOR2_X1 U742 ( .A1(n1035), .A2(n1036), .ZN(G75) );
XOR2_X1 U743 ( .A(KEYINPUT43), .B(n1037), .Z(n1036) );
NOR2_X1 U744 ( .A1(G952), .A2(n1038), .ZN(n1037) );
NOR4_X1 U745 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1038), .ZN(n1035) );
NAND2_X1 U746 ( .A1(n1042), .A2(n1043), .ZN(n1038) );
NAND4_X1 U747 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
NOR2_X1 U748 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XOR2_X1 U749 ( .A(n1050), .B(KEYINPUT1), .Z(n1048) );
NAND4_X1 U750 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1050) );
XOR2_X1 U751 ( .A(n1055), .B(n1056), .Z(n1052) );
NOR2_X1 U752 ( .A1(G469), .A2(KEYINPUT30), .ZN(n1056) );
XNOR2_X1 U753 ( .A(n1057), .B(n1058), .ZN(n1051) );
NAND2_X1 U754 ( .A1(KEYINPUT47), .A2(n1059), .ZN(n1057) );
XNOR2_X1 U755 ( .A(n1060), .B(n1061), .ZN(n1046) );
NAND2_X1 U756 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NAND2_X1 U757 ( .A1(KEYINPUT19), .A2(n1064), .ZN(n1063) );
OR2_X1 U758 ( .A1(KEYINPUT21), .A2(n1064), .ZN(n1062) );
NAND2_X1 U759 ( .A1(G478), .A2(n1065), .ZN(n1044) );
AND3_X1 U760 ( .A1(n1066), .A2(n1067), .A3(KEYINPUT42), .ZN(n1039) );
NAND2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NAND4_X1 U762 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
NAND2_X1 U763 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U764 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
INV_X1 U765 ( .A(n1078), .ZN(n1074) );
NAND3_X1 U766 ( .A1(n1079), .A2(n1053), .A3(n1077), .ZN(n1068) );
NAND2_X1 U767 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U768 ( .A1(n1072), .A2(n1082), .ZN(n1081) );
NAND2_X1 U769 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND3_X1 U770 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
INV_X1 U771 ( .A(KEYINPUT9), .ZN(n1086) );
NAND2_X1 U772 ( .A1(n1071), .A2(n1088), .ZN(n1083) );
NAND2_X1 U773 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U774 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U775 ( .A(KEYINPUT35), .B(n1093), .Z(n1092) );
NAND2_X1 U776 ( .A1(n1070), .A2(n1085), .ZN(n1080) );
NAND4_X1 U777 ( .A1(n1070), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1085) );
NAND2_X1 U778 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XNOR2_X1 U779 ( .A(KEYINPUT25), .B(n1049), .ZN(n1098) );
INV_X1 U780 ( .A(n1071), .ZN(n1049) );
NAND2_X1 U781 ( .A1(n1072), .A2(n1099), .ZN(n1095) );
NAND2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U783 ( .A1(KEYINPUT9), .A2(n1087), .ZN(n1101) );
INV_X1 U784 ( .A(n1102), .ZN(n1100) );
NAND2_X1 U785 ( .A1(n1103), .A2(n1071), .ZN(n1094) );
NAND2_X1 U786 ( .A1(n1104), .A2(n1105), .ZN(G72) );
NAND2_X1 U787 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U788 ( .A1(n1108), .A2(n1109), .ZN(n1104) );
NAND2_X1 U789 ( .A1(n1110), .A2(n1107), .ZN(n1109) );
NAND2_X1 U790 ( .A1(G953), .A2(n1111), .ZN(n1107) );
INV_X1 U791 ( .A(n1112), .ZN(n1110) );
INV_X1 U792 ( .A(n1106), .ZN(n1108) );
XNOR2_X1 U793 ( .A(n1113), .B(n1114), .ZN(n1106) );
NOR3_X1 U794 ( .A1(n1112), .A2(n1115), .A3(n1116), .ZN(n1114) );
NOR2_X1 U795 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U796 ( .A(KEYINPUT56), .B(n1119), .Z(n1117) );
NOR2_X1 U797 ( .A1(n1120), .A2(n1119), .ZN(n1115) );
XNOR2_X1 U798 ( .A(n1121), .B(n1122), .ZN(n1119) );
NOR2_X1 U799 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U800 ( .A(KEYINPUT31), .B(n1125), .Z(n1124) );
NOR2_X1 U801 ( .A1(G131), .A2(n1126), .ZN(n1125) );
XNOR2_X1 U802 ( .A(n1127), .B(KEYINPUT15), .ZN(n1126) );
NOR2_X1 U803 ( .A1(n1128), .A2(n1127), .ZN(n1123) );
XOR2_X1 U804 ( .A(G134), .B(n1129), .Z(n1127) );
NOR2_X1 U805 ( .A1(KEYINPUT29), .A2(n1130), .ZN(n1129) );
XOR2_X1 U806 ( .A(KEYINPUT55), .B(G137), .Z(n1130) );
NAND2_X1 U807 ( .A1(KEYINPUT39), .A2(n1131), .ZN(n1121) );
INV_X1 U808 ( .A(n1118), .ZN(n1120) );
NAND2_X1 U809 ( .A1(n1132), .A2(n1133), .ZN(n1118) );
NAND2_X1 U810 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U811 ( .A(KEYINPUT53), .B(n1136), .Z(n1132) );
NOR2_X1 U812 ( .A1(n1134), .A2(n1137), .ZN(n1136) );
XOR2_X1 U813 ( .A(KEYINPUT33), .B(n1135), .Z(n1137) );
XNOR2_X1 U814 ( .A(n1138), .B(KEYINPUT17), .ZN(n1135) );
XNOR2_X1 U815 ( .A(KEYINPUT28), .B(G125), .ZN(n1134) );
NAND3_X1 U816 ( .A1(n1139), .A2(n1042), .A3(KEYINPUT27), .ZN(n1113) );
NAND2_X1 U817 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U818 ( .A(n1142), .B(KEYINPUT23), .Z(n1140) );
XOR2_X1 U819 ( .A(n1143), .B(n1144), .Z(G69) );
XOR2_X1 U820 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR3_X1 U821 ( .A1(n1147), .A2(KEYINPUT48), .A3(G953), .ZN(n1146) );
NAND2_X1 U822 ( .A1(n1148), .A2(n1149), .ZN(n1145) );
INV_X1 U823 ( .A(n1150), .ZN(n1149) );
NAND2_X1 U824 ( .A1(G953), .A2(n1151), .ZN(n1143) );
NAND2_X1 U825 ( .A1(G898), .A2(G224), .ZN(n1151) );
NOR2_X1 U826 ( .A1(n1152), .A2(n1153), .ZN(G66) );
XOR2_X1 U827 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U828 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U829 ( .A1(KEYINPUT24), .A2(n1158), .ZN(n1154) );
NOR2_X1 U830 ( .A1(n1152), .A2(n1159), .ZN(G63) );
NOR2_X1 U831 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U832 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U833 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NOR2_X1 U834 ( .A1(n1166), .A2(n1157), .ZN(n1162) );
AND2_X1 U835 ( .A1(n1165), .A2(n1164), .ZN(n1160) );
INV_X1 U836 ( .A(KEYINPUT2), .ZN(n1165) );
NOR2_X1 U837 ( .A1(n1152), .A2(n1167), .ZN(G60) );
NOR3_X1 U838 ( .A1(n1064), .A2(n1168), .A3(n1169), .ZN(n1167) );
NOR3_X1 U839 ( .A1(n1170), .A2(n1061), .A3(n1157), .ZN(n1169) );
INV_X1 U840 ( .A(n1171), .ZN(n1170) );
NOR2_X1 U841 ( .A1(n1172), .A2(n1171), .ZN(n1168) );
AND2_X1 U842 ( .A1(n1041), .A2(G475), .ZN(n1172) );
XNOR2_X1 U843 ( .A(G104), .B(n1173), .ZN(G6) );
NOR2_X1 U844 ( .A1(n1152), .A2(n1174), .ZN(G57) );
XOR2_X1 U845 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U846 ( .A(n1177), .B(n1178), .Z(n1176) );
XNOR2_X1 U847 ( .A(G101), .B(n1179), .ZN(n1178) );
NOR2_X1 U848 ( .A1(KEYINPUT16), .A2(n1180), .ZN(n1177) );
XNOR2_X1 U849 ( .A(n1181), .B(n1182), .ZN(n1175) );
NOR2_X1 U850 ( .A1(n1183), .A2(n1157), .ZN(n1182) );
NOR2_X1 U851 ( .A1(n1152), .A2(n1184), .ZN(G54) );
XOR2_X1 U852 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U853 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U854 ( .A(n1189), .B(n1190), .Z(n1185) );
XOR2_X1 U855 ( .A(KEYINPUT41), .B(n1191), .Z(n1190) );
NOR2_X1 U856 ( .A1(n1157), .A2(n1192), .ZN(n1191) );
NAND2_X1 U857 ( .A1(KEYINPUT11), .A2(n1131), .ZN(n1189) );
NOR2_X1 U858 ( .A1(n1042), .A2(G952), .ZN(n1152) );
NOR2_X1 U859 ( .A1(n1193), .A2(n1194), .ZN(G51) );
XOR2_X1 U860 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U861 ( .A(n1197), .B(n1198), .Z(n1196) );
XNOR2_X1 U862 ( .A(n1199), .B(n1200), .ZN(n1195) );
NOR3_X1 U863 ( .A1(n1157), .A2(n1201), .A3(n1202), .ZN(n1200) );
INV_X1 U864 ( .A(G210), .ZN(n1202) );
NAND2_X1 U865 ( .A1(G902), .A2(n1041), .ZN(n1157) );
NAND3_X1 U866 ( .A1(n1141), .A2(n1142), .A3(n1147), .ZN(n1041) );
AND4_X1 U867 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1147) );
AND4_X1 U868 ( .A1(n1033), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1206) );
NAND3_X1 U869 ( .A1(n1071), .A2(n1210), .A3(n1103), .ZN(n1033) );
AND2_X1 U870 ( .A1(n1211), .A2(n1173), .ZN(n1205) );
NAND3_X1 U871 ( .A1(n1071), .A2(n1210), .A3(n1097), .ZN(n1173) );
NAND4_X1 U872 ( .A1(n1212), .A2(n1078), .A3(n1103), .A4(n1213), .ZN(n1142) );
NOR2_X1 U873 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XNOR2_X1 U874 ( .A(KEYINPUT58), .B(n1216), .ZN(n1215) );
AND4_X1 U875 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1141) );
NOR4_X1 U876 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1220) );
INV_X1 U877 ( .A(n1225), .ZN(n1224) );
NOR2_X1 U878 ( .A1(n1042), .A2(n1226), .ZN(n1193) );
XNOR2_X1 U879 ( .A(KEYINPUT46), .B(n1040), .ZN(n1226) );
INV_X1 U880 ( .A(G952), .ZN(n1040) );
NAND3_X1 U881 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(G48) );
OR2_X1 U882 ( .A1(n1219), .A2(G146), .ZN(n1229) );
NAND2_X1 U883 ( .A1(KEYINPUT44), .A2(n1230), .ZN(n1228) );
NAND2_X1 U884 ( .A1(G146), .A2(n1231), .ZN(n1230) );
XNOR2_X1 U885 ( .A(KEYINPUT52), .B(n1219), .ZN(n1231) );
NAND2_X1 U886 ( .A1(n1232), .A2(n1233), .ZN(n1227) );
INV_X1 U887 ( .A(KEYINPUT44), .ZN(n1233) );
NAND2_X1 U888 ( .A1(n1234), .A2(n1235), .ZN(n1232) );
NAND3_X1 U889 ( .A1(KEYINPUT52), .A2(G146), .A3(n1219), .ZN(n1235) );
OR2_X1 U890 ( .A1(n1219), .A2(KEYINPUT52), .ZN(n1234) );
NAND3_X1 U891 ( .A1(n1097), .A2(n1078), .A3(n1236), .ZN(n1219) );
XOR2_X1 U892 ( .A(n1217), .B(n1237), .Z(G45) );
XNOR2_X1 U893 ( .A(KEYINPUT38), .B(n1238), .ZN(n1237) );
NAND4_X1 U894 ( .A1(n1212), .A2(n1078), .A3(n1102), .A4(n1239), .ZN(n1217) );
NOR3_X1 U895 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1239) );
XNOR2_X1 U896 ( .A(G140), .B(n1218), .ZN(G42) );
NAND3_X1 U897 ( .A1(n1087), .A2(n1097), .A3(n1243), .ZN(n1218) );
XOR2_X1 U898 ( .A(G137), .B(n1223), .Z(G39) );
AND3_X1 U899 ( .A1(n1244), .A2(n1072), .A3(n1243), .ZN(n1223) );
XNOR2_X1 U900 ( .A(n1245), .B(n1222), .ZN(G36) );
AND3_X1 U901 ( .A1(n1102), .A2(n1103), .A3(n1243), .ZN(n1222) );
XNOR2_X1 U902 ( .A(n1128), .B(n1221), .ZN(G33) );
AND3_X1 U903 ( .A1(n1102), .A2(n1097), .A3(n1243), .ZN(n1221) );
NOR4_X1 U904 ( .A1(n1246), .A2(n1089), .A3(n1242), .A4(n1076), .ZN(n1243) );
XNOR2_X1 U905 ( .A(G128), .B(n1247), .ZN(G30) );
NAND2_X1 U906 ( .A1(n1078), .A2(n1248), .ZN(n1247) );
XOR2_X1 U907 ( .A(KEYINPUT22), .B(n1249), .Z(n1248) );
AND2_X1 U908 ( .A1(n1103), .A2(n1236), .ZN(n1249) );
NOR3_X1 U909 ( .A1(n1089), .A2(n1242), .A3(n1214), .ZN(n1236) );
INV_X1 U910 ( .A(n1216), .ZN(n1242) );
INV_X1 U911 ( .A(n1212), .ZN(n1089) );
XNOR2_X1 U912 ( .A(G101), .B(n1211), .ZN(G3) );
NAND3_X1 U913 ( .A1(n1210), .A2(n1072), .A3(n1102), .ZN(n1211) );
XNOR2_X1 U914 ( .A(G125), .B(n1225), .ZN(G27) );
NAND4_X1 U915 ( .A1(n1078), .A2(n1216), .A3(n1097), .A4(n1250), .ZN(n1225) );
NOR2_X1 U916 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U917 ( .A1(n1253), .A2(n1254), .ZN(n1216) );
NAND3_X1 U918 ( .A1(G902), .A2(n1067), .A3(n1112), .ZN(n1254) );
NOR2_X1 U919 ( .A1(G900), .A2(n1042), .ZN(n1112) );
XNOR2_X1 U920 ( .A(G122), .B(n1203), .ZN(G24) );
NAND4_X1 U921 ( .A1(n1255), .A2(n1071), .A3(n1256), .A4(n1257), .ZN(n1203) );
NOR2_X1 U922 ( .A1(n1258), .A2(n1259), .ZN(n1071) );
XNOR2_X1 U923 ( .A(G119), .B(n1260), .ZN(G21) );
NAND2_X1 U924 ( .A1(KEYINPUT0), .A2(n1261), .ZN(n1260) );
INV_X1 U925 ( .A(n1204), .ZN(n1261) );
NAND3_X1 U926 ( .A1(n1244), .A2(n1072), .A3(n1255), .ZN(n1204) );
INV_X1 U927 ( .A(n1214), .ZN(n1244) );
NAND2_X1 U928 ( .A1(n1259), .A2(n1258), .ZN(n1214) );
XNOR2_X1 U929 ( .A(G116), .B(n1209), .ZN(G18) );
NAND3_X1 U930 ( .A1(n1255), .A2(n1103), .A3(n1102), .ZN(n1209) );
NOR2_X1 U931 ( .A1(n1256), .A2(n1241), .ZN(n1103) );
INV_X1 U932 ( .A(n1257), .ZN(n1241) );
NAND2_X1 U933 ( .A1(n1262), .A2(n1263), .ZN(G15) );
NAND2_X1 U934 ( .A1(G113), .A2(n1208), .ZN(n1263) );
XOR2_X1 U935 ( .A(n1264), .B(KEYINPUT40), .Z(n1262) );
OR2_X1 U936 ( .A1(n1208), .A2(G113), .ZN(n1264) );
NAND3_X1 U937 ( .A1(n1255), .A2(n1097), .A3(n1102), .ZN(n1208) );
NOR2_X1 U938 ( .A1(n1259), .A2(n1265), .ZN(n1102) );
AND2_X1 U939 ( .A1(n1070), .A2(n1266), .ZN(n1255) );
INV_X1 U940 ( .A(n1252), .ZN(n1070) );
NAND2_X1 U941 ( .A1(n1093), .A2(n1054), .ZN(n1252) );
XOR2_X1 U942 ( .A(n1267), .B(G110), .Z(G12) );
NAND2_X1 U943 ( .A1(KEYINPUT7), .A2(n1207), .ZN(n1267) );
NAND3_X1 U944 ( .A1(n1210), .A2(n1072), .A3(n1087), .ZN(n1207) );
INV_X1 U945 ( .A(n1251), .ZN(n1087) );
NAND2_X1 U946 ( .A1(n1265), .A2(n1259), .ZN(n1251) );
XOR2_X1 U947 ( .A(n1268), .B(n1156), .Z(n1259) );
NAND2_X1 U948 ( .A1(G217), .A2(n1269), .ZN(n1156) );
NAND2_X1 U949 ( .A1(n1158), .A2(n1270), .ZN(n1268) );
XNOR2_X1 U950 ( .A(n1271), .B(n1272), .ZN(n1158) );
XNOR2_X1 U951 ( .A(G137), .B(n1273), .ZN(n1272) );
NAND3_X1 U952 ( .A1(n1274), .A2(n1042), .A3(G221), .ZN(n1273) );
NAND3_X1 U953 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1271) );
NAND2_X1 U954 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
OR3_X1 U955 ( .A1(n1279), .A2(n1278), .A3(KEYINPUT45), .ZN(n1276) );
XOR2_X1 U956 ( .A(n1280), .B(n1281), .Z(n1278) );
XNOR2_X1 U957 ( .A(G110), .B(G128), .ZN(n1280) );
OR2_X1 U958 ( .A1(KEYINPUT59), .A2(n1282), .ZN(n1279) );
NAND2_X1 U959 ( .A1(KEYINPUT45), .A2(n1282), .ZN(n1275) );
XNOR2_X1 U960 ( .A(G146), .B(n1283), .ZN(n1282) );
INV_X1 U961 ( .A(n1258), .ZN(n1265) );
XOR2_X1 U962 ( .A(n1284), .B(n1183), .Z(n1258) );
INV_X1 U963 ( .A(G472), .ZN(n1183) );
NAND2_X1 U964 ( .A1(n1285), .A2(n1270), .ZN(n1284) );
XOR2_X1 U965 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U966 ( .A(n1288), .B(n1180), .Z(n1287) );
XNOR2_X1 U967 ( .A(n1289), .B(n1281), .ZN(n1180) );
XNOR2_X1 U968 ( .A(n1290), .B(n1291), .ZN(n1288) );
INV_X1 U969 ( .A(n1181), .ZN(n1291) );
XOR2_X1 U970 ( .A(n1198), .B(n1188), .Z(n1181) );
NAND2_X1 U971 ( .A1(KEYINPUT63), .A2(G101), .ZN(n1290) );
XOR2_X1 U972 ( .A(n1179), .B(n1292), .Z(n1286) );
XOR2_X1 U973 ( .A(KEYINPUT4), .B(KEYINPUT18), .Z(n1292) );
NAND2_X1 U974 ( .A1(G210), .A2(n1293), .ZN(n1179) );
NAND2_X1 U975 ( .A1(n1294), .A2(n1295), .ZN(n1072) );
OR3_X1 U976 ( .A1(n1257), .A2(n1256), .A3(KEYINPUT3), .ZN(n1295) );
INV_X1 U977 ( .A(n1240), .ZN(n1256) );
NAND2_X1 U978 ( .A1(KEYINPUT3), .A2(n1097), .ZN(n1294) );
NOR2_X1 U979 ( .A1(n1257), .A2(n1240), .ZN(n1097) );
XOR2_X1 U980 ( .A(n1064), .B(n1061), .Z(n1240) );
INV_X1 U981 ( .A(G475), .ZN(n1061) );
NOR2_X1 U982 ( .A1(n1171), .A2(G902), .ZN(n1064) );
XNOR2_X1 U983 ( .A(n1296), .B(n1297), .ZN(n1171) );
XNOR2_X1 U984 ( .A(n1298), .B(n1299), .ZN(n1297) );
XOR2_X1 U985 ( .A(n1300), .B(n1301), .Z(n1299) );
AND2_X1 U986 ( .A1(n1293), .A2(G214), .ZN(n1301) );
NOR2_X1 U987 ( .A1(G953), .A2(G237), .ZN(n1293) );
NAND3_X1 U988 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1300) );
NAND2_X1 U989 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
OR3_X1 U990 ( .A1(n1306), .A2(n1305), .A3(KEYINPUT54), .ZN(n1303) );
INV_X1 U991 ( .A(n1283), .ZN(n1305) );
XNOR2_X1 U992 ( .A(G140), .B(n1199), .ZN(n1283) );
NAND2_X1 U993 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
XOR2_X1 U994 ( .A(KEYINPUT8), .B(KEYINPUT57), .Z(n1307) );
NAND2_X1 U995 ( .A1(KEYINPUT54), .A2(G146), .ZN(n1302) );
XNOR2_X1 U996 ( .A(G104), .B(n1309), .ZN(n1296) );
XNOR2_X1 U997 ( .A(n1128), .B(G113), .ZN(n1309) );
NAND3_X1 U998 ( .A1(n1310), .A2(n1311), .A3(n1045), .ZN(n1257) );
NAND2_X1 U999 ( .A1(n1312), .A2(n1166), .ZN(n1045) );
INV_X1 U1000 ( .A(G478), .ZN(n1166) );
OR2_X1 U1001 ( .A1(G478), .A2(KEYINPUT50), .ZN(n1311) );
NAND3_X1 U1002 ( .A1(G478), .A2(n1065), .A3(KEYINPUT50), .ZN(n1310) );
INV_X1 U1003 ( .A(n1312), .ZN(n1065) );
NOR2_X1 U1004 ( .A1(n1164), .A2(G902), .ZN(n1312) );
XNOR2_X1 U1005 ( .A(n1313), .B(n1314), .ZN(n1164) );
XOR2_X1 U1006 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1007 ( .A(n1317), .B(G116), .ZN(n1316) );
XNOR2_X1 U1008 ( .A(KEYINPUT10), .B(n1245), .ZN(n1315) );
INV_X1 U1009 ( .A(G134), .ZN(n1245) );
XOR2_X1 U1010 ( .A(n1318), .B(n1298), .Z(n1313) );
XNOR2_X1 U1011 ( .A(G122), .B(n1238), .ZN(n1298) );
XOR2_X1 U1012 ( .A(n1319), .B(G107), .Z(n1318) );
NAND3_X1 U1013 ( .A1(n1274), .A2(n1042), .A3(G217), .ZN(n1319) );
XOR2_X1 U1014 ( .A(G234), .B(KEYINPUT32), .Z(n1274) );
AND2_X1 U1015 ( .A1(n1212), .A2(n1266), .ZN(n1210) );
AND2_X1 U1016 ( .A1(n1078), .A2(n1320), .ZN(n1266) );
NAND2_X1 U1017 ( .A1(n1253), .A2(n1321), .ZN(n1320) );
NAND3_X1 U1018 ( .A1(G902), .A2(n1067), .A3(n1150), .ZN(n1321) );
NOR2_X1 U1019 ( .A1(n1042), .A2(G898), .ZN(n1150) );
NAND3_X1 U1020 ( .A1(n1067), .A2(n1042), .A3(G952), .ZN(n1253) );
NAND2_X1 U1021 ( .A1(G237), .A2(G234), .ZN(n1067) );
NOR2_X1 U1022 ( .A1(n1077), .A2(n1076), .ZN(n1078) );
INV_X1 U1023 ( .A(n1053), .ZN(n1076) );
NAND2_X1 U1024 ( .A1(G214), .A2(n1322), .ZN(n1053) );
INV_X1 U1025 ( .A(n1201), .ZN(n1322) );
INV_X1 U1026 ( .A(n1246), .ZN(n1077) );
XNOR2_X1 U1027 ( .A(n1058), .B(n1059), .ZN(n1246) );
AND2_X1 U1028 ( .A1(n1323), .A2(G210), .ZN(n1059) );
XNOR2_X1 U1029 ( .A(n1201), .B(KEYINPUT49), .ZN(n1323) );
NOR2_X1 U1030 ( .A1(n1324), .A2(G237), .ZN(n1201) );
XNOR2_X1 U1031 ( .A(n1270), .B(KEYINPUT26), .ZN(n1324) );
NAND2_X1 U1032 ( .A1(n1325), .A2(n1326), .ZN(n1058) );
XNOR2_X1 U1033 ( .A(KEYINPUT51), .B(n1270), .ZN(n1326) );
XOR2_X1 U1034 ( .A(n1197), .B(n1327), .Z(n1325) );
XNOR2_X1 U1035 ( .A(n1199), .B(n1328), .ZN(n1327) );
NOR2_X1 U1036 ( .A1(KEYINPUT5), .A2(n1198), .ZN(n1328) );
XNOR2_X1 U1037 ( .A(n1329), .B(n1330), .ZN(n1198) );
XNOR2_X1 U1038 ( .A(n1331), .B(n1238), .ZN(n1329) );
NAND2_X1 U1039 ( .A1(KEYINPUT6), .A2(n1308), .ZN(n1331) );
INV_X1 U1040 ( .A(G125), .ZN(n1199) );
XNOR2_X1 U1041 ( .A(n1332), .B(n1148), .ZN(n1197) );
XNOR2_X1 U1042 ( .A(n1333), .B(n1334), .ZN(n1148) );
XOR2_X1 U1043 ( .A(n1335), .B(n1336), .Z(n1334) );
NAND2_X1 U1044 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
NAND2_X1 U1045 ( .A1(n1289), .A2(n1281), .ZN(n1338) );
INV_X1 U1046 ( .A(n1339), .ZN(n1281) );
NAND2_X1 U1047 ( .A1(n1339), .A2(n1340), .ZN(n1337) );
XNOR2_X1 U1048 ( .A(n1289), .B(KEYINPUT12), .ZN(n1340) );
XOR2_X1 U1049 ( .A(G116), .B(G113), .Z(n1289) );
XOR2_X1 U1050 ( .A(G119), .B(KEYINPUT13), .Z(n1339) );
XOR2_X1 U1051 ( .A(n1341), .B(G122), .Z(n1333) );
NAND2_X1 U1052 ( .A1(KEYINPUT34), .A2(n1342), .ZN(n1341) );
INV_X1 U1053 ( .A(G101), .ZN(n1342) );
NAND2_X1 U1054 ( .A1(G224), .A2(n1042), .ZN(n1332) );
INV_X1 U1055 ( .A(G953), .ZN(n1042) );
NOR2_X1 U1056 ( .A1(n1093), .A2(n1091), .ZN(n1212) );
INV_X1 U1057 ( .A(n1054), .ZN(n1091) );
NAND2_X1 U1058 ( .A1(G221), .A2(n1269), .ZN(n1054) );
NAND2_X1 U1059 ( .A1(G234), .A2(n1270), .ZN(n1269) );
XNOR2_X1 U1060 ( .A(n1343), .B(n1055), .ZN(n1093) );
AND2_X1 U1061 ( .A1(n1344), .A2(n1270), .ZN(n1055) );
INV_X1 U1062 ( .A(G902), .ZN(n1270) );
XOR2_X1 U1063 ( .A(n1187), .B(n1345), .Z(n1344) );
XNOR2_X1 U1064 ( .A(n1346), .B(n1347), .ZN(n1345) );
NAND2_X1 U1065 ( .A1(KEYINPUT37), .A2(n1131), .ZN(n1347) );
XNOR2_X1 U1066 ( .A(n1348), .B(n1330), .ZN(n1131) );
XNOR2_X1 U1067 ( .A(n1317), .B(KEYINPUT61), .ZN(n1330) );
INV_X1 U1068 ( .A(G128), .ZN(n1317) );
XNOR2_X1 U1069 ( .A(n1349), .B(n1308), .ZN(n1348) );
INV_X1 U1070 ( .A(G146), .ZN(n1308) );
NAND2_X1 U1071 ( .A1(KEYINPUT62), .A2(n1238), .ZN(n1349) );
INV_X1 U1072 ( .A(G143), .ZN(n1238) );
NAND2_X1 U1073 ( .A1(KEYINPUT14), .A2(n1188), .ZN(n1346) );
XNOR2_X1 U1074 ( .A(n1128), .B(n1350), .ZN(n1188) );
NOR2_X1 U1075 ( .A1(KEYINPUT60), .A2(n1351), .ZN(n1350) );
XNOR2_X1 U1076 ( .A(G134), .B(G137), .ZN(n1351) );
INV_X1 U1077 ( .A(G131), .ZN(n1128) );
XOR2_X1 U1078 ( .A(n1352), .B(n1353), .Z(n1187) );
XNOR2_X1 U1079 ( .A(n1138), .B(G101), .ZN(n1353) );
INV_X1 U1080 ( .A(G140), .ZN(n1138) );
XOR2_X1 U1081 ( .A(n1335), .B(n1354), .Z(n1352) );
NOR2_X1 U1082 ( .A1(G953), .A2(n1111), .ZN(n1354) );
INV_X1 U1083 ( .A(G227), .ZN(n1111) );
XNOR2_X1 U1084 ( .A(G104), .B(n1355), .ZN(n1335) );
XOR2_X1 U1085 ( .A(G110), .B(G107), .Z(n1355) );
NAND2_X1 U1086 ( .A1(KEYINPUT36), .A2(n1192), .ZN(n1343) );
INV_X1 U1087 ( .A(G469), .ZN(n1192) );
endmodule


