//Key = 1011100111101001110011010010001101001010111001111001100110100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270;

XNOR2_X1 U702 ( .A(n961), .B(n962), .ZN(G9) );
NOR2_X1 U703 ( .A1(n963), .A2(n964), .ZN(G75) );
NOR4_X1 U704 ( .A1(n965), .A2(n966), .A3(n967), .A4(n968), .ZN(n964) );
INV_X1 U705 ( .A(G952), .ZN(n968) );
NOR2_X1 U706 ( .A1(KEYINPUT3), .A2(n969), .ZN(n967) );
NOR3_X1 U707 ( .A1(n970), .A2(n971), .A3(n972), .ZN(n969) );
NAND3_X1 U708 ( .A1(n973), .A2(n974), .A3(n975), .ZN(n970) );
NAND3_X1 U709 ( .A1(n976), .A2(n977), .A3(n978), .ZN(n965) );
NAND2_X1 U710 ( .A1(n979), .A2(n980), .ZN(n978) );
NAND2_X1 U711 ( .A1(n981), .A2(n982), .ZN(n980) );
NAND4_X1 U712 ( .A1(n974), .A2(n983), .A3(n984), .A4(n985), .ZN(n982) );
NAND2_X1 U713 ( .A1(n986), .A2(n987), .ZN(n984) );
NAND2_X1 U714 ( .A1(n988), .A2(n989), .ZN(n987) );
NAND2_X1 U715 ( .A1(n990), .A2(n991), .ZN(n989) );
NAND2_X1 U716 ( .A1(n975), .A2(n992), .ZN(n986) );
NAND2_X1 U717 ( .A1(n993), .A2(n994), .ZN(n992) );
NAND2_X1 U718 ( .A1(n995), .A2(n996), .ZN(n994) );
NAND3_X1 U719 ( .A1(n975), .A2(n997), .A3(n988), .ZN(n981) );
NAND2_X1 U720 ( .A1(n998), .A2(n999), .ZN(n997) );
NAND3_X1 U721 ( .A1(n973), .A2(n974), .A3(KEYINPUT3), .ZN(n999) );
NAND3_X1 U722 ( .A1(n1000), .A2(n1001), .A3(n983), .ZN(n998) );
NAND2_X1 U723 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
OR3_X1 U724 ( .A1(n1004), .A2(n1005), .A3(n1002), .ZN(n1000) );
INV_X1 U725 ( .A(n972), .ZN(n979) );
NOR3_X1 U726 ( .A1(n1006), .A2(G953), .A3(n1007), .ZN(n963) );
INV_X1 U727 ( .A(n976), .ZN(n1007) );
NAND4_X1 U728 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n976) );
NOR4_X1 U729 ( .A1(n996), .A2(n1002), .A3(n1012), .A4(n1013), .ZN(n1011) );
XOR2_X1 U730 ( .A(n1014), .B(KEYINPUT7), .Z(n1013) );
XOR2_X1 U731 ( .A(n1015), .B(n1016), .Z(n1012) );
NAND2_X1 U732 ( .A1(KEYINPUT8), .A2(n1017), .ZN(n1015) );
NOR2_X1 U733 ( .A1(n1018), .A2(n1019), .ZN(n1010) );
XNOR2_X1 U734 ( .A(n1020), .B(G478), .ZN(n1009) );
XNOR2_X1 U735 ( .A(n1021), .B(KEYINPUT34), .ZN(n1008) );
XNOR2_X1 U736 ( .A(G952), .B(KEYINPUT16), .ZN(n1006) );
XOR2_X1 U737 ( .A(n1022), .B(n1023), .Z(G72) );
NOR2_X1 U738 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
XOR2_X1 U739 ( .A(n1026), .B(n1027), .Z(n1025) );
XOR2_X1 U740 ( .A(n1028), .B(n1029), .Z(n1027) );
XOR2_X1 U741 ( .A(n1030), .B(n1031), .Z(n1026) );
XNOR2_X1 U742 ( .A(KEYINPUT35), .B(n1032), .ZN(n1031) );
NAND3_X1 U743 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1022) );
INV_X1 U744 ( .A(n1024), .ZN(n1035) );
NAND2_X1 U745 ( .A1(G953), .A2(n1036), .ZN(n1034) );
NAND2_X1 U746 ( .A1(n1037), .A2(n977), .ZN(n1033) );
NAND3_X1 U747 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
XNOR2_X1 U748 ( .A(n1041), .B(KEYINPUT22), .ZN(n1040) );
XOR2_X1 U749 ( .A(KEYINPUT62), .B(n1042), .Z(n1039) );
NAND2_X1 U750 ( .A1(n1043), .A2(n1044), .ZN(G69) );
NAND3_X1 U751 ( .A1(G953), .A2(n1045), .A3(n1046), .ZN(n1044) );
XOR2_X1 U752 ( .A(n1047), .B(KEYINPUT60), .Z(n1043) );
NAND2_X1 U753 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U754 ( .A1(G953), .A2(n1045), .ZN(n1049) );
NAND2_X1 U755 ( .A1(G224), .A2(G898), .ZN(n1045) );
XOR2_X1 U756 ( .A(n1046), .B(KEYINPUT17), .Z(n1048) );
XOR2_X1 U757 ( .A(n1050), .B(n1051), .Z(n1046) );
NOR2_X1 U758 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XOR2_X1 U759 ( .A(KEYINPUT6), .B(n1054), .Z(n1053) );
NAND2_X1 U760 ( .A1(n977), .A2(n1055), .ZN(n1050) );
NAND2_X1 U761 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U762 ( .A1(n1058), .A2(n1059), .ZN(G66) );
NOR3_X1 U763 ( .A1(n1016), .A2(n1060), .A3(n1061), .ZN(n1059) );
NOR3_X1 U764 ( .A1(n1062), .A2(n1017), .A3(n1063), .ZN(n1061) );
NOR2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1060) );
NOR2_X1 U766 ( .A1(n1066), .A2(n1017), .ZN(n1064) );
NOR2_X1 U767 ( .A1(n1058), .A2(n1067), .ZN(G63) );
NOR3_X1 U768 ( .A1(n1020), .A2(n1068), .A3(n1069), .ZN(n1067) );
NOR2_X1 U769 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR2_X1 U770 ( .A1(n1066), .A2(n1072), .ZN(n1070) );
INV_X1 U771 ( .A(n966), .ZN(n1066) );
NOR3_X1 U772 ( .A1(n1073), .A2(n1072), .A3(n1063), .ZN(n1068) );
INV_X1 U773 ( .A(G478), .ZN(n1072) );
NOR2_X1 U774 ( .A1(n1058), .A2(n1074), .ZN(G60) );
XOR2_X1 U775 ( .A(n1075), .B(n1076), .Z(n1074) );
NAND4_X1 U776 ( .A1(n1077), .A2(KEYINPUT26), .A3(G475), .A4(n966), .ZN(n1075) );
XNOR2_X1 U777 ( .A(G902), .B(KEYINPUT10), .ZN(n1077) );
XNOR2_X1 U778 ( .A(G104), .B(n1078), .ZN(G6) );
NOR2_X1 U779 ( .A1(n1058), .A2(n1079), .ZN(G57) );
XOR2_X1 U780 ( .A(n1080), .B(n1081), .Z(n1079) );
XNOR2_X1 U781 ( .A(G101), .B(n1082), .ZN(n1081) );
XNOR2_X1 U782 ( .A(KEYINPUT41), .B(KEYINPUT30), .ZN(n1082) );
XNOR2_X1 U783 ( .A(n1083), .B(n1084), .ZN(n1080) );
XOR2_X1 U784 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U785 ( .A1(n1087), .A2(n1063), .ZN(n1085) );
NOR2_X1 U786 ( .A1(n1058), .A2(n1088), .ZN(G54) );
XOR2_X1 U787 ( .A(n1089), .B(n1090), .Z(n1088) );
XOR2_X1 U788 ( .A(n1091), .B(n1092), .Z(n1090) );
XOR2_X1 U789 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U790 ( .A1(G140), .A2(KEYINPUT57), .ZN(n1094) );
XOR2_X1 U791 ( .A(G110), .B(n1095), .Z(n1091) );
NOR4_X1 U792 ( .A1(KEYINPUT63), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1095) );
XNOR2_X1 U793 ( .A(KEYINPUT5), .B(n966), .ZN(n1098) );
XOR2_X1 U794 ( .A(n1099), .B(n1100), .Z(n1089) );
XNOR2_X1 U795 ( .A(n1101), .B(n1102), .ZN(n1099) );
NOR2_X1 U796 ( .A1(KEYINPUT50), .A2(n1028), .ZN(n1102) );
NOR2_X1 U797 ( .A1(n1058), .A2(n1103), .ZN(G51) );
XOR2_X1 U798 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U799 ( .A1(n1106), .A2(n1063), .ZN(n1105) );
NAND2_X1 U800 ( .A1(G902), .A2(n966), .ZN(n1063) );
NAND4_X1 U801 ( .A1(n1107), .A2(n1056), .A3(n1108), .A4(n1038), .ZN(n966) );
AND4_X1 U802 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1038) );
NOR4_X1 U803 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1112) );
INV_X1 U804 ( .A(n1117), .ZN(n1116) );
INV_X1 U805 ( .A(n1118), .ZN(n1115) );
AND2_X1 U806 ( .A1(n1119), .A2(KEYINPUT23), .ZN(n1114) );
NOR4_X1 U807 ( .A1(KEYINPUT23), .A2(n1120), .A3(n990), .A4(n1121), .ZN(n1113) );
NAND3_X1 U808 ( .A1(n988), .A2(n973), .A3(n1004), .ZN(n1120) );
NOR2_X1 U809 ( .A1(n1042), .A2(n1041), .ZN(n1108) );
INV_X1 U810 ( .A(n1122), .ZN(n1041) );
AND4_X1 U811 ( .A1(n1123), .A2(n1078), .A3(n1124), .A4(n1125), .ZN(n1056) );
NOR4_X1 U812 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n962), .ZN(n1125) );
AND3_X1 U813 ( .A1(n975), .A2(n1129), .A3(n1005), .ZN(n962) );
NAND2_X1 U814 ( .A1(n1130), .A2(n1131), .ZN(n1124) );
XNOR2_X1 U815 ( .A(KEYINPUT14), .B(n1132), .ZN(n1131) );
NAND3_X1 U816 ( .A1(n975), .A2(n1129), .A3(n1004), .ZN(n1078) );
NAND3_X1 U817 ( .A1(n1129), .A2(n974), .A3(n1133), .ZN(n1123) );
INV_X1 U818 ( .A(n1134), .ZN(n1129) );
XNOR2_X1 U819 ( .A(n1135), .B(KEYINPUT32), .ZN(n1107) );
NAND2_X1 U820 ( .A1(n1136), .A2(KEYINPUT46), .ZN(n1104) );
XNOR2_X1 U821 ( .A(n1052), .B(n1137), .ZN(n1136) );
NOR2_X1 U822 ( .A1(KEYINPUT28), .A2(n1138), .ZN(n1137) );
XOR2_X1 U823 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U824 ( .A1(n977), .A2(G952), .ZN(n1058) );
XNOR2_X1 U825 ( .A(G146), .B(n1117), .ZN(G48) );
NAND4_X1 U826 ( .A1(n1141), .A2(n1004), .A3(n973), .A4(n1121), .ZN(n1117) );
XOR2_X1 U827 ( .A(G143), .B(n1142), .Z(G45) );
NOR2_X1 U828 ( .A1(KEYINPUT18), .A2(n1118), .ZN(n1142) );
NAND4_X1 U829 ( .A1(n1143), .A2(n1133), .A3(n973), .A4(n1121), .ZN(n1118) );
XOR2_X1 U830 ( .A(n1144), .B(n1042), .Z(G42) );
AND3_X1 U831 ( .A1(n1145), .A2(n1004), .A3(n1146), .ZN(n1042) );
XNOR2_X1 U832 ( .A(G140), .B(KEYINPUT38), .ZN(n1144) );
XNOR2_X1 U833 ( .A(G137), .B(n1111), .ZN(G39) );
NAND4_X1 U834 ( .A1(n1147), .A2(n1148), .A3(n1146), .A4(n974), .ZN(n1111) );
XNOR2_X1 U835 ( .A(KEYINPUT4), .B(n1149), .ZN(n1147) );
XNOR2_X1 U836 ( .A(G134), .B(n1109), .ZN(G36) );
NAND3_X1 U837 ( .A1(n1146), .A2(n1005), .A3(n1133), .ZN(n1109) );
NAND3_X1 U838 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(G33) );
OR2_X1 U839 ( .A1(n1119), .A2(KEYINPUT33), .ZN(n1152) );
NAND3_X1 U840 ( .A1(KEYINPUT33), .A2(n1119), .A3(n1153), .ZN(n1151) );
NAND2_X1 U841 ( .A1(G131), .A2(n1154), .ZN(n1150) );
NAND2_X1 U842 ( .A1(KEYINPUT33), .A2(n1155), .ZN(n1154) );
XOR2_X1 U843 ( .A(KEYINPUT54), .B(n1119), .Z(n1155) );
AND3_X1 U844 ( .A1(n1146), .A2(n1004), .A3(n1133), .ZN(n1119) );
AND3_X1 U845 ( .A1(n973), .A2(n1121), .A3(n988), .ZN(n1146) );
INV_X1 U846 ( .A(n971), .ZN(n988) );
NAND2_X1 U847 ( .A1(n995), .A2(n1156), .ZN(n971) );
INV_X1 U848 ( .A(n1021), .ZN(n995) );
XNOR2_X1 U849 ( .A(G128), .B(n1110), .ZN(G30) );
NAND4_X1 U850 ( .A1(n1141), .A2(n1005), .A3(n1157), .A4(n1121), .ZN(n1110) );
XNOR2_X1 U851 ( .A(n1158), .B(n1159), .ZN(G3) );
NOR4_X1 U852 ( .A1(KEYINPUT43), .A2(n1003), .A3(n1134), .A4(n990), .ZN(n1159) );
INV_X1 U853 ( .A(n1133), .ZN(n990) );
XNOR2_X1 U854 ( .A(G125), .B(n1122), .ZN(G27) );
NAND4_X1 U855 ( .A1(n1004), .A2(n1130), .A3(n1145), .A4(n1160), .ZN(n1122) );
AND3_X1 U856 ( .A1(n983), .A2(n985), .A3(n1121), .ZN(n1160) );
NAND2_X1 U857 ( .A1(n972), .A2(n1161), .ZN(n1121) );
NAND3_X1 U858 ( .A1(G902), .A2(n1162), .A3(n1024), .ZN(n1161) );
NOR2_X1 U859 ( .A1(G900), .A2(n977), .ZN(n1024) );
INV_X1 U860 ( .A(n991), .ZN(n1145) );
XNOR2_X1 U861 ( .A(G122), .B(n1163), .ZN(G24) );
NAND2_X1 U862 ( .A1(KEYINPUT21), .A2(n1135), .ZN(n1163) );
INV_X1 U863 ( .A(n1057), .ZN(n1135) );
NAND3_X1 U864 ( .A1(n1164), .A2(n975), .A3(n1143), .ZN(n1057) );
NOR3_X1 U865 ( .A1(n1165), .A2(n1166), .A3(n993), .ZN(n1143) );
NOR2_X1 U866 ( .A1(n1149), .A2(n1148), .ZN(n975) );
NAND2_X1 U867 ( .A1(n1167), .A2(n1168), .ZN(G21) );
NAND2_X1 U868 ( .A1(n1128), .A2(n1169), .ZN(n1168) );
XOR2_X1 U869 ( .A(KEYINPUT31), .B(n1170), .Z(n1167) );
NOR2_X1 U870 ( .A1(n1128), .A2(n1169), .ZN(n1170) );
AND3_X1 U871 ( .A1(n1164), .A2(n974), .A3(n1141), .ZN(n1128) );
AND3_X1 U872 ( .A1(n1171), .A2(n1172), .A3(n1130), .ZN(n1141) );
OR2_X1 U873 ( .A1(n1133), .A2(KEYINPUT4), .ZN(n1172) );
NAND2_X1 U874 ( .A1(KEYINPUT4), .A2(n1173), .ZN(n1171) );
NAND2_X1 U875 ( .A1(n1148), .A2(n1149), .ZN(n1173) );
INV_X1 U876 ( .A(n1174), .ZN(n1148) );
XNOR2_X1 U877 ( .A(n1175), .B(n1176), .ZN(G18) );
NOR2_X1 U878 ( .A1(n993), .A2(n1132), .ZN(n1176) );
NAND3_X1 U879 ( .A1(n1133), .A2(n1005), .A3(n1164), .ZN(n1132) );
XNOR2_X1 U880 ( .A(n1127), .B(n1177), .ZN(G15) );
XNOR2_X1 U881 ( .A(G113), .B(KEYINPUT1), .ZN(n1177) );
AND4_X1 U882 ( .A1(n1164), .A2(n1133), .A3(n1004), .A4(n1130), .ZN(n1127) );
NOR2_X1 U883 ( .A1(n1178), .A2(n1166), .ZN(n1004) );
INV_X1 U884 ( .A(n1019), .ZN(n1166) );
NOR2_X1 U885 ( .A1(n1174), .A2(n1149), .ZN(n1133) );
AND3_X1 U886 ( .A1(n985), .A2(n1179), .A3(n983), .ZN(n1164) );
XOR2_X1 U887 ( .A(G110), .B(n1126), .Z(G12) );
NOR3_X1 U888 ( .A1(n1134), .A2(n1003), .A3(n991), .ZN(n1126) );
NAND2_X1 U889 ( .A1(n1174), .A2(n1149), .ZN(n991) );
XNOR2_X1 U890 ( .A(n1016), .B(n1017), .ZN(n1149) );
NAND2_X1 U891 ( .A1(G217), .A2(n1180), .ZN(n1017) );
NOR2_X1 U892 ( .A1(n1065), .A2(G902), .ZN(n1016) );
INV_X1 U893 ( .A(n1062), .ZN(n1065) );
XNOR2_X1 U894 ( .A(n1181), .B(n1182), .ZN(n1062) );
XNOR2_X1 U895 ( .A(n1169), .B(n1183), .ZN(n1182) );
XOR2_X1 U896 ( .A(G137), .B(G128), .Z(n1183) );
INV_X1 U897 ( .A(G119), .ZN(n1169) );
XOR2_X1 U898 ( .A(n1184), .B(n1185), .Z(n1181) );
XNOR2_X1 U899 ( .A(G110), .B(n1186), .ZN(n1185) );
NAND3_X1 U900 ( .A1(n1187), .A2(n977), .A3(G221), .ZN(n1186) );
NAND3_X1 U901 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1184) );
OR2_X1 U902 ( .A1(n1029), .A2(G146), .ZN(n1190) );
NAND2_X1 U903 ( .A1(KEYINPUT59), .A2(n1191), .ZN(n1189) );
NAND2_X1 U904 ( .A1(n1192), .A2(n1029), .ZN(n1191) );
XNOR2_X1 U905 ( .A(KEYINPUT15), .B(G146), .ZN(n1192) );
NAND2_X1 U906 ( .A1(n1193), .A2(n1194), .ZN(n1188) );
INV_X1 U907 ( .A(KEYINPUT59), .ZN(n1194) );
NAND2_X1 U908 ( .A1(n1195), .A2(n1196), .ZN(n1193) );
OR2_X1 U909 ( .A1(G146), .A2(KEYINPUT15), .ZN(n1196) );
NAND3_X1 U910 ( .A1(G146), .A2(n1029), .A3(KEYINPUT15), .ZN(n1195) );
XOR2_X1 U911 ( .A(n1018), .B(KEYINPUT9), .Z(n1174) );
XOR2_X1 U912 ( .A(n1197), .B(n1087), .Z(n1018) );
INV_X1 U913 ( .A(G472), .ZN(n1087) );
NAND2_X1 U914 ( .A1(n1198), .A2(n1096), .ZN(n1197) );
XOR2_X1 U915 ( .A(n1199), .B(n1200), .Z(n1198) );
XNOR2_X1 U916 ( .A(n1201), .B(n1158), .ZN(n1200) );
INV_X1 U917 ( .A(G101), .ZN(n1158) );
NAND2_X1 U918 ( .A1(n1086), .A2(n1202), .ZN(n1201) );
XOR2_X1 U919 ( .A(KEYINPUT42), .B(KEYINPUT13), .Z(n1202) );
NOR2_X1 U920 ( .A1(n1203), .A2(n1204), .ZN(n1086) );
INV_X1 U921 ( .A(G210), .ZN(n1203) );
NAND2_X1 U922 ( .A1(KEYINPUT56), .A2(n1083), .ZN(n1199) );
XNOR2_X1 U923 ( .A(n1205), .B(n1206), .ZN(n1083) );
XOR2_X1 U924 ( .A(n1207), .B(n1208), .Z(n1206) );
XNOR2_X1 U925 ( .A(n1028), .B(G113), .ZN(n1205) );
INV_X1 U926 ( .A(n974), .ZN(n1003) );
NAND2_X1 U927 ( .A1(n1209), .A2(n1210), .ZN(n974) );
OR3_X1 U928 ( .A1(n1178), .A2(n1019), .A3(KEYINPUT53), .ZN(n1210) );
INV_X1 U929 ( .A(n1165), .ZN(n1178) );
NAND2_X1 U930 ( .A1(KEYINPUT53), .A2(n1005), .ZN(n1209) );
NOR2_X1 U931 ( .A1(n1019), .A2(n1165), .ZN(n1005) );
XOR2_X1 U932 ( .A(n1020), .B(n1211), .Z(n1165) );
NOR2_X1 U933 ( .A1(G478), .A2(KEYINPUT49), .ZN(n1211) );
NOR2_X1 U934 ( .A1(n1071), .A2(G902), .ZN(n1020) );
INV_X1 U935 ( .A(n1073), .ZN(n1071) );
XNOR2_X1 U936 ( .A(n1212), .B(n1213), .ZN(n1073) );
XOR2_X1 U937 ( .A(n1214), .B(n1215), .Z(n1213) );
NAND2_X1 U938 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U939 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XNOR2_X1 U940 ( .A(G107), .B(n1220), .ZN(n1218) );
XNOR2_X1 U941 ( .A(KEYINPUT48), .B(KEYINPUT45), .ZN(n1220) );
NAND2_X1 U942 ( .A1(n1221), .A2(n1222), .ZN(n1216) );
XNOR2_X1 U943 ( .A(G107), .B(KEYINPUT39), .ZN(n1222) );
INV_X1 U944 ( .A(n1219), .ZN(n1221) );
NAND2_X1 U945 ( .A1(n1223), .A2(n1224), .ZN(n1219) );
OR2_X1 U946 ( .A1(n1175), .A2(G122), .ZN(n1224) );
XOR2_X1 U947 ( .A(n1225), .B(KEYINPUT25), .Z(n1223) );
NAND2_X1 U948 ( .A1(G122), .A2(n1175), .ZN(n1225) );
XOR2_X1 U949 ( .A(n1226), .B(G134), .Z(n1212) );
NAND3_X1 U950 ( .A1(n1187), .A2(n977), .A3(G217), .ZN(n1226) );
XOR2_X1 U951 ( .A(G234), .B(KEYINPUT37), .Z(n1187) );
XNOR2_X1 U952 ( .A(n1227), .B(G475), .ZN(n1019) );
NAND2_X1 U953 ( .A1(n1076), .A2(n1096), .ZN(n1227) );
XNOR2_X1 U954 ( .A(n1228), .B(n1229), .ZN(n1076) );
XOR2_X1 U955 ( .A(n1230), .B(n1029), .Z(n1229) );
XNOR2_X1 U956 ( .A(G125), .B(n1231), .ZN(n1029) );
XOR2_X1 U957 ( .A(n1232), .B(n1233), .Z(n1228) );
NAND2_X1 U958 ( .A1(KEYINPUT2), .A2(n1234), .ZN(n1232) );
XOR2_X1 U959 ( .A(n1235), .B(n1236), .Z(n1234) );
XNOR2_X1 U960 ( .A(G143), .B(n1153), .ZN(n1236) );
INV_X1 U961 ( .A(G131), .ZN(n1153) );
NOR2_X1 U962 ( .A1(n1204), .A2(n1237), .ZN(n1235) );
INV_X1 U963 ( .A(G214), .ZN(n1237) );
NAND2_X1 U964 ( .A1(n1238), .A2(n977), .ZN(n1204) );
XNOR2_X1 U965 ( .A(KEYINPUT58), .B(n1239), .ZN(n1238) );
NAND3_X1 U966 ( .A1(n1157), .A2(n1179), .A3(n1130), .ZN(n1134) );
INV_X1 U967 ( .A(n993), .ZN(n1130) );
NAND2_X1 U968 ( .A1(n1156), .A2(n1021), .ZN(n993) );
XOR2_X1 U969 ( .A(n1240), .B(n1106), .Z(n1021) );
NAND2_X1 U970 ( .A1(G210), .A2(n1241), .ZN(n1106) );
NAND2_X1 U971 ( .A1(n1242), .A2(n1096), .ZN(n1240) );
XOR2_X1 U972 ( .A(n1243), .B(n1244), .Z(n1242) );
XNOR2_X1 U973 ( .A(n1245), .B(KEYINPUT19), .ZN(n1244) );
NAND2_X1 U974 ( .A1(KEYINPUT52), .A2(n1139), .ZN(n1245) );
AND2_X1 U975 ( .A1(G224), .A2(n977), .ZN(n1139) );
XOR2_X1 U976 ( .A(n1246), .B(n1140), .Z(n1243) );
XNOR2_X1 U977 ( .A(n1247), .B(n1207), .ZN(n1140) );
XNOR2_X1 U978 ( .A(n1248), .B(G128), .ZN(n1207) );
NAND2_X1 U979 ( .A1(KEYINPUT36), .A2(n1249), .ZN(n1248) );
XNOR2_X1 U980 ( .A(n1032), .B(G143), .ZN(n1249) );
INV_X1 U981 ( .A(G125), .ZN(n1247) );
NAND2_X1 U982 ( .A1(KEYINPUT47), .A2(n1250), .ZN(n1246) );
INV_X1 U983 ( .A(n1052), .ZN(n1250) );
XNOR2_X1 U984 ( .A(n1251), .B(n1252), .ZN(n1052) );
XNOR2_X1 U985 ( .A(G104), .B(n1253), .ZN(n1252) );
XNOR2_X1 U986 ( .A(KEYINPUT55), .B(KEYINPUT0), .ZN(n1253) );
XOR2_X1 U987 ( .A(n1254), .B(n1230), .Z(n1251) );
XNOR2_X1 U988 ( .A(n1255), .B(G122), .ZN(n1230) );
INV_X1 U989 ( .A(G113), .ZN(n1255) );
XOR2_X1 U990 ( .A(n1256), .B(n1257), .Z(n1254) );
NOR3_X1 U991 ( .A1(KEYINPUT24), .A2(n1258), .A3(n1259), .ZN(n1257) );
AND3_X1 U992 ( .A1(KEYINPUT27), .A2(n1175), .A3(G119), .ZN(n1259) );
NOR2_X1 U993 ( .A1(KEYINPUT27), .A2(n1208), .ZN(n1258) );
XNOR2_X1 U994 ( .A(n1175), .B(G119), .ZN(n1208) );
INV_X1 U995 ( .A(G116), .ZN(n1175) );
XNOR2_X1 U996 ( .A(n996), .B(KEYINPUT44), .ZN(n1156) );
AND2_X1 U997 ( .A1(G214), .A2(n1241), .ZN(n996) );
NAND2_X1 U998 ( .A1(n1239), .A2(n1096), .ZN(n1241) );
INV_X1 U999 ( .A(G237), .ZN(n1239) );
NAND2_X1 U1000 ( .A1(n972), .A2(n1260), .ZN(n1179) );
NAND3_X1 U1001 ( .A1(n1054), .A2(n1162), .A3(G902), .ZN(n1260) );
AND2_X1 U1002 ( .A1(G953), .A2(n1261), .ZN(n1054) );
XOR2_X1 U1003 ( .A(KEYINPUT12), .B(G898), .Z(n1261) );
NAND3_X1 U1004 ( .A1(n1162), .A2(n977), .A3(G952), .ZN(n972) );
INV_X1 U1005 ( .A(G953), .ZN(n977) );
NAND2_X1 U1006 ( .A1(G234), .A2(G237), .ZN(n1162) );
XOR2_X1 U1007 ( .A(n973), .B(KEYINPUT11), .Z(n1157) );
NOR2_X1 U1008 ( .A1(n983), .A2(n1002), .ZN(n973) );
INV_X1 U1009 ( .A(n985), .ZN(n1002) );
NAND2_X1 U1010 ( .A1(G221), .A2(n1180), .ZN(n985) );
NAND2_X1 U1011 ( .A1(G234), .A2(n1096), .ZN(n1180) );
XNOR2_X1 U1012 ( .A(n1014), .B(KEYINPUT20), .ZN(n983) );
XNOR2_X1 U1013 ( .A(n1262), .B(n1097), .ZN(n1014) );
INV_X1 U1014 ( .A(G469), .ZN(n1097) );
NAND2_X1 U1015 ( .A1(n1263), .A2(n1096), .ZN(n1262) );
INV_X1 U1016 ( .A(G902), .ZN(n1096) );
XOR2_X1 U1017 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U1018 ( .A(n1266), .B(n1028), .Z(n1265) );
XOR2_X1 U1019 ( .A(G131), .B(n1267), .Z(n1028) );
XOR2_X1 U1020 ( .A(G137), .B(G134), .Z(n1267) );
XOR2_X1 U1021 ( .A(n1256), .B(n1100), .Z(n1266) );
XOR2_X1 U1022 ( .A(n1233), .B(n1030), .Z(n1100) );
XNOR2_X1 U1023 ( .A(n1214), .B(KEYINPUT29), .ZN(n1030) );
XNOR2_X1 U1024 ( .A(G128), .B(G143), .ZN(n1214) );
XNOR2_X1 U1025 ( .A(G104), .B(n1032), .ZN(n1233) );
INV_X1 U1026 ( .A(G146), .ZN(n1032) );
XNOR2_X1 U1027 ( .A(G110), .B(n1101), .ZN(n1256) );
XNOR2_X1 U1028 ( .A(G101), .B(n961), .ZN(n1101) );
INV_X1 U1029 ( .A(G107), .ZN(n961) );
XOR2_X1 U1030 ( .A(n1268), .B(n1269), .Z(n1264) );
XOR2_X1 U1031 ( .A(KEYINPUT51), .B(KEYINPUT40), .Z(n1269) );
XNOR2_X1 U1032 ( .A(n1270), .B(n1231), .ZN(n1268) );
INV_X1 U1033 ( .A(G140), .ZN(n1231) );
NAND2_X1 U1034 ( .A1(KEYINPUT61), .A2(n1093), .ZN(n1270) );
NOR2_X1 U1035 ( .A1(n1036), .A2(G953), .ZN(n1093) );
INV_X1 U1036 ( .A(G227), .ZN(n1036) );
endmodule


