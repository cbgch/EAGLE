//Key = 0100000000110010000000000100000111001001010110010010110010101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315;

XOR2_X1 U720 ( .A(G107), .B(n1001), .Z(G9) );
NOR2_X1 U721 ( .A1(n1002), .A2(n1003), .ZN(G75) );
AND3_X1 U722 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1003) );
NOR4_X1 U723 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1002) );
NOR2_X1 U724 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR4_X1 U725 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1011) );
NAND4_X1 U726 ( .A1(n1004), .A2(n1017), .A3(n1018), .A4(n1005), .ZN(n1007) );
NAND4_X1 U727 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
NAND2_X1 U728 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U729 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
INV_X1 U730 ( .A(KEYINPUT33), .ZN(n1026) );
NAND4_X1 U731 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1021) );
NAND2_X1 U732 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NAND2_X1 U733 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U734 ( .A1(KEYINPUT33), .A2(n1025), .ZN(n1028) );
NAND2_X1 U735 ( .A1(n1035), .A2(n1036), .ZN(n1017) );
NAND3_X1 U736 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NAND2_X1 U737 ( .A1(n1019), .A2(n1040), .ZN(n1039) );
NAND2_X1 U738 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND3_X1 U739 ( .A1(n1043), .A2(n1012), .A3(n1044), .ZN(n1042) );
INV_X1 U740 ( .A(KEYINPUT54), .ZN(n1012) );
NAND3_X1 U741 ( .A1(n1020), .A2(n1045), .A3(n1046), .ZN(n1037) );
INV_X1 U742 ( .A(n1016), .ZN(n1035) );
NAND3_X1 U743 ( .A1(n1047), .A2(n1031), .A3(n1030), .ZN(n1016) );
INV_X1 U744 ( .A(n1024), .ZN(n1030) );
NAND4_X1 U745 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1004) );
NOR4_X1 U746 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1051) );
XNOR2_X1 U747 ( .A(n1056), .B(n1057), .ZN(n1055) );
XOR2_X1 U748 ( .A(n1058), .B(KEYINPUT55), .Z(n1057) );
XOR2_X1 U749 ( .A(G475), .B(n1059), .Z(n1054) );
NOR2_X1 U750 ( .A1(KEYINPUT17), .A2(n1060), .ZN(n1059) );
XOR2_X1 U751 ( .A(n1061), .B(n1062), .Z(n1053) );
XOR2_X1 U752 ( .A(n1063), .B(KEYINPUT41), .Z(n1062) );
NAND2_X1 U753 ( .A1(KEYINPUT58), .A2(n1064), .ZN(n1061) );
AND3_X1 U754 ( .A1(n1065), .A2(n1066), .A3(n1015), .ZN(n1050) );
OR2_X1 U755 ( .A1(n1067), .A2(n1068), .ZN(n1049) );
XOR2_X1 U756 ( .A(n1069), .B(n1070), .Z(n1048) );
XOR2_X1 U757 ( .A(n1071), .B(KEYINPUT47), .Z(n1070) );
XOR2_X1 U758 ( .A(n1072), .B(n1073), .Z(G72) );
XOR2_X1 U759 ( .A(n1074), .B(n1075), .Z(n1073) );
NOR2_X1 U760 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U761 ( .A(KEYINPUT46), .B(G953), .Z(n1077) );
INV_X1 U762 ( .A(n1008), .ZN(n1076) );
NAND2_X1 U763 ( .A1(n1078), .A2(n1079), .ZN(n1074) );
NAND2_X1 U764 ( .A1(G953), .A2(n1080), .ZN(n1079) );
XOR2_X1 U765 ( .A(n1081), .B(n1082), .Z(n1078) );
XOR2_X1 U766 ( .A(KEYINPUT14), .B(G128), .Z(n1082) );
XOR2_X1 U767 ( .A(n1083), .B(n1084), .Z(n1081) );
NOR2_X1 U768 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U769 ( .A(KEYINPUT18), .B(n1087), .Z(n1086) );
NOR2_X1 U770 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
AND2_X1 U771 ( .A1(n1088), .A2(n1089), .ZN(n1085) );
XOR2_X1 U772 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND2_X1 U773 ( .A1(G953), .A2(n1092), .ZN(n1072) );
NAND2_X1 U774 ( .A1(G900), .A2(G227), .ZN(n1092) );
XOR2_X1 U775 ( .A(n1093), .B(n1094), .Z(G69) );
NOR2_X1 U776 ( .A1(n1095), .A2(n1005), .ZN(n1094) );
NOR2_X1 U777 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U778 ( .A1(n1098), .A2(n1099), .ZN(n1093) );
NAND2_X1 U779 ( .A1(n1100), .A2(n1005), .ZN(n1099) );
XNOR2_X1 U780 ( .A(n1010), .B(n1101), .ZN(n1100) );
OR3_X1 U781 ( .A1(n1097), .A2(n1101), .A3(n1005), .ZN(n1098) );
XNOR2_X1 U782 ( .A(n1102), .B(n1103), .ZN(n1101) );
XNOR2_X1 U783 ( .A(n1104), .B(n1105), .ZN(n1103) );
XNOR2_X1 U784 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n1105) );
XOR2_X1 U785 ( .A(n1106), .B(n1107), .Z(n1102) );
NOR2_X1 U786 ( .A1(n1108), .A2(n1109), .ZN(G66) );
XOR2_X1 U787 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U788 ( .A1(n1067), .A2(n1112), .ZN(n1110) );
NOR2_X1 U789 ( .A1(n1108), .A2(n1113), .ZN(G63) );
XOR2_X1 U790 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U791 ( .A1(n1116), .A2(n1112), .ZN(n1115) );
NOR2_X1 U792 ( .A1(n1108), .A2(n1117), .ZN(G60) );
XNOR2_X1 U793 ( .A(n1118), .B(n1119), .ZN(n1117) );
NOR2_X1 U794 ( .A1(n1120), .A2(n1112), .ZN(n1119) );
INV_X1 U795 ( .A(G475), .ZN(n1120) );
XOR2_X1 U796 ( .A(G104), .B(n1121), .Z(G6) );
NOR2_X1 U797 ( .A1(n1108), .A2(n1122), .ZN(G57) );
XOR2_X1 U798 ( .A(n1123), .B(n1124), .Z(n1122) );
XNOR2_X1 U799 ( .A(n1125), .B(n1126), .ZN(n1124) );
NOR2_X1 U800 ( .A1(KEYINPUT42), .A2(n1127), .ZN(n1126) );
NAND2_X1 U801 ( .A1(KEYINPUT53), .A2(n1128), .ZN(n1125) );
XOR2_X1 U802 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U803 ( .A1(n1063), .A2(n1112), .ZN(n1129) );
INV_X1 U804 ( .A(G472), .ZN(n1063) );
NOR2_X1 U805 ( .A1(n1108), .A2(n1131), .ZN(G54) );
XOR2_X1 U806 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U807 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U808 ( .A1(n1058), .A2(n1112), .ZN(n1135) );
INV_X1 U809 ( .A(G469), .ZN(n1058) );
NOR2_X1 U810 ( .A1(n1136), .A2(n1137), .ZN(n1134) );
NOR2_X1 U811 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR2_X1 U812 ( .A1(KEYINPUT2), .A2(n1140), .ZN(n1139) );
NOR2_X1 U813 ( .A1(n1141), .A2(n1142), .ZN(n1138) );
AND2_X1 U814 ( .A1(n1140), .A2(KEYINPUT63), .ZN(n1141) );
NOR4_X1 U815 ( .A1(KEYINPUT63), .A2(KEYINPUT2), .A3(n1142), .A4(n1140), .ZN(n1136) );
XNOR2_X1 U816 ( .A(n1143), .B(n1144), .ZN(n1140) );
XOR2_X1 U817 ( .A(n1145), .B(G146), .Z(n1143) );
NOR2_X1 U818 ( .A1(n1146), .A2(n1147), .ZN(n1132) );
NOR2_X1 U819 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U820 ( .A(KEYINPUT44), .B(n1150), .Z(n1148) );
NOR2_X1 U821 ( .A1(n1150), .A2(n1151), .ZN(n1146) );
INV_X1 U822 ( .A(n1149), .ZN(n1151) );
XNOR2_X1 U823 ( .A(G140), .B(G110), .ZN(n1149) );
NOR2_X1 U824 ( .A1(n1108), .A2(n1152), .ZN(G51) );
XOR2_X1 U825 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U826 ( .A(n1155), .B(n1156), .Z(n1153) );
NOR2_X1 U827 ( .A1(n1071), .A2(n1112), .ZN(n1156) );
NAND2_X1 U828 ( .A1(G902), .A2(n1157), .ZN(n1112) );
OR2_X1 U829 ( .A1(n1008), .A2(n1010), .ZN(n1157) );
NAND2_X1 U830 ( .A1(n1158), .A2(n1159), .ZN(n1010) );
AND4_X1 U831 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1159) );
NOR4_X1 U832 ( .A1(n1001), .A2(n1164), .A3(n1121), .A4(n1165), .ZN(n1158) );
NOR2_X1 U833 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U834 ( .A(n1168), .B(KEYINPUT12), .Z(n1166) );
AND2_X1 U835 ( .A1(n1169), .A2(n1170), .ZN(n1121) );
NOR3_X1 U836 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1164) );
XOR2_X1 U837 ( .A(n1167), .B(KEYINPUT20), .Z(n1173) );
AND2_X1 U838 ( .A1(n1174), .A2(n1170), .ZN(n1001) );
AND4_X1 U839 ( .A1(n1175), .A2(n1031), .A3(n1176), .A4(n1177), .ZN(n1170) );
NAND4_X1 U840 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1008) );
NOR4_X1 U841 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181) );
INV_X1 U842 ( .A(n1186), .ZN(n1183) );
NAND3_X1 U843 ( .A1(n1169), .A2(n1187), .A3(n1019), .ZN(n1180) );
NAND2_X1 U844 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NAND3_X1 U845 ( .A1(n1190), .A2(n1176), .A3(n1191), .ZN(n1189) );
XNOR2_X1 U846 ( .A(KEYINPUT31), .B(n1192), .ZN(n1191) );
NAND2_X1 U847 ( .A1(n1193), .A2(n1194), .ZN(n1188) );
AND2_X1 U848 ( .A1(n1195), .A2(n1006), .ZN(n1108) );
INV_X1 U849 ( .A(G952), .ZN(n1006) );
XOR2_X1 U850 ( .A(KEYINPUT5), .B(G953), .Z(n1195) );
XNOR2_X1 U851 ( .A(G146), .B(n1196), .ZN(G48) );
NAND2_X1 U852 ( .A1(KEYINPUT61), .A2(n1185), .ZN(n1196) );
AND2_X1 U853 ( .A1(n1197), .A2(n1169), .ZN(n1185) );
XNOR2_X1 U854 ( .A(G143), .B(n1178), .ZN(G45) );
NAND4_X1 U855 ( .A1(n1190), .A2(n1176), .A3(n1175), .A4(n1198), .ZN(n1178) );
AND3_X1 U856 ( .A1(n1199), .A2(n1192), .A3(n1052), .ZN(n1198) );
XNOR2_X1 U857 ( .A(G140), .B(n1200), .ZN(G42) );
NAND4_X1 U858 ( .A1(n1193), .A2(n1169), .A3(n1194), .A4(n1201), .ZN(n1200) );
XOR2_X1 U859 ( .A(KEYINPUT51), .B(n1019), .Z(n1201) );
XNOR2_X1 U860 ( .A(n1179), .B(n1202), .ZN(G39) );
NOR2_X1 U861 ( .A1(KEYINPUT13), .A2(n1091), .ZN(n1202) );
NAND4_X1 U862 ( .A1(n1047), .A2(n1019), .A3(n1193), .A4(n1203), .ZN(n1179) );
XOR2_X1 U863 ( .A(G134), .B(n1184), .Z(G36) );
NOR2_X1 U864 ( .A1(n1204), .A2(n1034), .ZN(n1184) );
INV_X1 U865 ( .A(n1174), .ZN(n1034) );
XOR2_X1 U866 ( .A(n1205), .B(n1206), .Z(G33) );
NOR2_X1 U867 ( .A1(KEYINPUT28), .A2(n1207), .ZN(n1206) );
NOR2_X1 U868 ( .A1(n1033), .A2(n1204), .ZN(n1205) );
NAND4_X1 U869 ( .A1(n1019), .A2(n1190), .A3(n1176), .A4(n1192), .ZN(n1204) );
INV_X1 U870 ( .A(n1013), .ZN(n1019) );
NAND2_X1 U871 ( .A1(n1045), .A2(n1065), .ZN(n1013) );
XOR2_X1 U872 ( .A(n1208), .B(n1186), .Z(G30) );
NAND2_X1 U873 ( .A1(n1197), .A2(n1174), .ZN(n1186) );
AND3_X1 U874 ( .A1(n1175), .A2(n1203), .A3(n1193), .ZN(n1197) );
AND3_X1 U875 ( .A1(n1192), .A2(n1209), .A3(n1176), .ZN(n1193) );
XNOR2_X1 U876 ( .A(G101), .B(n1163), .ZN(G3) );
OR4_X1 U877 ( .A1(n1027), .A2(n1167), .A3(n1041), .A4(n1172), .ZN(n1163) );
INV_X1 U878 ( .A(n1176), .ZN(n1041) );
NAND2_X1 U879 ( .A1(n1047), .A2(n1190), .ZN(n1027) );
XNOR2_X1 U880 ( .A(G125), .B(n1210), .ZN(G27) );
NAND2_X1 U881 ( .A1(KEYINPUT56), .A2(n1182), .ZN(n1210) );
NOR3_X1 U882 ( .A1(n1038), .A2(n1033), .A3(n1211), .ZN(n1182) );
NAND3_X1 U883 ( .A1(n1194), .A2(n1209), .A3(n1192), .ZN(n1211) );
NAND2_X1 U884 ( .A1(n1024), .A2(n1212), .ZN(n1192) );
NAND2_X1 U885 ( .A1(n1213), .A2(n1080), .ZN(n1212) );
INV_X1 U886 ( .A(G900), .ZN(n1080) );
XOR2_X1 U887 ( .A(G122), .B(n1214), .Z(G24) );
NOR3_X1 U888 ( .A1(n1215), .A2(n1167), .A3(n1171), .ZN(n1214) );
NAND4_X1 U889 ( .A1(n1031), .A2(n1020), .A3(n1199), .A4(n1052), .ZN(n1171) );
XOR2_X1 U890 ( .A(KEYINPUT29), .B(n1172), .Z(n1215) );
XNOR2_X1 U891 ( .A(G119), .B(n1162), .ZN(G21) );
NAND4_X1 U892 ( .A1(n1216), .A2(n1047), .A3(n1203), .A4(n1209), .ZN(n1162) );
XNOR2_X1 U893 ( .A(n1161), .B(n1217), .ZN(G18) );
NOR2_X1 U894 ( .A1(KEYINPUT62), .A2(n1218), .ZN(n1217) );
NAND3_X1 U895 ( .A1(n1174), .A2(n1190), .A3(n1216), .ZN(n1161) );
NOR2_X1 U896 ( .A1(n1199), .A2(n1219), .ZN(n1174) );
XOR2_X1 U897 ( .A(n1220), .B(n1160), .Z(G15) );
NAND3_X1 U898 ( .A1(n1169), .A2(n1190), .A3(n1216), .ZN(n1160) );
NOR2_X1 U899 ( .A1(n1038), .A2(n1172), .ZN(n1216) );
INV_X1 U900 ( .A(n1177), .ZN(n1172) );
NAND2_X1 U901 ( .A1(n1175), .A2(n1020), .ZN(n1038) );
NAND2_X1 U902 ( .A1(n1221), .A2(n1222), .ZN(n1190) );
OR3_X1 U903 ( .A1(n1209), .A2(n1194), .A3(KEYINPUT15), .ZN(n1222) );
NAND2_X1 U904 ( .A1(KEYINPUT15), .A2(n1031), .ZN(n1221) );
NOR2_X1 U905 ( .A1(n1209), .A2(n1203), .ZN(n1031) );
INV_X1 U906 ( .A(n1194), .ZN(n1203) );
INV_X1 U907 ( .A(n1033), .ZN(n1169) );
NAND2_X1 U908 ( .A1(n1219), .A2(n1199), .ZN(n1033) );
XOR2_X1 U909 ( .A(G110), .B(n1223), .Z(G12) );
NOR2_X1 U910 ( .A1(n1167), .A2(n1168), .ZN(n1223) );
NAND3_X1 U911 ( .A1(n1176), .A2(n1177), .A3(n1025), .ZN(n1168) );
AND3_X1 U912 ( .A1(n1194), .A2(n1209), .A3(n1047), .ZN(n1025) );
NOR2_X1 U913 ( .A1(n1052), .A2(n1199), .ZN(n1047) );
XNOR2_X1 U914 ( .A(n1060), .B(G475), .ZN(n1199) );
NAND2_X1 U915 ( .A1(n1118), .A2(n1224), .ZN(n1060) );
XNOR2_X1 U916 ( .A(n1225), .B(n1226), .ZN(n1118) );
XOR2_X1 U917 ( .A(n1227), .B(n1228), .Z(n1226) );
XNOR2_X1 U918 ( .A(KEYINPUT43), .B(n1229), .ZN(n1228) );
NOR3_X1 U919 ( .A1(KEYINPUT27), .A2(n1230), .A3(n1231), .ZN(n1229) );
NOR2_X1 U920 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
INV_X1 U921 ( .A(G122), .ZN(n1233) );
XOR2_X1 U922 ( .A(KEYINPUT10), .B(n1234), .Z(n1232) );
NOR2_X1 U923 ( .A1(G122), .A2(n1235), .ZN(n1230) );
XNOR2_X1 U924 ( .A(n1234), .B(KEYINPUT36), .ZN(n1235) );
XNOR2_X1 U925 ( .A(n1220), .B(n1236), .ZN(n1234) );
NOR2_X1 U926 ( .A1(KEYINPUT21), .A2(n1237), .ZN(n1236) );
NAND2_X1 U927 ( .A1(G214), .A2(n1238), .ZN(n1227) );
XOR2_X1 U928 ( .A(n1083), .B(n1088), .Z(n1225) );
INV_X1 U929 ( .A(n1239), .ZN(n1088) );
XNOR2_X1 U930 ( .A(n1240), .B(n1241), .ZN(n1083) );
INV_X1 U931 ( .A(n1219), .ZN(n1052) );
XOR2_X1 U932 ( .A(n1116), .B(n1242), .Z(n1219) );
NOR2_X1 U933 ( .A1(G902), .A2(n1114), .ZN(n1242) );
XOR2_X1 U934 ( .A(n1243), .B(n1244), .Z(n1114) );
NOR2_X1 U935 ( .A1(KEYINPUT30), .A2(n1245), .ZN(n1244) );
XOR2_X1 U936 ( .A(n1246), .B(n1144), .Z(n1245) );
XOR2_X1 U937 ( .A(G128), .B(n1247), .Z(n1144) );
XOR2_X1 U938 ( .A(n1248), .B(G134), .Z(n1246) );
NAND2_X1 U939 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
NAND2_X1 U940 ( .A1(G107), .A2(n1251), .ZN(n1250) );
XOR2_X1 U941 ( .A(n1252), .B(KEYINPUT35), .Z(n1249) );
OR2_X1 U942 ( .A1(n1251), .A2(G107), .ZN(n1252) );
XNOR2_X1 U943 ( .A(n1218), .B(n1253), .ZN(n1251) );
XOR2_X1 U944 ( .A(KEYINPUT57), .B(G122), .Z(n1253) );
NAND2_X1 U945 ( .A1(G217), .A2(n1254), .ZN(n1243) );
INV_X1 U946 ( .A(G478), .ZN(n1116) );
NAND3_X1 U947 ( .A1(n1255), .A2(n1256), .A3(n1066), .ZN(n1209) );
NAND2_X1 U948 ( .A1(n1068), .A2(n1067), .ZN(n1066) );
OR3_X1 U949 ( .A1(n1067), .A2(n1068), .A3(KEYINPUT34), .ZN(n1256) );
NOR2_X1 U950 ( .A1(n1111), .A2(G902), .ZN(n1068) );
XNOR2_X1 U951 ( .A(n1257), .B(n1258), .ZN(n1111) );
XOR2_X1 U952 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U953 ( .A(n1208), .B(n1261), .Z(n1260) );
NOR2_X1 U954 ( .A1(KEYINPUT26), .A2(n1262), .ZN(n1261) );
XOR2_X1 U955 ( .A(n1263), .B(G137), .Z(n1262) );
NAND2_X1 U956 ( .A1(G221), .A2(n1254), .ZN(n1263) );
AND2_X1 U957 ( .A1(G234), .A2(n1005), .ZN(n1254) );
INV_X1 U958 ( .A(G128), .ZN(n1208) );
NAND2_X1 U959 ( .A1(KEYINPUT52), .A2(n1240), .ZN(n1259) );
XNOR2_X1 U960 ( .A(n1264), .B(n1107), .ZN(n1257) );
XOR2_X1 U961 ( .A(G110), .B(G119), .Z(n1107) );
NAND2_X1 U962 ( .A1(KEYINPUT34), .A2(n1067), .ZN(n1255) );
NAND2_X1 U963 ( .A1(G217), .A2(n1265), .ZN(n1067) );
XOR2_X1 U964 ( .A(n1064), .B(G472), .Z(n1194) );
NAND2_X1 U965 ( .A1(n1266), .A2(n1224), .ZN(n1064) );
XOR2_X1 U966 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U967 ( .A(n1130), .B(n1123), .Z(n1268) );
XNOR2_X1 U968 ( .A(n1269), .B(n1270), .ZN(n1130) );
XOR2_X1 U969 ( .A(n1142), .B(n1271), .Z(n1270) );
XOR2_X1 U970 ( .A(n1220), .B(n1272), .Z(n1269) );
NOR2_X1 U971 ( .A1(KEYINPUT38), .A2(n1273), .ZN(n1272) );
XOR2_X1 U972 ( .A(n1218), .B(G119), .Z(n1273) );
INV_X1 U973 ( .A(G116), .ZN(n1218) );
INV_X1 U974 ( .A(G113), .ZN(n1220) );
XOR2_X1 U975 ( .A(n1127), .B(KEYINPUT19), .Z(n1267) );
NAND2_X1 U976 ( .A1(G210), .A2(n1238), .ZN(n1127) );
NOR2_X1 U977 ( .A1(G953), .A2(G237), .ZN(n1238) );
NAND2_X1 U978 ( .A1(n1024), .A2(n1274), .ZN(n1177) );
NAND2_X1 U979 ( .A1(n1213), .A2(n1097), .ZN(n1274) );
INV_X1 U980 ( .A(G898), .ZN(n1097) );
AND3_X1 U981 ( .A1(G953), .A2(n1275), .A3(n1276), .ZN(n1213) );
XOR2_X1 U982 ( .A(n1224), .B(KEYINPUT11), .Z(n1276) );
NAND3_X1 U983 ( .A1(n1275), .A2(n1005), .A3(G952), .ZN(n1024) );
NAND2_X1 U984 ( .A1(G237), .A2(G234), .ZN(n1275) );
NAND2_X1 U985 ( .A1(n1277), .A2(n1278), .ZN(n1176) );
OR3_X1 U986 ( .A1(n1043), .A2(n1044), .A3(KEYINPUT16), .ZN(n1278) );
NAND2_X1 U987 ( .A1(KEYINPUT16), .A2(n1020), .ZN(n1277) );
NOR2_X1 U988 ( .A1(n1014), .A2(n1044), .ZN(n1020) );
INV_X1 U989 ( .A(n1015), .ZN(n1044) );
NAND2_X1 U990 ( .A1(G221), .A2(n1265), .ZN(n1015) );
NAND2_X1 U991 ( .A1(G234), .A2(n1224), .ZN(n1265) );
INV_X1 U992 ( .A(n1043), .ZN(n1014) );
XOR2_X1 U993 ( .A(n1279), .B(G469), .Z(n1043) );
NAND2_X1 U994 ( .A1(KEYINPUT1), .A2(n1056), .ZN(n1279) );
AND2_X1 U995 ( .A1(n1280), .A2(n1224), .ZN(n1056) );
XOR2_X1 U996 ( .A(n1281), .B(n1282), .Z(n1280) );
XOR2_X1 U997 ( .A(n1145), .B(n1283), .Z(n1282) );
XOR2_X1 U998 ( .A(n1150), .B(n1241), .Z(n1283) );
XOR2_X1 U999 ( .A(n1247), .B(n1264), .Z(n1241) );
XOR2_X1 U1000 ( .A(G140), .B(G146), .Z(n1264) );
AND2_X1 U1001 ( .A1(G227), .A2(n1005), .ZN(n1150) );
INV_X1 U1002 ( .A(G953), .ZN(n1005) );
XNOR2_X1 U1003 ( .A(n1284), .B(n1285), .ZN(n1145) );
XOR2_X1 U1004 ( .A(n1286), .B(n1287), .Z(n1281) );
XOR2_X1 U1005 ( .A(KEYINPUT25), .B(G128), .Z(n1287) );
XOR2_X1 U1006 ( .A(n1288), .B(G110), .Z(n1286) );
NAND2_X1 U1007 ( .A1(KEYINPUT50), .A2(n1142), .ZN(n1288) );
XOR2_X1 U1008 ( .A(n1289), .B(n1239), .Z(n1142) );
XOR2_X1 U1009 ( .A(n1207), .B(KEYINPUT59), .Z(n1239) );
INV_X1 U1010 ( .A(G131), .ZN(n1207) );
XOR2_X1 U1011 ( .A(n1290), .B(KEYINPUT6), .Z(n1289) );
NAND2_X1 U1012 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
NAND2_X1 U1013 ( .A1(G134), .A2(n1091), .ZN(n1292) );
INV_X1 U1014 ( .A(G137), .ZN(n1091) );
XOR2_X1 U1015 ( .A(n1293), .B(KEYINPUT4), .Z(n1291) );
NAND2_X1 U1016 ( .A1(G137), .A2(n1090), .ZN(n1293) );
INV_X1 U1017 ( .A(G134), .ZN(n1090) );
INV_X1 U1018 ( .A(n1175), .ZN(n1167) );
NOR2_X1 U1019 ( .A1(n1045), .A2(n1046), .ZN(n1175) );
INV_X1 U1020 ( .A(n1065), .ZN(n1046) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1294), .ZN(n1065) );
XNOR2_X1 U1022 ( .A(n1071), .B(n1295), .ZN(n1045) );
NOR2_X1 U1023 ( .A1(KEYINPUT45), .A2(n1296), .ZN(n1295) );
XNOR2_X1 U1024 ( .A(KEYINPUT8), .B(n1069), .ZN(n1296) );
NAND2_X1 U1025 ( .A1(n1297), .A2(n1224), .ZN(n1069) );
XOR2_X1 U1026 ( .A(n1155), .B(n1298), .Z(n1297) );
NOR2_X1 U1027 ( .A1(KEYINPUT7), .A2(n1154), .ZN(n1298) );
XOR2_X1 U1028 ( .A(n1240), .B(n1299), .Z(n1154) );
XOR2_X1 U1029 ( .A(n1300), .B(n1271), .Z(n1299) );
XNOR2_X1 U1030 ( .A(n1301), .B(n1302), .ZN(n1271) );
XOR2_X1 U1031 ( .A(G146), .B(n1303), .Z(n1302) );
NOR2_X1 U1032 ( .A1(KEYINPUT40), .A2(n1247), .ZN(n1303) );
XOR2_X1 U1033 ( .A(G143), .B(KEYINPUT48), .Z(n1247) );
NAND2_X1 U1034 ( .A1(KEYINPUT39), .A2(G128), .ZN(n1301) );
NOR2_X1 U1035 ( .A1(G953), .A2(n1096), .ZN(n1300) );
INV_X1 U1036 ( .A(G224), .ZN(n1096) );
XOR2_X1 U1037 ( .A(G125), .B(KEYINPUT60), .Z(n1240) );
XOR2_X1 U1038 ( .A(n1106), .B(n1304), .Z(n1155) );
XOR2_X1 U1039 ( .A(G119), .B(n1305), .Z(n1304) );
NOR2_X1 U1040 ( .A1(KEYINPUT24), .A2(n1306), .ZN(n1305) );
XNOR2_X1 U1041 ( .A(G110), .B(n1104), .ZN(n1306) );
NOR2_X1 U1042 ( .A1(KEYINPUT0), .A2(G122), .ZN(n1104) );
XOR2_X1 U1043 ( .A(n1307), .B(n1308), .Z(n1106) );
XOR2_X1 U1044 ( .A(G113), .B(n1309), .Z(n1308) );
NOR2_X1 U1045 ( .A1(G116), .A2(n1310), .ZN(n1309) );
XNOR2_X1 U1046 ( .A(KEYINPUT49), .B(KEYINPUT32), .ZN(n1310) );
NAND2_X1 U1047 ( .A1(n1311), .A2(n1312), .ZN(n1307) );
OR2_X1 U1048 ( .A1(n1284), .A2(n1285), .ZN(n1312) );
NAND2_X1 U1049 ( .A1(n1313), .A2(n1285), .ZN(n1311) );
XNOR2_X1 U1050 ( .A(n1237), .B(KEYINPUT9), .ZN(n1285) );
INV_X1 U1051 ( .A(G104), .ZN(n1237) );
XOR2_X1 U1052 ( .A(KEYINPUT37), .B(n1284), .Z(n1313) );
XOR2_X1 U1053 ( .A(G107), .B(n1314), .Z(n1284) );
INV_X1 U1054 ( .A(n1123), .ZN(n1314) );
XNOR2_X1 U1055 ( .A(G101), .B(KEYINPUT3), .ZN(n1123) );
NAND2_X1 U1056 ( .A1(G210), .A2(n1294), .ZN(n1071) );
NAND2_X1 U1057 ( .A1(n1315), .A2(n1224), .ZN(n1294) );
INV_X1 U1058 ( .A(G902), .ZN(n1224) );
INV_X1 U1059 ( .A(G237), .ZN(n1315) );
endmodule


