//Key = 0000111111001011101000100111101100001010000100111100100110111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318;

XNOR2_X1 U734 ( .A(G107), .B(n1003), .ZN(G9) );
NAND4_X1 U735 ( .A1(n1004), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n1003) );
AND2_X1 U736 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
XNOR2_X1 U737 ( .A(KEYINPUT43), .B(n1010), .ZN(n1004) );
NOR2_X1 U738 ( .A1(n1011), .A2(n1012), .ZN(G75) );
NOR4_X1 U739 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
XOR2_X1 U740 ( .A(n1017), .B(KEYINPUT63), .Z(n1015) );
NAND2_X1 U741 ( .A1(n1018), .A2(n1008), .ZN(n1017) );
XOR2_X1 U742 ( .A(n1019), .B(KEYINPUT56), .Z(n1018) );
NAND4_X1 U743 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1013) );
OR3_X1 U744 ( .A1(n1024), .A2(n1025), .A3(n1019), .ZN(n1021) );
NAND3_X1 U745 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1019) );
NAND3_X1 U746 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1020) );
NAND2_X1 U747 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NAND3_X1 U748 ( .A1(n1026), .A2(n1009), .A3(KEYINPUT13), .ZN(n1032) );
NAND3_X1 U749 ( .A1(n1034), .A2(n1035), .A3(n1028), .ZN(n1029) );
INV_X1 U750 ( .A(n1033), .ZN(n1028) );
NAND2_X1 U751 ( .A1(n1026), .A2(n1036), .ZN(n1035) );
NAND2_X1 U752 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U753 ( .A1(n1009), .A2(n1039), .ZN(n1038) );
INV_X1 U754 ( .A(KEYINPUT13), .ZN(n1039) );
NAND2_X1 U755 ( .A1(n1027), .A2(n1040), .ZN(n1034) );
NAND3_X1 U756 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NAND2_X1 U757 ( .A1(n1005), .A2(n1044), .ZN(n1043) );
NAND2_X1 U758 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U759 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U760 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1041) );
NOR3_X1 U761 ( .A1(n1052), .A2(G953), .A3(n1053), .ZN(n1011) );
INV_X1 U762 ( .A(n1022), .ZN(n1053) );
NAND4_X1 U763 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1022) );
NOR4_X1 U764 ( .A1(n1058), .A2(n1059), .A3(n1047), .A4(n1060), .ZN(n1057) );
NAND3_X1 U765 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1058) );
NAND2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND3_X1 U767 ( .A1(n1066), .A2(n1067), .A3(G217), .ZN(n1062) );
NAND2_X1 U768 ( .A1(n1068), .A2(G469), .ZN(n1061) );
NOR3_X1 U769 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1056) );
NOR2_X1 U770 ( .A1(KEYINPUT52), .A2(n1072), .ZN(n1071) );
XOR2_X1 U771 ( .A(n1073), .B(KEYINPUT18), .Z(n1070) );
NOR2_X1 U772 ( .A1(n1074), .A2(n1075), .ZN(n1055) );
NOR2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
INV_X1 U774 ( .A(KEYINPUT15), .ZN(n1077) );
NOR2_X1 U775 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NOR3_X1 U776 ( .A1(n1080), .A2(n1064), .A3(n1065), .ZN(n1079) );
NOR2_X1 U777 ( .A1(KEYINPUT4), .A2(n1081), .ZN(n1078) );
NOR2_X1 U778 ( .A1(KEYINPUT15), .A2(n1082), .ZN(n1074) );
NOR2_X1 U779 ( .A1(n1064), .A2(n1083), .ZN(n1082) );
XNOR2_X1 U780 ( .A(n1080), .B(n1081), .ZN(n1083) );
INV_X1 U781 ( .A(n1065), .ZN(n1081) );
INV_X1 U782 ( .A(KEYINPUT4), .ZN(n1080) );
NOR3_X1 U783 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1054) );
NOR2_X1 U784 ( .A1(G475), .A2(n1087), .ZN(n1086) );
NOR2_X1 U785 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XNOR2_X1 U786 ( .A(KEYINPUT53), .B(n1072), .ZN(n1089) );
INV_X1 U787 ( .A(n1090), .ZN(n1072) );
NOR3_X1 U788 ( .A1(n1091), .A2(n1090), .A3(n1088), .ZN(n1085) );
INV_X1 U789 ( .A(KEYINPUT52), .ZN(n1088) );
XOR2_X1 U790 ( .A(KEYINPUT33), .B(n1092), .Z(n1084) );
NOR2_X1 U791 ( .A1(G469), .A2(n1068), .ZN(n1092) );
XOR2_X1 U792 ( .A(n1093), .B(KEYINPUT35), .Z(n1068) );
XNOR2_X1 U793 ( .A(G952), .B(KEYINPUT25), .ZN(n1052) );
XOR2_X1 U794 ( .A(n1094), .B(n1095), .Z(G72) );
NOR2_X1 U795 ( .A1(n1096), .A2(n1023), .ZN(n1095) );
AND2_X1 U796 ( .A1(G227), .A2(G900), .ZN(n1096) );
NAND2_X1 U797 ( .A1(n1097), .A2(n1098), .ZN(n1094) );
NAND2_X1 U798 ( .A1(n1099), .A2(n1023), .ZN(n1098) );
XNOR2_X1 U799 ( .A(n1100), .B(n1101), .ZN(n1099) );
NAND3_X1 U800 ( .A1(G900), .A2(n1101), .A3(G953), .ZN(n1097) );
XOR2_X1 U801 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U802 ( .A(n1104), .B(n1105), .Z(G69) );
NOR2_X1 U803 ( .A1(n1106), .A2(n1023), .ZN(n1105) );
AND2_X1 U804 ( .A1(G224), .A2(G898), .ZN(n1106) );
NAND2_X1 U805 ( .A1(n1107), .A2(KEYINPUT8), .ZN(n1104) );
XOR2_X1 U806 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR3_X1 U807 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
NOR2_X1 U808 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U809 ( .A(KEYINPUT39), .B(n1115), .Z(n1114) );
XNOR2_X1 U810 ( .A(n1116), .B(n1117), .ZN(n1113) );
NOR2_X1 U811 ( .A1(n1118), .A2(n1119), .ZN(n1111) );
XOR2_X1 U812 ( .A(KEYINPUT49), .B(n1115), .Z(n1119) );
XNOR2_X1 U813 ( .A(n1120), .B(n1117), .ZN(n1118) );
NAND2_X1 U814 ( .A1(n1023), .A2(n1121), .ZN(n1108) );
NAND2_X1 U815 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR3_X1 U816 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(G66) );
NOR3_X1 U817 ( .A1(n1127), .A2(G953), .A3(G952), .ZN(n1126) );
AND2_X1 U818 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
INV_X1 U819 ( .A(KEYINPUT20), .ZN(n1127) );
XOR2_X1 U820 ( .A(n1129), .B(n1130), .Z(n1124) );
NAND3_X1 U821 ( .A1(n1131), .A2(n1066), .A3(n1132), .ZN(n1129) );
XOR2_X1 U822 ( .A(KEYINPUT2), .B(G217), .Z(n1131) );
NOR2_X1 U823 ( .A1(n1128), .A2(n1133), .ZN(G63) );
XOR2_X1 U824 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND3_X1 U825 ( .A1(G478), .A2(n1136), .A3(G902), .ZN(n1135) );
XNOR2_X1 U826 ( .A(KEYINPUT55), .B(n1014), .ZN(n1136) );
NOR2_X1 U827 ( .A1(n1128), .A2(n1137), .ZN(G60) );
NOR3_X1 U828 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1137) );
NOR2_X1 U829 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NOR2_X1 U830 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
INV_X1 U831 ( .A(KEYINPUT38), .ZN(n1144) );
XOR2_X1 U832 ( .A(KEYINPUT36), .B(n1145), .Z(n1143) );
AND3_X1 U833 ( .A1(n1141), .A2(n1145), .A3(KEYINPUT38), .ZN(n1139) );
NOR2_X1 U834 ( .A1(n1146), .A2(n1091), .ZN(n1141) );
NOR2_X1 U835 ( .A1(KEYINPUT38), .A2(n1145), .ZN(n1138) );
XNOR2_X1 U836 ( .A(G104), .B(n1147), .ZN(G6) );
NOR2_X1 U837 ( .A1(n1128), .A2(n1148), .ZN(G57) );
XOR2_X1 U838 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U839 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U840 ( .A(n1153), .B(KEYINPUT22), .Z(n1152) );
NAND2_X1 U841 ( .A1(n1132), .A2(G472), .ZN(n1151) );
XOR2_X1 U842 ( .A(n1154), .B(n1155), .Z(n1149) );
NOR2_X1 U843 ( .A1(G101), .A2(KEYINPUT50), .ZN(n1155) );
NOR2_X1 U844 ( .A1(n1128), .A2(n1156), .ZN(G54) );
NOR2_X1 U845 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XOR2_X1 U846 ( .A(n1159), .B(KEYINPUT5), .Z(n1158) );
NAND2_X1 U847 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR2_X1 U848 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
XNOR2_X1 U849 ( .A(n1162), .B(n1163), .ZN(n1161) );
AND2_X1 U850 ( .A1(n1132), .A2(G469), .ZN(n1160) );
INV_X1 U851 ( .A(n1146), .ZN(n1132) );
NOR2_X1 U852 ( .A1(n1164), .A2(n1165), .ZN(G51) );
XOR2_X1 U853 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U854 ( .A1(n1065), .A2(n1146), .ZN(n1167) );
NAND2_X1 U855 ( .A1(G902), .A2(n1014), .ZN(n1146) );
NAND3_X1 U856 ( .A1(n1122), .A2(n1168), .A3(n1100), .ZN(n1014) );
AND4_X1 U857 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1100) );
NOR4_X1 U858 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1172) );
NOR2_X1 U859 ( .A1(n1177), .A2(n1178), .ZN(n1171) );
NOR2_X1 U860 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XNOR2_X1 U861 ( .A(KEYINPUT60), .B(n1181), .ZN(n1180) );
NOR2_X1 U862 ( .A1(n1182), .A2(n1183), .ZN(n1177) );
XOR2_X1 U863 ( .A(KEYINPUT9), .B(n1184), .Z(n1183) );
XNOR2_X1 U864 ( .A(KEYINPUT16), .B(n1123), .ZN(n1168) );
AND4_X1 U865 ( .A1(n1185), .A2(n1186), .A3(n1147), .A4(n1187), .ZN(n1122) );
AND4_X1 U866 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187) );
NAND3_X1 U867 ( .A1(n1192), .A2(n1005), .A3(n1193), .ZN(n1147) );
NAND3_X1 U868 ( .A1(n1009), .A2(n1005), .A3(n1193), .ZN(n1186) );
NAND4_X1 U869 ( .A1(n1194), .A2(n1195), .A3(n1192), .A4(n1010), .ZN(n1185) );
XNOR2_X1 U870 ( .A(n1008), .B(KEYINPUT47), .ZN(n1194) );
NOR2_X1 U871 ( .A1(KEYINPUT1), .A2(n1196), .ZN(n1166) );
XOR2_X1 U872 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U873 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U874 ( .A1(KEYINPUT21), .A2(n1201), .ZN(n1199) );
XOR2_X1 U875 ( .A(n1202), .B(n1203), .Z(n1197) );
NOR3_X1 U876 ( .A1(n1204), .A2(KEYINPUT11), .A3(G953), .ZN(n1203) );
XOR2_X1 U877 ( .A(n1205), .B(KEYINPUT23), .Z(n1164) );
NAND2_X1 U878 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
OR3_X1 U879 ( .A1(n1016), .A2(n1023), .A3(KEYINPUT14), .ZN(n1207) );
INV_X1 U880 ( .A(G952), .ZN(n1016) );
NAND2_X1 U881 ( .A1(KEYINPUT14), .A2(n1128), .ZN(n1206) );
NOR2_X1 U882 ( .A1(n1023), .A2(G952), .ZN(n1128) );
XNOR2_X1 U883 ( .A(G146), .B(n1169), .ZN(G48) );
NAND3_X1 U884 ( .A1(n1192), .A2(n1008), .A3(n1208), .ZN(n1169) );
XNOR2_X1 U885 ( .A(G143), .B(n1170), .ZN(G45) );
NAND4_X1 U886 ( .A1(n1209), .A2(n1008), .A3(n1210), .A4(n1211), .ZN(n1170) );
XOR2_X1 U887 ( .A(G140), .B(n1173), .Z(G42) );
AND3_X1 U888 ( .A1(n1212), .A2(n1006), .A3(n1031), .ZN(n1173) );
XNOR2_X1 U889 ( .A(n1213), .B(n1176), .ZN(G39) );
AND3_X1 U890 ( .A1(n1208), .A2(n1031), .A3(n1027), .ZN(n1176) );
XOR2_X1 U891 ( .A(G134), .B(n1214), .Z(G36) );
NOR2_X1 U892 ( .A1(n1181), .A2(n1179), .ZN(n1214) );
NAND2_X1 U893 ( .A1(n1209), .A2(n1009), .ZN(n1179) );
INV_X1 U894 ( .A(n1031), .ZN(n1181) );
XOR2_X1 U895 ( .A(G131), .B(n1175), .Z(G33) );
AND3_X1 U896 ( .A1(n1031), .A2(n1192), .A3(n1209), .ZN(n1175) );
AND3_X1 U897 ( .A1(n1215), .A2(n1216), .A3(n1006), .ZN(n1209) );
NOR2_X1 U898 ( .A1(n1024), .A2(n1060), .ZN(n1031) );
INV_X1 U899 ( .A(n1025), .ZN(n1060) );
XNOR2_X1 U900 ( .A(G128), .B(n1217), .ZN(G30) );
NAND2_X1 U901 ( .A1(n1184), .A2(n1008), .ZN(n1217) );
AND2_X1 U902 ( .A1(n1208), .A2(n1009), .ZN(n1184) );
AND4_X1 U903 ( .A1(n1049), .A2(n1006), .A3(n1069), .A4(n1216), .ZN(n1208) );
XNOR2_X1 U904 ( .A(G101), .B(n1191), .ZN(G3) );
NAND3_X1 U905 ( .A1(n1027), .A2(n1215), .A3(n1193), .ZN(n1191) );
XOR2_X1 U906 ( .A(G125), .B(n1174), .Z(G27) );
AND3_X1 U907 ( .A1(n1212), .A2(n1008), .A3(n1051), .ZN(n1174) );
AND4_X1 U908 ( .A1(n1049), .A2(n1192), .A3(n1050), .A4(n1216), .ZN(n1212) );
NAND2_X1 U909 ( .A1(n1033), .A2(n1218), .ZN(n1216) );
NAND4_X1 U910 ( .A1(G953), .A2(G902), .A3(n1219), .A4(n1220), .ZN(n1218) );
INV_X1 U911 ( .A(G900), .ZN(n1220) );
INV_X1 U912 ( .A(n1037), .ZN(n1192) );
XNOR2_X1 U913 ( .A(G122), .B(n1190), .ZN(G24) );
NAND4_X1 U914 ( .A1(n1026), .A2(n1221), .A3(n1210), .A4(n1211), .ZN(n1190) );
AND2_X1 U915 ( .A1(n1051), .A2(n1005), .ZN(n1026) );
NAND2_X1 U916 ( .A1(n1222), .A2(n1223), .ZN(n1005) );
NAND2_X1 U917 ( .A1(n1215), .A2(n1224), .ZN(n1223) );
INV_X1 U918 ( .A(KEYINPUT62), .ZN(n1224) );
NAND3_X1 U919 ( .A1(n1225), .A2(n1050), .A3(KEYINPUT62), .ZN(n1222) );
XNOR2_X1 U920 ( .A(G119), .B(n1189), .ZN(G21) );
NAND3_X1 U921 ( .A1(n1221), .A2(n1027), .A3(n1226), .ZN(n1189) );
AND3_X1 U922 ( .A1(n1051), .A2(n1069), .A3(n1049), .ZN(n1226) );
XNOR2_X1 U923 ( .A(G116), .B(n1123), .ZN(G18) );
NAND3_X1 U924 ( .A1(n1221), .A2(n1009), .A3(n1195), .ZN(n1123) );
INV_X1 U925 ( .A(n1042), .ZN(n1195) );
NOR2_X1 U926 ( .A1(n1211), .A2(n1227), .ZN(n1009) );
INV_X1 U927 ( .A(n1228), .ZN(n1221) );
XNOR2_X1 U928 ( .A(n1229), .B(n1230), .ZN(G15) );
NOR4_X1 U929 ( .A1(KEYINPUT61), .A2(n1037), .A3(n1228), .A4(n1042), .ZN(n1230) );
NAND2_X1 U930 ( .A1(n1051), .A2(n1215), .ZN(n1042) );
AND2_X1 U931 ( .A1(n1225), .A2(n1069), .ZN(n1215) );
NOR2_X1 U932 ( .A1(n1231), .A2(n1047), .ZN(n1051) );
NAND2_X1 U933 ( .A1(n1227), .A2(n1211), .ZN(n1037) );
XNOR2_X1 U934 ( .A(n1232), .B(n1233), .ZN(G12) );
NOR2_X1 U935 ( .A1(KEYINPUT3), .A2(n1188), .ZN(n1233) );
NAND4_X1 U936 ( .A1(n1193), .A2(n1027), .A3(n1049), .A4(n1050), .ZN(n1188) );
INV_X1 U937 ( .A(n1069), .ZN(n1050) );
XNOR2_X1 U938 ( .A(n1234), .B(G472), .ZN(n1069) );
NAND2_X1 U939 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XOR2_X1 U940 ( .A(n1154), .B(n1237), .Z(n1235) );
XNOR2_X1 U941 ( .A(n1238), .B(n1153), .ZN(n1237) );
NAND3_X1 U942 ( .A1(n1239), .A2(n1023), .A3(G210), .ZN(n1153) );
XOR2_X1 U943 ( .A(n1240), .B(n1241), .Z(n1154) );
XOR2_X1 U944 ( .A(n1242), .B(n1243), .Z(n1241) );
XNOR2_X1 U945 ( .A(KEYINPUT30), .B(n1229), .ZN(n1243) );
XOR2_X1 U946 ( .A(n1244), .B(n1245), .Z(n1240) );
XNOR2_X1 U947 ( .A(n1246), .B(n1247), .ZN(n1245) );
XNOR2_X1 U948 ( .A(n1225), .B(KEYINPUT54), .ZN(n1049) );
NOR2_X1 U949 ( .A1(n1248), .A2(n1059), .ZN(n1225) );
NOR2_X1 U950 ( .A1(n1067), .A2(n1249), .ZN(n1059) );
AND2_X1 U951 ( .A1(G217), .A2(n1066), .ZN(n1249) );
AND3_X1 U952 ( .A1(G217), .A2(n1066), .A3(n1250), .ZN(n1248) );
XOR2_X1 U953 ( .A(n1067), .B(KEYINPUT24), .Z(n1250) );
NAND2_X1 U954 ( .A1(n1130), .A2(n1236), .ZN(n1067) );
XOR2_X1 U955 ( .A(n1251), .B(n1252), .Z(n1130) );
XNOR2_X1 U956 ( .A(n1213), .B(n1253), .ZN(n1252) );
AND3_X1 U957 ( .A1(n1254), .A2(G234), .A3(G221), .ZN(n1253) );
XNOR2_X1 U958 ( .A(KEYINPUT44), .B(G953), .ZN(n1254) );
INV_X1 U959 ( .A(G137), .ZN(n1213) );
NAND2_X1 U960 ( .A1(n1255), .A2(KEYINPUT28), .ZN(n1251) );
XOR2_X1 U961 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U962 ( .A(G119), .B(n1258), .Z(n1257) );
XOR2_X1 U963 ( .A(KEYINPUT41), .B(G146), .Z(n1258) );
XOR2_X1 U964 ( .A(n1259), .B(n1103), .Z(n1256) );
XNOR2_X1 U965 ( .A(G110), .B(n1260), .ZN(n1259) );
NOR2_X1 U966 ( .A1(KEYINPUT42), .A2(n1261), .ZN(n1260) );
INV_X1 U967 ( .A(G128), .ZN(n1261) );
NOR2_X1 U968 ( .A1(n1211), .A2(n1210), .ZN(n1027) );
INV_X1 U969 ( .A(n1227), .ZN(n1210) );
XNOR2_X1 U970 ( .A(n1073), .B(KEYINPUT7), .ZN(n1227) );
XOR2_X1 U971 ( .A(n1262), .B(G478), .Z(n1073) );
NAND2_X1 U972 ( .A1(n1236), .A2(n1134), .ZN(n1262) );
NAND2_X1 U973 ( .A1(n1263), .A2(n1264), .ZN(n1134) );
OR2_X1 U974 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
XOR2_X1 U975 ( .A(n1267), .B(KEYINPUT37), .Z(n1263) );
NAND2_X1 U976 ( .A1(n1266), .A2(n1265), .ZN(n1267) );
NAND3_X1 U977 ( .A1(G217), .A2(n1023), .A3(G234), .ZN(n1265) );
XNOR2_X1 U978 ( .A(n1268), .B(n1269), .ZN(n1266) );
XNOR2_X1 U979 ( .A(n1270), .B(n1271), .ZN(n1269) );
XNOR2_X1 U980 ( .A(G143), .B(n1272), .ZN(n1271) );
XNOR2_X1 U981 ( .A(G107), .B(n1273), .ZN(n1268) );
XNOR2_X1 U982 ( .A(n1090), .B(n1091), .ZN(n1211) );
INV_X1 U983 ( .A(G475), .ZN(n1091) );
NOR2_X1 U984 ( .A1(n1145), .A2(G902), .ZN(n1090) );
XNOR2_X1 U985 ( .A(n1274), .B(n1275), .ZN(n1145) );
XNOR2_X1 U986 ( .A(n1276), .B(n1277), .ZN(n1275) );
NAND2_X1 U987 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NAND2_X1 U988 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
XOR2_X1 U989 ( .A(KEYINPUT31), .B(n1282), .Z(n1280) );
NAND2_X1 U990 ( .A1(G104), .A2(n1283), .ZN(n1278) );
XNOR2_X1 U991 ( .A(n1282), .B(KEYINPUT48), .ZN(n1283) );
XNOR2_X1 U992 ( .A(G113), .B(n1272), .ZN(n1282) );
XNOR2_X1 U993 ( .A(n1284), .B(n1247), .ZN(n1274) );
XNOR2_X1 U994 ( .A(n1285), .B(n1286), .ZN(n1284) );
NOR2_X1 U995 ( .A1(KEYINPUT40), .A2(n1103), .ZN(n1286) );
XOR2_X1 U996 ( .A(G125), .B(G140), .Z(n1103) );
NOR4_X1 U997 ( .A1(KEYINPUT0), .A2(G953), .A3(G237), .A4(n1287), .ZN(n1285) );
INV_X1 U998 ( .A(G214), .ZN(n1287) );
NOR2_X1 U999 ( .A1(n1228), .A2(n1045), .ZN(n1193) );
INV_X1 U1000 ( .A(n1006), .ZN(n1045) );
NOR2_X1 U1001 ( .A1(n1048), .A2(n1047), .ZN(n1006) );
AND2_X1 U1002 ( .A1(G221), .A2(n1066), .ZN(n1047) );
NAND2_X1 U1003 ( .A1(G234), .A2(n1288), .ZN(n1066) );
XNOR2_X1 U1004 ( .A(KEYINPUT26), .B(n1236), .ZN(n1288) );
INV_X1 U1005 ( .A(n1231), .ZN(n1048) );
XNOR2_X1 U1006 ( .A(n1093), .B(G469), .ZN(n1231) );
NAND2_X1 U1007 ( .A1(n1289), .A2(n1236), .ZN(n1093) );
XOR2_X1 U1008 ( .A(n1162), .B(n1290), .Z(n1289) );
XNOR2_X1 U1009 ( .A(n1291), .B(KEYINPUT51), .ZN(n1290) );
NAND2_X1 U1010 ( .A1(KEYINPUT46), .A2(n1163), .ZN(n1291) );
XNOR2_X1 U1011 ( .A(n1292), .B(n1293), .ZN(n1163) );
XNOR2_X1 U1012 ( .A(G140), .B(n1232), .ZN(n1293) );
NAND2_X1 U1013 ( .A1(G227), .A2(n1023), .ZN(n1292) );
XOR2_X1 U1014 ( .A(n1294), .B(n1295), .Z(n1162) );
XOR2_X1 U1015 ( .A(n1296), .B(n1246), .Z(n1295) );
XOR2_X1 U1016 ( .A(KEYINPUT34), .B(KEYINPUT12), .Z(n1246) );
NOR2_X1 U1017 ( .A1(KEYINPUT17), .A2(n1238), .ZN(n1296) );
XOR2_X1 U1018 ( .A(n1102), .B(n1297), .Z(n1294) );
XOR2_X1 U1019 ( .A(n1244), .B(n1298), .Z(n1102) );
NOR2_X1 U1020 ( .A1(KEYINPUT29), .A2(n1247), .ZN(n1298) );
XOR2_X1 U1021 ( .A(n1299), .B(n1273), .Z(n1244) );
XOR2_X1 U1022 ( .A(G134), .B(G128), .Z(n1273) );
XNOR2_X1 U1023 ( .A(G137), .B(n1276), .ZN(n1299) );
XOR2_X1 U1024 ( .A(G131), .B(KEYINPUT45), .Z(n1276) );
NAND2_X1 U1025 ( .A1(n1008), .A2(n1010), .ZN(n1228) );
NAND2_X1 U1026 ( .A1(n1033), .A2(n1300), .ZN(n1010) );
NAND3_X1 U1027 ( .A1(G902), .A2(n1219), .A3(n1110), .ZN(n1300) );
NOR2_X1 U1028 ( .A1(n1023), .A2(G898), .ZN(n1110) );
NAND3_X1 U1029 ( .A1(n1219), .A2(n1023), .A3(G952), .ZN(n1033) );
INV_X1 U1030 ( .A(G953), .ZN(n1023) );
NAND2_X1 U1031 ( .A1(G237), .A2(G234), .ZN(n1219) );
INV_X1 U1032 ( .A(n1182), .ZN(n1008) );
NAND2_X1 U1033 ( .A1(n1024), .A2(n1025), .ZN(n1182) );
NAND2_X1 U1034 ( .A1(G214), .A2(n1301), .ZN(n1025) );
XNOR2_X1 U1035 ( .A(n1064), .B(n1065), .ZN(n1024) );
NAND2_X1 U1036 ( .A1(G210), .A2(n1301), .ZN(n1065) );
NAND2_X1 U1037 ( .A1(n1239), .A2(n1236), .ZN(n1301) );
INV_X1 U1038 ( .A(G237), .ZN(n1239) );
AND2_X1 U1039 ( .A1(n1302), .A2(n1236), .ZN(n1064) );
INV_X1 U1040 ( .A(G902), .ZN(n1236) );
XNOR2_X1 U1041 ( .A(n1303), .B(n1202), .ZN(n1302) );
NAND2_X1 U1042 ( .A1(n1304), .A2(n1305), .ZN(n1202) );
NAND2_X1 U1043 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XNOR2_X1 U1044 ( .A(KEYINPUT58), .B(n1120), .ZN(n1307) );
INV_X1 U1045 ( .A(n1116), .ZN(n1120) );
NAND2_X1 U1046 ( .A1(n1308), .A2(n1309), .ZN(n1304) );
XNOR2_X1 U1047 ( .A(n1310), .B(n1306), .ZN(n1309) );
XNOR2_X1 U1048 ( .A(n1115), .B(n1117), .ZN(n1306) );
XNOR2_X1 U1049 ( .A(n1229), .B(n1311), .ZN(n1117) );
NOR3_X1 U1050 ( .A1(KEYINPUT10), .A2(n1312), .A3(n1313), .ZN(n1311) );
NOR3_X1 U1051 ( .A1(n1314), .A2(G119), .A3(n1270), .ZN(n1313) );
INV_X1 U1052 ( .A(KEYINPUT57), .ZN(n1314) );
NOR2_X1 U1053 ( .A1(KEYINPUT57), .A2(n1242), .ZN(n1312) );
XNOR2_X1 U1054 ( .A(n1270), .B(G119), .ZN(n1242) );
INV_X1 U1055 ( .A(G116), .ZN(n1270) );
INV_X1 U1056 ( .A(G113), .ZN(n1229) );
XNOR2_X1 U1057 ( .A(G110), .B(n1272), .ZN(n1115) );
INV_X1 U1058 ( .A(G122), .ZN(n1272) );
XNOR2_X1 U1059 ( .A(KEYINPUT32), .B(KEYINPUT27), .ZN(n1310) );
XNOR2_X1 U1060 ( .A(KEYINPUT58), .B(n1116), .ZN(n1308) );
XOR2_X1 U1061 ( .A(n1315), .B(n1238), .Z(n1116) );
INV_X1 U1062 ( .A(G101), .ZN(n1238) );
NAND2_X1 U1063 ( .A1(KEYINPUT59), .A2(n1297), .ZN(n1315) );
XNOR2_X1 U1064 ( .A(G107), .B(n1281), .ZN(n1297) );
INV_X1 U1065 ( .A(G104), .ZN(n1281) );
NAND2_X1 U1066 ( .A1(n1316), .A2(KEYINPUT6), .ZN(n1303) );
XOR2_X1 U1067 ( .A(n1317), .B(n1200), .Z(n1316) );
XOR2_X1 U1068 ( .A(G125), .B(KEYINPUT19), .Z(n1200) );
XNOR2_X1 U1069 ( .A(n1201), .B(n1318), .ZN(n1317) );
NOR2_X1 U1070 ( .A1(G953), .A2(n1204), .ZN(n1318) );
INV_X1 U1071 ( .A(G224), .ZN(n1204) );
XNOR2_X1 U1072 ( .A(G128), .B(n1247), .ZN(n1201) );
XNOR2_X1 U1073 ( .A(G143), .B(G146), .ZN(n1247) );
INV_X1 U1074 ( .A(G110), .ZN(n1232) );
endmodule


