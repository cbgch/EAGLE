//Key = 0101011011111100101111101011001111011110100010111100000111010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395;

XNOR2_X1 U753 ( .A(G107), .B(n1058), .ZN(G9) );
NOR2_X1 U754 ( .A1(n1059), .A2(n1060), .ZN(G75) );
NOR4_X1 U755 ( .A1(G953), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1060) );
NOR2_X1 U756 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U757 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U758 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
INV_X1 U759 ( .A(n1070), .ZN(n1069) );
NOR2_X1 U760 ( .A1(n1071), .A2(n1072), .ZN(n1068) );
NOR2_X1 U761 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U762 ( .A1(n1075), .A2(n1076), .ZN(n1071) );
NOR2_X1 U763 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NOR2_X1 U764 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U765 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NOR3_X1 U766 ( .A1(n1083), .A2(n1073), .A3(n1084), .ZN(n1077) );
INV_X1 U767 ( .A(n1085), .ZN(n1084) );
AND3_X1 U768 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1073) );
NAND2_X1 U769 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
OR2_X1 U770 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U771 ( .A1(n1093), .A2(n1094), .ZN(n1086) );
NAND2_X1 U772 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U773 ( .A1(n1085), .A2(n1083), .ZN(n1096) );
NAND2_X1 U774 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
INV_X1 U775 ( .A(KEYINPUT28), .ZN(n1083) );
NOR4_X1 U776 ( .A1(n1099), .A2(n1074), .A3(n1076), .A4(n1080), .ZN(n1066) );
NOR2_X1 U777 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U778 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR3_X1 U779 ( .A1(n1061), .A2(G953), .A3(G952), .ZN(n1059) );
AND4_X1 U780 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1061) );
NOR4_X1 U781 ( .A1(n1108), .A2(n1109), .A3(n1097), .A4(n1110), .ZN(n1107) );
NOR2_X1 U782 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U783 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U784 ( .A1(n1115), .A2(KEYINPUT23), .ZN(n1113) );
NOR2_X1 U785 ( .A1(n1116), .A2(n1117), .ZN(n1111) );
XNOR2_X1 U786 ( .A(n1115), .B(KEYINPUT16), .ZN(n1117) );
NOR2_X1 U787 ( .A1(n1118), .A2(n1115), .ZN(n1116) );
NOR2_X1 U788 ( .A1(KEYINPUT23), .A2(G478), .ZN(n1118) );
NOR2_X1 U789 ( .A1(n1119), .A2(n1120), .ZN(n1108) );
NOR2_X1 U790 ( .A1(G469), .A2(n1121), .ZN(n1120) );
XNOR2_X1 U791 ( .A(KEYINPUT52), .B(n1122), .ZN(n1121) );
NOR2_X1 U792 ( .A1(n1123), .A2(n1124), .ZN(n1106) );
XNOR2_X1 U793 ( .A(n1125), .B(n1126), .ZN(n1124) );
NAND2_X1 U794 ( .A1(KEYINPUT12), .A2(n1127), .ZN(n1125) );
XNOR2_X1 U795 ( .A(n1102), .B(KEYINPUT6), .ZN(n1123) );
XOR2_X1 U796 ( .A(n1128), .B(n1129), .Z(n1105) );
XNOR2_X1 U797 ( .A(n1130), .B(KEYINPUT42), .ZN(n1128) );
XNOR2_X1 U798 ( .A(n1131), .B(n1132), .ZN(n1104) );
NAND2_X1 U799 ( .A1(n1133), .A2(n1134), .ZN(G72) );
NAND2_X1 U800 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U801 ( .A1(G953), .A2(n1137), .ZN(n1135) );
NAND2_X1 U802 ( .A1(G900), .A2(G227), .ZN(n1137) );
NAND2_X1 U803 ( .A1(n1138), .A2(n1139), .ZN(n1133) );
NAND2_X1 U804 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U805 ( .A1(G953), .A2(n1142), .ZN(n1141) );
INV_X1 U806 ( .A(n1143), .ZN(n1140) );
INV_X1 U807 ( .A(n1136), .ZN(n1138) );
NAND2_X1 U808 ( .A1(n1144), .A2(n1145), .ZN(n1136) );
NAND2_X1 U809 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U810 ( .A(KEYINPUT30), .B(n1148), .Z(n1144) );
NOR3_X1 U811 ( .A1(n1147), .A2(n1146), .A3(n1143), .ZN(n1148) );
AND2_X1 U812 ( .A1(n1149), .A2(n1150), .ZN(n1146) );
XOR2_X1 U813 ( .A(n1151), .B(n1152), .Z(n1147) );
NAND2_X1 U814 ( .A1(n1153), .A2(n1154), .ZN(G69) );
NAND2_X1 U815 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND2_X1 U816 ( .A1(G953), .A2(n1157), .ZN(n1155) );
NAND3_X1 U817 ( .A1(G953), .A2(n1158), .A3(n1159), .ZN(n1153) );
XOR2_X1 U818 ( .A(n1156), .B(KEYINPUT5), .Z(n1159) );
NAND2_X1 U819 ( .A1(n1160), .A2(n1161), .ZN(n1156) );
NAND4_X1 U820 ( .A1(n1162), .A2(n1150), .A3(n1163), .A4(n1164), .ZN(n1161) );
NAND2_X1 U821 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NAND2_X1 U822 ( .A1(KEYINPUT53), .A2(n1167), .ZN(n1163) );
NAND3_X1 U823 ( .A1(n1168), .A2(n1166), .A3(n1165), .ZN(n1160) );
INV_X1 U824 ( .A(n1167), .ZN(n1165) );
NAND2_X1 U825 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
NAND2_X1 U826 ( .A1(G953), .A2(n1171), .ZN(n1170) );
XOR2_X1 U827 ( .A(n1172), .B(n1173), .Z(n1169) );
INV_X1 U828 ( .A(KEYINPUT39), .ZN(n1166) );
NAND2_X1 U829 ( .A1(n1174), .A2(n1162), .ZN(n1168) );
INV_X1 U830 ( .A(KEYINPUT53), .ZN(n1174) );
NAND2_X1 U831 ( .A1(G898), .A2(G224), .ZN(n1158) );
NOR2_X1 U832 ( .A1(n1175), .A2(n1176), .ZN(G66) );
NOR3_X1 U833 ( .A1(n1130), .A2(n1177), .A3(n1178), .ZN(n1176) );
NOR4_X1 U834 ( .A1(n1179), .A2(n1180), .A3(KEYINPUT15), .A4(n1181), .ZN(n1178) );
NOR2_X1 U835 ( .A1(n1182), .A2(n1183), .ZN(n1177) );
NOR3_X1 U836 ( .A1(n1181), .A2(KEYINPUT15), .A3(n1184), .ZN(n1182) );
NOR2_X1 U837 ( .A1(n1175), .A2(n1185), .ZN(G63) );
NOR3_X1 U838 ( .A1(n1115), .A2(n1186), .A3(n1187), .ZN(n1185) );
NOR3_X1 U839 ( .A1(n1188), .A2(n1114), .A3(n1180), .ZN(n1187) );
NOR2_X1 U840 ( .A1(n1189), .A2(n1190), .ZN(n1186) );
NOR2_X1 U841 ( .A1(n1184), .A2(n1114), .ZN(n1189) );
NOR2_X1 U842 ( .A1(n1175), .A2(n1191), .ZN(G60) );
XOR2_X1 U843 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U844 ( .A(KEYINPUT59), .B(n1194), .Z(n1193) );
NOR2_X1 U845 ( .A1(n1126), .A2(n1180), .ZN(n1194) );
XNOR2_X1 U846 ( .A(n1195), .B(n1196), .ZN(G6) );
NOR2_X1 U847 ( .A1(n1175), .A2(n1197), .ZN(G57) );
XNOR2_X1 U848 ( .A(n1198), .B(n1199), .ZN(n1197) );
XOR2_X1 U849 ( .A(G101), .B(n1200), .Z(n1199) );
NOR2_X1 U850 ( .A1(KEYINPUT4), .A2(n1201), .ZN(n1200) );
XNOR2_X1 U851 ( .A(n1152), .B(n1202), .ZN(n1201) );
XOR2_X1 U852 ( .A(n1203), .B(n1204), .Z(n1202) );
NOR2_X1 U853 ( .A1(n1132), .A2(n1180), .ZN(n1204) );
NOR2_X1 U854 ( .A1(n1175), .A2(n1205), .ZN(G54) );
XOR2_X1 U855 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U856 ( .A(n1152), .B(n1208), .Z(n1207) );
XOR2_X1 U857 ( .A(n1209), .B(n1210), .Z(n1208) );
NOR2_X1 U858 ( .A1(KEYINPUT54), .A2(n1211), .ZN(n1210) );
NOR2_X1 U859 ( .A1(n1212), .A2(n1180), .ZN(n1209) );
XNOR2_X1 U860 ( .A(n1213), .B(n1214), .ZN(n1152) );
XOR2_X1 U861 ( .A(n1215), .B(n1216), .Z(n1206) );
XOR2_X1 U862 ( .A(n1217), .B(n1218), .Z(n1216) );
NOR2_X1 U863 ( .A1(KEYINPUT60), .A2(n1219), .ZN(n1218) );
XOR2_X1 U864 ( .A(KEYINPUT0), .B(G110), .Z(n1215) );
NOR2_X1 U865 ( .A1(n1175), .A2(n1220), .ZN(G51) );
XOR2_X1 U866 ( .A(n1221), .B(n1222), .Z(n1220) );
XOR2_X1 U867 ( .A(n1223), .B(n1224), .Z(n1222) );
XNOR2_X1 U868 ( .A(n1225), .B(n1226), .ZN(n1221) );
NOR2_X1 U869 ( .A1(n1227), .A2(n1180), .ZN(n1226) );
NAND2_X1 U870 ( .A1(G902), .A2(n1063), .ZN(n1180) );
INV_X1 U871 ( .A(n1184), .ZN(n1063) );
NOR2_X1 U872 ( .A1(n1162), .A2(n1149), .ZN(n1184) );
NAND4_X1 U873 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1149) );
NOR4_X1 U874 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1231) );
NOR2_X1 U875 ( .A1(n1236), .A2(n1237), .ZN(n1230) );
NAND2_X1 U876 ( .A1(n1070), .A2(n1238), .ZN(n1228) );
XOR2_X1 U877 ( .A(KEYINPUT58), .B(n1239), .Z(n1238) );
NAND4_X1 U878 ( .A1(n1240), .A2(n1058), .A3(n1241), .A4(n1242), .ZN(n1162) );
NOR4_X1 U879 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1242) );
NOR2_X1 U880 ( .A1(KEYINPUT34), .A2(n1247), .ZN(n1246) );
NOR2_X1 U881 ( .A1(n1248), .A2(n1249), .ZN(n1245) );
NOR2_X1 U882 ( .A1(n1250), .A2(n1251), .ZN(n1248) );
AND2_X1 U883 ( .A1(n1081), .A2(n1091), .ZN(n1251) );
NOR3_X1 U884 ( .A1(n1252), .A2(n1253), .A3(n1074), .ZN(n1250) );
INV_X1 U885 ( .A(n1088), .ZN(n1074) );
INV_X1 U886 ( .A(KEYINPUT34), .ZN(n1252) );
NOR2_X1 U887 ( .A1(n1254), .A2(n1196), .ZN(n1241) );
AND3_X1 U888 ( .A1(n1255), .A2(n1088), .A3(n1091), .ZN(n1196) );
NAND3_X1 U889 ( .A1(n1092), .A2(n1088), .A3(n1255), .ZN(n1058) );
NOR2_X1 U890 ( .A1(n1150), .A2(G952), .ZN(n1175) );
XOR2_X1 U891 ( .A(G146), .B(n1232), .Z(G48) );
AND3_X1 U892 ( .A1(n1091), .A2(n1101), .A3(n1256), .ZN(n1232) );
XNOR2_X1 U893 ( .A(G143), .B(n1229), .ZN(G45) );
NAND3_X1 U894 ( .A1(n1253), .A2(n1101), .A3(n1257), .ZN(n1229) );
XNOR2_X1 U895 ( .A(n1211), .B(n1237), .ZN(G42) );
AND3_X1 U896 ( .A1(n1258), .A2(n1085), .A3(n1070), .ZN(n1237) );
XOR2_X1 U897 ( .A(G137), .B(n1236), .Z(G39) );
AND3_X1 U898 ( .A1(n1256), .A2(n1093), .A3(n1070), .ZN(n1236) );
XOR2_X1 U899 ( .A(G134), .B(n1235), .Z(G36) );
AND3_X1 U900 ( .A1(n1070), .A2(n1092), .A3(n1257), .ZN(n1235) );
XNOR2_X1 U901 ( .A(G131), .B(n1259), .ZN(G33) );
NAND2_X1 U902 ( .A1(n1239), .A2(n1070), .ZN(n1259) );
NOR2_X1 U903 ( .A1(n1102), .A2(n1109), .ZN(n1070) );
AND2_X1 U904 ( .A1(n1257), .A2(n1091), .ZN(n1239) );
AND3_X1 U905 ( .A1(n1085), .A2(n1260), .A3(n1081), .ZN(n1257) );
NAND2_X1 U906 ( .A1(n1261), .A2(n1262), .ZN(G30) );
NAND2_X1 U907 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
NAND2_X1 U908 ( .A1(n1265), .A2(n1266), .ZN(n1263) );
OR2_X1 U909 ( .A1(n1234), .A2(KEYINPUT17), .ZN(n1266) );
NAND2_X1 U910 ( .A1(n1234), .A2(n1267), .ZN(n1265) );
OR2_X1 U911 ( .A1(KEYINPUT14), .A2(KEYINPUT17), .ZN(n1267) );
INV_X1 U912 ( .A(n1268), .ZN(n1234) );
OR3_X1 U913 ( .A1(n1268), .A2(KEYINPUT14), .A3(n1264), .ZN(n1261) );
XNOR2_X1 U914 ( .A(G128), .B(KEYINPUT27), .ZN(n1264) );
NAND3_X1 U915 ( .A1(n1092), .A2(n1101), .A3(n1256), .ZN(n1268) );
AND4_X1 U916 ( .A1(n1269), .A2(n1085), .A3(n1270), .A4(n1260), .ZN(n1256) );
XOR2_X1 U917 ( .A(G101), .B(n1254), .Z(G3) );
AND3_X1 U918 ( .A1(n1093), .A2(n1255), .A3(n1081), .ZN(n1254) );
XOR2_X1 U919 ( .A(G125), .B(n1233), .Z(G27) );
AND3_X1 U920 ( .A1(n1089), .A2(n1101), .A3(n1258), .ZN(n1233) );
AND3_X1 U921 ( .A1(n1091), .A2(n1260), .A3(n1082), .ZN(n1258) );
NAND2_X1 U922 ( .A1(n1065), .A2(n1271), .ZN(n1260) );
NAND3_X1 U923 ( .A1(G902), .A2(n1272), .A3(n1143), .ZN(n1271) );
NOR2_X1 U924 ( .A1(n1150), .A2(G900), .ZN(n1143) );
XNOR2_X1 U925 ( .A(G122), .B(n1247), .ZN(G24) );
NAND3_X1 U926 ( .A1(n1273), .A2(n1088), .A3(n1253), .ZN(n1247) );
NOR2_X1 U927 ( .A1(n1274), .A2(n1275), .ZN(n1253) );
NOR2_X1 U928 ( .A1(n1270), .A2(n1269), .ZN(n1088) );
XOR2_X1 U929 ( .A(G119), .B(n1244), .Z(G21) );
AND4_X1 U930 ( .A1(n1273), .A2(n1093), .A3(n1269), .A4(n1270), .ZN(n1244) );
INV_X1 U931 ( .A(n1276), .ZN(n1269) );
XOR2_X1 U932 ( .A(G116), .B(n1243), .Z(G18) );
AND3_X1 U933 ( .A1(n1081), .A2(n1092), .A3(n1273), .ZN(n1243) );
AND2_X1 U934 ( .A1(n1274), .A2(n1277), .ZN(n1092) );
XNOR2_X1 U935 ( .A(n1278), .B(n1279), .ZN(G15) );
NAND2_X1 U936 ( .A1(n1280), .A2(n1281), .ZN(n1278) );
NAND3_X1 U937 ( .A1(n1101), .A2(n1282), .A3(n1283), .ZN(n1281) );
INV_X1 U938 ( .A(KEYINPUT24), .ZN(n1283) );
NAND4_X1 U939 ( .A1(n1284), .A2(n1089), .A3(n1081), .A4(n1285), .ZN(n1282) );
NAND4_X1 U940 ( .A1(n1284), .A2(n1081), .A3(n1273), .A4(KEYINPUT24), .ZN(n1280) );
INV_X1 U941 ( .A(n1249), .ZN(n1273) );
NAND3_X1 U942 ( .A1(n1101), .A2(n1285), .A3(n1089), .ZN(n1249) );
INV_X1 U943 ( .A(n1080), .ZN(n1089) );
NAND2_X1 U944 ( .A1(n1286), .A2(n1098), .ZN(n1080) );
INV_X1 U945 ( .A(n1287), .ZN(n1286) );
NOR2_X1 U946 ( .A1(n1276), .A2(n1270), .ZN(n1081) );
XNOR2_X1 U947 ( .A(n1091), .B(KEYINPUT26), .ZN(n1284) );
NOR2_X1 U948 ( .A1(n1274), .A2(n1277), .ZN(n1091) );
INV_X1 U949 ( .A(n1275), .ZN(n1277) );
NAND2_X1 U950 ( .A1(n1288), .A2(n1289), .ZN(G12) );
NAND2_X1 U951 ( .A1(G110), .A2(n1240), .ZN(n1289) );
XOR2_X1 U952 ( .A(n1290), .B(KEYINPUT45), .Z(n1288) );
OR2_X1 U953 ( .A1(n1240), .A2(G110), .ZN(n1290) );
NAND3_X1 U954 ( .A1(n1093), .A2(n1255), .A3(n1082), .ZN(n1240) );
AND2_X1 U955 ( .A1(n1291), .A2(n1270), .ZN(n1082) );
XNOR2_X1 U956 ( .A(n1292), .B(n1293), .ZN(n1270) );
XOR2_X1 U957 ( .A(KEYINPUT62), .B(n1129), .Z(n1293) );
AND2_X1 U958 ( .A1(G217), .A2(n1294), .ZN(n1129) );
NAND2_X1 U959 ( .A1(KEYINPUT33), .A2(n1295), .ZN(n1292) );
INV_X1 U960 ( .A(n1130), .ZN(n1295) );
NOR2_X1 U961 ( .A1(n1183), .A2(G902), .ZN(n1130) );
INV_X1 U962 ( .A(n1179), .ZN(n1183) );
XNOR2_X1 U963 ( .A(n1296), .B(n1297), .ZN(n1179) );
XOR2_X1 U964 ( .A(n1298), .B(n1299), .Z(n1297) );
XOR2_X1 U965 ( .A(G137), .B(G128), .Z(n1299) );
XOR2_X1 U966 ( .A(KEYINPUT51), .B(G146), .Z(n1298) );
XOR2_X1 U967 ( .A(n1300), .B(n1301), .Z(n1296) );
XOR2_X1 U968 ( .A(n1302), .B(n1151), .Z(n1301) );
AND3_X1 U969 ( .A1(G221), .A2(n1150), .A3(G234), .ZN(n1302) );
XNOR2_X1 U970 ( .A(G119), .B(G110), .ZN(n1300) );
XNOR2_X1 U971 ( .A(KEYINPUT31), .B(n1276), .ZN(n1291) );
NAND3_X1 U972 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(n1276) );
NAND2_X1 U973 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U974 ( .A1(n1308), .A2(n1131), .ZN(n1307) );
XNOR2_X1 U975 ( .A(KEYINPUT41), .B(n1132), .ZN(n1306) );
INV_X1 U976 ( .A(G472), .ZN(n1132) );
OR2_X1 U977 ( .A1(n1131), .A2(KEYINPUT19), .ZN(n1304) );
NAND4_X1 U978 ( .A1(n1309), .A2(n1131), .A3(n1308), .A4(KEYINPUT19), .ZN(n1303) );
XOR2_X1 U979 ( .A(KEYINPUT50), .B(KEYINPUT21), .Z(n1308) );
NAND2_X1 U980 ( .A1(n1310), .A2(n1311), .ZN(n1131) );
XOR2_X1 U981 ( .A(n1312), .B(n1313), .Z(n1310) );
XOR2_X1 U982 ( .A(G101), .B(n1314), .Z(n1313) );
NOR2_X1 U983 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XOR2_X1 U984 ( .A(n1317), .B(KEYINPUT44), .Z(n1316) );
NAND2_X1 U985 ( .A1(n1318), .A2(n1203), .ZN(n1317) );
XNOR2_X1 U986 ( .A(n1319), .B(KEYINPUT56), .ZN(n1318) );
NOR2_X1 U987 ( .A1(n1203), .A2(n1319), .ZN(n1315) );
XOR2_X1 U988 ( .A(n1320), .B(n1321), .Z(n1319) );
NAND2_X1 U989 ( .A1(KEYINPUT40), .A2(n1214), .ZN(n1320) );
AND2_X1 U990 ( .A1(n1322), .A2(n1323), .ZN(n1203) );
NAND2_X1 U991 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
NAND2_X1 U992 ( .A1(KEYINPUT1), .A2(n1326), .ZN(n1325) );
NAND2_X1 U993 ( .A1(KEYINPUT46), .A2(n1279), .ZN(n1326) );
INV_X1 U994 ( .A(n1327), .ZN(n1324) );
NAND2_X1 U995 ( .A1(G113), .A2(n1328), .ZN(n1322) );
NAND2_X1 U996 ( .A1(KEYINPUT46), .A2(n1329), .ZN(n1328) );
NAND2_X1 U997 ( .A1(KEYINPUT1), .A2(n1327), .ZN(n1329) );
NOR2_X1 U998 ( .A1(KEYINPUT7), .A2(n1198), .ZN(n1312) );
NAND3_X1 U999 ( .A1(n1330), .A2(n1150), .A3(G210), .ZN(n1198) );
XNOR2_X1 U1000 ( .A(KEYINPUT41), .B(G472), .ZN(n1309) );
AND3_X1 U1001 ( .A1(n1085), .A2(n1285), .A3(n1101), .ZN(n1255) );
NOR2_X1 U1002 ( .A1(n1331), .A2(n1109), .ZN(n1101) );
INV_X1 U1003 ( .A(n1103), .ZN(n1109) );
NAND2_X1 U1004 ( .A1(G214), .A2(n1332), .ZN(n1103) );
INV_X1 U1005 ( .A(n1102), .ZN(n1331) );
XOR2_X1 U1006 ( .A(n1333), .B(n1227), .Z(n1102) );
NAND2_X1 U1007 ( .A1(G210), .A2(n1332), .ZN(n1227) );
NAND2_X1 U1008 ( .A1(n1334), .A2(n1311), .ZN(n1332) );
XNOR2_X1 U1009 ( .A(G237), .B(KEYINPUT29), .ZN(n1334) );
NAND2_X1 U1010 ( .A1(n1335), .A2(n1311), .ZN(n1333) );
XOR2_X1 U1011 ( .A(n1223), .B(n1336), .Z(n1335) );
XNOR2_X1 U1012 ( .A(n1337), .B(KEYINPUT48), .ZN(n1336) );
NAND3_X1 U1013 ( .A1(n1338), .A2(n1339), .A3(KEYINPUT9), .ZN(n1337) );
NAND2_X1 U1014 ( .A1(n1340), .A2(n1214), .ZN(n1339) );
XNOR2_X1 U1015 ( .A(n1224), .B(KEYINPUT35), .ZN(n1340) );
NAND2_X1 U1016 ( .A1(n1225), .A2(n1341), .ZN(n1338) );
XNOR2_X1 U1017 ( .A(n1224), .B(KEYINPUT2), .ZN(n1341) );
XOR2_X1 U1018 ( .A(G125), .B(n1342), .Z(n1224) );
NOR2_X1 U1019 ( .A1(G953), .A2(n1157), .ZN(n1342) );
INV_X1 U1020 ( .A(G224), .ZN(n1157) );
XOR2_X1 U1021 ( .A(n1343), .B(n1172), .Z(n1223) );
XNOR2_X1 U1022 ( .A(n1344), .B(n1345), .ZN(n1172) );
XOR2_X1 U1023 ( .A(n1346), .B(n1347), .Z(n1345) );
NAND2_X1 U1024 ( .A1(KEYINPUT8), .A2(G101), .ZN(n1347) );
NAND2_X1 U1025 ( .A1(n1348), .A2(n1349), .ZN(n1346) );
NAND2_X1 U1026 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
XOR2_X1 U1027 ( .A(KEYINPUT11), .B(n1352), .Z(n1350) );
XOR2_X1 U1028 ( .A(KEYINPUT38), .B(n1353), .Z(n1348) );
AND2_X1 U1029 ( .A1(n1352), .A2(G107), .ZN(n1353) );
XOR2_X1 U1030 ( .A(G104), .B(KEYINPUT57), .Z(n1352) );
XNOR2_X1 U1031 ( .A(G122), .B(G110), .ZN(n1344) );
NAND2_X1 U1032 ( .A1(KEYINPUT37), .A2(n1173), .ZN(n1343) );
XNOR2_X1 U1033 ( .A(n1354), .B(n1279), .ZN(n1173) );
NAND2_X1 U1034 ( .A1(KEYINPUT49), .A2(n1327), .ZN(n1354) );
XNOR2_X1 U1035 ( .A(G119), .B(G116), .ZN(n1327) );
NAND2_X1 U1036 ( .A1(n1065), .A2(n1355), .ZN(n1285) );
NAND4_X1 U1037 ( .A1(G953), .A2(G902), .A3(n1272), .A4(n1171), .ZN(n1355) );
INV_X1 U1038 ( .A(G898), .ZN(n1171) );
NAND3_X1 U1039 ( .A1(n1272), .A2(n1150), .A3(G952), .ZN(n1065) );
NAND2_X1 U1040 ( .A1(G234), .A2(G237), .ZN(n1272) );
NOR2_X1 U1041 ( .A1(n1098), .A2(n1287), .ZN(n1085) );
XNOR2_X1 U1042 ( .A(n1097), .B(KEYINPUT20), .ZN(n1287) );
AND2_X1 U1043 ( .A1(G221), .A2(n1294), .ZN(n1097) );
NAND2_X1 U1044 ( .A1(G234), .A2(n1311), .ZN(n1294) );
NAND3_X1 U1045 ( .A1(n1356), .A2(n1357), .A3(n1358), .ZN(n1098) );
INV_X1 U1046 ( .A(n1119), .ZN(n1358) );
NOR2_X1 U1047 ( .A1(n1212), .A2(n1122), .ZN(n1119) );
NAND3_X1 U1048 ( .A1(KEYINPUT63), .A2(n1122), .A3(n1212), .ZN(n1357) );
NAND2_X1 U1049 ( .A1(n1359), .A2(n1311), .ZN(n1122) );
XOR2_X1 U1050 ( .A(n1360), .B(n1361), .Z(n1359) );
XNOR2_X1 U1051 ( .A(n1321), .B(n1219), .ZN(n1361) );
XOR2_X1 U1052 ( .A(G101), .B(n1362), .Z(n1219) );
XNOR2_X1 U1053 ( .A(n1351), .B(G104), .ZN(n1362) );
INV_X1 U1054 ( .A(n1213), .ZN(n1321) );
XOR2_X1 U1055 ( .A(G131), .B(n1363), .Z(n1213) );
XOR2_X1 U1056 ( .A(G137), .B(G134), .Z(n1363) );
XOR2_X1 U1057 ( .A(n1364), .B(n1365), .Z(n1360) );
XNOR2_X1 U1058 ( .A(n1217), .B(n1366), .ZN(n1365) );
NAND2_X1 U1059 ( .A1(KEYINPUT32), .A2(n1367), .ZN(n1366) );
XNOR2_X1 U1060 ( .A(n1211), .B(G110), .ZN(n1367) );
NOR2_X1 U1061 ( .A1(n1142), .A2(G953), .ZN(n1217) );
INV_X1 U1062 ( .A(G227), .ZN(n1142) );
NAND2_X1 U1063 ( .A1(KEYINPUT55), .A2(n1368), .ZN(n1364) );
XNOR2_X1 U1064 ( .A(KEYINPUT13), .B(n1214), .ZN(n1368) );
INV_X1 U1065 ( .A(n1225), .ZN(n1214) );
XOR2_X1 U1066 ( .A(G146), .B(n1369), .Z(n1225) );
OR2_X1 U1067 ( .A1(n1212), .A2(KEYINPUT63), .ZN(n1356) );
INV_X1 U1068 ( .A(G469), .ZN(n1212) );
INV_X1 U1069 ( .A(n1076), .ZN(n1093) );
NAND2_X1 U1070 ( .A1(n1275), .A2(n1274), .ZN(n1076) );
XNOR2_X1 U1071 ( .A(n1127), .B(n1370), .ZN(n1274) );
XNOR2_X1 U1072 ( .A(KEYINPUT10), .B(n1126), .ZN(n1370) );
INV_X1 U1073 ( .A(G475), .ZN(n1126) );
NAND2_X1 U1074 ( .A1(n1192), .A2(n1311), .ZN(n1127) );
INV_X1 U1075 ( .A(G902), .ZN(n1311) );
XNOR2_X1 U1076 ( .A(n1371), .B(n1372), .ZN(n1192) );
XOR2_X1 U1077 ( .A(n1373), .B(n1374), .Z(n1372) );
XNOR2_X1 U1078 ( .A(n1375), .B(n1376), .ZN(n1374) );
NOR2_X1 U1079 ( .A1(KEYINPUT43), .A2(n1377), .ZN(n1376) );
XNOR2_X1 U1080 ( .A(n1195), .B(n1378), .ZN(n1377) );
XNOR2_X1 U1081 ( .A(G122), .B(n1279), .ZN(n1378) );
INV_X1 U1082 ( .A(G113), .ZN(n1279) );
INV_X1 U1083 ( .A(G104), .ZN(n1195) );
NAND2_X1 U1084 ( .A1(KEYINPUT18), .A2(n1151), .ZN(n1375) );
XNOR2_X1 U1085 ( .A(G125), .B(n1211), .ZN(n1151) );
INV_X1 U1086 ( .A(G140), .ZN(n1211) );
XOR2_X1 U1087 ( .A(G131), .B(n1379), .Z(n1373) );
AND3_X1 U1088 ( .A1(G214), .A2(n1150), .A3(n1330), .ZN(n1379) );
INV_X1 U1089 ( .A(G237), .ZN(n1330) );
INV_X1 U1090 ( .A(G953), .ZN(n1150) );
XOR2_X1 U1091 ( .A(n1380), .B(n1381), .Z(n1371) );
XOR2_X1 U1092 ( .A(G146), .B(G143), .Z(n1381) );
XNOR2_X1 U1093 ( .A(KEYINPUT25), .B(KEYINPUT22), .ZN(n1380) );
XOR2_X1 U1094 ( .A(n1115), .B(n1114), .Z(n1275) );
INV_X1 U1095 ( .A(G478), .ZN(n1114) );
NOR2_X1 U1096 ( .A1(n1190), .A2(G902), .ZN(n1115) );
INV_X1 U1097 ( .A(n1188), .ZN(n1190) );
XNOR2_X1 U1098 ( .A(n1382), .B(n1383), .ZN(n1188) );
NOR3_X1 U1099 ( .A1(n1384), .A2(G953), .A3(n1385), .ZN(n1383) );
INV_X1 U1100 ( .A(G234), .ZN(n1385) );
XNOR2_X1 U1101 ( .A(KEYINPUT47), .B(n1181), .ZN(n1384) );
INV_X1 U1102 ( .A(G217), .ZN(n1181) );
NAND3_X1 U1103 ( .A1(n1386), .A2(n1387), .A3(KEYINPUT36), .ZN(n1382) );
NAND2_X1 U1104 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
NAND2_X1 U1105 ( .A1(KEYINPUT3), .A2(n1390), .ZN(n1389) );
XOR2_X1 U1106 ( .A(n1391), .B(n1392), .Z(n1388) );
NOR2_X1 U1107 ( .A1(G107), .A2(n1393), .ZN(n1391) );
NAND3_X1 U1108 ( .A1(n1394), .A2(n1390), .A3(KEYINPUT3), .ZN(n1386) );
XOR2_X1 U1109 ( .A(G122), .B(G116), .Z(n1390) );
XOR2_X1 U1110 ( .A(n1395), .B(n1392), .Z(n1394) );
XOR2_X1 U1111 ( .A(G134), .B(n1369), .Z(n1392) );
XOR2_X1 U1112 ( .A(G128), .B(G143), .Z(n1369) );
NOR2_X1 U1113 ( .A1(n1351), .A2(n1393), .ZN(n1395) );
INV_X1 U1114 ( .A(KEYINPUT61), .ZN(n1393) );
INV_X1 U1115 ( .A(G107), .ZN(n1351) );
endmodule


