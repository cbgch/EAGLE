//Key = 1011000110110001100100110001000000011110000110101101100110010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323;

XNOR2_X1 U716 ( .A(G107), .B(n1006), .ZN(G9) );
NOR2_X1 U717 ( .A1(n1007), .A2(n1008), .ZN(G75) );
NOR4_X1 U718 ( .A1(n1009), .A2(n1010), .A3(G953), .A4(n1011), .ZN(n1008) );
NOR3_X1 U719 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1010) );
NOR2_X1 U720 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U721 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NOR2_X1 U722 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR2_X1 U723 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR3_X1 U724 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1021) );
NOR3_X1 U725 ( .A1(n1026), .A2(KEYINPUT28), .A3(n1027), .ZN(n1025) );
AND2_X1 U726 ( .A1(n1026), .A2(KEYINPUT28), .ZN(n1024) );
NOR3_X1 U727 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1019) );
NOR3_X1 U728 ( .A1(n1028), .A2(n1022), .A3(n1031), .ZN(n1015) );
INV_X1 U729 ( .A(n1032), .ZN(n1022) );
NAND3_X1 U730 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1009) );
NAND2_X1 U731 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NAND2_X1 U732 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND3_X1 U733 ( .A1(n1032), .A2(n1040), .A3(n1041), .ZN(n1039) );
INV_X1 U734 ( .A(n1012), .ZN(n1041) );
NAND2_X1 U735 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NAND2_X1 U736 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U737 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U738 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XNOR2_X1 U739 ( .A(KEYINPUT14), .B(n1050), .ZN(n1049) );
INV_X1 U740 ( .A(n1051), .ZN(n1046) );
NAND2_X1 U741 ( .A1(n1052), .A2(n1053), .ZN(n1042) );
XOR2_X1 U742 ( .A(KEYINPUT7), .B(n1054), .Z(n1038) );
NOR4_X1 U743 ( .A1(n1018), .A2(n1055), .A3(n1012), .A4(n1056), .ZN(n1054) );
XNOR2_X1 U744 ( .A(n1014), .B(KEYINPUT55), .ZN(n1056) );
INV_X1 U745 ( .A(n1053), .ZN(n1014) );
INV_X1 U746 ( .A(n1057), .ZN(n1055) );
NOR3_X1 U747 ( .A1(n1011), .A2(G953), .A3(G952), .ZN(n1007) );
AND4_X1 U748 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1011) );
NOR4_X1 U749 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1061) );
XNOR2_X1 U750 ( .A(n1066), .B(n1067), .ZN(n1065) );
NOR2_X1 U751 ( .A1(KEYINPUT9), .A2(n1068), .ZN(n1067) );
XNOR2_X1 U752 ( .A(n1069), .B(KEYINPUT15), .ZN(n1062) );
NOR3_X1 U753 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1060) );
NAND2_X1 U754 ( .A1(n1073), .A2(n1074), .ZN(n1059) );
XNOR2_X1 U755 ( .A(G469), .B(n1075), .ZN(n1058) );
NAND2_X1 U756 ( .A1(n1076), .A2(KEYINPUT36), .ZN(n1075) );
XOR2_X1 U757 ( .A(n1077), .B(KEYINPUT42), .Z(n1076) );
XOR2_X1 U758 ( .A(n1078), .B(n1079), .Z(G72) );
NOR2_X1 U759 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR2_X1 U760 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NAND2_X1 U761 ( .A1(n1084), .A2(n1085), .ZN(n1078) );
NAND2_X1 U762 ( .A1(n1086), .A2(n1081), .ZN(n1085) );
XNOR2_X1 U763 ( .A(n1087), .B(n1033), .ZN(n1086) );
NAND3_X1 U764 ( .A1(G900), .A2(n1087), .A3(G953), .ZN(n1084) );
XNOR2_X1 U765 ( .A(n1088), .B(n1089), .ZN(n1087) );
XNOR2_X1 U766 ( .A(KEYINPUT19), .B(n1090), .ZN(n1089) );
XNOR2_X1 U767 ( .A(n1091), .B(n1092), .ZN(n1088) );
INV_X1 U768 ( .A(n1093), .ZN(n1092) );
NAND2_X1 U769 ( .A1(KEYINPUT44), .A2(n1094), .ZN(n1091) );
XOR2_X1 U770 ( .A(n1095), .B(n1096), .Z(G69) );
NOR2_X1 U771 ( .A1(n1035), .A2(G953), .ZN(n1096) );
XOR2_X1 U772 ( .A(n1097), .B(n1098), .Z(n1095) );
NOR2_X1 U773 ( .A1(KEYINPUT50), .A2(n1099), .ZN(n1098) );
NOR2_X1 U774 ( .A1(n1100), .A2(n1081), .ZN(n1099) );
NOR2_X1 U775 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U776 ( .A1(n1103), .A2(n1104), .ZN(n1097) );
NAND2_X1 U777 ( .A1(G953), .A2(n1102), .ZN(n1104) );
XOR2_X1 U778 ( .A(n1105), .B(n1106), .Z(n1103) );
XNOR2_X1 U779 ( .A(n1107), .B(n1108), .ZN(n1106) );
XNOR2_X1 U780 ( .A(KEYINPUT24), .B(n1109), .ZN(n1105) );
NOR2_X1 U781 ( .A1(n1110), .A2(n1111), .ZN(G66) );
XOR2_X1 U782 ( .A(n1112), .B(n1113), .Z(n1111) );
OR2_X1 U783 ( .A1(n1114), .A2(n1068), .ZN(n1112) );
NOR2_X1 U784 ( .A1(n1110), .A2(n1115), .ZN(G63) );
XOR2_X1 U785 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR3_X1 U786 ( .A1(n1114), .A2(KEYINPUT41), .A3(n1118), .ZN(n1116) );
NOR2_X1 U787 ( .A1(n1110), .A2(n1119), .ZN(G60) );
XOR2_X1 U788 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U789 ( .A1(n1122), .A2(G475), .ZN(n1120) );
NAND3_X1 U790 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(G6) );
NAND2_X1 U791 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U792 ( .A1(n1128), .A2(n1129), .ZN(n1124) );
INV_X1 U793 ( .A(KEYINPUT0), .ZN(n1129) );
NAND2_X1 U794 ( .A1(n1130), .A2(G104), .ZN(n1128) );
XNOR2_X1 U795 ( .A(n1126), .B(KEYINPUT54), .ZN(n1130) );
NAND2_X1 U796 ( .A1(KEYINPUT0), .A2(n1131), .ZN(n1123) );
NAND2_X1 U797 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
OR3_X1 U798 ( .A1(n1127), .A2(n1126), .A3(KEYINPUT54), .ZN(n1133) );
NAND2_X1 U799 ( .A1(KEYINPUT54), .A2(n1126), .ZN(n1132) );
NOR3_X1 U800 ( .A1(n1134), .A2(n1110), .A3(n1135), .ZN(G57) );
NOR3_X1 U801 ( .A1(n1136), .A2(KEYINPUT34), .A3(n1137), .ZN(n1135) );
XOR2_X1 U802 ( .A(n1138), .B(n1139), .Z(n1136) );
NOR2_X1 U803 ( .A1(G101), .A2(n1140), .ZN(n1139) );
NOR2_X1 U804 ( .A1(n1141), .A2(n1142), .ZN(n1134) );
XOR2_X1 U805 ( .A(n1138), .B(n1143), .Z(n1142) );
NOR2_X1 U806 ( .A1(n1144), .A2(n1140), .ZN(n1143) );
INV_X1 U807 ( .A(KEYINPUT63), .ZN(n1140) );
XNOR2_X1 U808 ( .A(n1145), .B(n1109), .ZN(n1138) );
XOR2_X1 U809 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U810 ( .A1(n1122), .A2(G472), .ZN(n1146) );
NOR2_X1 U811 ( .A1(KEYINPUT34), .A2(n1137), .ZN(n1141) );
NOR2_X1 U812 ( .A1(n1148), .A2(n1149), .ZN(G54) );
XOR2_X1 U813 ( .A(KEYINPUT53), .B(n1110), .Z(n1149) );
XOR2_X1 U814 ( .A(n1150), .B(n1151), .Z(n1148) );
XNOR2_X1 U815 ( .A(n1152), .B(n1093), .ZN(n1151) );
XNOR2_X1 U816 ( .A(n1153), .B(n1154), .ZN(n1093) );
XOR2_X1 U817 ( .A(n1155), .B(n1156), .Z(n1150) );
XOR2_X1 U818 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U819 ( .A1(KEYINPUT10), .A2(G110), .ZN(n1157) );
NAND2_X1 U820 ( .A1(n1122), .A2(G469), .ZN(n1155) );
NOR2_X1 U821 ( .A1(n1110), .A2(n1159), .ZN(G51) );
XOR2_X1 U822 ( .A(n1160), .B(n1161), .Z(n1159) );
NAND2_X1 U823 ( .A1(n1122), .A2(n1073), .ZN(n1161) );
INV_X1 U824 ( .A(n1114), .ZN(n1122) );
NAND2_X1 U825 ( .A1(G902), .A2(n1162), .ZN(n1114) );
NAND2_X1 U826 ( .A1(n1163), .A2(n1033), .ZN(n1162) );
AND4_X1 U827 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1033) );
NOR4_X1 U828 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
NOR2_X1 U829 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XNOR2_X1 U830 ( .A(n1174), .B(KEYINPUT57), .ZN(n1172) );
INV_X1 U831 ( .A(n1175), .ZN(n1169) );
INV_X1 U832 ( .A(n1176), .ZN(n1168) );
NOR2_X1 U833 ( .A1(n1177), .A2(n1178), .ZN(n1166) );
INV_X1 U834 ( .A(n1179), .ZN(n1178) );
NOR2_X1 U835 ( .A1(n1180), .A2(n1028), .ZN(n1177) );
INV_X1 U836 ( .A(n1036), .ZN(n1028) );
XNOR2_X1 U837 ( .A(n1035), .B(KEYINPUT35), .ZN(n1163) );
AND4_X1 U838 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1035) );
AND4_X1 U839 ( .A1(n1006), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1184) );
NAND3_X1 U840 ( .A1(n1174), .A2(n1032), .A3(n1188), .ZN(n1006) );
NOR2_X1 U841 ( .A1(n1189), .A2(n1126), .ZN(n1183) );
AND3_X1 U842 ( .A1(n1188), .A2(n1032), .A3(n1052), .ZN(n1126) );
NAND2_X1 U843 ( .A1(n1190), .A2(n1191), .ZN(n1160) );
NAND2_X1 U844 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U845 ( .A(n1194), .B(KEYINPUT45), .Z(n1190) );
OR2_X1 U846 ( .A1(n1192), .A2(n1193), .ZN(n1194) );
XOR2_X1 U847 ( .A(G125), .B(n1195), .Z(n1192) );
NOR2_X1 U848 ( .A1(n1081), .A2(G952), .ZN(n1110) );
NAND2_X1 U849 ( .A1(n1196), .A2(n1197), .ZN(G48) );
NAND2_X1 U850 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XNOR2_X1 U851 ( .A(n1170), .B(KEYINPUT11), .ZN(n1198) );
NAND2_X1 U852 ( .A1(G146), .A2(n1200), .ZN(n1196) );
XNOR2_X1 U853 ( .A(n1170), .B(KEYINPUT20), .ZN(n1200) );
NOR2_X1 U854 ( .A1(n1173), .A2(n1201), .ZN(n1170) );
NAND2_X1 U855 ( .A1(n1202), .A2(n1203), .ZN(G45) );
NAND2_X1 U856 ( .A1(G143), .A2(n1175), .ZN(n1203) );
XOR2_X1 U857 ( .A(n1204), .B(KEYINPUT1), .Z(n1202) );
OR2_X1 U858 ( .A1(n1175), .A2(G143), .ZN(n1204) );
NAND4_X1 U859 ( .A1(n1205), .A2(n1023), .A3(n1064), .A4(n1069), .ZN(n1175) );
XNOR2_X1 U860 ( .A(G140), .B(n1176), .ZN(G42) );
NAND3_X1 U861 ( .A1(n1036), .A2(n1206), .A3(n1207), .ZN(n1176) );
XNOR2_X1 U862 ( .A(G137), .B(n1164), .ZN(G39) );
NAND4_X1 U863 ( .A1(n1036), .A2(n1206), .A3(n1208), .A4(n1044), .ZN(n1164) );
XOR2_X1 U864 ( .A(n1209), .B(n1210), .Z(G36) );
NAND2_X1 U865 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XNOR2_X1 U866 ( .A(G134), .B(KEYINPUT3), .ZN(n1212) );
XNOR2_X1 U867 ( .A(KEYINPUT56), .B(KEYINPUT51), .ZN(n1211) );
NAND2_X1 U868 ( .A1(n1036), .A2(n1213), .ZN(n1209) );
XNOR2_X1 U869 ( .A(KEYINPUT33), .B(n1180), .ZN(n1213) );
NAND2_X1 U870 ( .A1(n1205), .A2(n1174), .ZN(n1180) );
XNOR2_X1 U871 ( .A(G131), .B(n1165), .ZN(G33) );
NAND3_X1 U872 ( .A1(n1205), .A2(n1052), .A3(n1036), .ZN(n1165) );
NOR2_X1 U873 ( .A1(n1026), .A2(n1072), .ZN(n1036) );
INV_X1 U874 ( .A(n1214), .ZN(n1026) );
AND2_X1 U875 ( .A1(n1206), .A2(n1057), .ZN(n1205) );
XNOR2_X1 U876 ( .A(n1215), .B(n1216), .ZN(G30) );
NOR3_X1 U877 ( .A1(n1173), .A2(KEYINPUT39), .A3(n1031), .ZN(n1216) );
INV_X1 U878 ( .A(n1174), .ZN(n1031) );
NAND3_X1 U879 ( .A1(n1208), .A2(n1023), .A3(n1206), .ZN(n1173) );
AND2_X1 U880 ( .A1(n1051), .A2(n1217), .ZN(n1206) );
XNOR2_X1 U881 ( .A(G101), .B(n1218), .ZN(G3) );
NAND2_X1 U882 ( .A1(KEYINPUT48), .A2(n1189), .ZN(n1218) );
AND3_X1 U883 ( .A1(n1044), .A2(n1188), .A3(n1057), .ZN(n1189) );
XNOR2_X1 U884 ( .A(G125), .B(n1179), .ZN(G27) );
NAND4_X1 U885 ( .A1(n1207), .A2(n1023), .A3(n1053), .A4(n1217), .ZN(n1179) );
NAND2_X1 U886 ( .A1(n1219), .A2(n1220), .ZN(n1217) );
NAND4_X1 U887 ( .A1(G953), .A2(G902), .A3(n1221), .A4(n1083), .ZN(n1220) );
INV_X1 U888 ( .A(G900), .ZN(n1083) );
XNOR2_X1 U889 ( .A(KEYINPUT46), .B(n1012), .ZN(n1219) );
NOR3_X1 U890 ( .A1(n1030), .A2(n1029), .A3(n1201), .ZN(n1207) );
XNOR2_X1 U891 ( .A(G122), .B(n1181), .ZN(G24) );
NAND4_X1 U892 ( .A1(n1222), .A2(n1032), .A3(n1064), .A4(n1069), .ZN(n1181) );
NOR2_X1 U893 ( .A1(n1030), .A2(n1223), .ZN(n1032) );
XNOR2_X1 U894 ( .A(G119), .B(n1187), .ZN(G21) );
NAND3_X1 U895 ( .A1(n1222), .A2(n1044), .A3(n1208), .ZN(n1187) );
NOR2_X1 U896 ( .A1(n1029), .A2(n1224), .ZN(n1208) );
XNOR2_X1 U897 ( .A(G116), .B(n1186), .ZN(G18) );
NAND3_X1 U898 ( .A1(n1222), .A2(n1174), .A3(n1057), .ZN(n1186) );
NOR2_X1 U899 ( .A1(n1225), .A2(n1226), .ZN(n1174) );
XNOR2_X1 U900 ( .A(G113), .B(n1185), .ZN(G15) );
NAND3_X1 U901 ( .A1(n1057), .A2(n1222), .A3(n1052), .ZN(n1185) );
INV_X1 U902 ( .A(n1201), .ZN(n1052) );
NAND2_X1 U903 ( .A1(n1226), .A2(n1069), .ZN(n1201) );
AND3_X1 U904 ( .A1(n1053), .A2(n1227), .A3(n1023), .ZN(n1222) );
NAND2_X1 U905 ( .A1(n1228), .A2(n1229), .ZN(n1053) );
OR3_X1 U906 ( .A1(n1230), .A2(n1070), .A3(KEYINPUT5), .ZN(n1229) );
NAND2_X1 U907 ( .A1(KEYINPUT5), .A2(n1051), .ZN(n1228) );
NOR2_X1 U908 ( .A1(n1223), .A2(n1224), .ZN(n1057) );
XNOR2_X1 U909 ( .A(G110), .B(n1231), .ZN(G12) );
NAND2_X1 U910 ( .A1(KEYINPUT23), .A2(n1232), .ZN(n1231) );
INV_X1 U911 ( .A(n1182), .ZN(n1232) );
NAND4_X1 U912 ( .A1(n1044), .A2(n1188), .A3(n1224), .A4(n1223), .ZN(n1182) );
INV_X1 U913 ( .A(n1029), .ZN(n1223) );
XNOR2_X1 U914 ( .A(n1066), .B(n1068), .ZN(n1029) );
NAND2_X1 U915 ( .A1(G217), .A2(n1233), .ZN(n1068) );
NAND2_X1 U916 ( .A1(n1234), .A2(n1235), .ZN(n1066) );
XOR2_X1 U917 ( .A(KEYINPUT26), .B(n1113), .Z(n1234) );
XNOR2_X1 U918 ( .A(n1236), .B(n1237), .ZN(n1113) );
XOR2_X1 U919 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U920 ( .A(n1240), .B(n1241), .Z(n1239) );
NOR2_X1 U921 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U922 ( .A(n1244), .B(KEYINPUT27), .Z(n1243) );
NAND2_X1 U923 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
XOR2_X1 U924 ( .A(n1247), .B(KEYINPUT12), .Z(n1245) );
NOR2_X1 U925 ( .A1(n1246), .A2(n1247), .ZN(n1242) );
NAND2_X1 U926 ( .A1(n1248), .A2(G221), .ZN(n1247) );
NOR2_X1 U927 ( .A1(KEYINPUT13), .A2(n1249), .ZN(n1240) );
XNOR2_X1 U928 ( .A(G110), .B(n1250), .ZN(n1249) );
XNOR2_X1 U929 ( .A(n1215), .B(G119), .ZN(n1250) );
NOR2_X1 U930 ( .A1(G146), .A2(KEYINPUT4), .ZN(n1238) );
XNOR2_X1 U931 ( .A(G125), .B(n1251), .ZN(n1236) );
XNOR2_X1 U932 ( .A(KEYINPUT38), .B(n1252), .ZN(n1251) );
INV_X1 U933 ( .A(n1030), .ZN(n1224) );
XOR2_X1 U934 ( .A(n1063), .B(KEYINPUT60), .Z(n1030) );
XNOR2_X1 U935 ( .A(n1253), .B(G472), .ZN(n1063) );
NAND2_X1 U936 ( .A1(n1254), .A2(n1235), .ZN(n1253) );
XOR2_X1 U937 ( .A(n1147), .B(n1255), .Z(n1254) );
XOR2_X1 U938 ( .A(n1256), .B(n1257), .Z(n1255) );
NAND2_X1 U939 ( .A1(KEYINPUT16), .A2(n1109), .ZN(n1257) );
NAND3_X1 U940 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1256) );
OR2_X1 U941 ( .A1(n1137), .A2(KEYINPUT37), .ZN(n1260) );
INV_X1 U942 ( .A(n1261), .ZN(n1137) );
NAND3_X1 U943 ( .A1(KEYINPUT37), .A2(n1262), .A3(n1144), .ZN(n1259) );
OR2_X1 U944 ( .A1(n1144), .A2(n1262), .ZN(n1258) );
NOR2_X1 U945 ( .A1(KEYINPUT6), .A2(n1261), .ZN(n1262) );
NAND2_X1 U946 ( .A1(n1263), .A2(G210), .ZN(n1261) );
XOR2_X1 U947 ( .A(n1094), .B(n1264), .Z(n1147) );
XNOR2_X1 U948 ( .A(n1265), .B(n1266), .ZN(n1264) );
AND3_X1 U949 ( .A1(n1051), .A2(n1227), .A3(n1023), .ZN(n1188) );
NOR2_X1 U950 ( .A1(n1072), .A2(n1214), .ZN(n1023) );
NOR2_X1 U951 ( .A1(n1267), .A2(n1071), .ZN(n1214) );
NOR2_X1 U952 ( .A1(n1074), .A2(n1073), .ZN(n1071) );
XNOR2_X1 U953 ( .A(n1268), .B(KEYINPUT29), .ZN(n1267) );
NAND2_X1 U954 ( .A1(n1269), .A2(n1074), .ZN(n1268) );
NAND2_X1 U955 ( .A1(n1270), .A2(n1235), .ZN(n1074) );
XOR2_X1 U956 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U957 ( .A(n1273), .B(n1195), .Z(n1272) );
XNOR2_X1 U958 ( .A(n1266), .B(n1274), .ZN(n1195) );
XNOR2_X1 U959 ( .A(n1199), .B(n1275), .ZN(n1274) );
NOR2_X1 U960 ( .A1(G953), .A2(n1101), .ZN(n1275) );
INV_X1 U961 ( .A(G224), .ZN(n1101) );
XNOR2_X1 U962 ( .A(n1276), .B(n1277), .ZN(n1266) );
NOR2_X1 U963 ( .A1(KEYINPUT18), .A2(n1215), .ZN(n1277) );
NOR2_X1 U964 ( .A1(G143), .A2(KEYINPUT17), .ZN(n1276) );
NOR2_X1 U965 ( .A1(G125), .A2(KEYINPUT61), .ZN(n1273) );
XOR2_X1 U966 ( .A(n1193), .B(KEYINPUT31), .Z(n1271) );
NAND2_X1 U967 ( .A1(n1278), .A2(n1279), .ZN(n1193) );
NAND2_X1 U968 ( .A1(n1280), .A2(n1107), .ZN(n1279) );
XOR2_X1 U969 ( .A(KEYINPUT49), .B(n1281), .Z(n1278) );
NOR2_X1 U970 ( .A1(n1280), .A2(n1107), .ZN(n1281) );
XNOR2_X1 U971 ( .A(n1282), .B(G122), .ZN(n1107) );
XNOR2_X1 U972 ( .A(n1109), .B(n1283), .ZN(n1280) );
NOR2_X1 U973 ( .A1(KEYINPUT62), .A2(n1108), .ZN(n1283) );
XOR2_X1 U974 ( .A(n1284), .B(n1285), .Z(n1108) );
NOR2_X1 U975 ( .A1(KEYINPUT47), .A2(n1144), .ZN(n1285) );
INV_X1 U976 ( .A(G101), .ZN(n1144) );
XNOR2_X1 U977 ( .A(G107), .B(G104), .ZN(n1284) );
XOR2_X1 U978 ( .A(n1286), .B(n1287), .Z(n1109) );
XNOR2_X1 U979 ( .A(G116), .B(G119), .ZN(n1286) );
XOR2_X1 U980 ( .A(KEYINPUT32), .B(n1073), .Z(n1269) );
AND2_X1 U981 ( .A1(G210), .A2(n1288), .ZN(n1073) );
INV_X1 U982 ( .A(n1027), .ZN(n1072) );
NAND2_X1 U983 ( .A1(G214), .A2(n1288), .ZN(n1027) );
NAND2_X1 U984 ( .A1(n1235), .A2(n1289), .ZN(n1288) );
INV_X1 U985 ( .A(G237), .ZN(n1289) );
NAND2_X1 U986 ( .A1(n1012), .A2(n1290), .ZN(n1227) );
NAND4_X1 U987 ( .A1(G953), .A2(G902), .A3(n1221), .A4(n1102), .ZN(n1290) );
INV_X1 U988 ( .A(G898), .ZN(n1102) );
NAND3_X1 U989 ( .A1(n1221), .A2(n1081), .A3(G952), .ZN(n1012) );
NAND2_X1 U990 ( .A1(G237), .A2(G234), .ZN(n1221) );
NOR2_X1 U991 ( .A1(n1048), .A2(n1070), .ZN(n1051) );
INV_X1 U992 ( .A(n1050), .ZN(n1070) );
NAND2_X1 U993 ( .A1(G221), .A2(n1233), .ZN(n1050) );
NAND2_X1 U994 ( .A1(G234), .A2(n1235), .ZN(n1233) );
INV_X1 U995 ( .A(n1230), .ZN(n1048) );
XOR2_X1 U996 ( .A(G469), .B(n1291), .Z(n1230) );
NOR2_X1 U997 ( .A1(KEYINPUT25), .A2(n1077), .ZN(n1291) );
NAND2_X1 U998 ( .A1(n1292), .A2(n1235), .ZN(n1077) );
XOR2_X1 U999 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U1000 ( .A(n1152), .B(n1154), .Z(n1294) );
XNOR2_X1 U1001 ( .A(n1215), .B(KEYINPUT21), .ZN(n1154) );
INV_X1 U1002 ( .A(G128), .ZN(n1215) );
XOR2_X1 U1003 ( .A(n1295), .B(n1296), .Z(n1152) );
XNOR2_X1 U1004 ( .A(n1127), .B(G101), .ZN(n1296) );
INV_X1 U1005 ( .A(G104), .ZN(n1127) );
XOR2_X1 U1006 ( .A(n1297), .B(n1094), .Z(n1295) );
XNOR2_X1 U1007 ( .A(G134), .B(n1246), .ZN(n1094) );
INV_X1 U1008 ( .A(G137), .ZN(n1246) );
NAND2_X1 U1009 ( .A1(KEYINPUT52), .A2(n1298), .ZN(n1297) );
INV_X1 U1010 ( .A(G107), .ZN(n1298) );
XOR2_X1 U1011 ( .A(n1299), .B(n1300), .Z(n1293) );
NAND2_X1 U1012 ( .A1(n1301), .A2(n1302), .ZN(n1299) );
NAND2_X1 U1013 ( .A1(n1158), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1014 ( .A(n1304), .B(KEYINPUT58), .Z(n1301) );
OR2_X1 U1015 ( .A1(n1303), .A2(n1158), .ZN(n1304) );
NOR2_X1 U1016 ( .A1(n1082), .A2(G953), .ZN(n1158) );
INV_X1 U1017 ( .A(G227), .ZN(n1082) );
XNOR2_X1 U1018 ( .A(n1282), .B(n1252), .ZN(n1303) );
INV_X1 U1019 ( .A(G140), .ZN(n1252) );
INV_X1 U1020 ( .A(G110), .ZN(n1282) );
INV_X1 U1021 ( .A(n1018), .ZN(n1044) );
NAND2_X1 U1022 ( .A1(n1226), .A2(n1305), .ZN(n1018) );
XOR2_X1 U1023 ( .A(KEYINPUT22), .B(n1225), .Z(n1305) );
XOR2_X1 U1024 ( .A(n1069), .B(KEYINPUT40), .Z(n1225) );
XNOR2_X1 U1025 ( .A(n1306), .B(G475), .ZN(n1069) );
NAND2_X1 U1026 ( .A1(n1307), .A2(n1235), .ZN(n1306) );
INV_X1 U1027 ( .A(G902), .ZN(n1235) );
XNOR2_X1 U1028 ( .A(n1121), .B(KEYINPUT2), .ZN(n1307) );
XNOR2_X1 U1029 ( .A(n1308), .B(n1309), .ZN(n1121) );
XOR2_X1 U1030 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U1031 ( .A(G122), .B(G104), .ZN(n1311) );
NAND2_X1 U1032 ( .A1(KEYINPUT59), .A2(n1090), .ZN(n1310) );
INV_X1 U1033 ( .A(G125), .ZN(n1090) );
XOR2_X1 U1034 ( .A(n1153), .B(n1312), .Z(n1308) );
XNOR2_X1 U1035 ( .A(n1313), .B(n1287), .ZN(n1312) );
XOR2_X1 U1036 ( .A(G113), .B(KEYINPUT43), .Z(n1287) );
NAND2_X1 U1037 ( .A1(n1263), .A2(G214), .ZN(n1313) );
NOR2_X1 U1038 ( .A1(G953), .A2(G237), .ZN(n1263) );
XNOR2_X1 U1039 ( .A(n1300), .B(G140), .ZN(n1153) );
XOR2_X1 U1040 ( .A(G143), .B(n1265), .Z(n1300) );
XNOR2_X1 U1041 ( .A(G131), .B(n1199), .ZN(n1265) );
INV_X1 U1042 ( .A(G146), .ZN(n1199) );
INV_X1 U1043 ( .A(n1064), .ZN(n1226) );
XOR2_X1 U1044 ( .A(n1314), .B(n1118), .Z(n1064) );
INV_X1 U1045 ( .A(G478), .ZN(n1118) );
OR2_X1 U1046 ( .A1(n1117), .A2(G902), .ZN(n1314) );
XNOR2_X1 U1047 ( .A(n1315), .B(n1316), .ZN(n1117) );
XOR2_X1 U1048 ( .A(n1317), .B(n1318), .Z(n1316) );
NAND2_X1 U1049 ( .A1(G217), .A2(n1248), .ZN(n1318) );
AND2_X1 U1050 ( .A1(G234), .A2(n1081), .ZN(n1248) );
INV_X1 U1051 ( .A(G953), .ZN(n1081) );
NAND2_X1 U1052 ( .A1(KEYINPUT8), .A2(n1319), .ZN(n1317) );
XOR2_X1 U1053 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1054 ( .A(G143), .B(G134), .Z(n1321) );
NOR2_X1 U1055 ( .A1(G128), .A2(KEYINPUT30), .ZN(n1320) );
XNOR2_X1 U1056 ( .A(G107), .B(n1322), .ZN(n1315) );
XNOR2_X1 U1057 ( .A(n1323), .B(G116), .ZN(n1322) );
INV_X1 U1058 ( .A(G122), .ZN(n1323) );
endmodule


