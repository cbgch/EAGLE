//Key = 0101001101111101010000010001101001101110001111111010101010011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
n1480, n1481, n1482;

XNOR2_X1 U810 ( .A(G107), .B(n1130), .ZN(G9) );
NAND3_X1 U811 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1130) );
XNOR2_X1 U812 ( .A(n1134), .B(KEYINPUT56), .ZN(n1133) );
NOR2_X1 U813 ( .A1(n1135), .A2(n1136), .ZN(G75) );
NOR3_X1 U814 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
NOR3_X1 U815 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1138) );
NOR4_X1 U816 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1142) );
NOR2_X1 U817 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NOR2_X1 U818 ( .A1(n1149), .A2(n1150), .ZN(n1147) );
NOR3_X1 U819 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1145) );
NOR4_X1 U820 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1153) );
NOR2_X1 U821 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NOR2_X1 U822 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
NOR2_X1 U823 ( .A1(KEYINPUT57), .A2(n1162), .ZN(n1160) );
NOR3_X1 U824 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1156) );
NOR2_X1 U825 ( .A1(n1166), .A2(n1167), .ZN(n1155) );
INV_X1 U826 ( .A(KEYINPUT1), .ZN(n1167) );
NOR2_X1 U827 ( .A1(n1168), .A2(n1169), .ZN(n1152) );
NOR2_X1 U828 ( .A1(KEYINPUT1), .A2(n1166), .ZN(n1169) );
NOR2_X1 U829 ( .A1(n1170), .A2(n1171), .ZN(n1144) );
INV_X1 U830 ( .A(KEYINPUT57), .ZN(n1171) );
NOR4_X1 U831 ( .A1(n1151), .A2(n1162), .A3(n1159), .A4(n1154), .ZN(n1170) );
NOR2_X1 U832 ( .A1(n1172), .A2(n1173), .ZN(n1141) );
NOR2_X1 U833 ( .A1(n1148), .A2(n1174), .ZN(n1172) );
XNOR2_X1 U834 ( .A(KEYINPUT9), .B(n1151), .ZN(n1174) );
NAND3_X1 U835 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1137) );
OR3_X1 U836 ( .A1(n1151), .A2(n1178), .A3(n1148), .ZN(n1177) );
NAND3_X1 U837 ( .A1(n1179), .A2(n1180), .A3(n1168), .ZN(n1148) );
INV_X1 U838 ( .A(n1154), .ZN(n1168) );
INV_X1 U839 ( .A(n1134), .ZN(n1151) );
NOR3_X1 U840 ( .A1(n1181), .A2(G953), .A3(G952), .ZN(n1135) );
INV_X1 U841 ( .A(n1175), .ZN(n1181) );
NAND4_X1 U842 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1175) );
NOR4_X1 U843 ( .A1(n1186), .A2(n1143), .A3(n1187), .A4(n1188), .ZN(n1185) );
XOR2_X1 U844 ( .A(n1189), .B(KEYINPUT31), .Z(n1188) );
NAND3_X1 U845 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1189) );
OR2_X1 U846 ( .A1(n1193), .A2(KEYINPUT37), .ZN(n1191) );
NAND3_X1 U847 ( .A1(n1193), .A2(n1194), .A3(KEYINPUT37), .ZN(n1190) );
XNOR2_X1 U848 ( .A(n1195), .B(n1196), .ZN(n1187) );
NOR2_X1 U849 ( .A1(G478), .A2(KEYINPUT51), .ZN(n1196) );
NOR2_X1 U850 ( .A1(n1197), .A2(n1198), .ZN(n1184) );
XNOR2_X1 U851 ( .A(KEYINPUT19), .B(n1199), .ZN(n1198) );
XOR2_X1 U852 ( .A(n1200), .B(n1201), .Z(n1197) );
XNOR2_X1 U853 ( .A(KEYINPUT36), .B(n1202), .ZN(n1201) );
NOR2_X1 U854 ( .A1(KEYINPUT63), .A2(G469), .ZN(n1202) );
XOR2_X1 U855 ( .A(n1203), .B(n1204), .Z(G72) );
XOR2_X1 U856 ( .A(n1205), .B(n1206), .Z(n1204) );
NOR2_X1 U857 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XNOR2_X1 U858 ( .A(G953), .B(KEYINPUT45), .ZN(n1208) );
NAND2_X1 U859 ( .A1(n1209), .A2(n1210), .ZN(n1205) );
INV_X1 U860 ( .A(n1211), .ZN(n1210) );
XOR2_X1 U861 ( .A(n1212), .B(n1213), .Z(n1209) );
XOR2_X1 U862 ( .A(n1214), .B(n1215), .Z(n1213) );
NOR2_X1 U863 ( .A1(KEYINPUT0), .A2(n1216), .ZN(n1214) );
XNOR2_X1 U864 ( .A(G131), .B(n1217), .ZN(n1216) );
NOR2_X1 U865 ( .A1(KEYINPUT2), .A2(n1218), .ZN(n1217) );
XOR2_X1 U866 ( .A(KEYINPUT20), .B(n1219), .Z(n1218) );
NAND2_X1 U867 ( .A1(n1220), .A2(n1221), .ZN(n1212) );
NAND2_X1 U868 ( .A1(G125), .A2(n1222), .ZN(n1221) );
NAND2_X1 U869 ( .A1(G140), .A2(n1223), .ZN(n1222) );
NAND3_X1 U870 ( .A1(G140), .A2(n1223), .A3(n1224), .ZN(n1220) );
INV_X1 U871 ( .A(KEYINPUT8), .ZN(n1223) );
NAND2_X1 U872 ( .A1(G953), .A2(n1225), .ZN(n1203) );
NAND2_X1 U873 ( .A1(G900), .A2(G227), .ZN(n1225) );
XOR2_X1 U874 ( .A(n1226), .B(n1227), .Z(G69) );
NAND2_X1 U875 ( .A1(G953), .A2(n1228), .ZN(n1227) );
NAND2_X1 U876 ( .A1(G898), .A2(G224), .ZN(n1228) );
NAND2_X1 U877 ( .A1(KEYINPUT15), .A2(n1229), .ZN(n1226) );
XOR2_X1 U878 ( .A(n1230), .B(n1231), .Z(n1229) );
NOR2_X1 U879 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
INV_X1 U880 ( .A(n1234), .ZN(n1233) );
NOR2_X1 U881 ( .A1(n1235), .A2(n1236), .ZN(n1230) );
XNOR2_X1 U882 ( .A(G953), .B(KEYINPUT13), .ZN(n1236) );
NOR2_X1 U883 ( .A1(n1237), .A2(n1238), .ZN(G66) );
XOR2_X1 U884 ( .A(n1239), .B(n1240), .Z(n1238) );
NOR2_X1 U885 ( .A1(KEYINPUT18), .A2(n1241), .ZN(n1240) );
NOR2_X1 U886 ( .A1(n1242), .A2(n1243), .ZN(n1239) );
NOR2_X1 U887 ( .A1(n1237), .A2(n1244), .ZN(G63) );
NOR3_X1 U888 ( .A1(n1195), .A2(n1245), .A3(n1246), .ZN(n1244) );
AND4_X1 U889 ( .A1(n1247), .A2(KEYINPUT34), .A3(G478), .A4(n1248), .ZN(n1246) );
NOR2_X1 U890 ( .A1(n1249), .A2(n1247), .ZN(n1245) );
AND3_X1 U891 ( .A1(KEYINPUT34), .A2(n1139), .A3(G478), .ZN(n1249) );
NOR2_X1 U892 ( .A1(n1237), .A2(n1250), .ZN(G60) );
NOR2_X1 U893 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XOR2_X1 U894 ( .A(n1253), .B(n1254), .Z(n1252) );
NOR2_X1 U895 ( .A1(KEYINPUT21), .A2(n1255), .ZN(n1254) );
AND2_X1 U896 ( .A1(G475), .A2(n1248), .ZN(n1253) );
AND2_X1 U897 ( .A1(n1255), .A2(KEYINPUT21), .ZN(n1251) );
XOR2_X1 U898 ( .A(G104), .B(n1256), .Z(G6) );
NOR2_X1 U899 ( .A1(n1237), .A2(n1257), .ZN(G57) );
XOR2_X1 U900 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U901 ( .A(n1260), .B(n1261), .Z(n1258) );
AND2_X1 U902 ( .A1(G472), .A2(n1248), .ZN(n1261) );
NAND2_X1 U903 ( .A1(n1262), .A2(n1263), .ZN(n1260) );
NAND2_X1 U904 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
XOR2_X1 U905 ( .A(n1266), .B(KEYINPUT14), .Z(n1262) );
OR2_X1 U906 ( .A1(n1265), .A2(n1264), .ZN(n1266) );
NOR2_X1 U907 ( .A1(n1237), .A2(n1267), .ZN(G54) );
XOR2_X1 U908 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U909 ( .A(n1270), .B(n1271), .Z(n1269) );
XNOR2_X1 U910 ( .A(n1272), .B(n1273), .ZN(n1271) );
NOR2_X1 U911 ( .A1(G140), .A2(KEYINPUT4), .ZN(n1273) );
NAND2_X1 U912 ( .A1(KEYINPUT52), .A2(n1274), .ZN(n1272) );
AND2_X1 U913 ( .A1(G469), .A2(n1248), .ZN(n1270) );
INV_X1 U914 ( .A(n1243), .ZN(n1248) );
XNOR2_X1 U915 ( .A(n1275), .B(n1276), .ZN(n1268) );
NOR2_X1 U916 ( .A1(n1237), .A2(n1277), .ZN(G51) );
XOR2_X1 U917 ( .A(n1278), .B(n1279), .Z(n1277) );
NOR2_X1 U918 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NOR2_X1 U919 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
XOR2_X1 U920 ( .A(KEYINPUT62), .B(n1284), .Z(n1283) );
AND2_X1 U921 ( .A1(n1282), .A2(n1284), .ZN(n1280) );
XOR2_X1 U922 ( .A(G125), .B(n1285), .Z(n1284) );
NOR2_X1 U923 ( .A1(KEYINPUT39), .A2(n1234), .ZN(n1285) );
XNOR2_X1 U924 ( .A(n1286), .B(n1287), .ZN(n1278) );
NOR3_X1 U925 ( .A1(n1243), .A2(n1288), .A3(n1289), .ZN(n1287) );
NAND2_X1 U926 ( .A1(G902), .A2(n1139), .ZN(n1243) );
NAND2_X1 U927 ( .A1(n1207), .A2(n1235), .ZN(n1139) );
AND4_X1 U928 ( .A1(n1290), .A2(n1291), .A3(n1292), .A4(n1293), .ZN(n1235) );
NOR4_X1 U929 ( .A1(n1256), .A2(n1294), .A3(n1295), .A4(n1296), .ZN(n1293) );
NOR4_X1 U930 ( .A1(n1297), .A2(n1298), .A3(n1164), .A4(n1299), .ZN(n1296) );
INV_X1 U931 ( .A(n1149), .ZN(n1299) );
INV_X1 U932 ( .A(n1180), .ZN(n1164) );
NOR2_X1 U933 ( .A1(KEYINPUT23), .A2(n1300), .ZN(n1298) );
NOR2_X1 U934 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NOR2_X1 U935 ( .A1(n1132), .A2(n1303), .ZN(n1297) );
INV_X1 U936 ( .A(KEYINPUT23), .ZN(n1303) );
NOR2_X1 U937 ( .A1(n1304), .A2(n1178), .ZN(n1295) );
NOR3_X1 U938 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1304) );
XOR2_X1 U939 ( .A(n1308), .B(KEYINPUT17), .Z(n1307) );
NOR2_X1 U940 ( .A1(n1309), .A2(n1310), .ZN(n1306) );
NOR3_X1 U941 ( .A1(n1166), .A2(n1311), .A3(n1312), .ZN(n1309) );
NAND2_X1 U942 ( .A1(n1313), .A2(n1180), .ZN(n1166) );
XNOR2_X1 U943 ( .A(KEYINPUT32), .B(n1314), .ZN(n1305) );
AND3_X1 U944 ( .A1(n1132), .A2(n1134), .A3(n1161), .ZN(n1256) );
NAND2_X1 U945 ( .A1(KEYINPUT28), .A2(n1315), .ZN(n1292) );
NAND2_X1 U946 ( .A1(n1131), .A2(n1316), .ZN(n1291) );
NAND2_X1 U947 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND4_X1 U948 ( .A1(n1319), .A2(n1149), .A3(n1178), .A4(n1320), .ZN(n1318) );
INV_X1 U949 ( .A(KEYINPUT28), .ZN(n1320) );
NAND2_X1 U950 ( .A1(n1132), .A2(n1134), .ZN(n1317) );
NAND2_X1 U951 ( .A1(n1321), .A2(n1310), .ZN(n1290) );
INV_X1 U952 ( .A(KEYINPUT41), .ZN(n1310) );
AND4_X1 U953 ( .A1(n1322), .A2(n1323), .A3(n1324), .A4(n1325), .ZN(n1207) );
NOR4_X1 U954 ( .A1(n1326), .A2(n1327), .A3(n1328), .A4(n1329), .ZN(n1325) );
NOR3_X1 U955 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n1324) );
NOR3_X1 U956 ( .A1(n1333), .A2(n1334), .A3(n1335), .ZN(n1332) );
AND2_X1 U957 ( .A1(n1333), .A2(n1336), .ZN(n1331) );
INV_X1 U958 ( .A(KEYINPUT5), .ZN(n1333) );
NAND3_X1 U959 ( .A1(n1337), .A2(n1338), .A3(n1339), .ZN(n1323) );
OR2_X1 U960 ( .A1(n1340), .A2(KEYINPUT49), .ZN(n1338) );
NAND2_X1 U961 ( .A1(KEYINPUT49), .A2(n1341), .ZN(n1337) );
NAND4_X1 U962 ( .A1(n1199), .A2(n1342), .A3(n1313), .A4(n1173), .ZN(n1341) );
AND2_X1 U963 ( .A1(n1343), .A2(G953), .ZN(n1237) );
XNOR2_X1 U964 ( .A(G952), .B(KEYINPUT35), .ZN(n1343) );
XOR2_X1 U965 ( .A(G146), .B(n1329), .Z(G48) );
AND2_X1 U966 ( .A1(n1161), .A2(n1344), .ZN(n1329) );
XOR2_X1 U967 ( .A(G143), .B(n1330), .Z(G45) );
AND4_X1 U968 ( .A1(n1345), .A2(n1149), .A3(n1346), .A4(n1347), .ZN(n1330) );
NOR2_X1 U969 ( .A1(n1342), .A2(n1348), .ZN(n1346) );
XNOR2_X1 U970 ( .A(n1349), .B(n1328), .ZN(G42) );
AND3_X1 U971 ( .A1(n1161), .A2(n1340), .A3(n1150), .ZN(n1328) );
XOR2_X1 U972 ( .A(G137), .B(n1327), .Z(G39) );
AND4_X1 U973 ( .A1(n1340), .A2(n1180), .A3(n1350), .A4(n1351), .ZN(n1327) );
XNOR2_X1 U974 ( .A(G134), .B(n1322), .ZN(G36) );
NAND3_X1 U975 ( .A1(n1340), .A2(n1131), .A3(n1149), .ZN(n1322) );
NAND2_X1 U976 ( .A1(n1352), .A2(n1353), .ZN(G33) );
NAND3_X1 U977 ( .A1(n1354), .A2(n1355), .A3(n1339), .ZN(n1353) );
INV_X1 U978 ( .A(G131), .ZN(n1355) );
XOR2_X1 U979 ( .A(n1356), .B(KEYINPUT25), .Z(n1352) );
NAND2_X1 U980 ( .A1(G131), .A2(n1357), .ZN(n1356) );
NAND2_X1 U981 ( .A1(n1339), .A2(n1354), .ZN(n1357) );
NAND2_X1 U982 ( .A1(n1358), .A2(n1359), .ZN(n1354) );
NAND2_X1 U983 ( .A1(n1340), .A2(n1360), .ZN(n1359) );
INV_X1 U984 ( .A(KEYINPUT26), .ZN(n1360) );
NOR4_X1 U985 ( .A1(n1140), .A2(n1361), .A3(n1342), .A4(n1143), .ZN(n1340) );
NAND4_X1 U986 ( .A1(n1173), .A2(n1361), .A3(n1362), .A4(KEYINPUT26), .ZN(n1358) );
NOR2_X1 U987 ( .A1(n1342), .A2(n1140), .ZN(n1362) );
INV_X1 U988 ( .A(n1143), .ZN(n1173) );
AND2_X1 U989 ( .A1(n1149), .A2(n1161), .ZN(n1339) );
NAND2_X1 U990 ( .A1(n1363), .A2(n1364), .ZN(G30) );
NAND2_X1 U991 ( .A1(n1326), .A2(n1365), .ZN(n1364) );
XOR2_X1 U992 ( .A(KEYINPUT10), .B(n1366), .Z(n1363) );
NOR2_X1 U993 ( .A1(n1326), .A2(n1365), .ZN(n1366) );
AND2_X1 U994 ( .A1(n1344), .A2(n1131), .ZN(n1326) );
AND4_X1 U995 ( .A1(n1347), .A2(n1350), .A3(n1334), .A4(n1351), .ZN(n1344) );
NAND2_X1 U996 ( .A1(n1367), .A2(n1368), .ZN(G3) );
NAND2_X1 U997 ( .A1(G101), .A2(n1369), .ZN(n1368) );
XOR2_X1 U998 ( .A(KEYINPUT3), .B(n1370), .Z(n1367) );
NOR2_X1 U999 ( .A1(G101), .A2(n1369), .ZN(n1370) );
NAND3_X1 U1000 ( .A1(n1132), .A2(n1180), .A3(n1149), .ZN(n1369) );
XNOR2_X1 U1001 ( .A(n1224), .B(n1336), .ZN(G27) );
NOR2_X1 U1002 ( .A1(n1335), .A2(n1342), .ZN(n1336) );
INV_X1 U1003 ( .A(n1334), .ZN(n1342) );
NAND2_X1 U1004 ( .A1(n1154), .A2(n1371), .ZN(n1334) );
NAND3_X1 U1005 ( .A1(G902), .A2(n1372), .A3(n1211), .ZN(n1371) );
NOR2_X1 U1006 ( .A1(n1176), .A2(G900), .ZN(n1211) );
NAND4_X1 U1007 ( .A1(n1179), .A2(n1150), .A3(n1161), .A4(n1373), .ZN(n1335) );
NAND2_X1 U1008 ( .A1(n1374), .A2(n1375), .ZN(G24) );
OR3_X1 U1009 ( .A1(n1178), .A2(G122), .A3(n1314), .ZN(n1375) );
NAND2_X1 U1010 ( .A1(n1376), .A2(n1377), .ZN(n1374) );
XOR2_X1 U1011 ( .A(KEYINPUT48), .B(n1378), .Z(n1377) );
NOR2_X1 U1012 ( .A1(n1178), .A2(n1314), .ZN(n1378) );
NAND4_X1 U1013 ( .A1(n1345), .A2(n1319), .A3(n1134), .A4(n1379), .ZN(n1314) );
INV_X1 U1014 ( .A(n1348), .ZN(n1379) );
NOR2_X1 U1015 ( .A1(n1351), .A2(n1350), .ZN(n1134) );
XNOR2_X1 U1016 ( .A(G122), .B(KEYINPUT47), .ZN(n1376) );
XOR2_X1 U1017 ( .A(G119), .B(n1380), .Z(G21) );
NOR2_X1 U1018 ( .A1(n1178), .A2(n1308), .ZN(n1380) );
NAND4_X1 U1019 ( .A1(n1319), .A2(n1180), .A3(n1350), .A4(n1351), .ZN(n1308) );
XOR2_X1 U1020 ( .A(G116), .B(n1315), .Z(G18) );
AND2_X1 U1021 ( .A1(n1381), .A2(n1131), .ZN(n1315) );
XNOR2_X1 U1022 ( .A(n1382), .B(n1294), .ZN(G15) );
AND2_X1 U1023 ( .A1(n1381), .A2(n1161), .ZN(n1294) );
AND2_X1 U1024 ( .A1(n1345), .A2(n1383), .ZN(n1161) );
XNOR2_X1 U1025 ( .A(KEYINPUT50), .B(n1348), .ZN(n1383) );
AND3_X1 U1026 ( .A1(n1149), .A2(n1373), .A3(n1319), .ZN(n1381) );
NOR2_X1 U1027 ( .A1(n1159), .A2(n1311), .ZN(n1319) );
INV_X1 U1028 ( .A(n1179), .ZN(n1159) );
NOR2_X1 U1029 ( .A1(n1165), .A2(n1186), .ZN(n1179) );
NOR2_X1 U1030 ( .A1(n1351), .A2(n1183), .ZN(n1149) );
XNOR2_X1 U1031 ( .A(G110), .B(n1384), .ZN(G12) );
NAND2_X1 U1032 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
NAND2_X1 U1033 ( .A1(KEYINPUT16), .A2(n1321), .ZN(n1386) );
OR2_X1 U1034 ( .A1(KEYINPUT22), .A2(n1321), .ZN(n1385) );
AND3_X1 U1035 ( .A1(n1132), .A2(n1180), .A3(n1150), .ZN(n1321) );
INV_X1 U1036 ( .A(n1312), .ZN(n1150) );
NAND2_X1 U1037 ( .A1(n1183), .A2(n1351), .ZN(n1312) );
NAND2_X1 U1038 ( .A1(n1192), .A2(n1387), .ZN(n1351) );
NAND2_X1 U1039 ( .A1(n1193), .A2(n1194), .ZN(n1387) );
OR2_X1 U1040 ( .A1(n1194), .A2(n1193), .ZN(n1192) );
INV_X1 U1041 ( .A(n1242), .ZN(n1193) );
NAND2_X1 U1042 ( .A1(G217), .A2(n1388), .ZN(n1242) );
NAND2_X1 U1043 ( .A1(n1241), .A2(n1389), .ZN(n1194) );
XOR2_X1 U1044 ( .A(n1390), .B(n1391), .Z(n1241) );
XOR2_X1 U1045 ( .A(n1392), .B(n1393), .Z(n1391) );
NOR2_X1 U1046 ( .A1(n1394), .A2(n1395), .ZN(n1393) );
NOR3_X1 U1047 ( .A1(KEYINPUT7), .A2(G125), .A3(n1349), .ZN(n1395) );
NOR2_X1 U1048 ( .A1(n1396), .A2(n1397), .ZN(n1394) );
INV_X1 U1049 ( .A(KEYINPUT7), .ZN(n1397) );
XOR2_X1 U1050 ( .A(n1398), .B(n1399), .Z(n1390) );
XNOR2_X1 U1051 ( .A(G137), .B(n1400), .ZN(n1399) );
NAND2_X1 U1052 ( .A1(n1401), .A2(n1402), .ZN(n1400) );
OR2_X1 U1053 ( .A1(n1403), .A2(G110), .ZN(n1402) );
XOR2_X1 U1054 ( .A(n1404), .B(KEYINPUT29), .Z(n1401) );
NAND2_X1 U1055 ( .A1(G110), .A2(n1403), .ZN(n1404) );
XNOR2_X1 U1056 ( .A(G119), .B(n1365), .ZN(n1403) );
NAND4_X1 U1057 ( .A1(KEYINPUT43), .A2(G221), .A3(G234), .A4(n1176), .ZN(n1398) );
INV_X1 U1058 ( .A(n1350), .ZN(n1183) );
XNOR2_X1 U1059 ( .A(n1405), .B(G472), .ZN(n1350) );
NAND2_X1 U1060 ( .A1(n1406), .A2(n1389), .ZN(n1405) );
XOR2_X1 U1061 ( .A(n1407), .B(n1408), .Z(n1406) );
XNOR2_X1 U1062 ( .A(n1409), .B(n1259), .ZN(n1408) );
XNOR2_X1 U1063 ( .A(n1410), .B(G101), .ZN(n1259) );
NAND2_X1 U1064 ( .A1(G210), .A2(n1411), .ZN(n1410) );
NAND2_X1 U1065 ( .A1(KEYINPUT6), .A2(n1264), .ZN(n1409) );
XOR2_X1 U1066 ( .A(G113), .B(n1412), .Z(n1264) );
NAND2_X1 U1067 ( .A1(n1413), .A2(n1414), .ZN(n1407) );
NAND2_X1 U1068 ( .A1(n1265), .A2(n1415), .ZN(n1414) );
INV_X1 U1069 ( .A(KEYINPUT40), .ZN(n1415) );
XNOR2_X1 U1070 ( .A(n1282), .B(n1416), .ZN(n1265) );
NAND3_X1 U1071 ( .A1(n1275), .A2(n1282), .A3(KEYINPUT40), .ZN(n1413) );
NAND2_X1 U1072 ( .A1(n1417), .A2(n1418), .ZN(n1180) );
OR2_X1 U1073 ( .A1(n1162), .A2(KEYINPUT50), .ZN(n1418) );
INV_X1 U1074 ( .A(n1131), .ZN(n1162) );
NOR2_X1 U1075 ( .A1(n1345), .A2(n1348), .ZN(n1131) );
INV_X1 U1076 ( .A(n1419), .ZN(n1345) );
NAND3_X1 U1077 ( .A1(n1419), .A2(n1348), .A3(KEYINPUT50), .ZN(n1417) );
XNOR2_X1 U1078 ( .A(G478), .B(n1195), .ZN(n1348) );
NOR2_X1 U1079 ( .A1(n1247), .A2(G902), .ZN(n1195) );
NAND3_X1 U1080 ( .A1(n1420), .A2(n1421), .A3(n1422), .ZN(n1247) );
OR2_X1 U1081 ( .A1(n1423), .A2(KEYINPUT33), .ZN(n1422) );
NAND4_X1 U1082 ( .A1(KEYINPUT46), .A2(n1423), .A3(KEYINPUT33), .A4(n1424), .ZN(n1421) );
INV_X1 U1083 ( .A(n1425), .ZN(n1424) );
NAND2_X1 U1084 ( .A1(n1425), .A2(n1426), .ZN(n1420) );
NAND2_X1 U1085 ( .A1(KEYINPUT46), .A2(n1423), .ZN(n1426) );
AND3_X1 U1086 ( .A1(G217), .A2(n1176), .A3(G234), .ZN(n1423) );
XNOR2_X1 U1087 ( .A(n1427), .B(n1428), .ZN(n1425) );
XOR2_X1 U1088 ( .A(G116), .B(n1429), .Z(n1428) );
XOR2_X1 U1089 ( .A(KEYINPUT24), .B(G122), .Z(n1429) );
XOR2_X1 U1090 ( .A(n1430), .B(n1431), .Z(n1427) );
XNOR2_X1 U1091 ( .A(G107), .B(n1432), .ZN(n1431) );
NAND2_X1 U1092 ( .A1(n1433), .A2(n1434), .ZN(n1432) );
XNOR2_X1 U1093 ( .A(n1435), .B(KEYINPUT58), .ZN(n1433) );
NAND2_X1 U1094 ( .A1(KEYINPUT44), .A2(G134), .ZN(n1430) );
XNOR2_X1 U1095 ( .A(n1182), .B(KEYINPUT61), .ZN(n1419) );
XOR2_X1 U1096 ( .A(n1436), .B(G475), .Z(n1182) );
NAND2_X1 U1097 ( .A1(n1437), .A2(n1389), .ZN(n1436) );
XNOR2_X1 U1098 ( .A(n1255), .B(KEYINPUT55), .ZN(n1437) );
XNOR2_X1 U1099 ( .A(n1438), .B(n1439), .ZN(n1255) );
XOR2_X1 U1100 ( .A(n1396), .B(n1440), .Z(n1439) );
XNOR2_X1 U1101 ( .A(n1224), .B(G140), .ZN(n1396) );
INV_X1 U1102 ( .A(G125), .ZN(n1224) );
XOR2_X1 U1103 ( .A(n1441), .B(n1392), .Z(n1438) );
XNOR2_X1 U1104 ( .A(G104), .B(n1442), .ZN(n1441) );
NOR2_X1 U1105 ( .A1(KEYINPUT53), .A2(n1443), .ZN(n1442) );
NOR2_X1 U1106 ( .A1(n1444), .A2(n1445), .ZN(n1443) );
XOR2_X1 U1107 ( .A(n1446), .B(KEYINPUT42), .Z(n1445) );
NAND2_X1 U1108 ( .A1(G131), .A2(n1447), .ZN(n1446) );
NOR2_X1 U1109 ( .A1(G131), .A2(n1447), .ZN(n1444) );
XOR2_X1 U1110 ( .A(n1448), .B(G143), .Z(n1447) );
NAND2_X1 U1111 ( .A1(G214), .A2(n1411), .ZN(n1448) );
NOR2_X1 U1112 ( .A1(G953), .A2(G237), .ZN(n1411) );
NOR2_X1 U1113 ( .A1(n1301), .A2(n1311), .ZN(n1132) );
INV_X1 U1114 ( .A(n1302), .ZN(n1311) );
NAND2_X1 U1115 ( .A1(n1154), .A2(n1449), .ZN(n1302) );
NAND3_X1 U1116 ( .A1(G902), .A2(n1372), .A3(n1232), .ZN(n1449) );
NOR2_X1 U1117 ( .A1(n1176), .A2(G898), .ZN(n1232) );
NAND3_X1 U1118 ( .A1(n1372), .A2(n1176), .A3(G952), .ZN(n1154) );
NAND2_X1 U1119 ( .A1(G237), .A2(G234), .ZN(n1372) );
INV_X1 U1120 ( .A(n1347), .ZN(n1301) );
NOR2_X1 U1121 ( .A1(n1361), .A2(n1178), .ZN(n1347) );
INV_X1 U1122 ( .A(n1373), .ZN(n1178) );
NOR2_X1 U1123 ( .A1(n1199), .A2(n1143), .ZN(n1373) );
NOR2_X1 U1124 ( .A1(n1450), .A2(n1288), .ZN(n1143) );
INV_X1 U1125 ( .A(G214), .ZN(n1450) );
INV_X1 U1126 ( .A(n1140), .ZN(n1199) );
XNOR2_X1 U1127 ( .A(n1451), .B(n1452), .ZN(n1140) );
NOR2_X1 U1128 ( .A1(n1288), .A2(n1289), .ZN(n1452) );
INV_X1 U1129 ( .A(G210), .ZN(n1289) );
NOR2_X1 U1130 ( .A1(n1453), .A2(G237), .ZN(n1288) );
NAND2_X1 U1131 ( .A1(n1454), .A2(n1389), .ZN(n1451) );
XOR2_X1 U1132 ( .A(n1455), .B(n1456), .Z(n1454) );
XNOR2_X1 U1133 ( .A(G125), .B(n1457), .ZN(n1456) );
NAND2_X1 U1134 ( .A1(KEYINPUT27), .A2(n1286), .ZN(n1457) );
AND2_X1 U1135 ( .A1(G224), .A2(n1176), .ZN(n1286) );
XNOR2_X1 U1136 ( .A(n1234), .B(n1282), .ZN(n1455) );
XNOR2_X1 U1137 ( .A(n1458), .B(n1459), .ZN(n1282) );
NOR2_X1 U1138 ( .A1(n1435), .A2(n1460), .ZN(n1459) );
INV_X1 U1139 ( .A(n1434), .ZN(n1460) );
NAND2_X1 U1140 ( .A1(KEYINPUT54), .A2(n1392), .ZN(n1458) );
XNOR2_X1 U1141 ( .A(n1461), .B(n1462), .ZN(n1234) );
XOR2_X1 U1142 ( .A(n1463), .B(n1464), .Z(n1462) );
XNOR2_X1 U1143 ( .A(n1465), .B(G104), .ZN(n1464) );
XNOR2_X1 U1144 ( .A(KEYINPUT30), .B(n1466), .ZN(n1463) );
INV_X1 U1145 ( .A(G110), .ZN(n1466) );
XOR2_X1 U1146 ( .A(n1467), .B(n1440), .Z(n1461) );
XNOR2_X1 U1147 ( .A(n1382), .B(G122), .ZN(n1440) );
INV_X1 U1148 ( .A(G113), .ZN(n1382) );
XNOR2_X1 U1149 ( .A(G101), .B(n1412), .ZN(n1467) );
XOR2_X1 U1150 ( .A(G116), .B(G119), .Z(n1412) );
INV_X1 U1151 ( .A(n1313), .ZN(n1361) );
NOR2_X1 U1152 ( .A1(n1468), .A2(n1186), .ZN(n1313) );
INV_X1 U1153 ( .A(n1163), .ZN(n1186) );
NAND2_X1 U1154 ( .A1(G221), .A2(n1388), .ZN(n1163) );
NAND2_X1 U1155 ( .A1(G234), .A2(n1469), .ZN(n1388) );
INV_X1 U1156 ( .A(n1453), .ZN(n1469) );
XOR2_X1 U1157 ( .A(n1389), .B(KEYINPUT59), .Z(n1453) );
INV_X1 U1158 ( .A(n1165), .ZN(n1468) );
XNOR2_X1 U1159 ( .A(n1200), .B(G469), .ZN(n1165) );
NAND2_X1 U1160 ( .A1(n1470), .A2(n1389), .ZN(n1200) );
INV_X1 U1161 ( .A(G902), .ZN(n1389) );
XNOR2_X1 U1162 ( .A(n1276), .B(n1471), .ZN(n1470) );
XNOR2_X1 U1163 ( .A(n1472), .B(n1349), .ZN(n1471) );
INV_X1 U1164 ( .A(G140), .ZN(n1349) );
NAND2_X1 U1165 ( .A1(n1473), .A2(n1474), .ZN(n1472) );
NAND2_X1 U1166 ( .A1(n1416), .A2(n1274), .ZN(n1474) );
XOR2_X1 U1167 ( .A(KEYINPUT38), .B(n1475), .Z(n1473) );
NOR2_X1 U1168 ( .A1(n1416), .A2(n1274), .ZN(n1475) );
XNOR2_X1 U1169 ( .A(n1476), .B(n1477), .ZN(n1274) );
XNOR2_X1 U1170 ( .A(n1478), .B(n1215), .ZN(n1477) );
XNOR2_X1 U1171 ( .A(n1479), .B(n1392), .ZN(n1215) );
XOR2_X1 U1172 ( .A(G146), .B(KEYINPUT60), .Z(n1392) );
NAND3_X1 U1173 ( .A1(n1480), .A2(n1481), .A3(n1434), .ZN(n1479) );
NAND2_X1 U1174 ( .A1(G143), .A2(n1365), .ZN(n1434) );
OR2_X1 U1175 ( .A1(G128), .A2(KEYINPUT11), .ZN(n1481) );
NAND2_X1 U1176 ( .A1(n1435), .A2(KEYINPUT11), .ZN(n1480) );
NOR2_X1 U1177 ( .A1(n1365), .A2(G143), .ZN(n1435) );
INV_X1 U1178 ( .A(G128), .ZN(n1365) );
NAND2_X1 U1179 ( .A1(KEYINPUT12), .A2(n1465), .ZN(n1478) );
INV_X1 U1180 ( .A(G107), .ZN(n1465) );
XNOR2_X1 U1181 ( .A(G101), .B(G104), .ZN(n1476) );
INV_X1 U1182 ( .A(n1275), .ZN(n1416) );
XOR2_X1 U1183 ( .A(G131), .B(n1219), .Z(n1275) );
XOR2_X1 U1184 ( .A(G134), .B(G137), .Z(n1219) );
XOR2_X1 U1185 ( .A(G110), .B(n1482), .Z(n1276) );
AND2_X1 U1186 ( .A1(n1176), .A2(G227), .ZN(n1482) );
INV_X1 U1187 ( .A(G953), .ZN(n1176) );
endmodule


