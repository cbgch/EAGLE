//Key = 0101011101111010000100011101000111110001011100100100101000101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341;

XOR2_X1 U729 ( .A(G107), .B(n1015), .Z(G9) );
NOR2_X1 U730 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U731 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
NAND4_X1 U732 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1018) );
NAND2_X1 U733 ( .A1(n1026), .A2(n1027), .ZN(n1023) );
NAND2_X1 U734 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND3_X1 U735 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NAND2_X1 U736 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NAND2_X1 U737 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
OR2_X1 U738 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U739 ( .A1(n1039), .A2(n1040), .ZN(n1033) );
NAND2_X1 U740 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U741 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
INV_X1 U742 ( .A(n1045), .ZN(n1041) );
NAND3_X1 U743 ( .A1(n1035), .A2(n1046), .A3(n1039), .ZN(n1028) );
NAND2_X1 U744 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U745 ( .A1(n1032), .A2(n1049), .ZN(n1048) );
NAND2_X1 U746 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U747 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XOR2_X1 U748 ( .A(KEYINPUT26), .B(n1054), .Z(n1052) );
NAND2_X1 U749 ( .A1(KEYINPUT43), .A2(n1055), .ZN(n1050) );
NAND2_X1 U750 ( .A1(n1030), .A2(n1056), .ZN(n1047) );
NAND2_X1 U751 ( .A1(n1057), .A2(n1058), .ZN(n1022) );
INV_X1 U752 ( .A(KEYINPUT43), .ZN(n1058) );
NAND3_X1 U753 ( .A1(n1026), .A2(n1039), .A3(n1059), .ZN(n1057) );
NOR3_X1 U754 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
INV_X1 U755 ( .A(n1063), .ZN(n1026) );
NOR3_X1 U756 ( .A1(n1064), .A2(G953), .A3(n1065), .ZN(n1016) );
INV_X1 U757 ( .A(n1024), .ZN(n1065) );
NAND4_X1 U758 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1024) );
NOR3_X1 U759 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
XOR2_X1 U760 ( .A(n1073), .B(n1074), .Z(n1072) );
XOR2_X1 U761 ( .A(G475), .B(n1075), .Z(n1071) );
NAND3_X1 U762 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1070) );
XOR2_X1 U763 ( .A(n1079), .B(G472), .Z(n1078) );
NAND2_X1 U764 ( .A1(n1080), .A2(n1081), .ZN(n1077) );
INV_X1 U765 ( .A(KEYINPUT9), .ZN(n1081) );
NAND2_X1 U766 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
XNOR2_X1 U767 ( .A(n1084), .B(KEYINPUT34), .ZN(n1082) );
NAND2_X1 U768 ( .A1(KEYINPUT9), .A2(n1085), .ZN(n1076) );
NAND2_X1 U769 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
OR2_X1 U770 ( .A1(n1084), .A2(KEYINPUT34), .ZN(n1087) );
NAND3_X1 U771 ( .A1(n1084), .A2(n1083), .A3(KEYINPUT34), .ZN(n1086) );
NOR3_X1 U772 ( .A1(n1088), .A2(n1053), .A3(n1044), .ZN(n1068) );
XOR2_X1 U773 ( .A(n1089), .B(n1090), .Z(n1066) );
NOR2_X1 U774 ( .A1(KEYINPUT44), .A2(n1091), .ZN(n1090) );
XOR2_X1 U775 ( .A(n1020), .B(KEYINPUT42), .Z(n1064) );
INV_X1 U776 ( .A(G952), .ZN(n1020) );
XOR2_X1 U777 ( .A(n1092), .B(n1093), .Z(G72) );
NAND2_X1 U778 ( .A1(G953), .A2(n1094), .ZN(n1093) );
NAND2_X1 U779 ( .A1(G900), .A2(G227), .ZN(n1094) );
NAND2_X1 U780 ( .A1(KEYINPUT7), .A2(n1095), .ZN(n1092) );
XOR2_X1 U781 ( .A(n1096), .B(n1097), .Z(n1095) );
AND2_X1 U782 ( .A1(n1019), .A2(n1025), .ZN(n1097) );
NOR2_X1 U783 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
XNOR2_X1 U784 ( .A(n1100), .B(n1101), .ZN(n1099) );
XOR2_X1 U785 ( .A(n1102), .B(n1103), .Z(G69) );
XOR2_X1 U786 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U787 ( .A1(n1106), .A2(n1025), .ZN(n1105) );
AND2_X1 U788 ( .A1(G224), .A2(G898), .ZN(n1106) );
NAND3_X1 U789 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1104) );
NAND2_X1 U790 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U791 ( .A1(n1112), .A2(n1113), .ZN(n1108) );
NAND2_X1 U792 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U793 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U794 ( .A1(n1118), .A2(n1119), .ZN(n1107) );
INV_X1 U795 ( .A(n1112), .ZN(n1119) );
XOR2_X1 U796 ( .A(n1116), .B(n1117), .Z(n1118) );
INV_X1 U797 ( .A(n1120), .ZN(n1117) );
NAND2_X1 U798 ( .A1(n1025), .A2(n1021), .ZN(n1102) );
NOR2_X1 U799 ( .A1(n1121), .A2(n1122), .ZN(G66) );
XOR2_X1 U800 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR3_X1 U801 ( .A1(n1125), .A2(KEYINPUT59), .A3(n1126), .ZN(n1123) );
NOR2_X1 U802 ( .A1(n1121), .A2(n1127), .ZN(G63) );
XOR2_X1 U803 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND2_X1 U804 ( .A1(KEYINPUT5), .A2(n1130), .ZN(n1128) );
NAND2_X1 U805 ( .A1(n1131), .A2(G478), .ZN(n1130) );
NOR2_X1 U806 ( .A1(n1121), .A2(n1132), .ZN(G60) );
XOR2_X1 U807 ( .A(n1133), .B(n1134), .Z(n1132) );
AND2_X1 U808 ( .A1(G475), .A2(n1131), .ZN(n1133) );
XOR2_X1 U809 ( .A(G104), .B(n1135), .Z(G6) );
NOR3_X1 U810 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(G57) );
NOR2_X1 U811 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XNOR2_X1 U812 ( .A(n1141), .B(KEYINPUT29), .ZN(n1140) );
XOR2_X1 U813 ( .A(n1142), .B(KEYINPUT2), .Z(n1139) );
NOR2_X1 U814 ( .A1(n1141), .A2(n1143), .ZN(n1137) );
XNOR2_X1 U815 ( .A(KEYINPUT2), .B(n1142), .ZN(n1143) );
XNOR2_X1 U816 ( .A(n1144), .B(n1145), .ZN(n1141) );
NOR2_X1 U817 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U818 ( .A(n1148), .B(KEYINPUT31), .Z(n1147) );
NAND2_X1 U819 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U820 ( .A1(n1149), .A2(n1150), .ZN(n1146) );
AND2_X1 U821 ( .A1(n1131), .A2(G472), .ZN(n1149) );
INV_X1 U822 ( .A(n1125), .ZN(n1131) );
NOR2_X1 U823 ( .A1(n1025), .A2(n1151), .ZN(n1136) );
XOR2_X1 U824 ( .A(KEYINPUT13), .B(G952), .Z(n1151) );
NOR2_X1 U825 ( .A1(n1121), .A2(n1152), .ZN(G54) );
XOR2_X1 U826 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U827 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U828 ( .A(n1157), .B(n1100), .Z(n1156) );
NOR2_X1 U829 ( .A1(n1073), .A2(n1125), .ZN(n1157) );
INV_X1 U830 ( .A(G469), .ZN(n1073) );
XNOR2_X1 U831 ( .A(n1158), .B(n1159), .ZN(n1153) );
XOR2_X1 U832 ( .A(KEYINPUT3), .B(n1160), .Z(n1159) );
NOR2_X1 U833 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XOR2_X1 U834 ( .A(n1163), .B(KEYINPUT25), .Z(n1162) );
NAND2_X1 U835 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XOR2_X1 U836 ( .A(KEYINPUT0), .B(G140), .Z(n1164) );
INV_X1 U837 ( .A(n1166), .ZN(n1161) );
NOR2_X1 U838 ( .A1(n1121), .A2(n1167), .ZN(G51) );
XOR2_X1 U839 ( .A(n1168), .B(n1169), .Z(n1167) );
XNOR2_X1 U840 ( .A(n1170), .B(n1171), .ZN(n1169) );
XOR2_X1 U841 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U842 ( .A1(n1091), .A2(n1125), .ZN(n1173) );
NAND2_X1 U843 ( .A1(G902), .A2(n1174), .ZN(n1125) );
OR2_X1 U844 ( .A1(n1019), .A2(n1021), .ZN(n1174) );
NAND3_X1 U845 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1021) );
NOR3_X1 U846 ( .A1(n1015), .A2(n1178), .A3(n1135), .ZN(n1177) );
AND3_X1 U847 ( .A1(n1179), .A2(n1032), .A3(n1037), .ZN(n1135) );
AND3_X1 U848 ( .A1(n1038), .A2(n1032), .A3(n1179), .ZN(n1015) );
NAND3_X1 U849 ( .A1(n1179), .A2(n1056), .A3(n1039), .ZN(n1176) );
NAND2_X1 U850 ( .A1(n1180), .A2(n1181), .ZN(n1056) );
NAND2_X1 U851 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
INV_X1 U852 ( .A(n1184), .ZN(n1179) );
NAND2_X1 U853 ( .A1(n1185), .A2(n1186), .ZN(n1175) );
NAND2_X1 U854 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND4_X1 U855 ( .A1(n1032), .A2(n1055), .A3(n1189), .A4(n1190), .ZN(n1188) );
INV_X1 U856 ( .A(n1062), .ZN(n1032) );
NAND2_X1 U857 ( .A1(n1191), .A2(n1192), .ZN(n1187) );
NAND2_X1 U858 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NAND2_X1 U859 ( .A1(n1038), .A2(n1195), .ZN(n1194) );
XOR2_X1 U860 ( .A(KEYINPUT8), .B(n1055), .Z(n1195) );
NAND2_X1 U861 ( .A1(n1037), .A2(n1196), .ZN(n1193) );
NAND4_X1 U862 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1019) );
AND4_X1 U863 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
NOR2_X1 U864 ( .A1(n1205), .A2(n1206), .ZN(n1199) );
NOR2_X1 U865 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NOR2_X1 U866 ( .A1(KEYINPUT48), .A2(n1209), .ZN(n1172) );
XOR2_X1 U867 ( .A(n1210), .B(n1211), .Z(n1168) );
XOR2_X1 U868 ( .A(KEYINPUT20), .B(G125), .Z(n1211) );
NOR2_X1 U869 ( .A1(n1025), .A2(G952), .ZN(n1121) );
XOR2_X1 U870 ( .A(G146), .B(n1205), .Z(G48) );
AND4_X1 U871 ( .A1(n1045), .A2(n1037), .A3(n1212), .A4(n1213), .ZN(n1205) );
XNOR2_X1 U872 ( .A(G143), .B(n1197), .ZN(G45) );
NAND4_X1 U873 ( .A1(n1045), .A2(n1055), .A3(n1191), .A4(n1214), .ZN(n1197) );
AND3_X1 U874 ( .A1(n1189), .A2(n1190), .A3(n1215), .ZN(n1214) );
XOR2_X1 U875 ( .A(n1216), .B(n1198), .Z(G42) );
NAND4_X1 U876 ( .A1(n1217), .A2(n1037), .A3(n1182), .A4(n1183), .ZN(n1198) );
XOR2_X1 U877 ( .A(G137), .B(n1218), .Z(G39) );
NOR3_X1 U878 ( .A1(n1208), .A2(KEYINPUT22), .A3(n1207), .ZN(n1218) );
XNOR2_X1 U879 ( .A(G134), .B(n1204), .ZN(G36) );
NAND3_X1 U880 ( .A1(n1191), .A2(n1038), .A3(n1217), .ZN(n1204) );
XOR2_X1 U881 ( .A(n1203), .B(n1219), .Z(G33) );
NAND2_X1 U882 ( .A1(KEYINPUT54), .A2(G131), .ZN(n1219) );
NAND3_X1 U883 ( .A1(n1191), .A2(n1037), .A3(n1217), .ZN(n1203) );
INV_X1 U884 ( .A(n1207), .ZN(n1217) );
NAND3_X1 U885 ( .A1(n1030), .A2(n1215), .A3(n1045), .ZN(n1207) );
XNOR2_X1 U886 ( .A(n1220), .B(KEYINPUT10), .ZN(n1045) );
NAND2_X1 U887 ( .A1(n1221), .A2(n1222), .ZN(n1030) );
OR3_X1 U888 ( .A1(n1223), .A2(n1053), .A3(KEYINPUT26), .ZN(n1222) );
INV_X1 U889 ( .A(n1054), .ZN(n1223) );
NAND2_X1 U890 ( .A1(KEYINPUT26), .A2(n1055), .ZN(n1221) );
XNOR2_X1 U891 ( .A(G128), .B(n1202), .ZN(G30) );
NAND4_X1 U892 ( .A1(n1212), .A2(n1038), .A3(n1220), .A4(n1213), .ZN(n1202) );
XOR2_X1 U893 ( .A(G101), .B(n1224), .Z(G3) );
NOR4_X1 U894 ( .A1(KEYINPUT18), .A2(n1184), .A3(n1180), .A4(n1225), .ZN(n1224) );
XOR2_X1 U895 ( .A(G125), .B(n1226), .Z(G27) );
NOR2_X1 U896 ( .A1(KEYINPUT36), .A2(n1201), .ZN(n1226) );
NAND4_X1 U897 ( .A1(n1035), .A2(n1037), .A3(n1182), .A4(n1212), .ZN(n1201) );
AND3_X1 U898 ( .A1(n1183), .A2(n1215), .A3(n1055), .ZN(n1212) );
NAND2_X1 U899 ( .A1(n1063), .A2(n1227), .ZN(n1215) );
NAND3_X1 U900 ( .A1(G902), .A2(n1228), .A3(n1098), .ZN(n1227) );
NOR2_X1 U901 ( .A1(n1229), .A2(G900), .ZN(n1098) );
INV_X1 U902 ( .A(n1110), .ZN(n1229) );
XOR2_X1 U903 ( .A(n1230), .B(n1231), .Z(G24) );
NOR2_X1 U904 ( .A1(KEYINPUT15), .A2(n1232), .ZN(n1231) );
NOR4_X1 U905 ( .A1(n1233), .A2(n1234), .A3(n1062), .A4(n1235), .ZN(n1232) );
NAND2_X1 U906 ( .A1(n1067), .A2(n1182), .ZN(n1062) );
NAND2_X1 U907 ( .A1(n1189), .A2(n1190), .ZN(n1234) );
XOR2_X1 U908 ( .A(n1061), .B(KEYINPUT53), .Z(n1233) );
XOR2_X1 U909 ( .A(G119), .B(n1178), .Z(G21) );
NOR3_X1 U910 ( .A1(n1208), .A2(n1061), .A3(n1235), .ZN(n1178) );
NAND3_X1 U911 ( .A1(n1213), .A2(n1183), .A3(n1039), .ZN(n1208) );
INV_X1 U912 ( .A(n1067), .ZN(n1183) );
XNOR2_X1 U913 ( .A(G116), .B(n1236), .ZN(G18) );
NAND4_X1 U914 ( .A1(n1185), .A2(n1191), .A3(n1038), .A4(n1055), .ZN(n1236) );
NOR2_X1 U915 ( .A1(n1237), .A2(n1238), .ZN(n1038) );
INV_X1 U916 ( .A(n1190), .ZN(n1238) );
INV_X1 U917 ( .A(n1235), .ZN(n1185) );
XOR2_X1 U918 ( .A(n1239), .B(n1240), .Z(G15) );
NAND4_X1 U919 ( .A1(n1241), .A2(n1191), .A3(n1196), .A4(n1037), .ZN(n1240) );
NOR2_X1 U920 ( .A1(n1190), .A2(n1242), .ZN(n1037) );
INV_X1 U921 ( .A(n1180), .ZN(n1191) );
NAND2_X1 U922 ( .A1(n1067), .A2(n1213), .ZN(n1180) );
NOR2_X1 U923 ( .A1(n1243), .A2(n1244), .ZN(n1241) );
NOR2_X1 U924 ( .A1(KEYINPUT33), .A2(n1245), .ZN(n1244) );
NOR2_X1 U925 ( .A1(n1060), .A2(n1246), .ZN(n1245) );
AND2_X1 U926 ( .A1(n1235), .A2(KEYINPUT33), .ZN(n1243) );
NAND2_X1 U927 ( .A1(n1035), .A2(n1246), .ZN(n1235) );
INV_X1 U928 ( .A(n1060), .ZN(n1035) );
NAND2_X1 U929 ( .A1(n1043), .A2(n1247), .ZN(n1060) );
XOR2_X1 U930 ( .A(G110), .B(n1248), .Z(G12) );
NOR4_X1 U931 ( .A1(n1067), .A2(n1249), .A3(n1184), .A4(n1213), .ZN(n1248) );
INV_X1 U932 ( .A(n1182), .ZN(n1213) );
XNOR2_X1 U933 ( .A(n1250), .B(n1079), .ZN(n1182) );
NAND2_X1 U934 ( .A1(n1251), .A2(n1252), .ZN(n1079) );
XOR2_X1 U935 ( .A(n1253), .B(n1254), .Z(n1251) );
XNOR2_X1 U936 ( .A(n1142), .B(n1255), .ZN(n1254) );
NOR2_X1 U937 ( .A1(KEYINPUT16), .A2(n1256), .ZN(n1255) );
INV_X1 U938 ( .A(n1150), .ZN(n1256) );
XOR2_X1 U939 ( .A(n1257), .B(n1258), .Z(n1150) );
XNOR2_X1 U940 ( .A(n1259), .B(KEYINPUT57), .ZN(n1258) );
NAND2_X1 U941 ( .A1(KEYINPUT62), .A2(n1239), .ZN(n1259) );
XNOR2_X1 U942 ( .A(n1100), .B(n1260), .ZN(n1257) );
XOR2_X1 U943 ( .A(n1261), .B(n1262), .Z(n1100) );
NAND2_X1 U944 ( .A1(n1263), .A2(G210), .ZN(n1142) );
XOR2_X1 U945 ( .A(n1144), .B(KEYINPUT1), .Z(n1253) );
NAND2_X1 U946 ( .A1(KEYINPUT19), .A2(G472), .ZN(n1250) );
NAND3_X1 U947 ( .A1(n1196), .A2(n1246), .A3(n1220), .ZN(n1184) );
NOR2_X1 U948 ( .A1(n1264), .A2(n1043), .ZN(n1220) );
XOR2_X1 U949 ( .A(n1265), .B(G469), .Z(n1043) );
NAND2_X1 U950 ( .A1(KEYINPUT6), .A2(n1266), .ZN(n1265) );
XNOR2_X1 U951 ( .A(KEYINPUT37), .B(n1074), .ZN(n1266) );
NAND2_X1 U952 ( .A1(n1267), .A2(n1252), .ZN(n1074) );
XOR2_X1 U953 ( .A(n1268), .B(n1269), .Z(n1267) );
NOR2_X1 U954 ( .A1(KEYINPUT56), .A2(n1270), .ZN(n1269) );
XOR2_X1 U955 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U956 ( .A(n1158), .B(KEYINPUT50), .Z(n1272) );
NAND2_X1 U957 ( .A1(G227), .A2(n1025), .ZN(n1158) );
NAND2_X1 U958 ( .A1(n1273), .A2(n1166), .ZN(n1271) );
NAND2_X1 U959 ( .A1(G110), .A2(n1216), .ZN(n1166) );
XOR2_X1 U960 ( .A(n1274), .B(KEYINPUT28), .Z(n1273) );
NAND2_X1 U961 ( .A1(G140), .A2(n1165), .ZN(n1274) );
NAND2_X1 U962 ( .A1(n1275), .A2(n1276), .ZN(n1268) );
NAND2_X1 U963 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND2_X1 U964 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
OR2_X1 U965 ( .A1(n1261), .A2(KEYINPUT4), .ZN(n1280) );
INV_X1 U966 ( .A(KEYINPUT38), .ZN(n1279) );
NAND2_X1 U967 ( .A1(n1261), .A2(n1281), .ZN(n1275) );
NAND2_X1 U968 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
OR2_X1 U969 ( .A1(n1277), .A2(KEYINPUT38), .ZN(n1283) );
XNOR2_X1 U970 ( .A(n1262), .B(n1155), .ZN(n1277) );
XNOR2_X1 U971 ( .A(n1284), .B(n1285), .ZN(n1155) );
XOR2_X1 U972 ( .A(G107), .B(n1286), .Z(n1285) );
NOR2_X1 U973 ( .A1(KEYINPUT21), .A2(n1144), .ZN(n1286) );
INV_X1 U974 ( .A(G101), .ZN(n1144) );
NAND2_X1 U975 ( .A1(KEYINPUT39), .A2(n1287), .ZN(n1284) );
INV_X1 U976 ( .A(KEYINPUT4), .ZN(n1282) );
XNOR2_X1 U977 ( .A(G131), .B(n1288), .ZN(n1261) );
XOR2_X1 U978 ( .A(G137), .B(G134), .Z(n1288) );
XOR2_X1 U979 ( .A(n1247), .B(KEYINPUT24), .Z(n1264) );
XOR2_X1 U980 ( .A(n1044), .B(KEYINPUT41), .Z(n1247) );
AND2_X1 U981 ( .A1(G221), .A2(n1289), .ZN(n1044) );
NAND2_X1 U982 ( .A1(n1063), .A2(n1290), .ZN(n1246) );
NAND4_X1 U983 ( .A1(n1110), .A2(G902), .A3(n1228), .A4(n1111), .ZN(n1290) );
INV_X1 U984 ( .A(G898), .ZN(n1111) );
XOR2_X1 U985 ( .A(n1025), .B(KEYINPUT23), .Z(n1110) );
NAND3_X1 U986 ( .A1(n1228), .A2(n1025), .A3(G952), .ZN(n1063) );
NAND2_X1 U987 ( .A1(G237), .A2(G234), .ZN(n1228) );
XOR2_X1 U988 ( .A(n1061), .B(KEYINPUT49), .Z(n1196) );
INV_X1 U989 ( .A(n1055), .ZN(n1061) );
NOR2_X1 U990 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
AND2_X1 U991 ( .A1(n1291), .A2(G214), .ZN(n1053) );
XOR2_X1 U992 ( .A(n1292), .B(KEYINPUT47), .Z(n1291) );
XNOR2_X1 U993 ( .A(n1089), .B(n1091), .ZN(n1054) );
NAND2_X1 U994 ( .A1(G210), .A2(n1292), .ZN(n1091) );
NAND2_X1 U995 ( .A1(n1252), .A2(n1293), .ZN(n1292) );
INV_X1 U996 ( .A(G237), .ZN(n1293) );
NAND2_X1 U997 ( .A1(n1294), .A2(n1252), .ZN(n1089) );
XOR2_X1 U998 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U999 ( .A(n1209), .B(n1170), .Z(n1296) );
XNOR2_X1 U1000 ( .A(n1297), .B(n1298), .ZN(n1170) );
NOR2_X1 U1001 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XOR2_X1 U1002 ( .A(KEYINPUT45), .B(n1301), .Z(n1300) );
NOR2_X1 U1003 ( .A1(n1120), .A2(n1302), .ZN(n1301) );
XOR2_X1 U1004 ( .A(KEYINPUT40), .B(n1303), .Z(n1302) );
INV_X1 U1005 ( .A(n1114), .ZN(n1299) );
NAND2_X1 U1006 ( .A1(n1120), .A2(n1303), .ZN(n1114) );
INV_X1 U1007 ( .A(n1116), .ZN(n1303) );
XOR2_X1 U1008 ( .A(n1304), .B(n1305), .Z(n1116) );
XOR2_X1 U1009 ( .A(KEYINPUT63), .B(G101), .Z(n1305) );
NAND2_X1 U1010 ( .A1(n1306), .A2(n1307), .ZN(n1304) );
NAND2_X1 U1011 ( .A1(G107), .A2(n1287), .ZN(n1307) );
XOR2_X1 U1012 ( .A(KEYINPUT12), .B(n1308), .Z(n1306) );
NOR2_X1 U1013 ( .A1(G107), .A2(n1287), .ZN(n1308) );
INV_X1 U1014 ( .A(G104), .ZN(n1287) );
XOR2_X1 U1015 ( .A(n1309), .B(n1260), .Z(n1120) );
XOR2_X1 U1016 ( .A(G116), .B(G119), .Z(n1260) );
XOR2_X1 U1017 ( .A(n1239), .B(KEYINPUT46), .Z(n1309) );
INV_X1 U1018 ( .A(G113), .ZN(n1239) );
NAND2_X1 U1019 ( .A1(KEYINPUT14), .A2(n1112), .ZN(n1297) );
XNOR2_X1 U1020 ( .A(n1230), .B(G110), .ZN(n1112) );
INV_X1 U1021 ( .A(n1262), .ZN(n1209) );
XNOR2_X1 U1022 ( .A(G146), .B(n1310), .ZN(n1262) );
XNOR2_X1 U1023 ( .A(n1210), .B(n1311), .ZN(n1295) );
XOR2_X1 U1024 ( .A(KEYINPUT51), .B(G125), .Z(n1311) );
NAND2_X1 U1025 ( .A1(G224), .A2(n1025), .ZN(n1210) );
XOR2_X1 U1026 ( .A(n1225), .B(KEYINPUT30), .Z(n1249) );
INV_X1 U1027 ( .A(n1039), .ZN(n1225) );
NOR2_X1 U1028 ( .A1(n1190), .A2(n1237), .ZN(n1039) );
XNOR2_X1 U1029 ( .A(n1189), .B(KEYINPUT11), .ZN(n1237) );
INV_X1 U1030 ( .A(n1242), .ZN(n1189) );
XOR2_X1 U1031 ( .A(n1312), .B(G475), .Z(n1242) );
NAND2_X1 U1032 ( .A1(KEYINPUT27), .A2(n1075), .ZN(n1312) );
NOR2_X1 U1033 ( .A1(n1134), .A2(G902), .ZN(n1075) );
XNOR2_X1 U1034 ( .A(n1313), .B(n1314), .ZN(n1134) );
XOR2_X1 U1035 ( .A(G113), .B(G104), .Z(n1314) );
XOR2_X1 U1036 ( .A(n1315), .B(n1316), .Z(n1313) );
NOR2_X1 U1037 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
XOR2_X1 U1038 ( .A(n1319), .B(KEYINPUT52), .Z(n1318) );
NAND2_X1 U1039 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NOR2_X1 U1040 ( .A1(n1320), .A2(n1321), .ZN(n1317) );
XOR2_X1 U1041 ( .A(n1322), .B(G131), .Z(n1320) );
NAND2_X1 U1042 ( .A1(KEYINPUT35), .A2(n1323), .ZN(n1322) );
XOR2_X1 U1043 ( .A(n1324), .B(n1325), .Z(n1323) );
AND2_X1 U1044 ( .A1(G214), .A2(n1263), .ZN(n1325) );
NOR2_X1 U1045 ( .A1(G953), .A2(G237), .ZN(n1263) );
NOR2_X1 U1046 ( .A1(KEYINPUT55), .A2(G143), .ZN(n1324) );
NAND2_X1 U1047 ( .A1(KEYINPUT58), .A2(n1230), .ZN(n1315) );
INV_X1 U1048 ( .A(G122), .ZN(n1230) );
NAND2_X1 U1049 ( .A1(n1326), .A2(n1327), .ZN(n1190) );
NAND2_X1 U1050 ( .A1(n1084), .A2(n1083), .ZN(n1327) );
XOR2_X1 U1051 ( .A(KEYINPUT32), .B(n1088), .Z(n1326) );
NOR2_X1 U1052 ( .A1(n1084), .A2(n1083), .ZN(n1088) );
INV_X1 U1053 ( .A(G478), .ZN(n1083) );
NOR2_X1 U1054 ( .A1(n1129), .A2(G902), .ZN(n1084) );
XOR2_X1 U1055 ( .A(n1328), .B(n1329), .Z(n1129) );
XOR2_X1 U1056 ( .A(G116), .B(n1330), .Z(n1329) );
XOR2_X1 U1057 ( .A(G134), .B(G122), .Z(n1330) );
XOR2_X1 U1058 ( .A(n1331), .B(n1310), .Z(n1328) );
XOR2_X1 U1059 ( .A(G128), .B(G143), .Z(n1310) );
XOR2_X1 U1060 ( .A(n1332), .B(G107), .Z(n1331) );
NAND3_X1 U1061 ( .A1(n1333), .A2(n1025), .A3(n1334), .ZN(n1332) );
XNOR2_X1 U1062 ( .A(G217), .B(KEYINPUT60), .ZN(n1334) );
XNOR2_X1 U1063 ( .A(n1335), .B(n1126), .ZN(n1067) );
NAND2_X1 U1064 ( .A1(G217), .A2(n1289), .ZN(n1126) );
NAND2_X1 U1065 ( .A1(G234), .A2(n1252), .ZN(n1289) );
INV_X1 U1066 ( .A(G902), .ZN(n1252) );
OR2_X1 U1067 ( .A1(n1124), .A2(G902), .ZN(n1335) );
XNOR2_X1 U1068 ( .A(n1336), .B(n1337), .ZN(n1124) );
XOR2_X1 U1069 ( .A(n1338), .B(n1339), .Z(n1337) );
XOR2_X1 U1070 ( .A(G137), .B(n1165), .Z(n1339) );
INV_X1 U1071 ( .A(G110), .ZN(n1165) );
NAND3_X1 U1072 ( .A1(n1333), .A2(n1025), .A3(G221), .ZN(n1338) );
INV_X1 U1073 ( .A(G953), .ZN(n1025) );
XOR2_X1 U1074 ( .A(G234), .B(KEYINPUT17), .Z(n1333) );
XNOR2_X1 U1075 ( .A(n1321), .B(n1340), .ZN(n1336) );
NOR2_X1 U1076 ( .A1(KEYINPUT61), .A2(n1341), .ZN(n1340) );
XOR2_X1 U1077 ( .A(G128), .B(G119), .Z(n1341) );
XNOR2_X1 U1078 ( .A(G146), .B(n1101), .ZN(n1321) );
XOR2_X1 U1079 ( .A(G125), .B(n1216), .Z(n1101) );
INV_X1 U1080 ( .A(G140), .ZN(n1216) );
endmodule


