//Key = 0011100100100101110100100010110011011101001000111111010111100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350;

XOR2_X1 U743 ( .A(n1028), .B(n1029), .Z(G9) );
NAND2_X1 U744 ( .A1(KEYINPUT63), .A2(G107), .ZN(n1029) );
NOR2_X1 U745 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U746 ( .A1(G953), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1031) );
NOR2_X1 U747 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U748 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR3_X1 U749 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NOR2_X1 U750 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U751 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U752 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U753 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U754 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U756 ( .A1(n1054), .A2(n1055), .ZN(n1046) );
NOR2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR3_X1 U758 ( .A1(n1055), .A2(n1058), .A3(n1049), .ZN(n1042) );
NOR2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR2_X1 U760 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
XOR2_X1 U761 ( .A(KEYINPUT61), .B(n1063), .Z(n1062) );
NOR4_X1 U762 ( .A1(n1064), .A2(n1045), .A3(n1049), .A4(n1055), .ZN(n1037) );
INV_X1 U763 ( .A(n1065), .ZN(n1055) );
INV_X1 U764 ( .A(n1066), .ZN(n1049) );
NOR2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1064) );
NOR2_X1 U766 ( .A1(n1039), .A2(n1069), .ZN(n1067) );
NOR3_X1 U767 ( .A1(n1032), .A2(G953), .A3(G952), .ZN(n1030) );
AND4_X1 U768 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1032) );
AND4_X1 U769 ( .A1(n1053), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1073) );
XOR2_X1 U770 ( .A(n1077), .B(KEYINPUT23), .Z(n1072) );
XOR2_X1 U771 ( .A(n1078), .B(n1079), .Z(n1071) );
XOR2_X1 U772 ( .A(n1080), .B(G469), .Z(n1070) );
XOR2_X1 U773 ( .A(n1081), .B(n1082), .Z(G72) );
NOR2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U775 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NAND3_X1 U776 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1081) );
NAND2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND3_X1 U778 ( .A1(n1092), .A2(n1093), .A3(KEYINPUT42), .ZN(n1091) );
OR3_X1 U779 ( .A1(n1094), .A2(G953), .A3(KEYINPUT35), .ZN(n1093) );
NAND2_X1 U780 ( .A1(KEYINPUT35), .A2(n1095), .ZN(n1092) );
NAND2_X1 U781 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U782 ( .A1(n1094), .A2(n1084), .ZN(n1097) );
NAND2_X1 U783 ( .A1(G900), .A2(G953), .ZN(n1096) );
NAND3_X1 U784 ( .A1(KEYINPUT42), .A2(n1098), .A3(n1099), .ZN(n1088) );
INV_X1 U785 ( .A(n1090), .ZN(n1098) );
XOR2_X1 U786 ( .A(n1100), .B(n1101), .Z(n1090) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U788 ( .A(KEYINPUT56), .B(G131), .Z(n1103) );
NOR2_X1 U789 ( .A1(n1104), .A2(KEYINPUT6), .ZN(n1102) );
NOR2_X1 U790 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U791 ( .A(n1107), .B(KEYINPUT29), .Z(n1106) );
NAND2_X1 U792 ( .A1(G137), .A2(n1108), .ZN(n1107) );
NOR2_X1 U793 ( .A1(G137), .A2(n1108), .ZN(n1105) );
XOR2_X1 U794 ( .A(n1109), .B(n1110), .Z(n1100) );
NOR2_X1 U795 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U796 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XNOR2_X1 U797 ( .A(G140), .B(KEYINPUT38), .ZN(n1114) );
NOR2_X1 U798 ( .A1(G140), .A2(n1115), .ZN(n1111) );
INV_X1 U799 ( .A(n1113), .ZN(n1115) );
XNOR2_X1 U800 ( .A(G125), .B(KEYINPUT55), .ZN(n1113) );
OR2_X1 U801 ( .A1(n1099), .A2(KEYINPUT42), .ZN(n1087) );
NOR2_X1 U802 ( .A1(G953), .A2(n1094), .ZN(n1099) );
AND2_X1 U803 ( .A1(n1116), .A2(n1117), .ZN(n1094) );
XOR2_X1 U804 ( .A(n1118), .B(n1119), .Z(G69) );
NOR2_X1 U805 ( .A1(KEYINPUT40), .A2(n1120), .ZN(n1119) );
XOR2_X1 U806 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U807 ( .A1(G953), .A2(n1123), .ZN(n1122) );
NOR2_X1 U808 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U809 ( .A(n1028), .B(KEYINPUT2), .Z(n1124) );
NOR2_X1 U810 ( .A1(n1126), .A2(n1127), .ZN(n1121) );
XOR2_X1 U811 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND2_X1 U812 ( .A1(n1130), .A2(n1131), .ZN(n1118) );
NAND2_X1 U813 ( .A1(G898), .A2(G224), .ZN(n1131) );
XOR2_X1 U814 ( .A(n1084), .B(KEYINPUT49), .Z(n1130) );
NOR2_X1 U815 ( .A1(n1132), .A2(n1133), .ZN(G66) );
XOR2_X1 U816 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U817 ( .A1(KEYINPUT0), .A2(n1136), .ZN(n1135) );
NOR2_X1 U818 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U819 ( .A(n1139), .B(KEYINPUT20), .Z(n1137) );
NOR2_X1 U820 ( .A1(n1132), .A2(n1140), .ZN(G63) );
XOR2_X1 U821 ( .A(n1141), .B(n1142), .Z(n1140) );
AND2_X1 U822 ( .A1(G478), .A2(n1143), .ZN(n1141) );
NOR2_X1 U823 ( .A1(n1132), .A2(n1144), .ZN(G60) );
XOR2_X1 U824 ( .A(n1145), .B(n1146), .Z(n1144) );
AND2_X1 U825 ( .A1(G475), .A2(n1143), .ZN(n1145) );
XOR2_X1 U826 ( .A(n1147), .B(n1148), .Z(G6) );
XOR2_X1 U827 ( .A(KEYINPUT51), .B(G104), .Z(n1148) );
NOR2_X1 U828 ( .A1(n1132), .A2(n1149), .ZN(G57) );
XOR2_X1 U829 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U830 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U831 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U832 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U833 ( .A(n1158), .B(n1159), .Z(n1156) );
NAND2_X1 U834 ( .A1(n1160), .A2(n1161), .ZN(n1154) );
NAND2_X1 U835 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XNOR2_X1 U836 ( .A(n1164), .B(KEYINPUT46), .ZN(n1150) );
NAND3_X1 U837 ( .A1(n1143), .A2(G472), .A3(KEYINPUT17), .ZN(n1164) );
NOR2_X1 U838 ( .A1(n1132), .A2(n1165), .ZN(G54) );
XOR2_X1 U839 ( .A(n1166), .B(n1167), .Z(n1165) );
AND2_X1 U840 ( .A1(G469), .A2(n1143), .ZN(n1167) );
INV_X1 U841 ( .A(n1138), .ZN(n1143) );
NOR2_X1 U842 ( .A1(n1168), .A2(n1169), .ZN(n1166) );
XOR2_X1 U843 ( .A(KEYINPUT44), .B(n1170), .Z(n1169) );
AND2_X1 U844 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U845 ( .A1(n1172), .A2(n1171), .ZN(n1168) );
NAND2_X1 U846 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
NAND2_X1 U847 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XOR2_X1 U848 ( .A(KEYINPUT16), .B(n1177), .Z(n1173) );
NOR2_X1 U849 ( .A1(n1175), .A2(n1176), .ZN(n1177) );
XOR2_X1 U850 ( .A(KEYINPUT62), .B(n1178), .Z(n1176) );
XOR2_X1 U851 ( .A(n1179), .B(n1180), .Z(n1172) );
XNOR2_X1 U852 ( .A(n1109), .B(n1158), .ZN(n1179) );
NOR2_X1 U853 ( .A1(n1132), .A2(n1181), .ZN(G51) );
XOR2_X1 U854 ( .A(n1182), .B(n1183), .Z(n1181) );
NOR2_X1 U855 ( .A1(n1184), .A2(n1138), .ZN(n1183) );
NAND2_X1 U856 ( .A1(G902), .A2(n1034), .ZN(n1138) );
NAND4_X1 U857 ( .A1(n1185), .A2(n1116), .A3(n1186), .A4(n1028), .ZN(n1034) );
NAND2_X1 U858 ( .A1(n1056), .A2(n1187), .ZN(n1028) );
XNOR2_X1 U859 ( .A(KEYINPUT3), .B(n1117), .ZN(n1186) );
AND4_X1 U860 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1116) );
NOR4_X1 U861 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
NAND2_X1 U862 ( .A1(n1196), .A2(n1197), .ZN(n1190) );
INV_X1 U863 ( .A(KEYINPUT21), .ZN(n1197) );
NAND2_X1 U864 ( .A1(n1198), .A2(n1199), .ZN(n1188) );
NAND2_X1 U865 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND3_X1 U866 ( .A1(n1057), .A2(n1202), .A3(KEYINPUT21), .ZN(n1201) );
NAND3_X1 U867 ( .A1(n1203), .A2(n1204), .A3(n1068), .ZN(n1200) );
INV_X1 U868 ( .A(n1125), .ZN(n1185) );
NAND4_X1 U869 ( .A1(n1205), .A2(n1206), .A3(n1147), .A4(n1207), .ZN(n1125) );
NOR4_X1 U870 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1207) );
INV_X1 U871 ( .A(n1212), .ZN(n1211) );
NAND2_X1 U872 ( .A1(n1057), .A2(n1187), .ZN(n1147) );
AND3_X1 U873 ( .A1(n1075), .A2(n1069), .A3(n1213), .ZN(n1187) );
NOR2_X1 U874 ( .A1(KEYINPUT41), .A2(n1214), .ZN(n1182) );
XOR2_X1 U875 ( .A(n1215), .B(n1216), .Z(n1214) );
XNOR2_X1 U876 ( .A(G125), .B(n1217), .ZN(n1216) );
NOR2_X1 U877 ( .A1(n1084), .A2(G952), .ZN(n1132) );
XOR2_X1 U878 ( .A(G146), .B(n1196), .Z(G48) );
AND3_X1 U879 ( .A1(n1057), .A2(n1218), .A3(n1198), .ZN(n1196) );
XOR2_X1 U880 ( .A(n1219), .B(n1220), .Z(G45) );
NOR2_X1 U881 ( .A1(G143), .A2(KEYINPUT11), .ZN(n1220) );
NAND4_X1 U882 ( .A1(n1221), .A2(n1198), .A3(n1203), .A4(n1204), .ZN(n1219) );
XNOR2_X1 U883 ( .A(KEYINPUT32), .B(n1068), .ZN(n1221) );
XNOR2_X1 U884 ( .A(G140), .B(n1117), .ZN(G42) );
NAND2_X1 U885 ( .A1(n1222), .A2(n1223), .ZN(n1117) );
XOR2_X1 U886 ( .A(G137), .B(n1193), .Z(G39) );
AND3_X1 U887 ( .A1(n1218), .A2(n1066), .A3(n1223), .ZN(n1193) );
XOR2_X1 U888 ( .A(G134), .B(n1192), .Z(G36) );
AND3_X1 U889 ( .A1(n1056), .A2(n1068), .A3(n1223), .ZN(n1192) );
XOR2_X1 U890 ( .A(n1224), .B(n1189), .Z(G33) );
NAND3_X1 U891 ( .A1(n1057), .A2(n1068), .A3(n1223), .ZN(n1189) );
AND3_X1 U892 ( .A1(n1074), .A2(n1225), .A3(n1051), .ZN(n1223) );
INV_X1 U893 ( .A(n1045), .ZN(n1074) );
XOR2_X1 U894 ( .A(G128), .B(n1195), .Z(G30) );
AND3_X1 U895 ( .A1(n1218), .A2(n1056), .A3(n1198), .ZN(n1195) );
AND3_X1 U896 ( .A1(n1060), .A2(n1225), .A3(n1051), .ZN(n1198) );
XOR2_X1 U897 ( .A(n1205), .B(n1226), .Z(G3) );
NAND2_X1 U898 ( .A1(KEYINPUT36), .A2(G101), .ZN(n1226) );
NAND3_X1 U899 ( .A1(n1213), .A2(n1068), .A3(n1066), .ZN(n1205) );
XOR2_X1 U900 ( .A(G125), .B(n1194), .Z(G27) );
AND4_X1 U901 ( .A1(n1222), .A2(n1065), .A3(n1060), .A4(n1225), .ZN(n1194) );
NAND2_X1 U902 ( .A1(n1036), .A2(n1227), .ZN(n1225) );
NAND4_X1 U903 ( .A1(G902), .A2(G953), .A3(n1228), .A4(n1086), .ZN(n1227) );
INV_X1 U904 ( .A(G900), .ZN(n1086) );
AND3_X1 U905 ( .A1(n1075), .A2(n1041), .A3(n1057), .ZN(n1222) );
XOR2_X1 U906 ( .A(n1229), .B(G122), .Z(G24) );
NAND2_X1 U907 ( .A1(KEYINPUT4), .A2(n1212), .ZN(n1229) );
NAND4_X1 U908 ( .A1(n1203), .A2(n1204), .A3(n1069), .A4(n1230), .ZN(n1212) );
NOR2_X1 U909 ( .A1(n1231), .A2(n1039), .ZN(n1230) );
INV_X1 U910 ( .A(n1041), .ZN(n1069) );
NAND2_X1 U911 ( .A1(n1232), .A2(n1233), .ZN(G21) );
NAND2_X1 U912 ( .A1(G119), .A2(n1206), .ZN(n1233) );
XOR2_X1 U913 ( .A(KEYINPUT37), .B(n1234), .Z(n1232) );
NOR2_X1 U914 ( .A1(G119), .A2(n1206), .ZN(n1234) );
NAND3_X1 U915 ( .A1(n1218), .A2(n1066), .A3(n1235), .ZN(n1206) );
XOR2_X1 U916 ( .A(G116), .B(n1210), .Z(G18) );
AND3_X1 U917 ( .A1(n1056), .A2(n1068), .A3(n1235), .ZN(n1210) );
NOR2_X1 U918 ( .A1(n1203), .A2(n1076), .ZN(n1056) );
XOR2_X1 U919 ( .A(G113), .B(n1209), .Z(G15) );
AND3_X1 U920 ( .A1(n1057), .A2(n1068), .A3(n1235), .ZN(n1209) );
INV_X1 U921 ( .A(n1231), .ZN(n1235) );
NAND3_X1 U922 ( .A1(n1060), .A2(n1236), .A3(n1065), .ZN(n1231) );
NOR2_X1 U923 ( .A1(n1237), .A2(n1052), .ZN(n1065) );
INV_X1 U924 ( .A(n1238), .ZN(n1052) );
NAND2_X1 U925 ( .A1(n1239), .A2(n1240), .ZN(n1068) );
OR3_X1 U926 ( .A1(n1075), .A2(n1041), .A3(KEYINPUT60), .ZN(n1240) );
NAND2_X1 U927 ( .A1(KEYINPUT60), .A2(n1218), .ZN(n1239) );
INV_X1 U928 ( .A(n1202), .ZN(n1218) );
NAND2_X1 U929 ( .A1(n1041), .A2(n1039), .ZN(n1202) );
INV_X1 U930 ( .A(n1075), .ZN(n1039) );
AND2_X1 U931 ( .A1(n1076), .A2(n1203), .ZN(n1057) );
XOR2_X1 U932 ( .A(G110), .B(n1208), .Z(G12) );
AND4_X1 U933 ( .A1(n1041), .A2(n1066), .A3(n1075), .A4(n1213), .ZN(n1208) );
AND3_X1 U934 ( .A1(n1060), .A2(n1236), .A3(n1051), .ZN(n1213) );
NOR2_X1 U935 ( .A1(n1238), .A2(n1237), .ZN(n1051) );
XNOR2_X1 U936 ( .A(n1053), .B(KEYINPUT31), .ZN(n1237) );
NAND2_X1 U937 ( .A1(G221), .A2(n1241), .ZN(n1053) );
XNOR2_X1 U938 ( .A(n1080), .B(n1242), .ZN(n1238) );
NOR2_X1 U939 ( .A1(G469), .A2(KEYINPUT14), .ZN(n1242) );
NAND2_X1 U940 ( .A1(n1243), .A2(n1244), .ZN(n1080) );
XOR2_X1 U941 ( .A(n1245), .B(n1246), .Z(n1243) );
XOR2_X1 U942 ( .A(n1247), .B(n1175), .Z(n1246) );
XOR2_X1 U943 ( .A(n1248), .B(G140), .Z(n1175) );
NAND2_X1 U944 ( .A1(KEYINPUT48), .A2(n1158), .ZN(n1247) );
XNOR2_X1 U945 ( .A(n1249), .B(n1178), .ZN(n1245) );
NOR2_X1 U946 ( .A1(n1085), .A2(G953), .ZN(n1178) );
INV_X1 U947 ( .A(G227), .ZN(n1085) );
NAND3_X1 U948 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1249) );
NAND2_X1 U949 ( .A1(KEYINPUT1), .A2(n1109), .ZN(n1252) );
OR3_X1 U950 ( .A1(n1109), .A2(KEYINPUT1), .A3(n1180), .ZN(n1251) );
NAND2_X1 U951 ( .A1(n1180), .A2(n1253), .ZN(n1250) );
NAND2_X1 U952 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
INV_X1 U953 ( .A(KEYINPUT1), .ZN(n1255) );
XOR2_X1 U954 ( .A(n1109), .B(KEYINPUT19), .Z(n1254) );
XOR2_X1 U955 ( .A(n1256), .B(n1257), .Z(n1109) );
XOR2_X1 U956 ( .A(n1258), .B(n1259), .Z(n1180) );
XOR2_X1 U957 ( .A(G101), .B(n1260), .Z(n1258) );
NAND2_X1 U958 ( .A1(n1036), .A2(n1261), .ZN(n1236) );
NAND3_X1 U959 ( .A1(n1126), .A2(n1228), .A3(G902), .ZN(n1261) );
NOR2_X1 U960 ( .A1(n1084), .A2(G898), .ZN(n1126) );
NAND3_X1 U961 ( .A1(n1228), .A2(n1084), .A3(G952), .ZN(n1036) );
NAND2_X1 U962 ( .A1(G237), .A2(n1262), .ZN(n1228) );
NAND2_X1 U963 ( .A1(n1263), .A2(n1264), .ZN(n1060) );
OR2_X1 U964 ( .A1(n1045), .A2(KEYINPUT53), .ZN(n1264) );
NAND2_X1 U965 ( .A1(n1265), .A2(n1061), .ZN(n1045) );
NAND3_X1 U966 ( .A1(n1063), .A2(n1061), .A3(KEYINPUT53), .ZN(n1263) );
NAND2_X1 U967 ( .A1(G214), .A2(n1266), .ZN(n1061) );
INV_X1 U968 ( .A(n1265), .ZN(n1063) );
XNOR2_X1 U969 ( .A(n1267), .B(n1184), .ZN(n1265) );
NAND2_X1 U970 ( .A1(G210), .A2(n1266), .ZN(n1184) );
NAND2_X1 U971 ( .A1(n1268), .A2(n1244), .ZN(n1266) );
NAND2_X1 U972 ( .A1(n1269), .A2(n1244), .ZN(n1267) );
XOR2_X1 U973 ( .A(n1217), .B(n1270), .Z(n1269) );
XNOR2_X1 U974 ( .A(n1271), .B(n1272), .ZN(n1270) );
NOR2_X1 U975 ( .A1(G125), .A2(KEYINPUT45), .ZN(n1272) );
NAND2_X1 U976 ( .A1(KEYINPUT7), .A2(n1215), .ZN(n1271) );
XOR2_X1 U977 ( .A(n1273), .B(n1274), .Z(n1215) );
INV_X1 U978 ( .A(n1128), .ZN(n1274) );
XOR2_X1 U979 ( .A(n1275), .B(n1276), .Z(n1128) );
XOR2_X1 U980 ( .A(G122), .B(G110), .Z(n1276) );
NAND2_X1 U981 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
NAND2_X1 U982 ( .A1(G113), .A2(n1279), .ZN(n1278) );
XOR2_X1 U983 ( .A(KEYINPUT10), .B(n1280), .Z(n1277) );
NOR2_X1 U984 ( .A1(G113), .A2(n1279), .ZN(n1280) );
NAND2_X1 U985 ( .A1(n1281), .A2(n1282), .ZN(n1279) );
NAND2_X1 U986 ( .A1(G119), .A2(n1283), .ZN(n1282) );
XOR2_X1 U987 ( .A(n1284), .B(KEYINPUT5), .Z(n1281) );
OR2_X1 U988 ( .A1(n1283), .A2(G119), .ZN(n1284) );
XOR2_X1 U989 ( .A(G116), .B(KEYINPUT33), .Z(n1283) );
NAND2_X1 U990 ( .A1(KEYINPUT13), .A2(n1129), .ZN(n1273) );
XOR2_X1 U991 ( .A(n1285), .B(n1259), .Z(n1129) );
XOR2_X1 U992 ( .A(G104), .B(KEYINPUT12), .Z(n1259) );
XNOR2_X1 U993 ( .A(n1286), .B(n1287), .ZN(n1285) );
NAND2_X1 U994 ( .A1(KEYINPUT57), .A2(G101), .ZN(n1287) );
NAND2_X1 U995 ( .A1(KEYINPUT47), .A2(G107), .ZN(n1286) );
XOR2_X1 U996 ( .A(n1157), .B(n1288), .Z(n1217) );
AND2_X1 U997 ( .A1(n1084), .A2(G224), .ZN(n1288) );
XOR2_X1 U998 ( .A(n1289), .B(G472), .Z(n1075) );
NAND2_X1 U999 ( .A1(n1290), .A2(n1244), .ZN(n1289) );
XOR2_X1 U1000 ( .A(n1291), .B(n1152), .Z(n1290) );
XNOR2_X1 U1001 ( .A(G101), .B(n1292), .ZN(n1152) );
AND3_X1 U1002 ( .A1(G210), .A2(n1084), .A3(n1268), .ZN(n1292) );
INV_X1 U1003 ( .A(G237), .ZN(n1268) );
NAND2_X1 U1004 ( .A1(n1293), .A2(n1294), .ZN(n1291) );
NAND3_X1 U1005 ( .A1(n1295), .A2(n1296), .A3(n1160), .ZN(n1294) );
NAND3_X1 U1006 ( .A1(n1297), .A2(n1298), .A3(n1162), .ZN(n1295) );
OR2_X1 U1007 ( .A1(n1163), .A2(n1299), .ZN(n1298) );
NAND2_X1 U1008 ( .A1(n1159), .A2(n1299), .ZN(n1297) );
NAND4_X1 U1009 ( .A1(n1300), .A2(n1163), .A3(n1301), .A4(n1302), .ZN(n1293) );
NAND2_X1 U1010 ( .A1(n1303), .A2(n1299), .ZN(n1302) );
INV_X1 U1011 ( .A(n1159), .ZN(n1303) );
OR2_X1 U1012 ( .A1(n1162), .A2(n1299), .ZN(n1301) );
INV_X1 U1013 ( .A(KEYINPUT26), .ZN(n1299) );
NAND2_X1 U1014 ( .A1(n1159), .A2(n1158), .ZN(n1162) );
OR2_X1 U1015 ( .A1(n1159), .A2(n1158), .ZN(n1163) );
XOR2_X1 U1016 ( .A(n1304), .B(n1108), .Z(n1158) );
XOR2_X1 U1017 ( .A(G134), .B(KEYINPUT28), .Z(n1108) );
XOR2_X1 U1018 ( .A(n1224), .B(G137), .Z(n1304) );
INV_X1 U1019 ( .A(G131), .ZN(n1224) );
XOR2_X1 U1020 ( .A(n1305), .B(n1306), .Z(n1159) );
XOR2_X1 U1021 ( .A(KEYINPUT9), .B(G119), .Z(n1306) );
XNOR2_X1 U1022 ( .A(G113), .B(G116), .ZN(n1305) );
NAND2_X1 U1023 ( .A1(n1160), .A2(n1296), .ZN(n1300) );
INV_X1 U1024 ( .A(KEYINPUT27), .ZN(n1296) );
INV_X1 U1025 ( .A(n1157), .ZN(n1160) );
NAND2_X1 U1026 ( .A1(n1307), .A2(n1308), .ZN(n1157) );
NAND2_X1 U1027 ( .A1(n1256), .A2(G146), .ZN(n1308) );
NAND2_X1 U1028 ( .A1(n1309), .A2(n1257), .ZN(n1307) );
XNOR2_X1 U1029 ( .A(n1256), .B(KEYINPUT59), .ZN(n1309) );
XNOR2_X1 U1030 ( .A(n1310), .B(n1311), .ZN(n1256) );
XOR2_X1 U1031 ( .A(KEYINPUT8), .B(G143), .Z(n1311) );
INV_X1 U1032 ( .A(G128), .ZN(n1310) );
NOR2_X1 U1033 ( .A1(n1204), .A2(n1203), .ZN(n1066) );
XNOR2_X1 U1034 ( .A(n1077), .B(KEYINPUT43), .ZN(n1203) );
XOR2_X1 U1035 ( .A(n1312), .B(G475), .Z(n1077) );
OR2_X1 U1036 ( .A1(n1146), .A2(G902), .ZN(n1312) );
XNOR2_X1 U1037 ( .A(n1313), .B(n1314), .ZN(n1146) );
XOR2_X1 U1038 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1039 ( .A(G104), .B(n1317), .ZN(n1316) );
NOR4_X1 U1040 ( .A1(KEYINPUT24), .A2(G953), .A3(G237), .A4(n1318), .ZN(n1317) );
INV_X1 U1041 ( .A(G214), .ZN(n1318) );
NAND2_X1 U1042 ( .A1(n1319), .A2(KEYINPUT58), .ZN(n1315) );
XOR2_X1 U1043 ( .A(n1257), .B(n1320), .Z(n1319) );
NOR2_X1 U1044 ( .A1(KEYINPUT54), .A2(n1321), .ZN(n1320) );
INV_X1 U1045 ( .A(n1322), .ZN(n1321) );
XOR2_X1 U1046 ( .A(n1323), .B(n1324), .Z(n1313) );
XOR2_X1 U1047 ( .A(G143), .B(G131), .Z(n1324) );
XNOR2_X1 U1048 ( .A(G113), .B(G122), .ZN(n1323) );
INV_X1 U1049 ( .A(n1076), .ZN(n1204) );
XOR2_X1 U1050 ( .A(n1325), .B(G478), .Z(n1076) );
OR2_X1 U1051 ( .A1(n1142), .A2(G902), .ZN(n1325) );
XNOR2_X1 U1052 ( .A(n1326), .B(n1327), .ZN(n1142) );
XNOR2_X1 U1053 ( .A(n1328), .B(n1329), .ZN(n1327) );
NOR2_X1 U1054 ( .A1(G116), .A2(KEYINPUT30), .ZN(n1329) );
NAND2_X1 U1055 ( .A1(KEYINPUT22), .A2(n1330), .ZN(n1328) );
XOR2_X1 U1056 ( .A(n1331), .B(n1332), .Z(n1330) );
XOR2_X1 U1057 ( .A(G143), .B(G128), .Z(n1332) );
NOR2_X1 U1058 ( .A1(G134), .A2(KEYINPUT25), .ZN(n1331) );
XOR2_X1 U1059 ( .A(n1333), .B(n1334), .Z(n1326) );
XOR2_X1 U1060 ( .A(G122), .B(n1335), .Z(n1334) );
AND3_X1 U1061 ( .A1(G234), .A2(n1084), .A3(G217), .ZN(n1335) );
NAND2_X1 U1062 ( .A1(KEYINPUT50), .A2(n1260), .ZN(n1333) );
INV_X1 U1063 ( .A(G107), .ZN(n1260) );
XOR2_X1 U1064 ( .A(n1078), .B(n1336), .Z(n1041) );
NOR2_X1 U1065 ( .A1(n1079), .A2(KEYINPUT52), .ZN(n1336) );
INV_X1 U1066 ( .A(n1139), .ZN(n1079) );
NAND2_X1 U1067 ( .A1(G217), .A2(n1241), .ZN(n1139) );
NAND2_X1 U1068 ( .A1(n1262), .A2(n1244), .ZN(n1241) );
XNOR2_X1 U1069 ( .A(G234), .B(KEYINPUT15), .ZN(n1262) );
NAND2_X1 U1070 ( .A1(n1134), .A2(n1244), .ZN(n1078) );
INV_X1 U1071 ( .A(G902), .ZN(n1244) );
XOR2_X1 U1072 ( .A(n1337), .B(n1338), .Z(n1134) );
XNOR2_X1 U1073 ( .A(G137), .B(n1339), .ZN(n1338) );
NAND2_X1 U1074 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
OR2_X1 U1075 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
XOR2_X1 U1076 ( .A(n1344), .B(KEYINPUT18), .Z(n1340) );
NAND2_X1 U1077 ( .A1(n1343), .A2(n1342), .ZN(n1344) );
NAND3_X1 U1078 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1342) );
OR2_X1 U1079 ( .A1(n1322), .A2(KEYINPUT39), .ZN(n1347) );
NAND3_X1 U1080 ( .A1(KEYINPUT39), .A2(n1322), .A3(G146), .ZN(n1346) );
NAND2_X1 U1081 ( .A1(n1348), .A2(n1257), .ZN(n1345) );
INV_X1 U1082 ( .A(G146), .ZN(n1257) );
NAND2_X1 U1083 ( .A1(KEYINPUT39), .A2(n1349), .ZN(n1348) );
XOR2_X1 U1084 ( .A(KEYINPUT34), .B(n1322), .Z(n1349) );
XOR2_X1 U1085 ( .A(G125), .B(G140), .Z(n1322) );
XNOR2_X1 U1086 ( .A(n1248), .B(n1350), .ZN(n1343) );
XOR2_X1 U1087 ( .A(G128), .B(G119), .Z(n1350) );
INV_X1 U1088 ( .A(G110), .ZN(n1248) );
NAND3_X1 U1089 ( .A1(G234), .A2(n1084), .A3(G221), .ZN(n1337) );
INV_X1 U1090 ( .A(G953), .ZN(n1084) );
endmodule


