//Key = 0100100011111000100110000001000000110011001000101011001011010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407;

XOR2_X1 U779 ( .A(G107), .B(n1074), .Z(G9) );
NOR2_X1 U780 ( .A1(n1075), .A2(n1076), .ZN(G75) );
NOR4_X1 U781 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1076) );
XOR2_X1 U782 ( .A(n1081), .B(KEYINPUT59), .Z(n1079) );
NAND4_X1 U783 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1081) );
AND2_X1 U784 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND4_X1 U785 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1077) );
NAND4_X1 U786 ( .A1(n1087), .A2(n1092), .A3(n1083), .A4(n1093), .ZN(n1089) );
NAND3_X1 U787 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
NAND2_X1 U788 ( .A1(n1082), .A2(n1097), .ZN(n1096) );
NAND3_X1 U789 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1095) );
XOR2_X1 U790 ( .A(KEYINPUT0), .B(n1082), .Z(n1099) );
NAND2_X1 U791 ( .A1(n1086), .A2(n1101), .ZN(n1094) );
NAND2_X1 U792 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND2_X1 U793 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U794 ( .A1(n1086), .A2(n1106), .ZN(n1088) );
NAND2_X1 U795 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND3_X1 U796 ( .A1(n1082), .A2(n1109), .A3(n1087), .ZN(n1108) );
NAND2_X1 U797 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U798 ( .A1(n1112), .A2(n1083), .ZN(n1111) );
NAND2_X1 U799 ( .A1(n1113), .A2(n1092), .ZN(n1110) );
XOR2_X1 U800 ( .A(n1114), .B(KEYINPUT24), .Z(n1107) );
NAND4_X1 U801 ( .A1(n1087), .A2(n1082), .A3(n1115), .A4(n1092), .ZN(n1114) );
INV_X1 U802 ( .A(n1116), .ZN(n1087) );
NOR3_X1 U803 ( .A1(n1117), .A2(G953), .A3(G952), .ZN(n1075) );
INV_X1 U804 ( .A(n1090), .ZN(n1117) );
NAND4_X1 U805 ( .A1(n1083), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1090) );
NOR4_X1 U806 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1120) );
XNOR2_X1 U807 ( .A(G469), .B(n1125), .ZN(n1124) );
XNOR2_X1 U808 ( .A(G475), .B(n1126), .ZN(n1123) );
NOR2_X1 U809 ( .A1(n1127), .A2(n1128), .ZN(n1122) );
NOR2_X1 U810 ( .A1(G478), .A2(n1129), .ZN(n1121) );
NOR2_X1 U811 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
AND2_X1 U812 ( .A1(n1127), .A2(KEYINPUT50), .ZN(n1131) );
OR2_X1 U813 ( .A1(n1132), .A2(KEYINPUT40), .ZN(n1127) );
NOR2_X1 U814 ( .A1(KEYINPUT50), .A2(n1132), .ZN(n1130) );
NOR2_X1 U815 ( .A1(n1104), .A2(n1100), .ZN(n1119) );
XNOR2_X1 U816 ( .A(KEYINPUT63), .B(n1098), .ZN(n1118) );
NAND2_X1 U817 ( .A1(n1133), .A2(n1134), .ZN(G72) );
NAND2_X1 U818 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U819 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
NAND2_X1 U820 ( .A1(n1139), .A2(n1138), .ZN(n1133) );
NAND2_X1 U821 ( .A1(G953), .A2(n1140), .ZN(n1138) );
INV_X1 U822 ( .A(G227), .ZN(n1140) );
INV_X1 U823 ( .A(n1136), .ZN(n1139) );
NAND2_X1 U824 ( .A1(KEYINPUT46), .A2(n1141), .ZN(n1136) );
XOR2_X1 U825 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND2_X1 U826 ( .A1(n1091), .A2(n1080), .ZN(n1143) );
NAND2_X1 U827 ( .A1(n1144), .A2(n1137), .ZN(n1142) );
INV_X1 U828 ( .A(n1145), .ZN(n1137) );
XOR2_X1 U829 ( .A(n1146), .B(n1147), .Z(n1144) );
XOR2_X1 U830 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U831 ( .A(KEYINPUT6), .B(KEYINPUT11), .Z(n1149) );
NOR2_X1 U832 ( .A1(KEYINPUT15), .A2(n1150), .ZN(n1148) );
XOR2_X1 U833 ( .A(n1151), .B(n1152), .Z(n1146) );
XNOR2_X1 U834 ( .A(n1153), .B(n1154), .ZN(n1151) );
XOR2_X1 U835 ( .A(n1155), .B(n1156), .Z(G69) );
XOR2_X1 U836 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U837 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U838 ( .A(KEYINPUT28), .B(n1091), .ZN(n1160) );
INV_X1 U839 ( .A(n1078), .ZN(n1159) );
NAND3_X1 U840 ( .A1(G953), .A2(n1161), .A3(KEYINPUT19), .ZN(n1157) );
NAND2_X1 U841 ( .A1(G898), .A2(G224), .ZN(n1161) );
OR2_X1 U842 ( .A1(n1162), .A2(n1163), .ZN(n1155) );
NOR2_X1 U843 ( .A1(n1164), .A2(n1165), .ZN(G66) );
XOR2_X1 U844 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U845 ( .A1(n1168), .A2(n1169), .ZN(n1166) );
NOR2_X1 U846 ( .A1(n1164), .A2(n1170), .ZN(G63) );
NOR3_X1 U847 ( .A1(n1132), .A2(n1171), .A3(n1172), .ZN(n1170) );
NOR3_X1 U848 ( .A1(n1173), .A2(n1174), .A3(n1169), .ZN(n1172) );
NOR2_X1 U849 ( .A1(n1175), .A2(n1176), .ZN(n1171) );
NOR2_X1 U850 ( .A1(n1177), .A2(n1174), .ZN(n1176) );
XNOR2_X1 U851 ( .A(n1128), .B(KEYINPUT48), .ZN(n1174) );
NOR2_X1 U852 ( .A1(n1080), .A2(n1078), .ZN(n1177) );
NOR2_X1 U853 ( .A1(n1164), .A2(n1178), .ZN(G60) );
XOR2_X1 U854 ( .A(n1179), .B(n1180), .Z(n1178) );
NAND2_X1 U855 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
XNOR2_X1 U856 ( .A(KEYINPUT60), .B(n1183), .ZN(n1182) );
XOR2_X1 U857 ( .A(G104), .B(n1184), .Z(G6) );
NOR2_X1 U858 ( .A1(KEYINPUT47), .A2(n1185), .ZN(n1184) );
NOR2_X1 U859 ( .A1(n1164), .A2(n1186), .ZN(G57) );
XOR2_X1 U860 ( .A(n1187), .B(n1188), .Z(n1186) );
XNOR2_X1 U861 ( .A(n1189), .B(n1190), .ZN(n1188) );
XOR2_X1 U862 ( .A(n1191), .B(n1192), .Z(n1187) );
XOR2_X1 U863 ( .A(KEYINPUT54), .B(n1193), .Z(n1192) );
NOR2_X1 U864 ( .A1(KEYINPUT29), .A2(n1194), .ZN(n1193) );
AND2_X1 U865 ( .A1(G472), .A2(n1181), .ZN(n1191) );
NOR2_X1 U866 ( .A1(n1164), .A2(n1195), .ZN(G54) );
XOR2_X1 U867 ( .A(n1196), .B(n1197), .Z(n1195) );
NOR2_X1 U868 ( .A1(n1198), .A2(n1169), .ZN(n1197) );
NAND2_X1 U869 ( .A1(KEYINPUT1), .A2(n1199), .ZN(n1196) );
XNOR2_X1 U870 ( .A(n1200), .B(n1201), .ZN(n1199) );
NAND2_X1 U871 ( .A1(n1202), .A2(n1203), .ZN(n1200) );
OR2_X1 U872 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
XOR2_X1 U873 ( .A(n1206), .B(KEYINPUT3), .Z(n1202) );
NAND2_X1 U874 ( .A1(n1207), .A2(n1205), .ZN(n1206) );
NAND3_X1 U875 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1205) );
OR2_X1 U876 ( .A1(n1211), .A2(KEYINPUT56), .ZN(n1210) );
NAND3_X1 U877 ( .A1(KEYINPUT56), .A2(n1211), .A3(G110), .ZN(n1209) );
NAND2_X1 U878 ( .A1(n1212), .A2(n1213), .ZN(n1208) );
NAND2_X1 U879 ( .A1(KEYINPUT56), .A2(n1214), .ZN(n1212) );
XNOR2_X1 U880 ( .A(KEYINPUT39), .B(n1211), .ZN(n1214) );
XOR2_X1 U881 ( .A(n1204), .B(KEYINPUT36), .Z(n1207) );
NOR2_X1 U882 ( .A1(n1164), .A2(n1215), .ZN(G51) );
NOR2_X1 U883 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
XOR2_X1 U884 ( .A(KEYINPUT45), .B(n1218), .Z(n1217) );
NOR2_X1 U885 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
XOR2_X1 U886 ( .A(n1221), .B(n1222), .Z(n1219) );
XOR2_X1 U887 ( .A(KEYINPUT9), .B(KEYINPUT25), .Z(n1222) );
NOR2_X1 U888 ( .A1(n1223), .A2(n1221), .ZN(n1216) );
XOR2_X1 U889 ( .A(n1224), .B(n1225), .Z(n1221) );
XNOR2_X1 U890 ( .A(n1162), .B(n1194), .ZN(n1225) );
XNOR2_X1 U891 ( .A(n1226), .B(n1227), .ZN(n1224) );
INV_X1 U892 ( .A(n1220), .ZN(n1223) );
NAND2_X1 U893 ( .A1(n1181), .A2(n1228), .ZN(n1220) );
INV_X1 U894 ( .A(n1169), .ZN(n1181) );
NAND2_X1 U895 ( .A1(G902), .A2(n1229), .ZN(n1169) );
OR2_X1 U896 ( .A1(n1078), .A2(n1080), .ZN(n1229) );
NAND4_X1 U897 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1080) );
AND4_X1 U898 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1233) );
OR2_X1 U899 ( .A1(n1238), .A2(KEYINPUT22), .ZN(n1232) );
NAND4_X1 U900 ( .A1(n1239), .A2(n1240), .A3(n1097), .A4(n1241), .ZN(n1231) );
NOR2_X1 U901 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND2_X1 U902 ( .A1(n1244), .A2(n1245), .ZN(n1240) );
NAND3_X1 U903 ( .A1(n1112), .A2(n1102), .A3(KEYINPUT22), .ZN(n1245) );
NAND2_X1 U904 ( .A1(n1246), .A2(n1247), .ZN(n1239) );
NAND2_X1 U905 ( .A1(n1084), .A2(n1082), .ZN(n1247) );
NAND2_X1 U906 ( .A1(n1248), .A2(n1249), .ZN(n1230) );
NAND2_X1 U907 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NAND3_X1 U908 ( .A1(n1112), .A2(n1252), .A3(n1113), .ZN(n1251) );
XOR2_X1 U909 ( .A(KEYINPUT52), .B(n1086), .Z(n1252) );
NAND3_X1 U910 ( .A1(n1253), .A2(n1092), .A3(n1086), .ZN(n1250) );
NAND4_X1 U911 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1078) );
NOR4_X1 U912 ( .A1(n1258), .A2(n1259), .A3(n1074), .A4(n1260), .ZN(n1257) );
AND3_X1 U913 ( .A1(n1083), .A2(n1261), .A3(n1112), .ZN(n1074) );
AND2_X1 U914 ( .A1(n1262), .A2(n1185), .ZN(n1256) );
NAND3_X1 U915 ( .A1(n1083), .A2(n1261), .A3(n1084), .ZN(n1185) );
NOR2_X1 U916 ( .A1(n1091), .A2(G952), .ZN(n1164) );
XNOR2_X1 U917 ( .A(G146), .B(n1236), .ZN(G48) );
NAND3_X1 U918 ( .A1(n1253), .A2(n1097), .A3(n1263), .ZN(n1236) );
XNOR2_X1 U919 ( .A(G143), .B(n1237), .ZN(G45) );
NAND3_X1 U920 ( .A1(n1248), .A2(n1113), .A3(n1264), .ZN(n1237) );
AND3_X1 U921 ( .A1(n1097), .A2(n1265), .A3(n1266), .ZN(n1264) );
XNOR2_X1 U922 ( .A(G140), .B(n1235), .ZN(G42) );
NAND3_X1 U923 ( .A1(n1263), .A2(n1115), .A3(n1086), .ZN(n1235) );
XOR2_X1 U924 ( .A(n1267), .B(n1268), .Z(G39) );
NAND2_X1 U925 ( .A1(KEYINPUT12), .A2(G137), .ZN(n1268) );
NAND4_X1 U926 ( .A1(n1269), .A2(n1270), .A3(n1092), .A4(n1271), .ZN(n1267) );
AND2_X1 U927 ( .A1(n1253), .A2(n1086), .ZN(n1271) );
XNOR2_X1 U928 ( .A(KEYINPUT43), .B(n1102), .ZN(n1269) );
XNOR2_X1 U929 ( .A(G134), .B(n1272), .ZN(G36) );
NAND4_X1 U930 ( .A1(n1273), .A2(n1274), .A3(n1086), .A4(n1275), .ZN(n1272) );
AND2_X1 U931 ( .A1(n1112), .A2(n1113), .ZN(n1275) );
OR2_X1 U932 ( .A1(n1248), .A2(KEYINPUT33), .ZN(n1274) );
NAND2_X1 U933 ( .A1(KEYINPUT33), .A2(n1276), .ZN(n1273) );
NAND2_X1 U934 ( .A1(n1242), .A2(n1277), .ZN(n1276) );
XNOR2_X1 U935 ( .A(G131), .B(n1234), .ZN(G33) );
NAND3_X1 U936 ( .A1(n1263), .A2(n1113), .A3(n1086), .ZN(n1234) );
NOR2_X1 U937 ( .A1(n1278), .A2(n1100), .ZN(n1086) );
AND2_X1 U938 ( .A1(n1248), .A2(n1084), .ZN(n1263) );
XNOR2_X1 U939 ( .A(G128), .B(n1238), .ZN(G30) );
NAND4_X1 U940 ( .A1(n1248), .A2(n1253), .A3(n1112), .A4(n1097), .ZN(n1238) );
NOR2_X1 U941 ( .A1(n1102), .A2(n1242), .ZN(n1248) );
INV_X1 U942 ( .A(n1270), .ZN(n1242) );
INV_X1 U943 ( .A(n1277), .ZN(n1102) );
XNOR2_X1 U944 ( .A(n1279), .B(n1280), .ZN(G3) );
NOR2_X1 U945 ( .A1(KEYINPUT53), .A2(n1262), .ZN(n1280) );
NAND3_X1 U946 ( .A1(n1092), .A2(n1261), .A3(n1113), .ZN(n1262) );
NAND2_X1 U947 ( .A1(n1281), .A2(n1282), .ZN(G27) );
NAND2_X1 U948 ( .A1(n1283), .A2(n1226), .ZN(n1282) );
NAND2_X1 U949 ( .A1(G125), .A2(n1284), .ZN(n1281) );
NAND2_X1 U950 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
OR2_X1 U951 ( .A1(n1287), .A2(KEYINPUT20), .ZN(n1286) );
NAND2_X1 U952 ( .A1(KEYINPUT20), .A2(n1288), .ZN(n1285) );
INV_X1 U953 ( .A(n1283), .ZN(n1288) );
NOR2_X1 U954 ( .A1(KEYINPUT58), .A2(n1287), .ZN(n1283) );
NAND4_X1 U955 ( .A1(n1289), .A2(n1270), .A3(n1115), .A4(n1290), .ZN(n1287) );
AND2_X1 U956 ( .A1(n1082), .A2(n1084), .ZN(n1290) );
NAND2_X1 U957 ( .A1(n1116), .A2(n1291), .ZN(n1270) );
NAND3_X1 U958 ( .A1(G902), .A2(n1292), .A3(n1145), .ZN(n1291) );
NOR2_X1 U959 ( .A1(G900), .A2(n1091), .ZN(n1145) );
XOR2_X1 U960 ( .A(KEYINPUT31), .B(n1097), .Z(n1289) );
XNOR2_X1 U961 ( .A(G122), .B(n1254), .ZN(G24) );
NAND4_X1 U962 ( .A1(n1293), .A2(n1083), .A3(n1266), .A4(n1265), .ZN(n1254) );
NOR2_X1 U963 ( .A1(n1294), .A2(n1244), .ZN(n1083) );
XNOR2_X1 U964 ( .A(G119), .B(n1255), .ZN(G21) );
NAND3_X1 U965 ( .A1(n1293), .A2(n1092), .A3(n1253), .ZN(n1255) );
NOR2_X1 U966 ( .A1(n1246), .A2(n1243), .ZN(n1253) );
XOR2_X1 U967 ( .A(G116), .B(n1260), .Z(G18) );
AND3_X1 U968 ( .A1(n1293), .A2(n1112), .A3(n1113), .ZN(n1260) );
AND2_X1 U969 ( .A1(n1295), .A2(n1265), .ZN(n1112) );
NAND2_X1 U970 ( .A1(n1296), .A2(n1297), .ZN(G15) );
NAND2_X1 U971 ( .A1(n1259), .A2(n1298), .ZN(n1297) );
XOR2_X1 U972 ( .A(KEYINPUT42), .B(n1299), .Z(n1296) );
NOR2_X1 U973 ( .A1(n1259), .A2(n1298), .ZN(n1299) );
AND3_X1 U974 ( .A1(n1084), .A2(n1293), .A3(n1113), .ZN(n1259) );
NOR2_X1 U975 ( .A1(n1294), .A2(n1246), .ZN(n1113) );
INV_X1 U976 ( .A(n1244), .ZN(n1246) );
AND2_X1 U977 ( .A1(n1082), .A2(n1300), .ZN(n1293) );
AND2_X1 U978 ( .A1(n1105), .A2(n1301), .ZN(n1082) );
NOR2_X1 U979 ( .A1(n1265), .A2(n1295), .ZN(n1084) );
INV_X1 U980 ( .A(n1266), .ZN(n1295) );
XOR2_X1 U981 ( .A(n1258), .B(n1302), .Z(G12) );
NOR2_X1 U982 ( .A1(KEYINPUT21), .A2(n1213), .ZN(n1302) );
AND3_X1 U983 ( .A1(n1092), .A2(n1261), .A3(n1115), .ZN(n1258) );
NOR2_X1 U984 ( .A1(n1244), .A2(n1243), .ZN(n1115) );
INV_X1 U985 ( .A(n1294), .ZN(n1243) );
XOR2_X1 U986 ( .A(n1303), .B(n1168), .Z(n1294) );
NAND2_X1 U987 ( .A1(G217), .A2(n1304), .ZN(n1168) );
OR2_X1 U988 ( .A1(n1167), .A2(G902), .ZN(n1303) );
XNOR2_X1 U989 ( .A(n1305), .B(n1306), .ZN(n1167) );
XNOR2_X1 U990 ( .A(n1307), .B(n1152), .ZN(n1306) );
XOR2_X1 U991 ( .A(n1308), .B(n1309), .Z(n1305) );
NOR2_X1 U992 ( .A1(G110), .A2(KEYINPUT44), .ZN(n1309) );
XOR2_X1 U993 ( .A(n1310), .B(G119), .Z(n1308) );
NAND2_X1 U994 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NAND4_X1 U995 ( .A1(G221), .A2(G137), .A3(G234), .A4(n1091), .ZN(n1312) );
XOR2_X1 U996 ( .A(n1313), .B(KEYINPUT32), .Z(n1311) );
NAND2_X1 U997 ( .A1(n1150), .A2(n1314), .ZN(n1313) );
NAND3_X1 U998 ( .A1(G234), .A2(n1091), .A3(G221), .ZN(n1314) );
XNOR2_X1 U999 ( .A(n1315), .B(G472), .ZN(n1244) );
NAND2_X1 U1000 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XOR2_X1 U1001 ( .A(n1318), .B(n1319), .Z(n1316) );
XNOR2_X1 U1002 ( .A(n1190), .B(n1320), .ZN(n1319) );
INV_X1 U1003 ( .A(n1189), .ZN(n1320) );
XOR2_X1 U1004 ( .A(n1321), .B(n1279), .Z(n1189) );
INV_X1 U1005 ( .A(G101), .ZN(n1279) );
NAND2_X1 U1006 ( .A1(G210), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1007 ( .A(n1323), .B(n1324), .Z(n1190) );
XNOR2_X1 U1008 ( .A(n1325), .B(G113), .ZN(n1323) );
XNOR2_X1 U1009 ( .A(n1326), .B(KEYINPUT23), .ZN(n1318) );
AND2_X1 U1010 ( .A1(n1300), .A2(n1277), .ZN(n1261) );
NOR2_X1 U1011 ( .A1(n1105), .A2(n1104), .ZN(n1277) );
INV_X1 U1012 ( .A(n1301), .ZN(n1104) );
NAND2_X1 U1013 ( .A1(G221), .A2(n1304), .ZN(n1301) );
NAND2_X1 U1014 ( .A1(n1327), .A2(G234), .ZN(n1304) );
XOR2_X1 U1015 ( .A(n1328), .B(n1329), .Z(n1105) );
XNOR2_X1 U1016 ( .A(KEYINPUT27), .B(n1125), .ZN(n1329) );
NAND2_X1 U1017 ( .A1(n1330), .A2(n1317), .ZN(n1125) );
XOR2_X1 U1018 ( .A(n1331), .B(n1332), .Z(n1330) );
XNOR2_X1 U1019 ( .A(n1211), .B(n1333), .ZN(n1332) );
NOR2_X1 U1020 ( .A1(KEYINPUT41), .A2(n1334), .ZN(n1333) );
XNOR2_X1 U1021 ( .A(KEYINPUT30), .B(n1213), .ZN(n1334) );
INV_X1 U1022 ( .A(G110), .ZN(n1213) );
INV_X1 U1023 ( .A(G140), .ZN(n1211) );
XNOR2_X1 U1024 ( .A(n1335), .B(n1336), .ZN(n1331) );
INV_X1 U1025 ( .A(n1201), .ZN(n1336) );
XNOR2_X1 U1026 ( .A(n1337), .B(n1325), .ZN(n1201) );
XNOR2_X1 U1027 ( .A(n1150), .B(n1153), .ZN(n1325) );
XNOR2_X1 U1028 ( .A(G131), .B(n1338), .ZN(n1153) );
INV_X1 U1029 ( .A(G137), .ZN(n1150) );
XOR2_X1 U1030 ( .A(n1339), .B(n1154), .Z(n1337) );
XNOR2_X1 U1031 ( .A(n1307), .B(n1340), .ZN(n1154) );
NOR2_X1 U1032 ( .A1(G143), .A2(KEYINPUT7), .ZN(n1340) );
NAND2_X1 U1033 ( .A1(KEYINPUT57), .A2(n1204), .ZN(n1335) );
NAND2_X1 U1034 ( .A1(G227), .A2(n1091), .ZN(n1204) );
NAND2_X1 U1035 ( .A1(KEYINPUT34), .A2(n1198), .ZN(n1328) );
INV_X1 U1036 ( .A(G469), .ZN(n1198) );
AND2_X1 U1037 ( .A1(n1097), .A2(n1341), .ZN(n1300) );
NAND2_X1 U1038 ( .A1(n1116), .A2(n1342), .ZN(n1341) );
NAND3_X1 U1039 ( .A1(G902), .A2(n1292), .A3(n1163), .ZN(n1342) );
NOR2_X1 U1040 ( .A1(n1091), .A2(G898), .ZN(n1163) );
NAND3_X1 U1041 ( .A1(n1292), .A2(n1091), .A3(G952), .ZN(n1116) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1292) );
NOR2_X1 U1043 ( .A1(n1098), .A2(n1100), .ZN(n1097) );
AND2_X1 U1044 ( .A1(G214), .A2(n1343), .ZN(n1100) );
INV_X1 U1045 ( .A(n1278), .ZN(n1098) );
XNOR2_X1 U1046 ( .A(n1344), .B(n1228), .ZN(n1278) );
AND2_X1 U1047 ( .A1(G210), .A2(n1343), .ZN(n1228) );
NAND2_X1 U1048 ( .A1(n1345), .A2(n1327), .ZN(n1343) );
XNOR2_X1 U1049 ( .A(G902), .B(KEYINPUT13), .ZN(n1327) );
XNOR2_X1 U1050 ( .A(G237), .B(KEYINPUT26), .ZN(n1345) );
NAND2_X1 U1051 ( .A1(n1346), .A2(n1317), .ZN(n1344) );
XNOR2_X1 U1052 ( .A(n1347), .B(n1348), .ZN(n1346) );
INV_X1 U1053 ( .A(n1162), .ZN(n1348) );
XNOR2_X1 U1054 ( .A(n1349), .B(n1350), .ZN(n1162) );
XOR2_X1 U1055 ( .A(n1351), .B(n1352), .Z(n1350) );
NOR2_X1 U1056 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
XOR2_X1 U1057 ( .A(n1355), .B(KEYINPUT16), .Z(n1354) );
NAND2_X1 U1058 ( .A1(G110), .A2(n1356), .ZN(n1355) );
NOR2_X1 U1059 ( .A1(G110), .A2(n1356), .ZN(n1353) );
NOR2_X1 U1060 ( .A1(KEYINPUT61), .A2(n1357), .ZN(n1351) );
XNOR2_X1 U1061 ( .A(KEYINPUT14), .B(n1298), .ZN(n1357) );
XOR2_X1 U1062 ( .A(n1339), .B(n1324), .Z(n1349) );
XOR2_X1 U1063 ( .A(G116), .B(G119), .Z(n1324) );
XNOR2_X1 U1064 ( .A(G101), .B(n1358), .ZN(n1339) );
XOR2_X1 U1065 ( .A(G107), .B(G104), .Z(n1358) );
XOR2_X1 U1066 ( .A(n1359), .B(KEYINPUT49), .Z(n1347) );
NAND2_X1 U1067 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NAND2_X1 U1068 ( .A1(n1362), .A2(n1227), .ZN(n1361) );
XOR2_X1 U1069 ( .A(KEYINPUT62), .B(n1363), .Z(n1360) );
NOR2_X1 U1070 ( .A1(n1362), .A2(n1227), .ZN(n1363) );
NAND2_X1 U1071 ( .A1(G224), .A2(n1091), .ZN(n1227) );
XNOR2_X1 U1072 ( .A(G125), .B(n1364), .ZN(n1362) );
NOR2_X1 U1073 ( .A1(KEYINPUT55), .A2(n1326), .ZN(n1364) );
INV_X1 U1074 ( .A(n1194), .ZN(n1326) );
XOR2_X1 U1075 ( .A(G143), .B(n1307), .Z(n1194) );
XNOR2_X1 U1076 ( .A(G146), .B(G128), .ZN(n1307) );
NOR2_X1 U1077 ( .A1(n1265), .A2(n1266), .ZN(n1092) );
XOR2_X1 U1078 ( .A(n1365), .B(n1183), .Z(n1266) );
INV_X1 U1079 ( .A(G475), .ZN(n1183) );
NAND2_X1 U1080 ( .A1(KEYINPUT51), .A2(n1366), .ZN(n1365) );
INV_X1 U1081 ( .A(n1126), .ZN(n1366) );
NAND2_X1 U1082 ( .A1(n1180), .A2(n1317), .ZN(n1126) );
INV_X1 U1083 ( .A(G902), .ZN(n1317) );
XNOR2_X1 U1084 ( .A(n1367), .B(n1368), .ZN(n1180) );
XOR2_X1 U1085 ( .A(G104), .B(n1369), .Z(n1368) );
NOR2_X1 U1086 ( .A1(KEYINPUT17), .A2(n1370), .ZN(n1369) );
NOR2_X1 U1087 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
NOR2_X1 U1088 ( .A1(G122), .A2(n1373), .ZN(n1372) );
NOR2_X1 U1089 ( .A1(n1374), .A2(KEYINPUT2), .ZN(n1373) );
NOR2_X1 U1090 ( .A1(G113), .A2(n1375), .ZN(n1374) );
NOR2_X1 U1091 ( .A1(n1376), .A2(n1298), .ZN(n1371) );
INV_X1 U1092 ( .A(G113), .ZN(n1298) );
NOR2_X1 U1093 ( .A1(n1377), .A2(n1375), .ZN(n1376) );
INV_X1 U1094 ( .A(KEYINPUT8), .ZN(n1375) );
NOR2_X1 U1095 ( .A1(KEYINPUT2), .A2(n1356), .ZN(n1377) );
INV_X1 U1096 ( .A(G122), .ZN(n1356) );
NAND3_X1 U1097 ( .A1(n1378), .A2(n1379), .A3(n1380), .ZN(n1367) );
NAND2_X1 U1098 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
INV_X1 U1099 ( .A(KEYINPUT4), .ZN(n1382) );
NAND3_X1 U1100 ( .A1(KEYINPUT4), .A2(n1383), .A3(n1384), .ZN(n1379) );
OR2_X1 U1101 ( .A1(n1384), .A2(n1383), .ZN(n1378) );
NOR2_X1 U1102 ( .A1(n1385), .A2(n1381), .ZN(n1383) );
XOR2_X1 U1103 ( .A(G146), .B(n1152), .Z(n1381) );
XNOR2_X1 U1104 ( .A(n1226), .B(G140), .ZN(n1152) );
INV_X1 U1105 ( .A(G125), .ZN(n1226) );
INV_X1 U1106 ( .A(KEYINPUT35), .ZN(n1385) );
XNOR2_X1 U1107 ( .A(n1386), .B(n1387), .ZN(n1384) );
XNOR2_X1 U1108 ( .A(n1388), .B(G131), .ZN(n1387) );
NAND2_X1 U1109 ( .A1(n1322), .A2(n1389), .ZN(n1386) );
XOR2_X1 U1110 ( .A(KEYINPUT37), .B(G214), .Z(n1389) );
NOR2_X1 U1111 ( .A1(G953), .A2(G237), .ZN(n1322) );
XNOR2_X1 U1112 ( .A(n1132), .B(n1128), .ZN(n1265) );
INV_X1 U1113 ( .A(G478), .ZN(n1128) );
NOR2_X1 U1114 ( .A1(n1175), .A2(G902), .ZN(n1132) );
INV_X1 U1115 ( .A(n1173), .ZN(n1175) );
NAND2_X1 U1116 ( .A1(n1390), .A2(n1391), .ZN(n1173) );
NAND2_X1 U1117 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
XOR2_X1 U1118 ( .A(n1394), .B(KEYINPUT18), .Z(n1390) );
OR2_X1 U1119 ( .A1(n1393), .A2(n1392), .ZN(n1394) );
XNOR2_X1 U1120 ( .A(n1395), .B(n1396), .ZN(n1392) );
XOR2_X1 U1121 ( .A(n1397), .B(n1398), .Z(n1396) );
NAND2_X1 U1122 ( .A1(KEYINPUT38), .A2(G107), .ZN(n1398) );
NAND2_X1 U1123 ( .A1(n1399), .A2(n1400), .ZN(n1397) );
NAND3_X1 U1124 ( .A1(n1401), .A2(n1402), .A3(n1403), .ZN(n1400) );
XNOR2_X1 U1125 ( .A(n1404), .B(n1338), .ZN(n1403) );
INV_X1 U1126 ( .A(G134), .ZN(n1338) );
NAND2_X1 U1127 ( .A1(KEYINPUT10), .A2(G143), .ZN(n1404) );
NAND2_X1 U1128 ( .A1(n1405), .A2(n1406), .ZN(n1399) );
NAND2_X1 U1129 ( .A1(n1401), .A2(n1402), .ZN(n1406) );
INV_X1 U1130 ( .A(KEYINPUT5), .ZN(n1402) );
INV_X1 U1131 ( .A(G128), .ZN(n1401) );
XNOR2_X1 U1132 ( .A(G134), .B(n1407), .ZN(n1405) );
AND2_X1 U1133 ( .A1(n1388), .A2(KEYINPUT10), .ZN(n1407) );
INV_X1 U1134 ( .A(G143), .ZN(n1388) );
XNOR2_X1 U1135 ( .A(G116), .B(G122), .ZN(n1395) );
NAND3_X1 U1136 ( .A1(G217), .A2(n1091), .A3(G234), .ZN(n1393) );
INV_X1 U1137 ( .A(G953), .ZN(n1091) );
endmodule


