//Key = 0110101101100001110010100000011000010110110101100111011111100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421;

XOR2_X1 U777 ( .A(G107), .B(n1082), .Z(G9) );
NOR2_X1 U778 ( .A1(n1083), .A2(n1084), .ZN(G75) );
NOR3_X1 U779 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
NOR2_X1 U780 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR2_X1 U781 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
XOR2_X1 U782 ( .A(KEYINPUT52), .B(n1092), .Z(n1091) );
NOR4_X1 U783 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1092) );
NOR3_X1 U784 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1090) );
NOR2_X1 U785 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NOR2_X1 U786 ( .A1(n1101), .A2(n1095), .ZN(n1100) );
NOR2_X1 U787 ( .A1(n1102), .A2(n1094), .ZN(n1099) );
INV_X1 U788 ( .A(n1103), .ZN(n1094) );
NOR2_X1 U789 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NOR2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NAND3_X1 U791 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1085) );
NAND3_X1 U792 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1110) );
INV_X1 U793 ( .A(n1096), .ZN(n1113) );
NAND2_X1 U794 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NAND3_X1 U795 ( .A1(n1103), .A2(n1116), .A3(n1117), .ZN(n1115) );
NAND2_X1 U796 ( .A1(n1118), .A2(n1119), .ZN(n1114) );
NAND2_X1 U797 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U798 ( .A1(n1103), .A2(n1122), .ZN(n1121) );
NAND2_X1 U799 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
OR2_X1 U800 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U801 ( .A1(n1117), .A2(n1127), .ZN(n1120) );
NOR3_X1 U802 ( .A1(n1128), .A2(G953), .A3(G952), .ZN(n1083) );
INV_X1 U803 ( .A(n1108), .ZN(n1128) );
NAND4_X1 U804 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1108) );
NOR4_X1 U805 ( .A1(n1133), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n1132) );
XOR2_X1 U806 ( .A(KEYINPUT14), .B(n1137), .Z(n1136) );
XNOR2_X1 U807 ( .A(n1138), .B(n1139), .ZN(n1135) );
NAND2_X1 U808 ( .A1(KEYINPUT46), .A2(n1140), .ZN(n1138) );
XNOR2_X1 U809 ( .A(n1141), .B(n1142), .ZN(n1134) );
NAND2_X1 U810 ( .A1(KEYINPUT1), .A2(n1143), .ZN(n1141) );
XOR2_X1 U811 ( .A(n1144), .B(n1145), .Z(n1133) );
XOR2_X1 U812 ( .A(KEYINPUT28), .B(G478), .Z(n1145) );
NOR2_X1 U813 ( .A1(KEYINPUT13), .A2(n1146), .ZN(n1144) );
NOR2_X1 U814 ( .A1(n1147), .A2(n1148), .ZN(n1131) );
XOR2_X1 U815 ( .A(n1149), .B(n1150), .Z(n1130) );
NAND2_X1 U816 ( .A1(KEYINPUT61), .A2(n1151), .ZN(n1150) );
XNOR2_X1 U817 ( .A(n1152), .B(n1153), .ZN(n1129) );
NOR2_X1 U818 ( .A1(n1154), .A2(KEYINPUT25), .ZN(n1153) );
XOR2_X1 U819 ( .A(n1155), .B(n1156), .Z(G72) );
XOR2_X1 U820 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR3_X1 U821 ( .A1(n1159), .A2(KEYINPUT36), .A3(n1160), .ZN(n1158) );
AND2_X1 U822 ( .A1(G227), .A2(G900), .ZN(n1160) );
XNOR2_X1 U823 ( .A(G953), .B(KEYINPUT33), .ZN(n1159) );
NAND2_X1 U824 ( .A1(n1161), .A2(n1109), .ZN(n1157) );
NAND2_X1 U825 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XNOR2_X1 U826 ( .A(KEYINPUT7), .B(n1164), .ZN(n1163) );
NAND2_X1 U827 ( .A1(n1165), .A2(n1166), .ZN(n1155) );
INV_X1 U828 ( .A(n1167), .ZN(n1166) );
NAND3_X1 U829 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1165) );
NAND2_X1 U830 ( .A1(KEYINPUT44), .A2(n1171), .ZN(n1170) );
INV_X1 U831 ( .A(n1172), .ZN(n1171) );
OR3_X1 U832 ( .A1(n1173), .A2(KEYINPUT44), .A3(n1174), .ZN(n1169) );
NAND2_X1 U833 ( .A1(n1174), .A2(n1173), .ZN(n1168) );
NAND2_X1 U834 ( .A1(KEYINPUT20), .A2(n1172), .ZN(n1173) );
XOR2_X1 U835 ( .A(n1175), .B(n1176), .Z(n1172) );
INV_X1 U836 ( .A(n1177), .ZN(n1176) );
NAND2_X1 U837 ( .A1(KEYINPUT6), .A2(n1178), .ZN(n1175) );
XOR2_X1 U838 ( .A(n1179), .B(n1180), .Z(G69) );
XOR2_X1 U839 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U840 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XNOR2_X1 U841 ( .A(n1185), .B(n1186), .ZN(n1184) );
XNOR2_X1 U842 ( .A(n1187), .B(n1188), .ZN(n1186) );
NOR2_X1 U843 ( .A1(KEYINPUT62), .A2(n1189), .ZN(n1188) );
INV_X1 U844 ( .A(n1190), .ZN(n1189) );
NOR2_X1 U845 ( .A1(G898), .A2(n1109), .ZN(n1183) );
NAND2_X1 U846 ( .A1(G953), .A2(n1191), .ZN(n1181) );
NAND2_X1 U847 ( .A1(G224), .A2(n1192), .ZN(n1191) );
XNOR2_X1 U848 ( .A(KEYINPUT24), .B(n1193), .ZN(n1192) );
NAND2_X1 U849 ( .A1(n1109), .A2(n1194), .ZN(n1179) );
NOR2_X1 U850 ( .A1(n1195), .A2(n1196), .ZN(G66) );
NOR2_X1 U851 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
XOR2_X1 U852 ( .A(n1199), .B(KEYINPUT51), .Z(n1198) );
NAND2_X1 U853 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
OR2_X1 U854 ( .A1(n1202), .A2(n1151), .ZN(n1201) );
XNOR2_X1 U855 ( .A(KEYINPUT22), .B(n1203), .ZN(n1200) );
NOR3_X1 U856 ( .A1(n1202), .A2(n1203), .A3(n1151), .ZN(n1197) );
NOR2_X1 U857 ( .A1(n1195), .A2(n1204), .ZN(G63) );
XNOR2_X1 U858 ( .A(n1205), .B(n1206), .ZN(n1204) );
AND2_X1 U859 ( .A1(G478), .A2(n1207), .ZN(n1206) );
NOR2_X1 U860 ( .A1(n1195), .A2(n1208), .ZN(G60) );
NOR3_X1 U861 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1208) );
AND3_X1 U862 ( .A1(n1212), .A2(G475), .A3(n1207), .ZN(n1211) );
NOR2_X1 U863 ( .A1(n1213), .A2(n1212), .ZN(n1210) );
AND2_X1 U864 ( .A1(n1087), .A2(G475), .ZN(n1213) );
XNOR2_X1 U865 ( .A(G104), .B(n1214), .ZN(G6) );
NOR2_X1 U866 ( .A1(n1195), .A2(n1215), .ZN(G57) );
NOR3_X1 U867 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
NOR2_X1 U868 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NOR2_X1 U869 ( .A1(n1221), .A2(n1222), .ZN(n1219) );
XOR2_X1 U870 ( .A(KEYINPUT63), .B(n1223), .Z(n1222) );
NOR3_X1 U871 ( .A1(n1224), .A2(n1223), .A3(n1221), .ZN(n1217) );
INV_X1 U872 ( .A(n1220), .ZN(n1224) );
XOR2_X1 U873 ( .A(n1225), .B(n1226), .Z(n1220) );
AND2_X1 U874 ( .A1(n1221), .A2(n1223), .ZN(n1216) );
XNOR2_X1 U875 ( .A(n1227), .B(n1228), .ZN(n1223) );
XOR2_X1 U876 ( .A(n1229), .B(n1230), .Z(n1228) );
AND2_X1 U877 ( .A1(G472), .A2(n1207), .ZN(n1230) );
XNOR2_X1 U878 ( .A(n1177), .B(n1231), .ZN(n1227) );
INV_X1 U879 ( .A(KEYINPUT10), .ZN(n1221) );
NOR3_X1 U880 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(G54) );
AND2_X1 U881 ( .A1(KEYINPUT45), .A2(n1195), .ZN(n1234) );
NOR2_X1 U882 ( .A1(n1109), .A2(G952), .ZN(n1195) );
NOR3_X1 U883 ( .A1(KEYINPUT45), .A2(G953), .A3(G952), .ZN(n1233) );
XOR2_X1 U884 ( .A(n1235), .B(n1236), .Z(n1232) );
XOR2_X1 U885 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U886 ( .A(KEYINPUT59), .B(n1239), .Z(n1238) );
NOR2_X1 U887 ( .A1(KEYINPUT0), .A2(n1178), .ZN(n1237) );
XOR2_X1 U888 ( .A(n1240), .B(n1241), .Z(n1235) );
XNOR2_X1 U889 ( .A(n1242), .B(n1243), .ZN(n1240) );
AND2_X1 U890 ( .A1(G469), .A2(n1207), .ZN(n1243) );
INV_X1 U891 ( .A(n1202), .ZN(n1207) );
NOR2_X1 U892 ( .A1(n1244), .A2(n1245), .ZN(G51) );
XOR2_X1 U893 ( .A(n1246), .B(n1247), .Z(n1245) );
NOR2_X1 U894 ( .A1(n1152), .A2(n1202), .ZN(n1247) );
NAND2_X1 U895 ( .A1(G902), .A2(n1087), .ZN(n1202) );
NAND3_X1 U896 ( .A1(n1162), .A2(n1164), .A3(n1248), .ZN(n1087) );
INV_X1 U897 ( .A(n1194), .ZN(n1248) );
NAND4_X1 U898 ( .A1(n1249), .A2(n1214), .A3(n1250), .A4(n1251), .ZN(n1194) );
NOR4_X1 U899 ( .A1(n1252), .A2(n1253), .A3(n1254), .A4(n1082), .ZN(n1251) );
AND3_X1 U900 ( .A1(n1118), .A2(n1127), .A3(n1255), .ZN(n1082) );
NOR3_X1 U901 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1250) );
NOR2_X1 U902 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
INV_X1 U903 ( .A(KEYINPUT49), .ZN(n1259) );
NOR2_X1 U904 ( .A1(KEYINPUT49), .A2(n1261), .ZN(n1257) );
NAND4_X1 U905 ( .A1(n1262), .A2(n1123), .A3(n1263), .A4(n1264), .ZN(n1261) );
NOR3_X1 U906 ( .A1(n1095), .A2(n1265), .A3(n1098), .ZN(n1264) );
INV_X1 U907 ( .A(n1118), .ZN(n1098) );
INV_X1 U908 ( .A(n1111), .ZN(n1095) );
NAND3_X1 U909 ( .A1(n1255), .A2(n1118), .A3(n1266), .ZN(n1214) );
AND4_X1 U910 ( .A1(n1267), .A2(n1268), .A3(n1269), .A4(n1270), .ZN(n1162) );
NOR4_X1 U911 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1270) );
NOR4_X1 U912 ( .A1(n1275), .A2(n1276), .A3(n1117), .A4(n1277), .ZN(n1274) );
AND2_X1 U913 ( .A1(n1275), .A2(n1278), .ZN(n1273) );
INV_X1 U914 ( .A(KEYINPUT23), .ZN(n1275) );
NOR4_X1 U915 ( .A1(n1279), .A2(n1280), .A3(KEYINPUT15), .A4(n1281), .ZN(n1272) );
INV_X1 U916 ( .A(n1127), .ZN(n1281) );
NOR2_X1 U917 ( .A1(n1282), .A2(n1093), .ZN(n1271) );
NOR3_X1 U918 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1282) );
AND3_X1 U919 ( .A1(KEYINPUT15), .A2(n1127), .A3(n1286), .ZN(n1285) );
NOR3_X1 U920 ( .A1(n1101), .A2(n1287), .A3(n1288), .ZN(n1283) );
NOR2_X1 U921 ( .A1(KEYINPUT35), .A2(n1289), .ZN(n1288) );
NOR3_X1 U922 ( .A1(n1290), .A2(n1291), .A3(n1089), .ZN(n1289) );
AND2_X1 U923 ( .A1(n1280), .A2(KEYINPUT35), .ZN(n1287) );
NOR2_X1 U924 ( .A1(G952), .A2(n1292), .ZN(n1244) );
XNOR2_X1 U925 ( .A(G953), .B(KEYINPUT31), .ZN(n1292) );
XOR2_X1 U926 ( .A(n1293), .B(G146), .Z(G48) );
NAND2_X1 U927 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
OR2_X1 U928 ( .A1(n1164), .A2(KEYINPUT39), .ZN(n1295) );
NAND2_X1 U929 ( .A1(n1266), .A2(n1296), .ZN(n1164) );
NAND3_X1 U930 ( .A1(n1296), .A2(n1101), .A3(KEYINPUT39), .ZN(n1294) );
INV_X1 U931 ( .A(n1266), .ZN(n1101) );
XOR2_X1 U932 ( .A(G143), .B(n1297), .Z(G45) );
NOR2_X1 U933 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
INV_X1 U934 ( .A(n1284), .ZN(n1299) );
NOR4_X1 U935 ( .A1(n1300), .A2(n1277), .A3(n1123), .A4(n1265), .ZN(n1284) );
XNOR2_X1 U936 ( .A(n1279), .B(KEYINPUT19), .ZN(n1298) );
NAND2_X1 U937 ( .A1(n1301), .A2(n1302), .ZN(G42) );
NAND2_X1 U938 ( .A1(KEYINPUT42), .A2(n1303), .ZN(n1302) );
XOR2_X1 U939 ( .A(n1304), .B(n1278), .Z(n1301) );
NOR2_X1 U940 ( .A1(n1280), .A2(n1276), .ZN(n1278) );
OR2_X1 U941 ( .A1(n1303), .A2(KEYINPUT42), .ZN(n1304) );
XNOR2_X1 U942 ( .A(G137), .B(n1269), .ZN(G39) );
NAND3_X1 U943 ( .A1(n1103), .A2(n1305), .A3(n1286), .ZN(n1269) );
XNOR2_X1 U944 ( .A(G134), .B(n1306), .ZN(G36) );
NAND2_X1 U945 ( .A1(n1307), .A2(n1127), .ZN(n1306) );
XNOR2_X1 U946 ( .A(G131), .B(n1308), .ZN(G33) );
NAND2_X1 U947 ( .A1(n1307), .A2(n1266), .ZN(n1308) );
NOR2_X1 U948 ( .A1(n1280), .A2(n1093), .ZN(n1307) );
INV_X1 U949 ( .A(n1279), .ZN(n1093) );
INV_X1 U950 ( .A(n1286), .ZN(n1280) );
NOR2_X1 U951 ( .A1(n1089), .A2(n1277), .ZN(n1286) );
INV_X1 U952 ( .A(n1117), .ZN(n1089) );
NOR2_X1 U953 ( .A1(n1125), .A2(n1147), .ZN(n1117) );
XNOR2_X1 U954 ( .A(G128), .B(n1267), .ZN(G30) );
NAND2_X1 U955 ( .A1(n1296), .A2(n1127), .ZN(n1267) );
NOR3_X1 U956 ( .A1(n1123), .A2(n1309), .A3(n1277), .ZN(n1296) );
NAND2_X1 U957 ( .A1(n1105), .A2(n1290), .ZN(n1277) );
INV_X1 U958 ( .A(n1305), .ZN(n1309) );
XNOR2_X1 U959 ( .A(n1254), .B(n1310), .ZN(G3) );
NAND2_X1 U960 ( .A1(KEYINPUT2), .A2(G101), .ZN(n1310) );
AND3_X1 U961 ( .A1(n1279), .A2(n1255), .A3(n1103), .ZN(n1254) );
XNOR2_X1 U962 ( .A(G125), .B(n1268), .ZN(G27) );
NAND4_X1 U963 ( .A1(n1311), .A2(n1111), .A3(n1312), .A4(n1290), .ZN(n1268) );
NAND2_X1 U964 ( .A1(n1096), .A2(n1313), .ZN(n1290) );
NAND2_X1 U965 ( .A1(n1167), .A2(n1314), .ZN(n1313) );
NOR2_X1 U966 ( .A1(n1109), .A2(G900), .ZN(n1167) );
INV_X1 U967 ( .A(n1276), .ZN(n1311) );
NAND2_X1 U968 ( .A1(n1266), .A2(n1116), .ZN(n1276) );
XNOR2_X1 U969 ( .A(G122), .B(n1260), .ZN(G24) );
NAND4_X1 U970 ( .A1(n1263), .A2(n1315), .A3(n1118), .A4(n1316), .ZN(n1260) );
XOR2_X1 U971 ( .A(G119), .B(n1253), .Z(G21) );
AND3_X1 U972 ( .A1(n1103), .A2(n1305), .A3(n1315), .ZN(n1253) );
NAND2_X1 U973 ( .A1(n1317), .A2(n1318), .ZN(n1305) );
NAND2_X1 U974 ( .A1(n1279), .A2(n1319), .ZN(n1318) );
NAND3_X1 U975 ( .A1(n1320), .A2(n1321), .A3(KEYINPUT53), .ZN(n1317) );
XOR2_X1 U976 ( .A(G116), .B(n1256), .Z(G18) );
AND3_X1 U977 ( .A1(n1279), .A2(n1127), .A3(n1315), .ZN(n1256) );
NOR2_X1 U978 ( .A1(n1263), .A2(n1265), .ZN(n1127) );
INV_X1 U979 ( .A(n1316), .ZN(n1265) );
XNOR2_X1 U980 ( .A(G113), .B(n1249), .ZN(G15) );
NAND3_X1 U981 ( .A1(n1266), .A2(n1279), .A3(n1315), .ZN(n1249) );
AND3_X1 U982 ( .A1(n1312), .A2(n1262), .A3(n1111), .ZN(n1315) );
NOR2_X1 U983 ( .A1(n1106), .A2(n1148), .ZN(n1111) );
INV_X1 U984 ( .A(n1107), .ZN(n1148) );
NOR2_X1 U985 ( .A1(n1322), .A2(n1320), .ZN(n1279) );
NOR2_X1 U986 ( .A1(n1316), .A2(n1300), .ZN(n1266) );
XOR2_X1 U987 ( .A(G110), .B(n1252), .Z(G12) );
AND3_X1 U988 ( .A1(n1255), .A2(n1116), .A3(n1103), .ZN(n1252) );
NOR2_X1 U989 ( .A1(n1316), .A2(n1263), .ZN(n1103) );
INV_X1 U990 ( .A(n1300), .ZN(n1263) );
XOR2_X1 U991 ( .A(n1323), .B(n1143), .Z(n1300) );
INV_X1 U992 ( .A(n1209), .ZN(n1143) );
NOR2_X1 U993 ( .A1(n1212), .A2(G902), .ZN(n1209) );
XNOR2_X1 U994 ( .A(n1324), .B(n1325), .ZN(n1212) );
XOR2_X1 U995 ( .A(n1326), .B(n1327), .Z(n1325) );
XOR2_X1 U996 ( .A(G113), .B(G104), .Z(n1327) );
XNOR2_X1 U997 ( .A(KEYINPUT55), .B(n1328), .ZN(n1326) );
INV_X1 U998 ( .A(G131), .ZN(n1328) );
XOR2_X1 U999 ( .A(n1329), .B(n1330), .Z(n1324) );
XOR2_X1 U1000 ( .A(n1331), .B(n1332), .Z(n1330) );
AND2_X1 U1001 ( .A1(G214), .A2(n1333), .ZN(n1332) );
NOR2_X1 U1002 ( .A1(KEYINPUT12), .A2(n1334), .ZN(n1331) );
XOR2_X1 U1003 ( .A(KEYINPUT21), .B(G122), .Z(n1334) );
XNOR2_X1 U1004 ( .A(n1174), .B(n1335), .ZN(n1329) );
NAND2_X1 U1005 ( .A1(KEYINPUT41), .A2(n1142), .ZN(n1323) );
XOR2_X1 U1006 ( .A(G475), .B(KEYINPUT37), .Z(n1142) );
XNOR2_X1 U1007 ( .A(n1146), .B(G478), .ZN(n1316) );
NAND2_X1 U1008 ( .A1(n1205), .A2(n1336), .ZN(n1146) );
XNOR2_X1 U1009 ( .A(n1337), .B(n1338), .ZN(n1205) );
NOR2_X1 U1010 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
INV_X1 U1011 ( .A(G217), .ZN(n1340) );
NAND3_X1 U1012 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1337) );
NAND2_X1 U1013 ( .A1(KEYINPUT32), .A2(n1344), .ZN(n1343) );
NAND3_X1 U1014 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1342) );
INV_X1 U1015 ( .A(KEYINPUT32), .ZN(n1346) );
OR2_X1 U1016 ( .A1(n1347), .A2(n1345), .ZN(n1341) );
NOR2_X1 U1017 ( .A1(KEYINPUT47), .A2(n1344), .ZN(n1345) );
XNOR2_X1 U1018 ( .A(n1348), .B(n1349), .ZN(n1344) );
XOR2_X1 U1019 ( .A(KEYINPUT8), .B(G134), .Z(n1349) );
XNOR2_X1 U1020 ( .A(n1350), .B(n1351), .ZN(n1348) );
INV_X1 U1021 ( .A(G128), .ZN(n1351) );
NAND2_X1 U1022 ( .A1(KEYINPUT56), .A2(G143), .ZN(n1350) );
XNOR2_X1 U1023 ( .A(G107), .B(n1352), .ZN(n1347) );
XOR2_X1 U1024 ( .A(G122), .B(G116), .Z(n1352) );
NAND2_X1 U1025 ( .A1(n1353), .A2(n1354), .ZN(n1116) );
NAND2_X1 U1026 ( .A1(n1118), .A2(n1319), .ZN(n1354) );
INV_X1 U1027 ( .A(KEYINPUT53), .ZN(n1319) );
NOR2_X1 U1028 ( .A1(n1320), .A2(n1321), .ZN(n1118) );
INV_X1 U1029 ( .A(n1322), .ZN(n1321) );
NAND3_X1 U1030 ( .A1(n1322), .A2(n1320), .A3(KEYINPUT53), .ZN(n1353) );
XOR2_X1 U1031 ( .A(n1149), .B(n1151), .Z(n1320) );
NAND2_X1 U1032 ( .A1(G217), .A2(n1355), .ZN(n1151) );
NAND2_X1 U1033 ( .A1(n1203), .A2(n1336), .ZN(n1149) );
XOR2_X1 U1034 ( .A(n1356), .B(n1357), .Z(n1203) );
XOR2_X1 U1035 ( .A(n1358), .B(n1359), .Z(n1357) );
XOR2_X1 U1036 ( .A(G110), .B(n1360), .Z(n1359) );
NOR2_X1 U1037 ( .A1(KEYINPUT26), .A2(n1174), .ZN(n1360) );
XNOR2_X1 U1038 ( .A(G140), .B(n1361), .ZN(n1174) );
NOR2_X1 U1039 ( .A1(n1362), .A2(n1339), .ZN(n1358) );
NAND2_X1 U1040 ( .A1(G234), .A2(n1109), .ZN(n1339) );
INV_X1 U1041 ( .A(G221), .ZN(n1362) );
XOR2_X1 U1042 ( .A(n1363), .B(n1364), .Z(n1356) );
XOR2_X1 U1043 ( .A(G146), .B(G137), .Z(n1364) );
XNOR2_X1 U1044 ( .A(G119), .B(G128), .ZN(n1363) );
XOR2_X1 U1045 ( .A(n1140), .B(n1365), .Z(n1322) );
INV_X1 U1046 ( .A(n1139), .ZN(n1365) );
XOR2_X1 U1047 ( .A(G472), .B(KEYINPUT38), .Z(n1139) );
NAND3_X1 U1048 ( .A1(n1366), .A2(n1336), .A3(n1367), .ZN(n1140) );
NAND3_X1 U1049 ( .A1(KEYINPUT58), .A2(n1231), .A3(n1368), .ZN(n1367) );
XNOR2_X1 U1050 ( .A(n1369), .B(n1370), .ZN(n1368) );
NOR2_X1 U1051 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
INV_X1 U1052 ( .A(KEYINPUT54), .ZN(n1371) );
NAND2_X1 U1053 ( .A1(n1373), .A2(n1374), .ZN(n1366) );
NAND2_X1 U1054 ( .A1(KEYINPUT58), .A2(n1231), .ZN(n1374) );
XOR2_X1 U1055 ( .A(n1375), .B(n1376), .Z(n1231) );
NOR2_X1 U1056 ( .A1(G113), .A2(KEYINPUT11), .ZN(n1376) );
XNOR2_X1 U1057 ( .A(n1377), .B(n1378), .ZN(n1373) );
INV_X1 U1058 ( .A(n1369), .ZN(n1378) );
XNOR2_X1 U1059 ( .A(n1379), .B(n1380), .ZN(n1369) );
XNOR2_X1 U1060 ( .A(KEYINPUT17), .B(n1226), .ZN(n1380) );
INV_X1 U1061 ( .A(G101), .ZN(n1226) );
NAND2_X1 U1062 ( .A1(KEYINPUT29), .A2(n1225), .ZN(n1379) );
NAND2_X1 U1063 ( .A1(n1333), .A2(G210), .ZN(n1225) );
NOR2_X1 U1064 ( .A1(G953), .A2(G237), .ZN(n1333) );
NAND2_X1 U1065 ( .A1(KEYINPUT54), .A2(n1372), .ZN(n1377) );
XNOR2_X1 U1066 ( .A(n1381), .B(n1229), .ZN(n1372) );
NAND2_X1 U1067 ( .A1(KEYINPUT40), .A2(n1177), .ZN(n1381) );
AND3_X1 U1068 ( .A1(n1105), .A2(n1262), .A3(n1312), .ZN(n1255) );
INV_X1 U1069 ( .A(n1123), .ZN(n1312) );
NAND2_X1 U1070 ( .A1(n1382), .A2(n1125), .ZN(n1123) );
XNOR2_X1 U1071 ( .A(n1154), .B(n1152), .ZN(n1125) );
NAND2_X1 U1072 ( .A1(G210), .A2(n1383), .ZN(n1152) );
AND2_X1 U1073 ( .A1(n1384), .A2(n1336), .ZN(n1154) );
XOR2_X1 U1074 ( .A(n1246), .B(KEYINPUT9), .Z(n1384) );
XOR2_X1 U1075 ( .A(n1385), .B(n1386), .Z(n1246) );
XOR2_X1 U1076 ( .A(n1361), .B(n1185), .Z(n1386) );
XOR2_X1 U1077 ( .A(G110), .B(G122), .Z(n1185) );
XOR2_X1 U1078 ( .A(G125), .B(KEYINPUT43), .Z(n1361) );
XOR2_X1 U1079 ( .A(n1387), .B(n1388), .Z(n1385) );
XOR2_X1 U1080 ( .A(n1389), .B(n1229), .Z(n1388) );
AND2_X1 U1081 ( .A1(n1390), .A2(n1391), .ZN(n1229) );
NAND2_X1 U1082 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
NAND2_X1 U1083 ( .A1(KEYINPUT4), .A2(n1394), .ZN(n1393) );
NAND2_X1 U1084 ( .A1(KEYINPUT16), .A2(n1335), .ZN(n1394) );
INV_X1 U1085 ( .A(n1395), .ZN(n1335) );
NAND2_X1 U1086 ( .A1(n1395), .A2(n1396), .ZN(n1390) );
NAND2_X1 U1087 ( .A1(KEYINPUT16), .A2(n1397), .ZN(n1396) );
NAND2_X1 U1088 ( .A1(n1398), .A2(KEYINPUT4), .ZN(n1397) );
INV_X1 U1089 ( .A(n1392), .ZN(n1398) );
XOR2_X1 U1090 ( .A(G128), .B(KEYINPUT5), .Z(n1392) );
NOR2_X1 U1091 ( .A1(KEYINPUT48), .A2(n1399), .ZN(n1389) );
XNOR2_X1 U1092 ( .A(n1400), .B(n1401), .ZN(n1399) );
INV_X1 U1093 ( .A(n1187), .ZN(n1401) );
XOR2_X1 U1094 ( .A(G113), .B(n1375), .Z(n1187) );
XOR2_X1 U1095 ( .A(G116), .B(G119), .Z(n1375) );
NOR2_X1 U1096 ( .A1(KEYINPUT27), .A2(n1402), .ZN(n1400) );
XNOR2_X1 U1097 ( .A(n1190), .B(KEYINPUT50), .ZN(n1402) );
NAND2_X1 U1098 ( .A1(G224), .A2(n1109), .ZN(n1387) );
XNOR2_X1 U1099 ( .A(n1147), .B(KEYINPUT34), .ZN(n1382) );
INV_X1 U1100 ( .A(n1126), .ZN(n1147) );
NAND2_X1 U1101 ( .A1(G214), .A2(n1383), .ZN(n1126) );
NAND2_X1 U1102 ( .A1(n1403), .A2(n1336), .ZN(n1383) );
INV_X1 U1103 ( .A(G237), .ZN(n1403) );
NAND2_X1 U1104 ( .A1(n1096), .A2(n1404), .ZN(n1262) );
NAND3_X1 U1105 ( .A1(n1314), .A2(n1193), .A3(G953), .ZN(n1404) );
INV_X1 U1106 ( .A(G898), .ZN(n1193) );
AND2_X1 U1107 ( .A1(n1405), .A2(n1406), .ZN(n1314) );
XNOR2_X1 U1108 ( .A(KEYINPUT60), .B(n1336), .ZN(n1405) );
NAND3_X1 U1109 ( .A1(n1406), .A2(n1109), .A3(G952), .ZN(n1096) );
NAND2_X1 U1110 ( .A1(G237), .A2(G234), .ZN(n1406) );
INV_X1 U1111 ( .A(n1291), .ZN(n1105) );
NAND2_X1 U1112 ( .A1(n1106), .A2(n1107), .ZN(n1291) );
NAND2_X1 U1113 ( .A1(G221), .A2(n1355), .ZN(n1107) );
NAND2_X1 U1114 ( .A1(G234), .A2(n1336), .ZN(n1355) );
XNOR2_X1 U1115 ( .A(n1137), .B(KEYINPUT30), .ZN(n1106) );
XNOR2_X1 U1116 ( .A(n1407), .B(G469), .ZN(n1137) );
NAND2_X1 U1117 ( .A1(n1408), .A2(n1336), .ZN(n1407) );
INV_X1 U1118 ( .A(G902), .ZN(n1336) );
XOR2_X1 U1119 ( .A(n1242), .B(n1409), .Z(n1408) );
XOR2_X1 U1120 ( .A(n1410), .B(n1178), .Z(n1409) );
XNOR2_X1 U1121 ( .A(G128), .B(n1395), .ZN(n1178) );
XOR2_X1 U1122 ( .A(G143), .B(G146), .Z(n1395) );
NAND2_X1 U1123 ( .A1(n1411), .A2(n1412), .ZN(n1410) );
NAND2_X1 U1124 ( .A1(n1413), .A2(n1414), .ZN(n1412) );
NAND2_X1 U1125 ( .A1(n1415), .A2(n1416), .ZN(n1414) );
OR2_X1 U1126 ( .A1(n1241), .A2(KEYINPUT3), .ZN(n1416) );
INV_X1 U1127 ( .A(KEYINPUT18), .ZN(n1415) );
NAND2_X1 U1128 ( .A1(n1241), .A2(n1417), .ZN(n1411) );
NAND2_X1 U1129 ( .A1(n1418), .A2(n1419), .ZN(n1417) );
OR2_X1 U1130 ( .A1(n1413), .A2(KEYINPUT18), .ZN(n1419) );
XOR2_X1 U1131 ( .A(n1239), .B(KEYINPUT57), .Z(n1413) );
AND2_X1 U1132 ( .A1(G227), .A2(n1109), .ZN(n1239) );
INV_X1 U1133 ( .A(G953), .ZN(n1109) );
INV_X1 U1134 ( .A(KEYINPUT3), .ZN(n1418) );
XNOR2_X1 U1135 ( .A(G110), .B(n1303), .ZN(n1241) );
INV_X1 U1136 ( .A(G140), .ZN(n1303) );
XOR2_X1 U1137 ( .A(n1177), .B(n1190), .Z(n1242) );
XOR2_X1 U1138 ( .A(G101), .B(n1420), .Z(n1190) );
XOR2_X1 U1139 ( .A(G107), .B(G104), .Z(n1420) );
XOR2_X1 U1140 ( .A(G131), .B(n1421), .Z(n1177) );
XOR2_X1 U1141 ( .A(G137), .B(G134), .Z(n1421) );
endmodule


