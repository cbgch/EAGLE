//Key = 0001110000000110101010000000001011100101011001001100011111100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347;

XNOR2_X1 U730 ( .A(G107), .B(n1014), .ZN(G9) );
NOR2_X1 U731 ( .A1(n1015), .A2(n1016), .ZN(G75) );
NOR3_X1 U732 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1016) );
NOR2_X1 U733 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR2_X1 U734 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U735 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
INV_X1 U736 ( .A(KEYINPUT44), .ZN(n1025) );
NOR4_X1 U737 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n1024) );
NOR2_X1 U738 ( .A1(n1030), .A2(n1029), .ZN(n1022) );
NOR2_X1 U739 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U740 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR3_X1 U741 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1033) );
NOR2_X1 U742 ( .A1(n1038), .A2(n1027), .ZN(n1037) );
NOR2_X1 U743 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U744 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR3_X1 U745 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1036) );
XOR2_X1 U746 ( .A(n1028), .B(KEYINPUT47), .Z(n1043) );
NOR2_X1 U747 ( .A1(n1028), .A2(n1046), .ZN(n1035) );
NOR3_X1 U748 ( .A1(n1028), .A2(n1047), .A3(n1027), .ZN(n1031) );
NOR2_X1 U749 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U750 ( .A1(KEYINPUT44), .A2(n1026), .ZN(n1048) );
NAND3_X1 U751 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1017) );
NAND4_X1 U752 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
NOR2_X1 U753 ( .A1(n1057), .A2(n1027), .ZN(n1055) );
NOR2_X1 U754 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
AND2_X1 U755 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
INV_X1 U756 ( .A(n1029), .ZN(n1053) );
NOR3_X1 U757 ( .A1(n1062), .A2(G953), .A3(G952), .ZN(n1015) );
INV_X1 U758 ( .A(n1050), .ZN(n1062) );
NAND4_X1 U759 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1050) );
NOR4_X1 U760 ( .A1(n1067), .A2(n1060), .A3(n1068), .A4(n1069), .ZN(n1066) );
XOR2_X1 U761 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND2_X1 U762 ( .A1(KEYINPUT53), .A2(n1072), .ZN(n1070) );
NOR2_X1 U763 ( .A1(n1073), .A2(n1074), .ZN(n1068) );
NOR2_X1 U764 ( .A1(G902), .A2(n1075), .ZN(n1073) );
NOR2_X1 U765 ( .A1(n1028), .A2(n1076), .ZN(n1065) );
XOR2_X1 U766 ( .A(n1077), .B(n1078), .Z(n1064) );
NOR2_X1 U767 ( .A1(KEYINPUT51), .A2(n1079), .ZN(n1078) );
XOR2_X1 U768 ( .A(n1080), .B(KEYINPUT0), .Z(n1079) );
XOR2_X1 U769 ( .A(n1081), .B(KEYINPUT38), .Z(n1063) );
XOR2_X1 U770 ( .A(n1082), .B(n1083), .Z(G72) );
NOR2_X1 U771 ( .A1(n1084), .A2(n1051), .ZN(n1083) );
AND2_X1 U772 ( .A1(G227), .A2(G900), .ZN(n1084) );
NAND2_X1 U773 ( .A1(n1085), .A2(n1086), .ZN(n1082) );
NAND2_X1 U774 ( .A1(n1087), .A2(n1051), .ZN(n1086) );
XOR2_X1 U775 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND3_X1 U776 ( .A1(n1089), .A2(G900), .A3(G953), .ZN(n1085) );
AND2_X1 U777 ( .A1(n1090), .A2(KEYINPUT39), .ZN(n1089) );
XOR2_X1 U778 ( .A(n1091), .B(n1092), .Z(n1090) );
XOR2_X1 U779 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U780 ( .A(n1095), .B(G137), .Z(n1094) );
NAND2_X1 U781 ( .A1(KEYINPUT3), .A2(n1096), .ZN(n1095) );
XOR2_X1 U782 ( .A(KEYINPUT14), .B(G140), .Z(n1096) );
NAND2_X1 U783 ( .A1(KEYINPUT41), .A2(n1097), .ZN(n1093) );
INV_X1 U784 ( .A(G134), .ZN(n1097) );
XOR2_X1 U785 ( .A(n1098), .B(n1099), .Z(n1091) );
INV_X1 U786 ( .A(n1100), .ZN(n1099) );
NAND2_X1 U787 ( .A1(n1101), .A2(n1102), .ZN(G69) );
NAND3_X1 U788 ( .A1(n1103), .A2(n1104), .A3(G953), .ZN(n1102) );
XOR2_X1 U789 ( .A(n1105), .B(KEYINPUT25), .Z(n1101) );
NAND2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U791 ( .A1(n1108), .A2(n1104), .ZN(n1107) );
NAND2_X1 U792 ( .A1(n1109), .A2(n1110), .ZN(n1104) );
XOR2_X1 U793 ( .A(KEYINPUT32), .B(n1111), .Z(n1110) );
INV_X1 U794 ( .A(n1112), .ZN(n1109) );
NAND2_X1 U795 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
NAND3_X1 U796 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1112) );
NAND2_X1 U797 ( .A1(G953), .A2(n1116), .ZN(n1115) );
NAND2_X1 U798 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
NAND2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NAND2_X1 U800 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
INV_X1 U801 ( .A(KEYINPUT54), .ZN(n1122) );
NAND2_X1 U802 ( .A1(KEYINPUT54), .A2(n1123), .ZN(n1119) );
NAND2_X1 U803 ( .A1(n1121), .A2(n1124), .ZN(n1123) );
NAND3_X1 U804 ( .A1(n1121), .A2(n1124), .A3(n1125), .ZN(n1113) );
INV_X1 U805 ( .A(n1118), .ZN(n1125) );
XOR2_X1 U806 ( .A(n1126), .B(KEYINPUT37), .Z(n1118) );
INV_X1 U807 ( .A(KEYINPUT40), .ZN(n1124) );
NAND3_X1 U808 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1121) );
NAND2_X1 U809 ( .A1(KEYINPUT12), .A2(n1130), .ZN(n1128) );
NAND2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U811 ( .A(n1133), .B(n1134), .Z(n1131) );
NAND2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1127) );
INV_X1 U813 ( .A(KEYINPUT12), .ZN(n1136) );
NAND2_X1 U814 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
NAND2_X1 U815 ( .A1(KEYINPUT11), .A2(n1134), .ZN(n1138) );
NAND3_X1 U816 ( .A1(n1132), .A2(n1133), .A3(n1139), .ZN(n1137) );
INV_X1 U817 ( .A(KEYINPUT11), .ZN(n1133) );
AND2_X1 U818 ( .A1(n1051), .A2(n1140), .ZN(n1111) );
NAND2_X1 U819 ( .A1(G953), .A2(n1103), .ZN(n1106) );
NAND2_X1 U820 ( .A1(G898), .A2(G224), .ZN(n1103) );
NOR2_X1 U821 ( .A1(n1141), .A2(n1142), .ZN(G66) );
NOR3_X1 U822 ( .A1(n1071), .A2(n1143), .A3(n1144), .ZN(n1142) );
NOR3_X1 U823 ( .A1(n1145), .A2(n1072), .A3(n1146), .ZN(n1144) );
NOR2_X1 U824 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
NOR2_X1 U825 ( .A1(n1149), .A2(n1072), .ZN(n1147) );
NOR2_X1 U826 ( .A1(n1141), .A2(n1150), .ZN(G63) );
XNOR2_X1 U827 ( .A(n1151), .B(n1152), .ZN(n1150) );
NOR3_X1 U828 ( .A1(n1146), .A2(KEYINPUT24), .A3(n1153), .ZN(n1152) );
INV_X1 U829 ( .A(G478), .ZN(n1153) );
NOR2_X1 U830 ( .A1(n1141), .A2(n1154), .ZN(G60) );
XOR2_X1 U831 ( .A(n1155), .B(n1075), .Z(n1154) );
NOR2_X1 U832 ( .A1(n1074), .A2(n1146), .ZN(n1155) );
INV_X1 U833 ( .A(G475), .ZN(n1074) );
XNOR2_X1 U834 ( .A(G104), .B(n1156), .ZN(G6) );
NOR2_X1 U835 ( .A1(n1141), .A2(n1157), .ZN(G57) );
XOR2_X1 U836 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U837 ( .A1(KEYINPUT27), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U838 ( .A(n1161), .B(n1162), .ZN(n1160) );
XOR2_X1 U839 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U840 ( .A1(n1080), .A2(n1146), .ZN(n1164) );
NOR2_X1 U841 ( .A1(KEYINPUT19), .A2(n1165), .ZN(n1163) );
XNOR2_X1 U842 ( .A(n1166), .B(n1167), .ZN(n1165) );
XOR2_X1 U843 ( .A(n1168), .B(KEYINPUT56), .Z(n1167) );
NOR2_X1 U844 ( .A1(n1141), .A2(n1169), .ZN(G54) );
XOR2_X1 U845 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U846 ( .A(n1172), .B(n1166), .Z(n1171) );
XNOR2_X1 U847 ( .A(n1173), .B(n1174), .ZN(n1166) );
XOR2_X1 U848 ( .A(n1100), .B(n1175), .Z(n1172) );
XOR2_X1 U849 ( .A(n1176), .B(n1177), .Z(n1170) );
XOR2_X1 U850 ( .A(n1178), .B(n1179), .Z(n1176) );
NAND3_X1 U851 ( .A1(n1180), .A2(n1019), .A3(G469), .ZN(n1178) );
XOR2_X1 U852 ( .A(KEYINPUT36), .B(G902), .Z(n1180) );
NOR2_X1 U853 ( .A1(n1141), .A2(n1181), .ZN(G51) );
XOR2_X1 U854 ( .A(n1182), .B(n1183), .Z(n1181) );
XNOR2_X1 U855 ( .A(n1184), .B(n1185), .ZN(n1183) );
XNOR2_X1 U856 ( .A(n1186), .B(KEYINPUT63), .ZN(n1182) );
NAND3_X1 U857 ( .A1(n1187), .A2(n1188), .A3(KEYINPUT18), .ZN(n1186) );
INV_X1 U858 ( .A(n1146), .ZN(n1187) );
NAND2_X1 U859 ( .A1(G902), .A2(n1019), .ZN(n1146) );
INV_X1 U860 ( .A(n1149), .ZN(n1019) );
NOR2_X1 U861 ( .A1(n1140), .A2(n1088), .ZN(n1149) );
NAND2_X1 U862 ( .A1(n1189), .A2(n1190), .ZN(n1088) );
NOR4_X1 U863 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1190) );
AND4_X1 U864 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1189) );
NAND4_X1 U865 ( .A1(n1199), .A2(n1156), .A3(n1200), .A4(n1201), .ZN(n1140) );
AND4_X1 U866 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
NOR3_X1 U867 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1200) );
NOR4_X1 U868 ( .A1(n1209), .A2(n1210), .A3(n1027), .A4(n1211), .ZN(n1208) );
NAND3_X1 U869 ( .A1(n1040), .A2(n1212), .A3(n1213), .ZN(n1210) );
INV_X1 U870 ( .A(KEYINPUT17), .ZN(n1209) );
NOR2_X1 U871 ( .A1(KEYINPUT17), .A2(n1014), .ZN(n1207) );
NAND3_X1 U872 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1014) );
NOR2_X1 U873 ( .A1(n1216), .A2(n1046), .ZN(n1206) );
NAND3_X1 U874 ( .A1(n1215), .A2(n1214), .A3(n1049), .ZN(n1156) );
NAND2_X1 U875 ( .A1(n1217), .A2(n1218), .ZN(n1199) );
INV_X1 U876 ( .A(n1219), .ZN(n1217) );
NOR2_X1 U877 ( .A1(n1051), .A2(G952), .ZN(n1141) );
XOR2_X1 U878 ( .A(n1198), .B(n1220), .Z(G48) );
NOR2_X1 U879 ( .A1(G146), .A2(KEYINPUT15), .ZN(n1220) );
NAND3_X1 U880 ( .A1(n1049), .A2(n1059), .A3(n1221), .ZN(n1198) );
NAND2_X1 U881 ( .A1(n1222), .A2(n1223), .ZN(G45) );
NAND2_X1 U882 ( .A1(G143), .A2(n1197), .ZN(n1223) );
XOR2_X1 U883 ( .A(n1224), .B(KEYINPUT59), .Z(n1222) );
OR2_X1 U884 ( .A1(n1197), .A2(G143), .ZN(n1224) );
NAND2_X1 U885 ( .A1(n1225), .A2(n1226), .ZN(n1197) );
XOR2_X1 U886 ( .A(G140), .B(n1227), .Z(G42) );
NOR2_X1 U887 ( .A1(KEYINPUT21), .A2(n1196), .ZN(n1227) );
NAND3_X1 U888 ( .A1(n1228), .A2(n1040), .A3(n1229), .ZN(n1196) );
XOR2_X1 U889 ( .A(G137), .B(n1191), .Z(G39) );
AND3_X1 U890 ( .A1(n1228), .A2(n1054), .A3(n1221), .ZN(n1191) );
NAND2_X1 U891 ( .A1(n1230), .A2(n1231), .ZN(G36) );
NAND2_X1 U892 ( .A1(G134), .A2(n1195), .ZN(n1231) );
XOR2_X1 U893 ( .A(KEYINPUT20), .B(n1232), .Z(n1230) );
NOR2_X1 U894 ( .A1(G134), .A2(n1195), .ZN(n1232) );
NAND3_X1 U895 ( .A1(n1228), .A2(n1213), .A3(n1225), .ZN(n1195) );
XOR2_X1 U896 ( .A(G131), .B(n1194), .Z(G33) );
AND3_X1 U897 ( .A1(n1228), .A2(n1049), .A3(n1225), .ZN(n1194) );
AND3_X1 U898 ( .A1(n1040), .A2(n1233), .A3(n1234), .ZN(n1225) );
INV_X1 U899 ( .A(n1021), .ZN(n1228) );
NAND2_X1 U900 ( .A1(n1061), .A2(n1235), .ZN(n1021) );
XNOR2_X1 U901 ( .A(n1076), .B(KEYINPUT6), .ZN(n1061) );
NAND3_X1 U902 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(G30) );
NAND2_X1 U903 ( .A1(n1193), .A2(n1239), .ZN(n1238) );
NAND2_X1 U904 ( .A1(n1240), .A2(KEYINPUT33), .ZN(n1239) );
XOR2_X1 U905 ( .A(n1241), .B(KEYINPUT4), .Z(n1240) );
INV_X1 U906 ( .A(n1242), .ZN(n1193) );
NAND3_X1 U907 ( .A1(KEYINPUT33), .A2(n1242), .A3(G128), .ZN(n1237) );
NAND3_X1 U908 ( .A1(n1213), .A2(n1059), .A3(n1221), .ZN(n1242) );
AND4_X1 U909 ( .A1(n1045), .A2(n1040), .A3(n1243), .A4(n1233), .ZN(n1221) );
OR2_X1 U910 ( .A1(G128), .A2(KEYINPUT33), .ZN(n1236) );
XOR2_X1 U911 ( .A(G101), .B(n1244), .Z(G3) );
NOR2_X1 U912 ( .A1(n1245), .A2(n1216), .ZN(n1244) );
XOR2_X1 U913 ( .A(n1046), .B(KEYINPUT22), .Z(n1245) );
XOR2_X1 U914 ( .A(G125), .B(n1192), .Z(G27) );
AND3_X1 U915 ( .A1(n1056), .A2(n1059), .A3(n1229), .ZN(n1192) );
AND4_X1 U916 ( .A1(n1049), .A2(n1246), .A3(n1243), .A4(n1233), .ZN(n1229) );
NAND2_X1 U917 ( .A1(n1029), .A2(n1247), .ZN(n1233) );
NAND4_X1 U918 ( .A1(G953), .A2(G902), .A3(n1248), .A4(n1249), .ZN(n1247) );
INV_X1 U919 ( .A(G900), .ZN(n1249) );
XNOR2_X1 U920 ( .A(G122), .B(n1205), .ZN(G24) );
NAND3_X1 U921 ( .A1(n1218), .A2(n1215), .A3(n1226), .ZN(n1205) );
AND3_X1 U922 ( .A1(n1059), .A2(n1250), .A3(n1251), .ZN(n1226) );
XOR2_X1 U923 ( .A(KEYINPUT30), .B(n1252), .Z(n1251) );
INV_X1 U924 ( .A(n1027), .ZN(n1215) );
NAND2_X1 U925 ( .A1(n1044), .A2(n1246), .ZN(n1027) );
INV_X1 U926 ( .A(n1045), .ZN(n1246) );
NAND2_X1 U927 ( .A1(n1253), .A2(n1254), .ZN(G21) );
NAND2_X1 U928 ( .A1(G119), .A2(n1204), .ZN(n1254) );
XOR2_X1 U929 ( .A(KEYINPUT13), .B(n1255), .Z(n1253) );
NOR2_X1 U930 ( .A1(G119), .A2(n1204), .ZN(n1255) );
NAND3_X1 U931 ( .A1(n1045), .A2(n1218), .A3(n1256), .ZN(n1204) );
AND3_X1 U932 ( .A1(n1054), .A2(n1243), .A3(n1059), .ZN(n1256) );
INV_X1 U933 ( .A(n1044), .ZN(n1243) );
NAND2_X1 U934 ( .A1(n1257), .A2(n1258), .ZN(G18) );
OR2_X1 U935 ( .A1(n1259), .A2(G116), .ZN(n1258) );
NAND2_X1 U936 ( .A1(n1260), .A2(G116), .ZN(n1257) );
NAND2_X1 U937 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
OR2_X1 U938 ( .A1(n1203), .A2(KEYINPUT5), .ZN(n1262) );
NAND2_X1 U939 ( .A1(KEYINPUT5), .A2(n1259), .ZN(n1261) );
OR2_X1 U940 ( .A1(KEYINPUT50), .A2(n1203), .ZN(n1259) );
NAND4_X1 U941 ( .A1(n1234), .A2(n1218), .A3(n1213), .A4(n1059), .ZN(n1203) );
XOR2_X1 U942 ( .A(n1212), .B(KEYINPUT43), .Z(n1059) );
INV_X1 U943 ( .A(n1026), .ZN(n1213) );
NAND2_X1 U944 ( .A1(n1252), .A2(n1250), .ZN(n1026) );
AND2_X1 U945 ( .A1(n1056), .A2(n1211), .ZN(n1218) );
INV_X1 U946 ( .A(n1028), .ZN(n1056) );
XOR2_X1 U947 ( .A(n1263), .B(n1264), .Z(G15) );
NOR2_X1 U948 ( .A1(KEYINPUT28), .A2(n1265), .ZN(n1264) );
NOR3_X1 U949 ( .A1(n1266), .A2(n1028), .A3(n1219), .ZN(n1263) );
NAND3_X1 U950 ( .A1(n1234), .A2(n1212), .A3(n1049), .ZN(n1219) );
NOR2_X1 U951 ( .A1(n1250), .A2(n1252), .ZN(n1049) );
INV_X1 U952 ( .A(n1081), .ZN(n1250) );
INV_X1 U953 ( .A(n1046), .ZN(n1234) );
NAND2_X1 U954 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
NAND2_X1 U955 ( .A1(n1267), .A2(n1042), .ZN(n1028) );
XNOR2_X1 U956 ( .A(KEYINPUT46), .B(n1211), .ZN(n1266) );
XNOR2_X1 U957 ( .A(G110), .B(n1202), .ZN(G12) );
OR3_X1 U958 ( .A1(n1045), .A2(n1044), .A3(n1216), .ZN(n1202) );
NAND2_X1 U959 ( .A1(n1054), .A2(n1214), .ZN(n1216) );
AND3_X1 U960 ( .A1(n1212), .A2(n1211), .A3(n1040), .ZN(n1214) );
AND2_X1 U961 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U962 ( .A1(G221), .A2(n1268), .ZN(n1042) );
INV_X1 U963 ( .A(n1267), .ZN(n1041) );
XOR2_X1 U964 ( .A(n1269), .B(G469), .Z(n1267) );
NAND2_X1 U965 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XOR2_X1 U966 ( .A(n1272), .B(n1273), .Z(n1270) );
NOR2_X1 U967 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
NOR2_X1 U968 ( .A1(n1179), .A2(n1276), .ZN(n1275) );
XOR2_X1 U969 ( .A(KEYINPUT45), .B(n1177), .Z(n1276) );
INV_X1 U970 ( .A(n1277), .ZN(n1179) );
NOR2_X1 U971 ( .A1(n1177), .A2(n1277), .ZN(n1274) );
NAND2_X1 U972 ( .A1(G227), .A2(n1051), .ZN(n1277) );
XNOR2_X1 U973 ( .A(n1174), .B(n1278), .ZN(n1272) );
NOR2_X1 U974 ( .A1(KEYINPUT29), .A2(n1279), .ZN(n1278) );
XOR2_X1 U975 ( .A(n1100), .B(n1280), .Z(n1279) );
XOR2_X1 U976 ( .A(G146), .B(n1281), .Z(n1280) );
NOR2_X1 U977 ( .A1(KEYINPUT1), .A2(n1175), .ZN(n1281) );
XOR2_X1 U978 ( .A(G101), .B(n1282), .Z(n1175) );
NOR2_X1 U979 ( .A1(KEYINPUT35), .A2(n1283), .ZN(n1282) );
XOR2_X1 U980 ( .A(n1284), .B(G143), .Z(n1100) );
NAND2_X1 U981 ( .A1(KEYINPUT57), .A2(G128), .ZN(n1284) );
NAND2_X1 U982 ( .A1(n1285), .A2(n1029), .ZN(n1211) );
NAND3_X1 U983 ( .A1(n1248), .A2(n1051), .A3(G952), .ZN(n1029) );
NAND4_X1 U984 ( .A1(G953), .A2(G902), .A3(n1248), .A4(n1116), .ZN(n1285) );
INV_X1 U985 ( .A(G898), .ZN(n1116) );
NAND2_X1 U986 ( .A1(G237), .A2(G234), .ZN(n1248) );
AND2_X1 U987 ( .A1(n1235), .A2(n1076), .ZN(n1212) );
XNOR2_X1 U988 ( .A(n1286), .B(n1188), .ZN(n1076) );
AND2_X1 U989 ( .A1(G210), .A2(n1287), .ZN(n1188) );
NAND3_X1 U990 ( .A1(n1288), .A2(n1271), .A3(n1289), .ZN(n1286) );
XOR2_X1 U991 ( .A(n1290), .B(KEYINPUT31), .Z(n1289) );
NAND2_X1 U992 ( .A1(n1185), .A2(n1184), .ZN(n1290) );
OR2_X1 U993 ( .A1(n1184), .A2(n1185), .ZN(n1288) );
NAND2_X1 U994 ( .A1(n1291), .A2(n1292), .ZN(n1185) );
NAND2_X1 U995 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
NAND2_X1 U996 ( .A1(n1129), .A2(n1295), .ZN(n1294) );
NAND2_X1 U997 ( .A1(n1132), .A2(n1139), .ZN(n1295) );
OR2_X1 U998 ( .A1(n1139), .A2(n1132), .ZN(n1129) );
INV_X1 U999 ( .A(n1126), .ZN(n1293) );
NAND2_X1 U1000 ( .A1(n1296), .A2(n1126), .ZN(n1291) );
XNOR2_X1 U1001 ( .A(G110), .B(n1297), .ZN(n1126) );
XOR2_X1 U1002 ( .A(KEYINPUT61), .B(G122), .Z(n1297) );
XOR2_X1 U1003 ( .A(n1139), .B(n1132), .Z(n1296) );
XOR2_X1 U1004 ( .A(G101), .B(n1298), .Z(n1132) );
NOR2_X1 U1005 ( .A1(KEYINPUT26), .A2(n1283), .ZN(n1298) );
XNOR2_X1 U1006 ( .A(G104), .B(G107), .ZN(n1283) );
INV_X1 U1007 ( .A(n1134), .ZN(n1139) );
XOR2_X1 U1008 ( .A(n1299), .B(n1300), .Z(n1134) );
XOR2_X1 U1009 ( .A(G119), .B(G113), .Z(n1300) );
NAND2_X1 U1010 ( .A1(KEYINPUT48), .A2(G116), .ZN(n1299) );
XNOR2_X1 U1011 ( .A(n1301), .B(n1302), .ZN(n1184) );
XOR2_X1 U1012 ( .A(n1303), .B(n1304), .Z(n1301) );
NAND2_X1 U1013 ( .A1(G224), .A2(n1051), .ZN(n1303) );
XNOR2_X1 U1014 ( .A(n1060), .B(KEYINPUT23), .ZN(n1235) );
AND2_X1 U1015 ( .A1(G214), .A2(n1287), .ZN(n1060) );
OR2_X1 U1016 ( .A1(G902), .A2(G237), .ZN(n1287) );
INV_X1 U1017 ( .A(n1034), .ZN(n1054) );
NAND2_X1 U1018 ( .A1(n1081), .A2(n1252), .ZN(n1034) );
NOR2_X1 U1019 ( .A1(n1305), .A2(n1067), .ZN(n1252) );
NOR3_X1 U1020 ( .A1(G475), .A2(G902), .A3(n1075), .ZN(n1067) );
AND2_X1 U1021 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
OR2_X1 U1022 ( .A1(n1075), .A2(G902), .ZN(n1307) );
XNOR2_X1 U1023 ( .A(n1308), .B(n1309), .ZN(n1075) );
XOR2_X1 U1024 ( .A(n1098), .B(n1310), .Z(n1309) );
XOR2_X1 U1025 ( .A(n1311), .B(n1312), .Z(n1310) );
NOR2_X1 U1026 ( .A1(KEYINPUT8), .A2(n1313), .ZN(n1312) );
XNOR2_X1 U1027 ( .A(G104), .B(n1314), .ZN(n1313) );
XOR2_X1 U1028 ( .A(G122), .B(G113), .Z(n1314) );
NAND2_X1 U1029 ( .A1(G214), .A2(n1315), .ZN(n1311) );
XNOR2_X1 U1030 ( .A(G131), .B(n1304), .ZN(n1098) );
XNOR2_X1 U1031 ( .A(G140), .B(n1316), .ZN(n1308) );
XOR2_X1 U1032 ( .A(KEYINPUT16), .B(G143), .Z(n1316) );
XOR2_X1 U1033 ( .A(KEYINPUT10), .B(G475), .Z(n1306) );
XOR2_X1 U1034 ( .A(n1317), .B(G478), .Z(n1081) );
NAND2_X1 U1035 ( .A1(n1151), .A2(n1271), .ZN(n1317) );
XNOR2_X1 U1036 ( .A(n1318), .B(n1319), .ZN(n1151) );
XOR2_X1 U1037 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1038 ( .A(G128), .B(G122), .Z(n1321) );
XOR2_X1 U1039 ( .A(G143), .B(G134), .Z(n1320) );
XOR2_X1 U1040 ( .A(n1322), .B(n1323), .Z(n1318) );
XOR2_X1 U1041 ( .A(G116), .B(G107), .Z(n1323) );
NAND3_X1 U1042 ( .A1(n1324), .A2(G217), .A3(KEYINPUT55), .ZN(n1322) );
XNOR2_X1 U1043 ( .A(n1325), .B(n1072), .ZN(n1044) );
NAND2_X1 U1044 ( .A1(G217), .A2(n1268), .ZN(n1072) );
NAND2_X1 U1045 ( .A1(G234), .A2(n1271), .ZN(n1268) );
XNOR2_X1 U1046 ( .A(n1071), .B(KEYINPUT7), .ZN(n1325) );
NOR2_X1 U1047 ( .A1(n1148), .A2(G902), .ZN(n1071) );
INV_X1 U1048 ( .A(n1145), .ZN(n1148) );
XOR2_X1 U1049 ( .A(n1326), .B(n1327), .Z(n1145) );
XOR2_X1 U1050 ( .A(n1328), .B(n1329), .Z(n1327) );
XOR2_X1 U1051 ( .A(G128), .B(G119), .Z(n1329) );
XOR2_X1 U1052 ( .A(KEYINPUT42), .B(G137), .Z(n1328) );
XOR2_X1 U1053 ( .A(n1330), .B(n1177), .Z(n1326) );
XOR2_X1 U1054 ( .A(G110), .B(G140), .Z(n1177) );
XOR2_X1 U1055 ( .A(n1331), .B(n1304), .Z(n1330) );
XNOR2_X1 U1056 ( .A(G125), .B(n1173), .ZN(n1304) );
NAND2_X1 U1057 ( .A1(G221), .A2(n1324), .ZN(n1331) );
AND2_X1 U1058 ( .A1(G234), .A2(n1051), .ZN(n1324) );
INV_X1 U1059 ( .A(G953), .ZN(n1051) );
XNOR2_X1 U1060 ( .A(n1332), .B(n1077), .ZN(n1045) );
NAND2_X1 U1061 ( .A1(n1333), .A2(n1271), .ZN(n1077) );
INV_X1 U1062 ( .A(G902), .ZN(n1271) );
XOR2_X1 U1063 ( .A(n1334), .B(n1335), .Z(n1333) );
XNOR2_X1 U1064 ( .A(n1159), .B(n1174), .ZN(n1335) );
XNOR2_X1 U1065 ( .A(n1336), .B(n1337), .ZN(n1174) );
XOR2_X1 U1066 ( .A(G134), .B(n1338), .Z(n1337) );
NOR2_X1 U1067 ( .A1(G131), .A2(KEYINPUT52), .ZN(n1338) );
XNOR2_X1 U1068 ( .A(G137), .B(KEYINPUT9), .ZN(n1336) );
XNOR2_X1 U1069 ( .A(n1339), .B(G101), .ZN(n1159) );
NAND2_X1 U1070 ( .A1(G210), .A2(n1315), .ZN(n1339) );
NOR2_X1 U1071 ( .A1(G953), .A2(G237), .ZN(n1315) );
XNOR2_X1 U1072 ( .A(n1340), .B(n1341), .ZN(n1334) );
NAND2_X1 U1073 ( .A1(KEYINPUT58), .A2(n1161), .ZN(n1341) );
XOR2_X1 U1074 ( .A(n1342), .B(n1343), .Z(n1161) );
XOR2_X1 U1075 ( .A(KEYINPUT2), .B(G119), .Z(n1343) );
XOR2_X1 U1076 ( .A(n1265), .B(G116), .Z(n1342) );
INV_X1 U1077 ( .A(G113), .ZN(n1265) );
NAND2_X1 U1078 ( .A1(n1344), .A2(KEYINPUT34), .ZN(n1340) );
XOR2_X1 U1079 ( .A(n1173), .B(n1302), .Z(n1344) );
INV_X1 U1080 ( .A(n1168), .ZN(n1302) );
XOR2_X1 U1081 ( .A(n1241), .B(n1345), .Z(n1168) );
NOR2_X1 U1082 ( .A1(KEYINPUT60), .A2(n1346), .ZN(n1345) );
XOR2_X1 U1083 ( .A(n1347), .B(KEYINPUT62), .Z(n1346) );
INV_X1 U1084 ( .A(G143), .ZN(n1347) );
INV_X1 U1085 ( .A(G128), .ZN(n1241) );
INV_X1 U1086 ( .A(G146), .ZN(n1173) );
NAND2_X1 U1087 ( .A1(KEYINPUT49), .A2(n1080), .ZN(n1332) );
INV_X1 U1088 ( .A(G472), .ZN(n1080) );
endmodule


