//Key = 1000100011001111001011010111011100011001000000110011010011000011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360;

XOR2_X1 U753 ( .A(G107), .B(n1041), .Z(G9) );
NOR2_X1 U754 ( .A1(KEYINPUT1), .A2(n1042), .ZN(n1041) );
NOR2_X1 U755 ( .A1(n1043), .A2(n1044), .ZN(G75) );
NOR4_X1 U756 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1044) );
NOR2_X1 U757 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
XOR2_X1 U758 ( .A(KEYINPUT63), .B(n1051), .Z(n1050) );
AND4_X1 U759 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1051) );
XOR2_X1 U760 ( .A(KEYINPUT40), .B(n1056), .Z(n1046) );
NOR2_X1 U761 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U762 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U763 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U764 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U765 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U766 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR3_X1 U767 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1068) );
NOR3_X1 U768 ( .A1(n1049), .A2(n1072), .A3(n1073), .ZN(n1067) );
INV_X1 U769 ( .A(n1074), .ZN(n1049) );
NOR3_X1 U770 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1063) );
NOR3_X1 U771 ( .A1(n1076), .A2(n1078), .A3(n1066), .ZN(n1059) );
INV_X1 U772 ( .A(n1079), .ZN(n1066) );
NAND3_X1 U773 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1045) );
NAND3_X1 U774 ( .A1(n1079), .A2(n1083), .A3(n1055), .ZN(n1082) );
INV_X1 U775 ( .A(n1058), .ZN(n1055) );
NAND2_X1 U776 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U777 ( .A1(n1052), .A2(n1086), .ZN(n1085) );
NAND2_X1 U778 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U779 ( .A1(n1089), .A2(n1074), .ZN(n1088) );
NAND2_X1 U780 ( .A1(n1054), .A2(n1090), .ZN(n1087) );
NAND2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1084) );
INV_X1 U782 ( .A(n1076), .ZN(n1091) );
NAND2_X1 U783 ( .A1(n1074), .A2(n1054), .ZN(n1076) );
NOR3_X1 U784 ( .A1(n1093), .A2(G953), .A3(G952), .ZN(n1043) );
INV_X1 U785 ( .A(n1080), .ZN(n1093) );
NAND4_X1 U786 ( .A1(n1094), .A2(n1074), .A3(n1095), .A4(n1096), .ZN(n1080) );
NOR4_X1 U787 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
XOR2_X1 U788 ( .A(n1101), .B(n1102), .Z(n1100) );
NAND2_X1 U789 ( .A1(KEYINPUT12), .A2(n1103), .ZN(n1101) );
NOR2_X1 U790 ( .A1(n1104), .A2(n1105), .ZN(n1099) );
INV_X1 U791 ( .A(n1106), .ZN(n1097) );
NOR2_X1 U792 ( .A1(n1073), .A2(n1107), .ZN(n1095) );
INV_X1 U793 ( .A(n1108), .ZN(n1107) );
XOR2_X1 U794 ( .A(n1109), .B(KEYINPUT16), .Z(n1094) );
XOR2_X1 U795 ( .A(n1110), .B(n1111), .Z(G72) );
XOR2_X1 U796 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U797 ( .A1(n1114), .A2(n1081), .ZN(n1113) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U799 ( .A1(n1117), .A2(n1118), .ZN(n1112) );
NAND2_X1 U800 ( .A1(G953), .A2(n1116), .ZN(n1118) );
XOR2_X1 U801 ( .A(n1119), .B(n1120), .Z(n1117) );
XOR2_X1 U802 ( .A(n1121), .B(n1122), .Z(n1120) );
XNOR2_X1 U803 ( .A(G131), .B(G134), .ZN(n1122) );
XOR2_X1 U804 ( .A(n1123), .B(n1124), .Z(n1119) );
XOR2_X1 U805 ( .A(G140), .B(G137), .Z(n1124) );
XOR2_X1 U806 ( .A(KEYINPUT55), .B(KEYINPUT20), .Z(n1123) );
NAND2_X1 U807 ( .A1(n1081), .A2(n1125), .ZN(n1110) );
XOR2_X1 U808 ( .A(n1126), .B(n1127), .Z(G69) );
NOR2_X1 U809 ( .A1(n1128), .A2(n1081), .ZN(n1127) );
AND2_X1 U810 ( .A1(G224), .A2(G898), .ZN(n1128) );
NOR2_X1 U811 ( .A1(KEYINPUT19), .A2(n1129), .ZN(n1126) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U813 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NOR2_X1 U814 ( .A1(n1134), .A2(n1081), .ZN(n1132) );
XOR2_X1 U815 ( .A(n1135), .B(KEYINPUT53), .Z(n1134) );
NAND2_X1 U816 ( .A1(n1081), .A2(n1136), .ZN(n1130) );
NAND2_X1 U817 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U818 ( .A1(n1139), .A2(n1140), .ZN(G66) );
XOR2_X1 U819 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U820 ( .A1(n1105), .A2(n1143), .ZN(n1142) );
NOR2_X1 U821 ( .A1(n1139), .A2(n1144), .ZN(G63) );
XNOR2_X1 U822 ( .A(n1145), .B(n1146), .ZN(n1144) );
NOR2_X1 U823 ( .A1(n1147), .A2(n1143), .ZN(n1146) );
INV_X1 U824 ( .A(G478), .ZN(n1147) );
NOR2_X1 U825 ( .A1(n1139), .A2(n1148), .ZN(G60) );
NOR3_X1 U826 ( .A1(n1102), .A2(n1149), .A3(n1150), .ZN(n1148) );
NOR3_X1 U827 ( .A1(n1151), .A2(n1103), .A3(n1143), .ZN(n1150) );
INV_X1 U828 ( .A(G475), .ZN(n1103) );
INV_X1 U829 ( .A(n1152), .ZN(n1151) );
NOR2_X1 U830 ( .A1(n1153), .A2(n1152), .ZN(n1149) );
AND2_X1 U831 ( .A1(n1048), .A2(G475), .ZN(n1153) );
NAND2_X1 U832 ( .A1(n1154), .A2(n1155), .ZN(G6) );
NAND2_X1 U833 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U834 ( .A(KEYINPUT15), .B(n1158), .Z(n1154) );
NOR2_X1 U835 ( .A1(n1156), .A2(n1157), .ZN(n1158) );
INV_X1 U836 ( .A(G104), .ZN(n1157) );
AND2_X1 U837 ( .A1(n1159), .A2(n1090), .ZN(n1156) );
XNOR2_X1 U838 ( .A(n1160), .B(KEYINPUT13), .ZN(n1159) );
NOR2_X1 U839 ( .A1(n1139), .A2(n1161), .ZN(G57) );
XOR2_X1 U840 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U841 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR3_X1 U842 ( .A1(n1143), .A2(KEYINPUT11), .A3(n1166), .ZN(n1165) );
INV_X1 U843 ( .A(G472), .ZN(n1166) );
NOR2_X1 U844 ( .A1(n1139), .A2(n1167), .ZN(G54) );
XOR2_X1 U845 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U846 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U847 ( .A1(KEYINPUT56), .A2(n1172), .ZN(n1170) );
XOR2_X1 U848 ( .A(n1173), .B(n1174), .Z(n1168) );
NOR2_X1 U849 ( .A1(n1175), .A2(n1143), .ZN(n1174) );
INV_X1 U850 ( .A(G469), .ZN(n1175) );
XNOR2_X1 U851 ( .A(KEYINPUT7), .B(n1176), .ZN(n1173) );
NOR2_X1 U852 ( .A1(KEYINPUT24), .A2(n1177), .ZN(n1176) );
XOR2_X1 U853 ( .A(n1178), .B(n1179), .Z(n1177) );
XNOR2_X1 U854 ( .A(n1180), .B(n1181), .ZN(n1179) );
NOR2_X1 U855 ( .A1(KEYINPUT61), .A2(n1182), .ZN(n1180) );
XNOR2_X1 U856 ( .A(KEYINPUT31), .B(n1183), .ZN(n1182) );
NOR2_X1 U857 ( .A1(n1139), .A2(n1184), .ZN(G51) );
XNOR2_X1 U858 ( .A(n1133), .B(n1185), .ZN(n1184) );
XOR2_X1 U859 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U860 ( .A1(n1188), .A2(n1143), .ZN(n1187) );
NAND2_X1 U861 ( .A1(G902), .A2(n1048), .ZN(n1143) );
NAND3_X1 U862 ( .A1(n1137), .A2(n1189), .A3(n1190), .ZN(n1048) );
INV_X1 U863 ( .A(n1125), .ZN(n1190) );
NAND4_X1 U864 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1125) );
NOR4_X1 U865 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1194) );
NOR2_X1 U866 ( .A1(n1199), .A2(n1200), .ZN(n1193) );
NOR2_X1 U867 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
XNOR2_X1 U868 ( .A(KEYINPUT9), .B(n1138), .ZN(n1189) );
AND4_X1 U869 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1137) );
AND4_X1 U870 ( .A1(n1042), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1206) );
NAND3_X1 U871 ( .A1(n1210), .A2(n1054), .A3(n1211), .ZN(n1042) );
NAND2_X1 U872 ( .A1(n1160), .A2(n1090), .ZN(n1205) );
AND4_X1 U873 ( .A1(n1092), .A2(n1054), .A3(n1053), .A4(n1212), .ZN(n1160) );
NAND4_X1 U874 ( .A1(n1213), .A2(n1054), .A3(n1214), .A4(n1215), .ZN(n1203) );
INV_X1 U875 ( .A(n1070), .ZN(n1054) );
INV_X1 U876 ( .A(G210), .ZN(n1188) );
NOR2_X1 U877 ( .A1(KEYINPUT60), .A2(n1216), .ZN(n1186) );
XNOR2_X1 U878 ( .A(n1217), .B(n1218), .ZN(n1216) );
NAND2_X1 U879 ( .A1(n1219), .A2(KEYINPUT36), .ZN(n1217) );
XOR2_X1 U880 ( .A(n1121), .B(KEYINPUT47), .Z(n1219) );
NOR2_X1 U881 ( .A1(n1081), .A2(G952), .ZN(n1139) );
XOR2_X1 U882 ( .A(G146), .B(n1199), .Z(G48) );
AND3_X1 U883 ( .A1(n1053), .A2(n1073), .A3(n1220), .ZN(n1199) );
XOR2_X1 U884 ( .A(G143), .B(n1221), .Z(G45) );
NOR2_X1 U885 ( .A1(n1202), .A2(n1222), .ZN(n1221) );
XOR2_X1 U886 ( .A(KEYINPUT38), .B(n1201), .Z(n1222) );
NAND4_X1 U887 ( .A1(n1089), .A2(n1223), .A3(n1214), .A4(n1215), .ZN(n1202) );
INV_X1 U888 ( .A(n1224), .ZN(n1215) );
XOR2_X1 U889 ( .A(n1191), .B(n1225), .Z(G42) );
NAND2_X1 U890 ( .A1(KEYINPUT62), .A2(G140), .ZN(n1225) );
NAND4_X1 U891 ( .A1(n1092), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1191) );
XOR2_X1 U892 ( .A(n1229), .B(n1192), .Z(G39) );
NAND3_X1 U893 ( .A1(n1226), .A2(n1073), .A3(n1230), .ZN(n1192) );
XOR2_X1 U894 ( .A(G134), .B(n1196), .Z(G36) );
AND3_X1 U895 ( .A1(n1226), .A2(n1210), .A3(n1089), .ZN(n1196) );
XOR2_X1 U896 ( .A(G131), .B(n1198), .Z(G33) );
AND3_X1 U897 ( .A1(n1089), .A2(n1226), .A3(n1092), .ZN(n1198) );
AND3_X1 U898 ( .A1(n1053), .A2(n1231), .A3(n1074), .ZN(n1226) );
NOR2_X1 U899 ( .A1(n1071), .A2(n1232), .ZN(n1074) );
XOR2_X1 U900 ( .A(n1233), .B(n1234), .Z(G30) );
XOR2_X1 U901 ( .A(n1235), .B(KEYINPUT49), .Z(n1234) );
NAND2_X1 U902 ( .A1(KEYINPUT30), .A2(n1195), .ZN(n1233) );
AND3_X1 U903 ( .A1(n1210), .A2(n1223), .A3(n1236), .ZN(n1195) );
NOR3_X1 U904 ( .A1(n1227), .A2(n1072), .A3(n1201), .ZN(n1236) );
INV_X1 U905 ( .A(n1231), .ZN(n1201) );
NAND3_X1 U906 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(G3) );
OR2_X1 U907 ( .A1(n1204), .A2(G101), .ZN(n1239) );
NAND2_X1 U908 ( .A1(KEYINPUT32), .A2(n1240), .ZN(n1238) );
NAND2_X1 U909 ( .A1(G101), .A2(n1241), .ZN(n1240) );
XNOR2_X1 U910 ( .A(KEYINPUT50), .B(n1204), .ZN(n1241) );
NAND2_X1 U911 ( .A1(n1242), .A2(n1243), .ZN(n1237) );
INV_X1 U912 ( .A(KEYINPUT32), .ZN(n1243) );
NAND2_X1 U913 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
NAND3_X1 U914 ( .A1(KEYINPUT50), .A2(G101), .A3(n1204), .ZN(n1245) );
OR2_X1 U915 ( .A1(n1204), .A2(KEYINPUT50), .ZN(n1244) );
NAND3_X1 U916 ( .A1(n1211), .A2(n1052), .A3(n1089), .ZN(n1204) );
XOR2_X1 U917 ( .A(G125), .B(n1197), .Z(G27) );
AND3_X1 U918 ( .A1(n1227), .A2(n1220), .A3(n1079), .ZN(n1197) );
AND4_X1 U919 ( .A1(n1092), .A2(n1090), .A3(n1231), .A4(n1228), .ZN(n1220) );
NAND2_X1 U920 ( .A1(n1058), .A2(n1246), .ZN(n1231) );
NAND4_X1 U921 ( .A1(G953), .A2(G902), .A3(n1247), .A4(n1116), .ZN(n1246) );
INV_X1 U922 ( .A(G900), .ZN(n1116) );
XNOR2_X1 U923 ( .A(G122), .B(n1248), .ZN(G24) );
NAND3_X1 U924 ( .A1(n1249), .A2(n1213), .A3(n1250), .ZN(n1248) );
NOR3_X1 U925 ( .A1(n1251), .A2(n1224), .A3(n1109), .ZN(n1250) );
XNOR2_X1 U926 ( .A(KEYINPUT33), .B(KEYINPUT0), .ZN(n1251) );
XOR2_X1 U927 ( .A(n1070), .B(KEYINPUT51), .Z(n1249) );
NAND2_X1 U928 ( .A1(n1072), .A2(n1227), .ZN(n1070) );
NAND2_X1 U929 ( .A1(n1252), .A2(n1253), .ZN(G21) );
OR2_X1 U930 ( .A1(n1254), .A2(G119), .ZN(n1253) );
NAND2_X1 U931 ( .A1(G119), .A2(n1255), .ZN(n1252) );
NAND2_X1 U932 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
OR2_X1 U933 ( .A1(n1209), .A2(KEYINPUT23), .ZN(n1257) );
NAND2_X1 U934 ( .A1(KEYINPUT23), .A2(n1254), .ZN(n1256) );
OR2_X1 U935 ( .A1(KEYINPUT6), .A2(n1209), .ZN(n1254) );
NAND3_X1 U936 ( .A1(n1230), .A2(n1073), .A3(n1213), .ZN(n1209) );
INV_X1 U937 ( .A(n1227), .ZN(n1073) );
XNOR2_X1 U938 ( .A(G116), .B(n1208), .ZN(G18) );
NAND3_X1 U939 ( .A1(n1089), .A2(n1210), .A3(n1213), .ZN(n1208) );
INV_X1 U940 ( .A(n1078), .ZN(n1210) );
XOR2_X1 U941 ( .A(n1258), .B(n1207), .Z(G15) );
NAND3_X1 U942 ( .A1(n1092), .A2(n1089), .A3(n1213), .ZN(n1207) );
AND3_X1 U943 ( .A1(n1090), .A2(n1212), .A3(n1079), .ZN(n1213) );
NOR2_X1 U944 ( .A1(n1077), .A2(n1098), .ZN(n1079) );
XNOR2_X1 U945 ( .A(n1108), .B(KEYINPUT22), .ZN(n1077) );
NOR2_X1 U946 ( .A1(n1228), .A2(n1227), .ZN(n1089) );
NOR2_X1 U947 ( .A1(n1214), .A2(n1224), .ZN(n1092) );
XNOR2_X1 U948 ( .A(G110), .B(n1138), .ZN(G12) );
NAND3_X1 U949 ( .A1(n1227), .A2(n1211), .A3(n1230), .ZN(n1138) );
NOR2_X1 U950 ( .A1(n1062), .A2(n1072), .ZN(n1230) );
INV_X1 U951 ( .A(n1228), .ZN(n1072) );
NAND3_X1 U952 ( .A1(n1259), .A2(n1260), .A3(n1106), .ZN(n1228) );
NAND2_X1 U953 ( .A1(n1104), .A2(n1105), .ZN(n1106) );
NAND2_X1 U954 ( .A1(n1105), .A2(n1261), .ZN(n1260) );
OR3_X1 U955 ( .A1(n1105), .A2(n1104), .A3(n1261), .ZN(n1259) );
INV_X1 U956 ( .A(KEYINPUT46), .ZN(n1261) );
NOR2_X1 U957 ( .A1(n1141), .A2(G902), .ZN(n1104) );
XOR2_X1 U958 ( .A(n1262), .B(n1263), .Z(n1141) );
XOR2_X1 U959 ( .A(n1264), .B(n1265), .Z(n1263) );
XNOR2_X1 U960 ( .A(G110), .B(G146), .ZN(n1265) );
NAND2_X1 U961 ( .A1(KEYINPUT29), .A2(n1229), .ZN(n1264) );
INV_X1 U962 ( .A(G137), .ZN(n1229) );
XOR2_X1 U963 ( .A(n1266), .B(n1267), .Z(n1262) );
XOR2_X1 U964 ( .A(n1268), .B(n1269), .Z(n1267) );
NAND2_X1 U965 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U966 ( .A1(G140), .A2(n1272), .ZN(n1271) );
XOR2_X1 U967 ( .A(KEYINPUT57), .B(n1273), .Z(n1270) );
NOR2_X1 U968 ( .A1(G140), .A2(n1272), .ZN(n1273) );
NAND3_X1 U969 ( .A1(n1274), .A2(n1275), .A3(KEYINPUT14), .ZN(n1268) );
OR3_X1 U970 ( .A1(n1235), .A2(G119), .A3(KEYINPUT21), .ZN(n1275) );
NAND2_X1 U971 ( .A1(n1276), .A2(KEYINPUT21), .ZN(n1274) );
XOR2_X1 U972 ( .A(G119), .B(n1277), .Z(n1276) );
NOR2_X1 U973 ( .A1(G128), .A2(KEYINPUT52), .ZN(n1277) );
NAND2_X1 U974 ( .A1(n1278), .A2(G221), .ZN(n1266) );
NAND2_X1 U975 ( .A1(G217), .A2(n1279), .ZN(n1105) );
INV_X1 U976 ( .A(n1052), .ZN(n1062) );
NAND2_X1 U977 ( .A1(n1280), .A2(n1281), .ZN(n1052) );
OR2_X1 U978 ( .A1(n1078), .A2(KEYINPUT39), .ZN(n1281) );
NAND2_X1 U979 ( .A1(n1224), .A2(n1214), .ZN(n1078) );
INV_X1 U980 ( .A(n1109), .ZN(n1214) );
NAND3_X1 U981 ( .A1(n1224), .A2(n1109), .A3(KEYINPUT39), .ZN(n1280) );
XOR2_X1 U982 ( .A(n1282), .B(G478), .Z(n1109) );
NAND2_X1 U983 ( .A1(n1283), .A2(n1145), .ZN(n1282) );
NAND2_X1 U984 ( .A1(n1284), .A2(n1285), .ZN(n1145) );
NAND4_X1 U985 ( .A1(n1286), .A2(n1287), .A3(n1288), .A4(n1289), .ZN(n1285) );
NAND2_X1 U986 ( .A1(G217), .A2(n1278), .ZN(n1286) );
XOR2_X1 U987 ( .A(n1290), .B(KEYINPUT54), .Z(n1284) );
NAND3_X1 U988 ( .A1(n1278), .A2(n1291), .A3(G217), .ZN(n1290) );
NAND3_X1 U989 ( .A1(n1288), .A2(n1289), .A3(n1287), .ZN(n1291) );
OR2_X1 U990 ( .A1(n1292), .A2(KEYINPUT25), .ZN(n1287) );
NAND4_X1 U991 ( .A1(n1293), .A2(KEYINPUT25), .A3(n1292), .A4(n1294), .ZN(n1289) );
XNOR2_X1 U992 ( .A(G116), .B(n1295), .ZN(n1293) );
NAND2_X1 U993 ( .A1(n1296), .A2(n1297), .ZN(n1288) );
NAND2_X1 U994 ( .A1(n1292), .A2(n1294), .ZN(n1297) );
INV_X1 U995 ( .A(KEYINPUT41), .ZN(n1294) );
XNOR2_X1 U996 ( .A(G134), .B(n1298), .ZN(n1292) );
NOR2_X1 U997 ( .A1(KEYINPUT44), .A2(n1299), .ZN(n1298) );
XOR2_X1 U998 ( .A(G116), .B(n1295), .Z(n1296) );
AND2_X1 U999 ( .A1(G234), .A2(n1081), .ZN(n1278) );
XOR2_X1 U1000 ( .A(n1300), .B(KEYINPUT59), .Z(n1283) );
XNOR2_X1 U1001 ( .A(n1102), .B(n1301), .ZN(n1224) );
XOR2_X1 U1002 ( .A(KEYINPUT10), .B(G475), .Z(n1301) );
NOR2_X1 U1003 ( .A1(n1152), .A2(G902), .ZN(n1102) );
XOR2_X1 U1004 ( .A(n1302), .B(n1303), .Z(n1152) );
XOR2_X1 U1005 ( .A(n1304), .B(n1305), .Z(n1303) );
XOR2_X1 U1006 ( .A(G125), .B(G104), .Z(n1305) );
XOR2_X1 U1007 ( .A(G143), .B(G131), .Z(n1304) );
XOR2_X1 U1008 ( .A(n1306), .B(n1307), .Z(n1302) );
XOR2_X1 U1009 ( .A(n1308), .B(n1309), .Z(n1307) );
NOR2_X1 U1010 ( .A1(G140), .A2(KEYINPUT45), .ZN(n1309) );
NOR2_X1 U1011 ( .A1(G146), .A2(KEYINPUT3), .ZN(n1308) );
XOR2_X1 U1012 ( .A(n1310), .B(n1311), .Z(n1306) );
AND2_X1 U1013 ( .A1(G214), .A2(n1312), .ZN(n1311) );
NAND2_X1 U1014 ( .A1(n1313), .A2(KEYINPUT26), .ZN(n1310) );
XNOR2_X1 U1015 ( .A(G122), .B(n1314), .ZN(n1313) );
NOR2_X1 U1016 ( .A1(G113), .A2(KEYINPUT42), .ZN(n1314) );
AND2_X1 U1017 ( .A1(n1223), .A2(n1212), .ZN(n1211) );
NAND2_X1 U1018 ( .A1(n1058), .A2(n1315), .ZN(n1212) );
NAND4_X1 U1019 ( .A1(G953), .A2(G902), .A3(n1247), .A4(n1135), .ZN(n1315) );
INV_X1 U1020 ( .A(G898), .ZN(n1135) );
NAND3_X1 U1021 ( .A1(n1247), .A2(n1081), .A3(n1316), .ZN(n1058) );
XOR2_X1 U1022 ( .A(KEYINPUT2), .B(G952), .Z(n1316) );
NAND2_X1 U1023 ( .A1(G237), .A2(G234), .ZN(n1247) );
AND2_X1 U1024 ( .A1(n1090), .A2(n1053), .ZN(n1223) );
NOR2_X1 U1025 ( .A1(n1108), .A2(n1098), .ZN(n1053) );
INV_X1 U1026 ( .A(n1075), .ZN(n1098) );
NAND2_X1 U1027 ( .A1(G221), .A2(n1279), .ZN(n1075) );
NAND2_X1 U1028 ( .A1(G234), .A2(n1300), .ZN(n1279) );
XOR2_X1 U1029 ( .A(n1317), .B(G469), .Z(n1108) );
NAND2_X1 U1030 ( .A1(n1318), .A2(n1300), .ZN(n1317) );
XOR2_X1 U1031 ( .A(n1319), .B(n1320), .Z(n1318) );
XOR2_X1 U1032 ( .A(n1181), .B(n1321), .Z(n1320) );
NAND3_X1 U1033 ( .A1(n1322), .A2(n1323), .A3(n1324), .ZN(n1181) );
NAND2_X1 U1034 ( .A1(KEYINPUT17), .A2(n1325), .ZN(n1324) );
OR3_X1 U1035 ( .A1(n1326), .A2(KEYINPUT17), .A3(G101), .ZN(n1323) );
NAND2_X1 U1036 ( .A1(G101), .A2(n1326), .ZN(n1322) );
NAND2_X1 U1037 ( .A1(KEYINPUT8), .A2(n1327), .ZN(n1326) );
INV_X1 U1038 ( .A(n1325), .ZN(n1327) );
XOR2_X1 U1039 ( .A(n1328), .B(G107), .Z(n1325) );
NAND2_X1 U1040 ( .A1(KEYINPUT18), .A2(G104), .ZN(n1328) );
XOR2_X1 U1041 ( .A(n1329), .B(n1330), .Z(n1319) );
NOR2_X1 U1042 ( .A1(KEYINPUT5), .A2(n1171), .ZN(n1330) );
XNOR2_X1 U1043 ( .A(G110), .B(G140), .ZN(n1171) );
XNOR2_X1 U1044 ( .A(KEYINPUT31), .B(n1172), .ZN(n1329) );
NOR2_X1 U1045 ( .A1(n1115), .A2(G953), .ZN(n1172) );
INV_X1 U1046 ( .A(G227), .ZN(n1115) );
AND2_X1 U1047 ( .A1(n1071), .A2(n1069), .ZN(n1090) );
INV_X1 U1048 ( .A(n1232), .ZN(n1069) );
NOR2_X1 U1049 ( .A1(n1331), .A2(n1332), .ZN(n1232) );
INV_X1 U1050 ( .A(G214), .ZN(n1331) );
XNOR2_X1 U1051 ( .A(n1333), .B(n1334), .ZN(n1071) );
NOR2_X1 U1052 ( .A1(n1332), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1053 ( .A(KEYINPUT27), .B(G210), .Z(n1335) );
NOR2_X1 U1054 ( .A1(G902), .A2(G237), .ZN(n1332) );
NAND2_X1 U1055 ( .A1(n1336), .A2(n1300), .ZN(n1333) );
XNOR2_X1 U1056 ( .A(n1337), .B(n1133), .ZN(n1336) );
XNOR2_X1 U1057 ( .A(n1338), .B(n1339), .ZN(n1133) );
XOR2_X1 U1058 ( .A(G104), .B(n1340), .Z(n1339) );
XOR2_X1 U1059 ( .A(G113), .B(G110), .Z(n1340) );
XOR2_X1 U1060 ( .A(n1341), .B(n1295), .Z(n1338) );
XOR2_X1 U1061 ( .A(G107), .B(G122), .Z(n1295) );
XNOR2_X1 U1062 ( .A(G101), .B(n1342), .ZN(n1341) );
NOR2_X1 U1063 ( .A1(KEYINPUT48), .A2(n1343), .ZN(n1342) );
NAND2_X1 U1064 ( .A1(KEYINPUT4), .A2(n1344), .ZN(n1337) );
XOR2_X1 U1065 ( .A(n1121), .B(n1345), .Z(n1344) );
XNOR2_X1 U1066 ( .A(KEYINPUT37), .B(n1346), .ZN(n1345) );
NOR2_X1 U1067 ( .A1(KEYINPUT58), .A2(n1218), .ZN(n1346) );
NAND2_X1 U1068 ( .A1(G224), .A2(n1081), .ZN(n1218) );
INV_X1 U1069 ( .A(G953), .ZN(n1081) );
XOR2_X1 U1070 ( .A(n1178), .B(n1272), .Z(n1121) );
INV_X1 U1071 ( .A(G125), .ZN(n1272) );
XOR2_X1 U1072 ( .A(n1347), .B(G472), .Z(n1227) );
NAND2_X1 U1073 ( .A1(n1348), .A2(n1300), .ZN(n1347) );
INV_X1 U1074 ( .A(G902), .ZN(n1300) );
XOR2_X1 U1075 ( .A(n1162), .B(n1349), .Z(n1348) );
INV_X1 U1076 ( .A(n1164), .ZN(n1349) );
XOR2_X1 U1077 ( .A(n1321), .B(n1350), .Z(n1164) );
NOR2_X1 U1078 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
XOR2_X1 U1079 ( .A(KEYINPUT28), .B(n1353), .Z(n1352) );
NOR2_X1 U1080 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
XOR2_X1 U1081 ( .A(KEYINPUT34), .B(G113), .Z(n1355) );
NOR2_X1 U1082 ( .A1(n1343), .A2(n1356), .ZN(n1351) );
XOR2_X1 U1083 ( .A(KEYINPUT34), .B(n1258), .Z(n1356) );
INV_X1 U1084 ( .A(G113), .ZN(n1258) );
INV_X1 U1085 ( .A(n1354), .ZN(n1343) );
XOR2_X1 U1086 ( .A(G116), .B(G119), .Z(n1354) );
XNOR2_X1 U1087 ( .A(n1178), .B(n1183), .ZN(n1321) );
XNOR2_X1 U1088 ( .A(n1357), .B(n1358), .ZN(n1183) );
XOR2_X1 U1089 ( .A(G137), .B(n1359), .Z(n1358) );
NOR2_X1 U1090 ( .A1(G131), .A2(KEYINPUT43), .ZN(n1359) );
NAND2_X1 U1091 ( .A1(KEYINPUT35), .A2(G134), .ZN(n1357) );
XNOR2_X1 U1092 ( .A(G146), .B(n1299), .ZN(n1178) );
XOR2_X1 U1093 ( .A(G143), .B(n1235), .Z(n1299) );
INV_X1 U1094 ( .A(G128), .ZN(n1235) );
XOR2_X1 U1095 ( .A(n1360), .B(G101), .Z(n1162) );
NAND2_X1 U1096 ( .A1(n1312), .A2(G210), .ZN(n1360) );
NOR2_X1 U1097 ( .A1(G953), .A2(G237), .ZN(n1312) );
endmodule


