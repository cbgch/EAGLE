//Key = 0101111000000110010101001011010011011011001101100101001011011011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377;

XNOR2_X1 U748 ( .A(n1041), .B(n1042), .ZN(G9) );
NAND2_X1 U749 ( .A1(KEYINPUT33), .A2(n1043), .ZN(n1041) );
NOR2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(G75) );
XOR2_X1 U751 ( .A(n1046), .B(KEYINPUT51), .Z(n1045) );
NAND3_X1 U752 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
XNOR2_X1 U753 ( .A(G952), .B(KEYINPUT47), .ZN(n1049) );
NOR4_X1 U754 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1044) );
INV_X1 U755 ( .A(G952), .ZN(n1053) );
NOR3_X1 U756 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1052) );
NOR3_X1 U757 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1055) );
NOR3_X1 U758 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NOR2_X1 U759 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
INV_X1 U760 ( .A(n1065), .ZN(n1064) );
NOR2_X1 U761 ( .A1(n1066), .A2(n1067), .ZN(n1063) );
NOR3_X1 U762 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1058) );
NOR2_X1 U763 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U764 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U765 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
AND2_X1 U766 ( .A1(n1077), .A2(KEYINPUT43), .ZN(n1075) );
NOR2_X1 U767 ( .A1(n1078), .A2(n1062), .ZN(n1071) );
NOR2_X1 U768 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U769 ( .A1(n1081), .A2(KEYINPUT43), .ZN(n1057) );
NOR3_X1 U770 ( .A1(n1060), .A2(n1068), .A3(n1082), .ZN(n1081) );
INV_X1 U771 ( .A(n1083), .ZN(n1060) );
NAND3_X1 U772 ( .A1(n1047), .A2(n1048), .A3(n1084), .ZN(n1050) );
NAND4_X1 U773 ( .A1(n1083), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1084) );
NAND2_X1 U774 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U775 ( .A1(n1056), .A2(n1090), .ZN(n1089) );
NOR2_X1 U776 ( .A1(n1074), .A2(n1069), .ZN(n1083) );
INV_X1 U777 ( .A(n1091), .ZN(n1069) );
NAND4_X1 U778 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1047) );
NOR3_X1 U779 ( .A1(n1096), .A2(n1068), .A3(n1097), .ZN(n1095) );
XOR2_X1 U780 ( .A(G472), .B(n1098), .Z(n1097) );
NOR2_X1 U781 ( .A1(KEYINPUT16), .A2(n1099), .ZN(n1098) );
NAND3_X1 U782 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1096) );
XNOR2_X1 U783 ( .A(n1103), .B(KEYINPUT37), .ZN(n1102) );
OR2_X1 U784 ( .A1(G478), .A2(KEYINPUT13), .ZN(n1101) );
NAND3_X1 U785 ( .A1(G478), .A2(n1104), .A3(KEYINPUT13), .ZN(n1100) );
NOR3_X1 U786 ( .A1(n1105), .A2(n1106), .A3(n1056), .ZN(n1094) );
NOR2_X1 U787 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
XOR2_X1 U788 ( .A(n1109), .B(n1110), .Z(n1093) );
NAND2_X1 U789 ( .A1(KEYINPUT32), .A2(n1111), .ZN(n1110) );
XOR2_X1 U790 ( .A(KEYINPUT27), .B(n1112), .Z(n1092) );
AND2_X1 U791 ( .A1(n1108), .A2(n1107), .ZN(n1112) );
XOR2_X1 U792 ( .A(n1113), .B(KEYINPUT46), .Z(n1108) );
XOR2_X1 U793 ( .A(n1114), .B(n1115), .Z(G72) );
NOR2_X1 U794 ( .A1(KEYINPUT9), .A2(n1116), .ZN(n1115) );
XOR2_X1 U795 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U796 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XNOR2_X1 U797 ( .A(n1121), .B(n1122), .ZN(n1120) );
XOR2_X1 U798 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U799 ( .A1(KEYINPUT26), .A2(n1125), .ZN(n1123) );
XNOR2_X1 U800 ( .A(G131), .B(n1126), .ZN(n1125) );
NOR2_X1 U801 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR3_X1 U802 ( .A1(n1129), .A2(G137), .A3(n1130), .ZN(n1128) );
INV_X1 U803 ( .A(KEYINPUT7), .ZN(n1129) );
NOR2_X1 U804 ( .A1(KEYINPUT7), .A2(n1131), .ZN(n1127) );
NAND2_X1 U805 ( .A1(n1048), .A2(n1132), .ZN(n1117) );
NOR2_X1 U806 ( .A1(n1133), .A2(n1048), .ZN(n1114) );
XOR2_X1 U807 ( .A(n1134), .B(KEYINPUT59), .Z(n1133) );
NAND2_X1 U808 ( .A1(G900), .A2(G227), .ZN(n1134) );
XOR2_X1 U809 ( .A(n1135), .B(n1136), .Z(G69) );
XOR2_X1 U810 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR3_X1 U811 ( .A1(n1139), .A2(KEYINPUT23), .A3(n1140), .ZN(n1138) );
XOR2_X1 U812 ( .A(n1141), .B(n1142), .Z(n1139) );
XNOR2_X1 U813 ( .A(n1143), .B(n1144), .ZN(n1142) );
XOR2_X1 U814 ( .A(KEYINPUT25), .B(n1145), .Z(n1141) );
NAND2_X1 U815 ( .A1(n1146), .A2(n1147), .ZN(n1137) );
NAND2_X1 U816 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
INV_X1 U817 ( .A(n1150), .ZN(n1149) );
XOR2_X1 U818 ( .A(n1151), .B(KEYINPUT63), .Z(n1148) );
XNOR2_X1 U819 ( .A(G953), .B(KEYINPUT31), .ZN(n1146) );
NAND2_X1 U820 ( .A1(G953), .A2(n1152), .ZN(n1135) );
NAND2_X1 U821 ( .A1(G898), .A2(G224), .ZN(n1152) );
NOR2_X1 U822 ( .A1(n1153), .A2(n1154), .ZN(G66) );
XOR2_X1 U823 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND2_X1 U824 ( .A1(n1157), .A2(n1113), .ZN(n1155) );
INV_X1 U825 ( .A(n1158), .ZN(n1113) );
NOR3_X1 U826 ( .A1(n1153), .A2(n1159), .A3(n1160), .ZN(G63) );
AND4_X1 U827 ( .A1(n1161), .A2(KEYINPUT6), .A3(G478), .A4(n1157), .ZN(n1160) );
NOR2_X1 U828 ( .A1(n1161), .A2(n1162), .ZN(n1159) );
NOR3_X1 U829 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1162) );
INV_X1 U830 ( .A(G478), .ZN(n1165) );
NOR2_X1 U831 ( .A1(KEYINPUT6), .A2(n1166), .ZN(n1164) );
NOR2_X1 U832 ( .A1(n1167), .A2(KEYINPUT48), .ZN(n1161) );
INV_X1 U833 ( .A(n1166), .ZN(n1167) );
NOR2_X1 U834 ( .A1(n1153), .A2(n1168), .ZN(G60) );
XNOR2_X1 U835 ( .A(n1169), .B(n1170), .ZN(n1168) );
XOR2_X1 U836 ( .A(n1171), .B(KEYINPUT29), .Z(n1170) );
NAND2_X1 U837 ( .A1(n1157), .A2(G475), .ZN(n1171) );
XNOR2_X1 U838 ( .A(G104), .B(n1172), .ZN(G6) );
NOR2_X1 U839 ( .A1(n1153), .A2(n1173), .ZN(G57) );
XOR2_X1 U840 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U841 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U842 ( .A(KEYINPUT20), .B(n1178), .Z(n1177) );
AND2_X1 U843 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NAND2_X1 U844 ( .A1(n1181), .A2(n1182), .ZN(n1174) );
NAND4_X1 U845 ( .A1(n1183), .A2(G472), .A3(n1184), .A4(n1185), .ZN(n1182) );
XNOR2_X1 U846 ( .A(n1186), .B(n1187), .ZN(n1183) );
NAND2_X1 U847 ( .A1(n1188), .A2(n1189), .ZN(n1181) );
NAND3_X1 U848 ( .A1(n1184), .A2(n1185), .A3(G472), .ZN(n1189) );
NAND2_X1 U849 ( .A1(n1163), .A2(n1190), .ZN(n1185) );
INV_X1 U850 ( .A(KEYINPUT40), .ZN(n1190) );
NAND2_X1 U851 ( .A1(KEYINPUT40), .A2(n1191), .ZN(n1184) );
NAND2_X1 U852 ( .A1(n1192), .A2(n1051), .ZN(n1191) );
XNOR2_X1 U853 ( .A(n1187), .B(n1193), .ZN(n1188) );
NOR2_X1 U854 ( .A1(n1153), .A2(n1194), .ZN(G54) );
XOR2_X1 U855 ( .A(n1195), .B(n1196), .Z(n1194) );
XNOR2_X1 U856 ( .A(n1197), .B(n1198), .ZN(n1196) );
XOR2_X1 U857 ( .A(n1199), .B(n1200), .Z(n1195) );
XNOR2_X1 U858 ( .A(n1201), .B(n1202), .ZN(n1200) );
NAND2_X1 U859 ( .A1(n1157), .A2(G469), .ZN(n1201) );
NAND2_X1 U860 ( .A1(KEYINPUT14), .A2(n1203), .ZN(n1199) );
NOR2_X1 U861 ( .A1(n1153), .A2(n1204), .ZN(G51) );
XOR2_X1 U862 ( .A(n1205), .B(n1206), .Z(n1204) );
NAND2_X1 U863 ( .A1(n1157), .A2(n1207), .ZN(n1205) );
INV_X1 U864 ( .A(n1163), .ZN(n1157) );
NAND2_X1 U865 ( .A1(G902), .A2(n1051), .ZN(n1163) );
OR3_X1 U866 ( .A1(n1132), .A2(n1150), .A3(n1151), .ZN(n1051) );
NAND4_X1 U867 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1151) );
NAND4_X1 U868 ( .A1(n1212), .A2(n1213), .A3(n1042), .A4(n1172), .ZN(n1150) );
NAND2_X1 U869 ( .A1(n1080), .A2(n1214), .ZN(n1172) );
NAND2_X1 U870 ( .A1(n1079), .A2(n1214), .ZN(n1042) );
NOR3_X1 U871 ( .A1(n1062), .A2(n1215), .A3(n1216), .ZN(n1214) );
INV_X1 U872 ( .A(n1086), .ZN(n1062) );
NAND2_X1 U873 ( .A1(n1217), .A2(n1218), .ZN(n1213) );
INV_X1 U874 ( .A(n1219), .ZN(n1218) );
XOR2_X1 U875 ( .A(n1215), .B(KEYINPUT60), .Z(n1217) );
NAND2_X1 U876 ( .A1(n1220), .A2(n1221), .ZN(n1212) );
NAND4_X1 U877 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1132) );
NOR4_X1 U878 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1225) );
NAND2_X1 U879 ( .A1(KEYINPUT17), .A2(n1230), .ZN(n1224) );
NAND2_X1 U880 ( .A1(n1231), .A2(n1232), .ZN(n1222) );
NAND2_X1 U881 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND3_X1 U882 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1234) );
NAND2_X1 U883 ( .A1(n1103), .A2(n1238), .ZN(n1236) );
NAND3_X1 U884 ( .A1(n1239), .A2(n1240), .A3(n1077), .ZN(n1238) );
OR2_X1 U885 ( .A1(n1241), .A2(KEYINPUT55), .ZN(n1240) );
NAND2_X1 U886 ( .A1(KEYINPUT55), .A2(n1242), .ZN(n1239) );
NAND2_X1 U887 ( .A1(n1221), .A2(n1065), .ZN(n1242) );
NAND2_X1 U888 ( .A1(n1243), .A2(n1244), .ZN(n1235) );
OR3_X1 U889 ( .A1(n1245), .A2(KEYINPUT17), .A3(n1216), .ZN(n1244) );
INV_X1 U890 ( .A(n1241), .ZN(n1216) );
NOR2_X1 U891 ( .A1(n1048), .A2(G952), .ZN(n1153) );
XOR2_X1 U892 ( .A(G146), .B(n1229), .Z(G48) );
AND4_X1 U893 ( .A1(n1231), .A2(n1245), .A3(n1080), .A4(n1241), .ZN(n1229) );
XOR2_X1 U894 ( .A(G143), .B(n1246), .Z(G45) );
NOR4_X1 U895 ( .A1(KEYINPUT2), .A2(n1243), .A3(n1082), .A4(n1247), .ZN(n1246) );
XNOR2_X1 U896 ( .A(G140), .B(n1223), .ZN(G42) );
NAND3_X1 U897 ( .A1(n1248), .A2(n1080), .A3(n1076), .ZN(n1223) );
XOR2_X1 U898 ( .A(G137), .B(n1228), .Z(G39) );
AND3_X1 U899 ( .A1(n1249), .A2(n1245), .A3(n1248), .ZN(n1228) );
XNOR2_X1 U900 ( .A(n1130), .B(n1227), .ZN(G36) );
AND3_X1 U901 ( .A1(n1077), .A2(n1079), .A3(n1248), .ZN(n1227) );
XNOR2_X1 U902 ( .A(G131), .B(n1250), .ZN(G33) );
NAND2_X1 U903 ( .A1(KEYINPUT49), .A2(n1226), .ZN(n1250) );
AND3_X1 U904 ( .A1(n1080), .A2(n1077), .A3(n1248), .ZN(n1226) );
NOR4_X1 U905 ( .A1(n1054), .A2(n1251), .A3(n1065), .A4(n1056), .ZN(n1248) );
XOR2_X1 U906 ( .A(G128), .B(n1230), .Z(G30) );
NOR3_X1 U907 ( .A1(n1103), .A2(n1252), .A3(n1247), .ZN(n1230) );
NAND3_X1 U908 ( .A1(n1241), .A2(n1237), .A3(n1231), .ZN(n1247) );
XNOR2_X1 U909 ( .A(n1180), .B(n1253), .ZN(G3) );
NOR2_X1 U910 ( .A1(n1254), .A2(n1088), .ZN(n1253) );
XNOR2_X1 U911 ( .A(n1220), .B(KEYINPUT28), .ZN(n1254) );
NOR4_X1 U912 ( .A1(n1074), .A2(n1082), .A3(n1215), .A4(n1065), .ZN(n1220) );
INV_X1 U913 ( .A(n1249), .ZN(n1074) );
XNOR2_X1 U914 ( .A(G125), .B(n1255), .ZN(G27) );
NAND2_X1 U915 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
INV_X1 U916 ( .A(n1233), .ZN(n1257) );
NAND4_X1 U917 ( .A1(n1076), .A2(n1080), .A3(n1085), .A4(n1221), .ZN(n1233) );
INV_X1 U918 ( .A(n1068), .ZN(n1085) );
XNOR2_X1 U919 ( .A(n1231), .B(KEYINPUT54), .ZN(n1256) );
INV_X1 U920 ( .A(n1251), .ZN(n1231) );
NAND2_X1 U921 ( .A1(n1258), .A2(n1259), .ZN(n1251) );
NAND2_X1 U922 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
INV_X1 U923 ( .A(n1119), .ZN(n1260) );
NOR2_X1 U924 ( .A1(n1048), .A2(G900), .ZN(n1119) );
XNOR2_X1 U925 ( .A(G122), .B(n1209), .ZN(G24) );
NAND4_X1 U926 ( .A1(n1262), .A2(n1086), .A3(n1103), .A4(n1237), .ZN(n1209) );
NOR2_X1 U927 ( .A1(n1263), .A2(n1264), .ZN(n1086) );
XNOR2_X1 U928 ( .A(G119), .B(n1210), .ZN(G21) );
NAND3_X1 U929 ( .A1(n1245), .A2(n1262), .A3(n1249), .ZN(n1210) );
INV_X1 U930 ( .A(n1252), .ZN(n1245) );
NAND2_X1 U931 ( .A1(n1264), .A2(n1263), .ZN(n1252) );
INV_X1 U932 ( .A(n1265), .ZN(n1264) );
XNOR2_X1 U933 ( .A(G116), .B(n1266), .ZN(G18) );
NOR2_X1 U934 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NOR2_X1 U935 ( .A1(n1269), .A2(n1208), .ZN(n1268) );
NAND3_X1 U936 ( .A1(n1262), .A2(n1079), .A3(n1077), .ZN(n1208) );
INV_X1 U937 ( .A(KEYINPUT3), .ZN(n1269) );
NOR4_X1 U938 ( .A1(KEYINPUT3), .A2(n1270), .A3(n1068), .A4(n1082), .ZN(n1267) );
NAND3_X1 U939 ( .A1(n1221), .A2(n1215), .A3(n1079), .ZN(n1270) );
NOR2_X1 U940 ( .A1(n1103), .A2(n1271), .ZN(n1079) );
XNOR2_X1 U941 ( .A(G113), .B(n1211), .ZN(G15) );
NAND3_X1 U942 ( .A1(n1077), .A2(n1262), .A3(n1080), .ZN(n1211) );
NOR2_X1 U943 ( .A1(n1237), .A2(n1243), .ZN(n1080) );
INV_X1 U944 ( .A(n1103), .ZN(n1243) );
NOR3_X1 U945 ( .A1(n1215), .A2(n1088), .A3(n1068), .ZN(n1262) );
NAND2_X1 U946 ( .A1(n1272), .A2(n1067), .ZN(n1068) );
INV_X1 U947 ( .A(n1066), .ZN(n1272) );
INV_X1 U948 ( .A(n1082), .ZN(n1077) );
NAND2_X1 U949 ( .A1(n1263), .A2(n1265), .ZN(n1082) );
XNOR2_X1 U950 ( .A(n1203), .B(n1273), .ZN(G12) );
NOR2_X1 U951 ( .A1(n1215), .A2(n1219), .ZN(n1273) );
NAND3_X1 U952 ( .A1(n1249), .A2(n1241), .A3(n1076), .ZN(n1219) );
NOR2_X1 U953 ( .A1(n1265), .A2(n1263), .ZN(n1076) );
XNOR2_X1 U954 ( .A(n1099), .B(G472), .ZN(n1263) );
NAND2_X1 U955 ( .A1(n1274), .A2(n1192), .ZN(n1099) );
XOR2_X1 U956 ( .A(n1275), .B(n1276), .Z(n1274) );
NOR2_X1 U957 ( .A1(n1176), .A2(n1277), .ZN(n1276) );
NOR2_X1 U958 ( .A1(G101), .A2(n1278), .ZN(n1277) );
XOR2_X1 U959 ( .A(n1179), .B(KEYINPUT38), .Z(n1278) );
NOR2_X1 U960 ( .A1(n1179), .A2(n1180), .ZN(n1176) );
NAND3_X1 U961 ( .A1(n1279), .A2(n1048), .A3(G210), .ZN(n1179) );
NAND3_X1 U962 ( .A1(n1280), .A2(n1281), .A3(KEYINPUT56), .ZN(n1275) );
NAND2_X1 U963 ( .A1(n1193), .A2(n1197), .ZN(n1281) );
NAND2_X1 U964 ( .A1(n1282), .A2(n1187), .ZN(n1280) );
XNOR2_X1 U965 ( .A(KEYINPUT30), .B(n1193), .ZN(n1282) );
INV_X1 U966 ( .A(n1186), .ZN(n1193) );
XNOR2_X1 U967 ( .A(n1283), .B(n1284), .ZN(n1186) );
XNOR2_X1 U968 ( .A(n1285), .B(n1121), .ZN(n1284) );
XNOR2_X1 U969 ( .A(G113), .B(n1286), .ZN(n1283) );
NOR2_X1 U970 ( .A1(G119), .A2(KEYINPUT12), .ZN(n1286) );
XOR2_X1 U971 ( .A(n1287), .B(n1158), .Z(n1265) );
NAND2_X1 U972 ( .A1(G217), .A2(n1288), .ZN(n1158) );
XNOR2_X1 U973 ( .A(n1107), .B(KEYINPUT24), .ZN(n1287) );
AND2_X1 U974 ( .A1(n1289), .A2(n1192), .ZN(n1107) );
XOR2_X1 U975 ( .A(n1156), .B(KEYINPUT8), .Z(n1289) );
XNOR2_X1 U976 ( .A(n1290), .B(n1291), .ZN(n1156) );
XOR2_X1 U977 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U978 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U979 ( .A(n1296), .B(n1297), .Z(n1295) );
AND3_X1 U980 ( .A1(G221), .A2(n1048), .A3(G234), .ZN(n1297) );
NOR2_X1 U981 ( .A1(KEYINPUT18), .A2(G146), .ZN(n1296) );
XNOR2_X1 U982 ( .A(G119), .B(n1203), .ZN(n1294) );
XOR2_X1 U983 ( .A(n1298), .B(n1299), .Z(n1292) );
XOR2_X1 U984 ( .A(G137), .B(G128), .Z(n1299) );
XOR2_X1 U985 ( .A(KEYINPUT58), .B(KEYINPUT21), .Z(n1298) );
NOR2_X1 U986 ( .A1(n1088), .A2(n1065), .ZN(n1241) );
NAND2_X1 U987 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U988 ( .A1(G221), .A2(n1288), .ZN(n1067) );
NAND2_X1 U989 ( .A1(G234), .A2(n1192), .ZN(n1288) );
XNOR2_X1 U990 ( .A(n1300), .B(G469), .ZN(n1066) );
NAND2_X1 U991 ( .A1(n1301), .A2(n1192), .ZN(n1300) );
XOR2_X1 U992 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U993 ( .A(n1198), .B(n1304), .ZN(n1303) );
NOR2_X1 U994 ( .A1(KEYINPUT10), .A2(n1202), .ZN(n1304) );
INV_X1 U995 ( .A(G140), .ZN(n1202) );
XNOR2_X1 U996 ( .A(n1305), .B(n1306), .ZN(n1198) );
XNOR2_X1 U997 ( .A(n1307), .B(n1308), .ZN(n1306) );
AND2_X1 U998 ( .A1(n1048), .A2(G227), .ZN(n1307) );
XNOR2_X1 U999 ( .A(n1309), .B(n1180), .ZN(n1305) );
INV_X1 U1000 ( .A(G101), .ZN(n1180) );
NAND2_X1 U1001 ( .A1(KEYINPUT19), .A2(n1310), .ZN(n1309) );
XNOR2_X1 U1002 ( .A(n1043), .B(n1311), .ZN(n1310) );
NOR2_X1 U1003 ( .A1(KEYINPUT0), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U1004 ( .A(G110), .B(n1313), .ZN(n1302) );
NOR2_X1 U1005 ( .A1(KEYINPUT34), .A2(n1197), .ZN(n1313) );
INV_X1 U1006 ( .A(n1187), .ZN(n1197) );
XOR2_X1 U1007 ( .A(G131), .B(n1131), .Z(n1187) );
XNOR2_X1 U1008 ( .A(n1130), .B(G137), .ZN(n1131) );
INV_X1 U1009 ( .A(n1221), .ZN(n1088) );
NOR2_X1 U1010 ( .A1(n1090), .A2(n1056), .ZN(n1221) );
AND2_X1 U1011 ( .A1(G214), .A2(n1314), .ZN(n1056) );
INV_X1 U1012 ( .A(n1054), .ZN(n1090) );
NAND3_X1 U1013 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n1054) );
NAND2_X1 U1014 ( .A1(n1318), .A2(n1109), .ZN(n1317) );
NAND2_X1 U1015 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
NAND2_X1 U1016 ( .A1(n1207), .A2(n1321), .ZN(n1320) );
NAND3_X1 U1017 ( .A1(n1322), .A2(n1111), .A3(n1319), .ZN(n1316) );
INV_X1 U1018 ( .A(KEYINPUT15), .ZN(n1319) );
NAND2_X1 U1019 ( .A1(n1321), .A2(n1109), .ZN(n1322) );
NAND2_X1 U1020 ( .A1(n1323), .A2(n1192), .ZN(n1109) );
XNOR2_X1 U1021 ( .A(n1206), .B(KEYINPUT36), .ZN(n1323) );
XNOR2_X1 U1022 ( .A(n1324), .B(n1325), .ZN(n1206) );
XNOR2_X1 U1023 ( .A(n1308), .B(n1144), .ZN(n1325) );
XOR2_X1 U1024 ( .A(G110), .B(n1326), .Z(n1144) );
XOR2_X1 U1025 ( .A(KEYINPUT41), .B(G122), .Z(n1326) );
INV_X1 U1026 ( .A(n1121), .ZN(n1308) );
XOR2_X1 U1027 ( .A(G128), .B(n1327), .Z(n1121) );
XOR2_X1 U1028 ( .A(n1328), .B(n1329), .Z(n1324) );
AND2_X1 U1029 ( .A1(n1048), .A2(G224), .ZN(n1329) );
XNOR2_X1 U1030 ( .A(n1330), .B(n1331), .ZN(n1328) );
INV_X1 U1031 ( .A(G125), .ZN(n1331) );
NAND2_X1 U1032 ( .A1(n1332), .A2(n1333), .ZN(n1330) );
NAND2_X1 U1033 ( .A1(n1334), .A2(n1145), .ZN(n1333) );
XOR2_X1 U1034 ( .A(n1335), .B(KEYINPUT61), .Z(n1332) );
OR2_X1 U1035 ( .A1(n1145), .A2(n1334), .ZN(n1335) );
XNOR2_X1 U1036 ( .A(n1143), .B(KEYINPUT50), .ZN(n1334) );
XNOR2_X1 U1037 ( .A(n1336), .B(n1337), .ZN(n1143) );
NAND3_X1 U1038 ( .A1(n1338), .A2(n1339), .A3(KEYINPUT62), .ZN(n1336) );
NAND2_X1 U1039 ( .A1(KEYINPUT4), .A2(n1340), .ZN(n1339) );
XNOR2_X1 U1040 ( .A(G119), .B(n1341), .ZN(n1340) );
NAND3_X1 U1041 ( .A1(G119), .A2(n1285), .A3(n1342), .ZN(n1338) );
INV_X1 U1042 ( .A(KEYINPUT4), .ZN(n1342) );
XOR2_X1 U1043 ( .A(G101), .B(n1343), .Z(n1145) );
NOR2_X1 U1044 ( .A1(KEYINPUT11), .A2(n1344), .ZN(n1343) );
XNOR2_X1 U1045 ( .A(n1043), .B(n1312), .ZN(n1344) );
XOR2_X1 U1046 ( .A(KEYINPUT52), .B(KEYINPUT42), .Z(n1321) );
NAND2_X1 U1047 ( .A1(KEYINPUT15), .A2(n1207), .ZN(n1315) );
INV_X1 U1048 ( .A(n1111), .ZN(n1207) );
NAND2_X1 U1049 ( .A1(G210), .A2(n1314), .ZN(n1111) );
NAND2_X1 U1050 ( .A1(n1279), .A2(n1192), .ZN(n1314) );
NOR2_X1 U1051 ( .A1(n1237), .A2(n1103), .ZN(n1249) );
XNOR2_X1 U1052 ( .A(n1345), .B(G475), .ZN(n1103) );
NAND2_X1 U1053 ( .A1(n1169), .A2(n1192), .ZN(n1345) );
XNOR2_X1 U1054 ( .A(n1346), .B(n1347), .ZN(n1169) );
XOR2_X1 U1055 ( .A(n1348), .B(n1349), .Z(n1347) );
XNOR2_X1 U1056 ( .A(n1337), .B(n1350), .ZN(n1349) );
AND3_X1 U1057 ( .A1(G214), .A2(n1048), .A3(n1279), .ZN(n1350) );
INV_X1 U1058 ( .A(G237), .ZN(n1279) );
INV_X1 U1059 ( .A(G113), .ZN(n1337) );
XOR2_X1 U1060 ( .A(G131), .B(G122), .Z(n1348) );
XOR2_X1 U1061 ( .A(n1351), .B(n1312), .Z(n1346) );
XOR2_X1 U1062 ( .A(G104), .B(KEYINPUT5), .Z(n1312) );
XNOR2_X1 U1063 ( .A(n1327), .B(n1290), .ZN(n1351) );
XNOR2_X1 U1064 ( .A(n1124), .B(KEYINPUT57), .ZN(n1290) );
XNOR2_X1 U1065 ( .A(G125), .B(G140), .ZN(n1124) );
XOR2_X1 U1066 ( .A(G143), .B(G146), .Z(n1327) );
INV_X1 U1067 ( .A(n1271), .ZN(n1237) );
NOR2_X1 U1068 ( .A1(n1106), .A2(n1352), .ZN(n1271) );
AND2_X1 U1069 ( .A1(G478), .A2(n1104), .ZN(n1352) );
NOR2_X1 U1070 ( .A1(n1104), .A2(G478), .ZN(n1106) );
NAND2_X1 U1071 ( .A1(n1192), .A2(n1166), .ZN(n1104) );
NAND3_X1 U1072 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1166) );
NAND2_X1 U1073 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
NAND2_X1 U1074 ( .A1(n1358), .A2(n1359), .ZN(n1354) );
INV_X1 U1075 ( .A(KEYINPUT1), .ZN(n1359) );
NAND2_X1 U1076 ( .A1(n1360), .A2(n1361), .ZN(n1358) );
XNOR2_X1 U1077 ( .A(n1356), .B(KEYINPUT53), .ZN(n1360) );
NAND2_X1 U1078 ( .A1(KEYINPUT1), .A2(n1362), .ZN(n1353) );
NAND2_X1 U1079 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
OR3_X1 U1080 ( .A1(n1357), .A2(n1356), .A3(KEYINPUT53), .ZN(n1364) );
INV_X1 U1081 ( .A(n1361), .ZN(n1357) );
XNOR2_X1 U1082 ( .A(n1365), .B(n1366), .ZN(n1361) );
XNOR2_X1 U1083 ( .A(G122), .B(n1043), .ZN(n1366) );
INV_X1 U1084 ( .A(G107), .ZN(n1043) );
XNOR2_X1 U1085 ( .A(n1367), .B(n1285), .ZN(n1365) );
INV_X1 U1086 ( .A(n1341), .ZN(n1285) );
XOR2_X1 U1087 ( .A(G116), .B(KEYINPUT44), .Z(n1341) );
NAND2_X1 U1088 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
NAND2_X1 U1089 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
XNOR2_X1 U1090 ( .A(n1372), .B(n1130), .ZN(n1370) );
INV_X1 U1091 ( .A(G134), .ZN(n1130) );
XNOR2_X1 U1092 ( .A(KEYINPUT45), .B(KEYINPUT22), .ZN(n1372) );
XOR2_X1 U1093 ( .A(KEYINPUT39), .B(n1373), .Z(n1368) );
NOR2_X1 U1094 ( .A1(G134), .A2(n1371), .ZN(n1373) );
XOR2_X1 U1095 ( .A(G143), .B(G128), .Z(n1371) );
NAND2_X1 U1096 ( .A1(KEYINPUT53), .A2(n1356), .ZN(n1363) );
AND3_X1 U1097 ( .A1(G217), .A2(n1048), .A3(G234), .ZN(n1356) );
NAND2_X1 U1098 ( .A1(n1258), .A2(n1374), .ZN(n1215) );
NAND2_X1 U1099 ( .A1(n1375), .A2(n1261), .ZN(n1374) );
INV_X1 U1100 ( .A(n1140), .ZN(n1375) );
NOR2_X1 U1101 ( .A1(n1048), .A2(G898), .ZN(n1140) );
AND2_X1 U1102 ( .A1(n1091), .A2(n1376), .ZN(n1258) );
NAND2_X1 U1103 ( .A1(n1261), .A2(n1192), .ZN(n1376) );
INV_X1 U1104 ( .A(G902), .ZN(n1192) );
NAND2_X1 U1105 ( .A1(G952), .A2(n1377), .ZN(n1261) );
XNOR2_X1 U1106 ( .A(KEYINPUT35), .B(n1048), .ZN(n1377) );
INV_X1 U1107 ( .A(G953), .ZN(n1048) );
NAND2_X1 U1108 ( .A1(G237), .A2(G234), .ZN(n1091) );
INV_X1 U1109 ( .A(G110), .ZN(n1203) );
endmodule


