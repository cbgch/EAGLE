//Key = 0110000001001111100010001000111011110000010111010100000111100101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340;

XNOR2_X1 U733 ( .A(G107), .B(n1016), .ZN(G9) );
NOR2_X1 U734 ( .A1(n1017), .A2(n1018), .ZN(G75) );
NOR3_X1 U735 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NAND3_X1 U736 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1019) );
NAND2_X1 U737 ( .A1(n1025), .A2(n1026), .ZN(n1022) );
NAND2_X1 U738 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND3_X1 U739 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NAND3_X1 U740 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1030) );
NAND2_X1 U741 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND3_X1 U742 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1033) );
XNOR2_X1 U743 ( .A(n1036), .B(KEYINPUT41), .ZN(n1039) );
NAND2_X1 U744 ( .A1(n1040), .A2(n1041), .ZN(n1032) );
NAND2_X1 U745 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U746 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND4_X1 U747 ( .A1(n1036), .A2(n1040), .A3(n1046), .A4(n1047), .ZN(n1027) );
NAND2_X1 U748 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U749 ( .A1(n1029), .A2(n1050), .ZN(n1048) );
NAND2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
OR3_X1 U751 ( .A1(n1053), .A2(n1054), .A3(n1049), .ZN(n1046) );
INV_X1 U752 ( .A(n1031), .ZN(n1049) );
INV_X1 U753 ( .A(n1055), .ZN(n1025) );
AND3_X1 U754 ( .A1(n1024), .A2(n1056), .A3(n1023), .ZN(n1017) );
NAND4_X1 U755 ( .A1(n1057), .A2(n1036), .A3(n1058), .A4(n1059), .ZN(n1023) );
NOR4_X1 U756 ( .A1(n1051), .A2(n1060), .A3(n1061), .A4(n1038), .ZN(n1059) );
XOR2_X1 U757 ( .A(n1062), .B(n1063), .Z(n1061) );
XOR2_X1 U758 ( .A(KEYINPUT48), .B(G469), .Z(n1063) );
NAND2_X1 U759 ( .A1(KEYINPUT12), .A2(n1064), .ZN(n1062) );
NOR2_X1 U760 ( .A1(n1065), .A2(n1066), .ZN(n1060) );
NOR2_X1 U761 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U762 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
INV_X1 U763 ( .A(KEYINPUT33), .ZN(n1070) );
NOR2_X1 U764 ( .A1(KEYINPUT53), .A2(n1071), .ZN(n1069) );
NOR2_X1 U765 ( .A1(G472), .A2(n1072), .ZN(n1065) );
NOR2_X1 U766 ( .A1(n1073), .A2(KEYINPUT53), .ZN(n1072) );
AND2_X1 U767 ( .A1(n1068), .A2(KEYINPUT33), .ZN(n1073) );
XOR2_X1 U768 ( .A(n1074), .B(KEYINPUT32), .Z(n1058) );
NAND2_X1 U769 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U770 ( .A1(G478), .A2(n1077), .ZN(n1076) );
XNOR2_X1 U771 ( .A(n1078), .B(KEYINPUT54), .ZN(n1057) );
XOR2_X1 U772 ( .A(n1079), .B(n1080), .Z(G72) );
XOR2_X1 U773 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND3_X1 U774 ( .A1(n1020), .A2(n1083), .A3(KEYINPUT15), .ZN(n1082) );
NAND2_X1 U775 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
NAND2_X1 U776 ( .A1(G953), .A2(n1086), .ZN(n1085) );
XOR2_X1 U777 ( .A(n1087), .B(n1088), .Z(n1084) );
XNOR2_X1 U778 ( .A(n1089), .B(n1090), .ZN(n1088) );
XOR2_X1 U779 ( .A(KEYINPUT60), .B(KEYINPUT23), .Z(n1090) );
XNOR2_X1 U780 ( .A(n1091), .B(n1092), .ZN(n1087) );
NOR2_X1 U781 ( .A1(KEYINPUT6), .A2(n1093), .ZN(n1092) );
XOR2_X1 U782 ( .A(KEYINPUT34), .B(n1094), .Z(n1093) );
NOR3_X1 U783 ( .A1(n1083), .A2(KEYINPUT21), .A3(n1095), .ZN(n1079) );
NOR2_X1 U784 ( .A1(n1096), .A2(n1086), .ZN(n1095) );
XOR2_X1 U785 ( .A(n1097), .B(n1098), .Z(G69) );
NOR2_X1 U786 ( .A1(n1099), .A2(n1083), .ZN(n1098) );
NOR2_X1 U787 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U788 ( .A1(n1102), .A2(n1103), .ZN(n1097) );
NAND2_X1 U789 ( .A1(n1104), .A2(n1083), .ZN(n1103) );
XOR2_X1 U790 ( .A(n1105), .B(n1021), .Z(n1104) );
NAND3_X1 U791 ( .A1(n1105), .A2(G898), .A3(G953), .ZN(n1102) );
NOR2_X1 U792 ( .A1(KEYINPUT38), .A2(n1106), .ZN(n1105) );
NOR3_X1 U793 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(G66) );
AND3_X1 U794 ( .A1(KEYINPUT62), .A2(G953), .A3(G952), .ZN(n1109) );
NOR2_X1 U795 ( .A1(KEYINPUT62), .A2(n1110), .ZN(n1108) );
INV_X1 U796 ( .A(n1111), .ZN(n1110) );
XNOR2_X1 U797 ( .A(n1112), .B(n1113), .ZN(n1107) );
NOR2_X1 U798 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR3_X1 U799 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(G63) );
AND2_X1 U800 ( .A1(n1111), .A2(KEYINPUT45), .ZN(n1118) );
NOR3_X1 U801 ( .A1(KEYINPUT45), .A2(n1083), .A3(n1056), .ZN(n1117) );
INV_X1 U802 ( .A(G952), .ZN(n1056) );
NOR2_X1 U803 ( .A1(n1119), .A2(n1120), .ZN(n1116) );
XOR2_X1 U804 ( .A(n1121), .B(KEYINPUT43), .Z(n1120) );
NAND2_X1 U805 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XOR2_X1 U806 ( .A(KEYINPUT17), .B(n1124), .Z(n1123) );
NOR2_X1 U807 ( .A1(n1122), .A2(n1124), .ZN(n1119) );
INV_X1 U808 ( .A(n1125), .ZN(n1124) );
AND2_X1 U809 ( .A1(n1126), .A2(G478), .ZN(n1122) );
NOR2_X1 U810 ( .A1(n1111), .A2(n1127), .ZN(G60) );
XNOR2_X1 U811 ( .A(n1128), .B(n1129), .ZN(n1127) );
NOR3_X1 U812 ( .A1(n1115), .A2(KEYINPUT59), .A3(n1130), .ZN(n1128) );
XNOR2_X1 U813 ( .A(G104), .B(n1131), .ZN(G6) );
NAND4_X1 U814 ( .A1(n1132), .A2(n1053), .A3(n1040), .A4(n1133), .ZN(n1131) );
XOR2_X1 U815 ( .A(n1134), .B(KEYINPUT8), .Z(n1132) );
NOR2_X1 U816 ( .A1(n1111), .A2(n1135), .ZN(G57) );
XOR2_X1 U817 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U818 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U819 ( .A1(n1071), .A2(n1115), .ZN(n1139) );
NOR3_X1 U820 ( .A1(KEYINPUT37), .A2(n1140), .A3(n1141), .ZN(n1138) );
NOR2_X1 U821 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NOR2_X1 U822 ( .A1(n1144), .A2(n1145), .ZN(n1140) );
INV_X1 U823 ( .A(n1143), .ZN(n1145) );
XOR2_X1 U824 ( .A(KEYINPUT14), .B(n1142), .Z(n1144) );
NOR2_X1 U825 ( .A1(n1111), .A2(n1146), .ZN(G54) );
NOR2_X1 U826 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U827 ( .A(KEYINPUT26), .B(n1149), .Z(n1148) );
NOR2_X1 U828 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
AND2_X1 U829 ( .A1(n1151), .A2(n1150), .ZN(n1147) );
XOR2_X1 U830 ( .A(n1152), .B(n1153), .Z(n1150) );
XOR2_X1 U831 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U832 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
INV_X1 U833 ( .A(n1158), .ZN(n1157) );
NOR2_X1 U834 ( .A1(n1159), .A2(n1089), .ZN(n1156) );
NOR2_X1 U835 ( .A1(KEYINPUT22), .A2(n1160), .ZN(n1154) );
XOR2_X1 U836 ( .A(n1161), .B(n1162), .Z(n1152) );
NOR2_X1 U837 ( .A1(KEYINPUT36), .A2(n1163), .ZN(n1162) );
NAND2_X1 U838 ( .A1(n1126), .A2(G469), .ZN(n1151) );
NOR2_X1 U839 ( .A1(n1111), .A2(n1164), .ZN(G51) );
XOR2_X1 U840 ( .A(n1165), .B(n1166), .Z(n1164) );
XNOR2_X1 U841 ( .A(n1167), .B(n1106), .ZN(n1166) );
NAND2_X1 U842 ( .A1(n1126), .A2(n1168), .ZN(n1167) );
INV_X1 U843 ( .A(n1115), .ZN(n1126) );
NAND2_X1 U844 ( .A1(n1169), .A2(n1170), .ZN(n1115) );
OR2_X1 U845 ( .A1(n1021), .A2(n1020), .ZN(n1170) );
NAND4_X1 U846 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1020) );
AND4_X1 U847 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1174) );
OR2_X1 U848 ( .A1(n1179), .A2(n1180), .ZN(n1173) );
NAND4_X1 U849 ( .A1(n1037), .A2(n1038), .A3(n1181), .A4(n1182), .ZN(n1171) );
NAND2_X1 U850 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
INV_X1 U851 ( .A(n1053), .ZN(n1184) );
NAND2_X1 U852 ( .A1(KEYINPUT25), .A2(n1185), .ZN(n1183) );
NAND3_X1 U853 ( .A1(n1186), .A2(n1187), .A3(n1053), .ZN(n1181) );
NAND3_X1 U854 ( .A1(n1188), .A2(n1189), .A3(n1031), .ZN(n1187) );
OR2_X1 U855 ( .A1(n1190), .A2(KEYINPUT25), .ZN(n1186) );
NAND4_X1 U856 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1021) );
AND4_X1 U857 ( .A1(n1016), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1194) );
NAND3_X1 U858 ( .A1(n1040), .A2(n1198), .A3(n1054), .ZN(n1016) );
NOR2_X1 U859 ( .A1(n1199), .A2(n1200), .ZN(n1193) );
AND3_X1 U860 ( .A1(n1053), .A2(n1198), .A3(n1040), .ZN(n1200) );
INV_X1 U861 ( .A(n1201), .ZN(n1199) );
XNOR2_X1 U862 ( .A(KEYINPUT4), .B(n1202), .ZN(n1169) );
XOR2_X1 U863 ( .A(n1203), .B(n1204), .Z(n1165) );
NOR2_X1 U864 ( .A1(KEYINPUT52), .A2(n1091), .ZN(n1204) );
NOR2_X1 U865 ( .A1(n1083), .A2(G952), .ZN(n1111) );
XNOR2_X1 U866 ( .A(G146), .B(n1172), .ZN(G48) );
NAND2_X1 U867 ( .A1(n1205), .A2(n1053), .ZN(n1172) );
XNOR2_X1 U868 ( .A(G143), .B(n1178), .ZN(G45) );
NAND3_X1 U869 ( .A1(n1035), .A2(n1133), .A3(n1206), .ZN(n1178) );
NOR3_X1 U870 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1206) );
XNOR2_X1 U871 ( .A(n1089), .B(n1210), .ZN(G42) );
NOR2_X1 U872 ( .A1(n1190), .A2(n1211), .ZN(n1210) );
XNOR2_X1 U873 ( .A(G137), .B(n1177), .ZN(G39) );
NAND3_X1 U874 ( .A1(n1212), .A2(n1213), .A3(n1185), .ZN(n1177) );
XNOR2_X1 U875 ( .A(G134), .B(n1176), .ZN(G36) );
NAND3_X1 U876 ( .A1(n1035), .A2(n1054), .A3(n1185), .ZN(n1176) );
INV_X1 U877 ( .A(n1190), .ZN(n1185) );
NAND2_X1 U878 ( .A1(n1214), .A2(n1036), .ZN(n1190) );
INV_X1 U879 ( .A(n1180), .ZN(n1036) );
XNOR2_X1 U880 ( .A(n1215), .B(n1216), .ZN(G33) );
NOR2_X1 U881 ( .A1(n1217), .A2(n1180), .ZN(n1216) );
NAND2_X1 U882 ( .A1(n1045), .A2(n1218), .ZN(n1180) );
XOR2_X1 U883 ( .A(n1179), .B(KEYINPUT46), .Z(n1217) );
NAND3_X1 U884 ( .A1(n1035), .A2(n1053), .A3(n1214), .ZN(n1179) );
NOR3_X1 U885 ( .A1(n1209), .A2(n1051), .A3(n1219), .ZN(n1214) );
INV_X1 U886 ( .A(n1189), .ZN(n1209) );
XNOR2_X1 U887 ( .A(G128), .B(n1175), .ZN(G30) );
NAND2_X1 U888 ( .A1(n1205), .A2(n1054), .ZN(n1175) );
AND4_X1 U889 ( .A1(n1133), .A2(n1038), .A3(n1213), .A4(n1189), .ZN(n1205) );
XOR2_X1 U890 ( .A(n1220), .B(G101), .Z(G3) );
NAND2_X1 U891 ( .A1(KEYINPUT16), .A2(n1201), .ZN(n1220) );
NAND3_X1 U892 ( .A1(n1029), .A2(n1198), .A3(n1035), .ZN(n1201) );
XOR2_X1 U893 ( .A(n1221), .B(n1222), .Z(G27) );
XNOR2_X1 U894 ( .A(G125), .B(KEYINPUT40), .ZN(n1222) );
NAND4_X1 U895 ( .A1(n1223), .A2(n1224), .A3(n1031), .A4(n1189), .ZN(n1221) );
NAND2_X1 U896 ( .A1(n1055), .A2(n1225), .ZN(n1189) );
NAND4_X1 U897 ( .A1(G953), .A2(G902), .A3(n1226), .A4(n1086), .ZN(n1225) );
INV_X1 U898 ( .A(G900), .ZN(n1086) );
INV_X1 U899 ( .A(n1211), .ZN(n1224) );
NAND3_X1 U900 ( .A1(n1037), .A2(n1038), .A3(n1053), .ZN(n1211) );
XNOR2_X1 U901 ( .A(n1188), .B(KEYINPUT61), .ZN(n1223) );
XNOR2_X1 U902 ( .A(G122), .B(n1191), .ZN(G24) );
NAND4_X1 U903 ( .A1(n1227), .A2(n1040), .A3(n1078), .A4(n1228), .ZN(n1191) );
NOR2_X1 U904 ( .A1(n1213), .A2(n1038), .ZN(n1040) );
XNOR2_X1 U905 ( .A(G119), .B(n1192), .ZN(G21) );
NAND3_X1 U906 ( .A1(n1212), .A2(n1213), .A3(n1227), .ZN(n1192) );
XOR2_X1 U907 ( .A(n1197), .B(n1229), .Z(G18) );
XOR2_X1 U908 ( .A(KEYINPUT49), .B(G116), .Z(n1229) );
NAND3_X1 U909 ( .A1(n1227), .A2(n1054), .A3(n1035), .ZN(n1197) );
NOR2_X1 U910 ( .A1(n1078), .A2(n1208), .ZN(n1054) );
INV_X1 U911 ( .A(n1228), .ZN(n1208) );
XOR2_X1 U912 ( .A(n1196), .B(n1230), .Z(G15) );
XOR2_X1 U913 ( .A(KEYINPUT20), .B(G113), .Z(n1230) );
NAND3_X1 U914 ( .A1(n1227), .A2(n1053), .A3(n1035), .ZN(n1196) );
NOR2_X1 U915 ( .A1(n1038), .A2(n1037), .ZN(n1035) );
NOR2_X1 U916 ( .A1(n1228), .A2(n1207), .ZN(n1053) );
INV_X1 U917 ( .A(n1078), .ZN(n1207) );
AND3_X1 U918 ( .A1(n1188), .A2(n1134), .A3(n1031), .ZN(n1227) );
NOR2_X1 U919 ( .A1(n1052), .A2(n1051), .ZN(n1031) );
INV_X1 U920 ( .A(n1219), .ZN(n1052) );
XNOR2_X1 U921 ( .A(G110), .B(n1195), .ZN(G12) );
NAND3_X1 U922 ( .A1(n1037), .A2(n1198), .A3(n1212), .ZN(n1195) );
AND2_X1 U923 ( .A1(n1029), .A2(n1038), .ZN(n1212) );
XOR2_X1 U924 ( .A(n1231), .B(n1114), .Z(n1038) );
NAND2_X1 U925 ( .A1(G217), .A2(n1232), .ZN(n1114) );
NAND2_X1 U926 ( .A1(n1233), .A2(n1112), .ZN(n1231) );
NAND3_X1 U927 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1112) );
NAND2_X1 U928 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NAND2_X1 U929 ( .A1(n1239), .A2(n1240), .ZN(n1237) );
INV_X1 U930 ( .A(KEYINPUT50), .ZN(n1240) );
XOR2_X1 U931 ( .A(n1241), .B(KEYINPUT30), .Z(n1239) );
OR3_X1 U932 ( .A1(n1241), .A2(n1238), .A3(KEYINPUT50), .ZN(n1235) );
NAND2_X1 U933 ( .A1(n1242), .A2(n1243), .ZN(n1238) );
NAND2_X1 U934 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XOR2_X1 U935 ( .A(KEYINPUT28), .B(n1246), .Z(n1242) );
NOR2_X1 U936 ( .A1(n1245), .A2(n1244), .ZN(n1246) );
XNOR2_X1 U937 ( .A(n1247), .B(n1248), .ZN(n1244) );
XNOR2_X1 U938 ( .A(n1249), .B(n1250), .ZN(n1248) );
NOR2_X1 U939 ( .A1(G110), .A2(KEYINPUT7), .ZN(n1250) );
NAND2_X1 U940 ( .A1(KEYINPUT56), .A2(G128), .ZN(n1249) );
XNOR2_X1 U941 ( .A(G119), .B(KEYINPUT42), .ZN(n1247) );
NAND2_X1 U942 ( .A1(KEYINPUT50), .A2(n1241), .ZN(n1234) );
NAND2_X1 U943 ( .A1(n1251), .A2(n1252), .ZN(n1241) );
NAND3_X1 U944 ( .A1(n1253), .A2(n1254), .A3(G221), .ZN(n1252) );
NAND2_X1 U945 ( .A1(n1255), .A2(n1256), .ZN(n1251) );
NAND2_X1 U946 ( .A1(G221), .A2(n1253), .ZN(n1256) );
XOR2_X1 U947 ( .A(KEYINPUT35), .B(n1254), .Z(n1255) );
XNOR2_X1 U948 ( .A(n1257), .B(KEYINPUT3), .ZN(n1254) );
INV_X1 U949 ( .A(G137), .ZN(n1257) );
NOR2_X1 U950 ( .A1(n1228), .A2(n1078), .ZN(n1029) );
XOR2_X1 U951 ( .A(n1258), .B(n1130), .Z(n1078) );
INV_X1 U952 ( .A(G475), .ZN(n1130) );
NAND2_X1 U953 ( .A1(n1129), .A2(n1233), .ZN(n1258) );
XOR2_X1 U954 ( .A(n1259), .B(n1260), .Z(n1129) );
XOR2_X1 U955 ( .A(n1261), .B(n1262), .Z(n1260) );
XOR2_X1 U956 ( .A(n1263), .B(n1264), .Z(n1262) );
NOR2_X1 U957 ( .A1(KEYINPUT51), .A2(n1265), .ZN(n1264) );
NAND2_X1 U958 ( .A1(G214), .A2(n1266), .ZN(n1263) );
NAND2_X1 U959 ( .A1(KEYINPUT29), .A2(n1267), .ZN(n1261) );
INV_X1 U960 ( .A(n1245), .ZN(n1267) );
XOR2_X1 U961 ( .A(G125), .B(n1268), .Z(n1245) );
XNOR2_X1 U962 ( .A(G146), .B(n1089), .ZN(n1268) );
XOR2_X1 U963 ( .A(n1269), .B(n1270), .Z(n1259) );
XNOR2_X1 U964 ( .A(G143), .B(n1215), .ZN(n1270) );
XNOR2_X1 U965 ( .A(G113), .B(G104), .ZN(n1269) );
NAND3_X1 U966 ( .A1(n1271), .A2(n1272), .A3(n1075), .ZN(n1228) );
OR2_X1 U967 ( .A1(n1077), .A2(G478), .ZN(n1075) );
OR2_X1 U968 ( .A1(G478), .A2(KEYINPUT63), .ZN(n1272) );
NAND3_X1 U969 ( .A1(G478), .A2(n1077), .A3(KEYINPUT63), .ZN(n1271) );
NAND2_X1 U970 ( .A1(n1125), .A2(n1233), .ZN(n1077) );
XOR2_X1 U971 ( .A(n1273), .B(n1274), .Z(n1125) );
XNOR2_X1 U972 ( .A(n1275), .B(n1276), .ZN(n1274) );
NAND2_X1 U973 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
NAND2_X1 U974 ( .A1(G122), .A2(n1279), .ZN(n1278) );
XOR2_X1 U975 ( .A(n1280), .B(KEYINPUT10), .Z(n1277) );
NAND2_X1 U976 ( .A1(n1281), .A2(n1265), .ZN(n1280) );
XOR2_X1 U977 ( .A(n1282), .B(n1283), .Z(n1273) );
XOR2_X1 U978 ( .A(G134), .B(G107), .Z(n1283) );
NAND2_X1 U979 ( .A1(G217), .A2(n1253), .ZN(n1282) );
AND2_X1 U980 ( .A1(G234), .A2(n1083), .ZN(n1253) );
INV_X1 U981 ( .A(G953), .ZN(n1083) );
AND2_X1 U982 ( .A1(n1133), .A2(n1134), .ZN(n1198) );
NAND2_X1 U983 ( .A1(n1055), .A2(n1284), .ZN(n1134) );
NAND4_X1 U984 ( .A1(G953), .A2(G902), .A3(n1226), .A4(n1101), .ZN(n1284) );
INV_X1 U985 ( .A(G898), .ZN(n1101) );
NAND3_X1 U986 ( .A1(n1024), .A2(n1226), .A3(G952), .ZN(n1055) );
NAND2_X1 U987 ( .A1(G237), .A2(G234), .ZN(n1226) );
XOR2_X1 U988 ( .A(G953), .B(KEYINPUT47), .Z(n1024) );
NOR3_X1 U989 ( .A1(n1219), .A2(n1051), .A3(n1042), .ZN(n1133) );
INV_X1 U990 ( .A(n1188), .ZN(n1042) );
NOR2_X1 U991 ( .A1(n1045), .A2(n1044), .ZN(n1188) );
INV_X1 U992 ( .A(n1218), .ZN(n1044) );
NAND2_X1 U993 ( .A1(G214), .A2(n1285), .ZN(n1218) );
XOR2_X1 U994 ( .A(n1286), .B(n1168), .Z(n1045) );
AND2_X1 U995 ( .A1(G210), .A2(n1285), .ZN(n1168) );
NAND2_X1 U996 ( .A1(n1287), .A2(n1202), .ZN(n1285) );
INV_X1 U997 ( .A(G237), .ZN(n1287) );
NAND2_X1 U998 ( .A1(n1233), .A2(n1288), .ZN(n1286) );
XNOR2_X1 U999 ( .A(n1106), .B(n1289), .ZN(n1288) );
XOR2_X1 U1000 ( .A(n1290), .B(KEYINPUT27), .Z(n1289) );
NAND2_X1 U1001 ( .A1(KEYINPUT44), .A2(n1291), .ZN(n1290) );
XOR2_X1 U1002 ( .A(n1203), .B(n1091), .Z(n1291) );
XNOR2_X1 U1003 ( .A(n1292), .B(n1293), .ZN(n1091) );
INV_X1 U1004 ( .A(G125), .ZN(n1293) );
NOR2_X1 U1005 ( .A1(n1100), .A2(G953), .ZN(n1203) );
INV_X1 U1006 ( .A(G224), .ZN(n1100) );
XNOR2_X1 U1007 ( .A(n1294), .B(n1295), .ZN(n1106) );
XOR2_X1 U1008 ( .A(G101), .B(n1296), .Z(n1295) );
XNOR2_X1 U1009 ( .A(n1265), .B(G110), .ZN(n1296) );
INV_X1 U1010 ( .A(G122), .ZN(n1265) );
XOR2_X1 U1011 ( .A(n1297), .B(n1298), .Z(n1294) );
NOR2_X1 U1012 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
NOR2_X1 U1013 ( .A1(G107), .A2(n1301), .ZN(n1300) );
XNOR2_X1 U1014 ( .A(G104), .B(KEYINPUT58), .ZN(n1301) );
NAND2_X1 U1015 ( .A1(n1302), .A2(n1303), .ZN(n1297) );
OR2_X1 U1016 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
XOR2_X1 U1017 ( .A(n1306), .B(KEYINPUT18), .Z(n1302) );
NAND2_X1 U1018 ( .A1(n1304), .A2(n1305), .ZN(n1306) );
XNOR2_X1 U1019 ( .A(n1307), .B(KEYINPUT0), .ZN(n1304) );
AND2_X1 U1020 ( .A1(G221), .A2(n1232), .ZN(n1051) );
NAND2_X1 U1021 ( .A1(G234), .A2(n1202), .ZN(n1232) );
INV_X1 U1022 ( .A(G902), .ZN(n1202) );
XOR2_X1 U1023 ( .A(G469), .B(n1308), .Z(n1219) );
NOR2_X1 U1024 ( .A1(n1309), .A2(KEYINPUT11), .ZN(n1308) );
INV_X1 U1025 ( .A(n1064), .ZN(n1309) );
NAND2_X1 U1026 ( .A1(n1233), .A2(n1310), .ZN(n1064) );
XOR2_X1 U1027 ( .A(n1311), .B(n1312), .Z(n1310) );
XOR2_X1 U1028 ( .A(n1161), .B(n1160), .Z(n1312) );
XNOR2_X1 U1029 ( .A(n1143), .B(KEYINPUT55), .ZN(n1160) );
XOR2_X1 U1030 ( .A(n1313), .B(n1314), .Z(n1161) );
XOR2_X1 U1031 ( .A(G101), .B(n1315), .Z(n1314) );
XOR2_X1 U1032 ( .A(KEYINPUT60), .B(KEYINPUT1), .Z(n1315) );
XNOR2_X1 U1033 ( .A(n1292), .B(n1316), .ZN(n1313) );
NOR2_X1 U1034 ( .A1(n1317), .A2(n1299), .ZN(n1316) );
AND2_X1 U1035 ( .A1(G104), .A2(G107), .ZN(n1299) );
NOR2_X1 U1036 ( .A1(G107), .A2(G104), .ZN(n1317) );
NAND2_X1 U1037 ( .A1(n1318), .A2(n1319), .ZN(n1311) );
NAND2_X1 U1038 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
INV_X1 U1039 ( .A(n1322), .ZN(n1321) );
NAND2_X1 U1040 ( .A1(n1158), .A2(n1323), .ZN(n1320) );
NAND2_X1 U1041 ( .A1(G140), .A2(n1324), .ZN(n1323) );
NAND2_X1 U1042 ( .A1(n1159), .A2(n1089), .ZN(n1158) );
NAND2_X1 U1043 ( .A1(n1322), .A2(n1325), .ZN(n1318) );
NAND2_X1 U1044 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
NAND2_X1 U1045 ( .A1(n1324), .A2(n1089), .ZN(n1327) );
INV_X1 U1046 ( .A(G140), .ZN(n1089) );
XOR2_X1 U1047 ( .A(n1159), .B(KEYINPUT24), .Z(n1324) );
NAND2_X1 U1048 ( .A1(n1159), .A2(G140), .ZN(n1326) );
NOR2_X1 U1049 ( .A1(n1096), .A2(G953), .ZN(n1159) );
INV_X1 U1050 ( .A(G227), .ZN(n1096) );
NOR2_X1 U1051 ( .A1(KEYINPUT19), .A2(n1163), .ZN(n1322) );
INV_X1 U1052 ( .A(G110), .ZN(n1163) );
INV_X1 U1053 ( .A(n1213), .ZN(n1037) );
XOR2_X1 U1054 ( .A(n1068), .B(n1071), .Z(n1213) );
INV_X1 U1055 ( .A(G472), .ZN(n1071) );
NAND2_X1 U1056 ( .A1(n1233), .A2(n1328), .ZN(n1068) );
XNOR2_X1 U1057 ( .A(n1329), .B(n1136), .ZN(n1328) );
XNOR2_X1 U1058 ( .A(n1330), .B(G101), .ZN(n1136) );
NAND2_X1 U1059 ( .A1(G210), .A2(n1266), .ZN(n1330) );
NOR2_X1 U1060 ( .A1(G953), .A2(G237), .ZN(n1266) );
NAND2_X1 U1061 ( .A1(n1331), .A2(KEYINPUT2), .ZN(n1329) );
XNOR2_X1 U1062 ( .A(n1143), .B(n1142), .ZN(n1331) );
XNOR2_X1 U1063 ( .A(n1332), .B(n1305), .ZN(n1142) );
XNOR2_X1 U1064 ( .A(G119), .B(n1281), .ZN(n1305) );
INV_X1 U1065 ( .A(n1279), .ZN(n1281) );
XOR2_X1 U1066 ( .A(G116), .B(KEYINPUT13), .Z(n1279) );
XOR2_X1 U1067 ( .A(n1333), .B(n1292), .Z(n1332) );
XOR2_X1 U1068 ( .A(G146), .B(n1276), .Z(n1292) );
XOR2_X1 U1069 ( .A(G128), .B(G143), .Z(n1276) );
NAND2_X1 U1070 ( .A1(n1334), .A2(KEYINPUT57), .ZN(n1333) );
XOR2_X1 U1071 ( .A(n1307), .B(KEYINPUT31), .Z(n1334) );
XNOR2_X1 U1072 ( .A(G113), .B(KEYINPUT9), .ZN(n1307) );
NAND2_X1 U1073 ( .A1(n1335), .A2(n1336), .ZN(n1143) );
NAND2_X1 U1074 ( .A1(n1094), .A2(n1337), .ZN(n1336) );
INV_X1 U1075 ( .A(KEYINPUT5), .ZN(n1337) );
NOR2_X1 U1076 ( .A1(n1338), .A2(n1339), .ZN(n1094) );
AND2_X1 U1077 ( .A1(n1340), .A2(n1215), .ZN(n1338) );
NAND2_X1 U1078 ( .A1(n1339), .A2(KEYINPUT5), .ZN(n1335) );
NOR2_X1 U1079 ( .A1(n1215), .A2(n1340), .ZN(n1339) );
XNOR2_X1 U1080 ( .A(G134), .B(G137), .ZN(n1340) );
INV_X1 U1081 ( .A(G131), .ZN(n1215) );
XNOR2_X1 U1082 ( .A(G902), .B(KEYINPUT39), .ZN(n1233) );
endmodule


