//Key = 0011111001111101010101010110110010110110001010110011110111111111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304;

XNOR2_X1 U724 ( .A(G107), .B(n996), .ZN(G9) );
NOR2_X1 U725 ( .A1(n997), .A2(n998), .ZN(G75) );
NOR4_X1 U726 ( .A1(n999), .A2(n1000), .A3(n1001), .A4(n1002), .ZN(n998) );
NOR4_X1 U727 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1001) );
NOR3_X1 U728 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1004) );
NOR2_X1 U729 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NOR3_X1 U730 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1010) );
AND2_X1 U731 ( .A1(n1015), .A2(KEYINPUT45), .ZN(n1012) );
NOR2_X1 U732 ( .A1(n1016), .A2(n1017), .ZN(n1008) );
NOR2_X1 U733 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
AND2_X1 U734 ( .A1(n1020), .A2(KEYINPUT63), .ZN(n1019) );
NOR3_X1 U735 ( .A1(n1021), .A2(KEYINPUT45), .A3(n1022), .ZN(n1018) );
NOR2_X1 U736 ( .A1(n1023), .A2(n1024), .ZN(n1003) );
NOR3_X1 U737 ( .A1(n1017), .A2(KEYINPUT63), .A3(n1025), .ZN(n1024) );
NAND3_X1 U738 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n999) );
NAND4_X1 U739 ( .A1(n1023), .A2(n1029), .A3(n1015), .A4(n1030), .ZN(n1028) );
NAND2_X1 U740 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U741 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U742 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U743 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U744 ( .A1(n1039), .A2(n1040), .ZN(n1031) );
NAND2_X1 U745 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U746 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
INV_X1 U747 ( .A(n1007), .ZN(n1023) );
AND3_X1 U748 ( .A1(n1026), .A2(n1027), .A3(n1045), .ZN(n997) );
NAND4_X1 U749 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1026) );
NOR3_X1 U750 ( .A1(n1044), .A2(n1050), .A3(n1051), .ZN(n1049) );
XNOR2_X1 U751 ( .A(n1052), .B(KEYINPUT34), .ZN(n1051) );
INV_X1 U752 ( .A(n1053), .ZN(n1050) );
XOR2_X1 U753 ( .A(n1054), .B(KEYINPUT16), .Z(n1048) );
XOR2_X1 U754 ( .A(n1055), .B(KEYINPUT49), .Z(n1047) );
XOR2_X1 U755 ( .A(n1056), .B(KEYINPUT15), .Z(n1046) );
NAND4_X1 U756 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
NOR2_X1 U757 ( .A1(n1037), .A2(n1061), .ZN(n1059) );
NAND2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(n1058) );
XNOR2_X1 U759 ( .A(n1064), .B(n1065), .ZN(n1057) );
XOR2_X1 U760 ( .A(n1066), .B(n1067), .Z(G72) );
XOR2_X1 U761 ( .A(n1068), .B(n1069), .Z(n1067) );
NOR2_X1 U762 ( .A1(n1070), .A2(n1027), .ZN(n1069) );
AND2_X1 U763 ( .A1(G227), .A2(G900), .ZN(n1070) );
NAND3_X1 U764 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1068) );
XOR2_X1 U765 ( .A(KEYINPUT60), .B(n1074), .Z(n1073) );
NOR2_X1 U766 ( .A1(G900), .A2(n1027), .ZN(n1074) );
NAND2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(n1072) );
XOR2_X1 U768 ( .A(KEYINPUT38), .B(n1077), .Z(n1076) );
XNOR2_X1 U769 ( .A(n1078), .B(KEYINPUT44), .ZN(n1075) );
NAND2_X1 U770 ( .A1(n1079), .A2(n1077), .ZN(n1071) );
XNOR2_X1 U771 ( .A(KEYINPUT26), .B(n1080), .ZN(n1079) );
INV_X1 U772 ( .A(n1078), .ZN(n1080) );
XNOR2_X1 U773 ( .A(n1081), .B(n1082), .ZN(n1078) );
XNOR2_X1 U774 ( .A(KEYINPUT41), .B(n1083), .ZN(n1082) );
XOR2_X1 U775 ( .A(n1084), .B(n1085), .Z(n1081) );
NAND2_X1 U776 ( .A1(n1027), .A2(n1000), .ZN(n1066) );
XOR2_X1 U777 ( .A(n1086), .B(n1087), .Z(G69) );
XOR2_X1 U778 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U779 ( .A1(G953), .A2(n1090), .ZN(n1089) );
NAND2_X1 U780 ( .A1(G898), .A2(G224), .ZN(n1090) );
NAND3_X1 U781 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1088) );
XNOR2_X1 U782 ( .A(n1094), .B(KEYINPUT33), .ZN(n1093) );
NAND2_X1 U783 ( .A1(n1095), .A2(n1096), .ZN(n1091) );
XOR2_X1 U784 ( .A(KEYINPUT23), .B(n1097), .Z(n1095) );
NOR2_X1 U785 ( .A1(n1098), .A2(G953), .ZN(n1086) );
NOR2_X1 U786 ( .A1(n1099), .A2(n1100), .ZN(G66) );
XNOR2_X1 U787 ( .A(n1101), .B(n1102), .ZN(n1100) );
NOR2_X1 U788 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NOR2_X1 U789 ( .A1(n1099), .A2(n1105), .ZN(G63) );
XNOR2_X1 U790 ( .A(n1106), .B(n1107), .ZN(n1105) );
NOR2_X1 U791 ( .A1(n1108), .A2(n1104), .ZN(n1107) );
INV_X1 U792 ( .A(G478), .ZN(n1108) );
NOR3_X1 U793 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(G60) );
AND2_X1 U794 ( .A1(KEYINPUT6), .A2(n1099), .ZN(n1111) );
NOR3_X1 U795 ( .A1(KEYINPUT6), .A2(n1045), .A3(n1027), .ZN(n1110) );
INV_X1 U796 ( .A(G952), .ZN(n1045) );
XNOR2_X1 U797 ( .A(n1112), .B(n1113), .ZN(n1109) );
NOR2_X1 U798 ( .A1(n1114), .A2(n1104), .ZN(n1113) );
XNOR2_X1 U799 ( .A(G104), .B(n1115), .ZN(G6) );
NAND3_X1 U800 ( .A1(n1013), .A2(n1033), .A3(n1116), .ZN(n1115) );
NOR3_X1 U801 ( .A1(n1035), .A2(n1117), .A3(n1118), .ZN(n1116) );
XNOR2_X1 U802 ( .A(n1119), .B(KEYINPUT47), .ZN(n1118) );
NOR2_X1 U803 ( .A1(n1099), .A2(n1120), .ZN(G57) );
XOR2_X1 U804 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U805 ( .A(KEYINPUT5), .B(n1123), .Z(n1122) );
NOR2_X1 U806 ( .A1(n1124), .A2(n1104), .ZN(n1123) );
XOR2_X1 U807 ( .A(n1125), .B(n1126), .Z(n1121) );
NOR2_X1 U808 ( .A1(n1099), .A2(n1127), .ZN(G54) );
XOR2_X1 U809 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U810 ( .A1(n1065), .A2(n1104), .ZN(n1129) );
NAND2_X1 U811 ( .A1(n1130), .A2(KEYINPUT56), .ZN(n1128) );
XOR2_X1 U812 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U813 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U814 ( .A1(n1135), .A2(KEYINPUT57), .ZN(n1134) );
XNOR2_X1 U815 ( .A(n1084), .B(n1136), .ZN(n1135) );
XNOR2_X1 U816 ( .A(G143), .B(n1137), .ZN(n1084) );
XOR2_X1 U817 ( .A(n1138), .B(n1139), .Z(n1131) );
XNOR2_X1 U818 ( .A(n1140), .B(G110), .ZN(n1139) );
NOR2_X1 U819 ( .A1(n1099), .A2(n1141), .ZN(G51) );
XOR2_X1 U820 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U821 ( .A(n1144), .B(n1145), .Z(n1143) );
NAND2_X1 U822 ( .A1(KEYINPUT42), .A2(n1146), .ZN(n1144) );
XOR2_X1 U823 ( .A(n1147), .B(n1148), .Z(n1142) );
NOR2_X1 U824 ( .A1(n1063), .A2(n1104), .ZN(n1148) );
NAND2_X1 U825 ( .A1(G902), .A2(n1149), .ZN(n1104) );
NAND2_X1 U826 ( .A1(n1150), .A2(n1098), .ZN(n1149) );
INV_X1 U827 ( .A(n1002), .ZN(n1098) );
NAND4_X1 U828 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1002) );
AND4_X1 U829 ( .A1(n1155), .A2(n996), .A3(n1156), .A4(n1157), .ZN(n1154) );
NAND3_X1 U830 ( .A1(n1014), .A2(n1033), .A3(n1158), .ZN(n996) );
AND2_X1 U831 ( .A1(n1159), .A2(n1160), .ZN(n1153) );
NAND3_X1 U832 ( .A1(n1158), .A2(n1033), .A3(n1013), .ZN(n1151) );
XOR2_X1 U833 ( .A(n1000), .B(KEYINPUT55), .Z(n1150) );
NAND4_X1 U834 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1000) );
NOR4_X1 U835 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
NOR2_X1 U836 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
NOR3_X1 U837 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1169) );
NOR3_X1 U838 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1173) );
AND2_X1 U839 ( .A1(n1174), .A2(n1177), .ZN(n1172) );
INV_X1 U840 ( .A(KEYINPUT39), .ZN(n1174) );
INV_X1 U841 ( .A(n1178), .ZN(n1171) );
NOR3_X1 U842 ( .A1(n1020), .A2(KEYINPUT12), .A3(n1179), .ZN(n1166) );
NOR2_X1 U843 ( .A1(n1180), .A2(n1025), .ZN(n1165) );
NOR2_X1 U844 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NOR2_X1 U845 ( .A1(n1183), .A2(n1006), .ZN(n1182) );
NOR2_X1 U846 ( .A1(n1179), .A2(n1184), .ZN(n1181) );
INV_X1 U847 ( .A(KEYINPUT12), .ZN(n1184) );
OR3_X1 U848 ( .A1(n1011), .A2(n1035), .A3(n1183), .ZN(n1163) );
NAND2_X1 U849 ( .A1(KEYINPUT51), .A2(n1185), .ZN(n1147) );
NOR2_X1 U850 ( .A1(n1027), .A2(G952), .ZN(n1099) );
XNOR2_X1 U851 ( .A(G146), .B(n1161), .ZN(G48) );
NAND2_X1 U852 ( .A1(n1013), .A2(n1177), .ZN(n1161) );
XNOR2_X1 U853 ( .A(n1186), .B(n1187), .ZN(G45) );
NOR3_X1 U854 ( .A1(n1179), .A2(KEYINPUT18), .A3(n1025), .ZN(n1187) );
NAND3_X1 U855 ( .A1(n1052), .A2(n1188), .A3(n1189), .ZN(n1179) );
XOR2_X1 U856 ( .A(n1190), .B(n1191), .Z(G42) );
NOR3_X1 U857 ( .A1(n1192), .A2(n1011), .A3(n1183), .ZN(n1191) );
INV_X1 U858 ( .A(n1029), .ZN(n1011) );
XNOR2_X1 U859 ( .A(KEYINPUT4), .B(n1035), .ZN(n1192) );
NAND2_X1 U860 ( .A1(KEYINPUT32), .A2(n1140), .ZN(n1190) );
INV_X1 U861 ( .A(G140), .ZN(n1140) );
XNOR2_X1 U862 ( .A(G137), .B(n1162), .ZN(G39) );
NAND4_X1 U863 ( .A1(n1029), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1162) );
NOR2_X1 U864 ( .A1(n1196), .A2(n1035), .ZN(n1194) );
XOR2_X1 U865 ( .A(n1197), .B(n1198), .Z(G36) );
NOR2_X1 U866 ( .A1(n1178), .A2(n1199), .ZN(n1198) );
XNOR2_X1 U867 ( .A(KEYINPUT11), .B(n1170), .ZN(n1199) );
INV_X1 U868 ( .A(n1014), .ZN(n1170) );
XNOR2_X1 U869 ( .A(G134), .B(KEYINPUT13), .ZN(n1197) );
XNOR2_X1 U870 ( .A(n1083), .B(n1168), .ZN(G33) );
NOR2_X1 U871 ( .A1(n1200), .A2(n1178), .ZN(n1168) );
NAND2_X1 U872 ( .A1(n1189), .A2(n1029), .ZN(n1178) );
NOR2_X1 U873 ( .A1(n1022), .A2(n1061), .ZN(n1029) );
INV_X1 U874 ( .A(n1021), .ZN(n1061) );
NOR3_X1 U875 ( .A1(n1035), .A2(n1196), .A3(n1041), .ZN(n1189) );
XNOR2_X1 U876 ( .A(G128), .B(n1201), .ZN(G30) );
NAND2_X1 U877 ( .A1(n1177), .A2(n1014), .ZN(n1201) );
NOR2_X1 U878 ( .A1(n1175), .A2(n1196), .ZN(n1177) );
INV_X1 U879 ( .A(n1176), .ZN(n1196) );
NAND4_X1 U880 ( .A1(n1195), .A2(n1202), .A3(n1020), .A4(n1044), .ZN(n1175) );
XNOR2_X1 U881 ( .A(n1155), .B(n1203), .ZN(G3) );
XOR2_X1 U882 ( .A(KEYINPUT27), .B(G101), .Z(n1203) );
NAND3_X1 U883 ( .A1(n1015), .A2(n1158), .A3(n1204), .ZN(n1155) );
XNOR2_X1 U884 ( .A(n1205), .B(n1206), .ZN(G27) );
NOR4_X1 U885 ( .A1(n1025), .A2(n1183), .A3(n1207), .A4(n1208), .ZN(n1206) );
XNOR2_X1 U886 ( .A(KEYINPUT35), .B(n1006), .ZN(n1208) );
XOR2_X1 U887 ( .A(KEYINPUT43), .B(KEYINPUT31), .Z(n1207) );
NAND4_X1 U888 ( .A1(n1013), .A2(n1043), .A3(n1044), .A4(n1176), .ZN(n1183) );
NAND2_X1 U889 ( .A1(n1007), .A2(n1209), .ZN(n1176) );
NAND4_X1 U890 ( .A1(G902), .A2(G953), .A3(n1210), .A4(n1211), .ZN(n1209) );
INV_X1 U891 ( .A(G900), .ZN(n1211) );
INV_X1 U892 ( .A(n1200), .ZN(n1013) );
XNOR2_X1 U893 ( .A(G122), .B(n1152), .ZN(G24) );
NAND4_X1 U894 ( .A1(n1212), .A2(n1033), .A3(n1052), .A4(n1188), .ZN(n1152) );
INV_X1 U895 ( .A(n1005), .ZN(n1033) );
NAND2_X1 U896 ( .A1(n1213), .A2(n1043), .ZN(n1005) );
XNOR2_X1 U897 ( .A(G119), .B(n1160), .ZN(G21) );
NAND3_X1 U898 ( .A1(n1195), .A2(n1193), .A3(n1212), .ZN(n1160) );
XOR2_X1 U899 ( .A(n1159), .B(n1214), .Z(G18) );
NAND2_X1 U900 ( .A1(KEYINPUT25), .A2(G116), .ZN(n1214) );
NAND3_X1 U901 ( .A1(n1204), .A2(n1014), .A3(n1212), .ZN(n1159) );
NOR3_X1 U902 ( .A1(n1025), .A2(n1117), .A3(n1006), .ZN(n1212) );
NOR2_X1 U903 ( .A1(n1052), .A2(n1215), .ZN(n1014) );
XOR2_X1 U904 ( .A(n1157), .B(n1216), .Z(G15) );
XOR2_X1 U905 ( .A(KEYINPUT59), .B(G113), .Z(n1216) );
NAND3_X1 U906 ( .A1(n1039), .A2(n1204), .A3(n1217), .ZN(n1157) );
NOR3_X1 U907 ( .A1(n1200), .A2(n1117), .A3(n1119), .ZN(n1217) );
NAND2_X1 U908 ( .A1(n1215), .A2(n1052), .ZN(n1200) );
INV_X1 U909 ( .A(n1188), .ZN(n1215) );
INV_X1 U910 ( .A(n1041), .ZN(n1204) );
NAND2_X1 U911 ( .A1(n1213), .A2(n1195), .ZN(n1041) );
INV_X1 U912 ( .A(n1006), .ZN(n1039) );
NAND2_X1 U913 ( .A1(n1038), .A2(n1218), .ZN(n1006) );
XNOR2_X1 U914 ( .A(G110), .B(n1156), .ZN(G12) );
NAND3_X1 U915 ( .A1(n1158), .A2(n1043), .A3(n1193), .ZN(n1156) );
NOR2_X1 U916 ( .A1(n1017), .A2(n1213), .ZN(n1193) );
INV_X1 U917 ( .A(n1044), .ZN(n1213) );
XOR2_X1 U918 ( .A(n1219), .B(n1103), .Z(n1044) );
NAND2_X1 U919 ( .A1(G217), .A2(n1220), .ZN(n1103) );
NAND2_X1 U920 ( .A1(n1102), .A2(n1221), .ZN(n1219) );
XOR2_X1 U921 ( .A(n1222), .B(n1223), .Z(n1102) );
XOR2_X1 U922 ( .A(n1224), .B(n1225), .Z(n1223) );
XNOR2_X1 U923 ( .A(G119), .B(n1226), .ZN(n1225) );
XOR2_X1 U924 ( .A(KEYINPUT21), .B(G137), .Z(n1224) );
XOR2_X1 U925 ( .A(n1227), .B(n1077), .Z(n1222) );
XOR2_X1 U926 ( .A(n1228), .B(n1137), .Z(n1227) );
NAND3_X1 U927 ( .A1(n1229), .A2(G221), .A3(KEYINPUT9), .ZN(n1228) );
INV_X1 U928 ( .A(n1015), .ZN(n1017) );
NOR2_X1 U929 ( .A1(n1188), .A2(n1052), .ZN(n1015) );
XOR2_X1 U930 ( .A(n1230), .B(n1114), .Z(n1052) );
INV_X1 U931 ( .A(G475), .ZN(n1114) );
NAND2_X1 U932 ( .A1(n1221), .A2(n1112), .ZN(n1230) );
XNOR2_X1 U933 ( .A(n1231), .B(n1232), .ZN(n1112) );
XOR2_X1 U934 ( .A(n1077), .B(n1233), .Z(n1232) );
XOR2_X1 U935 ( .A(G104), .B(n1234), .Z(n1233) );
NOR2_X1 U936 ( .A1(KEYINPUT0), .A2(n1235), .ZN(n1234) );
XOR2_X1 U937 ( .A(n1236), .B(n1237), .Z(n1235) );
NAND2_X1 U938 ( .A1(KEYINPUT3), .A2(n1186), .ZN(n1237) );
INV_X1 U939 ( .A(G143), .ZN(n1186) );
NAND2_X1 U940 ( .A1(n1238), .A2(G214), .ZN(n1236) );
XNOR2_X1 U941 ( .A(n1205), .B(G140), .ZN(n1077) );
INV_X1 U942 ( .A(G125), .ZN(n1205) );
XOR2_X1 U943 ( .A(n1239), .B(n1240), .Z(n1231) );
XNOR2_X1 U944 ( .A(G146), .B(n1083), .ZN(n1240) );
XNOR2_X1 U945 ( .A(G113), .B(G122), .ZN(n1239) );
NAND2_X1 U946 ( .A1(n1055), .A2(n1053), .ZN(n1188) );
NAND2_X1 U947 ( .A1(n1241), .A2(n1242), .ZN(n1053) );
OR2_X1 U948 ( .A1(n1242), .A2(n1241), .ZN(n1055) );
AND2_X1 U949 ( .A1(n1221), .A2(n1106), .ZN(n1241) );
XNOR2_X1 U950 ( .A(n1243), .B(n1244), .ZN(n1106) );
XOR2_X1 U951 ( .A(n1245), .B(n1246), .Z(n1244) );
NAND2_X1 U952 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND2_X1 U953 ( .A1(G116), .A2(n1249), .ZN(n1248) );
XOR2_X1 U954 ( .A(n1250), .B(KEYINPUT24), .Z(n1247) );
OR2_X1 U955 ( .A1(n1249), .A2(G116), .ZN(n1250) );
NAND3_X1 U956 ( .A1(G217), .A2(n1229), .A3(KEYINPUT29), .ZN(n1245) );
AND2_X1 U957 ( .A1(G234), .A2(n1027), .ZN(n1229) );
XOR2_X1 U958 ( .A(n1251), .B(n1252), .Z(n1243) );
XNOR2_X1 U959 ( .A(n1253), .B(G107), .ZN(n1252) );
NAND2_X1 U960 ( .A1(n1254), .A2(KEYINPUT10), .ZN(n1251) );
XNOR2_X1 U961 ( .A(G128), .B(G143), .ZN(n1254) );
XOR2_X1 U962 ( .A(G478), .B(KEYINPUT37), .Z(n1242) );
XNOR2_X1 U963 ( .A(n1195), .B(KEYINPUT30), .ZN(n1043) );
XOR2_X1 U964 ( .A(n1054), .B(KEYINPUT28), .Z(n1195) );
XNOR2_X1 U965 ( .A(n1255), .B(n1124), .ZN(n1054) );
INV_X1 U966 ( .A(G472), .ZN(n1124) );
NAND3_X1 U967 ( .A1(n1256), .A2(n1257), .A3(n1221), .ZN(n1255) );
NAND2_X1 U968 ( .A1(KEYINPUT61), .A2(n1258), .ZN(n1257) );
XOR2_X1 U969 ( .A(n1259), .B(n1126), .Z(n1258) );
NAND3_X1 U970 ( .A1(n1126), .A2(n1259), .A3(n1260), .ZN(n1256) );
INV_X1 U971 ( .A(KEYINPUT61), .ZN(n1260) );
XOR2_X1 U972 ( .A(n1125), .B(KEYINPUT46), .Z(n1259) );
XOR2_X1 U973 ( .A(n1261), .B(n1262), .Z(n1125) );
XOR2_X1 U974 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U975 ( .A(n1265), .B(KEYINPUT36), .Z(n1261) );
XNOR2_X1 U976 ( .A(n1266), .B(G101), .ZN(n1126) );
NAND2_X1 U977 ( .A1(n1238), .A2(G210), .ZN(n1266) );
NOR2_X1 U978 ( .A1(G953), .A2(G237), .ZN(n1238) );
NOR3_X1 U979 ( .A1(n1119), .A2(n1117), .A3(n1035), .ZN(n1158) );
INV_X1 U980 ( .A(n1202), .ZN(n1035) );
NOR2_X1 U981 ( .A1(n1038), .A2(n1037), .ZN(n1202) );
INV_X1 U982 ( .A(n1218), .ZN(n1037) );
NAND2_X1 U983 ( .A1(G221), .A2(n1220), .ZN(n1218) );
NAND2_X1 U984 ( .A1(n1267), .A2(G234), .ZN(n1220) );
XNOR2_X1 U985 ( .A(G902), .B(KEYINPUT14), .ZN(n1267) );
XOR2_X1 U986 ( .A(n1064), .B(n1268), .Z(n1038) );
NOR2_X1 U987 ( .A1(KEYINPUT40), .A2(n1065), .ZN(n1268) );
INV_X1 U988 ( .A(G469), .ZN(n1065) );
NAND2_X1 U989 ( .A1(n1221), .A2(n1269), .ZN(n1064) );
XOR2_X1 U990 ( .A(n1270), .B(n1271), .Z(n1269) );
XNOR2_X1 U991 ( .A(n1272), .B(n1136), .ZN(n1271) );
XOR2_X1 U992 ( .A(n1273), .B(n1264), .Z(n1272) );
XNOR2_X1 U993 ( .A(n1133), .B(n1137), .ZN(n1264) );
NAND2_X1 U994 ( .A1(n1274), .A2(n1275), .ZN(n1133) );
NAND2_X1 U995 ( .A1(n1276), .A2(n1083), .ZN(n1275) );
XOR2_X1 U996 ( .A(KEYINPUT62), .B(n1277), .Z(n1274) );
NOR2_X1 U997 ( .A1(n1276), .A2(n1083), .ZN(n1277) );
INV_X1 U998 ( .A(G131), .ZN(n1083) );
NAND2_X1 U999 ( .A1(n1278), .A2(n1279), .ZN(n1276) );
OR2_X1 U1000 ( .A1(n1085), .A2(KEYINPUT8), .ZN(n1279) );
XNOR2_X1 U1001 ( .A(n1253), .B(G137), .ZN(n1085) );
NAND3_X1 U1002 ( .A1(G137), .A2(n1253), .A3(KEYINPUT8), .ZN(n1278) );
INV_X1 U1003 ( .A(G134), .ZN(n1253) );
NAND2_X1 U1004 ( .A1(n1280), .A2(KEYINPUT17), .ZN(n1273) );
XOR2_X1 U1005 ( .A(n1138), .B(KEYINPUT2), .Z(n1280) );
NAND2_X1 U1006 ( .A1(G227), .A2(n1027), .ZN(n1138) );
XOR2_X1 U1007 ( .A(n1281), .B(n1282), .Z(n1270) );
NOR2_X1 U1008 ( .A1(KEYINPUT48), .A2(n1226), .ZN(n1282) );
XNOR2_X1 U1009 ( .A(G140), .B(G143), .ZN(n1281) );
AND2_X1 U1010 ( .A1(n1283), .A2(n1007), .ZN(n1117) );
NAND3_X1 U1011 ( .A1(n1210), .A2(n1027), .A3(G952), .ZN(n1007) );
NAND3_X1 U1012 ( .A1(n1094), .A2(n1210), .A3(G902), .ZN(n1283) );
NAND2_X1 U1013 ( .A1(G237), .A2(G234), .ZN(n1210) );
NOR2_X1 U1014 ( .A1(n1027), .A2(G898), .ZN(n1094) );
XOR2_X1 U1015 ( .A(n1020), .B(KEYINPUT58), .Z(n1119) );
INV_X1 U1016 ( .A(n1025), .ZN(n1020) );
NAND2_X1 U1017 ( .A1(n1022), .A2(n1021), .ZN(n1025) );
NAND2_X1 U1018 ( .A1(G214), .A2(n1284), .ZN(n1021) );
NAND2_X1 U1019 ( .A1(n1060), .A2(n1285), .ZN(n1022) );
NAND2_X1 U1020 ( .A1(n1286), .A2(n1063), .ZN(n1285) );
XNOR2_X1 U1021 ( .A(n1062), .B(KEYINPUT53), .ZN(n1286) );
OR2_X1 U1022 ( .A1(n1063), .A2(n1062), .ZN(n1060) );
AND2_X1 U1023 ( .A1(n1287), .A2(n1221), .ZN(n1062) );
XNOR2_X1 U1024 ( .A(G902), .B(KEYINPUT22), .ZN(n1221) );
XOR2_X1 U1025 ( .A(n1145), .B(n1288), .Z(n1287) );
XNOR2_X1 U1026 ( .A(n1289), .B(n1290), .ZN(n1288) );
NOR2_X1 U1027 ( .A1(KEYINPUT20), .A2(n1185), .ZN(n1290) );
XOR2_X1 U1028 ( .A(n1265), .B(n1137), .Z(n1185) );
XNOR2_X1 U1029 ( .A(n1291), .B(G146), .ZN(n1137) );
INV_X1 U1030 ( .A(G128), .ZN(n1291) );
OR2_X1 U1031 ( .A1(G143), .A2(KEYINPUT7), .ZN(n1265) );
NAND2_X1 U1032 ( .A1(KEYINPUT19), .A2(n1146), .ZN(n1289) );
NAND2_X1 U1033 ( .A1(n1092), .A2(n1292), .ZN(n1146) );
NAND2_X1 U1034 ( .A1(n1293), .A2(n1096), .ZN(n1292) );
XOR2_X1 U1035 ( .A(KEYINPUT50), .B(n1097), .Z(n1293) );
NAND2_X1 U1036 ( .A1(n1136), .A2(n1097), .ZN(n1092) );
XNOR2_X1 U1037 ( .A(n1294), .B(n1263), .ZN(n1097) );
XOR2_X1 U1038 ( .A(G113), .B(n1295), .Z(n1263) );
XOR2_X1 U1039 ( .A(G119), .B(G116), .Z(n1295) );
XOR2_X1 U1040 ( .A(n1296), .B(KEYINPUT52), .Z(n1294) );
NAND2_X1 U1041 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
NAND2_X1 U1042 ( .A1(G110), .A2(n1249), .ZN(n1298) );
INV_X1 U1043 ( .A(G122), .ZN(n1249) );
XOR2_X1 U1044 ( .A(n1299), .B(KEYINPUT54), .Z(n1297) );
NAND2_X1 U1045 ( .A1(G122), .A2(n1226), .ZN(n1299) );
INV_X1 U1046 ( .A(G110), .ZN(n1226) );
INV_X1 U1047 ( .A(n1096), .ZN(n1136) );
XNOR2_X1 U1048 ( .A(n1300), .B(n1301), .ZN(n1096) );
XOR2_X1 U1049 ( .A(KEYINPUT1), .B(G107), .Z(n1301) );
XNOR2_X1 U1050 ( .A(G101), .B(G104), .ZN(n1300) );
XNOR2_X1 U1051 ( .A(G125), .B(n1302), .ZN(n1145) );
AND2_X1 U1052 ( .A1(n1027), .A2(G224), .ZN(n1302) );
INV_X1 U1053 ( .A(G953), .ZN(n1027) );
NAND2_X1 U1054 ( .A1(G210), .A2(n1284), .ZN(n1063) );
NAND2_X1 U1055 ( .A1(n1303), .A2(n1304), .ZN(n1284) );
INV_X1 U1056 ( .A(G902), .ZN(n1304) );
INV_X1 U1057 ( .A(G237), .ZN(n1303) );
endmodule


