//Key = 0010111111101011011101000110000011101110101010000111000111110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314;

XOR2_X1 U734 ( .A(n999), .B(n1000), .Z(G9) );
NAND2_X1 U735 ( .A1(KEYINPUT10), .A2(n1001), .ZN(n999) );
INV_X1 U736 ( .A(G107), .ZN(n1001) );
NOR2_X1 U737 ( .A1(n1002), .A2(n1003), .ZN(G75) );
NOR4_X1 U738 ( .A1(G953), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1003) );
NOR2_X1 U739 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR2_X1 U740 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U741 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NOR2_X1 U742 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
NOR3_X1 U743 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NOR2_X1 U744 ( .A1(n1018), .A2(n1019), .ZN(n1013) );
INV_X1 U745 ( .A(n1020), .ZN(n1019) );
NOR2_X1 U746 ( .A1(n1021), .A2(n1022), .ZN(n1018) );
NOR2_X1 U747 ( .A1(n1023), .A2(n1016), .ZN(n1022) );
NOR2_X1 U748 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NOR2_X1 U749 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U750 ( .A1(n1028), .A2(n1015), .ZN(n1021) );
INV_X1 U751 ( .A(n1029), .ZN(n1015) );
NOR2_X1 U752 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR2_X1 U753 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR3_X1 U754 ( .A1(n1034), .A2(n1016), .A3(n1035), .ZN(n1009) );
NAND3_X1 U755 ( .A1(n1036), .A2(n1037), .A3(n1029), .ZN(n1034) );
NAND2_X1 U756 ( .A1(n1038), .A2(n1012), .ZN(n1037) );
OR3_X1 U757 ( .A1(n1039), .A2(n1040), .A3(n1038), .ZN(n1036) );
NOR3_X1 U758 ( .A1(n1004), .A2(G953), .A3(G952), .ZN(n1002) );
AND4_X1 U759 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1004) );
NOR3_X1 U760 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NOR2_X1 U761 ( .A1(KEYINPUT2), .A2(n1048), .ZN(n1046) );
NAND3_X1 U762 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1045) );
NAND3_X1 U763 ( .A1(KEYINPUT2), .A2(n1048), .A3(n1052), .ZN(n1050) );
NAND2_X1 U764 ( .A1(n1053), .A2(n1054), .ZN(n1049) );
NAND2_X1 U765 ( .A1(KEYINPUT2), .A2(n1055), .ZN(n1053) );
XNOR2_X1 U766 ( .A(KEYINPUT21), .B(n1048), .ZN(n1055) );
NOR3_X1 U767 ( .A1(n1056), .A2(n1057), .A3(n1038), .ZN(n1043) );
XOR2_X1 U768 ( .A(n1058), .B(n1059), .Z(n1056) );
NOR2_X1 U769 ( .A1(G469), .A2(KEYINPUT48), .ZN(n1059) );
XOR2_X1 U770 ( .A(KEYINPUT7), .B(n1060), .Z(n1042) );
XOR2_X1 U771 ( .A(KEYINPUT26), .B(n1033), .Z(n1041) );
XOR2_X1 U772 ( .A(n1061), .B(n1062), .Z(G72) );
NOR2_X1 U773 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U774 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NAND2_X1 U775 ( .A1(n1067), .A2(n1068), .ZN(n1061) );
NAND2_X1 U776 ( .A1(n1069), .A2(n1064), .ZN(n1068) );
XOR2_X1 U777 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND2_X1 U778 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
XOR2_X1 U779 ( .A(n1074), .B(KEYINPUT34), .Z(n1072) );
NAND2_X1 U780 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND3_X1 U781 ( .A1(n1071), .A2(G900), .A3(G953), .ZN(n1067) );
NOR2_X1 U782 ( .A1(KEYINPUT43), .A2(n1077), .ZN(n1071) );
XOR2_X1 U783 ( .A(n1078), .B(n1079), .Z(n1077) );
XOR2_X1 U784 ( .A(G137), .B(n1080), .Z(n1079) );
NOR2_X1 U785 ( .A1(KEYINPUT47), .A2(n1081), .ZN(n1080) );
XOR2_X1 U786 ( .A(n1082), .B(n1083), .Z(n1078) );
XOR2_X1 U787 ( .A(n1084), .B(n1085), .Z(G69) );
NAND2_X1 U788 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
OR3_X1 U789 ( .A1(n1088), .A2(G953), .A3(n1089), .ZN(n1087) );
NAND3_X1 U790 ( .A1(n1090), .A2(n1091), .A3(n1089), .ZN(n1086) );
XOR2_X1 U791 ( .A(KEYINPUT31), .B(n1088), .Z(n1090) );
NAND2_X1 U792 ( .A1(n1091), .A2(n1092), .ZN(n1084) );
NAND2_X1 U793 ( .A1(G953), .A2(n1093), .ZN(n1092) );
INV_X1 U794 ( .A(n1094), .ZN(n1091) );
NOR2_X1 U795 ( .A1(n1095), .A2(n1096), .ZN(G66) );
XOR2_X1 U796 ( .A(n1097), .B(KEYINPUT25), .Z(n1096) );
XOR2_X1 U797 ( .A(n1098), .B(n1099), .Z(n1095) );
AND3_X1 U798 ( .A1(n1100), .A2(n1101), .A3(G217), .ZN(n1099) );
NAND2_X1 U799 ( .A1(KEYINPUT19), .A2(n1102), .ZN(n1098) );
NOR2_X1 U800 ( .A1(n1103), .A2(n1104), .ZN(G63) );
XOR2_X1 U801 ( .A(n1105), .B(n1106), .Z(n1104) );
AND2_X1 U802 ( .A1(G478), .A2(n1100), .ZN(n1106) );
NAND2_X1 U803 ( .A1(KEYINPUT36), .A2(n1107), .ZN(n1105) );
NOR2_X1 U804 ( .A1(n1103), .A2(n1108), .ZN(G60) );
XNOR2_X1 U805 ( .A(n1109), .B(n1110), .ZN(n1108) );
XOR2_X1 U806 ( .A(KEYINPUT9), .B(n1111), .Z(n1110) );
AND2_X1 U807 ( .A1(G475), .A2(n1100), .ZN(n1111) );
XNOR2_X1 U808 ( .A(n1112), .B(n1113), .ZN(G6) );
NAND2_X1 U809 ( .A1(KEYINPUT6), .A2(n1114), .ZN(n1112) );
NOR2_X1 U810 ( .A1(n1115), .A2(n1116), .ZN(G57) );
XOR2_X1 U811 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U812 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U813 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U814 ( .A(n1123), .B(n1124), .Z(n1117) );
XOR2_X1 U815 ( .A(KEYINPUT63), .B(n1125), .Z(n1124) );
NOR2_X1 U816 ( .A1(KEYINPUT11), .A2(n1126), .ZN(n1125) );
AND2_X1 U817 ( .A1(G472), .A2(n1100), .ZN(n1123) );
NOR2_X1 U818 ( .A1(n1127), .A2(n1064), .ZN(n1115) );
XNOR2_X1 U819 ( .A(G952), .B(KEYINPUT33), .ZN(n1127) );
NOR3_X1 U820 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(G54) );
AND3_X1 U821 ( .A1(KEYINPUT29), .A2(G953), .A3(G952), .ZN(n1130) );
NOR2_X1 U822 ( .A1(KEYINPUT29), .A2(n1097), .ZN(n1129) );
XOR2_X1 U823 ( .A(n1131), .B(n1132), .Z(n1128) );
XOR2_X1 U824 ( .A(n1126), .B(n1133), .Z(n1132) );
XOR2_X1 U825 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND3_X1 U826 ( .A1(n1136), .A2(n1006), .A3(G469), .ZN(n1135) );
XNOR2_X1 U827 ( .A(KEYINPUT37), .B(n1137), .ZN(n1136) );
NAND2_X1 U828 ( .A1(n1138), .A2(n1139), .ZN(n1134) );
NAND3_X1 U829 ( .A1(n1140), .A2(n1141), .A3(KEYINPUT4), .ZN(n1139) );
XOR2_X1 U830 ( .A(n1142), .B(n1143), .Z(n1140) );
AND2_X1 U831 ( .A1(G140), .A2(KEYINPUT40), .ZN(n1143) );
NAND2_X1 U832 ( .A1(n1144), .A2(n1145), .ZN(n1138) );
NAND2_X1 U833 ( .A1(KEYINPUT4), .A2(n1141), .ZN(n1145) );
XOR2_X1 U834 ( .A(n1142), .B(n1146), .Z(n1144) );
NOR2_X1 U835 ( .A1(G140), .A2(n1147), .ZN(n1146) );
INV_X1 U836 ( .A(KEYINPUT40), .ZN(n1147) );
XOR2_X1 U837 ( .A(n1082), .B(n1148), .Z(n1131) );
NOR3_X1 U838 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(G51) );
NOR3_X1 U839 ( .A1(n1152), .A2(G953), .A3(G952), .ZN(n1151) );
INV_X1 U840 ( .A(KEYINPUT28), .ZN(n1152) );
NOR2_X1 U841 ( .A1(KEYINPUT28), .A2(n1097), .ZN(n1150) );
INV_X1 U842 ( .A(n1103), .ZN(n1097) );
NOR2_X1 U843 ( .A1(n1064), .A2(G952), .ZN(n1103) );
NOR2_X1 U844 ( .A1(n1153), .A2(n1154), .ZN(n1149) );
XOR2_X1 U845 ( .A(n1155), .B(KEYINPUT17), .Z(n1154) );
NAND2_X1 U846 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U847 ( .A1(n1100), .A2(n1052), .ZN(n1157) );
INV_X1 U848 ( .A(n1158), .ZN(n1100) );
NOR3_X1 U849 ( .A1(n1156), .A2(n1054), .A3(n1158), .ZN(n1153) );
NAND2_X1 U850 ( .A1(n1137), .A2(n1006), .ZN(n1158) );
NAND4_X1 U851 ( .A1(n1159), .A2(n1088), .A3(n1075), .A4(n1073), .ZN(n1006) );
AND4_X1 U852 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1073) );
AND3_X1 U853 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1075) );
AND4_X1 U854 ( .A1(n1113), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1088) );
NOR4_X1 U855 ( .A1(n1000), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1169) );
INV_X1 U856 ( .A(n1173), .ZN(n1171) );
NOR3_X1 U857 ( .A1(n1174), .A2(n1016), .A3(n1175), .ZN(n1000) );
INV_X1 U858 ( .A(n1176), .ZN(n1016) );
NAND2_X1 U859 ( .A1(n1031), .A2(n1177), .ZN(n1168) );
NAND2_X1 U860 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND2_X1 U861 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U862 ( .A(n1174), .B(KEYINPUT18), .Z(n1180) );
NAND2_X1 U863 ( .A1(n1182), .A2(n1183), .ZN(n1178) );
NAND3_X1 U864 ( .A1(n1183), .A2(n1176), .A3(n1040), .ZN(n1113) );
XOR2_X1 U865 ( .A(n1076), .B(KEYINPUT22), .Z(n1159) );
XNOR2_X1 U866 ( .A(G902), .B(KEYINPUT32), .ZN(n1137) );
XNOR2_X1 U867 ( .A(n1184), .B(n1089), .ZN(n1156) );
NAND2_X1 U868 ( .A1(KEYINPUT15), .A2(n1185), .ZN(n1184) );
NAND2_X1 U869 ( .A1(n1186), .A2(n1187), .ZN(G48) );
NAND2_X1 U870 ( .A1(G146), .A2(n1160), .ZN(n1187) );
XOR2_X1 U871 ( .A(n1188), .B(KEYINPUT27), .Z(n1186) );
OR2_X1 U872 ( .A1(n1160), .A2(G146), .ZN(n1188) );
NAND3_X1 U873 ( .A1(n1040), .A2(n1025), .A3(n1189), .ZN(n1160) );
XOR2_X1 U874 ( .A(n1190), .B(n1161), .Z(G45) );
NAND4_X1 U875 ( .A1(n1191), .A2(n1192), .A3(n1025), .A4(n1193), .ZN(n1161) );
XNOR2_X1 U876 ( .A(G140), .B(n1162), .ZN(G42) );
NAND3_X1 U877 ( .A1(n1194), .A2(n1195), .A3(n1029), .ZN(n1162) );
XOR2_X1 U878 ( .A(n1196), .B(n1163), .Z(G39) );
NAND3_X1 U879 ( .A1(n1189), .A2(n1182), .A3(n1029), .ZN(n1163) );
XNOR2_X1 U880 ( .A(G134), .B(n1166), .ZN(G36) );
NAND3_X1 U881 ( .A1(n1192), .A2(n1039), .A3(n1029), .ZN(n1166) );
XNOR2_X1 U882 ( .A(G131), .B(n1076), .ZN(G33) );
NAND3_X1 U883 ( .A1(n1192), .A2(n1040), .A3(n1029), .ZN(n1076) );
NOR2_X1 U884 ( .A1(n1026), .A2(n1057), .ZN(n1029) );
INV_X1 U885 ( .A(n1027), .ZN(n1057) );
AND3_X1 U886 ( .A1(n1195), .A2(n1197), .A3(n1031), .ZN(n1192) );
XNOR2_X1 U887 ( .A(G128), .B(n1164), .ZN(G30) );
NAND3_X1 U888 ( .A1(n1039), .A2(n1025), .A3(n1189), .ZN(n1164) );
AND4_X1 U889 ( .A1(n1195), .A2(n1060), .A3(n1033), .A4(n1197), .ZN(n1189) );
INV_X1 U890 ( .A(n1174), .ZN(n1039) );
NAND2_X1 U891 ( .A1(n1198), .A2(n1199), .ZN(G3) );
NAND2_X1 U892 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U893 ( .A(KEYINPUT51), .B(n1202), .Z(n1198) );
NOR2_X1 U894 ( .A1(n1200), .A2(n1201), .ZN(n1202) );
INV_X1 U895 ( .A(G101), .ZN(n1201) );
AND4_X1 U896 ( .A1(n1182), .A2(n1031), .A3(n1203), .A4(n1204), .ZN(n1200) );
OR2_X1 U897 ( .A1(n1183), .A2(KEYINPUT0), .ZN(n1204) );
NAND2_X1 U898 ( .A1(KEYINPUT0), .A2(n1205), .ZN(n1203) );
NAND3_X1 U899 ( .A1(n1195), .A2(n1206), .A3(n1207), .ZN(n1205) );
INV_X1 U900 ( .A(n1017), .ZN(n1195) );
INV_X1 U901 ( .A(n1012), .ZN(n1182) );
XOR2_X1 U902 ( .A(G125), .B(n1208), .Z(G27) );
NOR2_X1 U903 ( .A1(KEYINPUT20), .A2(n1165), .ZN(n1208) );
NAND3_X1 U904 ( .A1(n1020), .A2(n1025), .A3(n1194), .ZN(n1165) );
AND4_X1 U905 ( .A1(n1209), .A2(n1040), .A3(n1060), .A4(n1197), .ZN(n1194) );
NAND2_X1 U906 ( .A1(n1008), .A2(n1210), .ZN(n1197) );
NAND4_X1 U907 ( .A1(G902), .A2(G953), .A3(n1211), .A4(n1066), .ZN(n1210) );
INV_X1 U908 ( .A(G900), .ZN(n1066) );
INV_X1 U909 ( .A(n1032), .ZN(n1060) );
XOR2_X1 U910 ( .A(n1212), .B(n1167), .Z(G24) );
NAND4_X1 U911 ( .A1(n1191), .A2(n1181), .A3(n1176), .A4(n1193), .ZN(n1167) );
NAND2_X1 U912 ( .A1(n1213), .A2(n1214), .ZN(n1176) );
NAND3_X1 U913 ( .A1(n1215), .A2(n1209), .A3(n1216), .ZN(n1214) );
INV_X1 U914 ( .A(KEYINPUT52), .ZN(n1216) );
NAND2_X1 U915 ( .A1(KEYINPUT52), .A2(n1031), .ZN(n1213) );
INV_X1 U916 ( .A(n1217), .ZN(n1031) );
INV_X1 U917 ( .A(n1218), .ZN(n1181) );
XNOR2_X1 U918 ( .A(n1172), .B(n1219), .ZN(G21) );
NAND2_X1 U919 ( .A1(G119), .A2(n1220), .ZN(n1219) );
XOR2_X1 U920 ( .A(KEYINPUT60), .B(KEYINPUT14), .Z(n1220) );
NOR4_X1 U921 ( .A1(n1218), .A2(n1012), .A3(n1032), .A4(n1209), .ZN(n1172) );
XOR2_X1 U922 ( .A(G116), .B(n1221), .Z(G18) );
NOR3_X1 U923 ( .A1(n1218), .A2(n1217), .A3(n1174), .ZN(n1221) );
NAND2_X1 U924 ( .A1(n1193), .A2(n1222), .ZN(n1174) );
NAND3_X1 U925 ( .A1(n1025), .A2(n1206), .A3(n1020), .ZN(n1218) );
XOR2_X1 U926 ( .A(G113), .B(n1223), .Z(G15) );
NOR2_X1 U927 ( .A1(KEYINPUT41), .A2(n1173), .ZN(n1223) );
NAND3_X1 U928 ( .A1(n1040), .A2(n1020), .A3(n1224), .ZN(n1173) );
NOR3_X1 U929 ( .A1(n1217), .A2(n1225), .A3(n1207), .ZN(n1224) );
NAND2_X1 U930 ( .A1(n1215), .A2(n1033), .ZN(n1217) );
XOR2_X1 U931 ( .A(n1032), .B(KEYINPUT16), .Z(n1215) );
NOR2_X1 U932 ( .A1(n1035), .A2(n1038), .ZN(n1020) );
INV_X1 U933 ( .A(n1226), .ZN(n1038) );
NOR2_X1 U934 ( .A1(n1222), .A2(n1193), .ZN(n1040) );
INV_X1 U935 ( .A(n1051), .ZN(n1193) );
XOR2_X1 U936 ( .A(G110), .B(n1170), .Z(G12) );
NOR4_X1 U937 ( .A1(n1012), .A2(n1175), .A3(n1033), .A4(n1032), .ZN(n1170) );
XOR2_X1 U938 ( .A(n1227), .B(n1228), .Z(n1032) );
NOR2_X1 U939 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
XNOR2_X1 U940 ( .A(KEYINPUT53), .B(n1101), .ZN(n1230) );
NAND2_X1 U941 ( .A1(n1102), .A2(n1231), .ZN(n1227) );
XOR2_X1 U942 ( .A(n1232), .B(n1233), .Z(n1102) );
XOR2_X1 U943 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U944 ( .A(n1236), .B(G110), .Z(n1235) );
NAND2_X1 U945 ( .A1(n1237), .A2(G221), .ZN(n1236) );
INV_X1 U946 ( .A(n1238), .ZN(n1237) );
XNOR2_X1 U947 ( .A(G119), .B(KEYINPUT1), .ZN(n1234) );
XNOR2_X1 U948 ( .A(n1239), .B(n1240), .ZN(n1232) );
XOR2_X1 U949 ( .A(n1241), .B(n1242), .Z(n1240) );
NOR2_X1 U950 ( .A1(G137), .A2(KEYINPUT13), .ZN(n1241) );
INV_X1 U951 ( .A(n1209), .ZN(n1033) );
XOR2_X1 U952 ( .A(n1243), .B(G472), .Z(n1209) );
NAND2_X1 U953 ( .A1(n1244), .A2(n1231), .ZN(n1243) );
XOR2_X1 U954 ( .A(n1245), .B(n1246), .Z(n1244) );
XOR2_X1 U955 ( .A(n1119), .B(n1126), .Z(n1246) );
INV_X1 U956 ( .A(n1247), .ZN(n1126) );
XOR2_X1 U957 ( .A(n1248), .B(n1249), .Z(n1245) );
NOR2_X1 U958 ( .A1(KEYINPUT39), .A2(n1250), .ZN(n1249) );
NAND2_X1 U959 ( .A1(KEYINPUT5), .A2(n1121), .ZN(n1248) );
XOR2_X1 U960 ( .A(n1251), .B(n1252), .Z(n1121) );
NAND2_X1 U961 ( .A1(n1253), .A2(G210), .ZN(n1251) );
INV_X1 U962 ( .A(n1183), .ZN(n1175) );
NOR3_X1 U963 ( .A1(n1207), .A2(n1225), .A3(n1017), .ZN(n1183) );
NAND2_X1 U964 ( .A1(n1035), .A2(n1226), .ZN(n1017) );
NAND2_X1 U965 ( .A1(G221), .A2(n1101), .ZN(n1226) );
NAND2_X1 U966 ( .A1(G234), .A2(n1231), .ZN(n1101) );
XNOR2_X1 U967 ( .A(n1058), .B(G469), .ZN(n1035) );
NAND2_X1 U968 ( .A1(n1254), .A2(n1231), .ZN(n1058) );
XOR2_X1 U969 ( .A(n1255), .B(n1256), .Z(n1254) );
XOR2_X1 U970 ( .A(n1257), .B(n1142), .Z(n1256) );
NOR2_X1 U971 ( .A1(n1065), .A2(G953), .ZN(n1142) );
INV_X1 U972 ( .A(G227), .ZN(n1065) );
NAND2_X1 U973 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NAND2_X1 U974 ( .A1(n1247), .A2(n1260), .ZN(n1259) );
XOR2_X1 U975 ( .A(KEYINPUT8), .B(n1261), .Z(n1258) );
NOR2_X1 U976 ( .A1(n1247), .A2(n1260), .ZN(n1261) );
XOR2_X1 U977 ( .A(n1262), .B(n1263), .Z(n1260) );
INV_X1 U978 ( .A(n1082), .ZN(n1263) );
XOR2_X1 U979 ( .A(n1190), .B(n1239), .Z(n1082) );
XOR2_X1 U980 ( .A(G128), .B(G146), .Z(n1239) );
NAND2_X1 U981 ( .A1(KEYINPUT62), .A2(n1264), .ZN(n1262) );
XNOR2_X1 U982 ( .A(G131), .B(n1265), .ZN(n1247) );
NOR2_X1 U983 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XOR2_X1 U984 ( .A(KEYINPUT61), .B(n1268), .Z(n1267) );
NOR2_X1 U985 ( .A1(n1081), .A2(n1196), .ZN(n1268) );
AND2_X1 U986 ( .A1(n1196), .A2(n1081), .ZN(n1266) );
XOR2_X1 U987 ( .A(G134), .B(KEYINPUT35), .Z(n1081) );
INV_X1 U988 ( .A(G137), .ZN(n1196) );
XOR2_X1 U989 ( .A(G140), .B(n1141), .Z(n1255) );
INV_X1 U990 ( .A(G110), .ZN(n1141) );
INV_X1 U991 ( .A(n1206), .ZN(n1225) );
NAND2_X1 U992 ( .A1(n1008), .A2(n1269), .ZN(n1206) );
NAND3_X1 U993 ( .A1(n1094), .A2(n1211), .A3(G902), .ZN(n1269) );
NOR2_X1 U994 ( .A1(G898), .A2(n1064), .ZN(n1094) );
NAND3_X1 U995 ( .A1(n1211), .A2(n1064), .A3(G952), .ZN(n1008) );
NAND2_X1 U996 ( .A1(G237), .A2(G234), .ZN(n1211) );
XNOR2_X1 U997 ( .A(n1025), .B(KEYINPUT46), .ZN(n1207) );
AND2_X1 U998 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U999 ( .A1(n1270), .A2(n1271), .ZN(n1027) );
XOR2_X1 U1000 ( .A(KEYINPUT3), .B(G214), .Z(n1270) );
XNOR2_X1 U1001 ( .A(n1048), .B(n1052), .ZN(n1026) );
INV_X1 U1002 ( .A(n1054), .ZN(n1052) );
NAND2_X1 U1003 ( .A1(G210), .A2(n1271), .ZN(n1054) );
NAND2_X1 U1004 ( .A1(n1272), .A2(n1231), .ZN(n1271) );
INV_X1 U1005 ( .A(G237), .ZN(n1272) );
NAND3_X1 U1006 ( .A1(n1273), .A2(n1231), .A3(n1274), .ZN(n1048) );
XOR2_X1 U1007 ( .A(n1275), .B(KEYINPUT23), .Z(n1274) );
OR2_X1 U1008 ( .A1(n1089), .A2(n1185), .ZN(n1275) );
NAND2_X1 U1009 ( .A1(n1185), .A2(n1089), .ZN(n1273) );
XNOR2_X1 U1010 ( .A(n1276), .B(n1277), .ZN(n1089) );
XOR2_X1 U1011 ( .A(n1250), .B(n1148), .Z(n1277) );
INV_X1 U1012 ( .A(n1264), .ZN(n1148) );
XOR2_X1 U1013 ( .A(n1278), .B(n1252), .Z(n1264) );
XOR2_X1 U1014 ( .A(G101), .B(KEYINPUT30), .Z(n1252) );
XOR2_X1 U1015 ( .A(n1114), .B(G107), .Z(n1278) );
INV_X1 U1016 ( .A(G104), .ZN(n1114) );
INV_X1 U1017 ( .A(n1122), .ZN(n1250) );
XOR2_X1 U1018 ( .A(n1279), .B(n1280), .Z(n1122) );
XOR2_X1 U1019 ( .A(KEYINPUT55), .B(G119), .Z(n1280) );
XOR2_X1 U1020 ( .A(n1281), .B(G116), .Z(n1279) );
INV_X1 U1021 ( .A(G113), .ZN(n1281) );
XOR2_X1 U1022 ( .A(n1212), .B(G110), .Z(n1276) );
XNOR2_X1 U1023 ( .A(n1282), .B(n1119), .ZN(n1185) );
XNOR2_X1 U1024 ( .A(n1283), .B(n1284), .ZN(n1119) );
NOR2_X1 U1025 ( .A1(G128), .A2(KEYINPUT24), .ZN(n1284) );
NAND2_X1 U1026 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
NAND2_X1 U1027 ( .A1(KEYINPUT12), .A2(n1287), .ZN(n1286) );
XOR2_X1 U1028 ( .A(n1190), .B(G146), .Z(n1287) );
OR3_X1 U1029 ( .A1(n1190), .A2(G146), .A3(KEYINPUT12), .ZN(n1285) );
XOR2_X1 U1030 ( .A(n1288), .B(n1289), .Z(n1282) );
NOR2_X1 U1031 ( .A1(G953), .A2(n1093), .ZN(n1289) );
INV_X1 U1032 ( .A(G224), .ZN(n1093) );
INV_X1 U1033 ( .A(G125), .ZN(n1288) );
NAND2_X1 U1034 ( .A1(n1051), .A2(n1222), .ZN(n1012) );
INV_X1 U1035 ( .A(n1191), .ZN(n1222) );
XNOR2_X1 U1036 ( .A(n1047), .B(KEYINPUT57), .ZN(n1191) );
XOR2_X1 U1037 ( .A(G475), .B(n1290), .Z(n1047) );
NOR2_X1 U1038 ( .A1(G902), .A2(n1109), .ZN(n1290) );
XNOR2_X1 U1039 ( .A(n1291), .B(n1292), .ZN(n1109) );
XOR2_X1 U1040 ( .A(G113), .B(n1293), .Z(n1292) );
XOR2_X1 U1041 ( .A(KEYINPUT38), .B(G122), .Z(n1293) );
XNOR2_X1 U1042 ( .A(n1294), .B(n1295), .ZN(n1291) );
NOR2_X1 U1043 ( .A1(G104), .A2(KEYINPUT45), .ZN(n1295) );
NOR2_X1 U1044 ( .A1(KEYINPUT54), .A2(n1296), .ZN(n1294) );
XNOR2_X1 U1045 ( .A(n1083), .B(n1297), .ZN(n1296) );
XNOR2_X1 U1046 ( .A(G146), .B(n1298), .ZN(n1297) );
NAND2_X1 U1047 ( .A1(n1299), .A2(KEYINPUT50), .ZN(n1298) );
XOR2_X1 U1048 ( .A(n1300), .B(G143), .Z(n1299) );
NAND2_X1 U1049 ( .A1(n1253), .A2(G214), .ZN(n1300) );
NOR2_X1 U1050 ( .A1(G953), .A2(G237), .ZN(n1253) );
XOR2_X1 U1051 ( .A(G131), .B(n1242), .Z(n1083) );
XOR2_X1 U1052 ( .A(G125), .B(G140), .Z(n1242) );
XOR2_X1 U1053 ( .A(n1301), .B(G478), .Z(n1051) );
NAND2_X1 U1054 ( .A1(n1107), .A2(n1231), .ZN(n1301) );
INV_X1 U1055 ( .A(G902), .ZN(n1231) );
XNOR2_X1 U1056 ( .A(n1302), .B(n1303), .ZN(n1107) );
NOR2_X1 U1057 ( .A1(n1238), .A2(n1229), .ZN(n1303) );
INV_X1 U1058 ( .A(G217), .ZN(n1229) );
NAND2_X1 U1059 ( .A1(G234), .A2(n1064), .ZN(n1238) );
INV_X1 U1060 ( .A(G953), .ZN(n1064) );
NAND3_X1 U1061 ( .A1(n1304), .A2(n1305), .A3(KEYINPUT59), .ZN(n1302) );
OR3_X1 U1062 ( .A1(n1306), .A2(n1307), .A3(KEYINPUT44), .ZN(n1305) );
NAND2_X1 U1063 ( .A1(n1308), .A2(KEYINPUT44), .ZN(n1304) );
XNOR2_X1 U1064 ( .A(n1309), .B(n1307), .ZN(n1308) );
XNOR2_X1 U1065 ( .A(n1310), .B(G134), .ZN(n1307) );
NAND2_X1 U1066 ( .A1(KEYINPUT49), .A2(n1311), .ZN(n1310) );
XNOR2_X1 U1067 ( .A(G128), .B(n1312), .ZN(n1311) );
NAND2_X1 U1068 ( .A1(KEYINPUT42), .A2(n1190), .ZN(n1312) );
INV_X1 U1069 ( .A(G143), .ZN(n1190) );
NAND2_X1 U1070 ( .A1(KEYINPUT58), .A2(n1306), .ZN(n1309) );
XOR2_X1 U1071 ( .A(n1313), .B(G107), .Z(n1306) );
NAND2_X1 U1072 ( .A1(n1314), .A2(KEYINPUT56), .ZN(n1313) );
XOR2_X1 U1073 ( .A(G116), .B(n1212), .Z(n1314) );
INV_X1 U1074 ( .A(G122), .ZN(n1212) );
endmodule


