//Key = 1010001000111101101111011110011110010110011011110101011011100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311;

XNOR2_X1 U720 ( .A(G107), .B(n998), .ZN(G9) );
NOR2_X1 U721 ( .A1(n999), .A2(n1000), .ZN(G75) );
NOR4_X1 U722 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n1000) );
XOR2_X1 U723 ( .A(KEYINPUT9), .B(n1005), .Z(n1002) );
NOR3_X1 U724 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n1005) );
XOR2_X1 U725 ( .A(KEYINPUT15), .B(n1009), .Z(n1008) );
NAND3_X1 U726 ( .A1(n1010), .A2(n1011), .A3(n1012), .ZN(n1006) );
NAND4_X1 U727 ( .A1(G952), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1001) );
NAND2_X1 U728 ( .A1(n1016), .A2(n1017), .ZN(n1013) );
NAND2_X1 U729 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND3_X1 U730 ( .A1(n1011), .A2(n1020), .A3(n1009), .ZN(n1019) );
NAND2_X1 U731 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U732 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U733 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U734 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
INV_X1 U735 ( .A(n1029), .ZN(n1025) );
NAND2_X1 U736 ( .A1(n1030), .A2(n1012), .ZN(n1021) );
NAND3_X1 U737 ( .A1(n1012), .A2(n1031), .A3(n1023), .ZN(n1018) );
NAND2_X1 U738 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U739 ( .A1(n1009), .A2(n1034), .ZN(n1033) );
NAND2_X1 U740 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U741 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U742 ( .A1(n1011), .A2(n1039), .ZN(n1032) );
NAND2_X1 U743 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U744 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
INV_X1 U745 ( .A(n1007), .ZN(n1016) );
NOR3_X1 U746 ( .A1(n1044), .A2(G953), .A3(n1045), .ZN(n999) );
INV_X1 U747 ( .A(n1014), .ZN(n1045) );
NAND4_X1 U748 ( .A1(n1046), .A2(n1012), .A3(n1047), .A4(n1048), .ZN(n1014) );
NOR4_X1 U749 ( .A1(n1042), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1048) );
XOR2_X1 U750 ( .A(n1052), .B(G478), .Z(n1050) );
NAND2_X1 U751 ( .A1(n1053), .A2(KEYINPUT26), .ZN(n1052) );
XOR2_X1 U752 ( .A(n1054), .B(KEYINPUT8), .Z(n1053) );
XOR2_X1 U753 ( .A(n1055), .B(n1056), .Z(n1049) );
XNOR2_X1 U754 ( .A(KEYINPUT18), .B(n1057), .ZN(n1056) );
XNOR2_X1 U755 ( .A(n1058), .B(n1059), .ZN(n1047) );
XOR2_X1 U756 ( .A(n1060), .B(KEYINPUT20), .Z(n1046) );
XOR2_X1 U757 ( .A(KEYINPUT17), .B(G952), .Z(n1044) );
NAND2_X1 U758 ( .A1(n1061), .A2(n1062), .ZN(G72) );
NAND2_X1 U759 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U760 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NAND2_X1 U761 ( .A1(KEYINPUT39), .A2(KEYINPUT6), .ZN(n1066) );
OR3_X1 U762 ( .A1(n1067), .A2(KEYINPUT39), .A3(n1064), .ZN(n1061) );
NAND2_X1 U763 ( .A1(G953), .A2(n1068), .ZN(n1064) );
NAND2_X1 U764 ( .A1(G900), .A2(G227), .ZN(n1068) );
XOR2_X1 U765 ( .A(KEYINPUT6), .B(n1065), .Z(n1067) );
XOR2_X1 U766 ( .A(n1069), .B(n1070), .Z(n1065) );
NOR2_X1 U767 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XOR2_X1 U768 ( .A(n1073), .B(n1074), .Z(n1072) );
XOR2_X1 U769 ( .A(n1075), .B(n1076), .Z(n1074) );
XOR2_X1 U770 ( .A(n1077), .B(n1078), .Z(n1073) );
XNOR2_X1 U771 ( .A(KEYINPUT33), .B(n1079), .ZN(n1077) );
NOR2_X1 U772 ( .A1(KEYINPUT7), .A2(n1080), .ZN(n1079) );
NOR2_X1 U773 ( .A1(G900), .A2(n1015), .ZN(n1071) );
NAND2_X1 U774 ( .A1(n1015), .A2(n1003), .ZN(n1069) );
XOR2_X1 U775 ( .A(n1081), .B(n1082), .Z(G69) );
XOR2_X1 U776 ( .A(n1083), .B(n1084), .Z(n1082) );
OR2_X1 U777 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U778 ( .A1(G953), .A2(n1087), .ZN(n1083) );
NAND2_X1 U779 ( .A1(G898), .A2(G224), .ZN(n1087) );
AND2_X1 U780 ( .A1(n1004), .A2(n1015), .ZN(n1081) );
NOR2_X1 U781 ( .A1(n1088), .A2(n1089), .ZN(G66) );
NOR3_X1 U782 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
NOR3_X1 U783 ( .A1(n1093), .A2(n1057), .A3(n1094), .ZN(n1092) );
NOR2_X1 U784 ( .A1(n1095), .A2(n1096), .ZN(n1091) );
NOR2_X1 U785 ( .A1(n1097), .A2(n1057), .ZN(n1095) );
NOR2_X1 U786 ( .A1(n1003), .A2(n1004), .ZN(n1097) );
NOR2_X1 U787 ( .A1(n1088), .A2(n1098), .ZN(G63) );
XOR2_X1 U788 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XNOR2_X1 U790 ( .A(KEYINPUT52), .B(KEYINPUT32), .ZN(n1102) );
XOR2_X1 U791 ( .A(n1103), .B(n1104), .Z(n1101) );
NAND2_X1 U792 ( .A1(n1105), .A2(G478), .ZN(n1099) );
NOR2_X1 U793 ( .A1(n1088), .A2(n1106), .ZN(G60) );
XOR2_X1 U794 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U795 ( .A(n1109), .B(KEYINPUT44), .Z(n1107) );
NAND2_X1 U796 ( .A1(n1105), .A2(G475), .ZN(n1109) );
XNOR2_X1 U797 ( .A(n1110), .B(n1111), .ZN(G6) );
NAND2_X1 U798 ( .A1(KEYINPUT42), .A2(n1112), .ZN(n1110) );
NOR2_X1 U799 ( .A1(n1088), .A2(n1113), .ZN(G57) );
XOR2_X1 U800 ( .A(n1114), .B(n1115), .Z(n1113) );
XNOR2_X1 U801 ( .A(n1116), .B(n1117), .ZN(n1115) );
NAND2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
XOR2_X1 U803 ( .A(n1120), .B(KEYINPUT63), .Z(n1118) );
XOR2_X1 U804 ( .A(n1121), .B(n1122), .Z(n1114) );
XOR2_X1 U805 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND3_X1 U806 ( .A1(n1105), .A2(G472), .A3(KEYINPUT23), .ZN(n1124) );
INV_X1 U807 ( .A(G101), .ZN(n1123) );
NAND2_X1 U808 ( .A1(n1125), .A2(KEYINPUT54), .ZN(n1121) );
XOR2_X1 U809 ( .A(n1126), .B(KEYINPUT29), .Z(n1125) );
NOR2_X1 U810 ( .A1(n1088), .A2(n1127), .ZN(G54) );
XOR2_X1 U811 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1129) );
XNOR2_X1 U813 ( .A(n1132), .B(n1133), .ZN(n1131) );
NAND2_X1 U814 ( .A1(KEYINPUT19), .A2(n1134), .ZN(n1132) );
XOR2_X1 U815 ( .A(n1135), .B(n1136), .Z(n1128) );
NOR2_X1 U816 ( .A1(KEYINPUT48), .A2(n1137), .ZN(n1136) );
XOR2_X1 U817 ( .A(n1138), .B(n1139), .Z(n1135) );
NAND2_X1 U818 ( .A1(n1105), .A2(G469), .ZN(n1138) );
INV_X1 U819 ( .A(n1094), .ZN(n1105) );
NOR2_X1 U820 ( .A1(n1140), .A2(n1141), .ZN(G51) );
XOR2_X1 U821 ( .A(KEYINPUT43), .B(n1088), .Z(n1141) );
NOR2_X1 U822 ( .A1(n1015), .A2(G952), .ZN(n1088) );
XOR2_X1 U823 ( .A(n1142), .B(n1143), .Z(n1140) );
XOR2_X1 U824 ( .A(n1144), .B(n1085), .Z(n1143) );
XOR2_X1 U825 ( .A(n1145), .B(n1146), .Z(n1142) );
NOR3_X1 U826 ( .A1(n1094), .A2(KEYINPUT50), .A3(n1058), .ZN(n1146) );
NAND2_X1 U827 ( .A1(G902), .A2(n1147), .ZN(n1094) );
OR2_X1 U828 ( .A1(n1004), .A2(n1003), .ZN(n1147) );
NAND4_X1 U829 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1003) );
NOR3_X1 U830 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
NAND2_X1 U831 ( .A1(n1155), .A2(n1156), .ZN(n1150) );
NAND2_X1 U832 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND2_X1 U833 ( .A1(n1159), .A2(n1010), .ZN(n1158) );
NAND2_X1 U834 ( .A1(n1009), .A2(n1160), .ZN(n1148) );
NAND2_X1 U835 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XOR2_X1 U836 ( .A(KEYINPUT0), .B(n1163), .Z(n1162) );
XOR2_X1 U837 ( .A(n1164), .B(KEYINPUT1), .Z(n1161) );
NAND4_X1 U838 ( .A1(n1111), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1004) );
AND4_X1 U839 ( .A1(n998), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1167) );
NAND3_X1 U840 ( .A1(n1010), .A2(n1011), .A3(n1171), .ZN(n998) );
NAND3_X1 U841 ( .A1(n1172), .A2(n1173), .A3(n1012), .ZN(n1166) );
NAND2_X1 U842 ( .A1(n1174), .A2(n1175), .ZN(n1172) );
NAND3_X1 U843 ( .A1(n1010), .A2(n1176), .A3(n1177), .ZN(n1175) );
XOR2_X1 U844 ( .A(KEYINPUT14), .B(n1155), .Z(n1176) );
NAND2_X1 U845 ( .A1(n1178), .A2(n1011), .ZN(n1174) );
NAND3_X1 U846 ( .A1(n1171), .A2(n1011), .A3(n1030), .ZN(n1111) );
XOR2_X1 U847 ( .A(G125), .B(n1179), .Z(n1145) );
XOR2_X1 U848 ( .A(n1180), .B(n1149), .Z(G48) );
NAND3_X1 U849 ( .A1(n1030), .A2(n1155), .A3(n1159), .ZN(n1149) );
XOR2_X1 U850 ( .A(G143), .B(n1152), .Z(G45) );
AND2_X1 U851 ( .A1(n1181), .A2(n1178), .ZN(n1152) );
NOR3_X1 U852 ( .A1(n1040), .A2(n1182), .A3(n1183), .ZN(n1178) );
XOR2_X1 U853 ( .A(n1184), .B(n1185), .Z(G42) );
XOR2_X1 U854 ( .A(KEYINPUT40), .B(G140), .Z(n1185) );
NOR3_X1 U855 ( .A1(n1164), .A2(KEYINPUT28), .A3(n1186), .ZN(n1184) );
NAND2_X1 U856 ( .A1(n1187), .A2(n1029), .ZN(n1164) );
XNOR2_X1 U857 ( .A(G137), .B(n1188), .ZN(G39) );
NAND2_X1 U858 ( .A1(n1163), .A2(n1009), .ZN(n1188) );
AND2_X1 U859 ( .A1(n1159), .A2(n1023), .ZN(n1163) );
INV_X1 U860 ( .A(n1189), .ZN(n1159) );
XOR2_X1 U861 ( .A(G134), .B(n1154), .Z(G36) );
AND3_X1 U862 ( .A1(n1009), .A2(n1010), .A3(n1181), .ZN(n1154) );
INV_X1 U863 ( .A(n1190), .ZN(n1010) );
XOR2_X1 U864 ( .A(G131), .B(n1153), .Z(G33) );
AND3_X1 U865 ( .A1(n1009), .A2(n1030), .A3(n1181), .ZN(n1153) );
AND3_X1 U866 ( .A1(n1029), .A2(n1191), .A3(n1177), .ZN(n1181) );
INV_X1 U867 ( .A(n1186), .ZN(n1009) );
NAND2_X1 U868 ( .A1(n1043), .A2(n1192), .ZN(n1186) );
XOR2_X1 U869 ( .A(G128), .B(n1193), .Z(G30) );
NOR3_X1 U870 ( .A1(n1194), .A2(n1190), .A3(n1189), .ZN(n1193) );
NAND4_X1 U871 ( .A1(n1037), .A2(n1029), .A3(n1051), .A4(n1191), .ZN(n1189) );
XOR2_X1 U872 ( .A(KEYINPUT13), .B(n1155), .Z(n1194) );
XOR2_X1 U873 ( .A(n1165), .B(n1195), .Z(G3) );
XOR2_X1 U874 ( .A(KEYINPUT35), .B(G101), .Z(n1195) );
NAND3_X1 U875 ( .A1(n1023), .A2(n1171), .A3(n1177), .ZN(n1165) );
XOR2_X1 U876 ( .A(G125), .B(n1196), .Z(G27) );
NOR2_X1 U877 ( .A1(n1040), .A2(n1197), .ZN(n1196) );
XNOR2_X1 U878 ( .A(KEYINPUT21), .B(n1157), .ZN(n1197) );
NAND2_X1 U879 ( .A1(n1187), .A2(n1012), .ZN(n1157) );
AND4_X1 U880 ( .A1(n1037), .A2(n1030), .A3(n1038), .A4(n1191), .ZN(n1187) );
NAND2_X1 U881 ( .A1(n1007), .A2(n1198), .ZN(n1191) );
NAND4_X1 U882 ( .A1(G953), .A2(G902), .A3(n1199), .A4(n1200), .ZN(n1198) );
INV_X1 U883 ( .A(G900), .ZN(n1200) );
XOR2_X1 U884 ( .A(n1201), .B(n1202), .Z(G24) );
XOR2_X1 U885 ( .A(KEYINPUT2), .B(G122), .Z(n1202) );
NAND4_X1 U886 ( .A1(n1060), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
XOR2_X1 U887 ( .A(KEYINPUT27), .B(n1011), .Z(n1204) );
NOR2_X1 U888 ( .A1(n1051), .A2(n1206), .ZN(n1011) );
XOR2_X1 U889 ( .A(n1170), .B(n1207), .Z(G21) );
XOR2_X1 U890 ( .A(KEYINPUT45), .B(G119), .Z(n1207) );
NAND4_X1 U891 ( .A1(n1203), .A2(n1023), .A3(n1037), .A4(n1051), .ZN(n1170) );
XOR2_X1 U892 ( .A(n1208), .B(n1209), .Z(G18) );
NAND4_X1 U893 ( .A1(n1210), .A2(n1177), .A3(n1211), .A4(n1012), .ZN(n1209) );
NOR2_X1 U894 ( .A1(n1040), .A2(n1190), .ZN(n1211) );
NAND2_X1 U895 ( .A1(n1183), .A2(n1205), .ZN(n1190) );
INV_X1 U896 ( .A(n1155), .ZN(n1040) );
XOR2_X1 U897 ( .A(n1173), .B(KEYINPUT4), .Z(n1210) );
NAND2_X1 U898 ( .A1(n1212), .A2(n1213), .ZN(G15) );
OR2_X1 U899 ( .A1(n1169), .A2(G113), .ZN(n1213) );
XOR2_X1 U900 ( .A(n1214), .B(KEYINPUT55), .Z(n1212) );
NAND2_X1 U901 ( .A1(G113), .A2(n1169), .ZN(n1214) );
NAND3_X1 U902 ( .A1(n1177), .A2(n1203), .A3(n1030), .ZN(n1169) );
NOR2_X1 U903 ( .A1(n1205), .A2(n1183), .ZN(n1030) );
INV_X1 U904 ( .A(n1060), .ZN(n1183) );
AND3_X1 U905 ( .A1(n1155), .A2(n1173), .A3(n1012), .ZN(n1203) );
NOR2_X1 U906 ( .A1(n1215), .A2(n1027), .ZN(n1012) );
INV_X1 U907 ( .A(n1028), .ZN(n1215) );
INV_X1 U908 ( .A(n1035), .ZN(n1177) );
NAND2_X1 U909 ( .A1(n1051), .A2(n1216), .ZN(n1035) );
INV_X1 U910 ( .A(n1206), .ZN(n1216) );
INV_X1 U911 ( .A(n1038), .ZN(n1051) );
XOR2_X1 U912 ( .A(n1217), .B(G110), .Z(G12) );
NAND2_X1 U913 ( .A1(KEYINPUT46), .A2(n1168), .ZN(n1217) );
NAND4_X1 U914 ( .A1(n1037), .A2(n1023), .A3(n1038), .A4(n1171), .ZN(n1168) );
AND3_X1 U915 ( .A1(n1029), .A2(n1173), .A3(n1155), .ZN(n1171) );
NOR2_X1 U916 ( .A1(n1043), .A2(n1042), .ZN(n1155) );
INV_X1 U917 ( .A(n1192), .ZN(n1042) );
NAND2_X1 U918 ( .A1(G214), .A2(n1218), .ZN(n1192) );
XNOR2_X1 U919 ( .A(n1059), .B(n1219), .ZN(n1043) );
NOR2_X1 U920 ( .A1(KEYINPUT62), .A2(n1220), .ZN(n1219) );
XOR2_X1 U921 ( .A(n1058), .B(KEYINPUT47), .Z(n1220) );
NAND2_X1 U922 ( .A1(G210), .A2(n1218), .ZN(n1058) );
NAND2_X1 U923 ( .A1(n1221), .A2(n1222), .ZN(n1218) );
INV_X1 U924 ( .A(G237), .ZN(n1221) );
NAND2_X1 U925 ( .A1(n1223), .A2(n1224), .ZN(n1059) );
XNOR2_X1 U926 ( .A(n1225), .B(n1085), .ZN(n1224) );
XOR2_X1 U927 ( .A(n1226), .B(n1227), .Z(n1085) );
XOR2_X1 U928 ( .A(n1228), .B(n1229), .Z(n1227) );
XOR2_X1 U929 ( .A(n1230), .B(n1231), .Z(n1226) );
XOR2_X1 U930 ( .A(G110), .B(G101), .Z(n1231) );
NAND2_X1 U931 ( .A1(n1232), .A2(n1233), .ZN(n1230) );
NAND2_X1 U932 ( .A1(G107), .A2(n1112), .ZN(n1233) );
XOR2_X1 U933 ( .A(KEYINPUT51), .B(n1234), .Z(n1232) );
NOR2_X1 U934 ( .A1(G107), .A2(n1112), .ZN(n1234) );
NOR2_X1 U935 ( .A1(n1235), .A2(n1236), .ZN(n1225) );
XOR2_X1 U936 ( .A(n1237), .B(KEYINPUT41), .Z(n1236) );
NAND2_X1 U937 ( .A1(n1238), .A2(n1179), .ZN(n1237) );
NOR2_X1 U938 ( .A1(n1179), .A2(n1238), .ZN(n1235) );
NAND2_X1 U939 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
NAND2_X1 U940 ( .A1(G125), .A2(n1241), .ZN(n1240) );
INV_X1 U941 ( .A(n1144), .ZN(n1241) );
XOR2_X1 U942 ( .A(n1242), .B(KEYINPUT22), .Z(n1239) );
NAND2_X1 U943 ( .A1(n1144), .A2(n1243), .ZN(n1242) );
INV_X1 U944 ( .A(G125), .ZN(n1243) );
NAND2_X1 U945 ( .A1(G224), .A2(n1015), .ZN(n1179) );
XOR2_X1 U946 ( .A(n1222), .B(KEYINPUT3), .Z(n1223) );
NAND2_X1 U947 ( .A1(n1007), .A2(n1244), .ZN(n1173) );
NAND3_X1 U948 ( .A1(G902), .A2(n1199), .A3(n1086), .ZN(n1244) );
NOR2_X1 U949 ( .A1(n1015), .A2(G898), .ZN(n1086) );
NAND3_X1 U950 ( .A1(n1199), .A2(n1015), .A3(G952), .ZN(n1007) );
NAND2_X1 U951 ( .A1(G237), .A2(G234), .ZN(n1199) );
NOR2_X1 U952 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
AND2_X1 U953 ( .A1(G221), .A2(n1245), .ZN(n1027) );
XOR2_X1 U954 ( .A(n1246), .B(G469), .Z(n1028) );
NAND2_X1 U955 ( .A1(n1247), .A2(n1222), .ZN(n1246) );
XOR2_X1 U956 ( .A(n1248), .B(n1249), .Z(n1247) );
XNOR2_X1 U957 ( .A(n1134), .B(n1137), .ZN(n1249) );
XOR2_X1 U958 ( .A(G140), .B(G110), .Z(n1137) );
XOR2_X1 U959 ( .A(n1250), .B(n1139), .Z(n1248) );
AND2_X1 U960 ( .A1(G227), .A2(n1015), .ZN(n1139) );
NAND3_X1 U961 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1250) );
NAND2_X1 U962 ( .A1(n1130), .A2(n1254), .ZN(n1253) );
NAND2_X1 U963 ( .A1(n1255), .A2(KEYINPUT12), .ZN(n1254) );
XNOR2_X1 U964 ( .A(n1133), .B(KEYINPUT37), .ZN(n1255) );
INV_X1 U965 ( .A(n1076), .ZN(n1130) );
NAND3_X1 U966 ( .A1(KEYINPUT12), .A2(n1076), .A3(n1133), .ZN(n1252) );
XOR2_X1 U967 ( .A(n1256), .B(n1257), .Z(n1076) );
XOR2_X1 U968 ( .A(G143), .B(n1180), .Z(n1256) );
OR2_X1 U969 ( .A1(n1133), .A2(KEYINPUT12), .ZN(n1251) );
XNOR2_X1 U970 ( .A(n1258), .B(G101), .ZN(n1133) );
NAND2_X1 U971 ( .A1(n1259), .A2(KEYINPUT10), .ZN(n1258) );
XOR2_X1 U972 ( .A(n1260), .B(G107), .Z(n1259) );
NAND2_X1 U973 ( .A1(KEYINPUT58), .A2(n1112), .ZN(n1260) );
INV_X1 U974 ( .A(G104), .ZN(n1112) );
XOR2_X1 U975 ( .A(n1261), .B(G472), .Z(n1038) );
NAND2_X1 U976 ( .A1(n1262), .A2(n1222), .ZN(n1261) );
XNOR2_X1 U977 ( .A(n1126), .B(n1263), .ZN(n1262) );
XOR2_X1 U978 ( .A(G101), .B(n1264), .Z(n1263) );
NOR2_X1 U979 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
XOR2_X1 U980 ( .A(n1267), .B(KEYINPUT11), .Z(n1266) );
NAND3_X1 U981 ( .A1(n1119), .A2(n1120), .A3(n1117), .ZN(n1267) );
NOR2_X1 U982 ( .A1(n1268), .A2(n1117), .ZN(n1265) );
XNOR2_X1 U983 ( .A(n1269), .B(n1228), .ZN(n1117) );
XOR2_X1 U984 ( .A(G116), .B(G119), .Z(n1228) );
XNOR2_X1 U985 ( .A(G113), .B(KEYINPUT36), .ZN(n1269) );
AND2_X1 U986 ( .A1(n1120), .A2(n1119), .ZN(n1268) );
OR2_X1 U987 ( .A1(n1134), .A2(n1144), .ZN(n1119) );
NAND2_X1 U988 ( .A1(n1134), .A2(n1144), .ZN(n1120) );
XOR2_X1 U989 ( .A(n1270), .B(n1257), .Z(n1144) );
XOR2_X1 U990 ( .A(G128), .B(KEYINPUT53), .Z(n1257) );
NAND3_X1 U991 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1270) );
NAND2_X1 U992 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
OR3_X1 U993 ( .A1(n1275), .A2(n1274), .A3(n1276), .ZN(n1272) );
XOR2_X1 U994 ( .A(G143), .B(KEYINPUT60), .Z(n1274) );
NAND2_X1 U995 ( .A1(KEYINPUT38), .A2(n1180), .ZN(n1275) );
INV_X1 U996 ( .A(G146), .ZN(n1180) );
NAND2_X1 U997 ( .A1(G146), .A2(n1276), .ZN(n1271) );
INV_X1 U998 ( .A(KEYINPUT30), .ZN(n1276) );
XOR2_X1 U999 ( .A(n1080), .B(n1075), .Z(n1134) );
XOR2_X1 U1000 ( .A(G134), .B(G137), .Z(n1075) );
NAND2_X1 U1001 ( .A1(n1277), .A2(G210), .ZN(n1126) );
NOR2_X1 U1002 ( .A1(n1205), .A2(n1060), .ZN(n1023) );
XOR2_X1 U1003 ( .A(n1278), .B(n1279), .Z(n1060) );
XOR2_X1 U1004 ( .A(KEYINPUT31), .B(G475), .Z(n1279) );
OR2_X1 U1005 ( .A1(n1108), .A2(G902), .ZN(n1278) );
XNOR2_X1 U1006 ( .A(n1280), .B(n1281), .ZN(n1108) );
XNOR2_X1 U1007 ( .A(n1229), .B(n1282), .ZN(n1281) );
XOR2_X1 U1008 ( .A(n1283), .B(n1284), .Z(n1282) );
INV_X1 U1009 ( .A(n1080), .ZN(n1284) );
XNOR2_X1 U1010 ( .A(G131), .B(KEYINPUT57), .ZN(n1080) );
NAND2_X1 U1011 ( .A1(n1277), .A2(G214), .ZN(n1283) );
NOR2_X1 U1012 ( .A1(G953), .A2(G237), .ZN(n1277) );
XOR2_X1 U1013 ( .A(G122), .B(G113), .Z(n1229) );
XOR2_X1 U1014 ( .A(n1285), .B(n1286), .Z(n1280) );
XOR2_X1 U1015 ( .A(G143), .B(G104), .Z(n1286) );
NAND2_X1 U1016 ( .A1(n1287), .A2(n1288), .ZN(n1285) );
NAND2_X1 U1017 ( .A1(G146), .A2(n1078), .ZN(n1288) );
XOR2_X1 U1018 ( .A(KEYINPUT61), .B(n1289), .Z(n1287) );
NOR2_X1 U1019 ( .A1(G146), .A2(n1290), .ZN(n1289) );
XNOR2_X1 U1020 ( .A(n1078), .B(KEYINPUT25), .ZN(n1290) );
INV_X1 U1021 ( .A(n1182), .ZN(n1205) );
XOR2_X1 U1022 ( .A(n1054), .B(G478), .Z(n1182) );
NAND2_X1 U1023 ( .A1(n1291), .A2(n1222), .ZN(n1054) );
XOR2_X1 U1024 ( .A(n1292), .B(n1104), .Z(n1291) );
XNOR2_X1 U1025 ( .A(n1293), .B(n1294), .ZN(n1104) );
XOR2_X1 U1026 ( .A(G107), .B(n1295), .Z(n1294) );
NOR2_X1 U1027 ( .A1(KEYINPUT34), .A2(n1296), .ZN(n1295) );
XOR2_X1 U1028 ( .A(n1208), .B(G122), .Z(n1296) );
INV_X1 U1029 ( .A(G116), .ZN(n1208) );
NAND2_X1 U1030 ( .A1(G217), .A2(n1297), .ZN(n1293) );
INV_X1 U1031 ( .A(n1103), .ZN(n1292) );
XNOR2_X1 U1032 ( .A(G128), .B(n1298), .ZN(n1103) );
XOR2_X1 U1033 ( .A(G143), .B(G134), .Z(n1298) );
XOR2_X1 U1034 ( .A(n1206), .B(KEYINPUT5), .Z(n1037) );
XOR2_X1 U1035 ( .A(n1299), .B(n1090), .Z(n1206) );
INV_X1 U1036 ( .A(n1055), .ZN(n1090) );
NAND2_X1 U1037 ( .A1(n1093), .A2(n1222), .ZN(n1055) );
INV_X1 U1038 ( .A(n1096), .ZN(n1093) );
XOR2_X1 U1039 ( .A(n1300), .B(n1301), .Z(n1096) );
XOR2_X1 U1040 ( .A(KEYINPUT24), .B(G137), .Z(n1301) );
XOR2_X1 U1041 ( .A(n1302), .B(n1303), .Z(n1300) );
AND2_X1 U1042 ( .A1(G221), .A2(n1297), .ZN(n1303) );
AND2_X1 U1043 ( .A1(G234), .A2(n1015), .ZN(n1297) );
INV_X1 U1044 ( .A(G953), .ZN(n1015) );
NAND2_X1 U1045 ( .A1(n1304), .A2(n1305), .ZN(n1302) );
NAND2_X1 U1046 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XOR2_X1 U1047 ( .A(KEYINPUT16), .B(n1308), .Z(n1304) );
NOR2_X1 U1048 ( .A1(n1306), .A2(n1307), .ZN(n1308) );
XOR2_X1 U1049 ( .A(G110), .B(n1309), .Z(n1307) );
XOR2_X1 U1050 ( .A(G128), .B(G119), .Z(n1309) );
XOR2_X1 U1051 ( .A(n1078), .B(n1310), .Z(n1306) );
NOR2_X1 U1052 ( .A1(G146), .A2(KEYINPUT59), .ZN(n1310) );
XOR2_X1 U1053 ( .A(G140), .B(G125), .Z(n1078) );
NAND2_X1 U1054 ( .A1(KEYINPUT49), .A2(n1311), .ZN(n1299) );
XNOR2_X1 U1055 ( .A(KEYINPUT56), .B(n1057), .ZN(n1311) );
NAND2_X1 U1056 ( .A1(G217), .A2(n1245), .ZN(n1057) );
NAND2_X1 U1057 ( .A1(G234), .A2(n1222), .ZN(n1245) );
INV_X1 U1058 ( .A(G902), .ZN(n1222) );
endmodule


