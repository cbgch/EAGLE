//Key = 0010011000100011110100001110011111011101110001000100100010000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397;

XOR2_X1 U759 ( .A(G107), .B(n1055), .Z(G9) );
NOR4_X1 U760 ( .A1(KEYINPUT58), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1055) );
NOR2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(G75) );
NOR3_X1 U762 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NAND3_X1 U763 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1061) );
NAND2_X1 U764 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U765 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND4_X1 U766 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1070) );
NAND2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NAND2_X1 U768 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U769 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
OR2_X1 U770 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
INV_X1 U771 ( .A(n1083), .ZN(n1079) );
NAND2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1075) );
NAND2_X1 U773 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U774 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
INV_X1 U775 ( .A(n1090), .ZN(n1088) );
NAND3_X1 U776 ( .A1(n1091), .A2(n1092), .A3(n1077), .ZN(n1069) );
NAND2_X1 U777 ( .A1(n1093), .A2(n1057), .ZN(n1092) );
INV_X1 U778 ( .A(n1084), .ZN(n1057) );
OR3_X1 U779 ( .A1(n1094), .A2(KEYINPUT17), .A3(n1095), .ZN(n1093) );
NAND3_X1 U780 ( .A1(n1096), .A2(n1097), .A3(n1084), .ZN(n1091) );
NAND3_X1 U781 ( .A1(n1072), .A2(n1098), .A3(KEYINPUT17), .ZN(n1097) );
NAND3_X1 U782 ( .A1(n1099), .A2(n1100), .A3(n1071), .ZN(n1096) );
NAND2_X1 U783 ( .A1(n1101), .A2(n1095), .ZN(n1100) );
NAND3_X1 U784 ( .A1(n1058), .A2(n1102), .A3(n1074), .ZN(n1099) );
INV_X1 U785 ( .A(n1103), .ZN(n1067) );
NOR3_X1 U786 ( .A1(n1104), .A2(G953), .A3(G952), .ZN(n1059) );
INV_X1 U787 ( .A(n1064), .ZN(n1104) );
NAND4_X1 U788 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1064) );
NOR3_X1 U789 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1108) );
NOR2_X1 U790 ( .A1(KEYINPUT37), .A2(n1112), .ZN(n1110) );
NAND3_X1 U791 ( .A1(n1074), .A2(n1090), .A3(n1113), .ZN(n1109) );
XOR2_X1 U792 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U793 ( .A(n1116), .B(KEYINPUT59), .Z(n1115) );
NAND2_X1 U794 ( .A1(KEYINPUT52), .A2(n1117), .ZN(n1114) );
NOR3_X1 U795 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1107) );
NOR2_X1 U796 ( .A1(G475), .A2(n1121), .ZN(n1120) );
NOR2_X1 U797 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XOR2_X1 U798 ( .A(KEYINPUT27), .B(n1124), .Z(n1123) );
NOR3_X1 U799 ( .A1(n1125), .A2(n1124), .A3(n1122), .ZN(n1119) );
INV_X1 U800 ( .A(KEYINPUT37), .ZN(n1122) );
XOR2_X1 U801 ( .A(n1126), .B(n1127), .Z(n1118) );
XOR2_X1 U802 ( .A(n1128), .B(G472), .Z(n1105) );
XOR2_X1 U803 ( .A(n1129), .B(n1130), .Z(G72) );
NOR2_X1 U804 ( .A1(n1131), .A2(n1065), .ZN(n1130) );
AND2_X1 U805 ( .A1(G227), .A2(G900), .ZN(n1131) );
XOR2_X1 U806 ( .A(n1132), .B(n1133), .Z(n1129) );
NOR2_X1 U807 ( .A1(n1134), .A2(KEYINPUT44), .ZN(n1133) );
AND2_X1 U808 ( .A1(n1065), .A2(n1063), .ZN(n1134) );
NAND2_X1 U809 ( .A1(n1135), .A2(n1136), .ZN(n1132) );
NAND2_X1 U810 ( .A1(G953), .A2(n1137), .ZN(n1136) );
XOR2_X1 U811 ( .A(n1138), .B(n1139), .Z(n1135) );
XOR2_X1 U812 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U813 ( .A(n1142), .B(n1143), .Z(n1138) );
NAND2_X1 U814 ( .A1(n1144), .A2(n1145), .ZN(G69) );
NAND2_X1 U815 ( .A1(n1146), .A2(n1065), .ZN(n1145) );
XNOR2_X1 U816 ( .A(n1062), .B(n1147), .ZN(n1146) );
NAND2_X1 U817 ( .A1(n1148), .A2(G953), .ZN(n1144) );
NAND2_X1 U818 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NAND2_X1 U819 ( .A1(n1147), .A2(n1151), .ZN(n1150) );
INV_X1 U820 ( .A(G224), .ZN(n1151) );
NAND2_X1 U821 ( .A1(G224), .A2(n1152), .ZN(n1149) );
NAND2_X1 U822 ( .A1(G898), .A2(n1147), .ZN(n1152) );
NAND2_X1 U823 ( .A1(n1153), .A2(n1154), .ZN(n1147) );
NAND2_X1 U824 ( .A1(G953), .A2(n1155), .ZN(n1154) );
XOR2_X1 U825 ( .A(n1156), .B(n1157), .Z(n1153) );
XOR2_X1 U826 ( .A(KEYINPUT41), .B(n1158), .Z(n1157) );
NOR2_X1 U827 ( .A1(n1159), .A2(n1160), .ZN(G66) );
XNOR2_X1 U828 ( .A(n1161), .B(n1162), .ZN(n1160) );
NOR2_X1 U829 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U830 ( .A1(n1159), .A2(n1165), .ZN(G63) );
XOR2_X1 U831 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U832 ( .A1(n1168), .A2(n1164), .ZN(n1167) );
INV_X1 U833 ( .A(G478), .ZN(n1168) );
NAND2_X1 U834 ( .A1(KEYINPUT6), .A2(n1169), .ZN(n1166) );
NOR2_X1 U835 ( .A1(n1159), .A2(n1170), .ZN(G60) );
XOR2_X1 U836 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U837 ( .A1(KEYINPUT13), .A2(n1173), .ZN(n1172) );
OR2_X1 U838 ( .A1(n1164), .A2(n1125), .ZN(n1171) );
XNOR2_X1 U839 ( .A(G104), .B(n1174), .ZN(G6) );
NOR3_X1 U840 ( .A1(n1159), .A2(n1175), .A3(n1176), .ZN(G57) );
NOR3_X1 U841 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1176) );
NOR2_X1 U842 ( .A1(KEYINPUT28), .A2(n1180), .ZN(n1178) );
INV_X1 U843 ( .A(KEYINPUT3), .ZN(n1180) );
NOR2_X1 U844 ( .A1(n1181), .A2(n1182), .ZN(n1175) );
NOR2_X1 U845 ( .A1(KEYINPUT3), .A2(n1183), .ZN(n1181) );
XOR2_X1 U846 ( .A(KEYINPUT28), .B(n1179), .Z(n1183) );
XNOR2_X1 U847 ( .A(n1184), .B(n1185), .ZN(n1179) );
NOR2_X1 U848 ( .A1(n1186), .A2(n1164), .ZN(n1185) );
INV_X1 U849 ( .A(G472), .ZN(n1186) );
NOR2_X1 U850 ( .A1(n1159), .A2(n1187), .ZN(G54) );
XOR2_X1 U851 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U852 ( .A(n1190), .B(n1191), .Z(n1189) );
XOR2_X1 U853 ( .A(n1192), .B(n1193), .Z(n1190) );
NAND3_X1 U854 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1192) );
OR2_X1 U855 ( .A1(n1197), .A2(KEYINPUT5), .ZN(n1196) );
NAND3_X1 U856 ( .A1(KEYINPUT5), .A2(n1197), .A3(n1198), .ZN(n1195) );
NAND2_X1 U857 ( .A1(n1143), .A2(n1199), .ZN(n1194) );
NAND2_X1 U858 ( .A1(KEYINPUT5), .A2(n1200), .ZN(n1199) );
XOR2_X1 U859 ( .A(KEYINPUT38), .B(n1197), .Z(n1200) );
XNOR2_X1 U860 ( .A(n1201), .B(KEYINPUT51), .ZN(n1197) );
XOR2_X1 U861 ( .A(n1202), .B(n1203), .Z(n1188) );
XOR2_X1 U862 ( .A(KEYINPUT20), .B(KEYINPUT12), .Z(n1203) );
XOR2_X1 U863 ( .A(n1204), .B(n1205), .Z(n1202) );
NOR2_X1 U864 ( .A1(n1116), .A2(n1164), .ZN(n1205) );
NOR2_X1 U865 ( .A1(n1159), .A2(n1206), .ZN(G51) );
XOR2_X1 U866 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR2_X1 U867 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NOR2_X1 U868 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NOR2_X1 U869 ( .A1(n1213), .A2(KEYINPUT1), .ZN(n1212) );
NOR2_X1 U870 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U871 ( .A(n1216), .B(KEYINPUT60), .Z(n1214) );
INV_X1 U872 ( .A(n1217), .ZN(n1211) );
NOR2_X1 U873 ( .A1(KEYINPUT1), .A2(n1217), .ZN(n1209) );
NAND2_X1 U874 ( .A1(n1215), .A2(n1216), .ZN(n1217) );
NAND3_X1 U875 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1216) );
NAND3_X1 U876 ( .A1(G125), .A2(n1221), .A3(n1222), .ZN(n1220) );
NAND2_X1 U877 ( .A1(n1223), .A2(n1224), .ZN(n1219) );
XOR2_X1 U878 ( .A(n1222), .B(n1221), .Z(n1223) );
NAND3_X1 U879 ( .A1(n1225), .A2(n1226), .A3(G125), .ZN(n1218) );
NOR2_X1 U880 ( .A1(n1126), .A2(n1164), .ZN(n1207) );
NAND2_X1 U881 ( .A1(G902), .A2(n1227), .ZN(n1164) );
OR2_X1 U882 ( .A1(n1063), .A2(n1062), .ZN(n1227) );
NAND4_X1 U883 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1062) );
AND4_X1 U884 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1174), .ZN(n1231) );
NAND3_X1 U885 ( .A1(n1084), .A2(n1235), .A3(n1236), .ZN(n1174) );
NOR2_X1 U886 ( .A1(n1237), .A2(n1238), .ZN(n1230) );
NOR2_X1 U887 ( .A1(KEYINPUT57), .A2(n1239), .ZN(n1238) );
NOR2_X1 U888 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
NOR2_X1 U889 ( .A1(n1242), .A2(n1243), .ZN(n1240) );
XOR2_X1 U890 ( .A(KEYINPUT34), .B(n1244), .Z(n1243) );
NOR2_X1 U891 ( .A1(n1102), .A2(n1245), .ZN(n1244) );
NOR3_X1 U892 ( .A1(n1246), .A2(n1095), .A3(n1247), .ZN(n1242) );
INV_X1 U893 ( .A(KEYINPUT57), .ZN(n1247) );
NAND3_X1 U894 ( .A1(n1248), .A2(n1094), .A3(n1083), .ZN(n1246) );
NAND3_X1 U895 ( .A1(n1084), .A2(n1235), .A3(n1249), .ZN(n1229) );
NAND2_X1 U896 ( .A1(n1250), .A2(n1251), .ZN(n1228) );
XOR2_X1 U897 ( .A(KEYINPUT43), .B(n1252), .Z(n1251) );
NAND2_X1 U898 ( .A1(n1253), .A2(n1254), .ZN(n1063) );
NOR4_X1 U899 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1254) );
INV_X1 U900 ( .A(n1259), .ZN(n1258) );
AND4_X1 U901 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(n1253) );
AND2_X1 U902 ( .A1(G953), .A2(n1264), .ZN(n1159) );
XOR2_X1 U903 ( .A(KEYINPUT31), .B(G952), .Z(n1264) );
NAND2_X1 U904 ( .A1(n1265), .A2(n1266), .ZN(G48) );
NAND2_X1 U905 ( .A1(G146), .A2(n1263), .ZN(n1266) );
XOR2_X1 U906 ( .A(KEYINPUT61), .B(n1267), .Z(n1265) );
NOR2_X1 U907 ( .A1(G146), .A2(n1263), .ZN(n1267) );
NAND4_X1 U908 ( .A1(n1236), .A2(n1268), .A3(n1082), .A4(n1250), .ZN(n1263) );
XOR2_X1 U909 ( .A(n1269), .B(n1262), .Z(G45) );
NAND4_X1 U910 ( .A1(n1098), .A2(n1250), .A3(n1083), .A4(n1270), .ZN(n1262) );
NOR3_X1 U911 ( .A1(n1106), .A2(n1271), .A3(n1272), .ZN(n1270) );
XOR2_X1 U912 ( .A(n1142), .B(n1261), .Z(G42) );
NAND4_X1 U913 ( .A1(n1236), .A2(n1077), .A3(n1268), .A4(n1273), .ZN(n1261) );
NAND3_X1 U914 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(G39) );
NAND2_X1 U915 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND3_X1 U916 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1278) );
NAND2_X1 U917 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U918 ( .A1(KEYINPUT7), .A2(G137), .ZN(n1280) );
NAND2_X1 U919 ( .A1(n1284), .A2(n1285), .ZN(n1279) );
INV_X1 U920 ( .A(KEYINPUT7), .ZN(n1285) );
NAND2_X1 U921 ( .A1(G137), .A2(n1286), .ZN(n1284) );
NAND2_X1 U922 ( .A1(KEYINPUT19), .A2(n1287), .ZN(n1286) );
INV_X1 U923 ( .A(n1260), .ZN(n1277) );
NAND4_X1 U924 ( .A1(n1282), .A2(n1260), .A3(G137), .A4(KEYINPUT19), .ZN(n1275) );
NAND2_X1 U925 ( .A1(n1288), .A2(n1283), .ZN(n1274) );
INV_X1 U926 ( .A(KEYINPUT19), .ZN(n1283) );
NAND2_X1 U927 ( .A1(G137), .A2(n1289), .ZN(n1288) );
NAND2_X1 U928 ( .A1(n1287), .A2(n1260), .ZN(n1289) );
NAND4_X1 U929 ( .A1(n1072), .A2(n1077), .A3(n1082), .A4(n1268), .ZN(n1260) );
INV_X1 U930 ( .A(n1282), .ZN(n1287) );
XNOR2_X1 U931 ( .A(KEYINPUT2), .B(KEYINPUT15), .ZN(n1282) );
XOR2_X1 U932 ( .A(G134), .B(n1257), .Z(G36) );
AND2_X1 U933 ( .A1(n1290), .A2(n1249), .ZN(n1257) );
XOR2_X1 U934 ( .A(G131), .B(n1256), .Z(G33) );
AND2_X1 U935 ( .A1(n1236), .A2(n1290), .ZN(n1256) );
AND4_X1 U936 ( .A1(n1083), .A2(n1077), .A3(n1098), .A4(n1291), .ZN(n1290) );
AND2_X1 U937 ( .A1(n1089), .A2(n1090), .ZN(n1077) );
XNOR2_X1 U938 ( .A(n1292), .B(KEYINPUT9), .ZN(n1089) );
XOR2_X1 U939 ( .A(G128), .B(n1255), .Z(G30) );
AND4_X1 U940 ( .A1(n1082), .A2(n1268), .A3(n1249), .A4(n1250), .ZN(n1255) );
INV_X1 U941 ( .A(n1058), .ZN(n1249) );
NOR3_X1 U942 ( .A1(n1081), .A2(n1272), .A3(n1094), .ZN(n1268) );
XOR2_X1 U943 ( .A(n1239), .B(n1293), .Z(G3) );
NAND2_X1 U944 ( .A1(KEYINPUT25), .A2(G101), .ZN(n1293) );
NAND3_X1 U945 ( .A1(n1083), .A2(n1235), .A3(n1072), .ZN(n1239) );
XOR2_X1 U946 ( .A(n1224), .B(n1259), .Z(G27) );
NAND3_X1 U947 ( .A1(n1294), .A2(n1236), .A3(n1295), .ZN(n1259) );
NOR3_X1 U948 ( .A1(n1081), .A2(n1272), .A3(n1082), .ZN(n1295) );
INV_X1 U949 ( .A(n1291), .ZN(n1272) );
NAND2_X1 U950 ( .A1(n1296), .A2(n1297), .ZN(n1291) );
NAND4_X1 U951 ( .A1(G953), .A2(G902), .A3(n1298), .A4(n1137), .ZN(n1297) );
INV_X1 U952 ( .A(G900), .ZN(n1137) );
XOR2_X1 U953 ( .A(n1103), .B(KEYINPUT47), .Z(n1296) );
INV_X1 U954 ( .A(n1102), .ZN(n1236) );
INV_X1 U955 ( .A(G125), .ZN(n1224) );
XNOR2_X1 U956 ( .A(G122), .B(n1234), .ZN(G24) );
NAND3_X1 U957 ( .A1(n1294), .A2(n1084), .A3(n1299), .ZN(n1234) );
NOR3_X1 U958 ( .A1(n1106), .A2(n1300), .A3(n1271), .ZN(n1299) );
NOR2_X1 U959 ( .A1(n1111), .A2(n1082), .ZN(n1084) );
XOR2_X1 U960 ( .A(n1233), .B(n1301), .Z(G21) );
NAND2_X1 U961 ( .A1(n1302), .A2(KEYINPUT26), .ZN(n1301) );
XOR2_X1 U962 ( .A(n1303), .B(KEYINPUT63), .Z(n1302) );
NAND3_X1 U963 ( .A1(n1072), .A2(n1294), .A3(n1304), .ZN(n1233) );
NOR3_X1 U964 ( .A1(n1273), .A2(n1300), .A3(n1081), .ZN(n1304) );
AND3_X1 U965 ( .A1(n1250), .A2(n1074), .A3(n1071), .ZN(n1294) );
INV_X1 U966 ( .A(n1095), .ZN(n1072) );
XNOR2_X1 U967 ( .A(G116), .B(n1305), .ZN(G18) );
NAND2_X1 U968 ( .A1(n1252), .A2(n1250), .ZN(n1305) );
INV_X1 U969 ( .A(n1086), .ZN(n1250) );
NOR2_X1 U970 ( .A1(n1245), .A2(n1058), .ZN(n1252) );
NAND2_X1 U971 ( .A1(n1271), .A2(n1306), .ZN(n1058) );
INV_X1 U972 ( .A(n1106), .ZN(n1306) );
XOR2_X1 U973 ( .A(n1307), .B(n1308), .Z(G15) );
NAND2_X1 U974 ( .A1(KEYINPUT16), .A2(G113), .ZN(n1308) );
OR3_X1 U975 ( .A1(n1241), .A2(n1309), .A3(n1245), .ZN(n1307) );
NAND4_X1 U976 ( .A1(n1071), .A2(n1083), .A3(n1074), .A4(n1248), .ZN(n1245) );
NOR2_X1 U977 ( .A1(n1273), .A2(n1111), .ZN(n1083) );
INV_X1 U978 ( .A(n1082), .ZN(n1273) );
XOR2_X1 U979 ( .A(KEYINPUT53), .B(n1102), .Z(n1309) );
NAND2_X1 U980 ( .A1(n1106), .A2(n1310), .ZN(n1102) );
XOR2_X1 U981 ( .A(n1232), .B(n1311), .Z(G12) );
NOR2_X1 U982 ( .A1(G110), .A2(KEYINPUT22), .ZN(n1311) );
OR4_X1 U983 ( .A1(n1095), .A2(n1056), .A3(n1081), .A4(n1082), .ZN(n1232) );
XNOR2_X1 U984 ( .A(n1312), .B(n1128), .ZN(n1082) );
NAND2_X1 U985 ( .A1(n1313), .A2(n1314), .ZN(n1128) );
XOR2_X1 U986 ( .A(n1184), .B(n1182), .Z(n1313) );
INV_X1 U987 ( .A(n1177), .ZN(n1182) );
XOR2_X1 U988 ( .A(n1315), .B(G101), .Z(n1177) );
NAND2_X1 U989 ( .A1(G210), .A2(n1316), .ZN(n1315) );
XOR2_X1 U990 ( .A(n1317), .B(n1318), .Z(n1184) );
XOR2_X1 U991 ( .A(G113), .B(n1319), .Z(n1318) );
NOR2_X1 U992 ( .A1(KEYINPUT46), .A2(n1320), .ZN(n1319) );
XOR2_X1 U993 ( .A(n1225), .B(n1191), .Z(n1317) );
NAND2_X1 U994 ( .A1(KEYINPUT49), .A2(n1321), .ZN(n1312) );
XOR2_X1 U995 ( .A(KEYINPUT24), .B(G472), .Z(n1321) );
XNOR2_X1 U996 ( .A(n1111), .B(KEYINPUT8), .ZN(n1081) );
XOR2_X1 U997 ( .A(n1322), .B(n1163), .Z(n1111) );
NAND2_X1 U998 ( .A1(G217), .A2(n1323), .ZN(n1163) );
NAND2_X1 U999 ( .A1(n1161), .A2(n1314), .ZN(n1322) );
XNOR2_X1 U1000 ( .A(n1324), .B(n1325), .ZN(n1161) );
XOR2_X1 U1001 ( .A(G119), .B(n1326), .Z(n1325) );
XOR2_X1 U1002 ( .A(G137), .B(G125), .Z(n1326) );
XOR2_X1 U1003 ( .A(n1327), .B(n1193), .Z(n1324) );
XNOR2_X1 U1004 ( .A(n1328), .B(n1329), .ZN(n1327) );
AND3_X1 U1005 ( .A1(G221), .A2(n1065), .A3(G234), .ZN(n1329) );
INV_X1 U1006 ( .A(n1235), .ZN(n1056) );
NOR3_X1 U1007 ( .A1(n1241), .A2(n1300), .A3(n1094), .ZN(n1235) );
INV_X1 U1008 ( .A(n1098), .ZN(n1094) );
NOR2_X1 U1009 ( .A1(n1071), .A2(n1101), .ZN(n1098) );
INV_X1 U1010 ( .A(n1074), .ZN(n1101) );
NAND2_X1 U1011 ( .A1(G221), .A2(n1323), .ZN(n1074) );
NAND2_X1 U1012 ( .A1(G234), .A2(n1330), .ZN(n1323) );
XNOR2_X1 U1013 ( .A(n1116), .B(n1331), .ZN(n1071) );
NOR2_X1 U1014 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
NOR2_X1 U1015 ( .A1(KEYINPUT30), .A2(n1334), .ZN(n1333) );
INV_X1 U1016 ( .A(n1117), .ZN(n1334) );
NOR2_X1 U1017 ( .A1(KEYINPUT18), .A2(n1117), .ZN(n1332) );
NAND2_X1 U1018 ( .A1(n1335), .A2(n1314), .ZN(n1117) );
XOR2_X1 U1019 ( .A(n1336), .B(n1337), .Z(n1335) );
XNOR2_X1 U1020 ( .A(n1201), .B(n1338), .ZN(n1337) );
NOR2_X1 U1021 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
NOR2_X1 U1022 ( .A1(KEYINPUT36), .A2(n1341), .ZN(n1340) );
INV_X1 U1023 ( .A(n1204), .ZN(n1341) );
NOR2_X1 U1024 ( .A1(KEYINPUT11), .A2(n1204), .ZN(n1339) );
NAND2_X1 U1025 ( .A1(G227), .A2(n1065), .ZN(n1204) );
XOR2_X1 U1026 ( .A(n1342), .B(n1343), .Z(n1201) );
XOR2_X1 U1027 ( .A(G104), .B(G101), .Z(n1343) );
NAND2_X1 U1028 ( .A1(KEYINPUT35), .A2(n1344), .ZN(n1342) );
XNOR2_X1 U1029 ( .A(n1193), .B(n1345), .ZN(n1336) );
XOR2_X1 U1030 ( .A(n1346), .B(n1198), .Z(n1345) );
INV_X1 U1031 ( .A(n1143), .ZN(n1198) );
XOR2_X1 U1032 ( .A(n1347), .B(n1348), .Z(n1143) );
NOR2_X1 U1033 ( .A1(KEYINPUT54), .A2(n1349), .ZN(n1348) );
XOR2_X1 U1034 ( .A(G146), .B(G143), .Z(n1349) );
NOR2_X1 U1035 ( .A1(KEYINPUT4), .A2(n1191), .ZN(n1346) );
AND2_X1 U1036 ( .A1(n1350), .A2(n1351), .ZN(n1191) );
NAND2_X1 U1037 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
INV_X1 U1038 ( .A(G131), .ZN(n1353) );
XOR2_X1 U1039 ( .A(n1354), .B(KEYINPUT33), .Z(n1352) );
NAND2_X1 U1040 ( .A1(n1355), .A2(G131), .ZN(n1350) );
XOR2_X1 U1041 ( .A(KEYINPUT29), .B(n1140), .Z(n1355) );
INV_X1 U1042 ( .A(n1354), .ZN(n1140) );
XNOR2_X1 U1043 ( .A(G134), .B(G137), .ZN(n1354) );
XNOR2_X1 U1044 ( .A(n1142), .B(n1356), .ZN(n1193) );
INV_X1 U1045 ( .A(G469), .ZN(n1116) );
INV_X1 U1046 ( .A(n1248), .ZN(n1300) );
NAND2_X1 U1047 ( .A1(n1103), .A2(n1357), .ZN(n1248) );
NAND4_X1 U1048 ( .A1(G953), .A2(G902), .A3(n1298), .A4(n1155), .ZN(n1357) );
INV_X1 U1049 ( .A(G898), .ZN(n1155) );
NAND3_X1 U1050 ( .A1(n1298), .A2(n1065), .A3(G952), .ZN(n1103) );
NAND2_X1 U1051 ( .A1(G237), .A2(G234), .ZN(n1298) );
XNOR2_X1 U1052 ( .A(n1086), .B(KEYINPUT14), .ZN(n1241) );
NAND2_X1 U1053 ( .A1(n1292), .A2(n1090), .ZN(n1086) );
NAND2_X1 U1054 ( .A1(G214), .A2(n1358), .ZN(n1090) );
XNOR2_X1 U1055 ( .A(n1359), .B(n1126), .ZN(n1292) );
NAND2_X1 U1056 ( .A1(G210), .A2(n1358), .ZN(n1126) );
NAND2_X1 U1057 ( .A1(n1360), .A2(n1330), .ZN(n1358) );
XOR2_X1 U1058 ( .A(G902), .B(KEYINPUT45), .Z(n1330) );
XNOR2_X1 U1059 ( .A(G237), .B(KEYINPUT21), .ZN(n1360) );
NAND2_X1 U1060 ( .A1(KEYINPUT39), .A2(n1127), .ZN(n1359) );
NAND2_X1 U1061 ( .A1(n1361), .A2(n1314), .ZN(n1127) );
XOR2_X1 U1062 ( .A(n1362), .B(n1363), .Z(n1361) );
XOR2_X1 U1063 ( .A(n1221), .B(n1215), .Z(n1363) );
XOR2_X1 U1064 ( .A(n1158), .B(n1364), .Z(n1215) );
NOR2_X1 U1065 ( .A1(KEYINPUT50), .A2(n1156), .ZN(n1364) );
XNOR2_X1 U1066 ( .A(n1365), .B(n1366), .ZN(n1156) );
XOR2_X1 U1067 ( .A(n1367), .B(n1320), .Z(n1366) );
XOR2_X1 U1068 ( .A(G116), .B(n1303), .Z(n1320) );
INV_X1 U1069 ( .A(G119), .ZN(n1303) );
NAND2_X1 U1070 ( .A1(KEYINPUT40), .A2(n1368), .ZN(n1367) );
XOR2_X1 U1071 ( .A(G107), .B(G104), .Z(n1368) );
XNOR2_X1 U1072 ( .A(G101), .B(G113), .ZN(n1365) );
XOR2_X1 U1073 ( .A(G122), .B(n1356), .Z(n1158) );
XOR2_X1 U1074 ( .A(G110), .B(KEYINPUT48), .Z(n1356) );
INV_X1 U1075 ( .A(n1225), .ZN(n1221) );
XOR2_X1 U1076 ( .A(n1269), .B(n1328), .Z(n1225) );
XOR2_X1 U1077 ( .A(G146), .B(n1369), .Z(n1328) );
INV_X1 U1078 ( .A(G143), .ZN(n1269) );
XOR2_X1 U1079 ( .A(n1222), .B(n1370), .Z(n1362) );
NOR2_X1 U1080 ( .A1(G125), .A2(KEYINPUT42), .ZN(n1370) );
INV_X1 U1081 ( .A(n1226), .ZN(n1222) );
NAND2_X1 U1082 ( .A1(G224), .A2(n1065), .ZN(n1226) );
NAND2_X1 U1083 ( .A1(n1106), .A2(n1271), .ZN(n1095) );
INV_X1 U1084 ( .A(n1310), .ZN(n1271) );
NAND3_X1 U1085 ( .A1(n1371), .A2(n1372), .A3(n1373), .ZN(n1310) );
NAND2_X1 U1086 ( .A1(G475), .A2(n1112), .ZN(n1373) );
NAND2_X1 U1087 ( .A1(KEYINPUT0), .A2(n1374), .ZN(n1372) );
NAND2_X1 U1088 ( .A1(n1375), .A2(n1125), .ZN(n1374) );
XOR2_X1 U1089 ( .A(n1112), .B(KEYINPUT56), .Z(n1375) );
INV_X1 U1090 ( .A(n1124), .ZN(n1112) );
NAND2_X1 U1091 ( .A1(n1376), .A2(n1377), .ZN(n1371) );
INV_X1 U1092 ( .A(KEYINPUT0), .ZN(n1377) );
NAND2_X1 U1093 ( .A1(n1378), .A2(n1379), .ZN(n1376) );
OR2_X1 U1094 ( .A1(n1124), .A2(KEYINPUT56), .ZN(n1379) );
NAND3_X1 U1095 ( .A1(n1124), .A2(n1125), .A3(KEYINPUT56), .ZN(n1378) );
INV_X1 U1096 ( .A(G475), .ZN(n1125) );
NOR2_X1 U1097 ( .A1(n1173), .A2(G902), .ZN(n1124) );
XOR2_X1 U1098 ( .A(n1380), .B(n1381), .Z(n1173) );
XOR2_X1 U1099 ( .A(n1382), .B(n1383), .Z(n1381) );
XOR2_X1 U1100 ( .A(n1384), .B(n1141), .Z(n1383) );
XOR2_X1 U1101 ( .A(G131), .B(G125), .Z(n1141) );
NAND2_X1 U1102 ( .A1(KEYINPUT10), .A2(n1142), .ZN(n1384) );
INV_X1 U1103 ( .A(G140), .ZN(n1142) );
XOR2_X1 U1104 ( .A(n1385), .B(n1386), .Z(n1382) );
NOR2_X1 U1105 ( .A1(G146), .A2(KEYINPUT23), .ZN(n1386) );
NAND2_X1 U1106 ( .A1(G214), .A2(n1316), .ZN(n1385) );
NOR2_X1 U1107 ( .A1(G953), .A2(G237), .ZN(n1316) );
XOR2_X1 U1108 ( .A(n1387), .B(n1388), .Z(n1380) );
XOR2_X1 U1109 ( .A(G143), .B(G122), .Z(n1388) );
XNOR2_X1 U1110 ( .A(G104), .B(G113), .ZN(n1387) );
XOR2_X1 U1111 ( .A(n1389), .B(G478), .Z(n1106) );
NAND2_X1 U1112 ( .A1(n1169), .A2(n1314), .ZN(n1389) );
INV_X1 U1113 ( .A(G902), .ZN(n1314) );
XNOR2_X1 U1114 ( .A(n1390), .B(n1391), .ZN(n1169) );
XOR2_X1 U1115 ( .A(n1392), .B(n1393), .Z(n1391) );
XOR2_X1 U1116 ( .A(G116), .B(n1344), .Z(n1393) );
INV_X1 U1117 ( .A(G107), .ZN(n1344) );
NAND3_X1 U1118 ( .A1(G217), .A2(n1065), .A3(G234), .ZN(n1392) );
INV_X1 U1119 ( .A(G953), .ZN(n1065) );
XNOR2_X1 U1120 ( .A(n1394), .B(n1395), .ZN(n1390) );
NAND2_X1 U1121 ( .A1(KEYINPUT62), .A2(n1396), .ZN(n1395) );
XOR2_X1 U1122 ( .A(n1369), .B(n1397), .Z(n1396) );
XOR2_X1 U1123 ( .A(G143), .B(G134), .Z(n1397) );
INV_X1 U1124 ( .A(n1347), .ZN(n1369) );
XNOR2_X1 U1125 ( .A(G128), .B(KEYINPUT55), .ZN(n1347) );
NAND2_X1 U1126 ( .A1(KEYINPUT32), .A2(G122), .ZN(n1394) );
endmodule


