//Key = 1011100100010001011000100011110101111101000110100100001011100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388;

XOR2_X1 U756 ( .A(n1048), .B(n1049), .Z(G9) );
NOR3_X1 U757 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
XNOR2_X1 U758 ( .A(n1053), .B(KEYINPUT8), .ZN(n1051) );
NAND2_X1 U759 ( .A1(n1054), .A2(KEYINPUT36), .ZN(n1048) );
XNOR2_X1 U760 ( .A(G107), .B(KEYINPUT32), .ZN(n1054) );
NOR2_X1 U761 ( .A1(n1055), .A2(n1056), .ZN(G75) );
NOR3_X1 U762 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
NAND3_X1 U763 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1057) );
NAND2_X1 U764 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U765 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND3_X1 U766 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
NAND2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NAND2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1070) );
NAND2_X1 U771 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U772 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND3_X1 U773 ( .A1(n1082), .A2(n1083), .A3(n1076), .ZN(n1065) );
NAND2_X1 U774 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
OR3_X1 U775 ( .A1(n1086), .A2(KEYINPUT34), .A3(n1052), .ZN(n1084) );
NAND4_X1 U776 ( .A1(n1087), .A2(n1088), .A3(n1089), .A4(n1072), .ZN(n1082) );
NAND2_X1 U777 ( .A1(n1069), .A2(n1090), .ZN(n1089) );
NAND2_X1 U778 ( .A1(n1067), .A2(n1091), .ZN(n1088) );
NAND2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U780 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U781 ( .A1(KEYINPUT34), .A2(n1096), .ZN(n1092) );
NAND2_X1 U782 ( .A1(n1097), .A2(n1098), .ZN(n1087) );
XNOR2_X1 U783 ( .A(n1069), .B(KEYINPUT39), .ZN(n1097) );
INV_X1 U784 ( .A(n1099), .ZN(n1063) );
AND3_X1 U785 ( .A1(n1060), .A2(n1061), .A3(n1100), .ZN(n1055) );
NAND4_X1 U786 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1060) );
NOR4_X1 U787 ( .A1(n1105), .A2(n1106), .A3(n1085), .A4(n1107), .ZN(n1104) );
XNOR2_X1 U788 ( .A(G472), .B(n1108), .ZN(n1107) );
XNOR2_X1 U789 ( .A(n1109), .B(KEYINPUT56), .ZN(n1105) );
NOR3_X1 U790 ( .A1(n1094), .A2(n1110), .A3(n1111), .ZN(n1103) );
NAND2_X1 U791 ( .A1(n1112), .A2(n1113), .ZN(n1102) );
XOR2_X1 U792 ( .A(KEYINPUT57), .B(n1114), .Z(n1101) );
NAND2_X1 U793 ( .A1(n1115), .A2(n1116), .ZN(G72) );
NAND2_X1 U794 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U795 ( .A1(n1119), .A2(n1120), .ZN(n1115) );
NAND2_X1 U796 ( .A1(n1121), .A2(n1118), .ZN(n1120) );
NAND2_X1 U797 ( .A1(G953), .A2(n1122), .ZN(n1118) );
INV_X1 U798 ( .A(n1117), .ZN(n1119) );
XNOR2_X1 U799 ( .A(n1123), .B(n1124), .ZN(n1117) );
AND2_X1 U800 ( .A1(n1058), .A2(n1061), .ZN(n1124) );
NAND4_X1 U801 ( .A1(n1121), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1123) );
NAND2_X1 U802 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
INV_X1 U803 ( .A(KEYINPUT47), .ZN(n1129) );
NAND2_X1 U804 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
NAND3_X1 U805 ( .A1(n1131), .A2(n1130), .A3(KEYINPUT47), .ZN(n1126) );
NAND3_X1 U806 ( .A1(n1132), .A2(n1133), .A3(KEYINPUT61), .ZN(n1130) );
NAND2_X1 U807 ( .A1(n1134), .A2(n1135), .ZN(n1131) );
INV_X1 U808 ( .A(KEYINPUT61), .ZN(n1135) );
INV_X1 U809 ( .A(n1133), .ZN(n1134) );
OR2_X1 U810 ( .A1(n1133), .A2(n1132), .ZN(n1125) );
NAND2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(n1133) );
OR2_X1 U812 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
XOR2_X1 U813 ( .A(n1140), .B(KEYINPUT41), .Z(n1136) );
NAND2_X1 U814 ( .A1(n1138), .A2(n1139), .ZN(n1140) );
XNOR2_X1 U815 ( .A(n1141), .B(n1142), .ZN(n1138) );
NOR2_X1 U816 ( .A1(G131), .A2(n1143), .ZN(n1142) );
XNOR2_X1 U817 ( .A(KEYINPUT42), .B(KEYINPUT2), .ZN(n1143) );
XNOR2_X1 U818 ( .A(G134), .B(G137), .ZN(n1141) );
INV_X1 U819 ( .A(n1144), .ZN(n1121) );
NAND2_X1 U820 ( .A1(n1145), .A2(n1146), .ZN(G69) );
NAND2_X1 U821 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U822 ( .A1(G953), .A2(n1149), .ZN(n1148) );
NAND2_X1 U823 ( .A1(G898), .A2(G224), .ZN(n1149) );
NAND2_X1 U824 ( .A1(n1150), .A2(n1151), .ZN(n1145) );
NAND2_X1 U825 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U826 ( .A1(G953), .A2(n1154), .ZN(n1153) );
INV_X1 U827 ( .A(n1155), .ZN(n1152) );
INV_X1 U828 ( .A(n1147), .ZN(n1150) );
XNOR2_X1 U829 ( .A(n1156), .B(n1157), .ZN(n1147) );
NOR2_X1 U830 ( .A1(n1155), .A2(n1158), .ZN(n1157) );
XOR2_X1 U831 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND2_X1 U832 ( .A1(n1161), .A2(n1162), .ZN(n1159) );
OR2_X1 U833 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U834 ( .A(n1165), .B(KEYINPUT14), .Z(n1161) );
NAND2_X1 U835 ( .A1(n1164), .A2(n1163), .ZN(n1165) );
NAND2_X1 U836 ( .A1(n1166), .A2(n1059), .ZN(n1156) );
XNOR2_X1 U837 ( .A(KEYINPUT27), .B(n1061), .ZN(n1166) );
NOR2_X1 U838 ( .A1(n1167), .A2(n1168), .ZN(G66) );
XOR2_X1 U839 ( .A(n1169), .B(n1170), .Z(n1168) );
AND2_X1 U840 ( .A1(G217), .A2(n1171), .ZN(n1169) );
NOR2_X1 U841 ( .A1(n1167), .A2(n1172), .ZN(G63) );
XOR2_X1 U842 ( .A(n1173), .B(n1174), .Z(n1172) );
AND2_X1 U843 ( .A1(G478), .A2(n1171), .ZN(n1173) );
NOR2_X1 U844 ( .A1(n1167), .A2(n1175), .ZN(G60) );
XNOR2_X1 U845 ( .A(n1176), .B(n1177), .ZN(n1175) );
AND2_X1 U846 ( .A1(G475), .A2(n1171), .ZN(n1177) );
XOR2_X1 U847 ( .A(n1178), .B(n1179), .Z(G6) );
NAND2_X1 U848 ( .A1(n1180), .A2(KEYINPUT31), .ZN(n1179) );
XNOR2_X1 U849 ( .A(G104), .B(KEYINPUT0), .ZN(n1180) );
NAND2_X1 U850 ( .A1(n1181), .A2(n1096), .ZN(n1178) );
XOR2_X1 U851 ( .A(n1182), .B(KEYINPUT49), .Z(n1181) );
NOR2_X1 U852 ( .A1(n1167), .A2(n1183), .ZN(G57) );
XOR2_X1 U853 ( .A(n1184), .B(n1185), .Z(n1183) );
XOR2_X1 U854 ( .A(n1186), .B(n1187), .Z(n1184) );
AND2_X1 U855 ( .A1(G472), .A2(n1171), .ZN(n1187) );
NAND2_X1 U856 ( .A1(KEYINPUT11), .A2(n1188), .ZN(n1186) );
NOR3_X1 U857 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(G54) );
NOR3_X1 U858 ( .A1(n1192), .A2(G952), .A3(n1193), .ZN(n1191) );
INV_X1 U859 ( .A(KEYINPUT13), .ZN(n1192) );
NOR2_X1 U860 ( .A1(KEYINPUT13), .A2(n1194), .ZN(n1190) );
XOR2_X1 U861 ( .A(n1195), .B(n1196), .Z(n1189) );
XOR2_X1 U862 ( .A(n1197), .B(n1198), .Z(n1196) );
AND2_X1 U863 ( .A1(G469), .A2(n1171), .ZN(n1198) );
XNOR2_X1 U864 ( .A(G110), .B(n1199), .ZN(n1195) );
XNOR2_X1 U865 ( .A(KEYINPUT12), .B(n1200), .ZN(n1199) );
NOR2_X1 U866 ( .A1(n1167), .A2(n1201), .ZN(G51) );
XOR2_X1 U867 ( .A(n1202), .B(n1203), .Z(n1201) );
NOR2_X1 U868 ( .A1(KEYINPUT45), .A2(n1204), .ZN(n1203) );
XOR2_X1 U869 ( .A(n1205), .B(n1206), .Z(n1204) );
NAND2_X1 U870 ( .A1(n1207), .A2(n1208), .ZN(n1205) );
NAND2_X1 U871 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XOR2_X1 U872 ( .A(KEYINPUT33), .B(n1211), .Z(n1207) );
NOR2_X1 U873 ( .A1(n1209), .A2(n1210), .ZN(n1211) );
NAND2_X1 U874 ( .A1(n1171), .A2(n1212), .ZN(n1202) );
AND2_X1 U875 ( .A1(G902), .A2(n1213), .ZN(n1171) );
OR2_X1 U876 ( .A1(n1059), .A2(n1058), .ZN(n1213) );
NAND2_X1 U877 ( .A1(n1214), .A2(n1215), .ZN(n1058) );
NOR4_X1 U878 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1215) );
INV_X1 U879 ( .A(n1220), .ZN(n1216) );
NOR4_X1 U880 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1214) );
NOR2_X1 U881 ( .A1(n1075), .A2(n1225), .ZN(n1224) );
NOR3_X1 U882 ( .A1(n1226), .A2(n1227), .A3(n1074), .ZN(n1223) );
INV_X1 U883 ( .A(n1228), .ZN(n1222) );
NAND4_X1 U884 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1059) );
NOR4_X1 U885 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1232) );
NOR2_X1 U886 ( .A1(n1237), .A2(n1238), .ZN(n1231) );
NOR2_X1 U887 ( .A1(n1086), .A2(n1182), .ZN(n1238) );
NAND4_X1 U888 ( .A1(n1239), .A2(n1067), .A3(n1240), .A4(n1241), .ZN(n1182) );
NOR3_X1 U889 ( .A1(n1050), .A2(n1075), .A3(n1052), .ZN(n1237) );
INV_X1 U890 ( .A(n1194), .ZN(n1167) );
NAND2_X1 U891 ( .A1(n1193), .A2(n1100), .ZN(n1194) );
INV_X1 U892 ( .A(G952), .ZN(n1100) );
XNOR2_X1 U893 ( .A(G953), .B(KEYINPUT54), .ZN(n1193) );
NAND2_X1 U894 ( .A1(n1242), .A2(n1243), .ZN(G48) );
NAND2_X1 U895 ( .A1(G146), .A2(n1244), .ZN(n1243) );
XOR2_X1 U896 ( .A(KEYINPUT18), .B(n1245), .Z(n1242) );
NOR2_X1 U897 ( .A1(G146), .A2(n1244), .ZN(n1245) );
INV_X1 U898 ( .A(n1221), .ZN(n1244) );
NOR2_X1 U899 ( .A1(n1225), .A2(n1074), .ZN(n1221) );
NAND3_X1 U900 ( .A1(n1246), .A2(n1240), .A3(n1247), .ZN(n1225) );
XNOR2_X1 U901 ( .A(G143), .B(n1228), .ZN(G45) );
NAND3_X1 U902 ( .A1(n1247), .A2(n1098), .A3(n1248), .ZN(n1228) );
AND3_X1 U903 ( .A1(n1249), .A2(n1106), .A3(n1240), .ZN(n1248) );
XNOR2_X1 U904 ( .A(n1200), .B(n1250), .ZN(G42) );
NOR3_X1 U905 ( .A1(n1226), .A2(n1251), .A3(n1227), .ZN(n1250) );
XNOR2_X1 U906 ( .A(n1239), .B(KEYINPUT19), .ZN(n1251) );
XNOR2_X1 U907 ( .A(n1252), .B(n1219), .ZN(G39) );
AND3_X1 U908 ( .A1(n1246), .A2(n1076), .A3(n1253), .ZN(n1219) );
XNOR2_X1 U909 ( .A(n1254), .B(n1218), .ZN(G36) );
AND3_X1 U910 ( .A1(n1098), .A2(n1053), .A3(n1253), .ZN(n1218) );
XOR2_X1 U911 ( .A(G131), .B(n1217), .Z(G33) );
AND3_X1 U912 ( .A1(n1098), .A2(n1239), .A3(n1253), .ZN(n1217) );
INV_X1 U913 ( .A(n1226), .ZN(n1253) );
NAND3_X1 U914 ( .A1(n1240), .A2(n1255), .A3(n1069), .ZN(n1226) );
AND2_X1 U915 ( .A1(n1095), .A2(n1256), .ZN(n1069) );
XOR2_X1 U916 ( .A(n1109), .B(KEYINPUT3), .Z(n1095) );
XNOR2_X1 U917 ( .A(G128), .B(n1257), .ZN(G30) );
NAND4_X1 U918 ( .A1(n1247), .A2(n1246), .A3(n1053), .A4(n1258), .ZN(n1257) );
XNOR2_X1 U919 ( .A(KEYINPUT21), .B(n1078), .ZN(n1258) );
INV_X1 U920 ( .A(n1240), .ZN(n1078) );
NAND2_X1 U921 ( .A1(n1259), .A2(n1260), .ZN(G3) );
NAND2_X1 U922 ( .A1(G101), .A2(n1229), .ZN(n1260) );
XOR2_X1 U923 ( .A(KEYINPUT43), .B(n1261), .Z(n1259) );
NOR2_X1 U924 ( .A1(G101), .A2(n1229), .ZN(n1261) );
NAND3_X1 U925 ( .A1(n1076), .A2(n1262), .A3(n1098), .ZN(n1229) );
XNOR2_X1 U926 ( .A(G125), .B(n1220), .ZN(G27) );
NAND4_X1 U927 ( .A1(n1247), .A2(n1239), .A3(n1090), .A4(n1072), .ZN(n1220) );
AND2_X1 U928 ( .A1(n1096), .A2(n1255), .ZN(n1247) );
NAND2_X1 U929 ( .A1(n1263), .A2(n1099), .ZN(n1255) );
NAND2_X1 U930 ( .A1(n1144), .A2(n1264), .ZN(n1263) );
NOR2_X1 U931 ( .A1(G900), .A2(n1061), .ZN(n1144) );
XOR2_X1 U932 ( .A(n1230), .B(n1265), .Z(G24) );
NAND2_X1 U933 ( .A1(KEYINPUT28), .A2(G122), .ZN(n1265) );
NAND4_X1 U934 ( .A1(n1266), .A2(n1067), .A3(n1249), .A4(n1106), .ZN(n1230) );
INV_X1 U935 ( .A(n1052), .ZN(n1067) );
NAND2_X1 U936 ( .A1(n1267), .A2(n1268), .ZN(n1052) );
XOR2_X1 U937 ( .A(G119), .B(n1236), .Z(G21) );
AND3_X1 U938 ( .A1(n1266), .A2(n1076), .A3(n1246), .ZN(n1236) );
AND2_X1 U939 ( .A1(n1269), .A2(n1270), .ZN(n1246) );
XNOR2_X1 U940 ( .A(n1268), .B(KEYINPUT20), .ZN(n1269) );
XOR2_X1 U941 ( .A(G116), .B(n1235), .Z(G18) );
AND3_X1 U942 ( .A1(n1098), .A2(n1053), .A3(n1266), .ZN(n1235) );
INV_X1 U943 ( .A(n1075), .ZN(n1053) );
NAND2_X1 U944 ( .A1(n1249), .A2(n1271), .ZN(n1075) );
XNOR2_X1 U945 ( .A(n1272), .B(KEYINPUT60), .ZN(n1249) );
XNOR2_X1 U946 ( .A(n1273), .B(n1234), .ZN(G15) );
AND3_X1 U947 ( .A1(n1098), .A2(n1239), .A3(n1266), .ZN(n1234) );
AND3_X1 U948 ( .A1(n1096), .A2(n1241), .A3(n1072), .ZN(n1266) );
INV_X1 U949 ( .A(n1085), .ZN(n1072) );
NAND2_X1 U950 ( .A1(n1081), .A2(n1274), .ZN(n1085) );
INV_X1 U951 ( .A(n1074), .ZN(n1239) );
NAND2_X1 U952 ( .A1(n1272), .A2(n1106), .ZN(n1074) );
AND2_X1 U953 ( .A1(n1275), .A2(n1267), .ZN(n1098) );
XNOR2_X1 U954 ( .A(KEYINPUT24), .B(n1270), .ZN(n1267) );
INV_X1 U955 ( .A(n1268), .ZN(n1275) );
XNOR2_X1 U956 ( .A(n1276), .B(n1233), .ZN(G12) );
AND3_X1 U957 ( .A1(n1076), .A2(n1262), .A3(n1090), .ZN(n1233) );
INV_X1 U958 ( .A(n1227), .ZN(n1090) );
NAND2_X1 U959 ( .A1(n1268), .A2(n1270), .ZN(n1227) );
NAND3_X1 U960 ( .A1(n1277), .A2(n1278), .A3(n1279), .ZN(n1270) );
INV_X1 U961 ( .A(n1111), .ZN(n1279) );
NOR2_X1 U962 ( .A1(n1113), .A2(n1112), .ZN(n1111) );
OR2_X1 U963 ( .A1(n1112), .A2(KEYINPUT37), .ZN(n1278) );
NAND3_X1 U964 ( .A1(n1112), .A2(n1113), .A3(KEYINPUT37), .ZN(n1277) );
OR2_X1 U965 ( .A1(n1170), .A2(G902), .ZN(n1113) );
XNOR2_X1 U966 ( .A(n1280), .B(n1281), .ZN(n1170) );
XOR2_X1 U967 ( .A(G119), .B(n1282), .Z(n1281) );
XNOR2_X1 U968 ( .A(n1252), .B(G128), .ZN(n1282) );
XOR2_X1 U969 ( .A(n1283), .B(n1284), .Z(n1280) );
AND3_X1 U970 ( .A1(G221), .A2(n1061), .A3(G234), .ZN(n1284) );
XNOR2_X1 U971 ( .A(n1285), .B(n1276), .ZN(n1283) );
NAND2_X1 U972 ( .A1(KEYINPUT22), .A2(n1286), .ZN(n1285) );
XOR2_X1 U973 ( .A(n1287), .B(n1132), .Z(n1286) );
XOR2_X1 U974 ( .A(G140), .B(G125), .Z(n1132) );
AND2_X1 U975 ( .A1(n1288), .A2(G217), .ZN(n1112) );
XOR2_X1 U976 ( .A(n1289), .B(KEYINPUT52), .Z(n1288) );
XNOR2_X1 U977 ( .A(n1108), .B(n1290), .ZN(n1268) );
NOR2_X1 U978 ( .A1(G472), .A2(KEYINPUT55), .ZN(n1290) );
NAND2_X1 U979 ( .A1(n1291), .A2(n1292), .ZN(n1108) );
XOR2_X1 U980 ( .A(n1188), .B(n1185), .Z(n1291) );
XNOR2_X1 U981 ( .A(n1293), .B(n1294), .ZN(n1185) );
XNOR2_X1 U982 ( .A(n1295), .B(n1209), .ZN(n1294) );
AND2_X1 U983 ( .A1(G210), .A2(n1296), .ZN(n1295) );
XOR2_X1 U984 ( .A(G113), .B(n1297), .Z(n1188) );
XOR2_X1 U985 ( .A(G119), .B(G116), .Z(n1297) );
INV_X1 U986 ( .A(n1050), .ZN(n1262) );
NAND3_X1 U987 ( .A1(n1096), .A2(n1241), .A3(n1240), .ZN(n1050) );
NOR2_X1 U988 ( .A1(n1081), .A2(n1080), .ZN(n1240) );
INV_X1 U989 ( .A(n1274), .ZN(n1080) );
NAND2_X1 U990 ( .A1(G221), .A2(n1289), .ZN(n1274) );
NAND2_X1 U991 ( .A1(G234), .A2(n1292), .ZN(n1289) );
XOR2_X1 U992 ( .A(n1298), .B(n1299), .Z(n1081) );
XOR2_X1 U993 ( .A(KEYINPUT30), .B(G469), .Z(n1299) );
NAND2_X1 U994 ( .A1(n1300), .A2(n1292), .ZN(n1298) );
XOR2_X1 U995 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U996 ( .A(n1303), .B(n1197), .Z(n1302) );
XOR2_X1 U997 ( .A(n1304), .B(n1305), .Z(n1197) );
XOR2_X1 U998 ( .A(n1306), .B(n1139), .Z(n1305) );
XNOR2_X1 U999 ( .A(n1307), .B(KEYINPUT35), .ZN(n1139) );
NAND3_X1 U1000 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1307) );
NAND2_X1 U1001 ( .A1(G128), .A2(n1311), .ZN(n1310) );
NAND2_X1 U1002 ( .A1(KEYINPUT25), .A2(n1312), .ZN(n1309) );
NAND2_X1 U1003 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XNOR2_X1 U1004 ( .A(KEYINPUT4), .B(n1315), .ZN(n1313) );
NAND2_X1 U1005 ( .A1(n1316), .A2(n1317), .ZN(n1308) );
INV_X1 U1006 ( .A(KEYINPUT25), .ZN(n1317) );
NAND2_X1 U1007 ( .A1(n1318), .A2(n1319), .ZN(n1316) );
NAND3_X1 U1008 ( .A1(KEYINPUT4), .A2(n1314), .A3(n1315), .ZN(n1319) );
OR2_X1 U1009 ( .A1(n1315), .A2(KEYINPUT4), .ZN(n1318) );
XOR2_X1 U1010 ( .A(n1293), .B(n1320), .Z(n1304) );
XOR2_X1 U1011 ( .A(G107), .B(n1321), .Z(n1320) );
NOR2_X1 U1012 ( .A1(G953), .A2(n1122), .ZN(n1321) );
INV_X1 U1013 ( .A(G227), .ZN(n1122) );
XOR2_X1 U1014 ( .A(n1322), .B(n1323), .Z(n1293) );
XNOR2_X1 U1015 ( .A(n1254), .B(G131), .ZN(n1323) );
XOR2_X1 U1016 ( .A(n1324), .B(G101), .Z(n1322) );
NAND2_X1 U1017 ( .A1(KEYINPUT29), .A2(n1252), .ZN(n1324) );
INV_X1 U1018 ( .A(G137), .ZN(n1252) );
NAND2_X1 U1019 ( .A1(KEYINPUT44), .A2(n1200), .ZN(n1303) );
XNOR2_X1 U1020 ( .A(KEYINPUT40), .B(n1276), .ZN(n1301) );
NAND2_X1 U1021 ( .A1(n1325), .A2(n1099), .ZN(n1241) );
NAND3_X1 U1022 ( .A1(n1326), .A2(n1061), .A3(G952), .ZN(n1099) );
XOR2_X1 U1023 ( .A(n1327), .B(KEYINPUT1), .Z(n1325) );
NAND2_X1 U1024 ( .A1(n1155), .A2(n1264), .ZN(n1327) );
AND2_X1 U1025 ( .A1(n1328), .A2(n1326), .ZN(n1264) );
NAND2_X1 U1026 ( .A1(G237), .A2(G234), .ZN(n1326) );
XNOR2_X1 U1027 ( .A(KEYINPUT59), .B(n1292), .ZN(n1328) );
NOR2_X1 U1028 ( .A1(n1061), .A2(G898), .ZN(n1155) );
INV_X1 U1029 ( .A(n1086), .ZN(n1096) );
NAND2_X1 U1030 ( .A1(n1329), .A2(n1109), .ZN(n1086) );
XNOR2_X1 U1031 ( .A(n1330), .B(n1212), .ZN(n1109) );
AND2_X1 U1032 ( .A1(G210), .A2(n1331), .ZN(n1212) );
NAND2_X1 U1033 ( .A1(n1332), .A2(n1292), .ZN(n1330) );
XOR2_X1 U1034 ( .A(n1333), .B(n1334), .Z(n1332) );
XNOR2_X1 U1035 ( .A(n1206), .B(n1209), .ZN(n1334) );
XNOR2_X1 U1036 ( .A(n1315), .B(n1311), .ZN(n1209) );
XOR2_X1 U1037 ( .A(n1335), .B(n1160), .Z(n1206) );
XOR2_X1 U1038 ( .A(G122), .B(n1336), .Z(n1160) );
NOR2_X1 U1039 ( .A1(G110), .A2(KEYINPUT50), .ZN(n1336) );
XOR2_X1 U1040 ( .A(n1337), .B(n1338), .Z(n1335) );
NOR2_X1 U1041 ( .A1(G953), .A2(n1154), .ZN(n1338) );
INV_X1 U1042 ( .A(G224), .ZN(n1154) );
NAND3_X1 U1043 ( .A1(n1339), .A2(n1340), .A3(n1341), .ZN(n1337) );
NAND2_X1 U1044 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
OR3_X1 U1045 ( .A1(n1343), .A2(n1342), .A3(KEYINPUT51), .ZN(n1340) );
INV_X1 U1046 ( .A(n1163), .ZN(n1342) );
NAND2_X1 U1047 ( .A1(n1344), .A2(n1345), .ZN(n1163) );
NAND2_X1 U1048 ( .A1(n1346), .A2(n1273), .ZN(n1345) );
XOR2_X1 U1049 ( .A(KEYINPUT15), .B(n1347), .Z(n1344) );
NOR2_X1 U1050 ( .A1(n1346), .A2(n1273), .ZN(n1347) );
INV_X1 U1051 ( .A(G113), .ZN(n1273) );
XOR2_X1 U1052 ( .A(G119), .B(n1348), .Z(n1346) );
NOR2_X1 U1053 ( .A1(G116), .A2(KEYINPUT38), .ZN(n1348) );
OR2_X1 U1054 ( .A1(KEYINPUT6), .A2(n1164), .ZN(n1343) );
NAND2_X1 U1055 ( .A1(KEYINPUT51), .A2(n1164), .ZN(n1339) );
XNOR2_X1 U1056 ( .A(G101), .B(n1349), .ZN(n1164) );
NOR2_X1 U1057 ( .A1(n1350), .A2(KEYINPUT10), .ZN(n1349) );
NOR2_X1 U1058 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
XOR2_X1 U1059 ( .A(n1353), .B(KEYINPUT62), .Z(n1352) );
NAND2_X1 U1060 ( .A1(G107), .A2(n1306), .ZN(n1353) );
NOR2_X1 U1061 ( .A1(G107), .A2(n1306), .ZN(n1351) );
XOR2_X1 U1062 ( .A(G104), .B(KEYINPUT46), .Z(n1306) );
XNOR2_X1 U1063 ( .A(G125), .B(KEYINPUT26), .ZN(n1333) );
XNOR2_X1 U1064 ( .A(n1094), .B(KEYINPUT9), .ZN(n1329) );
INV_X1 U1065 ( .A(n1256), .ZN(n1094) );
NAND2_X1 U1066 ( .A1(G214), .A2(n1331), .ZN(n1256) );
NAND2_X1 U1067 ( .A1(n1292), .A2(n1354), .ZN(n1331) );
INV_X1 U1068 ( .A(G237), .ZN(n1354) );
AND2_X1 U1069 ( .A1(n1271), .A2(n1272), .ZN(n1076) );
NOR2_X1 U1070 ( .A1(n1110), .A2(n1114), .ZN(n1272) );
AND2_X1 U1071 ( .A1(G478), .A2(n1355), .ZN(n1114) );
OR2_X1 U1072 ( .A1(n1174), .A2(G902), .ZN(n1355) );
NOR3_X1 U1073 ( .A1(G478), .A2(G902), .A3(n1174), .ZN(n1110) );
XNOR2_X1 U1074 ( .A(n1356), .B(n1357), .ZN(n1174) );
NOR2_X1 U1075 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
XOR2_X1 U1076 ( .A(KEYINPUT5), .B(n1360), .Z(n1359) );
NOR2_X1 U1077 ( .A1(G107), .A2(n1361), .ZN(n1360) );
AND2_X1 U1078 ( .A1(n1361), .A2(G107), .ZN(n1358) );
XOR2_X1 U1079 ( .A(G116), .B(G122), .Z(n1361) );
XOR2_X1 U1080 ( .A(n1362), .B(n1363), .Z(n1356) );
NOR2_X1 U1081 ( .A1(KEYINPUT48), .A2(n1364), .ZN(n1363) );
XNOR2_X1 U1082 ( .A(n1365), .B(n1254), .ZN(n1364) );
INV_X1 U1083 ( .A(G134), .ZN(n1254) );
NAND3_X1 U1084 ( .A1(n1366), .A2(n1367), .A3(n1368), .ZN(n1365) );
NAND2_X1 U1085 ( .A1(G128), .A2(n1369), .ZN(n1368) );
NAND2_X1 U1086 ( .A1(KEYINPUT53), .A2(n1370), .ZN(n1367) );
NAND2_X1 U1087 ( .A1(n1371), .A2(n1315), .ZN(n1370) );
INV_X1 U1088 ( .A(G128), .ZN(n1315) );
XNOR2_X1 U1089 ( .A(KEYINPUT16), .B(n1369), .ZN(n1371) );
NAND2_X1 U1090 ( .A1(n1372), .A2(n1373), .ZN(n1366) );
INV_X1 U1091 ( .A(KEYINPUT53), .ZN(n1373) );
NAND2_X1 U1092 ( .A1(n1374), .A2(n1375), .ZN(n1372) );
OR3_X1 U1093 ( .A1(n1369), .A2(G128), .A3(KEYINPUT16), .ZN(n1375) );
NAND2_X1 U1094 ( .A1(KEYINPUT16), .A2(n1369), .ZN(n1374) );
INV_X1 U1095 ( .A(G143), .ZN(n1369) );
NAND3_X1 U1096 ( .A1(G234), .A2(n1376), .A3(G217), .ZN(n1362) );
XNOR2_X1 U1097 ( .A(KEYINPUT17), .B(n1061), .ZN(n1376) );
INV_X1 U1098 ( .A(G953), .ZN(n1061) );
INV_X1 U1099 ( .A(n1106), .ZN(n1271) );
XNOR2_X1 U1100 ( .A(n1377), .B(G475), .ZN(n1106) );
NAND2_X1 U1101 ( .A1(n1176), .A2(n1292), .ZN(n1377) );
INV_X1 U1102 ( .A(G902), .ZN(n1292) );
XNOR2_X1 U1103 ( .A(n1378), .B(n1379), .ZN(n1176) );
XOR2_X1 U1104 ( .A(n1380), .B(n1381), .Z(n1379) );
XNOR2_X1 U1105 ( .A(n1382), .B(n1383), .ZN(n1381) );
INV_X1 U1106 ( .A(G104), .ZN(n1383) );
NAND2_X1 U1107 ( .A1(n1384), .A2(KEYINPUT63), .ZN(n1382) );
XNOR2_X1 U1108 ( .A(n1385), .B(n1210), .ZN(n1384) );
INV_X1 U1109 ( .A(G125), .ZN(n1210) );
NAND2_X1 U1110 ( .A1(KEYINPUT58), .A2(n1200), .ZN(n1385) );
INV_X1 U1111 ( .A(G140), .ZN(n1200) );
XNOR2_X1 U1112 ( .A(G122), .B(G131), .ZN(n1380) );
XNOR2_X1 U1113 ( .A(n1386), .B(n1311), .ZN(n1378) );
INV_X1 U1114 ( .A(n1314), .ZN(n1311) );
XOR2_X1 U1115 ( .A(G143), .B(n1287), .Z(n1314) );
XOR2_X1 U1116 ( .A(G146), .B(KEYINPUT7), .Z(n1287) );
XOR2_X1 U1117 ( .A(n1387), .B(n1388), .Z(n1386) );
NOR2_X1 U1118 ( .A1(G113), .A2(KEYINPUT23), .ZN(n1388) );
NAND2_X1 U1119 ( .A1(n1296), .A2(G214), .ZN(n1387) );
NOR2_X1 U1120 ( .A1(G953), .A2(G237), .ZN(n1296) );
INV_X1 U1121 ( .A(G110), .ZN(n1276) );
endmodule


