//Key = 0001010011001011110111111101011000000000001110001100101010111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398;

XOR2_X1 U762 ( .A(G107), .B(n1055), .Z(G9) );
NOR3_X1 U763 ( .A1(n1056), .A2(KEYINPUT0), .A3(n1057), .ZN(n1055) );
NOR2_X1 U764 ( .A1(n1058), .A2(n1059), .ZN(G75) );
NOR4_X1 U765 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1059) );
INV_X1 U766 ( .A(G952), .ZN(n1063) );
NOR2_X1 U767 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U768 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
XOR2_X1 U769 ( .A(KEYINPUT57), .B(n1068), .Z(n1067) );
NOR3_X1 U770 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1068) );
XOR2_X1 U771 ( .A(n1072), .B(KEYINPUT43), .Z(n1066) );
NAND4_X1 U772 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1072) );
NAND3_X1 U773 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1060) );
NAND2_X1 U774 ( .A1(n1073), .A2(n1080), .ZN(n1079) );
NAND2_X1 U775 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND3_X1 U776 ( .A1(n1074), .A2(n1083), .A3(n1084), .ZN(n1082) );
NAND2_X1 U777 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NAND2_X1 U778 ( .A1(n1087), .A2(n1076), .ZN(n1086) );
NAND2_X1 U779 ( .A1(n1088), .A2(n1089), .ZN(n1085) );
NAND3_X1 U780 ( .A1(n1076), .A2(n1090), .A3(n1088), .ZN(n1081) );
NAND4_X1 U781 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1090) );
NAND3_X1 U782 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1094) );
XOR2_X1 U783 ( .A(KEYINPUT18), .B(n1074), .Z(n1096) );
NAND3_X1 U784 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1093) );
XOR2_X1 U785 ( .A(n1065), .B(KEYINPUT23), .Z(n1100) );
XOR2_X1 U786 ( .A(KEYINPUT2), .B(n1101), .Z(n1099) );
NAND2_X1 U787 ( .A1(n1084), .A2(n1102), .ZN(n1092) );
NAND2_X1 U788 ( .A1(n1074), .A2(n1103), .ZN(n1091) );
INV_X1 U789 ( .A(n1069), .ZN(n1073) );
NOR3_X1 U790 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1058) );
NOR2_X1 U791 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
INV_X1 U792 ( .A(KEYINPUT44), .ZN(n1108) );
NOR2_X1 U793 ( .A1(G953), .A2(G952), .ZN(n1107) );
NOR2_X1 U794 ( .A1(KEYINPUT44), .A2(n1109), .ZN(n1105) );
INV_X1 U795 ( .A(n1077), .ZN(n1104) );
NAND4_X1 U796 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1077) );
NOR4_X1 U797 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1113) );
XOR2_X1 U798 ( .A(n1118), .B(n1119), .Z(n1117) );
INV_X1 U799 ( .A(n1095), .ZN(n1116) );
NOR3_X1 U800 ( .A1(n1120), .A2(n1101), .A3(n1097), .ZN(n1112) );
NOR2_X1 U801 ( .A1(G472), .A2(n1121), .ZN(n1120) );
XOR2_X1 U802 ( .A(KEYINPUT5), .B(n1122), .Z(n1111) );
AND2_X1 U803 ( .A1(n1121), .A2(G472), .ZN(n1122) );
XOR2_X1 U804 ( .A(KEYINPUT24), .B(n1123), .Z(n1110) );
INV_X1 U805 ( .A(n1098), .ZN(n1123) );
XOR2_X1 U806 ( .A(n1124), .B(n1125), .Z(G72) );
XOR2_X1 U807 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U808 ( .A1(n1128), .A2(G953), .ZN(n1127) );
NOR2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1126) );
XOR2_X1 U811 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U812 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U813 ( .A(n1137), .B(n1138), .Z(n1133) );
XNOR2_X1 U814 ( .A(n1139), .B(n1140), .ZN(n1138) );
NOR2_X1 U815 ( .A1(G131), .A2(KEYINPUT34), .ZN(n1140) );
NAND2_X1 U816 ( .A1(KEYINPUT8), .A2(n1141), .ZN(n1139) );
NOR2_X1 U817 ( .A1(G900), .A2(n1142), .ZN(n1131) );
XOR2_X1 U818 ( .A(n1078), .B(KEYINPUT26), .Z(n1142) );
NOR3_X1 U819 ( .A1(n1078), .A2(KEYINPUT46), .A3(n1143), .ZN(n1124) );
AND2_X1 U820 ( .A1(G227), .A2(G900), .ZN(n1143) );
NAND2_X1 U821 ( .A1(n1144), .A2(n1145), .ZN(G69) );
NAND2_X1 U822 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND2_X1 U823 ( .A1(G953), .A2(n1148), .ZN(n1147) );
INV_X1 U824 ( .A(n1149), .ZN(n1146) );
NAND3_X1 U825 ( .A1(G953), .A2(n1150), .A3(n1149), .ZN(n1144) );
XOR2_X1 U826 ( .A(n1151), .B(n1152), .Z(n1149) );
NOR2_X1 U827 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND2_X1 U829 ( .A1(KEYINPUT59), .A2(n1157), .ZN(n1155) );
NOR2_X1 U830 ( .A1(G898), .A2(n1078), .ZN(n1153) );
NAND2_X1 U831 ( .A1(n1078), .A2(n1158), .ZN(n1151) );
NAND3_X1 U832 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1158) );
NAND2_X1 U833 ( .A1(G898), .A2(G224), .ZN(n1150) );
NOR2_X1 U834 ( .A1(n1109), .A2(n1162), .ZN(G66) );
XOR2_X1 U835 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U836 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
NOR2_X1 U837 ( .A1(n1109), .A2(n1167), .ZN(G63) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1167) );
AND2_X1 U839 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NOR2_X1 U840 ( .A1(n1118), .A2(n1166), .ZN(n1168) );
INV_X1 U841 ( .A(G478), .ZN(n1118) );
NOR2_X1 U842 ( .A1(n1109), .A2(n1172), .ZN(G60) );
XNOR2_X1 U843 ( .A(n1173), .B(n1174), .ZN(n1172) );
AND2_X1 U844 ( .A1(G475), .A2(n1175), .ZN(n1174) );
XOR2_X1 U845 ( .A(n1176), .B(n1177), .Z(G6) );
NOR2_X1 U846 ( .A1(n1178), .A2(KEYINPUT55), .ZN(n1177) );
NOR2_X1 U847 ( .A1(n1057), .A2(n1179), .ZN(n1178) );
NOR2_X1 U848 ( .A1(n1109), .A2(n1180), .ZN(G57) );
XOR2_X1 U849 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U850 ( .A(n1183), .B(n1184), .Z(n1181) );
AND2_X1 U851 ( .A1(G472), .A2(n1175), .ZN(n1184) );
NAND3_X1 U852 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1183) );
XOR2_X1 U853 ( .A(KEYINPUT20), .B(n1188), .Z(n1187) );
NOR2_X1 U854 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XNOR2_X1 U855 ( .A(KEYINPUT14), .B(n1191), .ZN(n1190) );
XNOR2_X1 U856 ( .A(n1192), .B(n1193), .ZN(n1189) );
OR2_X1 U857 ( .A1(n1194), .A2(KEYINPUT50), .ZN(n1192) );
NAND3_X1 U858 ( .A1(n1195), .A2(n1196), .A3(n1191), .ZN(n1186) );
XNOR2_X1 U859 ( .A(KEYINPUT50), .B(n1193), .ZN(n1195) );
NOR2_X1 U860 ( .A1(n1109), .A2(n1197), .ZN(G54) );
XOR2_X1 U861 ( .A(n1198), .B(n1199), .Z(n1197) );
NOR2_X1 U862 ( .A1(KEYINPUT6), .A2(n1200), .ZN(n1199) );
XOR2_X1 U863 ( .A(n1201), .B(n1202), .Z(n1200) );
NAND3_X1 U864 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1202) );
INV_X1 U865 ( .A(n1206), .ZN(n1205) );
NAND2_X1 U866 ( .A1(KEYINPUT39), .A2(n1207), .ZN(n1204) );
XOR2_X1 U867 ( .A(n1208), .B(n1196), .Z(n1207) );
NAND2_X1 U868 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND2_X1 U869 ( .A1(n1211), .A2(n1212), .ZN(n1203) );
INV_X1 U870 ( .A(KEYINPUT39), .ZN(n1212) );
NAND2_X1 U871 ( .A1(n1213), .A2(n1214), .ZN(n1201) );
NAND2_X1 U872 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XOR2_X1 U873 ( .A(n1217), .B(n1218), .Z(n1215) );
XOR2_X1 U874 ( .A(n1219), .B(KEYINPUT10), .Z(n1213) );
NAND2_X1 U875 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
XOR2_X1 U876 ( .A(G140), .B(n1218), .Z(n1221) );
NOR2_X1 U877 ( .A1(G110), .A2(KEYINPUT41), .ZN(n1218) );
NAND2_X1 U878 ( .A1(n1175), .A2(G469), .ZN(n1198) );
NOR2_X1 U879 ( .A1(n1109), .A2(n1222), .ZN(G51) );
NOR2_X1 U880 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XOR2_X1 U881 ( .A(n1225), .B(n1226), .Z(n1224) );
AND2_X1 U882 ( .A1(G210), .A2(n1175), .ZN(n1226) );
INV_X1 U883 ( .A(n1166), .ZN(n1175) );
NAND2_X1 U884 ( .A1(G902), .A2(n1061), .ZN(n1166) );
NAND4_X1 U885 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1161), .ZN(n1061) );
AND2_X1 U886 ( .A1(n1230), .A2(n1231), .ZN(n1161) );
NAND2_X1 U887 ( .A1(n1232), .A2(n1233), .ZN(n1230) );
NAND2_X1 U888 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U889 ( .A1(n1089), .A2(n1075), .ZN(n1235) );
NOR2_X1 U890 ( .A1(n1236), .A2(n1130), .ZN(n1229) );
NAND4_X1 U891 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1130) );
NOR3_X1 U892 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1240) );
INV_X1 U893 ( .A(n1244), .ZN(n1243) );
NAND2_X1 U894 ( .A1(n1087), .A2(n1245), .ZN(n1239) );
NAND2_X1 U895 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
NAND2_X1 U896 ( .A1(n1248), .A2(n1103), .ZN(n1247) );
NAND3_X1 U897 ( .A1(n1075), .A2(n1249), .A3(n1250), .ZN(n1237) );
XOR2_X1 U898 ( .A(KEYINPUT37), .B(n1102), .Z(n1249) );
INV_X1 U899 ( .A(n1160), .ZN(n1236) );
XNOR2_X1 U900 ( .A(n1129), .B(KEYINPUT31), .ZN(n1228) );
AND2_X1 U901 ( .A1(n1251), .A2(n1252), .ZN(n1129) );
XNOR2_X1 U902 ( .A(n1102), .B(KEYINPUT9), .ZN(n1251) );
XNOR2_X1 U903 ( .A(n1159), .B(KEYINPUT58), .ZN(n1227) );
AND3_X1 U904 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1159) );
NAND2_X1 U905 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND2_X1 U906 ( .A1(n1179), .A2(n1056), .ZN(n1257) );
INV_X1 U907 ( .A(n1057), .ZN(n1256) );
NAND2_X1 U908 ( .A1(n1258), .A2(n1076), .ZN(n1057) );
NOR2_X1 U909 ( .A1(KEYINPUT7), .A2(n1259), .ZN(n1225) );
XOR2_X1 U910 ( .A(n1260), .B(KEYINPUT35), .Z(n1259) );
NOR2_X1 U911 ( .A1(n1261), .A2(n1262), .ZN(n1223) );
INV_X1 U912 ( .A(KEYINPUT7), .ZN(n1262) );
XOR2_X1 U913 ( .A(KEYINPUT35), .B(n1263), .Z(n1261) );
NOR2_X1 U914 ( .A1(n1078), .A2(G952), .ZN(n1109) );
XNOR2_X1 U915 ( .A(G146), .B(n1264), .ZN(G48) );
NAND3_X1 U916 ( .A1(KEYINPUT48), .A2(n1103), .A3(n1265), .ZN(n1264) );
XOR2_X1 U917 ( .A(n1266), .B(KEYINPUT21), .Z(n1265) );
NAND2_X1 U918 ( .A1(n1248), .A2(n1087), .ZN(n1266) );
XOR2_X1 U919 ( .A(n1267), .B(n1268), .Z(G45) );
NOR2_X1 U920 ( .A1(G143), .A2(KEYINPUT51), .ZN(n1268) );
NAND2_X1 U921 ( .A1(n1252), .A2(n1102), .ZN(n1267) );
AND3_X1 U922 ( .A1(n1089), .A2(n1103), .A3(n1269), .ZN(n1252) );
AND3_X1 U923 ( .A1(n1270), .A2(n1271), .A3(n1115), .ZN(n1269) );
XOR2_X1 U924 ( .A(n1217), .B(n1238), .Z(G42) );
NAND3_X1 U925 ( .A1(n1084), .A2(n1102), .A3(n1272), .ZN(n1238) );
XOR2_X1 U926 ( .A(n1242), .B(n1273), .Z(G39) );
NOR2_X1 U927 ( .A1(KEYINPUT4), .A2(n1141), .ZN(n1273) );
INV_X1 U928 ( .A(G137), .ZN(n1141) );
AND3_X1 U929 ( .A1(n1084), .A2(n1088), .A3(n1248), .ZN(n1242) );
XOR2_X1 U930 ( .A(n1274), .B(n1275), .Z(G36) );
NAND2_X1 U931 ( .A1(KEYINPUT17), .A2(G134), .ZN(n1275) );
OR2_X1 U932 ( .A1(n1246), .A2(n1056), .ZN(n1274) );
XOR2_X1 U933 ( .A(G131), .B(n1276), .Z(G33) );
NOR3_X1 U934 ( .A1(n1246), .A2(KEYINPUT62), .A3(n1179), .ZN(n1276) );
INV_X1 U935 ( .A(n1087), .ZN(n1179) );
NAND2_X1 U936 ( .A1(n1250), .A2(n1102), .ZN(n1246) );
AND3_X1 U937 ( .A1(n1089), .A2(n1271), .A3(n1084), .ZN(n1250) );
INV_X1 U938 ( .A(n1065), .ZN(n1084) );
NAND2_X1 U939 ( .A1(n1277), .A2(n1278), .ZN(n1065) );
XOR2_X1 U940 ( .A(n1095), .B(KEYINPUT47), .Z(n1277) );
XOR2_X1 U941 ( .A(G128), .B(n1241), .Z(G30) );
AND3_X1 U942 ( .A1(n1075), .A2(n1103), .A3(n1248), .ZN(n1241) );
AND4_X1 U943 ( .A1(n1102), .A2(n1114), .A3(n1279), .A4(n1271), .ZN(n1248) );
XOR2_X1 U944 ( .A(n1280), .B(n1253), .Z(G3) );
NAND3_X1 U945 ( .A1(n1089), .A2(n1258), .A3(n1088), .ZN(n1253) );
XOR2_X1 U946 ( .A(n1281), .B(n1244), .Z(G27) );
NAND3_X1 U947 ( .A1(n1074), .A2(n1103), .A3(n1272), .ZN(n1244) );
AND4_X1 U948 ( .A1(n1282), .A2(n1087), .A3(n1114), .A4(n1271), .ZN(n1272) );
NAND2_X1 U949 ( .A1(n1069), .A2(n1283), .ZN(n1271) );
NAND4_X1 U950 ( .A1(G902), .A2(G953), .A3(n1284), .A4(n1285), .ZN(n1283) );
INV_X1 U951 ( .A(G900), .ZN(n1285) );
XOR2_X1 U952 ( .A(n1286), .B(n1160), .Z(G24) );
NAND4_X1 U953 ( .A1(n1232), .A2(n1076), .A3(n1270), .A4(n1115), .ZN(n1160) );
NOR2_X1 U954 ( .A1(n1279), .A2(n1114), .ZN(n1076) );
NAND2_X1 U955 ( .A1(n1287), .A2(n1288), .ZN(G21) );
OR2_X1 U956 ( .A1(n1289), .A2(G119), .ZN(n1288) );
NAND2_X1 U957 ( .A1(G119), .A2(n1290), .ZN(n1287) );
NAND2_X1 U958 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
NAND2_X1 U959 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
INV_X1 U960 ( .A(KEYINPUT30), .ZN(n1294) );
NAND2_X1 U961 ( .A1(KEYINPUT30), .A2(n1289), .ZN(n1291) );
NAND2_X1 U962 ( .A1(KEYINPUT3), .A2(n1293), .ZN(n1289) );
AND4_X1 U963 ( .A1(n1295), .A2(n1074), .A3(n1103), .A4(n1296), .ZN(n1293) );
XOR2_X1 U964 ( .A(KEYINPUT29), .B(n1297), .Z(n1296) );
AND2_X1 U965 ( .A1(n1298), .A2(n1069), .ZN(n1297) );
INV_X1 U966 ( .A(n1234), .ZN(n1295) );
NAND3_X1 U967 ( .A1(n1114), .A2(n1279), .A3(n1088), .ZN(n1234) );
XOR2_X1 U968 ( .A(n1299), .B(n1300), .Z(G18) );
XOR2_X1 U969 ( .A(KEYINPUT60), .B(G116), .Z(n1300) );
NAND4_X1 U970 ( .A1(KEYINPUT42), .A2(n1089), .A3(n1232), .A4(n1075), .ZN(n1299) );
INV_X1 U971 ( .A(n1056), .ZN(n1075) );
NAND2_X1 U972 ( .A1(n1301), .A2(n1270), .ZN(n1056) );
XOR2_X1 U973 ( .A(n1302), .B(n1231), .Z(G15) );
NAND3_X1 U974 ( .A1(n1232), .A2(n1087), .A3(n1089), .ZN(n1231) );
NOR2_X1 U975 ( .A1(n1114), .A2(n1282), .ZN(n1089) );
NOR2_X1 U976 ( .A1(n1270), .A2(n1301), .ZN(n1087) );
AND2_X1 U977 ( .A1(n1074), .A2(n1303), .ZN(n1232) );
INV_X1 U978 ( .A(n1070), .ZN(n1074) );
NAND2_X1 U979 ( .A1(n1304), .A2(n1305), .ZN(n1070) );
XOR2_X1 U980 ( .A(n1098), .B(KEYINPUT28), .Z(n1304) );
XOR2_X1 U981 ( .A(n1254), .B(n1306), .Z(G12) );
NAND2_X1 U982 ( .A1(KEYINPUT52), .A2(G110), .ZN(n1306) );
NAND2_X1 U983 ( .A1(n1307), .A2(n1258), .ZN(n1254) );
AND2_X1 U984 ( .A1(n1102), .A2(n1303), .ZN(n1258) );
AND2_X1 U985 ( .A1(n1103), .A2(n1308), .ZN(n1303) );
NAND2_X1 U986 ( .A1(n1298), .A2(n1069), .ZN(n1308) );
NAND3_X1 U987 ( .A1(n1284), .A2(n1078), .A3(G952), .ZN(n1069) );
NAND4_X1 U988 ( .A1(n1309), .A2(G902), .A3(n1284), .A4(n1310), .ZN(n1298) );
INV_X1 U989 ( .A(G898), .ZN(n1310) );
NAND2_X1 U990 ( .A1(G237), .A2(G234), .ZN(n1284) );
XOR2_X1 U991 ( .A(n1078), .B(KEYINPUT63), .Z(n1309) );
NOR2_X1 U992 ( .A1(n1095), .A2(n1097), .ZN(n1103) );
INV_X1 U993 ( .A(n1278), .ZN(n1097) );
NAND2_X1 U994 ( .A1(G214), .A2(n1311), .ZN(n1278) );
XOR2_X1 U995 ( .A(n1312), .B(n1313), .Z(n1095) );
AND2_X1 U996 ( .A1(n1311), .A2(G210), .ZN(n1313) );
NAND2_X1 U997 ( .A1(n1314), .A2(n1315), .ZN(n1311) );
XNOR2_X1 U998 ( .A(G237), .B(KEYINPUT40), .ZN(n1314) );
NAND2_X1 U999 ( .A1(n1263), .A2(n1315), .ZN(n1312) );
INV_X1 U1000 ( .A(n1260), .ZN(n1263) );
XOR2_X1 U1001 ( .A(n1316), .B(n1317), .Z(n1260) );
XOR2_X1 U1002 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1003 ( .A(KEYINPUT25), .B(n1320), .Z(n1319) );
NOR2_X1 U1004 ( .A1(G953), .A2(n1148), .ZN(n1318) );
INV_X1 U1005 ( .A(G224), .ZN(n1148) );
XOR2_X1 U1006 ( .A(n1321), .B(n1322), .Z(n1316) );
NAND2_X1 U1007 ( .A1(n1323), .A2(n1324), .ZN(n1321) );
NAND2_X1 U1008 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
INV_X1 U1009 ( .A(n1156), .ZN(n1326) );
XOR2_X1 U1010 ( .A(KEYINPUT32), .B(n1157), .Z(n1325) );
NAND2_X1 U1011 ( .A1(n1156), .A2(n1327), .ZN(n1323) );
XOR2_X1 U1012 ( .A(KEYINPUT16), .B(n1157), .Z(n1327) );
XNOR2_X1 U1013 ( .A(n1328), .B(n1329), .ZN(n1157) );
XOR2_X1 U1014 ( .A(G113), .B(n1330), .Z(n1329) );
NOR2_X1 U1015 ( .A1(G101), .A2(KEYINPUT11), .ZN(n1330) );
XNOR2_X1 U1016 ( .A(n1331), .B(n1332), .ZN(n1328) );
NOR2_X1 U1017 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
NOR3_X1 U1018 ( .A1(KEYINPUT22), .A2(G107), .A3(n1176), .ZN(n1334) );
INV_X1 U1019 ( .A(G104), .ZN(n1176) );
NOR2_X1 U1020 ( .A1(n1335), .A2(n1336), .ZN(n1333) );
INV_X1 U1021 ( .A(KEYINPUT22), .ZN(n1336) );
XOR2_X1 U1022 ( .A(G110), .B(G122), .Z(n1156) );
NOR2_X1 U1023 ( .A1(n1098), .A2(n1101), .ZN(n1102) );
INV_X1 U1024 ( .A(n1305), .ZN(n1101) );
NAND2_X1 U1025 ( .A1(G221), .A2(n1337), .ZN(n1305) );
XOR2_X1 U1026 ( .A(n1338), .B(G469), .Z(n1098) );
NAND2_X1 U1027 ( .A1(n1339), .A2(n1315), .ZN(n1338) );
XOR2_X1 U1028 ( .A(n1340), .B(n1341), .Z(n1339) );
XOR2_X1 U1029 ( .A(n1342), .B(n1220), .Z(n1341) );
INV_X1 U1030 ( .A(n1216), .ZN(n1220) );
NAND2_X1 U1031 ( .A1(G227), .A2(n1078), .ZN(n1216) );
NOR2_X1 U1032 ( .A1(n1206), .A2(n1211), .ZN(n1342) );
NAND2_X1 U1033 ( .A1(n1343), .A2(n1344), .ZN(n1211) );
NAND3_X1 U1034 ( .A1(n1210), .A2(n1196), .A3(n1345), .ZN(n1344) );
NAND2_X1 U1035 ( .A1(n1346), .A2(n1209), .ZN(n1343) );
XOR2_X1 U1036 ( .A(n1196), .B(n1210), .Z(n1346) );
NOR3_X1 U1037 ( .A1(n1210), .A2(n1209), .A3(n1196), .ZN(n1206) );
INV_X1 U1038 ( .A(n1345), .ZN(n1209) );
XOR2_X1 U1039 ( .A(n1280), .B(n1335), .Z(n1345) );
XOR2_X1 U1040 ( .A(G104), .B(G107), .Z(n1335) );
INV_X1 U1041 ( .A(G101), .ZN(n1280) );
XNOR2_X1 U1042 ( .A(n1347), .B(n1135), .ZN(n1210) );
XOR2_X1 U1043 ( .A(G146), .B(KEYINPUT36), .Z(n1135) );
XNOR2_X1 U1044 ( .A(G128), .B(G143), .ZN(n1347) );
XOR2_X1 U1045 ( .A(G140), .B(G110), .Z(n1340) );
INV_X1 U1046 ( .A(n1071), .ZN(n1307) );
NAND3_X1 U1047 ( .A1(n1282), .A2(n1114), .A3(n1088), .ZN(n1071) );
NOR2_X1 U1048 ( .A1(n1115), .A2(n1270), .ZN(n1088) );
XOR2_X1 U1049 ( .A(n1348), .B(G478), .Z(n1270) );
NAND2_X1 U1050 ( .A1(KEYINPUT27), .A2(n1119), .ZN(n1348) );
NAND2_X1 U1051 ( .A1(n1315), .A2(n1349), .ZN(n1119) );
NAND2_X1 U1052 ( .A1(n1170), .A2(n1171), .ZN(n1349) );
NAND2_X1 U1053 ( .A1(n1350), .A2(n1351), .ZN(n1171) );
NAND3_X1 U1054 ( .A1(n1352), .A2(n1078), .A3(G217), .ZN(n1351) );
XOR2_X1 U1055 ( .A(n1353), .B(n1354), .Z(n1350) );
NAND4_X1 U1056 ( .A1(G217), .A2(n1355), .A3(n1352), .A4(n1078), .ZN(n1170) );
XOR2_X1 U1057 ( .A(G234), .B(KEYINPUT53), .Z(n1352) );
XOR2_X1 U1058 ( .A(n1356), .B(n1354), .Z(n1355) );
XOR2_X1 U1059 ( .A(n1136), .B(n1357), .Z(n1354) );
NOR2_X1 U1060 ( .A1(G128), .A2(KEYINPUT45), .ZN(n1357) );
XOR2_X1 U1061 ( .A(G134), .B(G143), .Z(n1136) );
INV_X1 U1062 ( .A(n1353), .ZN(n1356) );
XNOR2_X1 U1063 ( .A(G107), .B(n1358), .ZN(n1353) );
XOR2_X1 U1064 ( .A(G122), .B(G116), .Z(n1358) );
INV_X1 U1065 ( .A(n1301), .ZN(n1115) );
XOR2_X1 U1066 ( .A(n1359), .B(G475), .Z(n1301) );
NAND2_X1 U1067 ( .A1(n1173), .A2(n1315), .ZN(n1359) );
XNOR2_X1 U1068 ( .A(n1360), .B(n1361), .ZN(n1173) );
XOR2_X1 U1069 ( .A(n1362), .B(n1363), .Z(n1361) );
XOR2_X1 U1070 ( .A(n1364), .B(n1365), .Z(n1363) );
NOR2_X1 U1071 ( .A1(KEYINPUT38), .A2(G146), .ZN(n1365) );
NAND2_X1 U1072 ( .A1(n1366), .A2(n1367), .ZN(n1364) );
OR2_X1 U1073 ( .A1(n1368), .A2(G104), .ZN(n1367) );
XOR2_X1 U1074 ( .A(n1369), .B(KEYINPUT33), .Z(n1366) );
NAND2_X1 U1075 ( .A1(G104), .A2(n1368), .ZN(n1369) );
XOR2_X1 U1076 ( .A(n1302), .B(n1286), .Z(n1368) );
INV_X1 U1077 ( .A(G122), .ZN(n1286) );
NAND4_X1 U1078 ( .A1(KEYINPUT15), .A2(n1370), .A3(n1371), .A4(n1372), .ZN(n1362) );
NAND4_X1 U1079 ( .A1(n1373), .A2(n1374), .A3(KEYINPUT54), .A4(n1375), .ZN(n1372) );
INV_X1 U1080 ( .A(n1376), .ZN(n1375) );
NAND2_X1 U1081 ( .A1(n1376), .A2(n1377), .ZN(n1371) );
NAND3_X1 U1082 ( .A1(n1378), .A2(n1374), .A3(G214), .ZN(n1377) );
INV_X1 U1083 ( .A(KEYINPUT13), .ZN(n1374) );
XNOR2_X1 U1084 ( .A(G143), .B(KEYINPUT56), .ZN(n1376) );
OR2_X1 U1085 ( .A1(n1373), .A2(KEYINPUT54), .ZN(n1370) );
AND2_X1 U1086 ( .A1(G214), .A2(n1378), .ZN(n1373) );
XOR2_X1 U1087 ( .A(n1281), .B(n1379), .Z(n1360) );
XOR2_X1 U1088 ( .A(G140), .B(G131), .Z(n1379) );
INV_X1 U1089 ( .A(G125), .ZN(n1281) );
XNOR2_X1 U1090 ( .A(n1380), .B(n1381), .ZN(n1114) );
NOR2_X1 U1091 ( .A1(n1382), .A2(n1165), .ZN(n1381) );
INV_X1 U1092 ( .A(G217), .ZN(n1165) );
XOR2_X1 U1093 ( .A(n1337), .B(KEYINPUT19), .Z(n1382) );
NAND2_X1 U1094 ( .A1(G234), .A2(n1315), .ZN(n1337) );
OR2_X1 U1095 ( .A1(n1164), .A2(G902), .ZN(n1380) );
XNOR2_X1 U1096 ( .A(n1383), .B(n1384), .ZN(n1164) );
XOR2_X1 U1097 ( .A(G110), .B(n1385), .Z(n1384) );
XOR2_X1 U1098 ( .A(G137), .B(G119), .Z(n1385) );
XNOR2_X1 U1099 ( .A(n1137), .B(n1386), .ZN(n1383) );
XOR2_X1 U1100 ( .A(n1387), .B(n1388), .Z(n1386) );
AND3_X1 U1101 ( .A1(G221), .A2(n1078), .A3(G234), .ZN(n1388) );
INV_X1 U1102 ( .A(G953), .ZN(n1078) );
NOR2_X1 U1103 ( .A1(KEYINPUT1), .A2(G146), .ZN(n1387) );
XNOR2_X1 U1104 ( .A(n1217), .B(n1322), .ZN(n1137) );
XOR2_X1 U1105 ( .A(G125), .B(G128), .Z(n1322) );
INV_X1 U1106 ( .A(G140), .ZN(n1217) );
INV_X1 U1107 ( .A(n1279), .ZN(n1282) );
XNOR2_X1 U1108 ( .A(n1121), .B(G472), .ZN(n1279) );
NAND2_X1 U1109 ( .A1(n1389), .A2(n1315), .ZN(n1121) );
INV_X1 U1110 ( .A(G902), .ZN(n1315) );
XNOR2_X1 U1111 ( .A(n1390), .B(n1182), .ZN(n1389) );
XNOR2_X1 U1112 ( .A(n1391), .B(G101), .ZN(n1182) );
NAND2_X1 U1113 ( .A1(G210), .A2(n1378), .ZN(n1391) );
NOR2_X1 U1114 ( .A1(G953), .A2(G237), .ZN(n1378) );
NAND3_X1 U1115 ( .A1(n1392), .A2(n1393), .A3(n1185), .ZN(n1390) );
NAND3_X1 U1116 ( .A1(n1191), .A2(n1194), .A3(n1193), .ZN(n1185) );
OR3_X1 U1117 ( .A1(n1191), .A2(n1193), .A3(n1196), .ZN(n1393) );
NAND2_X1 U1118 ( .A1(n1394), .A2(n1196), .ZN(n1392) );
INV_X1 U1119 ( .A(n1194), .ZN(n1196) );
XOR2_X1 U1120 ( .A(n1395), .B(G131), .Z(n1194) );
NAND2_X1 U1121 ( .A1(KEYINPUT12), .A2(n1396), .ZN(n1395) );
XOR2_X1 U1122 ( .A(G137), .B(G134), .Z(n1396) );
XOR2_X1 U1123 ( .A(n1191), .B(n1193), .Z(n1394) );
XNOR2_X1 U1124 ( .A(G128), .B(n1320), .ZN(n1193) );
NOR2_X1 U1125 ( .A1(KEYINPUT61), .A2(n1397), .ZN(n1320) );
XOR2_X1 U1126 ( .A(G146), .B(G143), .Z(n1397) );
XOR2_X1 U1127 ( .A(n1398), .B(n1331), .Z(n1191) );
XOR2_X1 U1128 ( .A(G116), .B(G119), .Z(n1331) );
NAND2_X1 U1129 ( .A1(KEYINPUT49), .A2(n1302), .ZN(n1398) );
INV_X1 U1130 ( .A(G113), .ZN(n1302) );
endmodule


