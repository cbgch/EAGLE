//Key = 1101101111100010011010100011100111111000110110101100100011000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395;

XNOR2_X1 U763 ( .A(n1062), .B(n1063), .ZN(G9) );
NOR2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(G75) );
NOR3_X1 U765 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
NAND3_X1 U766 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1066) );
NAND2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U768 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND3_X1 U769 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NAND2_X1 U770 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NAND2_X1 U771 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U772 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U773 ( .A1(n1085), .A2(n1086), .ZN(n1079) );
OR2_X1 U774 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND3_X1 U775 ( .A1(n1081), .A2(n1089), .A3(n1085), .ZN(n1074) );
NAND3_X1 U776 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
NAND2_X1 U777 ( .A1(n1076), .A2(n1093), .ZN(n1092) );
NAND3_X1 U778 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1091) );
XNOR2_X1 U779 ( .A(n1076), .B(KEYINPUT56), .ZN(n1096) );
NAND2_X1 U780 ( .A1(n1078), .A2(n1097), .ZN(n1090) );
NAND2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
INV_X1 U783 ( .A(n1102), .ZN(n1072) );
AND3_X1 U784 ( .A1(n1069), .A2(n1070), .A3(n1103), .ZN(n1064) );
NAND4_X1 U785 ( .A1(n1094), .A2(n1076), .A3(n1104), .A4(n1105), .ZN(n1069) );
NOR4_X1 U786 ( .A1(n1095), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1105) );
XNOR2_X1 U787 ( .A(n1109), .B(n1110), .ZN(n1108) );
NAND2_X1 U788 ( .A1(KEYINPUT4), .A2(n1111), .ZN(n1109) );
NOR3_X1 U789 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1104) );
AND3_X1 U790 ( .A1(KEYINPUT62), .A2(n1115), .A3(n1116), .ZN(n1114) );
NOR2_X1 U791 ( .A1(KEYINPUT62), .A2(n1116), .ZN(n1113) );
XOR2_X1 U792 ( .A(KEYINPUT60), .B(n1117), .Z(n1112) );
XOR2_X1 U793 ( .A(n1118), .B(n1119), .Z(G72) );
NOR2_X1 U794 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U795 ( .A(n1122), .B(KEYINPUT57), .Z(n1121) );
NAND3_X1 U796 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1122) );
INV_X1 U797 ( .A(n1126), .ZN(n1123) );
NOR2_X1 U798 ( .A1(n1125), .A2(n1124), .ZN(n1120) );
NAND3_X1 U799 ( .A1(n1127), .A2(n1128), .A3(n1070), .ZN(n1124) );
OR4_X1 U800 ( .A1(n1129), .A2(n1083), .A3(n1130), .A4(KEYINPUT46), .ZN(n1128) );
NAND2_X1 U801 ( .A1(KEYINPUT46), .A2(n1131), .ZN(n1127) );
INV_X1 U802 ( .A(n1068), .ZN(n1131) );
XOR2_X1 U803 ( .A(n1132), .B(n1133), .Z(n1125) );
XOR2_X1 U804 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U805 ( .A1(KEYINPUT5), .A2(n1136), .ZN(n1134) );
XNOR2_X1 U806 ( .A(n1137), .B(n1138), .ZN(n1132) );
NAND2_X1 U807 ( .A1(n1139), .A2(KEYINPUT43), .ZN(n1138) );
XNOR2_X1 U808 ( .A(G134), .B(n1140), .ZN(n1139) );
XNOR2_X1 U809 ( .A(KEYINPUT31), .B(n1141), .ZN(n1140) );
INV_X1 U810 ( .A(G137), .ZN(n1141) );
NAND2_X1 U811 ( .A1(n1142), .A2(KEYINPUT33), .ZN(n1137) );
XNOR2_X1 U812 ( .A(G128), .B(n1143), .ZN(n1142) );
NAND2_X1 U813 ( .A1(G953), .A2(n1144), .ZN(n1118) );
NAND2_X1 U814 ( .A1(G900), .A2(G227), .ZN(n1144) );
XOR2_X1 U815 ( .A(n1145), .B(n1146), .Z(G69) );
XOR2_X1 U816 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U817 ( .A1(n1149), .A2(n1070), .ZN(n1148) );
NOR2_X1 U818 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND2_X1 U819 ( .A1(n1152), .A2(n1153), .ZN(n1147) );
NAND2_X1 U820 ( .A1(G953), .A2(n1151), .ZN(n1153) );
XNOR2_X1 U821 ( .A(n1154), .B(n1155), .ZN(n1152) );
NAND2_X1 U822 ( .A1(KEYINPUT6), .A2(n1156), .ZN(n1154) );
XOR2_X1 U823 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U824 ( .A1(KEYINPUT40), .A2(n1159), .ZN(n1157) );
NAND2_X1 U825 ( .A1(n1070), .A2(n1067), .ZN(n1145) );
NOR2_X1 U826 ( .A1(n1160), .A2(n1161), .ZN(G66) );
XNOR2_X1 U827 ( .A(n1162), .B(n1163), .ZN(n1161) );
NOR2_X1 U828 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NOR2_X1 U829 ( .A1(n1160), .A2(n1166), .ZN(G63) );
XOR2_X1 U830 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U831 ( .A1(n1110), .A2(n1165), .ZN(n1168) );
INV_X1 U832 ( .A(G478), .ZN(n1110) );
NAND2_X1 U833 ( .A1(n1169), .A2(KEYINPUT27), .ZN(n1167) );
XOR2_X1 U834 ( .A(n1170), .B(KEYINPUT14), .Z(n1169) );
NOR2_X1 U835 ( .A1(n1160), .A2(n1171), .ZN(G60) );
XOR2_X1 U836 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U837 ( .A1(n1174), .A2(n1165), .ZN(n1172) );
XOR2_X1 U838 ( .A(G104), .B(n1175), .Z(G6) );
NOR2_X1 U839 ( .A1(n1160), .A2(n1176), .ZN(G57) );
XOR2_X1 U840 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U841 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U842 ( .A(n1181), .B(n1182), .Z(n1177) );
NOR2_X1 U843 ( .A1(n1183), .A2(n1165), .ZN(n1182) );
NOR3_X1 U844 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(G54) );
AND2_X1 U845 ( .A1(KEYINPUT35), .A2(n1160), .ZN(n1186) );
NOR3_X1 U846 ( .A1(KEYINPUT35), .A2(n1070), .A3(n1103), .ZN(n1185) );
INV_X1 U847 ( .A(G952), .ZN(n1103) );
XOR2_X1 U848 ( .A(n1187), .B(n1188), .Z(n1184) );
XOR2_X1 U849 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U850 ( .A1(n1191), .A2(n1165), .ZN(n1190) );
INV_X1 U851 ( .A(G469), .ZN(n1191) );
NOR2_X1 U852 ( .A1(n1192), .A2(n1193), .ZN(n1189) );
XOR2_X1 U853 ( .A(n1194), .B(KEYINPUT1), .Z(n1193) );
INV_X1 U854 ( .A(n1195), .ZN(n1192) );
NOR2_X1 U855 ( .A1(n1160), .A2(n1196), .ZN(G51) );
XOR2_X1 U856 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U857 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U858 ( .A1(n1201), .A2(KEYINPUT53), .ZN(n1199) );
XOR2_X1 U859 ( .A(n1202), .B(n1203), .Z(n1197) );
NOR2_X1 U860 ( .A1(n1204), .A2(n1165), .ZN(n1203) );
NAND2_X1 U861 ( .A1(G902), .A2(n1205), .ZN(n1165) );
NAND2_X1 U862 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
INV_X1 U863 ( .A(n1067), .ZN(n1207) );
NAND4_X1 U864 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1067) );
NOR4_X1 U865 ( .A1(n1175), .A2(n1063), .A3(n1212), .A4(n1213), .ZN(n1211) );
AND3_X1 U866 ( .A1(n1081), .A2(n1214), .A3(n1215), .ZN(n1063) );
AND3_X1 U867 ( .A1(n1215), .A2(n1081), .A3(n1216), .ZN(n1175) );
NOR4_X1 U868 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1210) );
AND4_X1 U869 ( .A1(KEYINPUT47), .A2(n1221), .A3(n1222), .A4(n1081), .ZN(n1220) );
NOR2_X1 U870 ( .A1(KEYINPUT47), .A2(n1223), .ZN(n1219) );
NOR4_X1 U871 ( .A1(KEYINPUT36), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1218) );
NAND3_X1 U872 ( .A1(n1227), .A2(n1098), .A3(n1214), .ZN(n1224) );
AND2_X1 U873 ( .A1(KEYINPUT36), .A2(n1228), .ZN(n1217) );
XOR2_X1 U874 ( .A(n1068), .B(KEYINPUT49), .Z(n1206) );
NAND4_X1 U875 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1068) );
NOR2_X1 U876 ( .A1(n1233), .A2(n1130), .ZN(n1232) );
NAND4_X1 U877 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1130) );
NAND4_X1 U878 ( .A1(n1085), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1236) );
XNOR2_X1 U879 ( .A(KEYINPUT59), .B(n1241), .ZN(n1240) );
NAND2_X1 U880 ( .A1(n1242), .A2(n1243), .ZN(n1235) );
NAND2_X1 U881 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
NAND4_X1 U882 ( .A1(KEYINPUT19), .A2(n1216), .A3(n1246), .A4(n1239), .ZN(n1245) );
NOR2_X1 U883 ( .A1(n1093), .A2(n1247), .ZN(n1246) );
XNOR2_X1 U884 ( .A(KEYINPUT44), .B(n1248), .ZN(n1244) );
OR2_X1 U885 ( .A1(n1249), .A2(KEYINPUT19), .ZN(n1234) );
NOR2_X1 U886 ( .A1(n1083), .A2(n1129), .ZN(n1233) );
NOR3_X1 U887 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1202) );
NOR2_X1 U888 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NOR3_X1 U889 ( .A1(G125), .A2(KEYINPUT45), .A3(n1255), .ZN(n1251) );
INV_X1 U890 ( .A(n1253), .ZN(n1255) );
NOR2_X1 U891 ( .A1(KEYINPUT30), .A2(n1256), .ZN(n1253) );
AND2_X1 U892 ( .A1(n1256), .A2(KEYINPUT45), .ZN(n1250) );
NOR2_X1 U893 ( .A1(n1070), .A2(G952), .ZN(n1160) );
XNOR2_X1 U894 ( .A(G146), .B(n1249), .ZN(G48) );
NAND4_X1 U895 ( .A1(n1216), .A2(n1238), .A3(n1239), .A4(n1242), .ZN(n1249) );
XOR2_X1 U896 ( .A(G143), .B(n1257), .Z(G45) );
NOR2_X1 U897 ( .A1(n1098), .A2(n1248), .ZN(n1257) );
NAND3_X1 U898 ( .A1(n1087), .A2(n1238), .A3(n1258), .ZN(n1248) );
XNOR2_X1 U899 ( .A(G140), .B(n1237), .ZN(G42) );
NAND2_X1 U900 ( .A1(n1088), .A2(n1259), .ZN(n1237) );
XNOR2_X1 U901 ( .A(G137), .B(n1260), .ZN(G39) );
NAND3_X1 U902 ( .A1(n1261), .A2(n1085), .A3(n1262), .ZN(n1260) );
NOR3_X1 U903 ( .A1(n1263), .A2(KEYINPUT16), .A3(n1264), .ZN(n1262) );
XNOR2_X1 U904 ( .A(n1076), .B(KEYINPUT3), .ZN(n1261) );
XNOR2_X1 U905 ( .A(n1231), .B(n1265), .ZN(G36) );
NOR2_X1 U906 ( .A1(KEYINPUT37), .A2(n1266), .ZN(n1265) );
NAND4_X1 U907 ( .A1(n1087), .A2(n1238), .A3(n1076), .A4(n1214), .ZN(n1231) );
INV_X1 U908 ( .A(n1241), .ZN(n1076) );
INV_X1 U909 ( .A(n1263), .ZN(n1238) );
XNOR2_X1 U910 ( .A(G131), .B(n1229), .ZN(G33) );
NAND2_X1 U911 ( .A1(n1087), .A2(n1259), .ZN(n1229) );
NOR3_X1 U912 ( .A1(n1263), .A2(n1241), .A3(n1083), .ZN(n1259) );
NAND2_X1 U913 ( .A1(n1101), .A2(n1267), .ZN(n1241) );
NAND2_X1 U914 ( .A1(n1093), .A2(n1268), .ZN(n1263) );
XNOR2_X1 U915 ( .A(G128), .B(n1230), .ZN(G30) );
NAND4_X1 U916 ( .A1(n1239), .A2(n1214), .A3(n1269), .A4(n1242), .ZN(n1230) );
NOR2_X1 U917 ( .A1(n1247), .A2(n1270), .ZN(n1269) );
INV_X1 U918 ( .A(n1268), .ZN(n1247) );
INV_X1 U919 ( .A(n1084), .ZN(n1214) );
XNOR2_X1 U920 ( .A(G101), .B(n1208), .ZN(G3) );
NAND3_X1 U921 ( .A1(n1087), .A2(n1215), .A3(n1085), .ZN(n1208) );
INV_X1 U922 ( .A(n1225), .ZN(n1087) );
NAND3_X1 U923 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(G27) );
NAND2_X1 U924 ( .A1(n1274), .A2(n1254), .ZN(n1273) );
NAND2_X1 U925 ( .A1(KEYINPUT54), .A2(n1275), .ZN(n1272) );
NAND2_X1 U926 ( .A1(G125), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U927 ( .A(n1277), .B(n1274), .ZN(n1276) );
NAND2_X1 U928 ( .A1(n1278), .A2(n1279), .ZN(n1271) );
INV_X1 U929 ( .A(KEYINPUT54), .ZN(n1279) );
NAND2_X1 U930 ( .A1(n1280), .A2(n1281), .ZN(n1278) );
NAND2_X1 U931 ( .A1(n1274), .A2(n1277), .ZN(n1281) );
OR3_X1 U932 ( .A1(n1254), .A2(n1274), .A3(n1277), .ZN(n1280) );
INV_X1 U933 ( .A(KEYINPUT48), .ZN(n1277) );
NOR2_X1 U934 ( .A1(n1129), .A2(n1282), .ZN(n1274) );
XNOR2_X1 U935 ( .A(KEYINPUT21), .B(n1216), .ZN(n1282) );
NAND4_X1 U936 ( .A1(n1078), .A2(n1088), .A3(n1242), .A4(n1268), .ZN(n1129) );
NAND2_X1 U937 ( .A1(n1102), .A2(n1283), .ZN(n1268) );
NAND3_X1 U938 ( .A1(G902), .A2(n1284), .A3(n1126), .ZN(n1283) );
NOR2_X1 U939 ( .A1(n1070), .A2(G900), .ZN(n1126) );
INV_X1 U940 ( .A(n1226), .ZN(n1078) );
XNOR2_X1 U941 ( .A(G122), .B(n1223), .ZN(G24) );
NAND3_X1 U942 ( .A1(n1258), .A2(n1081), .A3(n1221), .ZN(n1223) );
NOR2_X1 U943 ( .A1(n1285), .A2(n1117), .ZN(n1081) );
INV_X1 U944 ( .A(n1222), .ZN(n1258) );
NAND2_X1 U945 ( .A1(n1286), .A2(n1287), .ZN(n1222) );
XNOR2_X1 U946 ( .A(KEYINPUT34), .B(n1288), .ZN(n1287) );
XNOR2_X1 U947 ( .A(G119), .B(n1209), .ZN(G21) );
NAND3_X1 U948 ( .A1(n1085), .A2(n1239), .A3(n1221), .ZN(n1209) );
INV_X1 U949 ( .A(n1264), .ZN(n1239) );
NAND2_X1 U950 ( .A1(n1117), .A2(n1285), .ZN(n1264) );
INV_X1 U951 ( .A(n1289), .ZN(n1285) );
XOR2_X1 U952 ( .A(n1228), .B(n1290), .Z(G18) );
NOR2_X1 U953 ( .A1(KEYINPUT23), .A2(n1291), .ZN(n1290) );
NOR3_X1 U954 ( .A1(n1225), .A2(n1084), .A3(n1292), .ZN(n1228) );
NAND2_X1 U955 ( .A1(n1293), .A2(n1294), .ZN(n1084) );
XOR2_X1 U956 ( .A(n1286), .B(KEYINPUT24), .Z(n1293) );
XOR2_X1 U957 ( .A(G113), .B(n1213), .Z(G15) );
NOR3_X1 U958 ( .A1(n1225), .A2(n1083), .A3(n1292), .ZN(n1213) );
INV_X1 U959 ( .A(n1221), .ZN(n1292) );
NOR3_X1 U960 ( .A1(n1098), .A2(n1295), .A3(n1226), .ZN(n1221) );
NAND2_X1 U961 ( .A1(n1094), .A2(n1296), .ZN(n1226) );
XOR2_X1 U962 ( .A(KEYINPUT28), .B(n1095), .Z(n1296) );
INV_X1 U963 ( .A(n1216), .ZN(n1083) );
NOR2_X1 U964 ( .A1(n1294), .A2(n1286), .ZN(n1216) );
NAND2_X1 U965 ( .A1(n1289), .A2(n1117), .ZN(n1225) );
XNOR2_X1 U966 ( .A(n1297), .B(n1212), .ZN(G12) );
AND3_X1 U967 ( .A1(n1088), .A2(n1215), .A3(n1085), .ZN(n1212) );
NOR2_X1 U968 ( .A1(n1286), .A2(n1288), .ZN(n1085) );
INV_X1 U969 ( .A(n1294), .ZN(n1288) );
XNOR2_X1 U970 ( .A(n1107), .B(KEYINPUT55), .ZN(n1294) );
XOR2_X1 U971 ( .A(n1298), .B(n1299), .Z(n1107) );
XNOR2_X1 U972 ( .A(KEYINPUT61), .B(n1174), .ZN(n1299) );
INV_X1 U973 ( .A(G475), .ZN(n1174) );
OR2_X1 U974 ( .A1(n1173), .A2(G902), .ZN(n1298) );
XNOR2_X1 U975 ( .A(n1300), .B(n1301), .ZN(n1173) );
XOR2_X1 U976 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U977 ( .A(G131), .B(G122), .Z(n1303) );
XNOR2_X1 U978 ( .A(n1304), .B(G143), .ZN(n1302) );
XOR2_X1 U979 ( .A(n1305), .B(n1306), .Z(n1300) );
XOR2_X1 U980 ( .A(G113), .B(G104), .Z(n1306) );
XNOR2_X1 U981 ( .A(n1136), .B(n1307), .ZN(n1305) );
AND2_X1 U982 ( .A1(G214), .A2(n1308), .ZN(n1307) );
XOR2_X1 U983 ( .A(G125), .B(n1309), .Z(n1136) );
XOR2_X1 U984 ( .A(n1111), .B(n1310), .Z(n1286) );
NOR2_X1 U985 ( .A1(G478), .A2(KEYINPUT12), .ZN(n1310) );
OR2_X1 U986 ( .A1(n1170), .A2(G902), .ZN(n1111) );
NAND3_X1 U987 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1170) );
NAND2_X1 U988 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
INV_X1 U989 ( .A(KEYINPUT63), .ZN(n1315) );
NAND3_X1 U990 ( .A1(KEYINPUT63), .A2(n1316), .A3(n1317), .ZN(n1312) );
OR2_X1 U991 ( .A1(n1317), .A2(n1316), .ZN(n1311) );
NOR2_X1 U992 ( .A1(KEYINPUT51), .A2(n1314), .ZN(n1316) );
NAND3_X1 U993 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1314) );
NAND2_X1 U994 ( .A1(KEYINPUT2), .A2(n1321), .ZN(n1320) );
OR3_X1 U995 ( .A1(n1321), .A2(KEYINPUT2), .A3(n1322), .ZN(n1319) );
NAND2_X1 U996 ( .A1(n1322), .A2(n1323), .ZN(n1318) );
NAND2_X1 U997 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
INV_X1 U998 ( .A(KEYINPUT2), .ZN(n1325) );
XOR2_X1 U999 ( .A(KEYINPUT41), .B(n1321), .Z(n1324) );
XOR2_X1 U1000 ( .A(G143), .B(n1326), .Z(n1321) );
XNOR2_X1 U1001 ( .A(G107), .B(n1327), .ZN(n1322) );
XNOR2_X1 U1002 ( .A(G122), .B(n1291), .ZN(n1327) );
NAND3_X1 U1003 ( .A1(G234), .A2(n1070), .A3(G217), .ZN(n1317) );
NOR3_X1 U1004 ( .A1(n1270), .A2(n1295), .A3(n1098), .ZN(n1215) );
INV_X1 U1005 ( .A(n1242), .ZN(n1098) );
NOR2_X1 U1006 ( .A1(n1101), .A2(n1100), .ZN(n1242) );
INV_X1 U1007 ( .A(n1267), .ZN(n1100) );
NAND2_X1 U1008 ( .A1(G214), .A2(n1328), .ZN(n1267) );
XNOR2_X1 U1009 ( .A(n1329), .B(n1204), .ZN(n1101) );
NAND2_X1 U1010 ( .A1(G210), .A2(n1328), .ZN(n1204) );
NAND2_X1 U1011 ( .A1(n1330), .A2(n1331), .ZN(n1328) );
INV_X1 U1012 ( .A(G237), .ZN(n1330) );
NAND2_X1 U1013 ( .A1(n1332), .A2(n1333), .ZN(n1329) );
XOR2_X1 U1014 ( .A(n1334), .B(n1335), .Z(n1333) );
XNOR2_X1 U1015 ( .A(n1254), .B(n1201), .ZN(n1335) );
NOR2_X1 U1016 ( .A1(n1150), .A2(G953), .ZN(n1201) );
INV_X1 U1017 ( .A(G224), .ZN(n1150) );
XOR2_X1 U1018 ( .A(n1336), .B(n1200), .Z(n1334) );
XNOR2_X1 U1019 ( .A(n1337), .B(n1338), .ZN(n1200) );
XNOR2_X1 U1020 ( .A(KEYINPUT26), .B(n1339), .ZN(n1338) );
INV_X1 U1021 ( .A(n1155), .ZN(n1339) );
XOR2_X1 U1022 ( .A(G110), .B(G122), .Z(n1155) );
XOR2_X1 U1023 ( .A(n1158), .B(n1159), .Z(n1337) );
XNOR2_X1 U1024 ( .A(n1340), .B(n1341), .ZN(n1159) );
NOR2_X1 U1025 ( .A1(KEYINPUT13), .A2(n1062), .ZN(n1341) );
XNOR2_X1 U1026 ( .A(G101), .B(G104), .ZN(n1340) );
XNOR2_X1 U1027 ( .A(n1342), .B(n1343), .ZN(n1158) );
NAND2_X1 U1028 ( .A1(KEYINPUT7), .A2(n1344), .ZN(n1336) );
INV_X1 U1029 ( .A(n1256), .ZN(n1344) );
XNOR2_X1 U1030 ( .A(n1345), .B(G128), .ZN(n1256) );
XNOR2_X1 U1031 ( .A(G902), .B(KEYINPUT50), .ZN(n1332) );
INV_X1 U1032 ( .A(n1227), .ZN(n1295) );
NAND2_X1 U1033 ( .A1(n1102), .A2(n1346), .ZN(n1227) );
NAND4_X1 U1034 ( .A1(G953), .A2(G902), .A3(n1284), .A4(n1151), .ZN(n1346) );
INV_X1 U1035 ( .A(G898), .ZN(n1151) );
NAND3_X1 U1036 ( .A1(n1284), .A2(n1070), .A3(G952), .ZN(n1102) );
NAND2_X1 U1037 ( .A1(G237), .A2(G234), .ZN(n1284) );
XOR2_X1 U1038 ( .A(n1093), .B(KEYINPUT18), .Z(n1270) );
NOR2_X1 U1039 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
AND2_X1 U1040 ( .A1(G221), .A2(n1347), .ZN(n1095) );
XOR2_X1 U1041 ( .A(n1348), .B(G469), .Z(n1094) );
NAND2_X1 U1042 ( .A1(n1349), .A2(n1331), .ZN(n1348) );
XOR2_X1 U1043 ( .A(n1350), .B(n1187), .Z(n1349) );
XOR2_X1 U1044 ( .A(n1351), .B(n1352), .Z(n1187) );
XOR2_X1 U1045 ( .A(n1353), .B(n1354), .Z(n1352) );
XNOR2_X1 U1046 ( .A(G101), .B(KEYINPUT8), .ZN(n1354) );
NAND2_X1 U1047 ( .A1(n1355), .A2(n1356), .ZN(n1353) );
NAND2_X1 U1048 ( .A1(G104), .A2(n1062), .ZN(n1356) );
XOR2_X1 U1049 ( .A(KEYINPUT32), .B(n1357), .Z(n1355) );
NOR2_X1 U1050 ( .A1(G104), .A2(n1062), .ZN(n1357) );
INV_X1 U1051 ( .A(G107), .ZN(n1062) );
XOR2_X1 U1052 ( .A(n1358), .B(n1143), .Z(n1351) );
XOR2_X1 U1053 ( .A(G143), .B(n1359), .Z(n1143) );
NOR2_X1 U1054 ( .A1(KEYINPUT39), .A2(n1360), .ZN(n1359) );
XNOR2_X1 U1055 ( .A(G146), .B(KEYINPUT10), .ZN(n1360) );
NAND2_X1 U1056 ( .A1(n1194), .A2(n1195), .ZN(n1350) );
NAND3_X1 U1057 ( .A1(n1361), .A2(n1070), .A3(G227), .ZN(n1195) );
XNOR2_X1 U1058 ( .A(n1297), .B(n1309), .ZN(n1361) );
NAND2_X1 U1059 ( .A1(n1362), .A2(n1363), .ZN(n1194) );
NAND2_X1 U1060 ( .A1(G227), .A2(n1070), .ZN(n1363) );
XNOR2_X1 U1061 ( .A(G110), .B(n1309), .ZN(n1362) );
NOR2_X1 U1062 ( .A1(n1117), .A2(n1289), .ZN(n1088) );
NOR2_X1 U1063 ( .A1(n1106), .A2(n1364), .ZN(n1289) );
AND2_X1 U1064 ( .A1(n1116), .A2(n1115), .ZN(n1364) );
NOR2_X1 U1065 ( .A1(n1115), .A2(n1116), .ZN(n1106) );
INV_X1 U1066 ( .A(n1164), .ZN(n1116) );
NAND2_X1 U1067 ( .A1(G217), .A2(n1347), .ZN(n1164) );
NAND2_X1 U1068 ( .A1(G234), .A2(n1331), .ZN(n1347) );
NAND2_X1 U1069 ( .A1(n1162), .A2(n1331), .ZN(n1115) );
XNOR2_X1 U1070 ( .A(n1365), .B(n1366), .ZN(n1162) );
XNOR2_X1 U1071 ( .A(n1367), .B(n1368), .ZN(n1366) );
XOR2_X1 U1072 ( .A(n1369), .B(n1370), .Z(n1368) );
AND3_X1 U1073 ( .A1(G221), .A2(n1070), .A3(G234), .ZN(n1370) );
INV_X1 U1074 ( .A(G953), .ZN(n1070) );
NOR2_X1 U1075 ( .A1(G137), .A2(KEYINPUT11), .ZN(n1369) );
XOR2_X1 U1076 ( .A(n1371), .B(n1372), .Z(n1365) );
XOR2_X1 U1077 ( .A(KEYINPUT0), .B(G128), .Z(n1372) );
XNOR2_X1 U1078 ( .A(n1373), .B(n1297), .ZN(n1371) );
NAND2_X1 U1079 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
NAND2_X1 U1080 ( .A1(n1376), .A2(n1304), .ZN(n1375) );
XOR2_X1 U1081 ( .A(n1377), .B(KEYINPUT38), .Z(n1374) );
OR2_X1 U1082 ( .A1(n1376), .A2(n1304), .ZN(n1377) );
XOR2_X1 U1083 ( .A(n1378), .B(n1254), .Z(n1376) );
INV_X1 U1084 ( .A(G125), .ZN(n1254) );
NAND2_X1 U1085 ( .A1(KEYINPUT9), .A2(n1309), .ZN(n1378) );
XOR2_X1 U1086 ( .A(G140), .B(KEYINPUT20), .Z(n1309) );
XNOR2_X1 U1087 ( .A(n1379), .B(n1380), .ZN(n1117) );
XNOR2_X1 U1088 ( .A(KEYINPUT29), .B(n1183), .ZN(n1380) );
INV_X1 U1089 ( .A(G472), .ZN(n1183) );
NAND2_X1 U1090 ( .A1(n1381), .A2(n1331), .ZN(n1379) );
INV_X1 U1091 ( .A(G902), .ZN(n1331) );
XOR2_X1 U1092 ( .A(n1382), .B(n1181), .Z(n1381) );
XOR2_X1 U1093 ( .A(n1383), .B(G101), .Z(n1181) );
NAND2_X1 U1094 ( .A1(n1308), .A2(G210), .ZN(n1383) );
NOR2_X1 U1095 ( .A1(G953), .A2(G237), .ZN(n1308) );
NAND2_X1 U1096 ( .A1(n1384), .A2(n1385), .ZN(n1382) );
NAND2_X1 U1097 ( .A1(n1180), .A2(n1179), .ZN(n1385) );
XOR2_X1 U1098 ( .A(KEYINPUT52), .B(n1386), .Z(n1384) );
NOR2_X1 U1099 ( .A1(n1180), .A2(n1179), .ZN(n1386) );
XNOR2_X1 U1100 ( .A(n1387), .B(n1388), .ZN(n1179) );
INV_X1 U1101 ( .A(n1342), .ZN(n1388) );
XOR2_X1 U1102 ( .A(G113), .B(n1389), .Z(n1342) );
XNOR2_X1 U1103 ( .A(KEYINPUT22), .B(n1291), .ZN(n1389) );
INV_X1 U1104 ( .A(G116), .ZN(n1291) );
NAND2_X1 U1105 ( .A1(KEYINPUT17), .A2(n1367), .ZN(n1387) );
INV_X1 U1106 ( .A(n1343), .ZN(n1367) );
XOR2_X1 U1107 ( .A(G119), .B(KEYINPUT58), .Z(n1343) );
XNOR2_X1 U1108 ( .A(n1358), .B(n1345), .ZN(n1180) );
NAND3_X1 U1109 ( .A1(n1390), .A2(n1391), .A3(n1392), .ZN(n1345) );
NAND2_X1 U1110 ( .A1(KEYINPUT25), .A2(G143), .ZN(n1392) );
NAND3_X1 U1111 ( .A1(n1393), .A2(n1394), .A3(n1304), .ZN(n1391) );
INV_X1 U1112 ( .A(KEYINPUT25), .ZN(n1394) );
OR2_X1 U1113 ( .A1(n1304), .A2(n1393), .ZN(n1390) );
NOR2_X1 U1114 ( .A1(G143), .A2(KEYINPUT15), .ZN(n1393) );
INV_X1 U1115 ( .A(G146), .ZN(n1304) );
XOR2_X1 U1116 ( .A(n1395), .B(n1135), .Z(n1358) );
XOR2_X1 U1117 ( .A(G131), .B(KEYINPUT42), .Z(n1135) );
XNOR2_X1 U1118 ( .A(G137), .B(n1326), .ZN(n1395) );
XNOR2_X1 U1119 ( .A(n1266), .B(G128), .ZN(n1326) );
INV_X1 U1120 ( .A(G134), .ZN(n1266) );
INV_X1 U1121 ( .A(G110), .ZN(n1297) );
endmodule


