//Key = 0011001111111111001100111011000100001010011101111001001111010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331;

XOR2_X1 U737 ( .A(n1009), .B(n1010), .Z(G9) );
XNOR2_X1 U738 ( .A(G107), .B(KEYINPUT17), .ZN(n1010) );
NOR2_X1 U739 ( .A1(n1011), .A2(n1012), .ZN(G75) );
NOR3_X1 U740 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NOR2_X1 U741 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NAND3_X1 U742 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1013) );
NAND2_X1 U743 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U744 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND4_X1 U745 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
NOR2_X1 U746 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND2_X1 U747 ( .A1(n1031), .A2(n1032), .ZN(n1027) );
NAND3_X1 U748 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1026) );
OR2_X1 U749 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U750 ( .A1(n1038), .A2(n1039), .ZN(n1033) );
NAND4_X1 U751 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NAND2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1025) );
INV_X1 U753 ( .A(n1046), .ZN(n1045) );
NAND2_X1 U754 ( .A1(n1038), .A2(n1047), .ZN(n1044) );
NAND2_X1 U755 ( .A1(n1041), .A2(n1043), .ZN(n1047) );
NAND2_X1 U756 ( .A1(n1048), .A2(n1049), .ZN(n1023) );
XOR2_X1 U757 ( .A(n1017), .B(KEYINPUT57), .Z(n1048) );
OR3_X1 U758 ( .A1(n1030), .A2(n1032), .A3(n1031), .ZN(n1017) );
NAND2_X1 U759 ( .A1(n1046), .A2(n1038), .ZN(n1031) );
NOR3_X1 U760 ( .A1(n1050), .A2(G953), .A3(G952), .ZN(n1011) );
INV_X1 U761 ( .A(n1018), .ZN(n1050) );
NAND4_X1 U762 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1018) );
NOR4_X1 U763 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1049), .ZN(n1054) );
INV_X1 U764 ( .A(n1058), .ZN(n1057) );
NOR2_X1 U765 ( .A1(n1059), .A2(n1060), .ZN(n1056) );
NAND3_X1 U766 ( .A1(n1061), .A2(n1036), .A3(n1062), .ZN(n1055) );
NOR3_X1 U767 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1053) );
XOR2_X1 U768 ( .A(n1066), .B(KEYINPUT59), .Z(n1065) );
NOR2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1064) );
XNOR2_X1 U770 ( .A(n1069), .B(n1070), .ZN(n1051) );
NAND2_X1 U771 ( .A1(KEYINPUT31), .A2(n1071), .ZN(n1069) );
XOR2_X1 U772 ( .A(n1072), .B(n1073), .Z(G72) );
XOR2_X1 U773 ( .A(n1074), .B(n1075), .Z(n1073) );
NAND2_X1 U774 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U775 ( .A1(G953), .A2(n1078), .ZN(n1077) );
XOR2_X1 U776 ( .A(n1079), .B(n1080), .Z(n1076) );
XOR2_X1 U777 ( .A(n1081), .B(n1082), .Z(n1080) );
XOR2_X1 U778 ( .A(n1083), .B(n1084), .Z(n1079) );
XNOR2_X1 U779 ( .A(G134), .B(n1085), .ZN(n1084) );
NAND2_X1 U780 ( .A1(KEYINPUT12), .A2(n1086), .ZN(n1083) );
NAND3_X1 U781 ( .A1(KEYINPUT38), .A2(n1087), .A3(n1088), .ZN(n1074) );
XNOR2_X1 U782 ( .A(G953), .B(KEYINPUT21), .ZN(n1088) );
NAND2_X1 U783 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR2_X1 U784 ( .A1(n1091), .A2(n1019), .ZN(n1072) );
NOR2_X1 U785 ( .A1(n1092), .A2(n1078), .ZN(n1091) );
NAND2_X1 U786 ( .A1(n1093), .A2(n1094), .ZN(G69) );
NAND2_X1 U787 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U788 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
NAND2_X1 U789 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U790 ( .A(n1101), .B(KEYINPUT4), .Z(n1093) );
NAND2_X1 U791 ( .A1(n1102), .A2(n1097), .ZN(n1101) );
OR2_X1 U792 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NAND2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(n1099) );
NAND2_X1 U794 ( .A1(G953), .A2(n1105), .ZN(n1104) );
XOR2_X1 U795 ( .A(n1106), .B(n1107), .Z(n1103) );
NOR2_X1 U796 ( .A1(KEYINPUT39), .A2(n1108), .ZN(n1107) );
NAND2_X1 U797 ( .A1(n1109), .A2(n1110), .ZN(n1106) );
NAND2_X1 U798 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U799 ( .A(KEYINPUT27), .B(n1113), .Z(n1109) );
NOR2_X1 U800 ( .A1(n1111), .A2(n1112), .ZN(n1113) );
XNOR2_X1 U801 ( .A(KEYINPUT24), .B(n1114), .ZN(n1112) );
XOR2_X1 U802 ( .A(n1096), .B(KEYINPUT46), .Z(n1102) );
NAND2_X1 U803 ( .A1(G953), .A2(n1115), .ZN(n1096) );
NAND2_X1 U804 ( .A1(G898), .A2(G224), .ZN(n1115) );
NOR2_X1 U805 ( .A1(n1116), .A2(n1117), .ZN(G66) );
XOR2_X1 U806 ( .A(n1118), .B(KEYINPUT54), .Z(n1117) );
NAND2_X1 U807 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U808 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
INV_X1 U809 ( .A(n1123), .ZN(n1122) );
XOR2_X1 U810 ( .A(n1124), .B(KEYINPUT63), .Z(n1119) );
NAND2_X1 U811 ( .A1(n1123), .A2(n1125), .ZN(n1124) );
XOR2_X1 U812 ( .A(KEYINPUT13), .B(n1121), .Z(n1125) );
NOR2_X1 U813 ( .A1(n1126), .A2(n1127), .ZN(n1123) );
NOR2_X1 U814 ( .A1(n1116), .A2(n1128), .ZN(G63) );
XOR2_X1 U815 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U816 ( .A1(n1131), .A2(n1126), .ZN(n1130) );
NOR2_X1 U817 ( .A1(n1116), .A2(n1132), .ZN(G60) );
XOR2_X1 U818 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U819 ( .A1(n1135), .A2(n1126), .ZN(n1133) );
XOR2_X1 U820 ( .A(n1136), .B(G104), .Z(G6) );
NAND2_X1 U821 ( .A1(KEYINPUT19), .A2(n1137), .ZN(n1136) );
NOR2_X1 U822 ( .A1(n1116), .A2(n1138), .ZN(G57) );
XOR2_X1 U823 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U824 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U825 ( .A1(n1143), .A2(n1126), .ZN(n1141) );
XOR2_X1 U826 ( .A(n1144), .B(n1145), .Z(n1139) );
NOR2_X1 U827 ( .A1(KEYINPUT60), .A2(n1146), .ZN(n1145) );
NOR2_X1 U828 ( .A1(KEYINPUT37), .A2(n1147), .ZN(n1144) );
XOR2_X1 U829 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U830 ( .A1(KEYINPUT15), .A2(n1150), .ZN(n1148) );
NOR2_X1 U831 ( .A1(n1116), .A2(n1151), .ZN(G54) );
XOR2_X1 U832 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U833 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND2_X1 U834 ( .A1(n1156), .A2(n1157), .ZN(n1154) );
NAND3_X1 U835 ( .A1(n1158), .A2(n1086), .A3(KEYINPUT7), .ZN(n1157) );
XOR2_X1 U836 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U837 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U838 ( .A1(n1163), .A2(n1164), .ZN(n1156) );
NAND2_X1 U839 ( .A1(KEYINPUT7), .A2(n1086), .ZN(n1164) );
XOR2_X1 U840 ( .A(n1159), .B(n1165), .Z(n1163) );
NOR2_X1 U841 ( .A1(G110), .A2(n1162), .ZN(n1165) );
INV_X1 U842 ( .A(KEYINPUT10), .ZN(n1162) );
XOR2_X1 U843 ( .A(n1166), .B(n1167), .Z(n1152) );
NOR2_X1 U844 ( .A1(n1070), .A2(n1126), .ZN(n1167) );
NAND2_X1 U845 ( .A1(n1168), .A2(KEYINPUT47), .ZN(n1166) );
XNOR2_X1 U846 ( .A(n1169), .B(n1170), .ZN(n1168) );
NOR2_X1 U847 ( .A1(KEYINPUT49), .A2(n1081), .ZN(n1170) );
XOR2_X1 U848 ( .A(n1171), .B(n1172), .Z(n1081) );
NOR2_X1 U849 ( .A1(n1116), .A2(n1173), .ZN(G51) );
XOR2_X1 U850 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR3_X1 U851 ( .A1(n1176), .A2(n1177), .A3(n1126), .ZN(n1175) );
NAND2_X1 U852 ( .A1(G902), .A2(n1015), .ZN(n1126) );
NAND3_X1 U853 ( .A1(n1178), .A2(n1179), .A3(n1089), .ZN(n1015) );
AND4_X1 U854 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1089) );
AND4_X1 U855 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1183) );
XNOR2_X1 U856 ( .A(KEYINPUT43), .B(n1090), .ZN(n1179) );
INV_X1 U857 ( .A(n1100), .ZN(n1178) );
NAND4_X1 U858 ( .A1(n1137), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1100) );
AND4_X1 U859 ( .A1(n1009), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1190) );
NAND3_X1 U860 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1009) );
NAND2_X1 U861 ( .A1(n1197), .A2(n1198), .ZN(n1189) );
NAND2_X1 U862 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND3_X1 U863 ( .A1(n1201), .A2(n1202), .A3(n1195), .ZN(n1200) );
NAND2_X1 U864 ( .A1(n1203), .A2(n1194), .ZN(n1199) );
NAND3_X1 U865 ( .A1(n1196), .A2(n1195), .A3(n1204), .ZN(n1137) );
XOR2_X1 U866 ( .A(KEYINPUT32), .B(n1205), .Z(n1176) );
NAND2_X1 U867 ( .A1(KEYINPUT26), .A2(n1206), .ZN(n1174) );
XOR2_X1 U868 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR2_X1 U869 ( .A1(KEYINPUT16), .A2(n1209), .ZN(n1207) );
NOR2_X1 U870 ( .A1(n1019), .A2(G952), .ZN(n1116) );
XNOR2_X1 U871 ( .A(n1210), .B(n1211), .ZN(G48) );
NAND2_X1 U872 ( .A1(n1212), .A2(n1213), .ZN(n1210) );
NAND3_X1 U873 ( .A1(n1214), .A2(n1041), .A3(n1215), .ZN(n1213) );
OR2_X1 U874 ( .A1(n1090), .A2(n1215), .ZN(n1212) );
INV_X1 U875 ( .A(KEYINPUT11), .ZN(n1215) );
NAND2_X1 U876 ( .A1(n1214), .A2(n1204), .ZN(n1090) );
XNOR2_X1 U877 ( .A(G143), .B(n1182), .ZN(G45) );
NAND4_X1 U878 ( .A1(n1201), .A2(n1202), .A3(n1216), .A4(n1217), .ZN(n1182) );
NOR2_X1 U879 ( .A1(n1218), .A2(n1040), .ZN(n1217) );
XNOR2_X1 U880 ( .A(G140), .B(n1180), .ZN(G42) );
NAND3_X1 U881 ( .A1(n1219), .A2(n1204), .A3(n1220), .ZN(n1180) );
XNOR2_X1 U882 ( .A(G137), .B(n1181), .ZN(G39) );
NAND2_X1 U883 ( .A1(n1221), .A2(n1220), .ZN(n1181) );
XOR2_X1 U884 ( .A(G134), .B(n1222), .Z(G36) );
NOR2_X1 U885 ( .A1(KEYINPUT29), .A2(n1187), .ZN(n1222) );
NAND3_X1 U886 ( .A1(n1203), .A2(n1194), .A3(n1220), .ZN(n1187) );
XOR2_X1 U887 ( .A(n1223), .B(n1224), .Z(G33) );
NOR2_X1 U888 ( .A1(KEYINPUT40), .A2(n1186), .ZN(n1224) );
NAND3_X1 U889 ( .A1(n1203), .A2(n1204), .A3(n1220), .ZN(n1186) );
AND4_X1 U890 ( .A1(n1021), .A2(n1216), .A3(n1225), .A4(n1226), .ZN(n1220) );
XNOR2_X1 U891 ( .A(G131), .B(KEYINPUT3), .ZN(n1223) );
XNOR2_X1 U892 ( .A(G128), .B(n1185), .ZN(G30) );
NAND2_X1 U893 ( .A1(n1214), .A2(n1194), .ZN(n1185) );
AND4_X1 U894 ( .A1(n1227), .A2(n1216), .A3(n1228), .A4(n1229), .ZN(n1214) );
NAND3_X1 U895 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(G3) );
NAND2_X1 U896 ( .A1(G101), .A2(n1188), .ZN(n1232) );
NAND2_X1 U897 ( .A1(n1233), .A2(n1234), .ZN(n1231) );
INV_X1 U898 ( .A(KEYINPUT51), .ZN(n1234) );
NAND2_X1 U899 ( .A1(n1235), .A2(n1236), .ZN(n1233) );
XNOR2_X1 U900 ( .A(KEYINPUT56), .B(n1150), .ZN(n1236) );
NAND2_X1 U901 ( .A1(KEYINPUT51), .A2(n1237), .ZN(n1230) );
NAND2_X1 U902 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND3_X1 U903 ( .A1(KEYINPUT56), .A2(n1235), .A3(n1150), .ZN(n1239) );
INV_X1 U904 ( .A(n1188), .ZN(n1235) );
NAND3_X1 U905 ( .A1(n1203), .A2(n1196), .A3(n1046), .ZN(n1188) );
OR2_X1 U906 ( .A1(n1150), .A2(KEYINPUT56), .ZN(n1238) );
INV_X1 U907 ( .A(G101), .ZN(n1150) );
XOR2_X1 U908 ( .A(n1240), .B(n1241), .Z(G27) );
NOR2_X1 U909 ( .A1(KEYINPUT25), .A2(n1085), .ZN(n1241) );
INV_X1 U910 ( .A(G125), .ZN(n1085) );
NAND2_X1 U911 ( .A1(n1242), .A2(n1243), .ZN(n1240) );
NAND4_X1 U912 ( .A1(n1038), .A2(n1227), .A3(n1244), .A4(n1245), .ZN(n1243) );
NOR2_X1 U913 ( .A1(n1219), .A2(n1041), .ZN(n1244) );
INV_X1 U914 ( .A(n1204), .ZN(n1041) );
OR2_X1 U915 ( .A1(n1184), .A2(n1245), .ZN(n1242) );
INV_X1 U916 ( .A(KEYINPUT6), .ZN(n1245) );
NAND4_X1 U917 ( .A1(n1038), .A2(n1227), .A3(n1219), .A4(n1204), .ZN(n1184) );
INV_X1 U918 ( .A(n1218), .ZN(n1227) );
NAND2_X1 U919 ( .A1(n1246), .A2(n1226), .ZN(n1218) );
NAND2_X1 U920 ( .A1(n1030), .A2(n1247), .ZN(n1226) );
NAND4_X1 U921 ( .A1(G953), .A2(G902), .A3(n1248), .A4(n1078), .ZN(n1247) );
INV_X1 U922 ( .A(G900), .ZN(n1078) );
XNOR2_X1 U923 ( .A(G122), .B(n1249), .ZN(G24) );
NAND4_X1 U924 ( .A1(n1250), .A2(n1251), .A3(n1195), .A4(n1252), .ZN(n1249) );
AND2_X1 U925 ( .A1(n1202), .A2(n1201), .ZN(n1252) );
XOR2_X1 U926 ( .A(n1063), .B(KEYINPUT1), .Z(n1201) );
INV_X1 U927 ( .A(n1032), .ZN(n1195) );
NAND2_X1 U928 ( .A1(n1052), .A2(n1253), .ZN(n1032) );
OR2_X1 U929 ( .A1(n1197), .A2(KEYINPUT53), .ZN(n1251) );
NAND2_X1 U930 ( .A1(KEYINPUT53), .A2(n1254), .ZN(n1250) );
NAND2_X1 U931 ( .A1(n1255), .A2(n1016), .ZN(n1254) );
XNOR2_X1 U932 ( .A(G119), .B(n1193), .ZN(G21) );
NAND2_X1 U933 ( .A1(n1197), .A2(n1221), .ZN(n1193) );
AND3_X1 U934 ( .A1(n1228), .A2(n1229), .A3(n1046), .ZN(n1221) );
XNOR2_X1 U935 ( .A(G116), .B(n1256), .ZN(G18) );
NAND3_X1 U936 ( .A1(n1197), .A2(n1203), .A3(n1257), .ZN(n1256) );
XNOR2_X1 U937 ( .A(n1194), .B(KEYINPUT9), .ZN(n1257) );
INV_X1 U938 ( .A(n1043), .ZN(n1194) );
NAND2_X1 U939 ( .A1(n1258), .A2(n1202), .ZN(n1043) );
AND2_X1 U940 ( .A1(n1255), .A2(n1246), .ZN(n1197) );
INV_X1 U941 ( .A(n1016), .ZN(n1246) );
XOR2_X1 U942 ( .A(n1259), .B(KEYINPUT14), .Z(n1016) );
XNOR2_X1 U943 ( .A(G113), .B(n1192), .ZN(G15) );
NAND4_X1 U944 ( .A1(n1255), .A2(n1203), .A3(n1204), .A4(n1259), .ZN(n1192) );
NOR2_X1 U945 ( .A1(n1202), .A2(n1258), .ZN(n1204) );
INV_X1 U946 ( .A(n1063), .ZN(n1258) );
INV_X1 U947 ( .A(n1040), .ZN(n1203) );
NAND2_X1 U948 ( .A1(n1052), .A2(n1229), .ZN(n1040) );
AND2_X1 U949 ( .A1(n1038), .A2(n1260), .ZN(n1255) );
NOR2_X1 U950 ( .A1(n1037), .A2(n1261), .ZN(n1038) );
INV_X1 U951 ( .A(n1036), .ZN(n1261) );
XNOR2_X1 U952 ( .A(G110), .B(n1191), .ZN(G12) );
NAND3_X1 U953 ( .A1(n1219), .A2(n1196), .A3(n1046), .ZN(n1191) );
NOR2_X1 U954 ( .A1(n1202), .A2(n1063), .ZN(n1046) );
XOR2_X1 U955 ( .A(n1262), .B(n1135), .Z(n1063) );
INV_X1 U956 ( .A(G475), .ZN(n1135) );
OR2_X1 U957 ( .A1(n1134), .A2(G902), .ZN(n1262) );
XNOR2_X1 U958 ( .A(n1263), .B(n1264), .ZN(n1134) );
XOR2_X1 U959 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U960 ( .A(n1267), .B(n1268), .Z(n1263) );
XNOR2_X1 U961 ( .A(G131), .B(n1269), .ZN(n1268) );
NAND3_X1 U962 ( .A1(G214), .A2(n1019), .A3(n1270), .ZN(n1269) );
NAND2_X1 U963 ( .A1(n1271), .A2(KEYINPUT48), .ZN(n1267) );
XNOR2_X1 U964 ( .A(G104), .B(n1272), .ZN(n1271) );
XOR2_X1 U965 ( .A(G122), .B(G113), .Z(n1272) );
NAND3_X1 U966 ( .A1(n1273), .A2(n1274), .A3(n1061), .ZN(n1202) );
NAND2_X1 U967 ( .A1(n1067), .A2(n1068), .ZN(n1061) );
OR3_X1 U968 ( .A1(n1068), .A2(n1067), .A3(KEYINPUT58), .ZN(n1274) );
XOR2_X1 U969 ( .A(n1131), .B(KEYINPUT33), .Z(n1068) );
INV_X1 U970 ( .A(G478), .ZN(n1131) );
NAND2_X1 U971 ( .A1(KEYINPUT58), .A2(n1067), .ZN(n1273) );
NOR2_X1 U972 ( .A1(n1129), .A2(G902), .ZN(n1067) );
XOR2_X1 U973 ( .A(n1275), .B(n1276), .Z(n1129) );
XNOR2_X1 U974 ( .A(n1277), .B(n1278), .ZN(n1276) );
XOR2_X1 U975 ( .A(n1279), .B(n1280), .Z(n1278) );
NOR2_X1 U976 ( .A1(KEYINPUT30), .A2(n1281), .ZN(n1280) );
XNOR2_X1 U977 ( .A(n1282), .B(n1283), .ZN(n1281) );
NAND2_X1 U978 ( .A1(KEYINPUT23), .A2(n1265), .ZN(n1282) );
NAND2_X1 U979 ( .A1(G217), .A2(n1284), .ZN(n1279) );
XNOR2_X1 U980 ( .A(G107), .B(n1285), .ZN(n1275) );
XOR2_X1 U981 ( .A(G134), .B(G122), .Z(n1285) );
AND3_X1 U982 ( .A1(n1259), .A2(n1260), .A3(n1216), .ZN(n1196) );
INV_X1 U983 ( .A(n1034), .ZN(n1216) );
NAND2_X1 U984 ( .A1(n1037), .A2(n1036), .ZN(n1034) );
NAND2_X1 U985 ( .A1(G221), .A2(n1286), .ZN(n1036) );
NAND3_X1 U986 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n1037) );
NAND2_X1 U987 ( .A1(n1290), .A2(n1070), .ZN(n1289) );
INV_X1 U988 ( .A(G469), .ZN(n1070) );
NAND2_X1 U989 ( .A1(n1291), .A2(KEYINPUT42), .ZN(n1290) );
XNOR2_X1 U990 ( .A(n1071), .B(KEYINPUT52), .ZN(n1291) );
INV_X1 U991 ( .A(n1292), .ZN(n1071) );
NAND3_X1 U992 ( .A1(KEYINPUT42), .A2(G469), .A3(n1292), .ZN(n1288) );
OR2_X1 U993 ( .A1(n1292), .A2(KEYINPUT42), .ZN(n1287) );
NAND2_X1 U994 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U995 ( .A(n1295), .B(n1296), .Z(n1293) );
XNOR2_X1 U996 ( .A(n1297), .B(n1114), .ZN(n1296) );
XNOR2_X1 U997 ( .A(n1298), .B(n1171), .ZN(n1295) );
NAND2_X1 U998 ( .A1(KEYINPUT22), .A2(n1299), .ZN(n1171) );
XNOR2_X1 U999 ( .A(KEYINPUT18), .B(n1211), .ZN(n1299) );
NOR2_X1 U1000 ( .A1(KEYINPUT44), .A2(n1300), .ZN(n1298) );
XOR2_X1 U1001 ( .A(n1301), .B(n1302), .Z(n1300) );
XNOR2_X1 U1002 ( .A(G110), .B(n1159), .ZN(n1302) );
NOR2_X1 U1003 ( .A1(n1092), .A2(G953), .ZN(n1159) );
INV_X1 U1004 ( .A(G227), .ZN(n1092) );
NAND2_X1 U1005 ( .A1(KEYINPUT55), .A2(n1303), .ZN(n1301) );
INV_X1 U1006 ( .A(n1086), .ZN(n1303) );
NAND2_X1 U1007 ( .A1(n1030), .A2(n1304), .ZN(n1260) );
NAND4_X1 U1008 ( .A1(G953), .A2(G902), .A3(n1248), .A4(n1105), .ZN(n1304) );
INV_X1 U1009 ( .A(G898), .ZN(n1105) );
NAND3_X1 U1010 ( .A1(n1248), .A2(n1019), .A3(G952), .ZN(n1030) );
NAND2_X1 U1011 ( .A1(G237), .A2(G234), .ZN(n1248) );
NOR2_X1 U1012 ( .A1(n1029), .A2(n1021), .ZN(n1259) );
AND3_X1 U1013 ( .A1(n1305), .A2(n1306), .A3(n1062), .ZN(n1021) );
NAND2_X1 U1014 ( .A1(n1059), .A2(n1060), .ZN(n1062) );
NAND2_X1 U1015 ( .A1(n1060), .A2(n1307), .ZN(n1306) );
OR3_X1 U1016 ( .A1(n1060), .A2(n1059), .A3(n1307), .ZN(n1305) );
INV_X1 U1017 ( .A(KEYINPUT8), .ZN(n1307) );
NOR2_X1 U1018 ( .A1(n1177), .A2(n1205), .ZN(n1059) );
INV_X1 U1019 ( .A(G210), .ZN(n1177) );
NAND2_X1 U1020 ( .A1(n1308), .A2(n1294), .ZN(n1060) );
XNOR2_X1 U1021 ( .A(n1208), .B(n1209), .ZN(n1308) );
XNOR2_X1 U1022 ( .A(n1114), .B(n1309), .ZN(n1209) );
XOR2_X1 U1023 ( .A(n1111), .B(n1108), .Z(n1309) );
XNOR2_X1 U1024 ( .A(G122), .B(G110), .ZN(n1108) );
INV_X1 U1025 ( .A(n1169), .ZN(n1114) );
XOR2_X1 U1026 ( .A(G101), .B(n1310), .Z(n1169) );
XNOR2_X1 U1027 ( .A(n1311), .B(G104), .ZN(n1310) );
INV_X1 U1028 ( .A(G107), .ZN(n1311) );
XNOR2_X1 U1029 ( .A(n1312), .B(n1313), .ZN(n1208) );
XOR2_X1 U1030 ( .A(n1314), .B(n1172), .Z(n1312) );
NAND2_X1 U1031 ( .A1(G224), .A2(n1019), .ZN(n1314) );
INV_X1 U1032 ( .A(n1225), .ZN(n1029) );
XOR2_X1 U1033 ( .A(n1049), .B(KEYINPUT2), .Z(n1225) );
NOR2_X1 U1034 ( .A1(n1315), .A2(n1205), .ZN(n1049) );
NOR2_X1 U1035 ( .A1(n1316), .A2(G237), .ZN(n1205) );
XNOR2_X1 U1036 ( .A(KEYINPUT36), .B(G902), .ZN(n1316) );
INV_X1 U1037 ( .A(G214), .ZN(n1315) );
INV_X1 U1038 ( .A(n1042), .ZN(n1219) );
NAND2_X1 U1039 ( .A1(n1228), .A2(n1253), .ZN(n1042) );
XNOR2_X1 U1040 ( .A(n1229), .B(KEYINPUT5), .ZN(n1253) );
NAND2_X1 U1041 ( .A1(n1317), .A2(n1058), .ZN(n1229) );
NAND3_X1 U1042 ( .A1(n1143), .A2(n1294), .A3(n1318), .ZN(n1058) );
INV_X1 U1043 ( .A(G472), .ZN(n1143) );
XOR2_X1 U1044 ( .A(n1066), .B(KEYINPUT35), .Z(n1317) );
NAND2_X1 U1045 ( .A1(G472), .A2(n1319), .ZN(n1066) );
NAND2_X1 U1046 ( .A1(n1318), .A2(n1294), .ZN(n1319) );
XOR2_X1 U1047 ( .A(n1320), .B(n1321), .Z(n1318) );
XOR2_X1 U1048 ( .A(n1149), .B(n1322), .Z(n1321) );
NOR2_X1 U1049 ( .A1(G101), .A2(KEYINPUT20), .ZN(n1322) );
AND3_X1 U1050 ( .A1(G210), .A2(n1019), .A3(n1270), .ZN(n1149) );
XNOR2_X1 U1051 ( .A(G237), .B(KEYINPUT28), .ZN(n1270) );
XOR2_X1 U1052 ( .A(n1142), .B(n1146), .Z(n1320) );
XOR2_X1 U1053 ( .A(n1111), .B(KEYINPUT50), .Z(n1146) );
XOR2_X1 U1054 ( .A(n1323), .B(n1277), .Z(n1111) );
XOR2_X1 U1055 ( .A(G116), .B(KEYINPUT62), .Z(n1277) );
XNOR2_X1 U1056 ( .A(G113), .B(G119), .ZN(n1323) );
XOR2_X1 U1057 ( .A(G146), .B(n1297), .Z(n1142) );
XOR2_X1 U1058 ( .A(n1155), .B(n1172), .Z(n1297) );
XOR2_X1 U1059 ( .A(n1265), .B(n1283), .Z(n1172) );
XOR2_X1 U1060 ( .A(G143), .B(KEYINPUT61), .Z(n1265) );
XOR2_X1 U1061 ( .A(n1082), .B(n1324), .Z(n1155) );
NOR2_X1 U1062 ( .A1(G134), .A2(KEYINPUT0), .ZN(n1324) );
XOR2_X1 U1063 ( .A(G131), .B(G137), .Z(n1082) );
INV_X1 U1064 ( .A(n1052), .ZN(n1228) );
XNOR2_X1 U1065 ( .A(n1325), .B(n1127), .ZN(n1052) );
NAND2_X1 U1066 ( .A1(G217), .A2(n1286), .ZN(n1127) );
NAND2_X1 U1067 ( .A1(G234), .A2(n1294), .ZN(n1286) );
NAND2_X1 U1068 ( .A1(n1121), .A2(n1294), .ZN(n1325) );
INV_X1 U1069 ( .A(G902), .ZN(n1294) );
XNOR2_X1 U1070 ( .A(n1326), .B(n1327), .ZN(n1121) );
XOR2_X1 U1071 ( .A(n1328), .B(n1329), .Z(n1327) );
XNOR2_X1 U1072 ( .A(G119), .B(n1161), .ZN(n1329) );
INV_X1 U1073 ( .A(G110), .ZN(n1161) );
XOR2_X1 U1074 ( .A(KEYINPUT45), .B(G137), .Z(n1328) );
XOR2_X1 U1075 ( .A(n1330), .B(n1266), .Z(n1326) );
XOR2_X1 U1076 ( .A(n1313), .B(n1086), .Z(n1266) );
XOR2_X1 U1077 ( .A(G140), .B(KEYINPUT41), .Z(n1086) );
XNOR2_X1 U1078 ( .A(G125), .B(n1211), .ZN(n1313) );
INV_X1 U1079 ( .A(G146), .ZN(n1211) );
XOR2_X1 U1080 ( .A(n1331), .B(n1283), .Z(n1330) );
XOR2_X1 U1081 ( .A(G128), .B(KEYINPUT34), .Z(n1283) );
NAND2_X1 U1082 ( .A1(n1284), .A2(G221), .ZN(n1331) );
AND2_X1 U1083 ( .A1(G234), .A2(n1019), .ZN(n1284) );
INV_X1 U1084 ( .A(G953), .ZN(n1019) );
endmodule


