//Key = 0100001111101010001011111100011001110111010100000000100010101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301;

NAND2_X1 U731 ( .A1(n1001), .A2(n1002), .ZN(G9) );
OR2_X1 U732 ( .A1(n1003), .A2(G107), .ZN(n1002) );
XOR2_X1 U733 ( .A(n1004), .B(KEYINPUT27), .Z(n1001) );
NAND2_X1 U734 ( .A1(G107), .A2(n1003), .ZN(n1004) );
NOR2_X1 U735 ( .A1(n1005), .A2(n1006), .ZN(G75) );
NOR4_X1 U736 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1006) );
NOR3_X1 U737 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1010) );
XNOR2_X1 U738 ( .A(n1014), .B(KEYINPUT12), .ZN(n1013) );
XNOR2_X1 U739 ( .A(n1015), .B(KEYINPUT61), .ZN(n1012) );
NOR4_X1 U740 ( .A1(n1016), .A2(n1017), .A3(n1018), .A4(n1014), .ZN(n1009) );
NOR2_X1 U741 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR2_X1 U742 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR3_X1 U743 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1021) );
NOR2_X1 U744 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
XNOR2_X1 U745 ( .A(n1028), .B(KEYINPUT31), .ZN(n1026) );
NOR2_X1 U746 ( .A1(n1029), .A2(n1030), .ZN(n1024) );
XNOR2_X1 U747 ( .A(n1031), .B(n1032), .ZN(n1029) );
NOR2_X1 U748 ( .A1(n1033), .A2(n1034), .ZN(n1023) );
NOR3_X1 U749 ( .A1(n1034), .A2(n1035), .A3(n1030), .ZN(n1019) );
NOR2_X1 U750 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
INV_X1 U751 ( .A(n1038), .ZN(n1008) );
NAND3_X1 U752 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1007) );
NAND2_X1 U753 ( .A1(n1015), .A2(n1042), .ZN(n1039) );
NOR4_X1 U754 ( .A1(n1017), .A2(n1034), .A3(n1030), .A4(n1022), .ZN(n1015) );
AND3_X1 U755 ( .A1(n1041), .A2(n1043), .A3(n1040), .ZN(n1005) );
NAND4_X1 U756 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1040) );
NOR4_X1 U757 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
XNOR2_X1 U758 ( .A(KEYINPUT51), .B(n1052), .ZN(n1051) );
XOR2_X1 U759 ( .A(KEYINPUT15), .B(n1053), .Z(n1050) );
XNOR2_X1 U760 ( .A(n1054), .B(n1055), .ZN(n1049) );
NOR2_X1 U761 ( .A1(KEYINPUT5), .A2(n1056), .ZN(n1055) );
NOR3_X1 U762 ( .A1(n1016), .A2(n1057), .A3(n1058), .ZN(n1046) );
XNOR2_X1 U763 ( .A(n1059), .B(n1060), .ZN(n1044) );
NOR2_X1 U764 ( .A1(n1061), .A2(KEYINPUT53), .ZN(n1060) );
XOR2_X1 U765 ( .A(n1062), .B(n1063), .Z(G72) );
NOR2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
AND2_X1 U767 ( .A1(G227), .A2(G900), .ZN(n1064) );
NAND2_X1 U768 ( .A1(n1066), .A2(n1067), .ZN(n1062) );
NAND2_X1 U769 ( .A1(n1068), .A2(n1065), .ZN(n1067) );
XNOR2_X1 U770 ( .A(n1069), .B(n1070), .ZN(n1068) );
NOR3_X1 U771 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1069) );
XOR2_X1 U772 ( .A(n1074), .B(KEYINPUT40), .Z(n1073) );
NAND3_X1 U773 ( .A1(n1075), .A2(n1070), .A3(G953), .ZN(n1066) );
NAND3_X1 U774 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1070) );
NAND2_X1 U775 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
INV_X1 U776 ( .A(KEYINPUT35), .ZN(n1080) );
NAND3_X1 U777 ( .A1(KEYINPUT35), .A2(n1081), .A3(n1082), .ZN(n1077) );
OR2_X1 U778 ( .A1(n1082), .A2(n1081), .ZN(n1076) );
NOR2_X1 U779 ( .A1(KEYINPUT59), .A2(n1079), .ZN(n1081) );
XNOR2_X1 U780 ( .A(n1083), .B(n1084), .ZN(n1079) );
XNOR2_X1 U781 ( .A(n1085), .B(n1086), .ZN(n1083) );
NOR2_X1 U782 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U783 ( .A(n1089), .B(KEYINPUT8), .Z(n1088) );
NOR2_X1 U784 ( .A1(G137), .A2(n1090), .ZN(n1087) );
XNOR2_X1 U785 ( .A(KEYINPUT1), .B(n1091), .ZN(n1090) );
XOR2_X1 U786 ( .A(n1092), .B(n1093), .Z(G69) );
XOR2_X1 U787 ( .A(n1094), .B(n1095), .Z(n1093) );
OR2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U789 ( .A1(G953), .A2(n1098), .ZN(n1094) );
NAND2_X1 U790 ( .A1(G898), .A2(G224), .ZN(n1098) );
AND2_X1 U791 ( .A1(n1099), .A2(n1065), .ZN(n1092) );
NOR2_X1 U792 ( .A1(n1100), .A2(n1101), .ZN(G66) );
NOR3_X1 U793 ( .A1(n1061), .A2(n1102), .A3(n1103), .ZN(n1101) );
NOR3_X1 U794 ( .A1(n1104), .A2(n1059), .A3(n1105), .ZN(n1103) );
NOR2_X1 U795 ( .A1(n1106), .A2(n1107), .ZN(n1102) );
NOR2_X1 U796 ( .A1(n1038), .A2(n1059), .ZN(n1106) );
NOR2_X1 U797 ( .A1(n1108), .A2(n1109), .ZN(G63) );
XOR2_X1 U798 ( .A(n1110), .B(n1111), .Z(n1109) );
AND2_X1 U799 ( .A1(G478), .A2(n1112), .ZN(n1111) );
NOR2_X1 U800 ( .A1(G952), .A2(n1113), .ZN(n1108) );
XNOR2_X1 U801 ( .A(KEYINPUT7), .B(n1065), .ZN(n1113) );
NOR2_X1 U802 ( .A1(n1100), .A2(n1114), .ZN(G60) );
XOR2_X1 U803 ( .A(n1115), .B(n1116), .Z(n1114) );
AND2_X1 U804 ( .A1(G475), .A2(n1112), .ZN(n1115) );
XNOR2_X1 U805 ( .A(G104), .B(n1117), .ZN(G6) );
NAND2_X1 U806 ( .A1(KEYINPUT23), .A2(n1118), .ZN(n1117) );
INV_X1 U807 ( .A(n1119), .ZN(n1118) );
NOR2_X1 U808 ( .A1(n1100), .A2(n1120), .ZN(G57) );
XOR2_X1 U809 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U810 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U811 ( .A1(n1056), .A2(n1105), .ZN(n1123) );
INV_X1 U812 ( .A(n1112), .ZN(n1105) );
XOR2_X1 U813 ( .A(n1125), .B(G101), .Z(n1121) );
NOR3_X1 U814 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(G54) );
AND2_X1 U815 ( .A1(KEYINPUT39), .A2(n1100), .ZN(n1128) );
NOR3_X1 U816 ( .A1(KEYINPUT39), .A2(n1065), .A3(n1043), .ZN(n1127) );
INV_X1 U817 ( .A(G952), .ZN(n1043) );
XOR2_X1 U818 ( .A(n1129), .B(n1130), .Z(n1126) );
XOR2_X1 U819 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U820 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U821 ( .A1(G953), .A2(n1135), .ZN(n1133) );
XOR2_X1 U822 ( .A(n1136), .B(n1137), .Z(n1129) );
XNOR2_X1 U823 ( .A(n1138), .B(n1139), .ZN(n1137) );
NAND3_X1 U824 ( .A1(n1112), .A2(G469), .A3(KEYINPUT24), .ZN(n1139) );
NAND2_X1 U825 ( .A1(KEYINPUT34), .A2(n1140), .ZN(n1138) );
XOR2_X1 U826 ( .A(n1141), .B(n1142), .Z(n1136) );
NOR2_X1 U827 ( .A1(KEYINPUT13), .A2(n1143), .ZN(n1142) );
XOR2_X1 U828 ( .A(n1084), .B(n1144), .Z(n1143) );
XNOR2_X1 U829 ( .A(n1145), .B(n1146), .ZN(n1144) );
NOR2_X1 U830 ( .A1(KEYINPUT19), .A2(n1147), .ZN(n1146) );
NOR2_X1 U831 ( .A1(n1100), .A2(n1148), .ZN(G51) );
XOR2_X1 U832 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U833 ( .A(n1151), .B(n1096), .Z(n1150) );
NAND2_X1 U834 ( .A1(KEYINPUT43), .A2(n1152), .ZN(n1151) );
XNOR2_X1 U835 ( .A(n1153), .B(n1154), .ZN(n1152) );
NAND2_X1 U836 ( .A1(KEYINPUT37), .A2(n1155), .ZN(n1153) );
XOR2_X1 U837 ( .A(KEYINPUT18), .B(n1156), .Z(n1155) );
XNOR2_X1 U838 ( .A(n1157), .B(n1158), .ZN(n1149) );
AND2_X1 U839 ( .A1(G210), .A2(n1112), .ZN(n1157) );
NOR2_X1 U840 ( .A1(n1159), .A2(n1038), .ZN(n1112) );
NOR4_X1 U841 ( .A1(n1074), .A2(n1099), .A3(n1071), .A4(n1160), .ZN(n1038) );
XNOR2_X1 U842 ( .A(KEYINPUT41), .B(n1072), .ZN(n1160) );
NAND3_X1 U843 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1071) );
NAND4_X1 U844 ( .A1(n1164), .A2(n1165), .A3(n1036), .A4(n1042), .ZN(n1163) );
NAND4_X1 U845 ( .A1(n1119), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1099) );
AND4_X1 U846 ( .A1(n1003), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1168) );
NAND3_X1 U847 ( .A1(n1172), .A2(n1036), .A3(n1173), .ZN(n1003) );
NAND3_X1 U848 ( .A1(n1174), .A2(n1175), .A3(n1173), .ZN(n1167) );
NAND2_X1 U849 ( .A1(n1033), .A2(n1027), .ZN(n1175) );
INV_X1 U850 ( .A(n1176), .ZN(n1033) );
NAND3_X1 U851 ( .A1(n1173), .A2(n1172), .A3(n1037), .ZN(n1119) );
NAND4_X1 U852 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1074) );
NOR2_X1 U853 ( .A1(n1065), .A2(G952), .ZN(n1100) );
XNOR2_X1 U854 ( .A(G146), .B(n1177), .ZN(G48) );
NAND4_X1 U855 ( .A1(n1037), .A2(n1164), .A3(n1165), .A4(n1042), .ZN(n1177) );
XNOR2_X1 U856 ( .A(G143), .B(n1178), .ZN(G45) );
NAND4_X1 U857 ( .A1(n1165), .A2(n1042), .A3(n1181), .A4(n1176), .ZN(n1178) );
AND2_X1 U858 ( .A1(n1182), .A2(n1048), .ZN(n1181) );
XNOR2_X1 U859 ( .A(G140), .B(n1179), .ZN(G42) );
NAND3_X1 U860 ( .A1(n1037), .A2(n1183), .A3(n1184), .ZN(n1179) );
XNOR2_X1 U861 ( .A(G137), .B(n1180), .ZN(G39) );
NAND3_X1 U862 ( .A1(n1183), .A2(n1174), .A3(n1164), .ZN(n1180) );
XNOR2_X1 U863 ( .A(G134), .B(n1161), .ZN(G36) );
NAND3_X1 U864 ( .A1(n1036), .A2(n1176), .A3(n1183), .ZN(n1161) );
XNOR2_X1 U865 ( .A(G131), .B(n1162), .ZN(G33) );
NAND3_X1 U866 ( .A1(n1183), .A2(n1176), .A3(n1037), .ZN(n1162) );
AND3_X1 U867 ( .A1(n1052), .A2(n1011), .A3(n1165), .ZN(n1183) );
XNOR2_X1 U868 ( .A(G128), .B(n1185), .ZN(G30) );
NAND4_X1 U869 ( .A1(n1186), .A2(n1187), .A3(n1165), .A4(n1036), .ZN(n1185) );
AND3_X1 U870 ( .A1(n1188), .A2(n1045), .A3(n1032), .ZN(n1165) );
XNOR2_X1 U871 ( .A(n1164), .B(KEYINPUT25), .ZN(n1187) );
XNOR2_X1 U872 ( .A(n1042), .B(KEYINPUT58), .ZN(n1186) );
XNOR2_X1 U873 ( .A(G101), .B(n1189), .ZN(G3) );
NAND4_X1 U874 ( .A1(n1174), .A2(n1176), .A3(n1190), .A4(n1191), .ZN(n1189) );
NOR3_X1 U875 ( .A1(n1192), .A2(n1031), .A3(n1193), .ZN(n1191) );
XNOR2_X1 U876 ( .A(KEYINPUT32), .B(n1194), .ZN(n1190) );
XOR2_X1 U877 ( .A(n1195), .B(G125), .Z(G27) );
NAND2_X1 U878 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND2_X1 U879 ( .A1(n1072), .A2(n1198), .ZN(n1197) );
INV_X1 U880 ( .A(KEYINPUT44), .ZN(n1198) );
AND2_X1 U881 ( .A1(n1199), .A2(n1028), .ZN(n1072) );
NAND3_X1 U882 ( .A1(n1199), .A2(n1034), .A3(KEYINPUT44), .ZN(n1196) );
AND4_X1 U883 ( .A1(n1184), .A2(n1037), .A3(n1042), .A4(n1188), .ZN(n1199) );
NAND2_X1 U884 ( .A1(n1017), .A2(n1200), .ZN(n1188) );
NAND4_X1 U885 ( .A1(G902), .A2(G953), .A3(n1201), .A4(n1202), .ZN(n1200) );
INV_X1 U886 ( .A(n1075), .ZN(n1201) );
XNOR2_X1 U887 ( .A(G900), .B(KEYINPUT60), .ZN(n1075) );
XOR2_X1 U888 ( .A(n1166), .B(n1203), .Z(G24) );
NAND2_X1 U889 ( .A1(KEYINPUT9), .A2(G122), .ZN(n1203) );
NAND4_X1 U890 ( .A1(n1204), .A2(n1172), .A3(n1048), .A4(n1182), .ZN(n1166) );
INV_X1 U891 ( .A(n1030), .ZN(n1172) );
XOR2_X1 U892 ( .A(n1171), .B(n1205), .Z(G21) );
NAND2_X1 U893 ( .A1(KEYINPUT22), .A2(G119), .ZN(n1205) );
NAND3_X1 U894 ( .A1(n1164), .A2(n1174), .A3(n1204), .ZN(n1171) );
NOR2_X1 U895 ( .A1(n1206), .A2(n1207), .ZN(n1164) );
XNOR2_X1 U896 ( .A(G116), .B(n1170), .ZN(G18) );
NAND3_X1 U897 ( .A1(n1036), .A2(n1176), .A3(n1204), .ZN(n1170) );
XNOR2_X1 U898 ( .A(G113), .B(n1169), .ZN(G15) );
NAND3_X1 U899 ( .A1(n1037), .A2(n1176), .A3(n1204), .ZN(n1169) );
NOR3_X1 U900 ( .A1(n1194), .A2(n1193), .A3(n1034), .ZN(n1204) );
INV_X1 U901 ( .A(n1028), .ZN(n1034) );
NOR2_X1 U902 ( .A1(n1032), .A2(n1031), .ZN(n1028) );
NAND2_X1 U903 ( .A1(n1208), .A2(n1209), .ZN(n1176) );
OR2_X1 U904 ( .A1(n1030), .A2(KEYINPUT14), .ZN(n1209) );
NAND2_X1 U905 ( .A1(n1207), .A2(n1206), .ZN(n1030) );
INV_X1 U906 ( .A(n1210), .ZN(n1207) );
NAND3_X1 U907 ( .A1(n1210), .A2(n1206), .A3(KEYINPUT14), .ZN(n1208) );
AND2_X1 U908 ( .A1(n1211), .A2(n1048), .ZN(n1037) );
XNOR2_X1 U909 ( .A(KEYINPUT17), .B(n1182), .ZN(n1211) );
XNOR2_X1 U910 ( .A(n1140), .B(n1212), .ZN(G12) );
NOR3_X1 U911 ( .A1(n1213), .A2(n1214), .A3(n1027), .ZN(n1212) );
INV_X1 U912 ( .A(n1184), .ZN(n1027) );
NOR2_X1 U913 ( .A1(n1210), .A2(n1206), .ZN(n1184) );
XNOR2_X1 U914 ( .A(n1215), .B(n1059), .ZN(n1206) );
NAND2_X1 U915 ( .A1(G217), .A2(n1216), .ZN(n1059) );
XNOR2_X1 U916 ( .A(n1061), .B(KEYINPUT55), .ZN(n1215) );
NOR2_X1 U917 ( .A1(n1107), .A2(G902), .ZN(n1061) );
INV_X1 U918 ( .A(n1104), .ZN(n1107) );
XNOR2_X1 U919 ( .A(n1217), .B(n1218), .ZN(n1104) );
XNOR2_X1 U920 ( .A(n1219), .B(n1082), .ZN(n1218) );
NOR2_X1 U921 ( .A1(KEYINPUT50), .A2(n1220), .ZN(n1219) );
XOR2_X1 U922 ( .A(n1221), .B(n1222), .Z(n1217) );
XNOR2_X1 U923 ( .A(n1140), .B(n1223), .ZN(n1222) );
NOR2_X1 U924 ( .A1(KEYINPUT48), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U925 ( .A(G137), .B(n1225), .ZN(n1224) );
AND3_X1 U926 ( .A1(G221), .A2(n1065), .A3(G234), .ZN(n1225) );
NAND2_X1 U927 ( .A1(n1226), .A2(KEYINPUT10), .ZN(n1221) );
XNOR2_X1 U928 ( .A(G128), .B(n1227), .ZN(n1226) );
XOR2_X1 U929 ( .A(n1054), .B(n1056), .Z(n1210) );
INV_X1 U930 ( .A(G472), .ZN(n1056) );
NAND3_X1 U931 ( .A1(n1228), .A2(n1229), .A3(n1159), .ZN(n1054) );
OR3_X1 U932 ( .A1(n1230), .A2(n1124), .A3(KEYINPUT21), .ZN(n1229) );
NAND2_X1 U933 ( .A1(n1231), .A2(KEYINPUT21), .ZN(n1228) );
XOR2_X1 U934 ( .A(n1124), .B(n1230), .Z(n1231) );
XNOR2_X1 U935 ( .A(G101), .B(n1232), .ZN(n1230) );
NOR2_X1 U936 ( .A1(KEYINPUT0), .A2(n1125), .ZN(n1232) );
NAND3_X1 U937 ( .A1(n1233), .A2(n1065), .A3(G210), .ZN(n1125) );
XOR2_X1 U938 ( .A(KEYINPUT30), .B(G237), .Z(n1233) );
XNOR2_X1 U939 ( .A(n1234), .B(n1235), .ZN(n1124) );
XOR2_X1 U940 ( .A(G113), .B(n1236), .Z(n1235) );
XOR2_X1 U941 ( .A(n1237), .B(n1238), .Z(n1234) );
NOR2_X1 U942 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
NOR2_X1 U943 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
AND3_X1 U944 ( .A1(n1241), .A2(n1227), .A3(G116), .ZN(n1239) );
INV_X1 U945 ( .A(KEYINPUT6), .ZN(n1241) );
INV_X1 U946 ( .A(n1173), .ZN(n1214) );
NOR4_X1 U947 ( .A1(n1194), .A2(n1192), .A3(n1193), .A4(n1031), .ZN(n1173) );
INV_X1 U948 ( .A(n1045), .ZN(n1031) );
NAND2_X1 U949 ( .A1(G221), .A2(n1216), .ZN(n1045) );
NAND2_X1 U950 ( .A1(G234), .A2(n1159), .ZN(n1216) );
AND2_X1 U951 ( .A1(n1017), .A2(n1243), .ZN(n1193) );
NAND3_X1 U952 ( .A1(n1097), .A2(n1202), .A3(G902), .ZN(n1243) );
NOR2_X1 U953 ( .A1(n1065), .A2(G898), .ZN(n1097) );
NAND3_X1 U954 ( .A1(n1041), .A2(n1202), .A3(G952), .ZN(n1017) );
NAND2_X1 U955 ( .A1(G234), .A2(G237), .ZN(n1202) );
XOR2_X1 U956 ( .A(G953), .B(KEYINPUT33), .Z(n1041) );
INV_X1 U957 ( .A(n1032), .ZN(n1192) );
XOR2_X1 U958 ( .A(n1053), .B(KEYINPUT49), .Z(n1032) );
XNOR2_X1 U959 ( .A(n1244), .B(G469), .ZN(n1053) );
NAND2_X1 U960 ( .A1(n1245), .A2(n1159), .ZN(n1244) );
XOR2_X1 U961 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U962 ( .A(n1147), .B(n1084), .Z(n1247) );
XNOR2_X1 U963 ( .A(n1248), .B(n1249), .ZN(n1084) );
XOR2_X1 U964 ( .A(KEYINPUT28), .B(n1250), .Z(n1249) );
NOR2_X1 U965 ( .A1(KEYINPUT16), .A2(n1220), .ZN(n1250) );
INV_X1 U966 ( .A(G146), .ZN(n1220) );
NAND2_X1 U967 ( .A1(KEYINPUT20), .A2(n1251), .ZN(n1248) );
XOR2_X1 U968 ( .A(n1237), .B(n1252), .Z(n1246) );
NOR2_X1 U969 ( .A1(KEYINPUT4), .A2(n1253), .ZN(n1252) );
XOR2_X1 U970 ( .A(n1131), .B(n1254), .Z(n1253) );
XNOR2_X1 U971 ( .A(n1140), .B(n1255), .ZN(n1254) );
NOR3_X1 U972 ( .A1(n1135), .A2(KEYINPUT57), .A3(G953), .ZN(n1255) );
INV_X1 U973 ( .A(G227), .ZN(n1135) );
XOR2_X1 U974 ( .A(G140), .B(KEYINPUT3), .Z(n1131) );
XNOR2_X1 U975 ( .A(n1141), .B(n1256), .ZN(n1237) );
INV_X1 U976 ( .A(n1085), .ZN(n1256) );
NAND2_X1 U977 ( .A1(n1257), .A2(n1258), .ZN(n1141) );
OR2_X1 U978 ( .A1(n1091), .A2(G137), .ZN(n1258) );
XOR2_X1 U979 ( .A(n1089), .B(KEYINPUT26), .Z(n1257) );
NAND2_X1 U980 ( .A1(G137), .A2(n1091), .ZN(n1089) );
INV_X1 U981 ( .A(n1042), .ZN(n1194) );
NOR2_X1 U982 ( .A1(n1052), .A2(n1016), .ZN(n1042) );
INV_X1 U983 ( .A(n1011), .ZN(n1016) );
NAND2_X1 U984 ( .A1(G214), .A2(n1259), .ZN(n1011) );
INV_X1 U985 ( .A(n1014), .ZN(n1052) );
XNOR2_X1 U986 ( .A(n1260), .B(n1261), .ZN(n1014) );
AND2_X1 U987 ( .A1(n1259), .A2(G210), .ZN(n1261) );
NAND2_X1 U988 ( .A1(n1262), .A2(n1159), .ZN(n1259) );
XOR2_X1 U989 ( .A(KEYINPUT62), .B(G237), .Z(n1262) );
NAND2_X1 U990 ( .A1(n1263), .A2(n1159), .ZN(n1260) );
INV_X1 U991 ( .A(G902), .ZN(n1159) );
XOR2_X1 U992 ( .A(n1264), .B(n1265), .Z(n1263) );
XNOR2_X1 U993 ( .A(n1156), .B(n1154), .ZN(n1265) );
XOR2_X1 U994 ( .A(G125), .B(KEYINPUT54), .Z(n1154) );
XNOR2_X1 U995 ( .A(n1236), .B(n1145), .ZN(n1156) );
XOR2_X1 U996 ( .A(G146), .B(n1251), .Z(n1236) );
XOR2_X1 U997 ( .A(G128), .B(KEYINPUT52), .Z(n1251) );
XOR2_X1 U998 ( .A(n1096), .B(n1266), .Z(n1264) );
NOR2_X1 U999 ( .A1(KEYINPUT42), .A2(n1158), .ZN(n1266) );
NAND2_X1 U1000 ( .A1(G224), .A2(n1065), .ZN(n1158) );
XOR2_X1 U1001 ( .A(n1267), .B(n1268), .Z(n1096) );
XNOR2_X1 U1002 ( .A(n1140), .B(n1269), .ZN(n1268) );
XOR2_X1 U1003 ( .A(n1242), .B(n1147), .Z(n1267) );
XOR2_X1 U1004 ( .A(G101), .B(n1270), .Z(n1147) );
XOR2_X1 U1005 ( .A(G107), .B(G104), .Z(n1270) );
XNOR2_X1 U1006 ( .A(G116), .B(n1227), .ZN(n1242) );
XOR2_X1 U1007 ( .A(G119), .B(KEYINPUT56), .Z(n1227) );
XNOR2_X1 U1008 ( .A(n1022), .B(KEYINPUT29), .ZN(n1213) );
INV_X1 U1009 ( .A(n1174), .ZN(n1022) );
NAND2_X1 U1010 ( .A1(n1271), .A2(n1272), .ZN(n1174) );
OR3_X1 U1011 ( .A1(n1182), .A2(n1048), .A3(KEYINPUT17), .ZN(n1272) );
INV_X1 U1012 ( .A(n1273), .ZN(n1182) );
NAND2_X1 U1013 ( .A1(KEYINPUT17), .A2(n1036), .ZN(n1271) );
NOR2_X1 U1014 ( .A1(n1048), .A2(n1273), .ZN(n1036) );
NOR2_X1 U1015 ( .A1(n1274), .A2(n1058), .ZN(n1273) );
NOR3_X1 U1016 ( .A1(G478), .A2(G902), .A3(n1110), .ZN(n1058) );
XOR2_X1 U1017 ( .A(n1057), .B(KEYINPUT47), .Z(n1274) );
AND2_X1 U1018 ( .A1(G478), .A2(n1275), .ZN(n1057) );
OR2_X1 U1019 ( .A1(n1110), .A2(G902), .ZN(n1275) );
NAND3_X1 U1020 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1110) );
OR2_X1 U1021 ( .A1(n1279), .A2(KEYINPUT63), .ZN(n1278) );
OR3_X1 U1022 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1277) );
INV_X1 U1023 ( .A(KEYINPUT63), .ZN(n1280) );
NAND2_X1 U1024 ( .A1(n1282), .A2(n1281), .ZN(n1276) );
NAND3_X1 U1025 ( .A1(n1283), .A2(n1065), .A3(G217), .ZN(n1281) );
INV_X1 U1026 ( .A(G953), .ZN(n1065) );
XOR2_X1 U1027 ( .A(KEYINPUT36), .B(G234), .Z(n1283) );
NAND2_X1 U1028 ( .A1(KEYINPUT38), .A2(n1279), .ZN(n1282) );
XNOR2_X1 U1029 ( .A(n1284), .B(n1285), .ZN(n1279) );
XOR2_X1 U1030 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U1031 ( .A(n1091), .B(G128), .ZN(n1287) );
INV_X1 U1032 ( .A(G134), .ZN(n1091) );
XNOR2_X1 U1033 ( .A(KEYINPUT2), .B(n1145), .ZN(n1286) );
INV_X1 U1034 ( .A(G143), .ZN(n1145) );
XNOR2_X1 U1035 ( .A(G107), .B(n1288), .ZN(n1284) );
XNOR2_X1 U1036 ( .A(G122), .B(n1289), .ZN(n1288) );
INV_X1 U1037 ( .A(G116), .ZN(n1289) );
XNOR2_X1 U1038 ( .A(n1290), .B(G475), .ZN(n1048) );
OR2_X1 U1039 ( .A1(n1116), .A2(G902), .ZN(n1290) );
XNOR2_X1 U1040 ( .A(n1291), .B(n1269), .ZN(n1116) );
XOR2_X1 U1041 ( .A(G113), .B(G122), .Z(n1269) );
XOR2_X1 U1042 ( .A(n1292), .B(G104), .Z(n1291) );
NAND3_X1 U1043 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(n1292) );
NAND2_X1 U1044 ( .A1(KEYINPUT46), .A2(n1296), .ZN(n1295) );
NAND3_X1 U1045 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1294) );
INV_X1 U1046 ( .A(KEYINPUT46), .ZN(n1298) );
OR2_X1 U1047 ( .A1(n1299), .A2(n1297), .ZN(n1293) );
NOR2_X1 U1048 ( .A1(KEYINPUT45), .A2(n1296), .ZN(n1297) );
XNOR2_X1 U1049 ( .A(G146), .B(n1082), .ZN(n1296) );
XNOR2_X1 U1050 ( .A(G125), .B(G140), .ZN(n1082) );
XOR2_X1 U1051 ( .A(n1085), .B(n1300), .Z(n1299) );
NOR3_X1 U1052 ( .A1(n1301), .A2(G953), .A3(G237), .ZN(n1300) );
INV_X1 U1053 ( .A(G214), .ZN(n1301) );
XOR2_X1 U1054 ( .A(G143), .B(n1134), .Z(n1085) );
XOR2_X1 U1055 ( .A(G131), .B(KEYINPUT11), .Z(n1134) );
INV_X1 U1056 ( .A(G110), .ZN(n1140) );
endmodule


