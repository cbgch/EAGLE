//Key = 1000111110111100101111100111001000111010010110111101000010000011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345;

XNOR2_X1 U744 ( .A(G107), .B(n1028), .ZN(G9) );
NOR2_X1 U745 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U746 ( .A1(n1031), .A2(n1032), .A3(G953), .A4(n1033), .ZN(n1030) );
NOR2_X1 U747 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U748 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR3_X1 U749 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NOR2_X1 U750 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR3_X1 U752 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1043) );
NOR2_X1 U753 ( .A1(KEYINPUT22), .A2(n1048), .ZN(n1047) );
XNOR2_X1 U754 ( .A(n1049), .B(KEYINPUT51), .ZN(n1045) );
NOR2_X1 U755 ( .A1(n1050), .A2(n1048), .ZN(n1041) );
NOR2_X1 U756 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U757 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1051) );
INV_X1 U758 ( .A(KEYINPUT22), .ZN(n1053) );
NOR3_X1 U759 ( .A1(n1044), .A2(n1056), .A3(n1048), .ZN(n1036) );
NOR2_X1 U760 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U761 ( .A1(n1059), .A2(n1038), .ZN(n1058) );
NOR2_X1 U762 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U764 ( .A1(n1064), .A2(n1040), .ZN(n1057) );
NOR2_X1 U765 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U766 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NAND3_X1 U767 ( .A1(n1069), .A2(G952), .A3(n1070), .ZN(n1031) );
NOR3_X1 U768 ( .A1(n1033), .A2(n1071), .A3(n1072), .ZN(n1029) );
NOR2_X1 U769 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
INV_X1 U770 ( .A(KEYINPUT10), .ZN(n1074) );
NOR2_X1 U771 ( .A1(G953), .A2(G952), .ZN(n1073) );
NOR2_X1 U772 ( .A1(KEYINPUT10), .A2(n1075), .ZN(n1071) );
AND4_X1 U773 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1033) );
NOR3_X1 U774 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
XOR2_X1 U775 ( .A(n1083), .B(KEYINPUT20), .Z(n1082) );
NOR2_X1 U776 ( .A1(G475), .A2(n1084), .ZN(n1081) );
NAND3_X1 U777 ( .A1(n1068), .A2(n1055), .A3(n1085), .ZN(n1080) );
NOR3_X1 U778 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1078) );
XOR2_X1 U779 ( .A(KEYINPUT45), .B(n1089), .Z(n1086) );
AND2_X1 U780 ( .A1(n1084), .A2(G475), .ZN(n1089) );
XNOR2_X1 U781 ( .A(n1090), .B(n1091), .ZN(n1077) );
XOR2_X1 U782 ( .A(n1092), .B(KEYINPUT29), .Z(n1076) );
XOR2_X1 U783 ( .A(n1093), .B(n1094), .Z(G72) );
NOR2_X1 U784 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U785 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
NOR2_X1 U786 ( .A1(KEYINPUT55), .A2(n1099), .ZN(n1093) );
XOR2_X1 U787 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR2_X1 U788 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U789 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U790 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U791 ( .A1(KEYINPUT54), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U792 ( .A(G131), .B(n1109), .ZN(n1104) );
NOR2_X1 U793 ( .A1(KEYINPUT3), .A2(n1110), .ZN(n1109) );
NAND3_X1 U794 ( .A1(n1111), .A2(n1096), .A3(KEYINPUT41), .ZN(n1100) );
XOR2_X1 U795 ( .A(n1112), .B(n1113), .Z(G69) );
XOR2_X1 U796 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U797 ( .A1(n1070), .A2(G953), .ZN(n1115) );
NOR2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
XOR2_X1 U799 ( .A(KEYINPUT44), .B(n1118), .Z(n1117) );
NOR3_X1 U800 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1118) );
NOR2_X1 U801 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U802 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
XOR2_X1 U803 ( .A(KEYINPUT58), .B(n1126), .Z(n1125) );
NOR3_X1 U804 ( .A1(n1127), .A2(n1126), .A3(n1124), .ZN(n1120) );
AND2_X1 U805 ( .A1(n1124), .A2(n1126), .ZN(n1119) );
XOR2_X1 U806 ( .A(n1128), .B(n1129), .Z(n1126) );
NOR2_X1 U807 ( .A1(KEYINPUT59), .A2(n1130), .ZN(n1129) );
INV_X1 U808 ( .A(KEYINPUT6), .ZN(n1124) );
NOR2_X1 U809 ( .A1(G898), .A2(n1131), .ZN(n1116) );
XOR2_X1 U810 ( .A(n1132), .B(KEYINPUT12), .Z(n1131) );
NOR2_X1 U811 ( .A1(n1133), .A2(n1096), .ZN(n1112) );
NOR2_X1 U812 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NOR2_X1 U813 ( .A1(n1136), .A2(n1137), .ZN(G66) );
XNOR2_X1 U814 ( .A(n1075), .B(KEYINPUT34), .ZN(n1137) );
XOR2_X1 U815 ( .A(n1138), .B(n1139), .Z(n1136) );
NAND2_X1 U816 ( .A1(n1140), .A2(n1141), .ZN(n1138) );
NOR2_X1 U817 ( .A1(n1075), .A2(n1142), .ZN(G63) );
XOR2_X1 U818 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U819 ( .A1(n1140), .A2(G478), .ZN(n1143) );
NOR3_X1 U820 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(G60) );
AND2_X1 U821 ( .A1(n1075), .A2(KEYINPUT4), .ZN(n1147) );
NOR3_X1 U822 ( .A1(KEYINPUT4), .A2(G953), .A3(G952), .ZN(n1146) );
XOR2_X1 U823 ( .A(n1148), .B(n1149), .Z(n1145) );
NAND2_X1 U824 ( .A1(n1140), .A2(G475), .ZN(n1148) );
XOR2_X1 U825 ( .A(n1150), .B(G104), .Z(G6) );
NAND2_X1 U826 ( .A1(KEYINPUT46), .A2(n1151), .ZN(n1150) );
NAND3_X1 U827 ( .A1(n1152), .A2(n1153), .A3(n1049), .ZN(n1151) );
NOR2_X1 U828 ( .A1(n1075), .A2(n1154), .ZN(G57) );
XOR2_X1 U829 ( .A(n1155), .B(n1156), .Z(n1154) );
XNOR2_X1 U830 ( .A(n1157), .B(n1158), .ZN(n1156) );
XOR2_X1 U831 ( .A(n1159), .B(n1160), .Z(n1155) );
NOR2_X1 U832 ( .A1(G101), .A2(KEYINPUT17), .ZN(n1160) );
NAND2_X1 U833 ( .A1(n1140), .A2(G472), .ZN(n1159) );
NOR2_X1 U834 ( .A1(n1075), .A2(n1161), .ZN(G54) );
XOR2_X1 U835 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U836 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U837 ( .A(n1166), .B(n1167), .Z(n1164) );
NAND3_X1 U838 ( .A1(n1140), .A2(G469), .A3(KEYINPUT56), .ZN(n1166) );
XOR2_X1 U839 ( .A(n1168), .B(n1169), .Z(n1162) );
XOR2_X1 U840 ( .A(KEYINPUT33), .B(KEYINPUT30), .Z(n1169) );
XNOR2_X1 U841 ( .A(n1170), .B(n1171), .ZN(n1168) );
NOR2_X1 U842 ( .A1(KEYINPUT2), .A2(n1172), .ZN(n1171) );
NOR2_X1 U843 ( .A1(KEYINPUT14), .A2(n1173), .ZN(n1170) );
XOR2_X1 U844 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U845 ( .A(n1176), .B(n1177), .Z(n1175) );
XNOR2_X1 U846 ( .A(n1178), .B(n1179), .ZN(n1174) );
NOR2_X1 U847 ( .A1(n1075), .A2(n1180), .ZN(G51) );
XOR2_X1 U848 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U849 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND2_X1 U850 ( .A1(KEYINPUT43), .A2(n1158), .ZN(n1184) );
NAND2_X1 U851 ( .A1(n1140), .A2(n1185), .ZN(n1183) );
XOR2_X1 U852 ( .A(KEYINPUT37), .B(G210), .Z(n1185) );
AND2_X1 U853 ( .A1(G902), .A2(n1186), .ZN(n1140) );
NAND2_X1 U854 ( .A1(n1187), .A2(n1069), .ZN(n1186) );
INV_X1 U855 ( .A(n1111), .ZN(n1069) );
NAND4_X1 U856 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1111) );
NOR4_X1 U857 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
NOR2_X1 U858 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NOR2_X1 U859 ( .A1(n1198), .A2(n1199), .ZN(n1194) );
AND2_X1 U860 ( .A1(n1200), .A2(n1201), .ZN(n1190) );
XNOR2_X1 U861 ( .A(n1070), .B(KEYINPUT27), .ZN(n1187) );
AND2_X1 U862 ( .A1(n1202), .A2(n1203), .ZN(n1070) );
AND4_X1 U863 ( .A1(n1028), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1203) );
NAND3_X1 U864 ( .A1(n1153), .A2(n1046), .A3(n1152), .ZN(n1028) );
NOR4_X1 U865 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1202) );
NOR2_X1 U866 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NOR2_X1 U867 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
XOR2_X1 U868 ( .A(n1215), .B(KEYINPUT21), .Z(n1214) );
NAND4_X1 U869 ( .A1(n1216), .A2(n1153), .A3(n1217), .A4(n1218), .ZN(n1215) );
XOR2_X1 U870 ( .A(KEYINPUT1), .B(n1219), .Z(n1217) );
NOR4_X1 U871 ( .A1(n1038), .A2(n1196), .A3(n1218), .A4(n1220), .ZN(n1213) );
INV_X1 U872 ( .A(KEYINPUT15), .ZN(n1220) );
INV_X1 U873 ( .A(n1216), .ZN(n1038) );
NOR3_X1 U874 ( .A1(n1196), .A2(KEYINPUT15), .A3(n1221), .ZN(n1209) );
NOR4_X1 U875 ( .A1(n1222), .A2(n1223), .A3(n1040), .A4(n1224), .ZN(n1208) );
INV_X1 U876 ( .A(n1153), .ZN(n1040) );
NAND2_X1 U877 ( .A1(n1225), .A2(n1218), .ZN(n1223) );
XNOR2_X1 U878 ( .A(KEYINPUT60), .B(n1226), .ZN(n1225) );
XNOR2_X1 U879 ( .A(n1052), .B(KEYINPUT57), .ZN(n1222) );
INV_X1 U880 ( .A(n1227), .ZN(n1207) );
NOR2_X1 U881 ( .A1(n1096), .A2(G952), .ZN(n1075) );
XNOR2_X1 U882 ( .A(n1228), .B(n1229), .ZN(G48) );
NOR2_X1 U883 ( .A1(n1199), .A2(n1230), .ZN(n1229) );
XNOR2_X1 U884 ( .A(KEYINPUT24), .B(n1231), .ZN(n1230) );
NAND4_X1 U885 ( .A1(n1062), .A2(n1049), .A3(n1232), .A4(n1088), .ZN(n1199) );
XNOR2_X1 U886 ( .A(G143), .B(n1189), .ZN(G45) );
NAND4_X1 U887 ( .A1(n1219), .A2(n1061), .A3(n1232), .A4(n1231), .ZN(n1189) );
XNOR2_X1 U888 ( .A(n1172), .B(n1193), .ZN(G42) );
AND2_X1 U889 ( .A1(n1233), .A2(n1234), .ZN(n1193) );
XOR2_X1 U890 ( .A(G137), .B(n1192), .Z(G39) );
AND3_X1 U891 ( .A1(n1062), .A2(n1235), .A3(n1233), .ZN(n1192) );
XOR2_X1 U892 ( .A(n1236), .B(n1237), .Z(G36) );
NOR2_X1 U893 ( .A1(KEYINPUT40), .A2(n1238), .ZN(n1237) );
NOR3_X1 U894 ( .A1(n1196), .A2(n1239), .A3(n1240), .ZN(n1236) );
NOR2_X1 U895 ( .A1(KEYINPUT0), .A2(n1241), .ZN(n1240) );
NOR3_X1 U896 ( .A1(n1044), .A2(n1066), .A3(n1198), .ZN(n1241) );
INV_X1 U897 ( .A(n1226), .ZN(n1066) );
AND2_X1 U898 ( .A1(n1197), .A2(KEYINPUT0), .ZN(n1239) );
INV_X1 U899 ( .A(n1233), .ZN(n1197) );
XNOR2_X1 U900 ( .A(G131), .B(n1201), .ZN(G33) );
NAND3_X1 U901 ( .A1(n1049), .A2(n1061), .A3(n1233), .ZN(n1201) );
NOR3_X1 U902 ( .A1(n1226), .A2(n1198), .A3(n1044), .ZN(n1233) );
NAND2_X1 U903 ( .A1(n1242), .A2(n1055), .ZN(n1044) );
XNOR2_X1 U904 ( .A(G128), .B(n1200), .ZN(G30) );
NAND4_X1 U905 ( .A1(n1062), .A2(n1046), .A3(n1243), .A4(n1232), .ZN(n1200) );
NOR2_X1 U906 ( .A1(n1198), .A2(n1063), .ZN(n1243) );
INV_X1 U907 ( .A(n1231), .ZN(n1198) );
XNOR2_X1 U908 ( .A(G101), .B(n1227), .ZN(G3) );
NAND3_X1 U909 ( .A1(n1244), .A2(n1152), .A3(n1061), .ZN(n1227) );
XNOR2_X1 U910 ( .A(G125), .B(n1188), .ZN(G27) );
NAND4_X1 U911 ( .A1(n1234), .A2(n1216), .A3(n1052), .A4(n1231), .ZN(n1188) );
NAND2_X1 U912 ( .A1(n1035), .A2(n1245), .ZN(n1231) );
NAND3_X1 U913 ( .A1(G902), .A2(n1246), .A3(n1102), .ZN(n1245) );
AND2_X1 U914 ( .A1(n1132), .A2(n1098), .ZN(n1102) );
INV_X1 U915 ( .A(G900), .ZN(n1098) );
NOR3_X1 U916 ( .A1(n1063), .A2(n1062), .A3(n1224), .ZN(n1234) );
XNOR2_X1 U917 ( .A(G122), .B(n1247), .ZN(G24) );
NAND3_X1 U918 ( .A1(n1248), .A2(n1153), .A3(n1219), .ZN(n1247) );
AND2_X1 U919 ( .A1(n1249), .A2(n1087), .ZN(n1219) );
NOR2_X1 U920 ( .A1(n1088), .A2(n1062), .ZN(n1153) );
XNOR2_X1 U921 ( .A(G119), .B(n1206), .ZN(G21) );
NAND3_X1 U922 ( .A1(n1062), .A2(n1235), .A3(n1248), .ZN(n1206) );
INV_X1 U923 ( .A(n1250), .ZN(n1062) );
XNOR2_X1 U924 ( .A(n1251), .B(n1252), .ZN(G18) );
NOR2_X1 U925 ( .A1(n1221), .A2(n1196), .ZN(n1252) );
NAND2_X1 U926 ( .A1(n1061), .A2(n1046), .ZN(n1196) );
NOR2_X1 U927 ( .A1(n1253), .A2(n1249), .ZN(n1046) );
XNOR2_X1 U928 ( .A(G113), .B(n1205), .ZN(G15) );
NAND3_X1 U929 ( .A1(n1248), .A2(n1061), .A3(n1049), .ZN(n1205) );
INV_X1 U930 ( .A(n1224), .ZN(n1049) );
NAND2_X1 U931 ( .A1(n1249), .A2(n1253), .ZN(n1224) );
INV_X1 U932 ( .A(n1087), .ZN(n1253) );
NOR2_X1 U933 ( .A1(n1250), .A2(n1088), .ZN(n1061) );
INV_X1 U934 ( .A(n1221), .ZN(n1248) );
NAND3_X1 U935 ( .A1(n1052), .A2(n1218), .A3(n1216), .ZN(n1221) );
NOR2_X1 U936 ( .A1(n1067), .A2(n1254), .ZN(n1216) );
INV_X1 U937 ( .A(n1068), .ZN(n1254) );
INV_X1 U938 ( .A(n1212), .ZN(n1052) );
XNOR2_X1 U939 ( .A(G110), .B(n1204), .ZN(G12) );
NAND3_X1 U940 ( .A1(n1152), .A2(n1250), .A3(n1235), .ZN(n1204) );
NOR2_X1 U941 ( .A1(n1048), .A2(n1063), .ZN(n1235) );
INV_X1 U942 ( .A(n1088), .ZN(n1063) );
XNOR2_X1 U943 ( .A(n1255), .B(n1141), .ZN(n1088) );
AND2_X1 U944 ( .A1(G217), .A2(n1256), .ZN(n1141) );
NAND2_X1 U945 ( .A1(n1139), .A2(n1257), .ZN(n1255) );
XNOR2_X1 U946 ( .A(n1258), .B(n1259), .ZN(n1139) );
XOR2_X1 U947 ( .A(G137), .B(n1260), .Z(n1259) );
NOR2_X1 U948 ( .A1(KEYINPUT42), .A2(n1261), .ZN(n1260) );
XOR2_X1 U949 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U950 ( .A(n1264), .B(n1167), .Z(n1263) );
XNOR2_X1 U951 ( .A(G119), .B(n1107), .ZN(n1264) );
XNOR2_X1 U952 ( .A(G128), .B(n1265), .ZN(n1262) );
XNOR2_X1 U953 ( .A(KEYINPUT52), .B(n1228), .ZN(n1265) );
NAND2_X1 U954 ( .A1(n1266), .A2(G221), .ZN(n1258) );
INV_X1 U955 ( .A(n1244), .ZN(n1048) );
NOR2_X1 U956 ( .A1(n1087), .A2(n1249), .ZN(n1244) );
XOR2_X1 U957 ( .A(n1084), .B(n1267), .Z(n1249) );
XOR2_X1 U958 ( .A(KEYINPUT63), .B(G475), .Z(n1267) );
NAND2_X1 U959 ( .A1(n1149), .A2(n1257), .ZN(n1084) );
XNOR2_X1 U960 ( .A(n1268), .B(n1269), .ZN(n1149) );
XOR2_X1 U961 ( .A(n1179), .B(n1107), .Z(n1269) );
XNOR2_X1 U962 ( .A(G125), .B(n1172), .ZN(n1107) );
XNOR2_X1 U963 ( .A(n1228), .B(n1270), .ZN(n1179) );
XNOR2_X1 U964 ( .A(n1271), .B(n1272), .ZN(n1268) );
NOR2_X1 U965 ( .A1(KEYINPUT31), .A2(n1273), .ZN(n1272) );
XNOR2_X1 U966 ( .A(G113), .B(n1274), .ZN(n1273) );
NAND2_X1 U967 ( .A1(KEYINPUT25), .A2(n1275), .ZN(n1274) );
NOR2_X1 U968 ( .A1(KEYINPUT50), .A2(n1276), .ZN(n1271) );
XOR2_X1 U969 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U970 ( .A(n1279), .B(G131), .ZN(n1278) );
INV_X1 U971 ( .A(G143), .ZN(n1279) );
NAND2_X1 U972 ( .A1(n1280), .A2(G214), .ZN(n1277) );
XNOR2_X1 U973 ( .A(n1281), .B(G478), .ZN(n1087) );
NAND2_X1 U974 ( .A1(n1144), .A2(n1257), .ZN(n1281) );
XNOR2_X1 U975 ( .A(n1282), .B(n1283), .ZN(n1144) );
XOR2_X1 U976 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U977 ( .A(G134), .B(G128), .ZN(n1285) );
NAND3_X1 U978 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1284) );
NAND2_X1 U979 ( .A1(G122), .A2(n1251), .ZN(n1288) );
NAND2_X1 U980 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
INV_X1 U981 ( .A(KEYINPUT26), .ZN(n1290) );
NAND2_X1 U982 ( .A1(n1291), .A2(n1275), .ZN(n1289) );
XNOR2_X1 U983 ( .A(KEYINPUT49), .B(G116), .ZN(n1291) );
NAND2_X1 U984 ( .A1(KEYINPUT26), .A2(n1292), .ZN(n1286) );
NAND2_X1 U985 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
OR2_X1 U986 ( .A1(G116), .A2(KEYINPUT49), .ZN(n1294) );
NAND3_X1 U987 ( .A1(G116), .A2(n1275), .A3(KEYINPUT49), .ZN(n1293) );
INV_X1 U988 ( .A(G122), .ZN(n1275) );
XNOR2_X1 U989 ( .A(n1176), .B(n1295), .ZN(n1282) );
AND2_X1 U990 ( .A1(G217), .A2(n1266), .ZN(n1295) );
AND2_X1 U991 ( .A1(G234), .A2(n1096), .ZN(n1266) );
XNOR2_X1 U992 ( .A(G143), .B(n1296), .ZN(n1176) );
XOR2_X1 U993 ( .A(n1297), .B(n1090), .Z(n1250) );
NAND2_X1 U994 ( .A1(n1298), .A2(n1257), .ZN(n1090) );
XOR2_X1 U995 ( .A(n1157), .B(n1299), .Z(n1298) );
XNOR2_X1 U996 ( .A(G101), .B(n1300), .ZN(n1299) );
NAND2_X1 U997 ( .A1(KEYINPUT38), .A2(n1158), .ZN(n1300) );
XOR2_X1 U998 ( .A(n1301), .B(n1302), .Z(n1157) );
XNOR2_X1 U999 ( .A(n1251), .B(n1303), .ZN(n1302) );
XNOR2_X1 U1000 ( .A(KEYINPUT9), .B(n1304), .ZN(n1303) );
INV_X1 U1001 ( .A(G116), .ZN(n1251) );
XOR2_X1 U1002 ( .A(n1305), .B(n1306), .Z(n1301) );
XNOR2_X1 U1003 ( .A(G113), .B(n1307), .ZN(n1306) );
NAND2_X1 U1004 ( .A1(n1280), .A2(G210), .ZN(n1307) );
NOR2_X1 U1005 ( .A1(G953), .A2(G237), .ZN(n1280) );
NAND2_X1 U1006 ( .A1(KEYINPUT5), .A2(n1091), .ZN(n1297) );
INV_X1 U1007 ( .A(G472), .ZN(n1091) );
AND2_X1 U1008 ( .A1(n1232), .A2(n1218), .ZN(n1152) );
NAND2_X1 U1009 ( .A1(n1035), .A2(n1308), .ZN(n1218) );
NAND4_X1 U1010 ( .A1(n1132), .A2(G902), .A3(n1246), .A4(n1135), .ZN(n1308) );
INV_X1 U1011 ( .A(G898), .ZN(n1135) );
XNOR2_X1 U1012 ( .A(G953), .B(KEYINPUT13), .ZN(n1132) );
NAND3_X1 U1013 ( .A1(n1246), .A2(n1096), .A3(G952), .ZN(n1035) );
INV_X1 U1014 ( .A(G953), .ZN(n1096) );
NAND2_X1 U1015 ( .A1(G237), .A2(G234), .ZN(n1246) );
NOR2_X1 U1016 ( .A1(n1212), .A2(n1226), .ZN(n1232) );
NAND2_X1 U1017 ( .A1(n1067), .A2(n1068), .ZN(n1226) );
NAND2_X1 U1018 ( .A1(G221), .A2(n1256), .ZN(n1068) );
NAND2_X1 U1019 ( .A1(G234), .A2(n1257), .ZN(n1256) );
NAND2_X1 U1020 ( .A1(n1083), .A2(n1085), .ZN(n1067) );
NAND2_X1 U1021 ( .A1(G469), .A2(n1309), .ZN(n1085) );
OR2_X1 U1022 ( .A1(n1309), .A2(G469), .ZN(n1083) );
NAND2_X1 U1023 ( .A1(n1310), .A2(n1257), .ZN(n1309) );
XOR2_X1 U1024 ( .A(n1311), .B(n1312), .Z(n1310) );
XNOR2_X1 U1025 ( .A(n1172), .B(n1313), .ZN(n1312) );
NOR2_X1 U1026 ( .A1(KEYINPUT32), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1027 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1028 ( .A(n1317), .B(n1270), .ZN(n1316) );
XNOR2_X1 U1029 ( .A(n1318), .B(n1178), .ZN(n1315) );
NAND2_X1 U1030 ( .A1(KEYINPUT11), .A2(n1108), .ZN(n1318) );
XNOR2_X1 U1031 ( .A(n1319), .B(n1177), .ZN(n1108) );
INV_X1 U1032 ( .A(G140), .ZN(n1172) );
XNOR2_X1 U1033 ( .A(n1165), .B(n1167), .ZN(n1311) );
XNOR2_X1 U1034 ( .A(n1305), .B(n1320), .ZN(n1165) );
NOR2_X1 U1035 ( .A1(G953), .A2(n1097), .ZN(n1320) );
INV_X1 U1036 ( .A(G227), .ZN(n1097) );
XOR2_X1 U1037 ( .A(G131), .B(n1110), .Z(n1305) );
XOR2_X1 U1038 ( .A(n1238), .B(G137), .Z(n1110) );
INV_X1 U1039 ( .A(G134), .ZN(n1238) );
NAND2_X1 U1040 ( .A1(n1054), .A2(n1055), .ZN(n1212) );
NAND2_X1 U1041 ( .A1(G214), .A2(n1321), .ZN(n1055) );
INV_X1 U1042 ( .A(n1242), .ZN(n1054) );
XNOR2_X1 U1043 ( .A(n1092), .B(KEYINPUT7), .ZN(n1242) );
XOR2_X1 U1044 ( .A(n1322), .B(n1323), .Z(n1092) );
AND2_X1 U1045 ( .A1(n1321), .A2(G210), .ZN(n1323) );
OR2_X1 U1046 ( .A1(G902), .A2(G237), .ZN(n1321) );
NAND2_X1 U1047 ( .A1(n1324), .A2(n1257), .ZN(n1322) );
INV_X1 U1048 ( .A(G902), .ZN(n1257) );
XNOR2_X1 U1049 ( .A(n1181), .B(n1325), .ZN(n1324) );
XNOR2_X1 U1050 ( .A(n1158), .B(KEYINPUT36), .ZN(n1325) );
XNOR2_X1 U1051 ( .A(n1326), .B(n1177), .ZN(n1158) );
XNOR2_X1 U1052 ( .A(n1327), .B(KEYINPUT8), .ZN(n1177) );
INV_X1 U1053 ( .A(G128), .ZN(n1327) );
NAND2_X1 U1054 ( .A1(KEYINPUT18), .A2(n1319), .ZN(n1326) );
XNOR2_X1 U1055 ( .A(G143), .B(n1228), .ZN(n1319) );
INV_X1 U1056 ( .A(G146), .ZN(n1228) );
XNOR2_X1 U1057 ( .A(n1328), .B(n1329), .ZN(n1181) );
XNOR2_X1 U1058 ( .A(n1330), .B(n1331), .ZN(n1329) );
XOR2_X1 U1059 ( .A(G125), .B(n1332), .Z(n1331) );
NOR2_X1 U1060 ( .A1(G953), .A2(n1134), .ZN(n1332) );
INV_X1 U1061 ( .A(G224), .ZN(n1134) );
INV_X1 U1062 ( .A(n1128), .ZN(n1330) );
XNOR2_X1 U1063 ( .A(n1333), .B(n1334), .ZN(n1128) );
NOR2_X1 U1064 ( .A1(KEYINPUT61), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1065 ( .A(n1336), .B(n1337), .Z(n1335) );
NOR2_X1 U1066 ( .A1(KEYINPUT53), .A2(n1338), .ZN(n1337) );
XNOR2_X1 U1067 ( .A(KEYINPUT47), .B(n1304), .ZN(n1338) );
INV_X1 U1068 ( .A(G119), .ZN(n1304) );
XNOR2_X1 U1069 ( .A(G116), .B(KEYINPUT35), .ZN(n1336) );
XNOR2_X1 U1070 ( .A(G113), .B(KEYINPUT16), .ZN(n1333) );
XNOR2_X1 U1071 ( .A(n1130), .B(n1127), .ZN(n1328) );
INV_X1 U1072 ( .A(n1123), .ZN(n1127) );
XOR2_X1 U1073 ( .A(G122), .B(n1167), .Z(n1123) );
XOR2_X1 U1074 ( .A(G110), .B(KEYINPUT19), .Z(n1167) );
XNOR2_X1 U1075 ( .A(n1339), .B(n1178), .ZN(n1130) );
INV_X1 U1076 ( .A(G101), .ZN(n1178) );
NAND2_X1 U1077 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
NAND2_X1 U1078 ( .A1(n1296), .A2(n1342), .ZN(n1341) );
INV_X1 U1079 ( .A(n1317), .ZN(n1296) );
XOR2_X1 U1080 ( .A(n1343), .B(KEYINPUT23), .Z(n1340) );
NAND2_X1 U1081 ( .A1(n1344), .A2(n1317), .ZN(n1343) );
XOR2_X1 U1082 ( .A(G107), .B(KEYINPUT62), .Z(n1317) );
XNOR2_X1 U1083 ( .A(n1345), .B(n1342), .ZN(n1344) );
INV_X1 U1084 ( .A(n1270), .ZN(n1342) );
XOR2_X1 U1085 ( .A(G104), .B(KEYINPUT39), .Z(n1270) );
XNOR2_X1 U1086 ( .A(KEYINPUT48), .B(KEYINPUT28), .ZN(n1345) );
endmodule


