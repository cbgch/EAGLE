//Key = 0000101100001111111111011000010011010100100111100111010011010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382;

XNOR2_X1 U742 ( .A(n1050), .B(n1051), .ZN(G9) );
NOR2_X1 U743 ( .A1(n1052), .A2(n1053), .ZN(G75) );
NOR4_X1 U744 ( .A1(n1054), .A2(n1055), .A3(G953), .A4(n1056), .ZN(n1053) );
NOR2_X1 U745 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U746 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U747 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U748 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR3_X1 U749 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NOR2_X1 U750 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U751 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR2_X1 U752 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR2_X1 U753 ( .A1(n1074), .A2(n1075), .ZN(n1068) );
NOR2_X1 U754 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U755 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
INV_X1 U756 ( .A(n1080), .ZN(n1065) );
NOR3_X1 U757 ( .A1(n1071), .A2(n1081), .A3(n1075), .ZN(n1063) );
NOR4_X1 U758 ( .A1(n1082), .A2(n1071), .A3(n1083), .A4(n1084), .ZN(n1059) );
NOR3_X1 U759 ( .A1(n1066), .A2(n1085), .A3(n1086), .ZN(n1084) );
NOR2_X1 U760 ( .A1(n1087), .A2(n1088), .ZN(n1083) );
NAND2_X1 U761 ( .A1(n1089), .A2(n1080), .ZN(n1082) );
NAND3_X1 U762 ( .A1(n1090), .A2(G952), .A3(n1091), .ZN(n1054) );
NOR3_X1 U763 ( .A1(n1092), .A2(G953), .A3(n1056), .ZN(n1052) );
AND4_X1 U764 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1056) );
NOR3_X1 U765 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
NAND3_X1 U766 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1097) );
XNOR2_X1 U767 ( .A(n1103), .B(n1104), .ZN(n1102) );
NAND2_X1 U768 ( .A1(n1105), .A2(n1106), .ZN(n1101) );
NAND2_X1 U769 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
NAND2_X1 U770 ( .A1(KEYINPUT10), .A2(n1109), .ZN(n1108) );
OR3_X1 U771 ( .A1(n1110), .A2(KEYINPUT10), .A3(n1106), .ZN(n1100) );
INV_X1 U772 ( .A(n1109), .ZN(n1110) );
XOR2_X1 U773 ( .A(n1107), .B(KEYINPUT26), .Z(n1109) );
NOR3_X1 U774 ( .A1(n1066), .A2(n1111), .A3(n1112), .ZN(n1095) );
NAND2_X1 U775 ( .A1(G475), .A2(n1113), .ZN(n1094) );
XOR2_X1 U776 ( .A(KEYINPUT11), .B(G952), .Z(n1092) );
XOR2_X1 U777 ( .A(n1114), .B(n1115), .Z(G72) );
NOR2_X1 U778 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NOR2_X1 U779 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XNOR2_X1 U780 ( .A(n1120), .B(KEYINPUT31), .ZN(n1119) );
NOR2_X1 U781 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
NOR3_X1 U782 ( .A1(n1122), .A2(n1121), .A3(n1120), .ZN(n1116) );
AND3_X1 U783 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1120) );
XNOR2_X1 U784 ( .A(G953), .B(KEYINPUT34), .ZN(n1125) );
NAND2_X1 U785 ( .A1(n1090), .A2(n1126), .ZN(n1124) );
INV_X1 U786 ( .A(KEYINPUT30), .ZN(n1126) );
NAND2_X1 U787 ( .A1(KEYINPUT30), .A2(n1127), .ZN(n1123) );
XOR2_X1 U788 ( .A(n1128), .B(n1129), .Z(n1122) );
XOR2_X1 U789 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U790 ( .A(n1132), .B(n1133), .Z(n1128) );
NOR2_X1 U791 ( .A1(G134), .A2(KEYINPUT55), .ZN(n1133) );
NAND2_X1 U792 ( .A1(G953), .A2(n1134), .ZN(n1114) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1134) );
XOR2_X1 U794 ( .A(n1135), .B(n1136), .Z(G69) );
XOR2_X1 U795 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U796 ( .A1(G953), .A2(n1139), .ZN(n1138) );
NAND2_X1 U797 ( .A1(G898), .A2(G224), .ZN(n1139) );
NAND2_X1 U798 ( .A1(n1140), .A2(n1141), .ZN(n1137) );
NAND2_X1 U799 ( .A1(G953), .A2(n1142), .ZN(n1141) );
XNOR2_X1 U800 ( .A(n1143), .B(n1144), .ZN(n1140) );
NAND2_X1 U801 ( .A1(n1145), .A2(n1146), .ZN(n1143) );
NAND2_X1 U802 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U803 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NAND2_X1 U804 ( .A1(KEYINPUT53), .A2(n1151), .ZN(n1150) );
INV_X1 U805 ( .A(n1152), .ZN(n1151) );
INV_X1 U806 ( .A(KEYINPUT5), .ZN(n1149) );
NAND2_X1 U807 ( .A1(n1152), .A2(n1153), .ZN(n1145) );
NAND2_X1 U808 ( .A1(KEYINPUT53), .A2(n1154), .ZN(n1153) );
OR2_X1 U809 ( .A1(n1147), .A2(KEYINPUT5), .ZN(n1154) );
NOR2_X1 U810 ( .A1(n1091), .A2(G953), .ZN(n1135) );
NOR2_X1 U811 ( .A1(n1155), .A2(n1156), .ZN(G66) );
NOR3_X1 U812 ( .A1(n1157), .A2(n1103), .A3(n1158), .ZN(n1156) );
NOR2_X1 U813 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U814 ( .A1(n1161), .A2(n1162), .ZN(n1159) );
XOR2_X1 U815 ( .A(KEYINPUT22), .B(n1163), .Z(n1157) );
NOR3_X1 U816 ( .A1(n1164), .A2(n1162), .A3(n1165), .ZN(n1163) );
NOR2_X1 U817 ( .A1(n1155), .A2(n1166), .ZN(G63) );
XOR2_X1 U818 ( .A(n1167), .B(n1168), .Z(n1166) );
NAND2_X1 U819 ( .A1(KEYINPUT23), .A2(n1169), .ZN(n1167) );
NAND2_X1 U820 ( .A1(n1170), .A2(G478), .ZN(n1169) );
NOR2_X1 U821 ( .A1(n1155), .A2(n1171), .ZN(G60) );
XOR2_X1 U822 ( .A(n1172), .B(n1173), .Z(n1171) );
NAND2_X1 U823 ( .A1(n1170), .A2(G475), .ZN(n1172) );
XOR2_X1 U824 ( .A(G104), .B(n1174), .Z(G6) );
NOR2_X1 U825 ( .A1(n1155), .A2(n1175), .ZN(G57) );
XOR2_X1 U826 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U827 ( .A1(KEYINPUT60), .A2(n1178), .ZN(n1177) );
NOR2_X1 U828 ( .A1(n1179), .A2(n1180), .ZN(n1176) );
XOR2_X1 U829 ( .A(n1181), .B(KEYINPUT35), .Z(n1180) );
NAND4_X1 U830 ( .A1(n1182), .A2(G472), .A3(G902), .A4(n1183), .ZN(n1181) );
XNOR2_X1 U831 ( .A(KEYINPUT2), .B(n1161), .ZN(n1182) );
NOR2_X1 U832 ( .A1(n1184), .A2(n1183), .ZN(n1179) );
NOR3_X1 U833 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
NOR2_X1 U834 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
INV_X1 U835 ( .A(KEYINPUT2), .ZN(n1189) );
NOR2_X1 U836 ( .A1(n1190), .A2(n1191), .ZN(n1188) );
NOR2_X1 U837 ( .A1(KEYINPUT2), .A2(n1170), .ZN(n1186) );
NOR2_X1 U838 ( .A1(n1155), .A2(n1192), .ZN(G54) );
XOR2_X1 U839 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U840 ( .A(n1195), .B(KEYINPUT29), .Z(n1194) );
NAND2_X1 U841 ( .A1(n1196), .A2(KEYINPUT49), .ZN(n1195) );
XOR2_X1 U842 ( .A(n1197), .B(n1198), .Z(n1196) );
XNOR2_X1 U843 ( .A(G110), .B(n1199), .ZN(n1198) );
NAND2_X1 U844 ( .A1(KEYINPUT13), .A2(n1200), .ZN(n1199) );
XOR2_X1 U845 ( .A(n1201), .B(n1202), .Z(n1197) );
NAND2_X1 U846 ( .A1(KEYINPUT20), .A2(G140), .ZN(n1201) );
NAND2_X1 U847 ( .A1(n1170), .A2(G469), .ZN(n1193) );
NOR2_X1 U848 ( .A1(n1155), .A2(n1203), .ZN(G51) );
XOR2_X1 U849 ( .A(n1204), .B(n1205), .Z(n1203) );
NOR2_X1 U850 ( .A1(n1106), .A2(n1164), .ZN(n1205) );
INV_X1 U851 ( .A(n1170), .ZN(n1164) );
NOR2_X1 U852 ( .A1(n1190), .A2(n1161), .ZN(n1170) );
INV_X1 U853 ( .A(n1191), .ZN(n1161) );
NAND2_X1 U854 ( .A1(n1091), .A2(n1206), .ZN(n1191) );
XOR2_X1 U855 ( .A(KEYINPUT1), .B(n1090), .Z(n1206) );
NOR3_X1 U856 ( .A1(n1127), .A2(n1207), .A3(n1208), .ZN(n1090) );
OR3_X1 U857 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1208) );
NAND4_X1 U858 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1127) );
NAND2_X1 U859 ( .A1(n1216), .A2(n1217), .ZN(n1212) );
AND4_X1 U860 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1091) );
NOR4_X1 U861 ( .A1(n1222), .A2(n1051), .A3(n1223), .A4(n1224), .ZN(n1221) );
AND2_X1 U862 ( .A1(n1073), .A2(n1225), .ZN(n1051) );
AND4_X1 U863 ( .A1(n1086), .A2(n1226), .A3(n1077), .A4(n1089), .ZN(n1222) );
NOR2_X1 U864 ( .A1(n1174), .A2(n1227), .ZN(n1220) );
NOR4_X1 U865 ( .A1(n1228), .A2(n1229), .A3(n1071), .A4(n1230), .ZN(n1227) );
XNOR2_X1 U866 ( .A(n1231), .B(KEYINPUT0), .ZN(n1229) );
AND2_X1 U867 ( .A1(n1058), .A2(n1232), .ZN(n1228) );
AND2_X1 U868 ( .A1(n1072), .A2(n1225), .ZN(n1174) );
NOR3_X1 U869 ( .A1(n1233), .A2(n1062), .A3(n1234), .ZN(n1225) );
INV_X1 U870 ( .A(n1087), .ZN(n1062) );
NAND2_X1 U871 ( .A1(n1235), .A2(KEYINPUT46), .ZN(n1204) );
XNOR2_X1 U872 ( .A(n1236), .B(n1237), .ZN(n1235) );
XOR2_X1 U873 ( .A(n1238), .B(n1239), .Z(n1237) );
NAND2_X1 U874 ( .A1(KEYINPUT50), .A2(n1240), .ZN(n1239) );
NOR2_X1 U875 ( .A1(n1241), .A2(G952), .ZN(n1155) );
XNOR2_X1 U876 ( .A(G146), .B(n1213), .ZN(G48) );
NAND2_X1 U877 ( .A1(n1242), .A2(n1072), .ZN(n1213) );
XNOR2_X1 U878 ( .A(G143), .B(n1243), .ZN(G45) );
NAND2_X1 U879 ( .A1(KEYINPUT32), .A2(n1244), .ZN(n1243) );
INV_X1 U880 ( .A(n1214), .ZN(n1244) );
NAND3_X1 U881 ( .A1(n1245), .A2(n1085), .A3(n1246), .ZN(n1214) );
NOR3_X1 U882 ( .A1(n1081), .A2(n1247), .A3(n1248), .ZN(n1246) );
XNOR2_X1 U883 ( .A(n1249), .B(n1215), .ZN(G42) );
NAND3_X1 U884 ( .A1(n1072), .A2(n1086), .A3(n1216), .ZN(n1215) );
XNOR2_X1 U885 ( .A(G140), .B(KEYINPUT4), .ZN(n1249) );
XOR2_X1 U886 ( .A(G137), .B(n1250), .Z(G39) );
NOR4_X1 U887 ( .A1(n1251), .A2(n1252), .A3(KEYINPUT38), .A4(n1253), .ZN(n1250) );
NOR2_X1 U888 ( .A1(KEYINPUT16), .A2(n1254), .ZN(n1252) );
NOR3_X1 U889 ( .A1(n1255), .A2(n1089), .A3(n1256), .ZN(n1254) );
AND2_X1 U890 ( .A1(n1230), .A2(KEYINPUT16), .ZN(n1251) );
INV_X1 U891 ( .A(n1217), .ZN(n1230) );
XNOR2_X1 U892 ( .A(G134), .B(n1257), .ZN(G36) );
NAND2_X1 U893 ( .A1(KEYINPUT24), .A2(n1209), .ZN(n1257) );
AND3_X1 U894 ( .A1(n1085), .A2(n1073), .A3(n1216), .ZN(n1209) );
XOR2_X1 U895 ( .A(G131), .B(n1211), .Z(G33) );
AND3_X1 U896 ( .A1(n1085), .A2(n1072), .A3(n1216), .ZN(n1211) );
INV_X1 U897 ( .A(n1253), .ZN(n1216) );
NAND3_X1 U898 ( .A1(n1080), .A2(n1088), .A3(n1245), .ZN(n1253) );
XNOR2_X1 U899 ( .A(n1258), .B(n1207), .ZN(G30) );
AND2_X1 U900 ( .A1(n1242), .A2(n1073), .ZN(n1207) );
AND4_X1 U901 ( .A1(n1245), .A2(n1231), .A3(n1259), .A4(n1098), .ZN(n1242) );
AND2_X1 U902 ( .A1(n1077), .A2(n1260), .ZN(n1245) );
XNOR2_X1 U903 ( .A(G101), .B(n1218), .ZN(G3) );
NAND4_X1 U904 ( .A1(n1085), .A2(n1089), .A3(n1077), .A4(n1226), .ZN(n1218) );
XNOR2_X1 U905 ( .A(n1261), .B(n1262), .ZN(G27) );
NAND2_X1 U906 ( .A1(n1263), .A2(n1264), .ZN(n1261) );
NAND2_X1 U907 ( .A1(n1210), .A2(n1265), .ZN(n1264) );
INV_X1 U908 ( .A(KEYINPUT25), .ZN(n1265) );
NOR2_X1 U909 ( .A1(n1266), .A2(n1081), .ZN(n1210) );
INV_X1 U910 ( .A(n1231), .ZN(n1081) );
NAND3_X1 U911 ( .A1(n1231), .A2(n1266), .A3(KEYINPUT25), .ZN(n1263) );
NAND4_X1 U912 ( .A1(n1072), .A2(n1267), .A3(n1086), .A4(n1260), .ZN(n1266) );
NAND2_X1 U913 ( .A1(n1058), .A2(n1268), .ZN(n1260) );
NAND3_X1 U914 ( .A1(G902), .A2(n1269), .A3(n1121), .ZN(n1268) );
NOR2_X1 U915 ( .A1(n1241), .A2(G900), .ZN(n1121) );
XNOR2_X1 U916 ( .A(G122), .B(n1219), .ZN(G24) );
NAND4_X1 U917 ( .A1(n1270), .A2(n1087), .A3(n1099), .A4(n1271), .ZN(n1219) );
XNOR2_X1 U918 ( .A(G119), .B(n1272), .ZN(G21) );
NOR2_X1 U919 ( .A1(n1273), .A2(KEYINPUT42), .ZN(n1272) );
AND2_X1 U920 ( .A1(n1270), .A2(n1217), .ZN(n1273) );
NOR3_X1 U921 ( .A1(n1255), .A2(n1256), .A3(n1075), .ZN(n1217) );
INV_X1 U922 ( .A(n1089), .ZN(n1075) );
INV_X1 U923 ( .A(n1098), .ZN(n1256) );
XOR2_X1 U924 ( .A(G116), .B(n1224), .Z(G18) );
AND3_X1 U925 ( .A1(n1270), .A2(n1073), .A3(n1085), .ZN(n1224) );
NOR2_X1 U926 ( .A1(n1271), .A2(n1248), .ZN(n1073) );
INV_X1 U927 ( .A(n1099), .ZN(n1248) );
NAND3_X1 U928 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(G15) );
NAND2_X1 U929 ( .A1(KEYINPUT39), .A2(n1277), .ZN(n1276) );
OR3_X1 U930 ( .A1(n1277), .A2(KEYINPUT39), .A3(G113), .ZN(n1275) );
NAND2_X1 U931 ( .A1(G113), .A2(n1278), .ZN(n1274) );
NAND2_X1 U932 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
INV_X1 U933 ( .A(KEYINPUT39), .ZN(n1280) );
XNOR2_X1 U934 ( .A(n1223), .B(KEYINPUT12), .ZN(n1279) );
INV_X1 U935 ( .A(n1277), .ZN(n1223) );
NAND3_X1 U936 ( .A1(n1072), .A2(n1270), .A3(n1085), .ZN(n1277) );
AND2_X1 U937 ( .A1(n1281), .A2(n1098), .ZN(n1085) );
XNOR2_X1 U938 ( .A(n1259), .B(KEYINPUT48), .ZN(n1281) );
NOR2_X1 U939 ( .A1(n1071), .A2(n1233), .ZN(n1270) );
INV_X1 U940 ( .A(n1267), .ZN(n1071) );
NOR2_X1 U941 ( .A1(n1078), .A2(n1112), .ZN(n1267) );
INV_X1 U942 ( .A(n1079), .ZN(n1112) );
NOR2_X1 U943 ( .A1(n1099), .A2(n1247), .ZN(n1072) );
INV_X1 U944 ( .A(n1271), .ZN(n1247) );
XNOR2_X1 U945 ( .A(G110), .B(n1282), .ZN(G12) );
NAND4_X1 U946 ( .A1(n1283), .A2(n1089), .A3(n1226), .A4(n1086), .ZN(n1282) );
NAND2_X1 U947 ( .A1(n1284), .A2(n1285), .ZN(n1086) );
OR3_X1 U948 ( .A1(n1255), .A2(n1098), .A3(KEYINPUT47), .ZN(n1285) );
INV_X1 U949 ( .A(n1259), .ZN(n1255) );
NAND2_X1 U950 ( .A1(KEYINPUT47), .A2(n1087), .ZN(n1284) );
NOR2_X1 U951 ( .A1(n1098), .A2(n1259), .ZN(n1087) );
XOR2_X1 U952 ( .A(n1286), .B(n1287), .Z(n1259) );
INV_X1 U953 ( .A(n1103), .ZN(n1287) );
NOR2_X1 U954 ( .A1(n1160), .A2(G902), .ZN(n1103) );
INV_X1 U955 ( .A(n1165), .ZN(n1160) );
XNOR2_X1 U956 ( .A(n1288), .B(n1289), .ZN(n1165) );
XNOR2_X1 U957 ( .A(G137), .B(n1290), .ZN(n1289) );
NAND2_X1 U958 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
NAND2_X1 U959 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U960 ( .A(KEYINPUT57), .B(n1295), .Z(n1291) );
NOR2_X1 U961 ( .A1(n1293), .A2(n1294), .ZN(n1295) );
INV_X1 U962 ( .A(G110), .ZN(n1294) );
XNOR2_X1 U963 ( .A(G119), .B(n1296), .ZN(n1293) );
NOR2_X1 U964 ( .A1(KEYINPUT54), .A2(n1258), .ZN(n1296) );
XOR2_X1 U965 ( .A(n1297), .B(n1298), .Z(n1288) );
NOR2_X1 U966 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
INV_X1 U967 ( .A(G221), .ZN(n1300) );
NAND2_X1 U968 ( .A1(n1301), .A2(n1302), .ZN(n1297) );
NAND2_X1 U969 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
XOR2_X1 U970 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U971 ( .A(KEYINPUT56), .B(KEYINPUT33), .Z(n1306) );
XOR2_X1 U972 ( .A(KEYINPUT44), .B(n1307), .Z(n1301) );
NOR2_X1 U973 ( .A1(n1303), .A2(n1305), .ZN(n1307) );
XOR2_X1 U974 ( .A(n1130), .B(KEYINPUT45), .Z(n1305) );
XNOR2_X1 U975 ( .A(G125), .B(n1308), .ZN(n1130) );
XNOR2_X1 U976 ( .A(G146), .B(KEYINPUT58), .ZN(n1303) );
NAND2_X1 U977 ( .A1(KEYINPUT17), .A2(n1104), .ZN(n1286) );
INV_X1 U978 ( .A(n1162), .ZN(n1104) );
NAND2_X1 U979 ( .A1(G217), .A2(n1309), .ZN(n1162) );
XOR2_X1 U980 ( .A(n1310), .B(n1185), .Z(n1098) );
INV_X1 U981 ( .A(G472), .ZN(n1185) );
NAND2_X1 U982 ( .A1(n1311), .A2(n1190), .ZN(n1310) );
XOR2_X1 U983 ( .A(n1178), .B(n1183), .Z(n1311) );
XNOR2_X1 U984 ( .A(n1312), .B(n1313), .ZN(n1183) );
XNOR2_X1 U985 ( .A(G113), .B(n1314), .ZN(n1313) );
NAND2_X1 U986 ( .A1(KEYINPUT21), .A2(n1315), .ZN(n1314) );
XOR2_X1 U987 ( .A(KEYINPUT52), .B(n1316), .Z(n1315) );
XNOR2_X1 U988 ( .A(n1200), .B(n1240), .ZN(n1312) );
AND2_X1 U989 ( .A1(n1317), .A2(n1318), .ZN(n1178) );
NAND2_X1 U990 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
NAND2_X1 U991 ( .A1(G210), .A2(n1321), .ZN(n1319) );
NAND3_X1 U992 ( .A1(G210), .A2(n1321), .A3(G101), .ZN(n1317) );
INV_X1 U993 ( .A(n1233), .ZN(n1226) );
NAND2_X1 U994 ( .A1(n1231), .A2(n1322), .ZN(n1233) );
NAND2_X1 U995 ( .A1(n1058), .A2(n1232), .ZN(n1322) );
NAND4_X1 U996 ( .A1(G953), .A2(G902), .A3(n1269), .A4(n1142), .ZN(n1232) );
INV_X1 U997 ( .A(G898), .ZN(n1142) );
NAND3_X1 U998 ( .A1(n1269), .A2(n1241), .A3(G952), .ZN(n1058) );
NAND2_X1 U999 ( .A1(n1323), .A2(G234), .ZN(n1269) );
XNOR2_X1 U1000 ( .A(G237), .B(KEYINPUT18), .ZN(n1323) );
NOR2_X1 U1001 ( .A1(n1080), .A2(n1066), .ZN(n1231) );
INV_X1 U1002 ( .A(n1088), .ZN(n1066) );
NAND2_X1 U1003 ( .A1(G214), .A2(n1324), .ZN(n1088) );
XOR2_X1 U1004 ( .A(n1325), .B(n1106), .Z(n1080) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1324), .ZN(n1106) );
NAND2_X1 U1006 ( .A1(n1326), .A2(n1190), .ZN(n1324) );
INV_X1 U1007 ( .A(G237), .ZN(n1326) );
NAND2_X1 U1008 ( .A1(KEYINPUT43), .A2(n1107), .ZN(n1325) );
NAND2_X1 U1009 ( .A1(n1327), .A2(n1190), .ZN(n1107) );
XNOR2_X1 U1010 ( .A(n1328), .B(n1238), .ZN(n1327) );
NAND2_X1 U1011 ( .A1(n1329), .A2(n1330), .ZN(n1238) );
NAND2_X1 U1012 ( .A1(n1331), .A2(n1144), .ZN(n1330) );
XOR2_X1 U1013 ( .A(n1332), .B(KEYINPUT41), .Z(n1329) );
NAND2_X1 U1014 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
INV_X1 U1015 ( .A(n1144), .ZN(n1334) );
XOR2_X1 U1016 ( .A(G110), .B(n1335), .Z(n1144) );
XOR2_X1 U1017 ( .A(KEYINPUT8), .B(G122), .Z(n1335) );
XOR2_X1 U1018 ( .A(n1331), .B(KEYINPUT14), .Z(n1333) );
XNOR2_X1 U1019 ( .A(n1152), .B(n1147), .ZN(n1331) );
XNOR2_X1 U1020 ( .A(n1336), .B(n1316), .ZN(n1147) );
XOR2_X1 U1021 ( .A(G116), .B(G119), .Z(n1316) );
XNOR2_X1 U1022 ( .A(G113), .B(KEYINPUT15), .ZN(n1336) );
XNOR2_X1 U1023 ( .A(n1337), .B(n1338), .ZN(n1152) );
XOR2_X1 U1024 ( .A(n1339), .B(KEYINPUT28), .Z(n1337) );
NAND2_X1 U1025 ( .A1(n1340), .A2(n1050), .ZN(n1339) );
XNOR2_X1 U1026 ( .A(KEYINPUT6), .B(KEYINPUT37), .ZN(n1340) );
NOR2_X1 U1027 ( .A1(KEYINPUT3), .A2(n1341), .ZN(n1328) );
XNOR2_X1 U1028 ( .A(n1240), .B(n1342), .ZN(n1341) );
INV_X1 U1029 ( .A(n1236), .ZN(n1342) );
XOR2_X1 U1030 ( .A(G125), .B(n1343), .Z(n1236) );
AND2_X1 U1031 ( .A1(n1241), .A2(G224), .ZN(n1343) );
XNOR2_X1 U1032 ( .A(n1344), .B(n1345), .ZN(n1240) );
XNOR2_X1 U1033 ( .A(G128), .B(KEYINPUT36), .ZN(n1344) );
NOR2_X1 U1034 ( .A1(n1099), .A2(n1271), .ZN(n1089) );
NAND3_X1 U1035 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1271) );
INV_X1 U1036 ( .A(n1111), .ZN(n1348) );
NOR2_X1 U1037 ( .A1(n1113), .A2(G475), .ZN(n1111) );
OR2_X1 U1038 ( .A1(n1349), .A2(G475), .ZN(n1347) );
NAND3_X1 U1039 ( .A1(n1113), .A2(n1349), .A3(G475), .ZN(n1346) );
INV_X1 U1040 ( .A(KEYINPUT9), .ZN(n1349) );
NAND2_X1 U1041 ( .A1(n1173), .A2(n1190), .ZN(n1113) );
XNOR2_X1 U1042 ( .A(n1350), .B(n1351), .ZN(n1173) );
XOR2_X1 U1043 ( .A(n1352), .B(n1353), .Z(n1351) );
XOR2_X1 U1044 ( .A(G122), .B(G113), .Z(n1353) );
XOR2_X1 U1045 ( .A(KEYINPUT61), .B(G131), .Z(n1352) );
XOR2_X1 U1046 ( .A(n1354), .B(n1355), .Z(n1350) );
XNOR2_X1 U1047 ( .A(n1356), .B(n1345), .ZN(n1355) );
NAND2_X1 U1048 ( .A1(G214), .A2(n1321), .ZN(n1356) );
NOR2_X1 U1049 ( .A1(G953), .A2(G237), .ZN(n1321) );
XOR2_X1 U1050 ( .A(n1357), .B(G104), .Z(n1354) );
NAND2_X1 U1051 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
NAND2_X1 U1052 ( .A1(G140), .A2(n1262), .ZN(n1359) );
XOR2_X1 U1053 ( .A(KEYINPUT62), .B(n1360), .Z(n1358) );
NOR2_X1 U1054 ( .A1(G140), .A2(n1262), .ZN(n1360) );
INV_X1 U1055 ( .A(G125), .ZN(n1262) );
XNOR2_X1 U1056 ( .A(n1361), .B(G478), .ZN(n1099) );
OR2_X1 U1057 ( .A1(n1168), .A2(G902), .ZN(n1361) );
XNOR2_X1 U1058 ( .A(n1362), .B(n1363), .ZN(n1168) );
XOR2_X1 U1059 ( .A(n1364), .B(n1365), .Z(n1363) );
XOR2_X1 U1060 ( .A(G122), .B(G116), .Z(n1365) );
XOR2_X1 U1061 ( .A(G143), .B(G134), .Z(n1364) );
XOR2_X1 U1062 ( .A(n1366), .B(n1367), .Z(n1362) );
NOR2_X1 U1063 ( .A1(n1299), .A2(n1368), .ZN(n1367) );
INV_X1 U1064 ( .A(G217), .ZN(n1368) );
NAND2_X1 U1065 ( .A1(G234), .A2(n1241), .ZN(n1299) );
XNOR2_X1 U1066 ( .A(n1369), .B(n1050), .ZN(n1366) );
NAND2_X1 U1067 ( .A1(KEYINPUT7), .A2(n1258), .ZN(n1369) );
INV_X1 U1068 ( .A(G128), .ZN(n1258) );
XNOR2_X1 U1069 ( .A(n1077), .B(KEYINPUT51), .ZN(n1283) );
INV_X1 U1070 ( .A(n1234), .ZN(n1077) );
NAND2_X1 U1071 ( .A1(n1078), .A2(n1079), .ZN(n1234) );
NAND2_X1 U1072 ( .A1(G221), .A2(n1309), .ZN(n1079) );
NAND2_X1 U1073 ( .A1(G234), .A2(n1190), .ZN(n1309) );
XOR2_X1 U1074 ( .A(n1093), .B(KEYINPUT63), .Z(n1078) );
XOR2_X1 U1075 ( .A(n1370), .B(G469), .Z(n1093) );
NAND2_X1 U1076 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
XNOR2_X1 U1077 ( .A(KEYINPUT40), .B(n1190), .ZN(n1372) );
INV_X1 U1078 ( .A(G902), .ZN(n1190) );
XOR2_X1 U1079 ( .A(n1373), .B(n1374), .Z(n1371) );
XNOR2_X1 U1080 ( .A(n1308), .B(G110), .ZN(n1374) );
INV_X1 U1081 ( .A(G140), .ZN(n1308) );
XNOR2_X1 U1082 ( .A(n1202), .B(n1200), .ZN(n1373) );
XOR2_X1 U1083 ( .A(G134), .B(n1131), .Z(n1200) );
XOR2_X1 U1084 ( .A(G131), .B(G137), .Z(n1131) );
XNOR2_X1 U1085 ( .A(n1375), .B(n1376), .ZN(n1202) );
XOR2_X1 U1086 ( .A(n1377), .B(n1338), .Z(n1376) );
XNOR2_X1 U1087 ( .A(G104), .B(n1320), .ZN(n1338) );
INV_X1 U1088 ( .A(G101), .ZN(n1320) );
AND2_X1 U1089 ( .A1(n1241), .A2(G227), .ZN(n1377) );
INV_X1 U1090 ( .A(G953), .ZN(n1241) );
XOR2_X1 U1091 ( .A(n1132), .B(n1378), .Z(n1375) );
XNOR2_X1 U1092 ( .A(KEYINPUT59), .B(n1050), .ZN(n1378) );
INV_X1 U1093 ( .A(G107), .ZN(n1050) );
NAND2_X1 U1094 ( .A1(n1379), .A2(n1380), .ZN(n1132) );
NAND2_X1 U1095 ( .A1(G128), .A2(n1381), .ZN(n1380) );
XOR2_X1 U1096 ( .A(KEYINPUT19), .B(n1382), .Z(n1379) );
NOR2_X1 U1097 ( .A1(G128), .A2(n1381), .ZN(n1382) );
XOR2_X1 U1098 ( .A(KEYINPUT27), .B(n1345), .Z(n1381) );
XOR2_X1 U1099 ( .A(G143), .B(G146), .Z(n1345) );
endmodule


