//Key = 1100011110100011001000000010100101110101101010011111110101010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392;

XOR2_X1 U761 ( .A(n1055), .B(n1056), .Z(G9) );
NOR3_X1 U762 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
XOR2_X1 U763 ( .A(KEYINPUT1), .B(n1060), .Z(n1059) );
NAND3_X1 U764 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1057) );
XOR2_X1 U765 ( .A(KEYINPUT63), .B(n1064), .Z(n1061) );
NAND2_X1 U766 ( .A1(KEYINPUT6), .A2(n1065), .ZN(n1055) );
NOR2_X1 U767 ( .A1(n1066), .A2(n1067), .ZN(G75) );
NOR4_X1 U768 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1067) );
NOR2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U770 ( .A(n1074), .B(KEYINPUT56), .Z(n1072) );
NOR3_X1 U771 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1070) );
NAND4_X1 U772 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1074) );
NAND3_X1 U773 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1068) );
NAND3_X1 U774 ( .A1(n1084), .A2(n1085), .A3(n1077), .ZN(n1083) );
INV_X1 U775 ( .A(n1086), .ZN(n1077) );
NAND2_X1 U776 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NAND3_X1 U777 ( .A1(n1080), .A2(n1089), .A3(n1078), .ZN(n1088) );
OR2_X1 U778 ( .A1(n1090), .A2(n1063), .ZN(n1089) );
NAND2_X1 U779 ( .A1(n1079), .A2(n1091), .ZN(n1087) );
NAND2_X1 U780 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U781 ( .A1(n1078), .A2(n1094), .ZN(n1093) );
OR2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U783 ( .A1(n1080), .A2(n1097), .ZN(n1092) );
NAND2_X1 U784 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
OR2_X1 U785 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
AND3_X1 U786 ( .A1(n1081), .A2(n1082), .A3(n1102), .ZN(n1066) );
NAND4_X1 U787 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1081) );
AND4_X1 U788 ( .A1(n1107), .A2(n1108), .A3(n1101), .A4(n1075), .ZN(n1106) );
AND3_X1 U789 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1107) );
NAND3_X1 U790 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
INV_X1 U791 ( .A(KEYINPUT54), .ZN(n1114) );
OR2_X1 U792 ( .A1(G469), .A2(KEYINPUT39), .ZN(n1113) );
NAND2_X1 U793 ( .A1(KEYINPUT39), .A2(n1115), .ZN(n1112) );
OR2_X1 U794 ( .A1(n1116), .A2(G469), .ZN(n1115) );
NAND2_X1 U795 ( .A1(n1117), .A2(n1118), .ZN(n1110) );
NAND2_X1 U796 ( .A1(n1119), .A2(n1116), .ZN(n1109) );
NAND2_X1 U797 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U798 ( .A1(KEYINPUT54), .A2(KEYINPUT39), .ZN(n1121) );
NOR3_X1 U799 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1105) );
XOR2_X1 U800 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U801 ( .A1(n1127), .A2(KEYINPUT19), .ZN(n1126) );
NOR2_X1 U802 ( .A1(n1128), .A2(n1129), .ZN(n1123) );
XOR2_X1 U803 ( .A(n1130), .B(n1131), .Z(n1122) );
XOR2_X1 U804 ( .A(KEYINPUT42), .B(G472), .Z(n1131) );
XOR2_X1 U805 ( .A(KEYINPUT52), .B(n1132), .Z(n1104) );
NOR2_X1 U806 ( .A1(n1117), .A2(n1118), .ZN(n1132) );
XOR2_X1 U807 ( .A(KEYINPUT37), .B(n1133), .Z(n1117) );
XOR2_X1 U808 ( .A(n1134), .B(n1135), .Z(G72) );
NOR2_X1 U809 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XOR2_X1 U810 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U811 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U812 ( .A(n1142), .B(G131), .Z(n1138) );
NAND4_X1 U813 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1134) );
INV_X1 U814 ( .A(n1136), .ZN(n1146) );
NAND2_X1 U815 ( .A1(G953), .A2(n1147), .ZN(n1144) );
XOR2_X1 U816 ( .A(n1148), .B(n1149), .Z(G69) );
XOR2_X1 U817 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U818 ( .A1(G953), .A2(n1152), .ZN(n1151) );
NAND2_X1 U819 ( .A1(G898), .A2(G224), .ZN(n1152) );
NAND2_X1 U820 ( .A1(n1153), .A2(n1154), .ZN(n1150) );
NAND2_X1 U821 ( .A1(G953), .A2(n1155), .ZN(n1154) );
XOR2_X1 U822 ( .A(n1156), .B(n1157), .Z(n1153) );
NAND2_X1 U823 ( .A1(KEYINPUT50), .A2(n1158), .ZN(n1156) );
NOR2_X1 U824 ( .A1(n1159), .A2(G953), .ZN(n1148) );
NOR2_X1 U825 ( .A1(n1160), .A2(n1161), .ZN(G66) );
NOR2_X1 U826 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U827 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U828 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NOR2_X1 U829 ( .A1(KEYINPUT61), .A2(n1168), .ZN(n1164) );
AND2_X1 U830 ( .A1(n1168), .A2(KEYINPUT61), .ZN(n1162) );
NOR2_X1 U831 ( .A1(n1160), .A2(n1169), .ZN(G63) );
NOR3_X1 U832 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1169) );
NOR3_X1 U833 ( .A1(n1173), .A2(n1133), .A3(n1167), .ZN(n1172) );
NOR2_X1 U834 ( .A1(n1174), .A2(n1175), .ZN(n1171) );
AND2_X1 U835 ( .A1(n1069), .A2(G478), .ZN(n1174) );
NOR3_X1 U836 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(G60) );
NOR3_X1 U837 ( .A1(n1179), .A2(n1082), .A3(n1102), .ZN(n1178) );
INV_X1 U838 ( .A(G952), .ZN(n1102) );
AND2_X1 U839 ( .A1(n1179), .A2(n1160), .ZN(n1177) );
INV_X1 U840 ( .A(KEYINPUT9), .ZN(n1179) );
XOR2_X1 U841 ( .A(n1180), .B(n1181), .Z(n1176) );
NOR2_X1 U842 ( .A1(n1182), .A2(n1167), .ZN(n1180) );
INV_X1 U843 ( .A(G475), .ZN(n1182) );
XNOR2_X1 U844 ( .A(G104), .B(n1183), .ZN(G6) );
NOR2_X1 U845 ( .A1(n1160), .A2(n1184), .ZN(G57) );
XOR2_X1 U846 ( .A(n1185), .B(n1186), .Z(n1184) );
XNOR2_X1 U847 ( .A(n1187), .B(n1188), .ZN(n1186) );
XNOR2_X1 U848 ( .A(n1189), .B(G101), .ZN(n1188) );
XOR2_X1 U849 ( .A(n1190), .B(n1191), .Z(n1185) );
XOR2_X1 U850 ( .A(n1192), .B(n1193), .Z(n1191) );
NOR2_X1 U851 ( .A1(n1194), .A2(n1167), .ZN(n1193) );
INV_X1 U852 ( .A(G472), .ZN(n1194) );
NOR2_X1 U853 ( .A1(KEYINPUT12), .A2(n1195), .ZN(n1192) );
XOR2_X1 U854 ( .A(KEYINPUT16), .B(n1196), .Z(n1195) );
NOR2_X1 U855 ( .A1(n1160), .A2(n1197), .ZN(G54) );
XOR2_X1 U856 ( .A(n1198), .B(n1199), .Z(n1197) );
XOR2_X1 U857 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U858 ( .A(n1202), .B(n1203), .Z(n1201) );
NOR2_X1 U859 ( .A1(G140), .A2(KEYINPUT30), .ZN(n1203) );
NOR2_X1 U860 ( .A1(n1120), .A2(n1167), .ZN(n1202) );
INV_X1 U861 ( .A(G469), .ZN(n1120) );
XOR2_X1 U862 ( .A(n1204), .B(n1205), .Z(n1198) );
NOR2_X1 U863 ( .A1(KEYINPUT21), .A2(n1206), .ZN(n1205) );
XOR2_X1 U864 ( .A(n1207), .B(n1208), .Z(n1206) );
NAND2_X1 U865 ( .A1(KEYINPUT28), .A2(n1209), .ZN(n1207) );
XNOR2_X1 U866 ( .A(n1189), .B(KEYINPUT2), .ZN(n1204) );
NOR2_X1 U867 ( .A1(n1160), .A2(n1210), .ZN(G51) );
XOR2_X1 U868 ( .A(n1211), .B(n1212), .Z(n1210) );
XNOR2_X1 U869 ( .A(n1213), .B(n1214), .ZN(n1212) );
NOR2_X1 U870 ( .A1(n1215), .A2(n1167), .ZN(n1214) );
NAND2_X1 U871 ( .A1(G902), .A2(n1069), .ZN(n1167) );
NAND3_X1 U872 ( .A1(n1143), .A2(n1159), .A3(n1216), .ZN(n1069) );
XOR2_X1 U873 ( .A(n1145), .B(KEYINPUT4), .Z(n1216) );
NAND2_X1 U874 ( .A1(n1217), .A2(n1084), .ZN(n1145) );
AND4_X1 U875 ( .A1(n1218), .A2(n1183), .A3(n1219), .A4(n1220), .ZN(n1159) );
NOR4_X1 U876 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1220) );
NOR2_X1 U877 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
INV_X1 U878 ( .A(KEYINPUT31), .ZN(n1226) );
NOR2_X1 U879 ( .A1(KEYINPUT41), .A2(n1227), .ZN(n1223) );
NOR2_X1 U880 ( .A1(n1228), .A2(n1229), .ZN(n1222) );
NOR2_X1 U881 ( .A1(n1230), .A2(n1231), .ZN(n1228) );
AND2_X1 U882 ( .A1(n1232), .A2(n1079), .ZN(n1231) );
NOR3_X1 U883 ( .A1(n1233), .A2(KEYINPUT31), .A3(n1096), .ZN(n1230) );
NOR3_X1 U884 ( .A1(n1234), .A2(n1235), .A3(n1073), .ZN(n1221) );
AND4_X1 U885 ( .A1(n1062), .A2(n1060), .A3(n1063), .A4(n1236), .ZN(n1235) );
NOR3_X1 U886 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1219) );
NAND4_X1 U887 ( .A1(n1090), .A2(n1240), .A3(n1080), .A4(n1062), .ZN(n1183) );
NAND3_X1 U888 ( .A1(n1241), .A2(n1062), .A3(n1063), .ZN(n1218) );
NAND2_X1 U889 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND4_X1 U890 ( .A1(KEYINPUT41), .A2(n1078), .A3(n1096), .A4(n1073), .ZN(n1243) );
NAND3_X1 U891 ( .A1(n1240), .A2(n1234), .A3(n1236), .ZN(n1242) );
XOR2_X1 U892 ( .A(n1058), .B(KEYINPUT5), .Z(n1236) );
INV_X1 U893 ( .A(KEYINPUT36), .ZN(n1234) );
AND4_X1 U894 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1247), .ZN(n1143) );
AND4_X1 U895 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1247) );
NAND3_X1 U896 ( .A1(n1252), .A2(n1063), .A3(n1084), .ZN(n1246) );
NAND2_X1 U897 ( .A1(n1253), .A2(n1254), .ZN(n1244) );
INV_X1 U898 ( .A(n1255), .ZN(n1254) );
XOR2_X1 U899 ( .A(n1256), .B(KEYINPUT7), .Z(n1253) );
XOR2_X1 U900 ( .A(n1257), .B(n1258), .Z(n1211) );
NOR2_X1 U901 ( .A1(n1082), .A2(G952), .ZN(n1160) );
XNOR2_X1 U902 ( .A(n1245), .B(n1259), .ZN(G48) );
NOR2_X1 U903 ( .A1(KEYINPUT43), .A2(n1260), .ZN(n1259) );
NAND2_X1 U904 ( .A1(n1090), .A2(n1261), .ZN(n1245) );
XOR2_X1 U905 ( .A(n1262), .B(n1251), .Z(G45) );
NAND3_X1 U906 ( .A1(n1240), .A2(n1096), .A3(n1263), .ZN(n1251) );
AND3_X1 U907 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1263) );
XOR2_X1 U908 ( .A(G140), .B(n1267), .Z(G42) );
NOR3_X1 U909 ( .A1(n1268), .A2(KEYINPUT45), .A3(n1269), .ZN(n1267) );
XOR2_X1 U910 ( .A(KEYINPUT14), .B(n1217), .Z(n1268) );
AND4_X1 U911 ( .A1(n1090), .A2(n1060), .A3(n1095), .A4(n1265), .ZN(n1217) );
XOR2_X1 U912 ( .A(n1270), .B(n1250), .Z(G39) );
NAND4_X1 U913 ( .A1(n1232), .A2(n1265), .A3(n1060), .A4(n1271), .ZN(n1250) );
NOR2_X1 U914 ( .A1(n1269), .A2(n1272), .ZN(n1271) );
XNOR2_X1 U915 ( .A(G134), .B(n1273), .ZN(G36) );
NAND3_X1 U916 ( .A1(n1252), .A2(n1063), .A3(n1274), .ZN(n1273) );
XOR2_X1 U917 ( .A(n1269), .B(KEYINPUT10), .Z(n1274) );
INV_X1 U918 ( .A(n1084), .ZN(n1269) );
XOR2_X1 U919 ( .A(n1275), .B(n1249), .Z(G33) );
NAND3_X1 U920 ( .A1(n1084), .A2(n1252), .A3(n1090), .ZN(n1249) );
AND3_X1 U921 ( .A1(n1060), .A2(n1265), .A3(n1096), .ZN(n1252) );
INV_X1 U922 ( .A(n1098), .ZN(n1060) );
NOR2_X1 U923 ( .A1(n1076), .A2(n1276), .ZN(n1084) );
XOR2_X1 U924 ( .A(n1277), .B(n1248), .Z(G30) );
NAND2_X1 U925 ( .A1(n1261), .A2(n1063), .ZN(n1248) );
AND3_X1 U926 ( .A1(n1232), .A2(n1265), .A3(n1240), .ZN(n1261) );
XOR2_X1 U927 ( .A(G101), .B(n1237), .Z(G3) );
AND2_X1 U928 ( .A1(n1278), .A2(n1096), .ZN(n1237) );
XOR2_X1 U929 ( .A(G125), .B(n1279), .Z(G27) );
NOR2_X1 U930 ( .A1(n1256), .A2(n1255), .ZN(n1279) );
NAND4_X1 U931 ( .A1(n1090), .A2(n1064), .A3(n1095), .A4(n1265), .ZN(n1255) );
NAND2_X1 U932 ( .A1(n1086), .A2(n1280), .ZN(n1265) );
NAND3_X1 U933 ( .A1(G902), .A2(n1281), .A3(n1136), .ZN(n1280) );
NOR2_X1 U934 ( .A1(G900), .A2(n1082), .ZN(n1136) );
XOR2_X1 U935 ( .A(G122), .B(n1239), .Z(G24) );
NOR4_X1 U936 ( .A1(n1229), .A2(n1058), .A3(n1282), .A4(n1283), .ZN(n1239) );
XNOR2_X1 U937 ( .A(G119), .B(n1284), .ZN(G21) );
NAND4_X1 U938 ( .A1(n1232), .A2(n1062), .A3(n1285), .A4(n1286), .ZN(n1284) );
NOR2_X1 U939 ( .A1(n1272), .A2(n1256), .ZN(n1286) );
INV_X1 U940 ( .A(n1079), .ZN(n1272) );
XOR2_X1 U941 ( .A(KEYINPUT11), .B(n1064), .Z(n1285) );
NAND2_X1 U942 ( .A1(n1287), .A2(n1288), .ZN(n1232) );
NAND3_X1 U943 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1288) );
NAND2_X1 U944 ( .A1(KEYINPUT20), .A2(n1096), .ZN(n1287) );
XNOR2_X1 U945 ( .A(G116), .B(n1227), .ZN(G18) );
NAND3_X1 U946 ( .A1(n1096), .A2(n1063), .A3(n1292), .ZN(n1227) );
NOR2_X1 U947 ( .A1(n1293), .A2(n1282), .ZN(n1063) );
XNOR2_X1 U948 ( .A(G113), .B(n1225), .ZN(G15) );
NAND3_X1 U949 ( .A1(n1090), .A2(n1096), .A3(n1292), .ZN(n1225) );
INV_X1 U950 ( .A(n1229), .ZN(n1292) );
NAND3_X1 U951 ( .A1(n1064), .A2(n1062), .A3(n1078), .ZN(n1229) );
INV_X1 U952 ( .A(n1256), .ZN(n1078) );
NAND2_X1 U953 ( .A1(n1294), .A2(n1295), .ZN(n1256) );
INV_X1 U954 ( .A(n1100), .ZN(n1294) );
INV_X1 U955 ( .A(n1073), .ZN(n1064) );
NOR2_X1 U956 ( .A1(n1296), .A2(n1289), .ZN(n1096) );
INV_X1 U957 ( .A(n1233), .ZN(n1090) );
NAND2_X1 U958 ( .A1(n1266), .A2(n1282), .ZN(n1233) );
INV_X1 U959 ( .A(n1264), .ZN(n1282) );
INV_X1 U960 ( .A(n1283), .ZN(n1266) );
XOR2_X1 U961 ( .A(n1293), .B(KEYINPUT44), .Z(n1283) );
XOR2_X1 U962 ( .A(G110), .B(n1238), .Z(G12) );
AND2_X1 U963 ( .A1(n1278), .A2(n1095), .ZN(n1238) );
NAND2_X1 U964 ( .A1(n1297), .A2(n1298), .ZN(n1095) );
NAND3_X1 U965 ( .A1(n1296), .A2(n1289), .A3(n1291), .ZN(n1298) );
INV_X1 U966 ( .A(KEYINPUT20), .ZN(n1291) );
INV_X1 U967 ( .A(n1103), .ZN(n1289) );
NAND2_X1 U968 ( .A1(KEYINPUT20), .A2(n1080), .ZN(n1297) );
INV_X1 U969 ( .A(n1058), .ZN(n1080) );
NAND2_X1 U970 ( .A1(n1103), .A2(n1296), .ZN(n1058) );
INV_X1 U971 ( .A(n1290), .ZN(n1296) );
XOR2_X1 U972 ( .A(n1130), .B(n1299), .Z(n1290) );
NOR2_X1 U973 ( .A1(G472), .A2(KEYINPUT24), .ZN(n1299) );
NAND2_X1 U974 ( .A1(n1300), .A2(n1301), .ZN(n1130) );
XOR2_X1 U975 ( .A(n1302), .B(n1303), .Z(n1300) );
XOR2_X1 U976 ( .A(n1304), .B(G101), .Z(n1303) );
NAND2_X1 U977 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
OR2_X1 U978 ( .A1(n1307), .A2(n1190), .ZN(n1306) );
XOR2_X1 U979 ( .A(n1308), .B(KEYINPUT3), .Z(n1305) );
NAND2_X1 U980 ( .A1(n1190), .A2(n1307), .ZN(n1308) );
XOR2_X1 U981 ( .A(n1189), .B(n1196), .Z(n1307) );
XOR2_X1 U982 ( .A(n1309), .B(KEYINPUT8), .Z(n1190) );
NAND2_X1 U983 ( .A1(KEYINPUT33), .A2(n1187), .ZN(n1302) );
AND3_X1 U984 ( .A1(G210), .A2(n1082), .A3(n1310), .ZN(n1187) );
XOR2_X1 U985 ( .A(n1311), .B(KEYINPUT23), .Z(n1310) );
XOR2_X1 U986 ( .A(n1312), .B(n1313), .Z(n1103) );
NOR2_X1 U987 ( .A1(n1166), .A2(n1314), .ZN(n1313) );
XNOR2_X1 U988 ( .A(KEYINPUT13), .B(n1315), .ZN(n1314) );
INV_X1 U989 ( .A(G217), .ZN(n1166) );
OR2_X1 U990 ( .A1(n1168), .A2(G902), .ZN(n1312) );
XOR2_X1 U991 ( .A(n1316), .B(n1317), .Z(n1168) );
XOR2_X1 U992 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U993 ( .A(n1270), .B(G110), .Z(n1319) );
INV_X1 U994 ( .A(G137), .ZN(n1270) );
NAND3_X1 U995 ( .A1(G221), .A2(n1082), .A3(n1320), .ZN(n1318) );
XNOR2_X1 U996 ( .A(G234), .B(KEYINPUT53), .ZN(n1320) );
XOR2_X1 U997 ( .A(n1321), .B(n1322), .Z(n1316) );
NAND2_X1 U998 ( .A1(KEYINPUT40), .A2(n1323), .ZN(n1321) );
XOR2_X1 U999 ( .A(G128), .B(G119), .Z(n1323) );
AND3_X1 U1000 ( .A1(n1240), .A2(n1062), .A3(n1079), .ZN(n1278) );
NOR2_X1 U1001 ( .A1(n1293), .A2(n1264), .ZN(n1079) );
XOR2_X1 U1002 ( .A(n1324), .B(n1170), .Z(n1264) );
INV_X1 U1003 ( .A(n1118), .ZN(n1170) );
NAND2_X1 U1004 ( .A1(n1173), .A2(n1301), .ZN(n1118) );
INV_X1 U1005 ( .A(n1175), .ZN(n1173) );
XOR2_X1 U1006 ( .A(n1325), .B(n1326), .Z(n1175) );
XOR2_X1 U1007 ( .A(n1327), .B(n1328), .Z(n1326) );
XOR2_X1 U1008 ( .A(G122), .B(G116), .Z(n1328) );
XOR2_X1 U1009 ( .A(KEYINPUT29), .B(G134), .Z(n1327) );
XOR2_X1 U1010 ( .A(n1329), .B(n1330), .Z(n1325) );
AND3_X1 U1011 ( .A1(G217), .A2(n1082), .A3(G234), .ZN(n1330) );
XOR2_X1 U1012 ( .A(n1065), .B(n1331), .Z(n1329) );
NOR2_X1 U1013 ( .A1(KEYINPUT60), .A2(n1332), .ZN(n1331) );
XOR2_X1 U1014 ( .A(n1277), .B(G143), .Z(n1332) );
INV_X1 U1015 ( .A(G128), .ZN(n1277) );
NAND2_X1 U1016 ( .A1(KEYINPUT0), .A2(n1133), .ZN(n1324) );
INV_X1 U1017 ( .A(G478), .ZN(n1133) );
NAND3_X1 U1018 ( .A1(n1333), .A2(n1334), .A3(n1108), .ZN(n1293) );
NAND2_X1 U1019 ( .A1(n1128), .A2(n1129), .ZN(n1108) );
NAND2_X1 U1020 ( .A1(n1129), .A2(n1335), .ZN(n1334) );
OR3_X1 U1021 ( .A1(n1129), .A2(n1128), .A3(n1335), .ZN(n1333) );
INV_X1 U1022 ( .A(KEYINPUT59), .ZN(n1335) );
NOR2_X1 U1023 ( .A1(n1181), .A2(G902), .ZN(n1128) );
XNOR2_X1 U1024 ( .A(n1336), .B(n1337), .ZN(n1181) );
XOR2_X1 U1025 ( .A(n1338), .B(n1339), .Z(n1337) );
XOR2_X1 U1026 ( .A(G122), .B(G113), .Z(n1339) );
XOR2_X1 U1027 ( .A(G143), .B(G131), .Z(n1338) );
XNOR2_X1 U1028 ( .A(n1322), .B(n1340), .ZN(n1336) );
XNOR2_X1 U1029 ( .A(n1341), .B(n1342), .ZN(n1340) );
AND3_X1 U1030 ( .A1(G214), .A2(n1082), .A3(n1311), .ZN(n1341) );
XNOR2_X1 U1031 ( .A(n1260), .B(n1141), .ZN(n1322) );
XOR2_X1 U1032 ( .A(G125), .B(G140), .Z(n1141) );
XNOR2_X1 U1033 ( .A(G475), .B(KEYINPUT32), .ZN(n1129) );
NAND2_X1 U1034 ( .A1(n1086), .A2(n1343), .ZN(n1062) );
NAND4_X1 U1035 ( .A1(G953), .A2(G902), .A3(n1281), .A4(n1155), .ZN(n1343) );
INV_X1 U1036 ( .A(G898), .ZN(n1155) );
NAND3_X1 U1037 ( .A1(n1281), .A2(n1082), .A3(G952), .ZN(n1086) );
NAND2_X1 U1038 ( .A1(G237), .A2(G234), .ZN(n1281) );
NOR2_X1 U1039 ( .A1(n1098), .A2(n1073), .ZN(n1240) );
NAND2_X1 U1040 ( .A1(n1344), .A2(n1076), .ZN(n1073) );
XNOR2_X1 U1041 ( .A(n1125), .B(n1127), .ZN(n1076) );
INV_X1 U1042 ( .A(n1215), .ZN(n1127) );
NAND2_X1 U1043 ( .A1(G210), .A2(n1345), .ZN(n1215) );
NAND2_X1 U1044 ( .A1(n1346), .A2(n1301), .ZN(n1125) );
XOR2_X1 U1045 ( .A(n1347), .B(n1348), .Z(n1346) );
INV_X1 U1046 ( .A(n1257), .ZN(n1348) );
XNOR2_X1 U1047 ( .A(n1158), .B(n1157), .ZN(n1257) );
AND2_X1 U1048 ( .A1(n1349), .A2(n1350), .ZN(n1157) );
NAND2_X1 U1049 ( .A1(G110), .A2(n1351), .ZN(n1350) );
XOR2_X1 U1050 ( .A(KEYINPUT49), .B(n1352), .Z(n1349) );
NOR2_X1 U1051 ( .A1(G110), .A2(n1351), .ZN(n1352) );
INV_X1 U1052 ( .A(G122), .ZN(n1351) );
XNOR2_X1 U1053 ( .A(n1353), .B(n1354), .ZN(n1158) );
XNOR2_X1 U1054 ( .A(KEYINPUT27), .B(n1342), .ZN(n1354) );
XOR2_X1 U1055 ( .A(n1309), .B(n1355), .Z(n1353) );
INV_X1 U1056 ( .A(n1356), .ZN(n1355) );
XNOR2_X1 U1057 ( .A(G113), .B(n1357), .ZN(n1309) );
XOR2_X1 U1058 ( .A(G119), .B(G116), .Z(n1357) );
NAND3_X1 U1059 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1347) );
NAND2_X1 U1060 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
NAND2_X1 U1061 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
XNOR2_X1 U1062 ( .A(KEYINPUT57), .B(n1213), .ZN(n1363) );
NAND3_X1 U1063 ( .A1(n1365), .A2(n1213), .A3(n1364), .ZN(n1359) );
INV_X1 U1064 ( .A(n1361), .ZN(n1365) );
XNOR2_X1 U1065 ( .A(n1258), .B(KEYINPUT25), .ZN(n1361) );
XOR2_X1 U1066 ( .A(n1196), .B(G125), .Z(n1258) );
XNOR2_X1 U1067 ( .A(n1366), .B(G128), .ZN(n1196) );
NAND4_X1 U1068 ( .A1(n1367), .A2(n1368), .A3(n1369), .A4(n1370), .ZN(n1366) );
NAND3_X1 U1069 ( .A1(n1371), .A2(n1262), .A3(n1372), .ZN(n1370) );
INV_X1 U1070 ( .A(KEYINPUT15), .ZN(n1372) );
OR2_X1 U1071 ( .A1(KEYINPUT48), .A2(G146), .ZN(n1371) );
NAND3_X1 U1072 ( .A1(G143), .A2(n1373), .A3(KEYINPUT15), .ZN(n1369) );
NAND2_X1 U1073 ( .A1(KEYINPUT48), .A2(n1260), .ZN(n1373) );
NAND3_X1 U1074 ( .A1(n1374), .A2(n1260), .A3(n1375), .ZN(n1368) );
INV_X1 U1075 ( .A(KEYINPUT58), .ZN(n1375) );
XOR2_X1 U1076 ( .A(KEYINPUT48), .B(G143), .Z(n1374) );
NAND2_X1 U1077 ( .A1(KEYINPUT58), .A2(G146), .ZN(n1367) );
OR2_X1 U1078 ( .A1(n1213), .A2(n1364), .ZN(n1358) );
INV_X1 U1079 ( .A(KEYINPUT22), .ZN(n1364) );
NAND2_X1 U1080 ( .A1(G224), .A2(n1082), .ZN(n1213) );
INV_X1 U1081 ( .A(G953), .ZN(n1082) );
XOR2_X1 U1082 ( .A(KEYINPUT51), .B(n1276), .Z(n1344) );
XNOR2_X1 U1083 ( .A(n1075), .B(KEYINPUT46), .ZN(n1276) );
NAND2_X1 U1084 ( .A1(G214), .A2(n1345), .ZN(n1075) );
NAND2_X1 U1085 ( .A1(n1311), .A2(n1301), .ZN(n1345) );
INV_X1 U1086 ( .A(G237), .ZN(n1311) );
NAND2_X1 U1087 ( .A1(n1100), .A2(n1295), .ZN(n1098) );
XNOR2_X1 U1088 ( .A(n1101), .B(KEYINPUT47), .ZN(n1295) );
NAND2_X1 U1089 ( .A1(G221), .A2(n1315), .ZN(n1101) );
NAND2_X1 U1090 ( .A1(G234), .A2(n1301), .ZN(n1315) );
XNOR2_X1 U1091 ( .A(n1116), .B(G469), .ZN(n1100) );
NAND2_X1 U1092 ( .A1(n1376), .A2(n1301), .ZN(n1116) );
INV_X1 U1093 ( .A(G902), .ZN(n1301) );
XOR2_X1 U1094 ( .A(n1377), .B(n1378), .Z(n1376) );
XNOR2_X1 U1095 ( .A(n1209), .B(n1200), .ZN(n1378) );
XOR2_X1 U1096 ( .A(G110), .B(n1379), .Z(n1200) );
NOR2_X1 U1097 ( .A1(G953), .A2(n1147), .ZN(n1379) );
INV_X1 U1098 ( .A(G227), .ZN(n1147) );
XOR2_X1 U1099 ( .A(n1356), .B(n1380), .Z(n1209) );
NOR2_X1 U1100 ( .A1(KEYINPUT38), .A2(n1342), .ZN(n1380) );
XNOR2_X1 U1101 ( .A(G104), .B(KEYINPUT55), .ZN(n1342) );
XOR2_X1 U1102 ( .A(n1065), .B(G101), .Z(n1356) );
INV_X1 U1103 ( .A(G107), .ZN(n1065) );
XOR2_X1 U1104 ( .A(n1381), .B(n1208), .Z(n1377) );
INV_X1 U1105 ( .A(n1142), .ZN(n1208) );
XOR2_X1 U1106 ( .A(n1382), .B(n1383), .Z(n1142) );
XOR2_X1 U1107 ( .A(G128), .B(n1384), .Z(n1383) );
NOR2_X1 U1108 ( .A1(KEYINPUT17), .A2(n1260), .ZN(n1384) );
INV_X1 U1109 ( .A(G146), .ZN(n1260) );
XOR2_X1 U1110 ( .A(n1262), .B(KEYINPUT34), .Z(n1382) );
INV_X1 U1111 ( .A(G143), .ZN(n1262) );
XNOR2_X1 U1112 ( .A(n1385), .B(n1386), .ZN(n1381) );
NAND2_X1 U1113 ( .A1(KEYINPUT18), .A2(n1189), .ZN(n1386) );
AND3_X1 U1114 ( .A1(n1387), .A2(n1388), .A3(n1389), .ZN(n1189) );
OR2_X1 U1115 ( .A1(n1140), .A2(KEYINPUT26), .ZN(n1389) );
NAND3_X1 U1116 ( .A1(KEYINPUT26), .A2(n1140), .A3(G131), .ZN(n1388) );
NAND2_X1 U1117 ( .A1(n1390), .A2(n1275), .ZN(n1387) );
INV_X1 U1118 ( .A(G131), .ZN(n1275) );
NAND2_X1 U1119 ( .A1(n1391), .A2(KEYINPUT26), .ZN(n1390) );
XNOR2_X1 U1120 ( .A(n1140), .B(KEYINPUT62), .ZN(n1391) );
XOR2_X1 U1121 ( .A(G134), .B(G137), .Z(n1140) );
NAND2_X1 U1122 ( .A1(KEYINPUT35), .A2(n1392), .ZN(n1385) );
INV_X1 U1123 ( .A(G140), .ZN(n1392) );
endmodule


