//Key = 1010011110010011000100110000011011101000011010000000001000001010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336;

XOR2_X1 U748 ( .A(n1021), .B(n1022), .Z(G9) );
NOR3_X1 U749 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
XNOR2_X1 U750 ( .A(n1026), .B(KEYINPUT28), .ZN(n1024) );
NAND2_X1 U751 ( .A1(KEYINPUT2), .A2(n1027), .ZN(n1021) );
NOR2_X1 U752 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR3_X1 U753 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NAND3_X1 U754 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1030) );
NAND2_X1 U755 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U756 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND4_X1 U757 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NAND2_X1 U758 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U759 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
XOR2_X1 U760 ( .A(n1048), .B(KEYINPUT59), .Z(n1046) );
XNOR2_X1 U761 ( .A(n1026), .B(KEYINPUT9), .ZN(n1044) );
NAND3_X1 U762 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1038) );
NAND2_X1 U763 ( .A1(n1052), .A2(n1053), .ZN(n1049) );
NAND3_X1 U764 ( .A1(n1042), .A2(n1054), .A3(n1041), .ZN(n1053) );
NAND2_X1 U765 ( .A1(n1040), .A2(n1055), .ZN(n1052) );
NAND2_X1 U766 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U767 ( .A1(n1042), .A2(n1058), .ZN(n1057) );
NAND2_X1 U768 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U769 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U770 ( .A1(n1041), .A2(n1063), .ZN(n1056) );
NAND2_X1 U771 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
INV_X1 U772 ( .A(n1066), .ZN(n1036) );
NOR3_X1 U773 ( .A1(n1067), .A2(G953), .A3(G952), .ZN(n1028) );
INV_X1 U774 ( .A(n1033), .ZN(n1067) );
NAND4_X1 U775 ( .A1(n1068), .A2(n1050), .A3(n1069), .A4(n1070), .ZN(n1033) );
NOR4_X1 U776 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1070) );
NOR2_X1 U777 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NAND3_X1 U778 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1071) );
XOR2_X1 U779 ( .A(n1080), .B(G472), .Z(n1079) );
NAND3_X1 U780 ( .A1(G475), .A2(n1076), .A3(n1075), .ZN(n1078) );
INV_X1 U781 ( .A(KEYINPUT55), .ZN(n1076) );
OR2_X1 U782 ( .A1(n1075), .A2(G475), .ZN(n1077) );
NOR3_X1 U783 ( .A1(n1061), .A2(n1081), .A3(n1082), .ZN(n1069) );
INV_X1 U784 ( .A(n1083), .ZN(n1082) );
XOR2_X1 U785 ( .A(n1084), .B(n1085), .Z(n1068) );
NOR2_X1 U786 ( .A1(n1086), .A2(KEYINPUT26), .ZN(n1085) );
NAND2_X1 U787 ( .A1(n1087), .A2(n1088), .ZN(G72) );
NAND3_X1 U788 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
NAND2_X1 U789 ( .A1(G953), .A2(n1092), .ZN(n1089) );
NAND2_X1 U790 ( .A1(G953), .A2(n1093), .ZN(n1087) );
NAND2_X1 U791 ( .A1(G900), .A2(n1094), .ZN(n1093) );
NAND2_X1 U792 ( .A1(n1095), .A2(n1092), .ZN(n1094) );
NAND2_X1 U793 ( .A1(n1091), .A2(n1090), .ZN(n1095) );
INV_X1 U794 ( .A(KEYINPUT13), .ZN(n1090) );
XNOR2_X1 U795 ( .A(n1096), .B(n1032), .ZN(n1091) );
NAND2_X1 U796 ( .A1(KEYINPUT0), .A2(n1097), .ZN(n1096) );
XNOR2_X1 U797 ( .A(n1098), .B(n1099), .ZN(n1097) );
XNOR2_X1 U798 ( .A(n1100), .B(n1101), .ZN(n1099) );
NOR2_X1 U799 ( .A1(KEYINPUT35), .A2(n1102), .ZN(n1101) );
XNOR2_X1 U800 ( .A(G131), .B(n1103), .ZN(n1102) );
NAND2_X1 U801 ( .A1(KEYINPUT41), .A2(n1104), .ZN(n1103) );
XOR2_X1 U802 ( .A(n1105), .B(n1106), .Z(G69) );
NAND2_X1 U803 ( .A1(G953), .A2(n1107), .ZN(n1106) );
NAND2_X1 U804 ( .A1(G898), .A2(G224), .ZN(n1107) );
NAND4_X1 U805 ( .A1(KEYINPUT33), .A2(n1108), .A3(n1109), .A4(n1110), .ZN(n1105) );
NAND3_X1 U806 ( .A1(n1111), .A2(n1034), .A3(n1031), .ZN(n1110) );
OR2_X1 U807 ( .A1(n1111), .A2(n1031), .ZN(n1109) );
NAND2_X1 U808 ( .A1(G953), .A2(n1112), .ZN(n1108) );
NAND2_X1 U809 ( .A1(G898), .A2(n1111), .ZN(n1112) );
XNOR2_X1 U810 ( .A(n1113), .B(n1114), .ZN(n1111) );
NAND3_X1 U811 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1113) );
OR2_X1 U812 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND3_X1 U813 ( .A1(n1119), .A2(n1118), .A3(KEYINPUT30), .ZN(n1116) );
NOR2_X1 U814 ( .A1(KEYINPUT63), .A2(n1120), .ZN(n1119) );
NAND2_X1 U815 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
INV_X1 U816 ( .A(KEYINPUT30), .ZN(n1121) );
NOR2_X1 U817 ( .A1(n1122), .A2(n1123), .ZN(G66) );
NOR3_X1 U818 ( .A1(n1084), .A2(n1124), .A3(n1125), .ZN(n1123) );
AND3_X1 U819 ( .A1(n1126), .A2(n1127), .A3(n1086), .ZN(n1125) );
INV_X1 U820 ( .A(n1128), .ZN(n1086) );
NOR2_X1 U821 ( .A1(n1129), .A2(n1126), .ZN(n1124) );
NOR2_X1 U822 ( .A1(n1130), .A2(n1128), .ZN(n1129) );
NOR2_X1 U823 ( .A1(n1031), .A2(n1032), .ZN(n1130) );
NOR2_X1 U824 ( .A1(n1122), .A2(n1131), .ZN(G63) );
XOR2_X1 U825 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U826 ( .A1(n1127), .A2(G478), .ZN(n1132) );
NOR2_X1 U827 ( .A1(n1122), .A2(n1134), .ZN(G60) );
XNOR2_X1 U828 ( .A(n1135), .B(n1136), .ZN(n1134) );
NOR3_X1 U829 ( .A1(n1137), .A2(KEYINPUT12), .A3(n1138), .ZN(n1136) );
INV_X1 U830 ( .A(G475), .ZN(n1138) );
XOR2_X1 U831 ( .A(G104), .B(n1139), .Z(G6) );
NOR2_X1 U832 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR2_X1 U833 ( .A1(n1122), .A2(n1142), .ZN(G57) );
XOR2_X1 U834 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U835 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND2_X1 U836 ( .A1(KEYINPUT5), .A2(n1147), .ZN(n1146) );
NAND2_X1 U837 ( .A1(n1127), .A2(G472), .ZN(n1145) );
XOR2_X1 U838 ( .A(n1148), .B(n1149), .Z(n1143) );
NAND2_X1 U839 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
XOR2_X1 U840 ( .A(n1152), .B(KEYINPUT58), .Z(n1150) );
OR2_X1 U841 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U842 ( .A1(n1155), .A2(n1156), .ZN(G54) );
XOR2_X1 U843 ( .A(KEYINPUT38), .B(n1157), .Z(n1156) );
NOR2_X1 U844 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XNOR2_X1 U845 ( .A(G953), .B(KEYINPUT50), .ZN(n1159) );
XOR2_X1 U846 ( .A(n1160), .B(n1161), .Z(n1155) );
XOR2_X1 U847 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U848 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U849 ( .A1(n1127), .A2(G469), .ZN(n1165) );
NAND2_X1 U850 ( .A1(KEYINPUT19), .A2(n1166), .ZN(n1164) );
XOR2_X1 U851 ( .A(n1167), .B(n1168), .Z(n1160) );
XNOR2_X1 U852 ( .A(n1169), .B(G110), .ZN(n1168) );
NOR2_X1 U853 ( .A1(KEYINPUT48), .A2(n1170), .ZN(n1167) );
XNOR2_X1 U854 ( .A(n1118), .B(n1171), .ZN(n1170) );
NOR2_X1 U855 ( .A1(n1122), .A2(n1172), .ZN(G51) );
XOR2_X1 U856 ( .A(n1173), .B(n1174), .Z(n1172) );
XNOR2_X1 U857 ( .A(G125), .B(n1175), .ZN(n1174) );
XNOR2_X1 U858 ( .A(KEYINPUT20), .B(KEYINPUT18), .ZN(n1175) );
XOR2_X1 U859 ( .A(n1176), .B(n1177), .Z(n1173) );
XOR2_X1 U860 ( .A(n1178), .B(n1179), .Z(n1176) );
NAND2_X1 U861 ( .A1(n1127), .A2(n1180), .ZN(n1178) );
INV_X1 U862 ( .A(n1137), .ZN(n1127) );
NAND2_X1 U863 ( .A1(G902), .A2(n1181), .ZN(n1137) );
OR2_X1 U864 ( .A1(n1032), .A2(n1031), .ZN(n1181) );
NAND4_X1 U865 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1031) );
NOR2_X1 U866 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NOR2_X1 U867 ( .A1(KEYINPUT45), .A2(n1188), .ZN(n1187) );
NOR2_X1 U868 ( .A1(n1189), .A2(n1140), .ZN(n1186) );
NOR3_X1 U869 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1189) );
NOR2_X1 U870 ( .A1(n1025), .A2(n1023), .ZN(n1192) );
NOR3_X1 U871 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1191) );
NOR2_X1 U872 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
AND2_X1 U873 ( .A1(n1041), .A2(n1198), .ZN(n1197) );
AND3_X1 U874 ( .A1(KEYINPUT45), .A2(n1059), .A3(n1199), .ZN(n1196) );
XOR2_X1 U875 ( .A(n1141), .B(KEYINPUT34), .Z(n1190) );
OR2_X1 U876 ( .A1(n1200), .A2(n1025), .ZN(n1141) );
NAND3_X1 U877 ( .A1(n1042), .A2(n1201), .A3(n1202), .ZN(n1025) );
NAND2_X1 U878 ( .A1(n1203), .A2(n1054), .ZN(n1184) );
NAND2_X1 U879 ( .A1(n1200), .A2(n1023), .ZN(n1054) );
NAND4_X1 U880 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1032) );
NOR4_X1 U881 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1207) );
NOR3_X1 U882 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1206) );
NOR2_X1 U883 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
INV_X1 U884 ( .A(KEYINPUT7), .ZN(n1215) );
NOR4_X1 U885 ( .A1(KEYINPUT7), .A2(n1217), .A3(n1198), .A4(n1023), .ZN(n1213) );
NOR3_X1 U886 ( .A1(n1218), .A2(n1219), .A3(n1193), .ZN(n1212) );
XNOR2_X1 U887 ( .A(KEYINPUT22), .B(n1220), .ZN(n1218) );
NOR2_X1 U888 ( .A1(n1034), .A2(n1158), .ZN(n1122) );
XNOR2_X1 U889 ( .A(G952), .B(KEYINPUT23), .ZN(n1158) );
XNOR2_X1 U890 ( .A(G146), .B(n1204), .ZN(G48) );
NAND3_X1 U891 ( .A1(n1221), .A2(n1222), .A3(n1198), .ZN(n1204) );
XOR2_X1 U892 ( .A(n1205), .B(n1223), .Z(G45) );
XNOR2_X1 U893 ( .A(G143), .B(KEYINPUT49), .ZN(n1223) );
NAND4_X1 U894 ( .A1(n1221), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1205) );
XNOR2_X1 U895 ( .A(n1169), .B(n1211), .ZN(G42) );
NOR3_X1 U896 ( .A1(n1200), .A2(n1064), .A3(n1219), .ZN(n1211) );
XOR2_X1 U897 ( .A(G137), .B(n1227), .Z(G39) );
NOR3_X1 U898 ( .A1(n1193), .A2(n1219), .A3(n1220), .ZN(n1227) );
NAND2_X1 U899 ( .A1(n1228), .A2(n1229), .ZN(G36) );
NAND2_X1 U900 ( .A1(n1210), .A2(n1230), .ZN(n1229) );
XOR2_X1 U901 ( .A(n1231), .B(KEYINPUT52), .Z(n1228) );
OR2_X1 U902 ( .A1(n1230), .A2(n1210), .ZN(n1231) );
NOR3_X1 U903 ( .A1(n1065), .A2(n1023), .A3(n1219), .ZN(n1210) );
INV_X1 U904 ( .A(G134), .ZN(n1230) );
XNOR2_X1 U905 ( .A(n1232), .B(n1209), .ZN(G33) );
NOR3_X1 U906 ( .A1(n1065), .A2(n1200), .A3(n1219), .ZN(n1209) );
NAND4_X1 U907 ( .A1(n1051), .A2(n1202), .A3(n1233), .A4(n1050), .ZN(n1219) );
XOR2_X1 U908 ( .A(n1048), .B(KEYINPUT4), .Z(n1051) );
XNOR2_X1 U909 ( .A(n1072), .B(KEYINPUT46), .ZN(n1048) );
XNOR2_X1 U910 ( .A(G128), .B(n1216), .ZN(G30) );
NAND3_X1 U911 ( .A1(n1221), .A2(n1234), .A3(n1198), .ZN(n1216) );
INV_X1 U912 ( .A(n1220), .ZN(n1198) );
INV_X1 U913 ( .A(n1217), .ZN(n1221) );
NAND3_X1 U914 ( .A1(n1202), .A2(n1233), .A3(n1026), .ZN(n1217) );
XNOR2_X1 U915 ( .A(G101), .B(n1182), .ZN(G3) );
NAND2_X1 U916 ( .A1(n1235), .A2(n1224), .ZN(n1182) );
INV_X1 U917 ( .A(n1065), .ZN(n1224) );
XNOR2_X1 U918 ( .A(n1208), .B(n1236), .ZN(G27) );
NAND2_X1 U919 ( .A1(KEYINPUT14), .A2(G125), .ZN(n1236) );
AND4_X1 U920 ( .A1(n1026), .A2(n1233), .A3(n1041), .A4(n1237), .ZN(n1208) );
NOR2_X1 U921 ( .A1(n1064), .A2(n1200), .ZN(n1237) );
NAND2_X1 U922 ( .A1(n1066), .A2(n1238), .ZN(n1233) );
NAND4_X1 U923 ( .A1(G953), .A2(G902), .A3(n1239), .A4(n1240), .ZN(n1238) );
INV_X1 U924 ( .A(G900), .ZN(n1240) );
XNOR2_X1 U925 ( .A(G122), .B(n1183), .ZN(G24) );
NAND4_X1 U926 ( .A1(n1241), .A2(n1042), .A3(n1225), .A4(n1226), .ZN(n1183) );
AND2_X1 U927 ( .A1(n1242), .A2(n1243), .ZN(n1042) );
INV_X1 U928 ( .A(n1244), .ZN(n1241) );
XOR2_X1 U929 ( .A(G119), .B(n1245), .Z(G21) );
NOR4_X1 U930 ( .A1(KEYINPUT39), .A2(n1220), .A3(n1193), .A4(n1244), .ZN(n1245) );
NAND2_X1 U931 ( .A1(n1246), .A2(n1247), .ZN(n1220) );
XOR2_X1 U932 ( .A(G116), .B(n1248), .Z(G18) );
NOR3_X1 U933 ( .A1(n1249), .A2(KEYINPUT25), .A3(n1250), .ZN(n1248) );
INV_X1 U934 ( .A(n1203), .ZN(n1250) );
XNOR2_X1 U935 ( .A(KEYINPUT8), .B(n1023), .ZN(n1249) );
INV_X1 U936 ( .A(n1234), .ZN(n1023) );
NOR2_X1 U937 ( .A1(n1226), .A2(n1251), .ZN(n1234) );
XNOR2_X1 U938 ( .A(G113), .B(n1252), .ZN(G15) );
NAND2_X1 U939 ( .A1(n1203), .A2(n1222), .ZN(n1252) );
INV_X1 U940 ( .A(n1200), .ZN(n1222) );
NAND2_X1 U941 ( .A1(n1251), .A2(n1226), .ZN(n1200) );
INV_X1 U942 ( .A(n1225), .ZN(n1251) );
NOR2_X1 U943 ( .A1(n1244), .A2(n1065), .ZN(n1203) );
NAND2_X1 U944 ( .A1(n1246), .A2(n1243), .ZN(n1065) );
XNOR2_X1 U945 ( .A(n1247), .B(KEYINPUT57), .ZN(n1243) );
INV_X1 U946 ( .A(n1242), .ZN(n1246) );
NAND3_X1 U947 ( .A1(n1026), .A2(n1201), .A3(n1041), .ZN(n1244) );
NOR2_X1 U948 ( .A1(n1253), .A2(n1061), .ZN(n1041) );
XNOR2_X1 U949 ( .A(G110), .B(n1188), .ZN(G12) );
NAND2_X1 U950 ( .A1(n1235), .A2(n1199), .ZN(n1188) );
INV_X1 U951 ( .A(n1064), .ZN(n1199) );
NAND2_X1 U952 ( .A1(n1247), .A2(n1242), .ZN(n1064) );
XNOR2_X1 U953 ( .A(n1254), .B(G472), .ZN(n1242) );
NAND2_X1 U954 ( .A1(KEYINPUT11), .A2(n1080), .ZN(n1254) );
NAND2_X1 U955 ( .A1(n1255), .A2(n1256), .ZN(n1080) );
XOR2_X1 U956 ( .A(n1257), .B(n1149), .Z(n1256) );
XNOR2_X1 U957 ( .A(n1258), .B(KEYINPUT16), .ZN(n1149) );
XOR2_X1 U958 ( .A(n1259), .B(n1147), .Z(n1257) );
XOR2_X1 U959 ( .A(n1162), .B(n1179), .Z(n1147) );
NAND3_X1 U960 ( .A1(n1260), .A2(n1261), .A3(KEYINPUT44), .ZN(n1259) );
NAND2_X1 U961 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XNOR2_X1 U962 ( .A(n1153), .B(n1264), .ZN(n1262) );
NOR2_X1 U963 ( .A1(KEYINPUT3), .A2(n1154), .ZN(n1264) );
OR2_X1 U964 ( .A1(n1151), .A2(n1263), .ZN(n1260) );
INV_X1 U965 ( .A(KEYINPUT37), .ZN(n1263) );
NAND2_X1 U966 ( .A1(n1154), .A2(n1153), .ZN(n1151) );
NAND2_X1 U967 ( .A1(G210), .A2(n1265), .ZN(n1153) );
INV_X1 U968 ( .A(G101), .ZN(n1154) );
XNOR2_X1 U969 ( .A(G902), .B(KEYINPUT61), .ZN(n1255) );
XOR2_X1 U970 ( .A(n1266), .B(n1084), .Z(n1247) );
NOR2_X1 U971 ( .A1(n1126), .A2(G902), .ZN(n1084) );
XNOR2_X1 U972 ( .A(n1267), .B(n1268), .ZN(n1126) );
XOR2_X1 U973 ( .A(n1269), .B(n1270), .Z(n1268) );
XOR2_X1 U974 ( .A(G128), .B(G119), .Z(n1270) );
XOR2_X1 U975 ( .A(G146), .B(G137), .Z(n1269) );
XOR2_X1 U976 ( .A(n1271), .B(n1272), .Z(n1267) );
NOR2_X1 U977 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XOR2_X1 U978 ( .A(n1275), .B(KEYINPUT15), .Z(n1274) );
NAND2_X1 U979 ( .A1(G125), .A2(n1169), .ZN(n1275) );
NOR2_X1 U980 ( .A1(G125), .A2(n1169), .ZN(n1273) );
INV_X1 U981 ( .A(G140), .ZN(n1169) );
XOR2_X1 U982 ( .A(n1276), .B(G110), .Z(n1271) );
NAND3_X1 U983 ( .A1(G221), .A2(n1277), .A3(KEYINPUT60), .ZN(n1276) );
NAND2_X1 U984 ( .A1(KEYINPUT36), .A2(n1128), .ZN(n1266) );
NAND2_X1 U985 ( .A1(G217), .A2(n1278), .ZN(n1128) );
NOR4_X1 U986 ( .A1(n1193), .A2(n1140), .A3(n1059), .A4(n1194), .ZN(n1235) );
INV_X1 U987 ( .A(n1201), .ZN(n1194) );
NAND2_X1 U988 ( .A1(n1066), .A2(n1279), .ZN(n1201) );
NAND4_X1 U989 ( .A1(G953), .A2(G902), .A3(n1239), .A4(n1280), .ZN(n1279) );
INV_X1 U990 ( .A(G898), .ZN(n1280) );
NAND3_X1 U991 ( .A1(n1239), .A2(n1034), .A3(G952), .ZN(n1066) );
NAND2_X1 U992 ( .A1(G237), .A2(G234), .ZN(n1239) );
INV_X1 U993 ( .A(n1202), .ZN(n1059) );
NOR2_X1 U994 ( .A1(n1061), .A2(n1062), .ZN(n1202) );
INV_X1 U995 ( .A(n1253), .ZN(n1062) );
NAND2_X1 U996 ( .A1(n1281), .A2(n1083), .ZN(n1253) );
NAND2_X1 U997 ( .A1(G469), .A2(n1282), .ZN(n1083) );
OR2_X1 U998 ( .A1(n1283), .A2(G902), .ZN(n1282) );
XNOR2_X1 U999 ( .A(n1081), .B(KEYINPUT17), .ZN(n1281) );
NOR3_X1 U1000 ( .A1(G469), .A2(G902), .A3(n1283), .ZN(n1081) );
XOR2_X1 U1001 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U1002 ( .A(n1162), .B(n1171), .ZN(n1285) );
INV_X1 U1003 ( .A(n1100), .ZN(n1171) );
XOR2_X1 U1004 ( .A(n1286), .B(n1287), .Z(n1100) );
XNOR2_X1 U1005 ( .A(G128), .B(KEYINPUT10), .ZN(n1286) );
XOR2_X1 U1006 ( .A(G131), .B(n1104), .Z(n1162) );
XOR2_X1 U1007 ( .A(G137), .B(G134), .Z(n1104) );
XOR2_X1 U1008 ( .A(n1288), .B(n1289), .Z(n1284) );
NOR2_X1 U1009 ( .A1(KEYINPUT27), .A2(n1118), .ZN(n1289) );
NAND2_X1 U1010 ( .A1(n1290), .A2(n1291), .ZN(n1288) );
NAND2_X1 U1011 ( .A1(n1166), .A2(n1292), .ZN(n1291) );
INV_X1 U1012 ( .A(n1293), .ZN(n1292) );
XOR2_X1 U1013 ( .A(n1294), .B(KEYINPUT40), .Z(n1290) );
NAND2_X1 U1014 ( .A1(n1295), .A2(n1293), .ZN(n1294) );
XOR2_X1 U1015 ( .A(G140), .B(n1296), .Z(n1293) );
NOR2_X1 U1016 ( .A1(KEYINPUT31), .A2(n1297), .ZN(n1296) );
XOR2_X1 U1017 ( .A(KEYINPUT29), .B(G110), .Z(n1297) );
XNOR2_X1 U1018 ( .A(n1166), .B(KEYINPUT24), .ZN(n1295) );
NOR2_X1 U1019 ( .A1(n1092), .A2(G953), .ZN(n1166) );
INV_X1 U1020 ( .A(G227), .ZN(n1092) );
AND2_X1 U1021 ( .A1(G221), .A2(n1278), .ZN(n1061) );
NAND2_X1 U1022 ( .A1(G234), .A2(n1298), .ZN(n1278) );
INV_X1 U1023 ( .A(n1026), .ZN(n1140) );
NOR2_X1 U1024 ( .A1(n1299), .A2(n1047), .ZN(n1026) );
INV_X1 U1025 ( .A(n1050), .ZN(n1047) );
NAND2_X1 U1026 ( .A1(G214), .A2(n1300), .ZN(n1050) );
INV_X1 U1027 ( .A(n1072), .ZN(n1299) );
XNOR2_X1 U1028 ( .A(n1301), .B(n1180), .ZN(n1072) );
AND2_X1 U1029 ( .A1(G210), .A2(n1300), .ZN(n1180) );
NAND2_X1 U1030 ( .A1(n1302), .A2(n1298), .ZN(n1300) );
INV_X1 U1031 ( .A(G237), .ZN(n1302) );
NAND3_X1 U1032 ( .A1(n1303), .A2(n1304), .A3(n1298), .ZN(n1301) );
NAND2_X1 U1033 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
INV_X1 U1034 ( .A(G125), .ZN(n1306) );
XNOR2_X1 U1035 ( .A(n1307), .B(KEYINPUT43), .ZN(n1305) );
NAND2_X1 U1036 ( .A1(n1308), .A2(G125), .ZN(n1303) );
XNOR2_X1 U1037 ( .A(KEYINPUT51), .B(n1309), .ZN(n1308) );
INV_X1 U1038 ( .A(n1307), .ZN(n1309) );
XOR2_X1 U1039 ( .A(n1179), .B(n1177), .Z(n1307) );
XNOR2_X1 U1040 ( .A(n1310), .B(n1114), .ZN(n1177) );
XOR2_X1 U1041 ( .A(G110), .B(G122), .Z(n1114) );
XOR2_X1 U1042 ( .A(n1311), .B(n1312), .Z(n1310) );
NOR2_X1 U1043 ( .A1(KEYINPUT56), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1044 ( .A(n1118), .B(n1120), .Z(n1313) );
XOR2_X1 U1045 ( .A(n1258), .B(KEYINPUT1), .Z(n1120) );
XOR2_X1 U1046 ( .A(n1314), .B(n1315), .Z(n1258) );
XNOR2_X1 U1047 ( .A(G113), .B(G119), .ZN(n1314) );
XOR2_X1 U1048 ( .A(G101), .B(n1316), .Z(n1118) );
XNOR2_X1 U1049 ( .A(n1027), .B(G104), .ZN(n1316) );
NAND2_X1 U1050 ( .A1(G224), .A2(n1034), .ZN(n1311) );
XOR2_X1 U1051 ( .A(n1317), .B(n1318), .Z(n1179) );
NOR2_X1 U1052 ( .A1(G128), .A2(KEYINPUT47), .ZN(n1318) );
INV_X1 U1053 ( .A(n1287), .ZN(n1317) );
INV_X1 U1054 ( .A(n1040), .ZN(n1193) );
NOR2_X1 U1055 ( .A1(n1225), .A2(n1226), .ZN(n1040) );
XNOR2_X1 U1056 ( .A(n1075), .B(G475), .ZN(n1226) );
NAND2_X1 U1057 ( .A1(n1135), .A2(n1298), .ZN(n1075) );
XNOR2_X1 U1058 ( .A(n1319), .B(n1320), .ZN(n1135) );
XOR2_X1 U1059 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1060 ( .A(G113), .B(G104), .Z(n1322) );
XNOR2_X1 U1061 ( .A(n1232), .B(G122), .ZN(n1321) );
INV_X1 U1062 ( .A(G131), .ZN(n1232) );
XOR2_X1 U1063 ( .A(n1323), .B(n1098), .Z(n1319) );
XOR2_X1 U1064 ( .A(G125), .B(G140), .Z(n1098) );
XNOR2_X1 U1065 ( .A(n1324), .B(n1287), .ZN(n1323) );
XNOR2_X1 U1066 ( .A(G143), .B(G146), .ZN(n1287) );
NAND2_X1 U1067 ( .A1(G214), .A2(n1265), .ZN(n1324) );
NOR2_X1 U1068 ( .A1(G953), .A2(G237), .ZN(n1265) );
XOR2_X1 U1069 ( .A(n1074), .B(KEYINPUT53), .Z(n1225) );
XNOR2_X1 U1070 ( .A(n1325), .B(G478), .ZN(n1074) );
NAND2_X1 U1071 ( .A1(n1133), .A2(n1298), .ZN(n1325) );
INV_X1 U1072 ( .A(G902), .ZN(n1298) );
XNOR2_X1 U1073 ( .A(n1326), .B(n1327), .ZN(n1133) );
XOR2_X1 U1074 ( .A(n1328), .B(n1329), .Z(n1327) );
NAND2_X1 U1075 ( .A1(G217), .A2(n1277), .ZN(n1329) );
AND2_X1 U1076 ( .A1(n1330), .A2(n1034), .ZN(n1277) );
INV_X1 U1077 ( .A(G953), .ZN(n1034) );
XNOR2_X1 U1078 ( .A(G234), .B(KEYINPUT62), .ZN(n1330) );
NAND2_X1 U1079 ( .A1(KEYINPUT32), .A2(n1331), .ZN(n1328) );
XOR2_X1 U1080 ( .A(n1332), .B(n1333), .Z(n1331) );
XNOR2_X1 U1081 ( .A(n1027), .B(n1315), .ZN(n1333) );
XOR2_X1 U1082 ( .A(G116), .B(KEYINPUT54), .Z(n1315) );
INV_X1 U1083 ( .A(G107), .ZN(n1027) );
XNOR2_X1 U1084 ( .A(G122), .B(n1334), .ZN(n1332) );
XNOR2_X1 U1085 ( .A(KEYINPUT6), .B(KEYINPUT42), .ZN(n1334) );
XOR2_X1 U1086 ( .A(n1335), .B(n1336), .Z(n1326) );
NOR2_X1 U1087 ( .A1(KEYINPUT21), .A2(G128), .ZN(n1336) );
XNOR2_X1 U1088 ( .A(G143), .B(G134), .ZN(n1335) );
endmodule


