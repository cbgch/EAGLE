//Key = 1011110100011011101000000101010010100100010001100000111100111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322;

NAND2_X1 U730 ( .A1(n1008), .A2(n1009), .ZN(G9) );
NAND2_X1 U731 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
XOR2_X1 U732 ( .A(n1012), .B(KEYINPUT44), .Z(n1008) );
NAND2_X1 U733 ( .A1(G107), .A2(n1013), .ZN(n1012) );
NOR2_X1 U734 ( .A1(n1014), .A2(n1015), .ZN(G75) );
NOR3_X1 U735 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1015) );
NAND3_X1 U736 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1016) );
NAND2_X1 U737 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U738 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND4_X1 U739 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n1025) );
NAND2_X1 U740 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NAND2_X1 U741 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U742 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U743 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
XNOR2_X1 U744 ( .A(KEYINPUT35), .B(n1038), .ZN(n1036) );
NAND3_X1 U745 ( .A1(n1039), .A2(n1040), .A3(n1032), .ZN(n1024) );
NAND2_X1 U746 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND3_X1 U747 ( .A1(n1043), .A2(n1029), .A3(n1027), .ZN(n1042) );
NAND2_X1 U748 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U749 ( .A1(n1046), .A2(n1047), .A3(n1026), .ZN(n1041) );
NAND2_X1 U750 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U751 ( .A1(n1030), .A2(n1027), .ZN(n1046) );
INV_X1 U752 ( .A(n1049), .ZN(n1027) );
AND3_X1 U753 ( .A1(n1050), .A2(n1029), .A3(n1051), .ZN(n1030) );
NAND2_X1 U754 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XNOR2_X1 U755 ( .A(KEYINPUT59), .B(n1039), .ZN(n1052) );
NAND2_X1 U756 ( .A1(n1054), .A2(n1055), .ZN(n1050) );
XOR2_X1 U757 ( .A(n1039), .B(KEYINPUT9), .Z(n1055) );
INV_X1 U758 ( .A(n1056), .ZN(n1022) );
NOR3_X1 U759 ( .A1(n1057), .A2(G953), .A3(G952), .ZN(n1014) );
INV_X1 U760 ( .A(n1019), .ZN(n1057) );
NAND2_X1 U761 ( .A1(n1058), .A2(n1059), .ZN(n1019) );
NOR4_X1 U762 ( .A1(n1037), .A2(n1048), .A3(n1060), .A4(n1061), .ZN(n1059) );
XNOR2_X1 U763 ( .A(n1062), .B(n1063), .ZN(n1061) );
NAND2_X1 U764 ( .A1(KEYINPUT52), .A2(n1064), .ZN(n1062) );
XOR2_X1 U765 ( .A(n1065), .B(n1066), .Z(n1060) );
NAND2_X1 U766 ( .A1(KEYINPUT16), .A2(n1067), .ZN(n1065) );
NOR4_X1 U767 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1058) );
XNOR2_X1 U768 ( .A(n1072), .B(n1073), .ZN(n1071) );
NOR2_X1 U769 ( .A1(KEYINPUT30), .A2(n1074), .ZN(n1073) );
XOR2_X1 U770 ( .A(n1075), .B(KEYINPUT0), .Z(n1068) );
XOR2_X1 U771 ( .A(n1076), .B(n1077), .Z(G72) );
XOR2_X1 U772 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U773 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U774 ( .A(n1082), .B(n1083), .Z(n1081) );
XOR2_X1 U775 ( .A(n1084), .B(n1085), .Z(n1083) );
XOR2_X1 U776 ( .A(G131), .B(n1086), .Z(n1085) );
NOR2_X1 U777 ( .A1(KEYINPUT49), .A2(n1087), .ZN(n1086) );
XOR2_X1 U778 ( .A(n1088), .B(n1089), .Z(n1082) );
AND2_X1 U779 ( .A1(n1090), .A2(n1091), .ZN(n1080) );
NAND2_X1 U780 ( .A1(n1020), .A2(n1017), .ZN(n1078) );
NAND2_X1 U781 ( .A1(G953), .A2(n1092), .ZN(n1076) );
NAND2_X1 U782 ( .A1(G900), .A2(G227), .ZN(n1092) );
NAND3_X1 U783 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(G69) );
XOR2_X1 U784 ( .A(n1096), .B(KEYINPUT43), .Z(n1095) );
NAND3_X1 U785 ( .A1(n1097), .A2(n1098), .A3(G953), .ZN(n1096) );
NAND2_X1 U786 ( .A1(G898), .A2(G224), .ZN(n1097) );
NAND2_X1 U787 ( .A1(n1099), .A2(n1020), .ZN(n1094) );
XOR2_X1 U788 ( .A(n1100), .B(n1018), .Z(n1099) );
NAND4_X1 U789 ( .A1(G898), .A2(G224), .A3(n1100), .A4(G953), .ZN(n1093) );
INV_X1 U790 ( .A(n1098), .ZN(n1100) );
NAND2_X1 U791 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
NAND2_X1 U792 ( .A1(n1103), .A2(n1091), .ZN(n1102) );
NOR2_X1 U793 ( .A1(n1104), .A2(n1105), .ZN(G66) );
XOR2_X1 U794 ( .A(n1106), .B(n1107), .Z(n1105) );
NAND2_X1 U795 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NOR2_X1 U796 ( .A1(n1104), .A2(n1110), .ZN(G63) );
XOR2_X1 U797 ( .A(n1111), .B(n1112), .Z(n1110) );
NAND2_X1 U798 ( .A1(n1108), .A2(G478), .ZN(n1111) );
NOR2_X1 U799 ( .A1(n1104), .A2(n1113), .ZN(G60) );
XOR2_X1 U800 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U801 ( .A1(n1108), .A2(G475), .ZN(n1114) );
XOR2_X1 U802 ( .A(G104), .B(n1116), .Z(G6) );
NOR2_X1 U803 ( .A1(n1104), .A2(n1117), .ZN(G57) );
XNOR2_X1 U804 ( .A(n1118), .B(n1119), .ZN(n1117) );
XOR2_X1 U805 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U806 ( .A1(n1108), .A2(G472), .ZN(n1120) );
NOR2_X1 U807 ( .A1(n1104), .A2(n1122), .ZN(G54) );
XOR2_X1 U808 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U809 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U810 ( .A(n1088), .B(n1127), .Z(n1126) );
XOR2_X1 U811 ( .A(n1128), .B(n1129), .Z(n1123) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND3_X1 U813 ( .A1(G469), .A2(n1108), .A3(KEYINPUT15), .ZN(n1131) );
INV_X1 U814 ( .A(n1132), .ZN(n1108) );
NAND2_X1 U815 ( .A1(KEYINPUT12), .A2(n1133), .ZN(n1128) );
XOR2_X1 U816 ( .A(G140), .B(G110), .Z(n1133) );
NOR2_X1 U817 ( .A1(n1104), .A2(n1134), .ZN(G51) );
XOR2_X1 U818 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR3_X1 U819 ( .A1(n1132), .A2(KEYINPUT62), .A3(n1074), .ZN(n1136) );
NAND2_X1 U820 ( .A1(G902), .A2(n1137), .ZN(n1132) );
OR2_X1 U821 ( .A1(n1018), .A2(n1017), .ZN(n1137) );
NAND4_X1 U822 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1017) );
AND4_X1 U823 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1141) );
NAND2_X1 U824 ( .A1(n1146), .A2(n1147), .ZN(n1140) );
NAND2_X1 U825 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND2_X1 U826 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND2_X1 U827 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U828 ( .A1(n1054), .A2(n1154), .ZN(n1153) );
INV_X1 U829 ( .A(KEYINPUT50), .ZN(n1154) );
NAND2_X1 U830 ( .A1(KEYINPUT50), .A2(n1155), .ZN(n1148) );
NAND4_X1 U831 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1018) );
NOR4_X1 U832 ( .A1(n1160), .A2(n1161), .A3(n1116), .A4(n1162), .ZN(n1159) );
NOR2_X1 U833 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
AND2_X1 U834 ( .A1(n1053), .A2(n1165), .ZN(n1116) );
NOR2_X1 U835 ( .A1(n1034), .A2(n1166), .ZN(n1161) );
XOR2_X1 U836 ( .A(KEYINPUT37), .B(n1167), .Z(n1166) );
NOR2_X1 U837 ( .A1(n1168), .A2(n1044), .ZN(n1167) );
NOR2_X1 U838 ( .A1(n1010), .A2(n1169), .ZN(n1158) );
INV_X1 U839 ( .A(n1013), .ZN(n1010) );
NAND2_X1 U840 ( .A1(n1054), .A2(n1165), .ZN(n1013) );
AND3_X1 U841 ( .A1(n1170), .A2(n1026), .A3(n1146), .ZN(n1165) );
NAND2_X1 U842 ( .A1(n1171), .A2(n1172), .ZN(n1135) );
NAND2_X1 U843 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NAND2_X1 U844 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
OR2_X1 U845 ( .A1(n1177), .A2(KEYINPUT10), .ZN(n1176) );
INV_X1 U846 ( .A(KEYINPUT40), .ZN(n1175) );
NAND2_X1 U847 ( .A1(n1177), .A2(n1178), .ZN(n1171) );
NAND2_X1 U848 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
OR2_X1 U849 ( .A1(n1173), .A2(KEYINPUT40), .ZN(n1180) );
XNOR2_X1 U850 ( .A(n1181), .B(n1182), .ZN(n1173) );
NOR2_X1 U851 ( .A1(KEYINPUT28), .A2(n1183), .ZN(n1182) );
XOR2_X1 U852 ( .A(G125), .B(n1184), .Z(n1181) );
INV_X1 U853 ( .A(KEYINPUT10), .ZN(n1179) );
NOR2_X1 U854 ( .A1(n1020), .A2(G952), .ZN(n1104) );
XOR2_X1 U855 ( .A(G146), .B(n1185), .Z(G48) );
NOR3_X1 U856 ( .A1(n1186), .A2(n1187), .A3(n1152), .ZN(n1185) );
XOR2_X1 U857 ( .A(n1034), .B(KEYINPUT51), .Z(n1187) );
XOR2_X1 U858 ( .A(n1188), .B(n1138), .Z(G45) );
NAND4_X1 U859 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1146), .ZN(n1138) );
NOR2_X1 U860 ( .A1(n1075), .A2(n1192), .ZN(n1191) );
XOR2_X1 U861 ( .A(n1193), .B(n1139), .Z(G42) );
NAND2_X1 U862 ( .A1(n1194), .A2(n1195), .ZN(n1139) );
XOR2_X1 U863 ( .A(n1087), .B(n1145), .Z(G39) );
NAND3_X1 U864 ( .A1(n1032), .A2(n1039), .A3(n1150), .ZN(n1145) );
INV_X1 U865 ( .A(G137), .ZN(n1087) );
XNOR2_X1 U866 ( .A(G134), .B(n1144), .ZN(G36) );
NAND3_X1 U867 ( .A1(n1196), .A2(n1039), .A3(n1189), .ZN(n1144) );
XNOR2_X1 U868 ( .A(G131), .B(n1143), .ZN(G33) );
NAND2_X1 U869 ( .A1(n1194), .A2(n1190), .ZN(n1143) );
AND3_X1 U870 ( .A1(n1053), .A2(n1039), .A3(n1189), .ZN(n1194) );
NAND2_X1 U871 ( .A1(n1197), .A2(n1198), .ZN(n1039) );
OR3_X1 U872 ( .A1(n1038), .A2(n1037), .A3(KEYINPUT35), .ZN(n1198) );
INV_X1 U873 ( .A(n1199), .ZN(n1037) );
NAND2_X1 U874 ( .A1(KEYINPUT35), .A2(n1146), .ZN(n1197) );
XNOR2_X1 U875 ( .A(G128), .B(n1200), .ZN(G30) );
NAND3_X1 U876 ( .A1(n1201), .A2(n1146), .A3(KEYINPUT53), .ZN(n1200) );
INV_X1 U877 ( .A(n1034), .ZN(n1146) );
INV_X1 U878 ( .A(n1155), .ZN(n1201) );
NAND2_X1 U879 ( .A1(n1150), .A2(n1054), .ZN(n1155) );
INV_X1 U880 ( .A(n1186), .ZN(n1150) );
NAND3_X1 U881 ( .A1(n1202), .A2(n1203), .A3(n1189), .ZN(n1186) );
AND3_X1 U882 ( .A1(n1204), .A2(n1029), .A3(n1049), .ZN(n1189) );
XOR2_X1 U883 ( .A(G101), .B(n1160), .Z(G3) );
NOR3_X1 U884 ( .A1(n1045), .A2(n1034), .A3(n1168), .ZN(n1160) );
XOR2_X1 U885 ( .A(n1142), .B(n1205), .Z(G27) );
NOR2_X1 U886 ( .A1(G125), .A2(KEYINPUT20), .ZN(n1205) );
NAND4_X1 U887 ( .A1(n1195), .A2(n1053), .A3(n1206), .A4(n1204), .ZN(n1142) );
NAND2_X1 U888 ( .A1(n1056), .A2(n1207), .ZN(n1204) );
NAND4_X1 U889 ( .A1(G902), .A2(n1091), .A3(n1208), .A4(n1090), .ZN(n1207) );
INV_X1 U890 ( .A(G900), .ZN(n1090) );
INV_X1 U891 ( .A(n1152), .ZN(n1053) );
XNOR2_X1 U892 ( .A(G122), .B(n1156), .ZN(G24) );
NAND4_X1 U893 ( .A1(n1209), .A2(n1026), .A3(n1210), .A4(n1211), .ZN(n1156) );
NOR2_X1 U894 ( .A1(n1203), .A2(n1202), .ZN(n1026) );
XNOR2_X1 U895 ( .A(G119), .B(n1157), .ZN(G21) );
NAND4_X1 U896 ( .A1(n1202), .A2(n1032), .A3(n1209), .A4(n1203), .ZN(n1157) );
INV_X1 U897 ( .A(n1163), .ZN(n1209) );
NAND2_X1 U898 ( .A1(n1212), .A2(n1213), .ZN(G18) );
NAND2_X1 U899 ( .A1(G116), .A2(n1214), .ZN(n1213) );
XOR2_X1 U900 ( .A(KEYINPUT3), .B(n1215), .Z(n1212) );
NOR2_X1 U901 ( .A1(G116), .A2(n1214), .ZN(n1215) );
NAND3_X1 U902 ( .A1(n1206), .A2(n1216), .A3(n1196), .ZN(n1214) );
INV_X1 U903 ( .A(n1164), .ZN(n1196) );
NAND2_X1 U904 ( .A1(n1190), .A2(n1054), .ZN(n1164) );
NOR2_X1 U905 ( .A1(n1211), .A2(n1192), .ZN(n1054) );
INV_X1 U906 ( .A(n1045), .ZN(n1190) );
XNOR2_X1 U907 ( .A(KEYINPUT55), .B(n1217), .ZN(n1216) );
XOR2_X1 U908 ( .A(G113), .B(n1169), .Z(G15) );
NOR3_X1 U909 ( .A1(n1152), .A2(n1045), .A3(n1163), .ZN(n1169) );
NAND2_X1 U910 ( .A1(n1206), .A2(n1217), .ZN(n1163) );
NOR3_X1 U911 ( .A1(n1049), .A2(n1048), .A3(n1034), .ZN(n1206) );
INV_X1 U912 ( .A(n1029), .ZN(n1048) );
NAND2_X1 U913 ( .A1(n1203), .A2(n1218), .ZN(n1045) );
NAND2_X1 U914 ( .A1(n1192), .A2(n1211), .ZN(n1152) );
INV_X1 U915 ( .A(n1210), .ZN(n1192) );
XOR2_X1 U916 ( .A(n1219), .B(n1220), .Z(G12) );
NAND3_X1 U917 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1220) );
XOR2_X1 U918 ( .A(n1044), .B(KEYINPUT2), .Z(n1223) );
INV_X1 U919 ( .A(n1195), .ZN(n1044) );
NOR2_X1 U920 ( .A1(n1218), .A2(n1203), .ZN(n1195) );
XOR2_X1 U921 ( .A(n1063), .B(n1064), .Z(n1203) );
INV_X1 U922 ( .A(G472), .ZN(n1064) );
NAND2_X1 U923 ( .A1(n1224), .A2(n1225), .ZN(n1063) );
XOR2_X1 U924 ( .A(n1121), .B(n1226), .Z(n1224) );
NOR2_X1 U925 ( .A1(KEYINPUT42), .A2(n1118), .ZN(n1226) );
XNOR2_X1 U926 ( .A(n1183), .B(n1227), .ZN(n1118) );
XOR2_X1 U927 ( .A(n1228), .B(n1229), .Z(n1121) );
XOR2_X1 U928 ( .A(G101), .B(n1230), .Z(n1229) );
XOR2_X1 U929 ( .A(KEYINPUT24), .B(G113), .Z(n1230) );
XOR2_X1 U930 ( .A(n1231), .B(n1232), .Z(n1228) );
NOR2_X1 U931 ( .A1(KEYINPUT8), .A2(n1233), .ZN(n1232) );
NAND2_X1 U932 ( .A1(G210), .A2(n1234), .ZN(n1231) );
INV_X1 U933 ( .A(n1202), .ZN(n1218) );
XNOR2_X1 U934 ( .A(n1070), .B(KEYINPUT46), .ZN(n1202) );
XNOR2_X1 U935 ( .A(n1235), .B(n1109), .ZN(n1070) );
AND2_X1 U936 ( .A1(G217), .A2(n1236), .ZN(n1109) );
NAND2_X1 U937 ( .A1(n1107), .A2(n1225), .ZN(n1235) );
XNOR2_X1 U938 ( .A(n1237), .B(n1238), .ZN(n1107) );
XOR2_X1 U939 ( .A(G110), .B(n1239), .Z(n1238) );
XOR2_X1 U940 ( .A(G128), .B(G119), .Z(n1239) );
XNOR2_X1 U941 ( .A(n1240), .B(n1241), .ZN(n1237) );
NOR2_X1 U942 ( .A1(KEYINPUT39), .A2(n1242), .ZN(n1241) );
XOR2_X1 U943 ( .A(n1243), .B(n1084), .Z(n1242) );
XOR2_X1 U944 ( .A(G125), .B(G140), .Z(n1084) );
XOR2_X1 U945 ( .A(n1244), .B(KEYINPUT57), .Z(n1243) );
NOR2_X1 U946 ( .A1(KEYINPUT19), .A2(n1245), .ZN(n1240) );
XOR2_X1 U947 ( .A(n1246), .B(G137), .Z(n1245) );
NAND2_X1 U948 ( .A1(G221), .A2(n1247), .ZN(n1246) );
INV_X1 U949 ( .A(n1168), .ZN(n1222) );
NAND2_X1 U950 ( .A1(n1032), .A2(n1170), .ZN(n1168) );
AND3_X1 U951 ( .A1(n1217), .A2(n1029), .A3(n1049), .ZN(n1170) );
XOR2_X1 U952 ( .A(n1248), .B(n1066), .Z(n1049) );
AND2_X1 U953 ( .A1(n1249), .A2(n1225), .ZN(n1066) );
XOR2_X1 U954 ( .A(n1250), .B(n1251), .Z(n1249) );
XOR2_X1 U955 ( .A(n1252), .B(n1253), .Z(n1251) );
NOR2_X1 U956 ( .A1(KEYINPUT21), .A2(n1254), .ZN(n1253) );
XOR2_X1 U957 ( .A(n1130), .B(n1255), .Z(n1254) );
NOR2_X1 U958 ( .A1(KEYINPUT1), .A2(n1256), .ZN(n1255) );
XOR2_X1 U959 ( .A(n1219), .B(G140), .Z(n1256) );
NAND2_X1 U960 ( .A1(G227), .A2(n1020), .ZN(n1130) );
NAND2_X1 U961 ( .A1(n1257), .A2(n1258), .ZN(n1252) );
OR2_X1 U962 ( .A1(n1259), .A2(n1088), .ZN(n1258) );
XOR2_X1 U963 ( .A(n1260), .B(KEYINPUT23), .Z(n1257) );
NAND2_X1 U964 ( .A1(n1088), .A2(n1259), .ZN(n1260) );
XNOR2_X1 U965 ( .A(n1127), .B(KEYINPUT58), .ZN(n1259) );
XOR2_X1 U966 ( .A(n1261), .B(n1262), .Z(n1127) );
XOR2_X1 U967 ( .A(G107), .B(n1263), .Z(n1262) );
NOR2_X1 U968 ( .A1(KEYINPUT47), .A2(n1264), .ZN(n1263) );
NAND2_X1 U969 ( .A1(KEYINPUT41), .A2(n1265), .ZN(n1261) );
INV_X1 U970 ( .A(G101), .ZN(n1265) );
XOR2_X1 U971 ( .A(n1266), .B(n1267), .Z(n1088) );
XOR2_X1 U972 ( .A(n1244), .B(n1268), .Z(n1267) );
NAND2_X1 U973 ( .A1(KEYINPUT11), .A2(n1269), .ZN(n1268) );
XOR2_X1 U974 ( .A(KEYINPUT22), .B(G128), .Z(n1269) );
INV_X1 U975 ( .A(G146), .ZN(n1244) );
NAND2_X1 U976 ( .A1(KEYINPUT29), .A2(n1188), .ZN(n1266) );
INV_X1 U977 ( .A(G143), .ZN(n1188) );
NAND2_X1 U978 ( .A1(KEYINPUT25), .A2(n1125), .ZN(n1250) );
XOR2_X1 U979 ( .A(n1227), .B(KEYINPUT5), .Z(n1125) );
XOR2_X1 U980 ( .A(n1089), .B(n1270), .Z(n1227) );
XOR2_X1 U981 ( .A(G137), .B(n1271), .Z(n1270) );
NOR2_X1 U982 ( .A1(G131), .A2(KEYINPUT13), .ZN(n1271) );
XOR2_X1 U983 ( .A(G134), .B(KEYINPUT36), .Z(n1089) );
NAND2_X1 U984 ( .A1(KEYINPUT34), .A2(n1067), .ZN(n1248) );
INV_X1 U985 ( .A(G469), .ZN(n1067) );
NAND2_X1 U986 ( .A1(G221), .A2(n1236), .ZN(n1029) );
NAND2_X1 U987 ( .A1(n1272), .A2(G234), .ZN(n1236) );
NAND2_X1 U988 ( .A1(n1056), .A2(n1273), .ZN(n1217) );
NAND4_X1 U989 ( .A1(n1103), .A2(G902), .A3(n1091), .A4(n1208), .ZN(n1273) );
XNOR2_X1 U990 ( .A(n1020), .B(KEYINPUT26), .ZN(n1091) );
XNOR2_X1 U991 ( .A(KEYINPUT48), .B(G898), .ZN(n1103) );
NAND3_X1 U992 ( .A1(n1208), .A2(n1020), .A3(G952), .ZN(n1056) );
NAND2_X1 U993 ( .A1(G237), .A2(G234), .ZN(n1208) );
NOR2_X1 U994 ( .A1(n1211), .A2(n1210), .ZN(n1032) );
XNOR2_X1 U995 ( .A(n1069), .B(KEYINPUT45), .ZN(n1210) );
XOR2_X1 U996 ( .A(G478), .B(n1274), .Z(n1069) );
AND2_X1 U997 ( .A1(n1225), .A2(n1112), .ZN(n1274) );
XNOR2_X1 U998 ( .A(n1275), .B(n1276), .ZN(n1112) );
XOR2_X1 U999 ( .A(n1277), .B(n1278), .Z(n1276) );
NAND2_X1 U1000 ( .A1(G217), .A2(n1247), .ZN(n1277) );
AND2_X1 U1001 ( .A1(G234), .A2(n1020), .ZN(n1247) );
XOR2_X1 U1002 ( .A(n1279), .B(n1280), .Z(n1275) );
NOR2_X1 U1003 ( .A1(KEYINPUT56), .A2(n1281), .ZN(n1280) );
XOR2_X1 U1004 ( .A(n1282), .B(n1283), .Z(n1281) );
XOR2_X1 U1005 ( .A(KEYINPUT54), .B(G134), .Z(n1283) );
XOR2_X1 U1006 ( .A(G116), .B(n1011), .Z(n1279) );
INV_X1 U1007 ( .A(n1075), .ZN(n1211) );
XOR2_X1 U1008 ( .A(n1284), .B(G475), .Z(n1075) );
NAND2_X1 U1009 ( .A1(n1115), .A2(n1225), .ZN(n1284) );
XNOR2_X1 U1010 ( .A(n1285), .B(n1286), .ZN(n1115) );
XOR2_X1 U1011 ( .A(G131), .B(n1287), .Z(n1286) );
XOR2_X1 U1012 ( .A(G146), .B(G143), .Z(n1287) );
XOR2_X1 U1013 ( .A(n1288), .B(n1289), .Z(n1285) );
XOR2_X1 U1014 ( .A(n1290), .B(n1291), .Z(n1289) );
NAND2_X1 U1015 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND2_X1 U1016 ( .A1(G125), .A2(n1193), .ZN(n1293) );
XOR2_X1 U1017 ( .A(KEYINPUT14), .B(n1294), .Z(n1292) );
NOR2_X1 U1018 ( .A1(G125), .A2(n1193), .ZN(n1294) );
INV_X1 U1019 ( .A(G140), .ZN(n1193) );
NAND2_X1 U1020 ( .A1(n1295), .A2(KEYINPUT61), .ZN(n1290) );
XOR2_X1 U1021 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U1022 ( .A(KEYINPUT38), .B(G104), .Z(n1297) );
XOR2_X1 U1023 ( .A(n1298), .B(n1299), .Z(n1296) );
INV_X1 U1024 ( .A(n1278), .ZN(n1299) );
NAND2_X1 U1025 ( .A1(KEYINPUT27), .A2(G113), .ZN(n1298) );
NAND2_X1 U1026 ( .A1(G214), .A2(n1234), .ZN(n1288) );
NOR2_X1 U1027 ( .A1(G953), .A2(G237), .ZN(n1234) );
XOR2_X1 U1028 ( .A(n1034), .B(KEYINPUT7), .Z(n1221) );
NAND2_X1 U1029 ( .A1(n1038), .A2(n1199), .ZN(n1034) );
NAND2_X1 U1030 ( .A1(G214), .A2(n1300), .ZN(n1199) );
XOR2_X1 U1031 ( .A(n1072), .B(n1074), .Z(n1038) );
NAND2_X1 U1032 ( .A1(G210), .A2(n1300), .ZN(n1074) );
NAND2_X1 U1033 ( .A1(n1272), .A2(n1301), .ZN(n1300) );
INV_X1 U1034 ( .A(G237), .ZN(n1301) );
XOR2_X1 U1035 ( .A(n1225), .B(KEYINPUT33), .Z(n1272) );
NAND2_X1 U1036 ( .A1(n1302), .A2(n1225), .ZN(n1072) );
INV_X1 U1037 ( .A(G902), .ZN(n1225) );
XOR2_X1 U1038 ( .A(n1303), .B(n1177), .Z(n1302) );
XOR2_X1 U1039 ( .A(n1101), .B(KEYINPUT4), .Z(n1177) );
XOR2_X1 U1040 ( .A(n1304), .B(n1305), .Z(n1101) );
XOR2_X1 U1041 ( .A(n1233), .B(n1278), .Z(n1305) );
XNOR2_X1 U1042 ( .A(G122), .B(KEYINPUT6), .ZN(n1278) );
XNOR2_X1 U1043 ( .A(G119), .B(G116), .ZN(n1233) );
XOR2_X1 U1044 ( .A(n1306), .B(n1307), .Z(n1304) );
XOR2_X1 U1045 ( .A(G113), .B(G110), .Z(n1307) );
NAND2_X1 U1046 ( .A1(n1308), .A2(n1309), .ZN(n1306) );
NAND2_X1 U1047 ( .A1(G101), .A2(n1310), .ZN(n1309) );
XOR2_X1 U1048 ( .A(KEYINPUT18), .B(n1311), .Z(n1308) );
NOR2_X1 U1049 ( .A1(G101), .A2(n1310), .ZN(n1311) );
NAND2_X1 U1050 ( .A1(n1312), .A2(n1313), .ZN(n1310) );
NAND2_X1 U1051 ( .A1(G107), .A2(n1264), .ZN(n1313) );
INV_X1 U1052 ( .A(G104), .ZN(n1264) );
XOR2_X1 U1053 ( .A(n1314), .B(KEYINPUT31), .Z(n1312) );
NAND2_X1 U1054 ( .A1(G104), .A2(n1011), .ZN(n1314) );
INV_X1 U1055 ( .A(G107), .ZN(n1011) );
NAND2_X1 U1056 ( .A1(n1315), .A2(n1316), .ZN(n1303) );
OR2_X1 U1057 ( .A1(n1184), .A2(n1317), .ZN(n1316) );
XOR2_X1 U1058 ( .A(n1318), .B(KEYINPUT17), .Z(n1315) );
NAND2_X1 U1059 ( .A1(n1317), .A2(n1184), .ZN(n1318) );
NAND2_X1 U1060 ( .A1(G224), .A2(n1020), .ZN(n1184) );
INV_X1 U1061 ( .A(G953), .ZN(n1020) );
XOR2_X1 U1062 ( .A(n1319), .B(n1183), .Z(n1317) );
XOR2_X1 U1063 ( .A(n1320), .B(n1282), .Z(n1183) );
XOR2_X1 U1064 ( .A(G128), .B(G143), .Z(n1282) );
NAND2_X1 U1065 ( .A1(KEYINPUT32), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1066 ( .A(KEYINPUT63), .B(G146), .Z(n1321) );
NAND2_X1 U1067 ( .A1(KEYINPUT60), .A2(n1322), .ZN(n1319) );
INV_X1 U1068 ( .A(G125), .ZN(n1322) );
INV_X1 U1069 ( .A(G110), .ZN(n1219) );
endmodule


