//Key = 1000101101101011110011110101100100001010000111110111000001100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351;

NAND2_X1 U737 ( .A1(n1027), .A2(n1028), .ZN(G9) );
NAND2_X1 U738 ( .A1(G107), .A2(n1029), .ZN(n1028) );
XOR2_X1 U739 ( .A(n1030), .B(KEYINPUT52), .Z(n1027) );
OR2_X1 U740 ( .A1(n1029), .A2(G107), .ZN(n1030) );
NOR2_X1 U741 ( .A1(n1031), .A2(n1032), .ZN(G75) );
NOR4_X1 U742 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1032) );
XOR2_X1 U743 ( .A(n1037), .B(KEYINPUT20), .Z(n1035) );
NAND3_X1 U744 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
XNOR2_X1 U745 ( .A(KEYINPUT56), .B(n1041), .ZN(n1039) );
NAND4_X1 U746 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1033) );
NAND3_X1 U747 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1043) );
INV_X1 U748 ( .A(n1049), .ZN(n1048) );
NAND2_X1 U749 ( .A1(n1050), .A2(n1051), .ZN(n1047) );
NAND3_X1 U750 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1051) );
NAND2_X1 U751 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NAND2_X1 U752 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U753 ( .A1(n1059), .A2(n1060), .ZN(n1050) );
NAND3_X1 U754 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NAND2_X1 U755 ( .A1(n1054), .A2(n1064), .ZN(n1063) );
NAND2_X1 U756 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U757 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U758 ( .A1(n1052), .A2(n1069), .ZN(n1062) );
NAND2_X1 U759 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
OR2_X1 U760 ( .A1(n1072), .A2(KEYINPUT5), .ZN(n1071) );
NAND3_X1 U761 ( .A1(KEYINPUT5), .A2(n1073), .A3(n1041), .ZN(n1061) );
XOR2_X1 U762 ( .A(KEYINPUT50), .B(n1074), .Z(n1042) );
AND3_X1 U763 ( .A1(n1040), .A2(n1075), .A3(n1052), .ZN(n1074) );
NOR3_X1 U764 ( .A1(n1076), .A2(n1077), .A3(n1049), .ZN(n1040) );
AND3_X1 U765 ( .A1(n1044), .A2(n1045), .A3(n1078), .ZN(n1031) );
NAND4_X1 U766 ( .A1(n1079), .A2(n1080), .A3(n1052), .A4(n1081), .ZN(n1044) );
NOR3_X1 U767 ( .A1(n1082), .A2(n1077), .A3(n1083), .ZN(n1081) );
XOR2_X1 U768 ( .A(n1084), .B(n1085), .Z(n1083) );
XOR2_X1 U769 ( .A(n1086), .B(KEYINPUT8), .Z(n1085) );
XOR2_X1 U770 ( .A(n1087), .B(n1088), .Z(n1082) );
XNOR2_X1 U771 ( .A(KEYINPUT4), .B(n1089), .ZN(n1088) );
NOR2_X1 U772 ( .A1(n1090), .A2(KEYINPUT2), .ZN(n1087) );
XOR2_X1 U773 ( .A(G472), .B(n1091), .Z(n1079) );
NOR2_X1 U774 ( .A1(n1092), .A2(KEYINPUT30), .ZN(n1091) );
XOR2_X1 U775 ( .A(n1093), .B(n1094), .Z(G72) );
NOR2_X1 U776 ( .A1(n1095), .A2(n1045), .ZN(n1094) );
NOR2_X1 U777 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U778 ( .A1(n1098), .A2(n1099), .ZN(n1093) );
NAND2_X1 U779 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XOR2_X1 U780 ( .A(KEYINPUT59), .B(n1102), .Z(n1100) );
AND2_X1 U781 ( .A1(n1036), .A2(n1045), .ZN(n1102) );
OR2_X1 U782 ( .A1(n1101), .A2(n1036), .ZN(n1098) );
NAND2_X1 U783 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NAND2_X1 U784 ( .A1(G953), .A2(n1097), .ZN(n1104) );
XOR2_X1 U785 ( .A(n1105), .B(n1106), .Z(n1103) );
XNOR2_X1 U786 ( .A(G125), .B(n1107), .ZN(n1106) );
XNOR2_X1 U787 ( .A(KEYINPUT23), .B(KEYINPUT18), .ZN(n1107) );
XOR2_X1 U788 ( .A(n1108), .B(n1109), .Z(n1105) );
XOR2_X1 U789 ( .A(n1110), .B(n1111), .Z(n1108) );
NAND2_X1 U790 ( .A1(KEYINPUT15), .A2(n1112), .ZN(n1110) );
XOR2_X1 U791 ( .A(n1113), .B(n1114), .Z(G69) );
NOR3_X1 U792 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
NOR2_X1 U793 ( .A1(G953), .A2(n1118), .ZN(n1117) );
XOR2_X1 U794 ( .A(n1034), .B(KEYINPUT0), .Z(n1118) );
NOR2_X1 U795 ( .A1(G224), .A2(n1045), .ZN(n1116) );
NAND2_X1 U796 ( .A1(n1119), .A2(n1120), .ZN(n1113) );
INV_X1 U797 ( .A(n1115), .ZN(n1120) );
NOR2_X1 U798 ( .A1(n1121), .A2(n1122), .ZN(G66) );
XOR2_X1 U799 ( .A(n1123), .B(n1124), .Z(n1122) );
OR2_X1 U800 ( .A1(n1125), .A2(n1089), .ZN(n1123) );
NOR2_X1 U801 ( .A1(n1121), .A2(n1126), .ZN(G63) );
NOR2_X1 U802 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U803 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U804 ( .A1(n1131), .A2(G478), .ZN(n1130) );
NAND2_X1 U805 ( .A1(KEYINPUT51), .A2(n1132), .ZN(n1129) );
NOR2_X1 U806 ( .A1(KEYINPUT51), .A2(n1132), .ZN(n1127) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1133), .ZN(G60) );
XOR2_X1 U808 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U809 ( .A1(n1131), .A2(G475), .ZN(n1134) );
XOR2_X1 U810 ( .A(n1136), .B(n1137), .Z(G6) );
XNOR2_X1 U811 ( .A(G104), .B(KEYINPUT29), .ZN(n1137) );
NOR3_X1 U812 ( .A1(n1121), .A2(n1138), .A3(n1139), .ZN(G57) );
NOR2_X1 U813 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR2_X1 U814 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NOR2_X1 U815 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NOR2_X1 U816 ( .A1(n1146), .A2(n1147), .ZN(n1142) );
NOR2_X1 U817 ( .A1(G101), .A2(n1148), .ZN(n1138) );
NOR2_X1 U818 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U819 ( .A1(n1147), .A2(n1145), .ZN(n1150) );
XNOR2_X1 U820 ( .A(n1146), .B(KEYINPUT35), .ZN(n1145) );
NOR2_X1 U821 ( .A1(n1144), .A2(n1146), .ZN(n1149) );
XNOR2_X1 U822 ( .A(n1151), .B(n1152), .ZN(n1146) );
NAND2_X1 U823 ( .A1(n1131), .A2(G472), .ZN(n1151) );
NOR3_X1 U824 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(G54) );
NOR3_X1 U825 ( .A1(n1156), .A2(n1045), .A3(n1078), .ZN(n1155) );
INV_X1 U826 ( .A(G952), .ZN(n1078) );
AND2_X1 U827 ( .A1(n1156), .A2(n1121), .ZN(n1154) );
INV_X1 U828 ( .A(KEYINPUT37), .ZN(n1156) );
XOR2_X1 U829 ( .A(n1157), .B(KEYINPUT25), .Z(n1153) );
XOR2_X1 U830 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U831 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U832 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U833 ( .A1(KEYINPUT6), .A2(n1164), .ZN(n1162) );
XNOR2_X1 U834 ( .A(KEYINPUT26), .B(KEYINPUT27), .ZN(n1160) );
XOR2_X1 U835 ( .A(n1165), .B(n1166), .Z(n1158) );
XNOR2_X1 U836 ( .A(n1167), .B(n1109), .ZN(n1166) );
XOR2_X1 U837 ( .A(n1168), .B(n1169), .Z(n1109) );
XOR2_X1 U838 ( .A(n1170), .B(n1171), .Z(n1165) );
NOR2_X1 U839 ( .A1(KEYINPUT1), .A2(n1172), .ZN(n1171) );
NAND2_X1 U840 ( .A1(n1131), .A2(G469), .ZN(n1170) );
INV_X1 U841 ( .A(n1125), .ZN(n1131) );
NOR3_X1 U842 ( .A1(n1173), .A2(n1121), .A3(n1174), .ZN(G51) );
NOR4_X1 U843 ( .A1(n1175), .A2(n1176), .A3(n1084), .A4(n1125), .ZN(n1174) );
NOR2_X1 U844 ( .A1(KEYINPUT63), .A2(n1177), .ZN(n1176) );
NOR2_X1 U845 ( .A1(n1178), .A2(n1179), .ZN(n1175) );
NOR2_X1 U846 ( .A1(KEYINPUT63), .A2(n1180), .ZN(n1178) );
NOR2_X1 U847 ( .A1(n1045), .A2(G952), .ZN(n1121) );
NOR2_X1 U848 ( .A1(n1181), .A2(n1182), .ZN(n1173) );
NOR2_X1 U849 ( .A1(n1179), .A2(n1180), .ZN(n1182) );
INV_X1 U850 ( .A(KEYINPUT7), .ZN(n1180) );
INV_X1 U851 ( .A(n1177), .ZN(n1179) );
XNOR2_X1 U852 ( .A(n1183), .B(n1184), .ZN(n1177) );
XOR2_X1 U853 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U854 ( .A1(KEYINPUT48), .A2(n1187), .ZN(n1185) );
NOR2_X1 U855 ( .A1(n1084), .A2(n1125), .ZN(n1181) );
NAND2_X1 U856 ( .A1(n1188), .A2(n1189), .ZN(n1125) );
OR2_X1 U857 ( .A1(n1034), .A2(n1036), .ZN(n1189) );
NAND2_X1 U858 ( .A1(n1190), .A2(n1191), .ZN(n1036) );
NOR4_X1 U859 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
NOR4_X1 U860 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1190) );
NOR2_X1 U861 ( .A1(n1076), .A2(n1200), .ZN(n1199) );
NOR4_X1 U862 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1198) );
XNOR2_X1 U863 ( .A(KEYINPUT16), .B(n1065), .ZN(n1204) );
INV_X1 U864 ( .A(n1205), .ZN(n1197) );
NAND4_X1 U865 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1034) );
AND3_X1 U866 ( .A1(n1136), .A2(n1029), .A3(n1210), .ZN(n1209) );
NAND3_X1 U867 ( .A1(n1046), .A2(n1073), .A3(n1211), .ZN(n1029) );
NAND3_X1 U868 ( .A1(n1211), .A2(n1046), .A3(n1212), .ZN(n1136) );
NAND2_X1 U869 ( .A1(n1054), .A2(n1213), .ZN(n1208) );
NAND2_X1 U870 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND3_X1 U871 ( .A1(KEYINPUT3), .A2(n1038), .A3(n1216), .ZN(n1215) );
NOR3_X1 U872 ( .A1(n1217), .A2(n1065), .A3(n1055), .ZN(n1216) );
NAND2_X1 U873 ( .A1(n1211), .A2(n1218), .ZN(n1214) );
NAND2_X1 U874 ( .A1(n1202), .A2(n1219), .ZN(n1218) );
OR2_X1 U875 ( .A1(n1220), .A2(KEYINPUT3), .ZN(n1219) );
INV_X1 U876 ( .A(n1038), .ZN(n1220) );
INV_X1 U877 ( .A(n1075), .ZN(n1202) );
NAND2_X1 U878 ( .A1(n1221), .A2(n1222), .ZN(n1207) );
XNOR2_X1 U879 ( .A(n1223), .B(KEYINPUT61), .ZN(n1221) );
NAND2_X1 U880 ( .A1(n1224), .A2(n1225), .ZN(n1206) );
NAND2_X1 U881 ( .A1(n1226), .A2(n1070), .ZN(n1225) );
XNOR2_X1 U882 ( .A(n1073), .B(KEYINPUT11), .ZN(n1226) );
INV_X1 U883 ( .A(n1227), .ZN(n1224) );
XNOR2_X1 U884 ( .A(KEYINPUT60), .B(n1228), .ZN(n1188) );
XNOR2_X1 U885 ( .A(n1229), .B(n1194), .ZN(G48) );
AND3_X1 U886 ( .A1(n1230), .A2(n1212), .A3(n1231), .ZN(n1194) );
XOR2_X1 U887 ( .A(G143), .B(n1232), .Z(G45) );
NOR3_X1 U888 ( .A1(n1233), .A2(KEYINPUT32), .A3(n1203), .ZN(n1232) );
INV_X1 U889 ( .A(n1234), .ZN(n1203) );
XNOR2_X1 U890 ( .A(G140), .B(n1235), .ZN(G42) );
NAND2_X1 U891 ( .A1(n1236), .A2(n1059), .ZN(n1235) );
XOR2_X1 U892 ( .A(n1200), .B(KEYINPUT14), .Z(n1236) );
NAND3_X1 U893 ( .A1(n1038), .A2(n1212), .A3(n1230), .ZN(n1200) );
XOR2_X1 U894 ( .A(G137), .B(n1237), .Z(G39) );
NOR2_X1 U895 ( .A1(KEYINPUT55), .A2(n1205), .ZN(n1237) );
NAND3_X1 U896 ( .A1(n1230), .A2(n1238), .A3(n1059), .ZN(n1205) );
INV_X1 U897 ( .A(n1076), .ZN(n1059) );
XOR2_X1 U898 ( .A(G134), .B(n1196), .Z(G36) );
NOR3_X1 U899 ( .A1(n1233), .A2(n1072), .A3(n1076), .ZN(n1196) );
XNOR2_X1 U900 ( .A(n1112), .B(n1195), .ZN(G33) );
NOR3_X1 U901 ( .A1(n1233), .A2(n1070), .A3(n1076), .ZN(n1195) );
NAND2_X1 U902 ( .A1(n1058), .A2(n1080), .ZN(n1076) );
NAND2_X1 U903 ( .A1(n1230), .A2(n1075), .ZN(n1233) );
XOR2_X1 U904 ( .A(G128), .B(n1193), .Z(G30) );
AND3_X1 U905 ( .A1(n1230), .A2(n1073), .A3(n1231), .ZN(n1193) );
NOR3_X1 U906 ( .A1(n1055), .A2(n1239), .A3(n1240), .ZN(n1231) );
NOR2_X1 U907 ( .A1(n1065), .A2(n1201), .ZN(n1230) );
INV_X1 U908 ( .A(n1241), .ZN(n1065) );
NAND2_X1 U909 ( .A1(n1242), .A2(n1243), .ZN(G3) );
NAND2_X1 U910 ( .A1(G101), .A2(n1244), .ZN(n1243) );
XOR2_X1 U911 ( .A(KEYINPUT22), .B(n1245), .Z(n1242) );
NOR2_X1 U912 ( .A1(G101), .A2(n1244), .ZN(n1245) );
NAND4_X1 U913 ( .A1(n1075), .A2(n1217), .A3(n1241), .A4(n1246), .ZN(n1244) );
NOR2_X1 U914 ( .A1(n1077), .A2(n1247), .ZN(n1246) );
XNOR2_X1 U915 ( .A(KEYINPUT47), .B(n1055), .ZN(n1247) );
XNOR2_X1 U916 ( .A(n1192), .B(n1248), .ZN(G27) );
XNOR2_X1 U917 ( .A(KEYINPUT31), .B(n1187), .ZN(n1248) );
INV_X1 U918 ( .A(G125), .ZN(n1187) );
AND3_X1 U919 ( .A1(n1038), .A2(n1212), .A3(n1249), .ZN(n1192) );
NOR3_X1 U920 ( .A1(n1041), .A2(n1201), .A3(n1055), .ZN(n1249) );
AND2_X1 U921 ( .A1(n1049), .A2(n1250), .ZN(n1201) );
NAND4_X1 U922 ( .A1(G902), .A2(G953), .A3(n1251), .A4(n1097), .ZN(n1250) );
INV_X1 U923 ( .A(G900), .ZN(n1097) );
XNOR2_X1 U924 ( .A(G122), .B(n1210), .ZN(G24) );
NAND4_X1 U925 ( .A1(n1234), .A2(n1052), .A3(n1046), .A4(n1217), .ZN(n1210) );
NOR3_X1 U926 ( .A1(n1055), .A2(n1252), .A3(n1253), .ZN(n1234) );
INV_X1 U927 ( .A(n1222), .ZN(n1055) );
XNOR2_X1 U928 ( .A(G119), .B(n1254), .ZN(G21) );
NAND2_X1 U929 ( .A1(n1223), .A2(n1222), .ZN(n1254) );
AND3_X1 U930 ( .A1(n1052), .A2(n1217), .A3(n1238), .ZN(n1223) );
NOR3_X1 U931 ( .A1(n1077), .A2(n1239), .A3(n1240), .ZN(n1238) );
INV_X1 U932 ( .A(n1255), .ZN(n1239) );
INV_X1 U933 ( .A(n1054), .ZN(n1077) );
XOR2_X1 U934 ( .A(G116), .B(n1256), .Z(G18) );
NOR2_X1 U935 ( .A1(n1072), .A2(n1227), .ZN(n1256) );
INV_X1 U936 ( .A(n1073), .ZN(n1072) );
NOR2_X1 U937 ( .A1(n1257), .A2(n1252), .ZN(n1073) );
INV_X1 U938 ( .A(n1258), .ZN(n1252) );
XOR2_X1 U939 ( .A(G113), .B(n1259), .Z(G15) );
NOR2_X1 U940 ( .A1(n1070), .A2(n1227), .ZN(n1259) );
NAND4_X1 U941 ( .A1(n1052), .A2(n1222), .A3(n1075), .A4(n1217), .ZN(n1227) );
NAND2_X1 U942 ( .A1(n1260), .A2(n1261), .ZN(n1075) );
NAND2_X1 U943 ( .A1(n1046), .A2(n1262), .ZN(n1261) );
INV_X1 U944 ( .A(KEYINPUT49), .ZN(n1262) );
NOR2_X1 U945 ( .A1(n1255), .A2(n1263), .ZN(n1046) );
INV_X1 U946 ( .A(n1240), .ZN(n1263) );
NAND3_X1 U947 ( .A1(n1240), .A2(n1255), .A3(KEYINPUT49), .ZN(n1260) );
INV_X1 U948 ( .A(n1041), .ZN(n1052) );
NAND2_X1 U949 ( .A1(n1068), .A2(n1264), .ZN(n1041) );
INV_X1 U950 ( .A(n1212), .ZN(n1070) );
NOR2_X1 U951 ( .A1(n1253), .A2(n1258), .ZN(n1212) );
XNOR2_X1 U952 ( .A(G110), .B(n1265), .ZN(G12) );
NAND3_X1 U953 ( .A1(n1054), .A2(n1211), .A3(n1266), .ZN(n1265) );
XNOR2_X1 U954 ( .A(n1038), .B(KEYINPUT45), .ZN(n1266) );
NOR2_X1 U955 ( .A1(n1240), .A2(n1255), .ZN(n1038) );
XOR2_X1 U956 ( .A(n1092), .B(G472), .Z(n1255) );
AND3_X1 U957 ( .A1(n1267), .A2(n1268), .A3(n1228), .ZN(n1092) );
NAND2_X1 U958 ( .A1(n1269), .A2(n1144), .ZN(n1268) );
INV_X1 U959 ( .A(n1147), .ZN(n1144) );
NAND2_X1 U960 ( .A1(n1270), .A2(n1147), .ZN(n1267) );
NAND2_X1 U961 ( .A1(n1271), .A2(G210), .ZN(n1147) );
XNOR2_X1 U962 ( .A(n1269), .B(KEYINPUT41), .ZN(n1270) );
XNOR2_X1 U963 ( .A(n1152), .B(n1140), .ZN(n1269) );
INV_X1 U964 ( .A(G101), .ZN(n1140) );
XNOR2_X1 U965 ( .A(n1272), .B(n1273), .ZN(n1152) );
XOR2_X1 U966 ( .A(n1274), .B(n1164), .Z(n1273) );
NOR2_X1 U967 ( .A1(G113), .A2(KEYINPUT39), .ZN(n1274) );
XNOR2_X1 U968 ( .A(n1186), .B(n1275), .ZN(n1272) );
XNOR2_X1 U969 ( .A(n1276), .B(n1090), .ZN(n1240) );
AND2_X1 U970 ( .A1(n1124), .A2(n1228), .ZN(n1090) );
XOR2_X1 U971 ( .A(n1277), .B(n1278), .Z(n1124) );
XOR2_X1 U972 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U973 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR2_X1 U974 ( .A1(KEYINPUT19), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U975 ( .A(G125), .B(n1168), .ZN(n1283) );
XNOR2_X1 U976 ( .A(G140), .B(n1229), .ZN(n1168) );
NAND2_X1 U977 ( .A1(n1284), .A2(G221), .ZN(n1281) );
XOR2_X1 U978 ( .A(n1285), .B(n1286), .Z(n1277) );
XOR2_X1 U979 ( .A(KEYINPUT17), .B(G128), .Z(n1286) );
XNOR2_X1 U980 ( .A(G119), .B(G110), .ZN(n1285) );
NAND2_X1 U981 ( .A1(KEYINPUT57), .A2(n1089), .ZN(n1276) );
NAND2_X1 U982 ( .A1(G217), .A2(n1287), .ZN(n1089) );
AND3_X1 U983 ( .A1(n1241), .A2(n1217), .A3(n1222), .ZN(n1211) );
NOR2_X1 U984 ( .A1(n1058), .A2(n1057), .ZN(n1222) );
INV_X1 U985 ( .A(n1080), .ZN(n1057) );
NAND2_X1 U986 ( .A1(G214), .A2(n1288), .ZN(n1080) );
XNOR2_X1 U987 ( .A(n1086), .B(n1289), .ZN(n1058) );
NOR2_X1 U988 ( .A1(KEYINPUT34), .A2(n1290), .ZN(n1289) );
XNOR2_X1 U989 ( .A(KEYINPUT24), .B(n1084), .ZN(n1290) );
NAND2_X1 U990 ( .A1(G210), .A2(n1288), .ZN(n1084) );
NAND2_X1 U991 ( .A1(n1291), .A2(n1228), .ZN(n1288) );
XNOR2_X1 U992 ( .A(G237), .B(KEYINPUT53), .ZN(n1291) );
NAND2_X1 U993 ( .A1(n1292), .A2(n1228), .ZN(n1086) );
XOR2_X1 U994 ( .A(n1293), .B(n1183), .Z(n1292) );
XNOR2_X1 U995 ( .A(n1119), .B(n1294), .ZN(n1183) );
AND2_X1 U996 ( .A1(n1045), .A2(G224), .ZN(n1294) );
XNOR2_X1 U997 ( .A(n1295), .B(n1296), .ZN(n1119) );
XNOR2_X1 U998 ( .A(G110), .B(n1297), .ZN(n1296) );
XNOR2_X1 U999 ( .A(KEYINPUT54), .B(KEYINPUT44), .ZN(n1297) );
XNOR2_X1 U1000 ( .A(n1298), .B(n1299), .ZN(n1295) );
XOR2_X1 U1001 ( .A(n1300), .B(n1275), .Z(n1299) );
XOR2_X1 U1002 ( .A(G116), .B(G119), .Z(n1275) );
NAND2_X1 U1003 ( .A1(n1301), .A2(n1302), .ZN(n1293) );
NAND2_X1 U1004 ( .A1(G125), .A2(n1186), .ZN(n1302) );
XOR2_X1 U1005 ( .A(n1303), .B(KEYINPUT42), .Z(n1301) );
OR2_X1 U1006 ( .A1(n1186), .A2(G125), .ZN(n1303) );
XNOR2_X1 U1007 ( .A(n1304), .B(G128), .ZN(n1186) );
NAND3_X1 U1008 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1304) );
NAND2_X1 U1009 ( .A1(n1229), .A2(n1308), .ZN(n1307) );
OR3_X1 U1010 ( .A1(n1308), .A2(n1229), .A3(G143), .ZN(n1306) );
INV_X1 U1011 ( .A(KEYINPUT21), .ZN(n1308) );
NAND2_X1 U1012 ( .A1(G143), .A2(n1309), .ZN(n1305) );
NAND2_X1 U1013 ( .A1(n1310), .A2(KEYINPUT21), .ZN(n1309) );
XNOR2_X1 U1014 ( .A(G146), .B(KEYINPUT9), .ZN(n1310) );
NAND2_X1 U1015 ( .A1(n1049), .A2(n1311), .ZN(n1217) );
NAND3_X1 U1016 ( .A1(n1115), .A2(n1251), .A3(G902), .ZN(n1311) );
NOR2_X1 U1017 ( .A1(G898), .A2(n1045), .ZN(n1115) );
NAND3_X1 U1018 ( .A1(n1251), .A2(n1045), .A3(G952), .ZN(n1049) );
NAND2_X1 U1019 ( .A1(G234), .A2(G237), .ZN(n1251) );
NOR2_X1 U1020 ( .A1(n1068), .A2(n1067), .ZN(n1241) );
INV_X1 U1021 ( .A(n1264), .ZN(n1067) );
NAND2_X1 U1022 ( .A1(G221), .A2(n1287), .ZN(n1264) );
NAND2_X1 U1023 ( .A1(G234), .A2(n1228), .ZN(n1287) );
XOR2_X1 U1024 ( .A(n1312), .B(G469), .Z(n1068) );
NAND3_X1 U1025 ( .A1(n1313), .A2(n1314), .A3(n1228), .ZN(n1312) );
NAND2_X1 U1026 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
INV_X1 U1027 ( .A(n1317), .ZN(n1316) );
XOR2_X1 U1028 ( .A(KEYINPUT43), .B(n1318), .Z(n1315) );
NAND2_X1 U1029 ( .A1(n1317), .A2(n1319), .ZN(n1313) );
XNOR2_X1 U1030 ( .A(n1318), .B(KEYINPUT38), .ZN(n1319) );
XNOR2_X1 U1031 ( .A(n1320), .B(n1163), .ZN(n1318) );
NOR2_X1 U1032 ( .A1(n1096), .A2(G953), .ZN(n1163) );
INV_X1 U1033 ( .A(G227), .ZN(n1096) );
NAND2_X1 U1034 ( .A1(n1321), .A2(KEYINPUT10), .ZN(n1320) );
XNOR2_X1 U1035 ( .A(n1322), .B(n1172), .ZN(n1321) );
INV_X1 U1036 ( .A(G110), .ZN(n1172) );
NAND2_X1 U1037 ( .A1(KEYINPUT46), .A2(n1323), .ZN(n1322) );
XNOR2_X1 U1038 ( .A(KEYINPUT25), .B(n1324), .ZN(n1323) );
XOR2_X1 U1039 ( .A(n1325), .B(n1167), .Z(n1317) );
INV_X1 U1040 ( .A(n1298), .ZN(n1167) );
XOR2_X1 U1041 ( .A(G101), .B(n1326), .Z(n1298) );
XOR2_X1 U1042 ( .A(G107), .B(G104), .Z(n1326) );
XOR2_X1 U1043 ( .A(n1327), .B(n1164), .Z(n1325) );
XOR2_X1 U1044 ( .A(n1111), .B(G131), .Z(n1164) );
XNOR2_X1 U1045 ( .A(G134), .B(n1279), .ZN(n1111) );
XNOR2_X1 U1046 ( .A(G137), .B(KEYINPUT13), .ZN(n1279) );
NAND2_X1 U1047 ( .A1(KEYINPUT62), .A2(n1328), .ZN(n1327) );
XOR2_X1 U1048 ( .A(n1169), .B(n1329), .Z(n1328) );
XNOR2_X1 U1049 ( .A(KEYINPUT26), .B(n1229), .ZN(n1329) );
NOR2_X1 U1050 ( .A1(n1258), .A2(n1257), .ZN(n1054) );
INV_X1 U1051 ( .A(n1253), .ZN(n1257) );
XNOR2_X1 U1052 ( .A(n1330), .B(n1331), .ZN(n1253) );
XOR2_X1 U1053 ( .A(KEYINPUT12), .B(G475), .Z(n1331) );
NAND2_X1 U1054 ( .A1(n1332), .A2(n1135), .ZN(n1330) );
XNOR2_X1 U1055 ( .A(n1333), .B(n1334), .ZN(n1135) );
XNOR2_X1 U1056 ( .A(n1300), .B(n1335), .ZN(n1334) );
XOR2_X1 U1057 ( .A(n1336), .B(n1337), .Z(n1335) );
NOR2_X1 U1058 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
XOR2_X1 U1059 ( .A(n1340), .B(KEYINPUT36), .Z(n1339) );
NAND2_X1 U1060 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
NOR2_X1 U1061 ( .A1(n1342), .A2(n1341), .ZN(n1338) );
XNOR2_X1 U1062 ( .A(KEYINPUT40), .B(n1229), .ZN(n1341) );
INV_X1 U1063 ( .A(G146), .ZN(n1229) );
XNOR2_X1 U1064 ( .A(n1324), .B(G125), .ZN(n1342) );
INV_X1 U1065 ( .A(G140), .ZN(n1324) );
NAND2_X1 U1066 ( .A1(n1271), .A2(G214), .ZN(n1336) );
NOR2_X1 U1067 ( .A1(G953), .A2(G237), .ZN(n1271) );
XOR2_X1 U1068 ( .A(G113), .B(G122), .Z(n1300) );
XNOR2_X1 U1069 ( .A(G104), .B(n1343), .ZN(n1333) );
XNOR2_X1 U1070 ( .A(G143), .B(n1112), .ZN(n1343) );
INV_X1 U1071 ( .A(G131), .ZN(n1112) );
XNOR2_X1 U1072 ( .A(KEYINPUT28), .B(n1228), .ZN(n1332) );
XOR2_X1 U1073 ( .A(G478), .B(n1344), .Z(n1258) );
AND2_X1 U1074 ( .A1(n1228), .A2(n1132), .ZN(n1344) );
XNOR2_X1 U1075 ( .A(n1345), .B(n1346), .ZN(n1132) );
XOR2_X1 U1076 ( .A(G134), .B(n1347), .Z(n1346) );
NOR2_X1 U1077 ( .A1(KEYINPUT33), .A2(n1348), .ZN(n1347) );
XOR2_X1 U1078 ( .A(n1349), .B(n1350), .Z(n1348) );
XOR2_X1 U1079 ( .A(G116), .B(G107), .Z(n1350) );
XOR2_X1 U1080 ( .A(KEYINPUT58), .B(G122), .Z(n1349) );
XOR2_X1 U1081 ( .A(n1351), .B(n1169), .Z(n1345) );
XOR2_X1 U1082 ( .A(G128), .B(G143), .Z(n1169) );
NAND2_X1 U1083 ( .A1(G217), .A2(n1284), .ZN(n1351) );
AND2_X1 U1084 ( .A1(G234), .A2(n1045), .ZN(n1284) );
INV_X1 U1085 ( .A(G953), .ZN(n1045) );
INV_X1 U1086 ( .A(G902), .ZN(n1228) );
endmodule


