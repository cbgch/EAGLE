//Key = 0010010100100001011010000010010010010111010000000111110001110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341;

XNOR2_X1 U736 ( .A(G107), .B(n1017), .ZN(G9) );
NOR2_X1 U737 ( .A1(n1018), .A2(n1019), .ZN(G75) );
NOR3_X1 U738 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1019) );
NOR2_X1 U739 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR3_X1 U740 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1023) );
NOR2_X1 U741 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR2_X1 U742 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR3_X1 U743 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1026) );
NOR2_X1 U744 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
AND2_X1 U745 ( .A1(n1029), .A2(n1036), .ZN(n1035) );
INV_X1 U746 ( .A(KEYINPUT56), .ZN(n1029) );
NOR2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(n1034) );
NOR2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1025) );
NOR2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U750 ( .A1(n1043), .A2(n1031), .ZN(n1042) );
INV_X1 U751 ( .A(n1044), .ZN(n1031) );
NOR2_X1 U752 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U753 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
XNOR2_X1 U754 ( .A(n1049), .B(KEYINPUT23), .ZN(n1047) );
NOR3_X1 U755 ( .A1(n1033), .A2(n1050), .A3(n1051), .ZN(n1041) );
NOR2_X1 U756 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U757 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
INV_X1 U758 ( .A(n1056), .ZN(n1033) );
NAND3_X1 U759 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1020) );
NAND3_X1 U760 ( .A1(n1056), .A2(n1060), .A3(n1044), .ZN(n1059) );
NOR2_X1 U761 ( .A1(n1061), .A2(n1051), .ZN(n1044) );
INV_X1 U762 ( .A(n1062), .ZN(n1061) );
NAND2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1060) );
NAND3_X1 U764 ( .A1(n1024), .A2(n1038), .A3(n1065), .ZN(n1064) );
INV_X1 U765 ( .A(KEYINPUT20), .ZN(n1038) );
NAND2_X1 U766 ( .A1(n1066), .A2(n1067), .ZN(n1063) );
XOR2_X1 U767 ( .A(n1068), .B(n1069), .Z(n1066) );
AND2_X1 U768 ( .A1(KEYINPUT39), .A2(n1070), .ZN(n1069) );
NOR3_X1 U769 ( .A1(n1071), .A2(G953), .A3(G952), .ZN(n1018) );
INV_X1 U770 ( .A(n1057), .ZN(n1071) );
NAND4_X1 U771 ( .A1(n1072), .A2(n1067), .A3(n1073), .A4(n1074), .ZN(n1057) );
NOR4_X1 U772 ( .A1(n1070), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1074) );
XNOR2_X1 U773 ( .A(n1078), .B(n1079), .ZN(n1076) );
XNOR2_X1 U774 ( .A(KEYINPUT35), .B(n1080), .ZN(n1079) );
XNOR2_X1 U775 ( .A(n1081), .B(n1082), .ZN(n1073) );
XNOR2_X1 U776 ( .A(KEYINPUT55), .B(n1083), .ZN(n1082) );
XNOR2_X1 U777 ( .A(n1084), .B(n1085), .ZN(n1072) );
XOR2_X1 U778 ( .A(n1086), .B(n1087), .Z(G72) );
NOR2_X1 U779 ( .A1(n1088), .A2(n1058), .ZN(n1087) );
AND2_X1 U780 ( .A1(G227), .A2(G900), .ZN(n1088) );
NAND2_X1 U781 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NAND3_X1 U782 ( .A1(n1091), .A2(n1058), .A3(n1092), .ZN(n1090) );
XOR2_X1 U783 ( .A(n1093), .B(KEYINPUT62), .Z(n1089) );
NAND2_X1 U784 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U785 ( .A1(n1092), .A2(n1058), .ZN(n1095) );
NAND2_X1 U786 ( .A1(n1096), .A2(n1097), .ZN(n1092) );
INV_X1 U787 ( .A(n1091), .ZN(n1094) );
NAND4_X1 U788 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1091) );
OR3_X1 U789 ( .A1(n1102), .A2(KEYINPUT54), .A3(n1103), .ZN(n1101) );
NAND2_X1 U790 ( .A1(n1103), .A2(n1104), .ZN(n1100) );
NAND2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
INV_X1 U792 ( .A(KEYINPUT54), .ZN(n1106) );
XOR2_X1 U793 ( .A(KEYINPUT57), .B(n1102), .Z(n1105) );
XOR2_X1 U794 ( .A(n1107), .B(KEYINPUT41), .Z(n1103) );
NAND2_X1 U795 ( .A1(G953), .A2(n1108), .ZN(n1099) );
NAND2_X1 U796 ( .A1(KEYINPUT54), .A2(n1102), .ZN(n1098) );
XNOR2_X1 U797 ( .A(n1109), .B(n1110), .ZN(n1102) );
XOR2_X1 U798 ( .A(KEYINPUT3), .B(n1111), .Z(n1110) );
NOR2_X1 U799 ( .A1(KEYINPUT19), .A2(n1112), .ZN(n1111) );
XOR2_X1 U800 ( .A(KEYINPUT14), .B(G137), .Z(n1112) );
XOR2_X1 U801 ( .A(n1113), .B(n1114), .Z(G69) );
XOR2_X1 U802 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U803 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U804 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U805 ( .A(n1121), .B(n1122), .Z(n1119) );
NAND2_X1 U806 ( .A1(KEYINPUT61), .A2(n1123), .ZN(n1121) );
NOR2_X1 U807 ( .A1(G898), .A2(n1058), .ZN(n1117) );
NAND2_X1 U808 ( .A1(n1058), .A2(n1124), .ZN(n1115) );
NAND2_X1 U809 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XNOR2_X1 U810 ( .A(KEYINPUT50), .B(n1127), .ZN(n1126) );
NAND2_X1 U811 ( .A1(G953), .A2(n1128), .ZN(n1113) );
NAND2_X1 U812 ( .A1(G898), .A2(G224), .ZN(n1128) );
NOR2_X1 U813 ( .A1(n1129), .A2(n1130), .ZN(G66) );
XNOR2_X1 U814 ( .A(n1131), .B(n1132), .ZN(n1130) );
NOR2_X1 U815 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U816 ( .A1(n1135), .A2(n1136), .ZN(G63) );
XOR2_X1 U817 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U818 ( .A1(n1139), .A2(n1134), .ZN(n1137) );
NOR2_X1 U819 ( .A1(n1140), .A2(n1058), .ZN(n1135) );
XNOR2_X1 U820 ( .A(G952), .B(KEYINPUT53), .ZN(n1140) );
NOR2_X1 U821 ( .A1(n1129), .A2(n1141), .ZN(G60) );
XNOR2_X1 U822 ( .A(n1142), .B(n1143), .ZN(n1141) );
NOR2_X1 U823 ( .A1(n1144), .A2(n1134), .ZN(n1143) );
XNOR2_X1 U824 ( .A(G104), .B(n1127), .ZN(G6) );
NOR2_X1 U825 ( .A1(n1129), .A2(n1145), .ZN(G57) );
XOR2_X1 U826 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U827 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U828 ( .A1(KEYINPUT4), .A2(n1150), .ZN(n1149) );
NOR2_X1 U829 ( .A1(n1083), .A2(n1134), .ZN(n1148) );
INV_X1 U830 ( .A(G472), .ZN(n1083) );
XNOR2_X1 U831 ( .A(n1151), .B(n1152), .ZN(n1146) );
NOR2_X1 U832 ( .A1(n1129), .A2(n1153), .ZN(G54) );
XOR2_X1 U833 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U834 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR2_X1 U835 ( .A1(n1080), .A2(n1134), .ZN(n1156) );
XOR2_X1 U836 ( .A(n1158), .B(n1159), .Z(n1154) );
XOR2_X1 U837 ( .A(G137), .B(n1160), .Z(n1159) );
NOR2_X1 U838 ( .A1(KEYINPUT47), .A2(n1161), .ZN(n1160) );
XOR2_X1 U839 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U840 ( .A1(n1164), .A2(n1165), .ZN(n1158) );
NAND2_X1 U841 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XNOR2_X1 U842 ( .A(KEYINPUT7), .B(n1168), .ZN(n1167) );
XOR2_X1 U843 ( .A(KEYINPUT18), .B(n1169), .Z(n1164) );
NOR2_X1 U844 ( .A1(n1166), .A2(n1168), .ZN(n1169) );
XNOR2_X1 U845 ( .A(n1170), .B(n1171), .ZN(n1166) );
NOR2_X1 U846 ( .A1(G110), .A2(KEYINPUT44), .ZN(n1171) );
NOR2_X1 U847 ( .A1(n1129), .A2(n1172), .ZN(G51) );
XOR2_X1 U848 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U849 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U850 ( .A1(KEYINPUT24), .A2(n1177), .ZN(n1175) );
XOR2_X1 U851 ( .A(n1178), .B(n1179), .Z(n1173) );
NOR4_X1 U852 ( .A1(n1180), .A2(n1181), .A3(KEYINPUT34), .A4(n1085), .ZN(n1179) );
NOR2_X1 U853 ( .A1(KEYINPUT5), .A2(n1182), .ZN(n1181) );
AND2_X1 U854 ( .A1(n1183), .A2(n1022), .ZN(n1182) );
AND2_X1 U855 ( .A1(n1134), .A2(KEYINPUT5), .ZN(n1180) );
NAND2_X1 U856 ( .A1(G902), .A2(n1022), .ZN(n1134) );
NAND4_X1 U857 ( .A1(n1184), .A2(n1096), .A3(n1125), .A4(n1127), .ZN(n1022) );
NAND3_X1 U858 ( .A1(n1185), .A2(n1062), .A3(n1036), .ZN(n1127) );
AND4_X1 U859 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1125) );
AND4_X1 U860 ( .A1(n1017), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1189) );
NAND3_X1 U861 ( .A1(n1065), .A2(n1062), .A3(n1185), .ZN(n1017) );
AND4_X1 U862 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1096) );
NOR4_X1 U863 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1196) );
INV_X1 U864 ( .A(n1201), .ZN(n1200) );
INV_X1 U865 ( .A(n1202), .ZN(n1198) );
XOR2_X1 U866 ( .A(n1097), .B(KEYINPUT45), .Z(n1184) );
NOR2_X1 U867 ( .A1(n1058), .A2(G952), .ZN(n1129) );
XNOR2_X1 U868 ( .A(G146), .B(n1195), .ZN(G48) );
NAND4_X1 U869 ( .A1(n1055), .A2(n1203), .A3(n1036), .A4(n1046), .ZN(n1195) );
XNOR2_X1 U870 ( .A(G143), .B(n1193), .ZN(G45) );
NAND4_X1 U871 ( .A1(n1068), .A2(n1046), .A3(n1053), .A4(n1204), .ZN(n1193) );
NOR4_X1 U872 ( .A1(n1070), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1204) );
INV_X1 U873 ( .A(n1208), .ZN(n1070) );
XNOR2_X1 U874 ( .A(G140), .B(n1194), .ZN(G42) );
NAND4_X1 U875 ( .A1(n1209), .A2(n1036), .A3(n1210), .A4(n1077), .ZN(n1194) );
NAND2_X1 U876 ( .A1(n1211), .A2(n1212), .ZN(G39) );
OR2_X1 U877 ( .A1(n1201), .A2(G137), .ZN(n1212) );
XOR2_X1 U878 ( .A(n1213), .B(KEYINPUT48), .Z(n1211) );
NAND2_X1 U879 ( .A1(G137), .A2(n1201), .ZN(n1213) );
NAND3_X1 U880 ( .A1(n1055), .A2(n1209), .A3(n1214), .ZN(n1201) );
XNOR2_X1 U881 ( .A(G134), .B(n1215), .ZN(G36) );
NAND2_X1 U882 ( .A1(KEYINPUT2), .A2(n1199), .ZN(n1215) );
AND3_X1 U883 ( .A1(n1209), .A2(n1065), .A3(n1053), .ZN(n1199) );
XNOR2_X1 U884 ( .A(G131), .B(n1097), .ZN(G33) );
NAND3_X1 U885 ( .A1(n1209), .A2(n1036), .A3(n1053), .ZN(n1097) );
NOR3_X1 U886 ( .A1(n1216), .A2(n1205), .A3(n1024), .ZN(n1209) );
NAND2_X1 U887 ( .A1(n1217), .A2(n1208), .ZN(n1024) );
XOR2_X1 U888 ( .A(n1068), .B(KEYINPUT39), .Z(n1217) );
INV_X1 U889 ( .A(n1218), .ZN(n1205) );
XNOR2_X1 U890 ( .A(G128), .B(n1202), .ZN(G30) );
NAND4_X1 U891 ( .A1(n1055), .A2(n1203), .A3(n1065), .A4(n1219), .ZN(n1202) );
XNOR2_X1 U892 ( .A(KEYINPUT60), .B(n1216), .ZN(n1219) );
INV_X1 U893 ( .A(n1046), .ZN(n1216) );
INV_X1 U894 ( .A(n1220), .ZN(n1203) );
XNOR2_X1 U895 ( .A(G101), .B(n1186), .ZN(G3) );
NAND3_X1 U896 ( .A1(n1067), .A2(n1185), .A3(n1053), .ZN(n1186) );
XOR2_X1 U897 ( .A(G125), .B(n1197), .Z(G27) );
NOR3_X1 U898 ( .A1(n1030), .A2(n1055), .A3(n1220), .ZN(n1197) );
NAND4_X1 U899 ( .A1(n1068), .A2(n1077), .A3(n1218), .A4(n1208), .ZN(n1220) );
NAND2_X1 U900 ( .A1(n1221), .A2(n1222), .ZN(n1218) );
NAND4_X1 U901 ( .A1(G953), .A2(n1223), .A3(n1224), .A4(n1108), .ZN(n1222) );
INV_X1 U902 ( .A(G900), .ZN(n1108) );
XNOR2_X1 U903 ( .A(KEYINPUT8), .B(n1183), .ZN(n1223) );
XOR2_X1 U904 ( .A(n1051), .B(KEYINPUT40), .Z(n1221) );
NAND2_X1 U905 ( .A1(n1056), .A2(n1036), .ZN(n1030) );
XNOR2_X1 U906 ( .A(G122), .B(n1187), .ZN(G24) );
NAND4_X1 U907 ( .A1(n1225), .A2(n1062), .A3(n1226), .A4(n1227), .ZN(n1187) );
NOR2_X1 U908 ( .A1(n1077), .A2(n1055), .ZN(n1062) );
XNOR2_X1 U909 ( .A(G119), .B(n1192), .ZN(G21) );
NAND3_X1 U910 ( .A1(n1055), .A2(n1214), .A3(n1225), .ZN(n1192) );
INV_X1 U911 ( .A(n1210), .ZN(n1055) );
XNOR2_X1 U912 ( .A(n1228), .B(n1229), .ZN(G18) );
NAND2_X1 U913 ( .A1(n1230), .A2(n1231), .ZN(n1228) );
NAND4_X1 U914 ( .A1(n1053), .A2(n1037), .A3(n1225), .A4(n1232), .ZN(n1231) );
INV_X1 U915 ( .A(n1065), .ZN(n1037) );
OR2_X1 U916 ( .A1(n1188), .A2(n1232), .ZN(n1230) );
INV_X1 U917 ( .A(KEYINPUT15), .ZN(n1232) );
NAND3_X1 U918 ( .A1(n1053), .A2(n1065), .A3(n1225), .ZN(n1188) );
NOR2_X1 U919 ( .A1(n1227), .A2(n1207), .ZN(n1065) );
INV_X1 U920 ( .A(n1226), .ZN(n1207) );
XNOR2_X1 U921 ( .A(G113), .B(n1191), .ZN(G15) );
NAND3_X1 U922 ( .A1(n1053), .A2(n1036), .A3(n1225), .ZN(n1191) );
AND2_X1 U923 ( .A1(n1056), .A2(n1233), .ZN(n1225) );
NOR2_X1 U924 ( .A1(n1234), .A2(n1075), .ZN(n1056) );
NOR2_X1 U925 ( .A1(n1226), .A2(n1206), .ZN(n1036) );
INV_X1 U926 ( .A(n1227), .ZN(n1206) );
NOR2_X1 U927 ( .A1(n1210), .A2(n1077), .ZN(n1053) );
XNOR2_X1 U928 ( .A(G110), .B(n1190), .ZN(G12) );
NAND3_X1 U929 ( .A1(n1185), .A2(n1210), .A3(n1214), .ZN(n1190) );
NOR2_X1 U930 ( .A1(n1040), .A2(n1054), .ZN(n1214) );
INV_X1 U931 ( .A(n1077), .ZN(n1054) );
XNOR2_X1 U932 ( .A(n1235), .B(n1236), .ZN(n1077) );
NOR2_X1 U933 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XOR2_X1 U934 ( .A(n1133), .B(KEYINPUT31), .Z(n1238) );
INV_X1 U935 ( .A(G217), .ZN(n1133) );
INV_X1 U936 ( .A(n1239), .ZN(n1237) );
NAND2_X1 U937 ( .A1(n1131), .A2(n1183), .ZN(n1235) );
XNOR2_X1 U938 ( .A(n1240), .B(n1241), .ZN(n1131) );
XOR2_X1 U939 ( .A(n1107), .B(n1242), .Z(n1241) );
XOR2_X1 U940 ( .A(n1243), .B(n1244), .Z(n1242) );
NOR2_X1 U941 ( .A1(G128), .A2(KEYINPUT30), .ZN(n1243) );
XNOR2_X1 U942 ( .A(G125), .B(n1245), .ZN(n1107) );
XOR2_X1 U943 ( .A(n1246), .B(n1247), .Z(n1240) );
XOR2_X1 U944 ( .A(KEYINPUT17), .B(G119), .Z(n1247) );
XOR2_X1 U945 ( .A(n1248), .B(G110), .Z(n1246) );
NAND2_X1 U946 ( .A1(n1249), .A2(G221), .ZN(n1248) );
INV_X1 U947 ( .A(n1067), .ZN(n1040) );
NOR2_X1 U948 ( .A1(n1226), .A2(n1227), .ZN(n1067) );
XOR2_X1 U949 ( .A(n1250), .B(n1144), .Z(n1227) );
INV_X1 U950 ( .A(G475), .ZN(n1144) );
NAND2_X1 U951 ( .A1(n1142), .A2(n1183), .ZN(n1250) );
XNOR2_X1 U952 ( .A(n1251), .B(n1252), .ZN(n1142) );
XOR2_X1 U953 ( .A(n1253), .B(n1254), .Z(n1252) );
XNOR2_X1 U954 ( .A(n1255), .B(n1256), .ZN(n1254) );
NOR2_X1 U955 ( .A1(KEYINPUT16), .A2(n1257), .ZN(n1256) );
XNOR2_X1 U956 ( .A(n1170), .B(n1258), .ZN(n1257) );
XNOR2_X1 U957 ( .A(n1259), .B(n1260), .ZN(n1258) );
NOR2_X1 U958 ( .A1(G146), .A2(KEYINPUT27), .ZN(n1260) );
NAND2_X1 U959 ( .A1(KEYINPUT52), .A2(G125), .ZN(n1259) );
NAND2_X1 U960 ( .A1(n1261), .A2(KEYINPUT51), .ZN(n1255) );
XNOR2_X1 U961 ( .A(n1262), .B(n1263), .ZN(n1261) );
NAND2_X1 U962 ( .A1(n1264), .A2(G214), .ZN(n1262) );
NOR2_X1 U963 ( .A1(G122), .A2(KEYINPUT11), .ZN(n1253) );
XOR2_X1 U964 ( .A(n1265), .B(n1266), .Z(n1251) );
XOR2_X1 U965 ( .A(G113), .B(G104), .Z(n1266) );
XNOR2_X1 U966 ( .A(G131), .B(KEYINPUT38), .ZN(n1265) );
XOR2_X1 U967 ( .A(n1267), .B(n1139), .Z(n1226) );
INV_X1 U968 ( .A(G478), .ZN(n1139) );
OR2_X1 U969 ( .A1(n1138), .A2(G902), .ZN(n1267) );
XNOR2_X1 U970 ( .A(n1268), .B(n1269), .ZN(n1138) );
XNOR2_X1 U971 ( .A(n1229), .B(n1270), .ZN(n1269) );
XOR2_X1 U972 ( .A(KEYINPUT59), .B(G122), .Z(n1270) );
XOR2_X1 U973 ( .A(n1271), .B(n1272), .Z(n1268) );
XNOR2_X1 U974 ( .A(G107), .B(n1273), .ZN(n1272) );
NAND2_X1 U975 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
NAND2_X1 U976 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XNOR2_X1 U977 ( .A(n1278), .B(n1279), .ZN(n1277) );
INV_X1 U978 ( .A(G128), .ZN(n1278) );
XNOR2_X1 U979 ( .A(KEYINPUT42), .B(n1280), .ZN(n1276) );
XOR2_X1 U980 ( .A(n1281), .B(KEYINPUT36), .Z(n1274) );
NAND2_X1 U981 ( .A1(n1282), .A2(n1280), .ZN(n1281) );
INV_X1 U982 ( .A(G134), .ZN(n1280) );
XNOR2_X1 U983 ( .A(G128), .B(n1279), .ZN(n1282) );
NOR2_X1 U984 ( .A1(KEYINPUT0), .A2(n1263), .ZN(n1279) );
INV_X1 U985 ( .A(G143), .ZN(n1263) );
NAND2_X1 U986 ( .A1(G217), .A2(n1249), .ZN(n1271) );
AND2_X1 U987 ( .A1(G234), .A2(n1058), .ZN(n1249) );
XOR2_X1 U988 ( .A(G472), .B(n1283), .Z(n1210) );
NOR2_X1 U989 ( .A1(n1081), .A2(KEYINPUT1), .ZN(n1283) );
AND2_X1 U990 ( .A1(n1284), .A2(n1183), .ZN(n1081) );
XOR2_X1 U991 ( .A(n1285), .B(n1286), .Z(n1284) );
XOR2_X1 U992 ( .A(n1152), .B(n1150), .Z(n1286) );
AND2_X1 U993 ( .A1(n1287), .A2(n1288), .ZN(n1150) );
NAND2_X1 U994 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
NAND2_X1 U995 ( .A1(n1264), .A2(G210), .ZN(n1289) );
NAND3_X1 U996 ( .A1(n1264), .A2(G210), .A3(G101), .ZN(n1287) );
NOR2_X1 U997 ( .A1(G953), .A2(G237), .ZN(n1264) );
XOR2_X1 U998 ( .A(G113), .B(n1291), .Z(n1152) );
XNOR2_X1 U999 ( .A(KEYINPUT32), .B(n1292), .ZN(n1285) );
NOR2_X1 U1000 ( .A1(KEYINPUT13), .A2(n1151), .ZN(n1292) );
XNOR2_X1 U1001 ( .A(n1293), .B(n1294), .ZN(n1151) );
XOR2_X1 U1002 ( .A(n1157), .B(n1244), .Z(n1294) );
XNOR2_X1 U1003 ( .A(G137), .B(n1295), .ZN(n1244) );
AND2_X1 U1004 ( .A1(n1233), .A2(n1296), .ZN(n1185) );
XOR2_X1 U1005 ( .A(KEYINPUT60), .B(n1046), .Z(n1296) );
NOR2_X1 U1006 ( .A1(n1049), .A2(n1075), .ZN(n1046) );
INV_X1 U1007 ( .A(n1048), .ZN(n1075) );
NAND2_X1 U1008 ( .A1(G221), .A2(n1239), .ZN(n1048) );
NAND2_X1 U1009 ( .A1(G234), .A2(n1183), .ZN(n1239) );
INV_X1 U1010 ( .A(n1234), .ZN(n1049) );
NAND2_X1 U1011 ( .A1(n1297), .A2(n1298), .ZN(n1234) );
NAND2_X1 U1012 ( .A1(n1078), .A2(n1080), .ZN(n1298) );
XOR2_X1 U1013 ( .A(KEYINPUT49), .B(n1299), .Z(n1297) );
NOR2_X1 U1014 ( .A1(n1078), .A2(n1080), .ZN(n1299) );
INV_X1 U1015 ( .A(G469), .ZN(n1080) );
AND2_X1 U1016 ( .A1(n1300), .A2(n1183), .ZN(n1078) );
XOR2_X1 U1017 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1018 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U1019 ( .A(G110), .B(n1168), .ZN(n1304) );
NAND2_X1 U1020 ( .A1(G227), .A2(n1058), .ZN(n1168) );
XOR2_X1 U1021 ( .A(KEYINPUT46), .B(G137), .Z(n1303) );
XOR2_X1 U1022 ( .A(n1109), .B(n1305), .Z(n1301) );
XNOR2_X1 U1023 ( .A(n1245), .B(n1163), .ZN(n1305) );
XNOR2_X1 U1024 ( .A(n1290), .B(n1306), .ZN(n1163) );
XNOR2_X1 U1025 ( .A(n1307), .B(G104), .ZN(n1306) );
INV_X1 U1026 ( .A(G101), .ZN(n1290) );
INV_X1 U1027 ( .A(n1170), .ZN(n1245) );
XOR2_X1 U1028 ( .A(G140), .B(KEYINPUT12), .Z(n1170) );
XOR2_X1 U1029 ( .A(n1162), .B(n1157), .Z(n1109) );
XOR2_X1 U1030 ( .A(G131), .B(G134), .Z(n1157) );
NAND3_X1 U1031 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1162) );
NAND2_X1 U1032 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
INV_X1 U1033 ( .A(KEYINPUT10), .ZN(n1312) );
NAND3_X1 U1034 ( .A1(KEYINPUT10), .A2(n1313), .A3(G128), .ZN(n1309) );
OR2_X1 U1035 ( .A1(n1313), .A2(G128), .ZN(n1308) );
NOR2_X1 U1036 ( .A1(KEYINPUT25), .A2(n1311), .ZN(n1313) );
NAND2_X1 U1037 ( .A1(n1314), .A2(n1315), .ZN(n1311) );
OR2_X1 U1038 ( .A1(n1316), .A2(n1295), .ZN(n1315) );
XOR2_X1 U1039 ( .A(n1317), .B(KEYINPUT28), .Z(n1314) );
NAND2_X1 U1040 ( .A1(n1316), .A2(n1295), .ZN(n1317) );
XOR2_X1 U1041 ( .A(n1318), .B(KEYINPUT37), .Z(n1316) );
AND3_X1 U1042 ( .A1(n1319), .A2(n1208), .A3(n1068), .ZN(n1233) );
XOR2_X1 U1043 ( .A(n1084), .B(n1320), .Z(n1068) );
NOR2_X1 U1044 ( .A1(n1321), .A2(KEYINPUT22), .ZN(n1320) );
INV_X1 U1045 ( .A(n1085), .ZN(n1321) );
NAND2_X1 U1046 ( .A1(G210), .A2(n1322), .ZN(n1085) );
NAND2_X1 U1047 ( .A1(n1323), .A2(n1183), .ZN(n1084) );
XOR2_X1 U1048 ( .A(n1324), .B(n1176), .Z(n1323) );
XNOR2_X1 U1049 ( .A(n1325), .B(n1122), .ZN(n1176) );
XNOR2_X1 U1050 ( .A(n1326), .B(G101), .ZN(n1122) );
NAND2_X1 U1051 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
NAND2_X1 U1052 ( .A1(G104), .A2(n1307), .ZN(n1328) );
XOR2_X1 U1053 ( .A(n1329), .B(KEYINPUT33), .Z(n1327) );
OR2_X1 U1054 ( .A1(n1307), .A2(G104), .ZN(n1329) );
INV_X1 U1055 ( .A(G107), .ZN(n1307) );
XNOR2_X1 U1056 ( .A(n1123), .B(n1330), .ZN(n1325) );
NOR2_X1 U1057 ( .A1(KEYINPUT9), .A2(n1331), .ZN(n1330) );
XOR2_X1 U1058 ( .A(KEYINPUT43), .B(n1120), .Z(n1331) );
XNOR2_X1 U1059 ( .A(n1332), .B(G113), .ZN(n1120) );
NAND3_X1 U1060 ( .A1(n1333), .A2(n1334), .A3(KEYINPUT29), .ZN(n1332) );
OR2_X1 U1061 ( .A1(n1291), .A2(KEYINPUT6), .ZN(n1334) );
XOR2_X1 U1062 ( .A(G116), .B(G119), .Z(n1291) );
NAND3_X1 U1063 ( .A1(G119), .A2(n1229), .A3(KEYINPUT6), .ZN(n1333) );
INV_X1 U1064 ( .A(G116), .ZN(n1229) );
XOR2_X1 U1065 ( .A(G110), .B(G122), .Z(n1123) );
NAND2_X1 U1066 ( .A1(n1335), .A2(KEYINPUT26), .ZN(n1324) );
XOR2_X1 U1067 ( .A(n1178), .B(n1336), .Z(n1335) );
NOR2_X1 U1068 ( .A1(KEYINPUT21), .A2(n1177), .ZN(n1336) );
XNOR2_X1 U1069 ( .A(n1293), .B(n1337), .ZN(n1177) );
XNOR2_X1 U1070 ( .A(n1295), .B(G125), .ZN(n1337) );
INV_X1 U1071 ( .A(G146), .ZN(n1295) );
XNOR2_X1 U1072 ( .A(G128), .B(n1318), .ZN(n1293) );
XOR2_X1 U1073 ( .A(G143), .B(KEYINPUT58), .Z(n1318) );
NAND2_X1 U1074 ( .A1(G224), .A2(n1058), .ZN(n1178) );
NAND2_X1 U1075 ( .A1(G214), .A2(n1322), .ZN(n1208) );
NAND2_X1 U1076 ( .A1(n1338), .A2(n1183), .ZN(n1322) );
INV_X1 U1077 ( .A(G902), .ZN(n1183) );
INV_X1 U1078 ( .A(G237), .ZN(n1338) );
NAND2_X1 U1079 ( .A1(n1339), .A2(n1340), .ZN(n1319) );
NAND4_X1 U1080 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1341), .ZN(n1340) );
INV_X1 U1081 ( .A(G898), .ZN(n1341) );
XNOR2_X1 U1082 ( .A(KEYINPUT63), .B(n1051), .ZN(n1339) );
NAND3_X1 U1083 ( .A1(n1224), .A2(n1058), .A3(G952), .ZN(n1051) );
INV_X1 U1084 ( .A(G953), .ZN(n1058) );
NAND2_X1 U1085 ( .A1(G237), .A2(G234), .ZN(n1224) );
endmodule


