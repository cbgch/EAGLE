//Key = 1001100100110000110100100011110001011101100001001000110000111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388;

NAND2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(G9) );
OR2_X1 U753 ( .A1(n1053), .A2(G107), .ZN(n1052) );
NAND2_X1 U754 ( .A1(G107), .A2(n1054), .ZN(n1051) );
NAND2_X1 U755 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
OR2_X1 U756 ( .A1(n1057), .A2(KEYINPUT63), .ZN(n1056) );
NAND2_X1 U757 ( .A1(KEYINPUT63), .A2(n1053), .ZN(n1055) );
OR2_X1 U758 ( .A1(KEYINPUT24), .A2(n1057), .ZN(n1053) );
NAND3_X1 U759 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
XOR2_X1 U760 ( .A(KEYINPUT23), .B(n1061), .Z(n1059) );
NAND4_X1 U761 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(G75) );
NAND2_X1 U762 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U763 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NAND4_X1 U764 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
NAND2_X1 U765 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND3_X1 U766 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NAND2_X1 U767 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NAND3_X1 U768 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1076) );
NAND2_X1 U769 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
NAND2_X1 U770 ( .A1(n1086), .A2(n1087), .ZN(n1074) );
INV_X1 U771 ( .A(n1088), .ZN(n1071) );
NAND4_X1 U772 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1068) );
NOR3_X1 U773 ( .A1(n1080), .A2(n1093), .A3(n1079), .ZN(n1092) );
XOR2_X1 U774 ( .A(n1094), .B(n1095), .Z(n1091) );
NAND2_X1 U775 ( .A1(n1096), .A2(n1097), .ZN(n1090) );
XNOR2_X1 U776 ( .A(KEYINPUT1), .B(n1098), .ZN(n1096) );
NAND2_X1 U777 ( .A1(n1099), .A2(G469), .ZN(n1089) );
XOR2_X1 U778 ( .A(n1098), .B(KEYINPUT5), .Z(n1099) );
NOR2_X1 U779 ( .A1(G953), .A2(n1100), .ZN(n1064) );
NOR3_X1 U780 ( .A1(n1101), .A2(n1080), .A3(n1088), .ZN(n1100) );
INV_X1 U781 ( .A(n1086), .ZN(n1080) );
NAND3_X1 U782 ( .A1(n1078), .A2(n1102), .A3(n1083), .ZN(n1101) );
NAND2_X1 U783 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND3_X1 U784 ( .A1(n1105), .A2(n1106), .A3(n1070), .ZN(n1103) );
NAND2_X1 U785 ( .A1(n1107), .A2(n1093), .ZN(n1106) );
NAND3_X1 U786 ( .A1(n1108), .A2(n1109), .A3(n1067), .ZN(n1105) );
XOR2_X1 U787 ( .A(n1110), .B(n1111), .Z(G72) );
XOR2_X1 U788 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND2_X1 U789 ( .A1(G953), .A2(n1114), .ZN(n1113) );
NAND2_X1 U790 ( .A1(G900), .A2(G227), .ZN(n1114) );
NAND3_X1 U791 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1112) );
NAND2_X1 U792 ( .A1(G953), .A2(n1118), .ZN(n1117) );
NAND2_X1 U793 ( .A1(n1119), .A2(n1120), .ZN(n1116) );
XOR2_X1 U794 ( .A(n1121), .B(n1122), .Z(n1119) );
XOR2_X1 U795 ( .A(KEYINPUT30), .B(KEYINPUT26), .Z(n1122) );
NAND2_X1 U796 ( .A1(n1121), .A2(n1123), .ZN(n1115) );
INV_X1 U797 ( .A(n1120), .ZN(n1123) );
XOR2_X1 U798 ( .A(n1124), .B(G131), .Z(n1120) );
NAND2_X1 U799 ( .A1(KEYINPUT19), .A2(n1125), .ZN(n1124) );
XOR2_X1 U800 ( .A(G134), .B(n1126), .Z(n1125) );
XOR2_X1 U801 ( .A(KEYINPUT34), .B(G137), .Z(n1126) );
XNOR2_X1 U802 ( .A(n1127), .B(n1128), .ZN(n1121) );
XOR2_X1 U803 ( .A(G140), .B(G125), .Z(n1128) );
NOR2_X1 U804 ( .A1(n1063), .A2(G953), .ZN(n1110) );
NAND2_X1 U805 ( .A1(n1129), .A2(n1130), .ZN(G69) );
NAND3_X1 U806 ( .A1(KEYINPUT59), .A2(n1131), .A3(n1132), .ZN(n1130) );
NAND2_X1 U807 ( .A1(n1133), .A2(n1134), .ZN(n1129) );
NAND2_X1 U808 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U809 ( .A1(n1131), .A2(n1137), .ZN(n1136) );
INV_X1 U810 ( .A(KEYINPUT53), .ZN(n1137) );
NAND2_X1 U811 ( .A1(KEYINPUT53), .A2(n1138), .ZN(n1135) );
NAND2_X1 U812 ( .A1(KEYINPUT59), .A2(n1131), .ZN(n1138) );
AND2_X1 U813 ( .A1(n1139), .A2(G953), .ZN(n1131) );
XOR2_X1 U814 ( .A(n1140), .B(KEYINPUT31), .Z(n1139) );
NAND2_X1 U815 ( .A1(G898), .A2(G224), .ZN(n1140) );
INV_X1 U816 ( .A(n1132), .ZN(n1133) );
XOR2_X1 U817 ( .A(n1141), .B(n1142), .Z(n1132) );
NOR2_X1 U818 ( .A1(n1062), .A2(G953), .ZN(n1142) );
NAND3_X1 U819 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1141) );
NAND2_X1 U820 ( .A1(G953), .A2(n1146), .ZN(n1145) );
NAND2_X1 U821 ( .A1(n1147), .A2(n1148), .ZN(n1144) );
XOR2_X1 U822 ( .A(n1149), .B(KEYINPUT43), .Z(n1148) );
NAND2_X1 U823 ( .A1(n1150), .A2(n1151), .ZN(n1143) );
NOR2_X1 U824 ( .A1(n1152), .A2(n1153), .ZN(G66) );
XOR2_X1 U825 ( .A(KEYINPUT49), .B(n1154), .Z(n1153) );
XOR2_X1 U826 ( .A(n1155), .B(n1156), .Z(n1152) );
NOR2_X1 U827 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND2_X1 U828 ( .A1(KEYINPUT16), .A2(n1159), .ZN(n1155) );
XOR2_X1 U829 ( .A(KEYINPUT7), .B(n1160), .Z(n1159) );
NOR2_X1 U830 ( .A1(n1154), .A2(n1161), .ZN(G63) );
XOR2_X1 U831 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U832 ( .A1(n1164), .A2(n1158), .ZN(n1162) );
INV_X1 U833 ( .A(G478), .ZN(n1164) );
NOR2_X1 U834 ( .A1(n1154), .A2(n1165), .ZN(G60) );
NOR2_X1 U835 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U836 ( .A(KEYINPUT2), .B(n1168), .Z(n1167) );
NOR3_X1 U837 ( .A1(n1169), .A2(n1170), .A3(n1158), .ZN(n1168) );
XOR2_X1 U838 ( .A(KEYINPUT58), .B(n1171), .Z(n1169) );
NOR2_X1 U839 ( .A1(n1172), .A2(n1171), .ZN(n1166) );
NOR2_X1 U840 ( .A1(n1170), .A2(n1158), .ZN(n1172) );
INV_X1 U841 ( .A(G475), .ZN(n1170) );
XOR2_X1 U842 ( .A(n1173), .B(G104), .Z(G6) );
NAND2_X1 U843 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NAND2_X1 U844 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
OR3_X1 U845 ( .A1(n1178), .A2(n1179), .A3(n1177), .ZN(n1174) );
INV_X1 U846 ( .A(KEYINPUT15), .ZN(n1177) );
NOR2_X1 U847 ( .A1(n1154), .A2(n1180), .ZN(G57) );
XOR2_X1 U848 ( .A(n1181), .B(n1182), .Z(n1180) );
XNOR2_X1 U849 ( .A(n1183), .B(n1184), .ZN(n1182) );
NAND2_X1 U850 ( .A1(n1185), .A2(KEYINPUT39), .ZN(n1183) );
XOR2_X1 U851 ( .A(n1186), .B(G101), .Z(n1185) );
XOR2_X1 U852 ( .A(n1187), .B(n1188), .Z(n1181) );
NOR2_X1 U853 ( .A1(n1095), .A2(n1158), .ZN(n1188) );
NOR2_X1 U854 ( .A1(KEYINPUT61), .A2(n1189), .ZN(n1187) );
XOR2_X1 U855 ( .A(n1190), .B(n1191), .Z(n1189) );
NOR2_X1 U856 ( .A1(n1154), .A2(n1192), .ZN(G54) );
XOR2_X1 U857 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U858 ( .A(n1195), .B(n1196), .Z(n1193) );
NOR2_X1 U859 ( .A1(n1097), .A2(n1158), .ZN(n1196) );
INV_X1 U860 ( .A(G469), .ZN(n1097) );
NAND2_X1 U861 ( .A1(KEYINPUT48), .A2(n1197), .ZN(n1195) );
NOR2_X1 U862 ( .A1(n1154), .A2(n1198), .ZN(G51) );
XOR2_X1 U863 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U864 ( .A1(n1201), .A2(n1158), .ZN(n1199) );
NAND2_X1 U865 ( .A1(G902), .A2(n1202), .ZN(n1158) );
NAND2_X1 U866 ( .A1(n1062), .A2(n1203), .ZN(n1202) );
XOR2_X1 U867 ( .A(KEYINPUT13), .B(n1063), .Z(n1203) );
AND4_X1 U868 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1063) );
NOR4_X1 U869 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1207) );
NOR2_X1 U870 ( .A1(n1212), .A2(n1213), .ZN(n1206) );
INV_X1 U871 ( .A(n1214), .ZN(n1213) );
NAND3_X1 U872 ( .A1(n1215), .A2(n1216), .A3(n1086), .ZN(n1204) );
XOR2_X1 U873 ( .A(KEYINPUT51), .B(n1217), .Z(n1216) );
AND4_X1 U874 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1062) );
AND4_X1 U875 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1221) );
OR2_X1 U876 ( .A1(n1109), .A2(n1178), .ZN(n1222) );
AND2_X1 U877 ( .A1(n1226), .A2(n1227), .ZN(n1220) );
INV_X1 U878 ( .A(n1176), .ZN(n1218) );
NOR2_X1 U879 ( .A1(n1108), .A2(n1178), .ZN(n1176) );
NAND2_X1 U880 ( .A1(n1058), .A2(n1061), .ZN(n1178) );
NOR4_X1 U881 ( .A1(n1079), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1058) );
INV_X1 U882 ( .A(G210), .ZN(n1201) );
NOR2_X1 U883 ( .A1(n1231), .A2(G952), .ZN(n1154) );
XOR2_X1 U884 ( .A(G146), .B(n1212), .Z(G48) );
AND3_X1 U885 ( .A1(n1179), .A2(n1061), .A3(n1232), .ZN(n1212) );
XOR2_X1 U886 ( .A(n1233), .B(n1205), .Z(G45) );
NAND4_X1 U887 ( .A1(n1234), .A2(n1061), .A3(n1235), .A4(n1236), .ZN(n1205) );
XOR2_X1 U888 ( .A(G140), .B(n1237), .Z(G42) );
NOR3_X1 U889 ( .A1(n1238), .A2(n1228), .A3(n1239), .ZN(n1237) );
XOR2_X1 U890 ( .A(KEYINPUT40), .B(n1086), .Z(n1238) );
XOR2_X1 U891 ( .A(G137), .B(n1211), .Z(G39) );
AND3_X1 U892 ( .A1(n1232), .A2(n1072), .A3(n1086), .ZN(n1211) );
XOR2_X1 U893 ( .A(G134), .B(n1210), .Z(G36) );
AND3_X1 U894 ( .A1(n1234), .A2(n1060), .A3(n1086), .ZN(n1210) );
XOR2_X1 U895 ( .A(n1240), .B(n1214), .Z(G33) );
NAND3_X1 U896 ( .A1(n1234), .A2(n1179), .A3(n1086), .ZN(n1214) );
NOR2_X1 U897 ( .A1(n1241), .A2(n1084), .ZN(n1086) );
AND3_X1 U898 ( .A1(n1217), .A2(n1242), .A3(n1087), .ZN(n1234) );
XOR2_X1 U899 ( .A(G128), .B(n1209), .Z(G30) );
AND3_X1 U900 ( .A1(n1060), .A2(n1061), .A3(n1232), .ZN(n1209) );
AND4_X1 U901 ( .A1(n1229), .A2(n1217), .A3(n1079), .A4(n1242), .ZN(n1232) );
XOR2_X1 U902 ( .A(n1243), .B(n1244), .Z(G3) );
NAND2_X1 U903 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND4_X1 U904 ( .A1(n1230), .A2(n1087), .A3(n1247), .A4(n1248), .ZN(n1246) );
NOR2_X1 U905 ( .A1(n1082), .A2(n1104), .ZN(n1247) );
OR2_X1 U906 ( .A1(n1219), .A2(n1248), .ZN(n1245) );
INV_X1 U907 ( .A(KEYINPUT29), .ZN(n1248) );
NAND2_X1 U908 ( .A1(n1087), .A2(n1249), .ZN(n1219) );
NAND2_X1 U909 ( .A1(KEYINPUT27), .A2(n1250), .ZN(n1243) );
XNOR2_X1 U910 ( .A(n1208), .B(n1251), .ZN(G27) );
NAND2_X1 U911 ( .A1(KEYINPUT3), .A2(G125), .ZN(n1251) );
AND2_X1 U912 ( .A1(n1215), .A2(n1252), .ZN(n1208) );
INV_X1 U913 ( .A(n1239), .ZN(n1215) );
NAND4_X1 U914 ( .A1(n1179), .A2(n1078), .A3(n1079), .A4(n1242), .ZN(n1239) );
NAND2_X1 U915 ( .A1(n1088), .A2(n1253), .ZN(n1242) );
NAND4_X1 U916 ( .A1(G953), .A2(G902), .A3(n1254), .A4(n1118), .ZN(n1253) );
INV_X1 U917 ( .A(G900), .ZN(n1118) );
XOR2_X1 U918 ( .A(n1255), .B(n1227), .Z(G24) );
NAND4_X1 U919 ( .A1(n1083), .A2(n1256), .A3(n1257), .A4(n1078), .ZN(n1227) );
NOR2_X1 U920 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XNOR2_X1 U921 ( .A(G119), .B(n1226), .ZN(G21) );
NAND4_X1 U922 ( .A1(n1229), .A2(n1256), .A3(n1072), .A4(n1079), .ZN(n1226) );
NAND2_X1 U923 ( .A1(n1260), .A2(n1261), .ZN(G18) );
OR2_X1 U924 ( .A1(n1225), .A2(G116), .ZN(n1261) );
XOR2_X1 U925 ( .A(n1262), .B(KEYINPUT42), .Z(n1260) );
NAND2_X1 U926 ( .A1(G116), .A2(n1225), .ZN(n1262) );
NAND3_X1 U927 ( .A1(n1256), .A2(n1060), .A3(n1087), .ZN(n1225) );
INV_X1 U928 ( .A(n1109), .ZN(n1060) );
NAND2_X1 U929 ( .A1(n1259), .A2(n1236), .ZN(n1109) );
INV_X1 U930 ( .A(n1258), .ZN(n1236) );
XOR2_X1 U931 ( .A(n1263), .B(n1224), .Z(G15) );
NAND3_X1 U932 ( .A1(n1256), .A2(n1179), .A3(n1087), .ZN(n1224) );
NOR2_X1 U933 ( .A1(n1078), .A2(n1079), .ZN(n1087) );
INV_X1 U934 ( .A(n1108), .ZN(n1179) );
NAND2_X1 U935 ( .A1(n1258), .A2(n1235), .ZN(n1108) );
INV_X1 U936 ( .A(n1259), .ZN(n1235) );
AND2_X1 U937 ( .A1(n1252), .A2(n1264), .ZN(n1256) );
NOR3_X1 U938 ( .A1(n1082), .A2(n1107), .A3(n1265), .ZN(n1252) );
INV_X1 U939 ( .A(n1067), .ZN(n1107) );
XNOR2_X1 U940 ( .A(G110), .B(n1223), .ZN(G12) );
NAND3_X1 U941 ( .A1(n1078), .A2(n1079), .A3(n1249), .ZN(n1223) );
NOR3_X1 U942 ( .A1(n1082), .A2(n1230), .A3(n1104), .ZN(n1249) );
NAND2_X1 U943 ( .A1(n1072), .A2(n1217), .ZN(n1104) );
INV_X1 U944 ( .A(n1228), .ZN(n1217) );
NAND2_X1 U945 ( .A1(n1265), .A2(n1067), .ZN(n1228) );
NAND2_X1 U946 ( .A1(G221), .A2(n1266), .ZN(n1067) );
INV_X1 U947 ( .A(n1070), .ZN(n1265) );
XOR2_X1 U948 ( .A(n1098), .B(G469), .Z(n1070) );
NAND2_X1 U949 ( .A1(n1267), .A2(n1268), .ZN(n1098) );
XOR2_X1 U950 ( .A(n1269), .B(n1270), .Z(n1267) );
XNOR2_X1 U951 ( .A(n1194), .B(n1197), .ZN(n1270) );
XOR2_X1 U952 ( .A(n1191), .B(KEYINPUT18), .Z(n1197) );
XNOR2_X1 U953 ( .A(n1271), .B(n1272), .ZN(n1194) );
XOR2_X1 U954 ( .A(n1273), .B(n1274), .Z(n1272) );
NAND2_X1 U955 ( .A1(n1275), .A2(n1231), .ZN(n1274) );
XOR2_X1 U956 ( .A(KEYINPUT47), .B(G227), .Z(n1275) );
NAND2_X1 U957 ( .A1(n1276), .A2(n1277), .ZN(n1273) );
NAND3_X1 U958 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1277) );
NAND3_X1 U959 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1278) );
OR2_X1 U960 ( .A1(n1284), .A2(KEYINPUT14), .ZN(n1282) );
NAND2_X1 U961 ( .A1(KEYINPUT14), .A2(G101), .ZN(n1281) );
NAND4_X1 U962 ( .A1(n1285), .A2(n1284), .A3(n1286), .A4(n1287), .ZN(n1276) );
NAND2_X1 U963 ( .A1(KEYINPUT14), .A2(n1250), .ZN(n1287) );
OR2_X1 U964 ( .A1(n1283), .A2(KEYINPUT14), .ZN(n1286) );
NAND2_X1 U965 ( .A1(n1280), .A2(n1279), .ZN(n1285) );
INV_X1 U966 ( .A(KEYINPUT55), .ZN(n1279) );
XOR2_X1 U967 ( .A(n1127), .B(n1288), .Z(n1271) );
XOR2_X1 U968 ( .A(n1289), .B(n1290), .Z(n1127) );
NAND2_X1 U969 ( .A1(KEYINPUT33), .A2(n1291), .ZN(n1289) );
XOR2_X1 U970 ( .A(G143), .B(n1292), .Z(n1291) );
NOR2_X1 U971 ( .A1(KEYINPUT25), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U972 ( .A(KEYINPUT38), .B(KEYINPUT32), .ZN(n1269) );
INV_X1 U973 ( .A(n1093), .ZN(n1072) );
NAND2_X1 U974 ( .A1(n1258), .A2(n1259), .ZN(n1093) );
XOR2_X1 U975 ( .A(n1294), .B(G475), .Z(n1259) );
OR2_X1 U976 ( .A1(n1171), .A2(G902), .ZN(n1294) );
XNOR2_X1 U977 ( .A(n1295), .B(n1296), .ZN(n1171) );
XOR2_X1 U978 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U979 ( .A(n1299), .B(n1300), .Z(n1298) );
NAND2_X1 U980 ( .A1(n1301), .A2(KEYINPUT52), .ZN(n1300) );
XOR2_X1 U981 ( .A(n1302), .B(G143), .Z(n1301) );
NAND2_X1 U982 ( .A1(G214), .A2(n1303), .ZN(n1302) );
NAND2_X1 U983 ( .A1(n1304), .A2(n1305), .ZN(n1299) );
NAND2_X1 U984 ( .A1(G113), .A2(n1255), .ZN(n1305) );
XOR2_X1 U985 ( .A(KEYINPUT35), .B(n1306), .Z(n1304) );
NOR2_X1 U986 ( .A1(G113), .A2(n1255), .ZN(n1306) );
XOR2_X1 U987 ( .A(n1307), .B(n1308), .Z(n1295) );
XOR2_X1 U988 ( .A(G131), .B(G104), .Z(n1308) );
NAND2_X1 U989 ( .A1(KEYINPUT45), .A2(n1309), .ZN(n1307) );
INV_X1 U990 ( .A(G140), .ZN(n1309) );
XOR2_X1 U991 ( .A(n1310), .B(G478), .Z(n1258) );
OR2_X1 U992 ( .A1(n1163), .A2(G902), .ZN(n1310) );
XNOR2_X1 U993 ( .A(n1311), .B(n1312), .ZN(n1163) );
AND2_X1 U994 ( .A1(n1313), .A2(G217), .ZN(n1312) );
NAND2_X1 U995 ( .A1(KEYINPUT22), .A2(n1314), .ZN(n1311) );
XOR2_X1 U996 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U997 ( .A(n1317), .B(n1318), .ZN(n1316) );
NOR2_X1 U998 ( .A1(KEYINPUT46), .A2(n1319), .ZN(n1318) );
XOR2_X1 U999 ( .A(n1320), .B(n1321), .Z(n1319) );
NAND2_X1 U1000 ( .A1(n1322), .A2(KEYINPUT36), .ZN(n1320) );
XOR2_X1 U1001 ( .A(G116), .B(n1255), .Z(n1322) );
INV_X1 U1002 ( .A(G122), .ZN(n1255) );
NAND2_X1 U1003 ( .A1(KEYINPUT37), .A2(n1323), .ZN(n1317) );
XOR2_X1 U1004 ( .A(G143), .B(G134), .Z(n1315) );
INV_X1 U1005 ( .A(n1264), .ZN(n1230) );
NAND2_X1 U1006 ( .A1(n1088), .A2(n1324), .ZN(n1264) );
NAND4_X1 U1007 ( .A1(G953), .A2(G902), .A3(n1254), .A4(n1146), .ZN(n1324) );
INV_X1 U1008 ( .A(G898), .ZN(n1146) );
NAND3_X1 U1009 ( .A1(n1254), .A2(n1231), .A3(G952), .ZN(n1088) );
NAND2_X1 U1010 ( .A1(G237), .A2(n1325), .ZN(n1254) );
XOR2_X1 U1011 ( .A(KEYINPUT41), .B(G234), .Z(n1325) );
INV_X1 U1012 ( .A(n1061), .ZN(n1082) );
NOR2_X1 U1013 ( .A1(n1085), .A2(n1084), .ZN(n1061) );
AND2_X1 U1014 ( .A1(G214), .A2(n1326), .ZN(n1084) );
NAND2_X1 U1015 ( .A1(n1268), .A2(n1327), .ZN(n1326) );
INV_X1 U1016 ( .A(n1241), .ZN(n1085) );
NAND2_X1 U1017 ( .A1(n1328), .A2(n1329), .ZN(n1241) );
NAND2_X1 U1018 ( .A1(G210), .A2(n1330), .ZN(n1329) );
NAND2_X1 U1019 ( .A1(n1268), .A2(n1331), .ZN(n1330) );
OR2_X1 U1020 ( .A1(n1327), .A2(n1332), .ZN(n1331) );
INV_X1 U1021 ( .A(G237), .ZN(n1327) );
NAND3_X1 U1022 ( .A1(n1333), .A2(n1268), .A3(n1332), .ZN(n1328) );
XOR2_X1 U1023 ( .A(n1200), .B(KEYINPUT11), .Z(n1332) );
XNOR2_X1 U1024 ( .A(n1334), .B(n1335), .ZN(n1200) );
XOR2_X1 U1025 ( .A(n1150), .B(n1151), .Z(n1335) );
INV_X1 U1026 ( .A(n1147), .ZN(n1151) );
NAND2_X1 U1027 ( .A1(n1336), .A2(n1337), .ZN(n1147) );
NAND2_X1 U1028 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
NAND2_X1 U1029 ( .A1(n1283), .A2(n1284), .ZN(n1339) );
NAND2_X1 U1030 ( .A1(n1321), .A2(n1250), .ZN(n1284) );
NAND2_X1 U1031 ( .A1(G101), .A2(n1340), .ZN(n1283) );
NAND2_X1 U1032 ( .A1(n1341), .A2(n1280), .ZN(n1336) );
INV_X1 U1033 ( .A(n1338), .ZN(n1280) );
XNOR2_X1 U1034 ( .A(G104), .B(KEYINPUT28), .ZN(n1338) );
XOR2_X1 U1035 ( .A(G101), .B(n1340), .Z(n1341) );
INV_X1 U1036 ( .A(n1321), .ZN(n1340) );
XNOR2_X1 U1037 ( .A(G107), .B(KEYINPUT12), .ZN(n1321) );
INV_X1 U1038 ( .A(n1149), .ZN(n1150) );
XOR2_X1 U1039 ( .A(n1342), .B(n1343), .Z(n1149) );
XOR2_X1 U1040 ( .A(n1344), .B(n1345), .Z(n1343) );
XOR2_X1 U1041 ( .A(G113), .B(G110), .Z(n1345) );
NOR2_X1 U1042 ( .A1(G119), .A2(KEYINPUT8), .ZN(n1344) );
XNOR2_X1 U1043 ( .A(G116), .B(n1346), .ZN(n1342) );
XOR2_X1 U1044 ( .A(KEYINPUT4), .B(G122), .Z(n1346) );
XOR2_X1 U1045 ( .A(n1347), .B(n1297), .Z(n1334) );
XOR2_X1 U1046 ( .A(n1348), .B(n1349), .Z(n1347) );
AND2_X1 U1047 ( .A1(n1231), .A2(G224), .ZN(n1349) );
NAND2_X1 U1048 ( .A1(G210), .A2(G237), .ZN(n1333) );
INV_X1 U1049 ( .A(n1083), .ZN(n1079) );
XNOR2_X1 U1050 ( .A(n1350), .B(n1157), .ZN(n1083) );
NAND2_X1 U1051 ( .A1(G217), .A2(n1266), .ZN(n1157) );
NAND2_X1 U1052 ( .A1(G234), .A2(n1268), .ZN(n1266) );
OR2_X1 U1053 ( .A1(n1160), .A2(G902), .ZN(n1350) );
XNOR2_X1 U1054 ( .A(n1351), .B(n1352), .ZN(n1160) );
XOR2_X1 U1055 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1056 ( .A(n1355), .B(G119), .Z(n1354) );
NAND2_X1 U1057 ( .A1(G221), .A2(n1313), .ZN(n1355) );
AND2_X1 U1058 ( .A1(G234), .A2(n1231), .ZN(n1313) );
INV_X1 U1059 ( .A(G953), .ZN(n1231) );
XNOR2_X1 U1060 ( .A(G137), .B(KEYINPUT54), .ZN(n1353) );
XNOR2_X1 U1061 ( .A(n1288), .B(n1356), .ZN(n1351) );
XOR2_X1 U1062 ( .A(n1323), .B(n1297), .Z(n1356) );
XNOR2_X1 U1063 ( .A(G125), .B(n1293), .ZN(n1297) );
INV_X1 U1064 ( .A(G146), .ZN(n1293) );
XOR2_X1 U1065 ( .A(G110), .B(G140), .Z(n1288) );
INV_X1 U1066 ( .A(n1229), .ZN(n1078) );
XOR2_X1 U1067 ( .A(n1095), .B(n1357), .Z(n1229) );
NOR2_X1 U1068 ( .A1(n1094), .A2(KEYINPUT20), .ZN(n1357) );
AND2_X1 U1069 ( .A1(n1358), .A2(n1268), .ZN(n1094) );
INV_X1 U1070 ( .A(G902), .ZN(n1268) );
XOR2_X1 U1071 ( .A(n1359), .B(n1360), .Z(n1358) );
NAND3_X1 U1072 ( .A1(KEYINPUT62), .A2(n1361), .A3(n1362), .ZN(n1360) );
XOR2_X1 U1073 ( .A(n1363), .B(KEYINPUT21), .Z(n1362) );
NAND2_X1 U1074 ( .A1(n1184), .A2(n1364), .ZN(n1363) );
OR2_X1 U1075 ( .A1(n1364), .A2(n1184), .ZN(n1361) );
XNOR2_X1 U1076 ( .A(n1365), .B(n1366), .ZN(n1184) );
XOR2_X1 U1077 ( .A(G119), .B(G116), .Z(n1366) );
NAND2_X1 U1078 ( .A1(KEYINPUT17), .A2(n1263), .ZN(n1365) );
INV_X1 U1079 ( .A(G113), .ZN(n1263) );
NAND3_X1 U1080 ( .A1(n1367), .A2(n1368), .A3(n1369), .ZN(n1364) );
NAND2_X1 U1081 ( .A1(KEYINPUT6), .A2(n1190), .ZN(n1369) );
NAND3_X1 U1082 ( .A1(n1370), .A2(n1371), .A3(n1372), .ZN(n1368) );
INV_X1 U1083 ( .A(n1190), .ZN(n1370) );
NAND2_X1 U1084 ( .A1(n1191), .A2(n1373), .ZN(n1367) );
NAND2_X1 U1085 ( .A1(n1374), .A2(n1371), .ZN(n1373) );
INV_X1 U1086 ( .A(KEYINPUT6), .ZN(n1371) );
XOR2_X1 U1087 ( .A(n1190), .B(KEYINPUT60), .Z(n1374) );
XOR2_X1 U1088 ( .A(n1348), .B(n1375), .Z(n1190) );
XOR2_X1 U1089 ( .A(KEYINPUT44), .B(G146), .Z(n1375) );
XOR2_X1 U1090 ( .A(n1376), .B(n1290), .Z(n1348) );
XOR2_X1 U1091 ( .A(n1323), .B(KEYINPUT57), .Z(n1290) );
XOR2_X1 U1092 ( .A(G128), .B(KEYINPUT0), .Z(n1323) );
XOR2_X1 U1093 ( .A(n1233), .B(KEYINPUT10), .Z(n1376) );
INV_X1 U1094 ( .A(G143), .ZN(n1233) );
INV_X1 U1095 ( .A(n1372), .ZN(n1191) );
XOR2_X1 U1096 ( .A(n1377), .B(n1378), .Z(n1372) );
NOR2_X1 U1097 ( .A1(G137), .A2(KEYINPUT56), .ZN(n1378) );
XOR2_X1 U1098 ( .A(n1240), .B(G134), .Z(n1377) );
INV_X1 U1099 ( .A(G131), .ZN(n1240) );
NAND3_X1 U1100 ( .A1(n1379), .A2(n1380), .A3(n1381), .ZN(n1359) );
NAND2_X1 U1101 ( .A1(n1186), .A2(n1250), .ZN(n1381) );
NAND2_X1 U1102 ( .A1(KEYINPUT9), .A2(n1382), .ZN(n1380) );
NAND2_X1 U1103 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
XOR2_X1 U1104 ( .A(KEYINPUT50), .B(G101), .Z(n1384) );
INV_X1 U1105 ( .A(n1186), .ZN(n1383) );
NAND2_X1 U1106 ( .A1(n1385), .A2(n1386), .ZN(n1379) );
INV_X1 U1107 ( .A(KEYINPUT9), .ZN(n1386) );
NAND2_X1 U1108 ( .A1(n1387), .A2(n1388), .ZN(n1385) );
NAND2_X1 U1109 ( .A1(KEYINPUT50), .A2(n1250), .ZN(n1388) );
OR3_X1 U1110 ( .A1(n1186), .A2(KEYINPUT50), .A3(n1250), .ZN(n1387) );
INV_X1 U1111 ( .A(G101), .ZN(n1250) );
NAND2_X1 U1112 ( .A1(G210), .A2(n1303), .ZN(n1186) );
NOR2_X1 U1113 ( .A1(G953), .A2(G237), .ZN(n1303) );
INV_X1 U1114 ( .A(G472), .ZN(n1095) );
endmodule


