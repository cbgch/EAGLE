//Key = 1010100100101000011010000111111000000010001100000011111001001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378;

XOR2_X1 U743 ( .A(G107), .B(n1047), .Z(G9) );
NOR4_X1 U744 ( .A1(KEYINPUT44), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1047) );
NOR2_X1 U745 ( .A1(n1051), .A2(n1052), .ZN(G75) );
NOR3_X1 U746 ( .A1(n1053), .A2(G953), .A3(G952), .ZN(n1052) );
NOR4_X1 U747 ( .A1(n1054), .A2(n1055), .A3(n1053), .A4(n1056), .ZN(n1051) );
AND4_X1 U748 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1053) );
NOR3_X1 U749 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NOR2_X1 U750 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
INV_X1 U751 ( .A(n1066), .ZN(n1062) );
NAND3_X1 U752 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1061) );
NOR3_X1 U753 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1059) );
XOR2_X1 U754 ( .A(n1073), .B(KEYINPUT2), .Z(n1071) );
XNOR2_X1 U755 ( .A(n1074), .B(n1075), .ZN(n1070) );
NOR2_X1 U756 ( .A1(KEYINPUT6), .A2(n1076), .ZN(n1075) );
XOR2_X1 U757 ( .A(n1077), .B(n1078), .Z(n1058) );
XOR2_X1 U758 ( .A(KEYINPUT38), .B(G469), .Z(n1078) );
NAND2_X1 U759 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
XOR2_X1 U760 ( .A(KEYINPUT7), .B(KEYINPUT46), .Z(n1079) );
XOR2_X1 U761 ( .A(n1081), .B(G472), .Z(n1057) );
NAND4_X1 U762 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1054) );
NAND4_X1 U763 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1084) );
NOR2_X1 U764 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U765 ( .A1(n1092), .A2(n1049), .ZN(n1087) );
NAND3_X1 U766 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1083) );
INV_X1 U767 ( .A(n1090), .ZN(n1095) );
NAND2_X1 U768 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NAND3_X1 U769 ( .A1(n1086), .A2(n1098), .A3(n1088), .ZN(n1097) );
NAND2_X1 U770 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U771 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
INV_X1 U772 ( .A(n1103), .ZN(n1099) );
NAND2_X1 U773 ( .A1(n1104), .A2(n1105), .ZN(n1096) );
NAND2_X1 U774 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U775 ( .A1(n1088), .A2(n1108), .ZN(n1107) );
OR2_X1 U776 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U777 ( .A1(n1086), .A2(n1111), .ZN(n1106) );
NAND2_X1 U778 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
OR2_X1 U779 ( .A1(n1114), .A2(n1069), .ZN(n1113) );
XOR2_X1 U780 ( .A(n1115), .B(n1116), .Z(G72) );
XOR2_X1 U781 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U782 ( .A1(G953), .A2(n1119), .ZN(n1118) );
NAND2_X1 U783 ( .A1(G900), .A2(G227), .ZN(n1119) );
NAND2_X1 U784 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
NAND2_X1 U785 ( .A1(G953), .A2(n1122), .ZN(n1121) );
XOR2_X1 U786 ( .A(n1123), .B(KEYINPUT12), .Z(n1120) );
NAND3_X1 U787 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
NAND2_X1 U788 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
OR3_X1 U789 ( .A1(n1128), .A2(n1127), .A3(n1129), .ZN(n1125) );
INV_X1 U790 ( .A(KEYINPUT53), .ZN(n1128) );
NAND2_X1 U791 ( .A1(n1129), .A2(n1130), .ZN(n1124) );
NAND2_X1 U792 ( .A1(n1131), .A2(KEYINPUT53), .ZN(n1130) );
XNOR2_X1 U793 ( .A(n1127), .B(KEYINPUT48), .ZN(n1131) );
XOR2_X1 U794 ( .A(n1132), .B(n1133), .Z(n1127) );
XOR2_X1 U795 ( .A(n1134), .B(n1135), .Z(n1129) );
XOR2_X1 U796 ( .A(n1136), .B(n1137), .Z(n1135) );
NOR2_X1 U797 ( .A1(KEYINPUT55), .A2(n1138), .ZN(n1136) );
INV_X1 U798 ( .A(G134), .ZN(n1138) );
XOR2_X1 U799 ( .A(n1139), .B(G137), .Z(n1134) );
NOR2_X1 U800 ( .A1(n1140), .A2(G953), .ZN(n1115) );
XOR2_X1 U801 ( .A(n1141), .B(n1142), .Z(G69) );
NOR2_X1 U802 ( .A1(n1143), .A2(n1085), .ZN(n1142) );
NOR2_X1 U803 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND2_X1 U804 ( .A1(n1146), .A2(n1147), .ZN(n1141) );
NAND2_X1 U805 ( .A1(n1148), .A2(n1085), .ZN(n1147) );
XNOR2_X1 U806 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR2_X1 U807 ( .A1(n1151), .A2(n1055), .ZN(n1150) );
XOR2_X1 U808 ( .A(n1082), .B(KEYINPUT4), .Z(n1151) );
NAND3_X1 U809 ( .A1(G898), .A2(n1149), .A3(G953), .ZN(n1146) );
NOR2_X1 U810 ( .A1(n1152), .A2(n1153), .ZN(G66) );
XOR2_X1 U811 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND3_X1 U812 ( .A1(G217), .A2(n1156), .A3(n1157), .ZN(n1154) );
NOR2_X1 U813 ( .A1(n1152), .A2(n1158), .ZN(G63) );
NOR2_X1 U814 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U815 ( .A(KEYINPUT34), .B(n1161), .Z(n1160) );
AND2_X1 U816 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NOR2_X1 U817 ( .A1(n1163), .A2(n1162), .ZN(n1159) );
NOR2_X1 U818 ( .A1(n1164), .A2(n1065), .ZN(n1163) );
NOR2_X1 U819 ( .A1(n1152), .A2(n1165), .ZN(G60) );
XOR2_X1 U820 ( .A(n1166), .B(n1167), .Z(n1165) );
NAND2_X1 U821 ( .A1(n1157), .A2(G475), .ZN(n1166) );
XOR2_X1 U822 ( .A(n1168), .B(n1169), .Z(G6) );
NAND2_X1 U823 ( .A1(n1170), .A2(G104), .ZN(n1168) );
XNOR2_X1 U824 ( .A(KEYINPUT9), .B(KEYINPUT19), .ZN(n1170) );
NOR2_X1 U825 ( .A1(n1152), .A2(n1171), .ZN(G57) );
XNOR2_X1 U826 ( .A(n1172), .B(n1173), .ZN(n1171) );
NAND2_X1 U827 ( .A1(n1174), .A2(n1175), .ZN(n1172) );
NAND2_X1 U828 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U829 ( .A(n1178), .B(KEYINPUT11), .Z(n1177) );
NAND2_X1 U830 ( .A1(n1157), .A2(G472), .ZN(n1178) );
INV_X1 U831 ( .A(n1164), .ZN(n1157) );
OR3_X1 U832 ( .A1(n1164), .A2(n1179), .A3(n1176), .ZN(n1174) );
XNOR2_X1 U833 ( .A(n1180), .B(n1181), .ZN(n1176) );
NOR2_X1 U834 ( .A1(n1152), .A2(n1182), .ZN(G54) );
XOR2_X1 U835 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U836 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U837 ( .A(n1187), .B(n1188), .Z(n1186) );
NOR2_X1 U838 ( .A1(n1189), .A2(n1164), .ZN(n1188) );
NAND2_X1 U839 ( .A1(KEYINPUT0), .A2(n1190), .ZN(n1187) );
XOR2_X1 U840 ( .A(n1191), .B(n1192), .Z(n1183) );
NOR2_X1 U841 ( .A1(n1152), .A2(n1193), .ZN(G51) );
XOR2_X1 U842 ( .A(n1194), .B(n1195), .Z(n1193) );
OR2_X1 U843 ( .A1(n1164), .A2(n1074), .ZN(n1195) );
NAND2_X1 U844 ( .A1(n1196), .A2(n1197), .ZN(n1164) );
NAND3_X1 U845 ( .A1(n1198), .A2(n1082), .A3(n1199), .ZN(n1197) );
XOR2_X1 U846 ( .A(KEYINPUT42), .B(n1056), .Z(n1199) );
AND2_X1 U847 ( .A1(n1200), .A2(n1201), .ZN(n1056) );
NAND2_X1 U848 ( .A1(n1140), .A2(n1202), .ZN(n1201) );
INV_X1 U849 ( .A(KEYINPUT37), .ZN(n1202) );
AND2_X1 U850 ( .A1(n1203), .A2(n1204), .ZN(n1140) );
NOR4_X1 U851 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
INV_X1 U852 ( .A(n1209), .ZN(n1207) );
AND4_X1 U853 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1203) );
NAND2_X1 U854 ( .A1(n1205), .A2(KEYINPUT37), .ZN(n1200) );
INV_X1 U855 ( .A(n1055), .ZN(n1198) );
NAND4_X1 U856 ( .A1(n1214), .A2(n1215), .A3(n1169), .A4(n1216), .ZN(n1055) );
NOR3_X1 U857 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1216) );
NOR3_X1 U858 ( .A1(n1050), .A2(n1048), .A3(n1049), .ZN(n1219) );
INV_X1 U859 ( .A(n1086), .ZN(n1048) );
NOR3_X1 U860 ( .A1(n1091), .A2(n1220), .A3(n1221), .ZN(n1218) );
NOR2_X1 U861 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
NOR2_X1 U862 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NOR2_X1 U863 ( .A1(n1049), .A2(n1226), .ZN(n1222) );
NOR2_X1 U864 ( .A1(n1112), .A2(n1227), .ZN(n1217) );
NAND3_X1 U865 ( .A1(n1086), .A2(n1228), .A3(n1229), .ZN(n1169) );
XOR2_X1 U866 ( .A(KEYINPUT35), .B(G902), .Z(n1196) );
NAND2_X1 U867 ( .A1(n1230), .A2(n1231), .ZN(n1194) );
NAND2_X1 U868 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
XOR2_X1 U869 ( .A(KEYINPUT43), .B(n1234), .Z(n1230) );
NOR2_X1 U870 ( .A1(n1233), .A2(n1232), .ZN(n1234) );
XNOR2_X1 U871 ( .A(n1235), .B(KEYINPUT57), .ZN(n1232) );
NOR2_X1 U872 ( .A1(n1085), .A2(G952), .ZN(n1152) );
XNOR2_X1 U873 ( .A(G146), .B(n1210), .ZN(G48) );
NAND3_X1 U874 ( .A1(n1236), .A2(n1228), .A3(n1237), .ZN(n1210) );
XOR2_X1 U875 ( .A(n1238), .B(n1213), .Z(G45) );
NAND4_X1 U876 ( .A1(n1239), .A2(n1236), .A3(n1072), .A4(n1240), .ZN(n1213) );
INV_X1 U877 ( .A(n1241), .ZN(n1072) );
XOR2_X1 U878 ( .A(n1133), .B(n1212), .Z(G42) );
NAND4_X1 U879 ( .A1(n1228), .A2(n1242), .A3(n1109), .A4(n1243), .ZN(n1212) );
AND2_X1 U880 ( .A1(n1103), .A2(n1088), .ZN(n1243) );
XOR2_X1 U881 ( .A(n1208), .B(n1244), .Z(G39) );
NOR2_X1 U882 ( .A1(KEYINPUT5), .A2(n1245), .ZN(n1244) );
INV_X1 U883 ( .A(G137), .ZN(n1245) );
AND3_X1 U884 ( .A1(n1088), .A2(n1093), .A3(n1237), .ZN(n1208) );
XOR2_X1 U885 ( .A(n1246), .B(G134), .Z(G36) );
NAND2_X1 U886 ( .A1(KEYINPUT28), .A2(n1211), .ZN(n1246) );
NAND3_X1 U887 ( .A1(n1088), .A2(n1247), .A3(n1239), .ZN(n1211) );
XOR2_X1 U888 ( .A(n1139), .B(n1209), .Z(G33) );
NAND3_X1 U889 ( .A1(n1088), .A2(n1228), .A3(n1239), .ZN(n1209) );
AND3_X1 U890 ( .A1(n1103), .A2(n1242), .A3(n1110), .ZN(n1239) );
NOR2_X1 U891 ( .A1(n1114), .A2(n1248), .ZN(n1088) );
XOR2_X1 U892 ( .A(G128), .B(n1206), .Z(G30) );
AND3_X1 U893 ( .A1(n1247), .A2(n1236), .A3(n1237), .ZN(n1206) );
AND3_X1 U894 ( .A1(n1103), .A2(n1242), .A3(n1249), .ZN(n1237) );
INV_X1 U895 ( .A(n1049), .ZN(n1247) );
XOR2_X1 U896 ( .A(n1250), .B(n1214), .Z(G3) );
NAND3_X1 U897 ( .A1(n1093), .A2(n1229), .A3(n1110), .ZN(n1214) );
XOR2_X1 U898 ( .A(n1251), .B(G125), .Z(G27) );
NAND2_X1 U899 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND3_X1 U900 ( .A1(n1254), .A2(n1092), .A3(n1255), .ZN(n1253) );
INV_X1 U901 ( .A(KEYINPUT51), .ZN(n1255) );
INV_X1 U902 ( .A(n1228), .ZN(n1092) );
NAND2_X1 U903 ( .A1(KEYINPUT51), .A2(n1205), .ZN(n1252) );
AND2_X1 U904 ( .A1(n1254), .A2(n1228), .ZN(n1205) );
AND4_X1 U905 ( .A1(n1104), .A2(n1236), .A3(n1109), .A4(n1242), .ZN(n1254) );
NAND2_X1 U906 ( .A1(n1090), .A2(n1256), .ZN(n1242) );
NAND4_X1 U907 ( .A1(G902), .A2(G953), .A3(n1257), .A4(n1122), .ZN(n1256) );
INV_X1 U908 ( .A(G900), .ZN(n1122) );
XNOR2_X1 U909 ( .A(G122), .B(n1215), .ZN(G24) );
NAND4_X1 U910 ( .A1(n1104), .A2(n1086), .A3(n1258), .A4(n1259), .ZN(n1215) );
NOR2_X1 U911 ( .A1(n1260), .A2(n1241), .ZN(n1258) );
NOR2_X1 U912 ( .A1(n1261), .A2(n1262), .ZN(n1086) );
XNOR2_X1 U913 ( .A(G119), .B(n1263), .ZN(G21) );
NAND4_X1 U914 ( .A1(KEYINPUT50), .A2(n1249), .A3(n1264), .A4(n1104), .ZN(n1263) );
NOR2_X1 U915 ( .A1(n1221), .A2(n1224), .ZN(n1264) );
XOR2_X1 U916 ( .A(n1265), .B(n1266), .Z(G18) );
NOR2_X1 U917 ( .A1(KEYINPUT23), .A2(n1267), .ZN(n1266) );
NOR4_X1 U918 ( .A1(n1268), .A2(n1221), .A3(n1049), .A4(n1226), .ZN(n1265) );
NAND2_X1 U919 ( .A1(n1241), .A2(n1240), .ZN(n1049) );
XOR2_X1 U920 ( .A(n1091), .B(KEYINPUT13), .Z(n1268) );
XOR2_X1 U921 ( .A(G113), .B(n1269), .Z(G15) );
NOR2_X1 U922 ( .A1(n1270), .A2(n1112), .ZN(n1269) );
XOR2_X1 U923 ( .A(n1227), .B(KEYINPUT32), .Z(n1270) );
NAND4_X1 U924 ( .A1(n1110), .A2(n1104), .A3(n1228), .A4(n1271), .ZN(n1227) );
NAND2_X1 U925 ( .A1(n1272), .A2(n1273), .ZN(n1228) );
OR3_X1 U926 ( .A1(n1240), .A2(n1241), .A3(KEYINPUT41), .ZN(n1273) );
NAND2_X1 U927 ( .A1(KEYINPUT41), .A2(n1093), .ZN(n1272) );
INV_X1 U928 ( .A(n1091), .ZN(n1104) );
NAND2_X1 U929 ( .A1(n1102), .A2(n1067), .ZN(n1091) );
INV_X1 U930 ( .A(n1226), .ZN(n1110) );
NAND2_X1 U931 ( .A1(n1274), .A2(n1262), .ZN(n1226) );
XNOR2_X1 U932 ( .A(G110), .B(n1082), .ZN(G12) );
NAND3_X1 U933 ( .A1(n1229), .A2(n1109), .A3(n1093), .ZN(n1082) );
INV_X1 U934 ( .A(n1224), .ZN(n1093) );
NAND2_X1 U935 ( .A1(n1260), .A2(n1241), .ZN(n1224) );
XOR2_X1 U936 ( .A(n1275), .B(G475), .Z(n1241) );
NAND2_X1 U937 ( .A1(n1167), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U938 ( .A(n1277), .B(n1278), .ZN(n1167) );
XOR2_X1 U939 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U940 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR2_X1 U941 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
XOR2_X1 U942 ( .A(n1285), .B(KEYINPUT20), .Z(n1284) );
NAND2_X1 U943 ( .A1(n1286), .A2(n1139), .ZN(n1285) );
NOR2_X1 U944 ( .A1(n1139), .A2(n1286), .ZN(n1283) );
XOR2_X1 U945 ( .A(n1287), .B(n1238), .Z(n1286) );
INV_X1 U946 ( .A(G143), .ZN(n1238) );
NAND2_X1 U947 ( .A1(n1288), .A2(G214), .ZN(n1287) );
NAND2_X1 U948 ( .A1(KEYINPUT27), .A2(n1289), .ZN(n1281) );
XOR2_X1 U949 ( .A(n1290), .B(n1291), .Z(n1277) );
XOR2_X1 U950 ( .A(KEYINPUT45), .B(G140), .Z(n1291) );
XNOR2_X1 U951 ( .A(G104), .B(G113), .ZN(n1290) );
INV_X1 U952 ( .A(n1240), .ZN(n1260) );
NAND3_X1 U953 ( .A1(n1292), .A2(n1293), .A3(n1068), .ZN(n1240) );
NAND2_X1 U954 ( .A1(n1064), .A2(n1065), .ZN(n1068) );
NAND2_X1 U955 ( .A1(KEYINPUT1), .A2(n1065), .ZN(n1293) );
OR3_X1 U956 ( .A1(n1064), .A2(KEYINPUT1), .A3(n1065), .ZN(n1292) );
INV_X1 U957 ( .A(G478), .ZN(n1065) );
NOR2_X1 U958 ( .A1(n1162), .A2(G902), .ZN(n1064) );
XOR2_X1 U959 ( .A(n1294), .B(n1295), .Z(n1162) );
XOR2_X1 U960 ( .A(G128), .B(n1296), .Z(n1295) );
XOR2_X1 U961 ( .A(G143), .B(G134), .Z(n1296) );
XOR2_X1 U962 ( .A(n1297), .B(n1298), .Z(n1294) );
XOR2_X1 U963 ( .A(n1299), .B(G107), .Z(n1297) );
NAND2_X1 U964 ( .A1(G217), .A2(n1300), .ZN(n1299) );
NAND2_X1 U965 ( .A1(n1301), .A2(n1302), .ZN(n1109) );
NAND2_X1 U966 ( .A1(n1249), .A2(n1303), .ZN(n1302) );
INV_X1 U967 ( .A(n1225), .ZN(n1249) );
NAND2_X1 U968 ( .A1(n1262), .A2(n1261), .ZN(n1225) );
OR3_X1 U969 ( .A1(n1262), .A2(n1274), .A3(n1303), .ZN(n1301) );
INV_X1 U970 ( .A(KEYINPUT25), .ZN(n1303) );
INV_X1 U971 ( .A(n1261), .ZN(n1274) );
NAND2_X1 U972 ( .A1(n1066), .A2(n1073), .ZN(n1261) );
NAND3_X1 U973 ( .A1(n1304), .A2(n1276), .A3(n1305), .ZN(n1073) );
NAND2_X1 U974 ( .A1(G217), .A2(n1156), .ZN(n1304) );
NAND3_X1 U975 ( .A1(n1306), .A2(n1156), .A3(G217), .ZN(n1066) );
NAND2_X1 U976 ( .A1(n1305), .A2(n1276), .ZN(n1306) );
XNOR2_X1 U977 ( .A(n1155), .B(KEYINPUT63), .ZN(n1305) );
XNOR2_X1 U978 ( .A(n1307), .B(n1308), .ZN(n1155) );
XOR2_X1 U979 ( .A(n1309), .B(n1310), .Z(n1308) );
XNOR2_X1 U980 ( .A(n1311), .B(n1312), .ZN(n1310) );
NOR2_X1 U981 ( .A1(KEYINPUT58), .A2(n1133), .ZN(n1312) );
NOR2_X1 U982 ( .A1(KEYINPUT59), .A2(n1313), .ZN(n1311) );
XOR2_X1 U983 ( .A(KEYINPUT54), .B(G137), .Z(n1313) );
XNOR2_X1 U984 ( .A(G128), .B(KEYINPUT21), .ZN(n1309) );
XNOR2_X1 U985 ( .A(n1314), .B(n1315), .ZN(n1307) );
XOR2_X1 U986 ( .A(n1316), .B(n1279), .Z(n1315) );
XOR2_X1 U987 ( .A(G146), .B(n1132), .Z(n1279) );
INV_X1 U988 ( .A(G125), .ZN(n1132) );
NAND2_X1 U989 ( .A1(n1300), .A2(G221), .ZN(n1316) );
AND2_X1 U990 ( .A1(G234), .A2(n1085), .ZN(n1300) );
XNOR2_X1 U991 ( .A(n1081), .B(n1317), .ZN(n1262) );
NOR2_X1 U992 ( .A1(KEYINPUT16), .A2(n1179), .ZN(n1317) );
INV_X1 U993 ( .A(G472), .ZN(n1179) );
NAND2_X1 U994 ( .A1(n1318), .A2(n1319), .ZN(n1081) );
XOR2_X1 U995 ( .A(n1320), .B(n1321), .Z(n1319) );
NOR2_X1 U996 ( .A1(KEYINPUT3), .A2(n1173), .ZN(n1321) );
XNOR2_X1 U997 ( .A(n1322), .B(n1250), .ZN(n1173) );
INV_X1 U998 ( .A(G101), .ZN(n1250) );
NAND2_X1 U999 ( .A1(n1288), .A2(G210), .ZN(n1322) );
NOR2_X1 U1000 ( .A1(G953), .A2(G237), .ZN(n1288) );
NAND3_X1 U1001 ( .A1(n1323), .A2(n1324), .A3(n1325), .ZN(n1320) );
NAND2_X1 U1002 ( .A1(KEYINPUT8), .A2(n1181), .ZN(n1325) );
NAND3_X1 U1003 ( .A1(n1326), .A2(n1327), .A3(n1180), .ZN(n1324) );
INV_X1 U1004 ( .A(KEYINPUT8), .ZN(n1327) );
OR2_X1 U1005 ( .A1(n1180), .A2(n1326), .ZN(n1323) );
NOR2_X1 U1006 ( .A1(KEYINPUT14), .A2(n1181), .ZN(n1326) );
XOR2_X1 U1007 ( .A(n1328), .B(G113), .Z(n1181) );
NAND3_X1 U1008 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1328) );
NAND2_X1 U1009 ( .A1(n1332), .A2(G116), .ZN(n1331) );
NAND2_X1 U1010 ( .A1(KEYINPUT39), .A2(n1333), .ZN(n1330) );
NAND2_X1 U1011 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
XOR2_X1 U1012 ( .A(KEYINPUT15), .B(n1267), .Z(n1334) );
NAND2_X1 U1013 ( .A1(n1336), .A2(n1337), .ZN(n1329) );
INV_X1 U1014 ( .A(KEYINPUT39), .ZN(n1337) );
NAND2_X1 U1015 ( .A1(n1338), .A2(n1339), .ZN(n1336) );
OR3_X1 U1016 ( .A1(n1332), .A2(G116), .A3(KEYINPUT15), .ZN(n1339) );
NAND2_X1 U1017 ( .A1(KEYINPUT15), .A2(G116), .ZN(n1338) );
XNOR2_X1 U1018 ( .A(n1340), .B(n1341), .ZN(n1180) );
XOR2_X1 U1019 ( .A(n1276), .B(KEYINPUT62), .Z(n1318) );
INV_X1 U1020 ( .A(n1050), .ZN(n1229) );
NAND2_X1 U1021 ( .A1(n1103), .A2(n1259), .ZN(n1050) );
INV_X1 U1022 ( .A(n1221), .ZN(n1259) );
NAND2_X1 U1023 ( .A1(n1236), .A2(n1271), .ZN(n1221) );
NAND2_X1 U1024 ( .A1(n1090), .A2(n1342), .ZN(n1271) );
NAND4_X1 U1025 ( .A1(G902), .A2(G953), .A3(n1257), .A4(n1145), .ZN(n1342) );
INV_X1 U1026 ( .A(G898), .ZN(n1145) );
NAND3_X1 U1027 ( .A1(n1257), .A2(n1085), .A3(G952), .ZN(n1090) );
INV_X1 U1028 ( .A(G953), .ZN(n1085) );
NAND2_X1 U1029 ( .A1(G237), .A2(G234), .ZN(n1257) );
INV_X1 U1030 ( .A(n1112), .ZN(n1236) );
NAND2_X1 U1031 ( .A1(n1343), .A2(n1114), .ZN(n1112) );
XNOR2_X1 U1032 ( .A(n1076), .B(n1344), .ZN(n1114) );
NOR2_X1 U1033 ( .A1(KEYINPUT47), .A2(n1074), .ZN(n1344) );
NAND2_X1 U1034 ( .A1(G210), .A2(n1345), .ZN(n1074) );
NAND2_X1 U1035 ( .A1(n1346), .A2(n1276), .ZN(n1076) );
XNOR2_X1 U1036 ( .A(n1233), .B(n1235), .ZN(n1346) );
XOR2_X1 U1037 ( .A(n1149), .B(KEYINPUT10), .Z(n1235) );
XNOR2_X1 U1038 ( .A(n1347), .B(n1348), .ZN(n1149) );
XOR2_X1 U1039 ( .A(n1314), .B(n1298), .Z(n1348) );
XOR2_X1 U1040 ( .A(n1267), .B(n1289), .Z(n1298) );
XNOR2_X1 U1041 ( .A(G122), .B(KEYINPUT22), .ZN(n1289) );
INV_X1 U1042 ( .A(G116), .ZN(n1267) );
XOR2_X1 U1043 ( .A(G110), .B(n1335), .Z(n1314) );
INV_X1 U1044 ( .A(n1332), .ZN(n1335) );
XNOR2_X1 U1045 ( .A(G119), .B(KEYINPUT24), .ZN(n1332) );
XOR2_X1 U1046 ( .A(n1349), .B(n1350), .Z(n1347) );
XNOR2_X1 U1047 ( .A(G113), .B(n1351), .ZN(n1350) );
NAND2_X1 U1048 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
NAND2_X1 U1049 ( .A1(G104), .A2(n1354), .ZN(n1353) );
XOR2_X1 U1050 ( .A(KEYINPUT52), .B(n1355), .Z(n1352) );
NOR2_X1 U1051 ( .A1(G104), .A2(n1354), .ZN(n1355) );
INV_X1 U1052 ( .A(G107), .ZN(n1354) );
NAND2_X1 U1053 ( .A1(KEYINPUT30), .A2(G101), .ZN(n1349) );
XOR2_X1 U1054 ( .A(n1340), .B(n1356), .Z(n1233) );
XOR2_X1 U1055 ( .A(G125), .B(n1357), .Z(n1356) );
NOR2_X1 U1056 ( .A1(G953), .A2(n1144), .ZN(n1357) );
INV_X1 U1057 ( .A(G224), .ZN(n1144) );
XOR2_X1 U1058 ( .A(n1358), .B(n1359), .Z(n1340) );
XOR2_X1 U1059 ( .A(KEYINPUT40), .B(n1360), .Z(n1359) );
INV_X1 U1060 ( .A(n1248), .ZN(n1343) );
XNOR2_X1 U1061 ( .A(n1069), .B(KEYINPUT56), .ZN(n1248) );
NAND2_X1 U1062 ( .A1(G214), .A2(n1345), .ZN(n1069) );
NAND2_X1 U1063 ( .A1(n1361), .A2(n1276), .ZN(n1345) );
INV_X1 U1064 ( .A(G237), .ZN(n1361) );
NOR2_X1 U1065 ( .A1(n1102), .A2(n1101), .ZN(n1103) );
INV_X1 U1066 ( .A(n1067), .ZN(n1101) );
NAND2_X1 U1067 ( .A1(G221), .A2(n1156), .ZN(n1067) );
NAND2_X1 U1068 ( .A1(n1362), .A2(n1276), .ZN(n1156) );
XOR2_X1 U1069 ( .A(KEYINPUT33), .B(G234), .Z(n1362) );
XOR2_X1 U1070 ( .A(n1363), .B(n1080), .Z(n1102) );
NAND2_X1 U1071 ( .A1(n1364), .A2(n1276), .ZN(n1080) );
INV_X1 U1072 ( .A(G902), .ZN(n1276) );
XOR2_X1 U1073 ( .A(n1365), .B(n1366), .Z(n1364) );
XNOR2_X1 U1074 ( .A(n1190), .B(n1192), .ZN(n1366) );
XOR2_X1 U1075 ( .A(n1137), .B(KEYINPUT60), .Z(n1192) );
XOR2_X1 U1076 ( .A(n1360), .B(n1367), .Z(n1137) );
NOR2_X1 U1077 ( .A1(KEYINPUT61), .A2(n1358), .ZN(n1367) );
XNOR2_X1 U1078 ( .A(G128), .B(KEYINPUT36), .ZN(n1358) );
XOR2_X1 U1079 ( .A(G146), .B(G143), .Z(n1360) );
XNOR2_X1 U1080 ( .A(n1368), .B(n1369), .ZN(n1190) );
XOR2_X1 U1081 ( .A(KEYINPUT29), .B(G107), .Z(n1369) );
XOR2_X1 U1082 ( .A(n1370), .B(G101), .Z(n1368) );
NAND2_X1 U1083 ( .A1(KEYINPUT26), .A2(G104), .ZN(n1370) );
XOR2_X1 U1084 ( .A(n1371), .B(n1372), .Z(n1365) );
INV_X1 U1085 ( .A(n1191), .ZN(n1372) );
XOR2_X1 U1086 ( .A(n1373), .B(n1374), .Z(n1191) );
NOR2_X1 U1087 ( .A1(n1375), .A2(n1376), .ZN(n1374) );
XOR2_X1 U1088 ( .A(KEYINPUT31), .B(G953), .Z(n1376) );
INV_X1 U1089 ( .A(G227), .ZN(n1375) );
XOR2_X1 U1090 ( .A(G110), .B(n1133), .Z(n1373) );
INV_X1 U1091 ( .A(G140), .ZN(n1133) );
NAND2_X1 U1092 ( .A1(KEYINPUT17), .A2(n1341), .ZN(n1371) );
INV_X1 U1093 ( .A(n1185), .ZN(n1341) );
XOR2_X1 U1094 ( .A(n1377), .B(n1378), .Z(n1185) );
XOR2_X1 U1095 ( .A(KEYINPUT49), .B(G137), .Z(n1378) );
XOR2_X1 U1096 ( .A(n1139), .B(G134), .Z(n1377) );
INV_X1 U1097 ( .A(G131), .ZN(n1139) );
NAND2_X1 U1098 ( .A1(KEYINPUT18), .A2(n1189), .ZN(n1363) );
INV_X1 U1099 ( .A(G469), .ZN(n1189) );
endmodule


