//Key = 0110010000011111000010100001111101000111010010111000110110001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389;

NAND2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(G9) );
OR2_X1 U761 ( .A1(n1058), .A2(G107), .ZN(n1057) );
XOR2_X1 U762 ( .A(n1059), .B(KEYINPUT9), .Z(n1056) );
NAND2_X1 U763 ( .A1(G107), .A2(n1058), .ZN(n1059) );
NOR2_X1 U764 ( .A1(n1060), .A2(n1061), .ZN(G75) );
NOR4_X1 U765 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1061) );
NAND3_X1 U766 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1062) );
NAND2_X1 U767 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U768 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U769 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
NAND2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NAND3_X1 U771 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
XNOR2_X1 U772 ( .A(n1081), .B(KEYINPUT38), .ZN(n1080) );
NAND2_X1 U773 ( .A1(n1082), .A2(n1083), .ZN(n1076) );
NAND2_X1 U774 ( .A1(n1081), .A2(n1084), .ZN(n1071) );
NAND2_X1 U775 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U776 ( .A1(n1075), .A2(n1087), .ZN(n1086) );
NAND2_X1 U777 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U778 ( .A1(n1090), .A2(n1091), .A3(KEYINPUT49), .ZN(n1089) );
NAND2_X1 U779 ( .A1(n1073), .A2(n1092), .ZN(n1088) );
NAND2_X1 U780 ( .A1(n1082), .A2(n1091), .ZN(n1085) );
NAND4_X1 U781 ( .A1(n1082), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1091) );
NAND3_X1 U782 ( .A1(n1096), .A2(n1073), .A3(n1097), .ZN(n1094) );
NAND2_X1 U783 ( .A1(n1075), .A2(n1098), .ZN(n1093) );
NAND2_X1 U784 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U785 ( .A1(n1090), .A2(n1101), .ZN(n1100) );
INV_X1 U786 ( .A(KEYINPUT49), .ZN(n1101) );
NAND2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1099) );
INV_X1 U788 ( .A(n1104), .ZN(n1069) );
AND3_X1 U789 ( .A1(n1066), .A2(n1067), .A3(n1105), .ZN(n1060) );
NAND4_X1 U790 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1066) );
NOR2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U792 ( .A(n1078), .B(KEYINPUT12), .Z(n1111) );
XOR2_X1 U793 ( .A(n1112), .B(KEYINPUT26), .Z(n1110) );
NAND4_X1 U794 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1112) );
XNOR2_X1 U795 ( .A(n1117), .B(n1118), .ZN(n1114) );
XNOR2_X1 U796 ( .A(G475), .B(n1119), .ZN(n1113) );
XOR2_X1 U797 ( .A(n1120), .B(n1121), .Z(n1108) );
NAND2_X1 U798 ( .A1(KEYINPUT27), .A2(n1122), .ZN(n1121) );
XOR2_X1 U799 ( .A(n1123), .B(n1124), .Z(G72) );
XOR2_X1 U800 ( .A(n1125), .B(n1126), .Z(n1124) );
AND2_X1 U801 ( .A1(n1064), .A2(n1067), .ZN(n1126) );
NOR2_X1 U802 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
XOR2_X1 U803 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U804 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U805 ( .A(n1133), .B(n1134), .ZN(n1129) );
INV_X1 U806 ( .A(G128), .ZN(n1134) );
NAND2_X1 U807 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
OR2_X1 U808 ( .A1(n1137), .A2(G131), .ZN(n1136) );
XOR2_X1 U809 ( .A(n1138), .B(KEYINPUT35), .Z(n1135) );
NAND2_X1 U810 ( .A1(G131), .A2(n1137), .ZN(n1138) );
XOR2_X1 U811 ( .A(G134), .B(G137), .Z(n1137) );
NOR2_X1 U812 ( .A1(G900), .A2(n1139), .ZN(n1127) );
XNOR2_X1 U813 ( .A(G953), .B(KEYINPUT10), .ZN(n1139) );
NOR3_X1 U814 ( .A1(n1067), .A2(KEYINPUT54), .A3(n1140), .ZN(n1123) );
AND2_X1 U815 ( .A1(G227), .A2(G900), .ZN(n1140) );
NAND2_X1 U816 ( .A1(n1141), .A2(n1142), .ZN(G69) );
NAND2_X1 U817 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
OR2_X1 U818 ( .A1(n1067), .A2(G224), .ZN(n1144) );
NAND3_X1 U819 ( .A1(G953), .A2(n1145), .A3(n1146), .ZN(n1141) );
INV_X1 U820 ( .A(n1143), .ZN(n1146) );
XNOR2_X1 U821 ( .A(n1147), .B(n1148), .ZN(n1143) );
NOR2_X1 U822 ( .A1(n1149), .A2(G953), .ZN(n1148) );
NOR2_X1 U823 ( .A1(n1150), .A2(n1063), .ZN(n1149) );
NAND3_X1 U824 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1147) );
NAND2_X1 U825 ( .A1(G953), .A2(n1154), .ZN(n1153) );
OR2_X1 U826 ( .A1(n1155), .A2(n1156), .ZN(n1152) );
NAND2_X1 U827 ( .A1(n1155), .A2(n1157), .ZN(n1151) );
XNOR2_X1 U828 ( .A(n1156), .B(KEYINPUT22), .ZN(n1157) );
NAND2_X1 U829 ( .A1(G898), .A2(G224), .ZN(n1145) );
NOR2_X1 U830 ( .A1(n1158), .A2(n1159), .ZN(G66) );
XNOR2_X1 U831 ( .A(n1160), .B(n1161), .ZN(n1159) );
NOR2_X1 U832 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NOR2_X1 U833 ( .A1(n1158), .A2(n1164), .ZN(G63) );
XOR2_X1 U834 ( .A(n1165), .B(n1166), .Z(n1164) );
XNOR2_X1 U835 ( .A(KEYINPUT61), .B(n1167), .ZN(n1166) );
NAND3_X1 U836 ( .A1(n1168), .A2(G478), .A3(KEYINPUT55), .ZN(n1165) );
NOR2_X1 U837 ( .A1(n1158), .A2(n1169), .ZN(G60) );
XOR2_X1 U838 ( .A(n1170), .B(n1171), .Z(n1169) );
AND2_X1 U839 ( .A1(G475), .A2(n1168), .ZN(n1171) );
NAND2_X1 U840 ( .A1(KEYINPUT29), .A2(n1172), .ZN(n1170) );
XNOR2_X1 U841 ( .A(G104), .B(n1173), .ZN(G6) );
NOR2_X1 U842 ( .A1(n1158), .A2(n1174), .ZN(G57) );
XNOR2_X1 U843 ( .A(n1175), .B(n1176), .ZN(n1174) );
XOR2_X1 U844 ( .A(KEYINPUT57), .B(n1177), .Z(n1176) );
AND2_X1 U845 ( .A1(G472), .A2(n1168), .ZN(n1177) );
INV_X1 U846 ( .A(n1163), .ZN(n1168) );
NOR2_X1 U847 ( .A1(n1158), .A2(n1178), .ZN(G54) );
NOR2_X1 U848 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XOR2_X1 U849 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U850 ( .A1(n1183), .A2(KEYINPUT40), .ZN(n1182) );
NOR2_X1 U851 ( .A1(n1122), .A2(n1163), .ZN(n1181) );
AND2_X1 U852 ( .A1(n1183), .A2(KEYINPUT40), .ZN(n1179) );
AND2_X1 U853 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NAND2_X1 U854 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
INV_X1 U855 ( .A(n1188), .ZN(n1187) );
XNOR2_X1 U856 ( .A(n1189), .B(n1190), .ZN(n1186) );
XOR2_X1 U857 ( .A(n1191), .B(KEYINPUT42), .Z(n1184) );
NAND2_X1 U858 ( .A1(n1192), .A2(n1188), .ZN(n1191) );
XNOR2_X1 U859 ( .A(n1193), .B(n1194), .ZN(n1188) );
NOR2_X1 U860 ( .A1(G140), .A2(KEYINPUT36), .ZN(n1194) );
XNOR2_X1 U861 ( .A(n1195), .B(n1196), .ZN(n1193) );
XNOR2_X1 U862 ( .A(n1197), .B(n1190), .ZN(n1192) );
XNOR2_X1 U863 ( .A(n1198), .B(n1199), .ZN(n1190) );
NAND2_X1 U864 ( .A1(KEYINPUT39), .A2(n1200), .ZN(n1198) );
NOR2_X1 U865 ( .A1(n1158), .A2(n1201), .ZN(G51) );
XOR2_X1 U866 ( .A(n1202), .B(n1203), .Z(n1201) );
XOR2_X1 U867 ( .A(n1204), .B(n1205), .Z(n1203) );
NOR2_X1 U868 ( .A1(n1206), .A2(n1163), .ZN(n1204) );
NAND2_X1 U869 ( .A1(G902), .A2(n1207), .ZN(n1163) );
OR3_X1 U870 ( .A1(n1065), .A2(n1064), .A3(n1063), .ZN(n1207) );
NAND3_X1 U871 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1063) );
NAND2_X1 U872 ( .A1(n1211), .A2(n1083), .ZN(n1210) );
OR2_X1 U873 ( .A1(n1212), .A2(n1213), .ZN(n1083) );
NAND2_X1 U874 ( .A1(n1214), .A2(n1215), .ZN(n1064) );
NOR4_X1 U875 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1215) );
INV_X1 U876 ( .A(n1220), .ZN(n1216) );
AND4_X1 U877 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1214) );
XNOR2_X1 U878 ( .A(n1150), .B(KEYINPUT2), .ZN(n1065) );
NAND4_X1 U879 ( .A1(n1225), .A2(n1173), .A3(n1226), .A4(n1058), .ZN(n1150) );
NAND3_X1 U880 ( .A1(n1213), .A2(n1227), .A3(n1228), .ZN(n1058) );
NAND3_X1 U881 ( .A1(n1228), .A2(n1227), .A3(n1212), .ZN(n1173) );
INV_X1 U882 ( .A(n1095), .ZN(n1227) );
NAND2_X1 U883 ( .A1(n1229), .A2(n1073), .ZN(n1095) );
NOR2_X1 U884 ( .A1(n1230), .A2(n1103), .ZN(n1073) );
NAND2_X1 U885 ( .A1(n1231), .A2(n1232), .ZN(n1225) );
XOR2_X1 U886 ( .A(KEYINPUT34), .B(n1090), .Z(n1232) );
AND2_X1 U887 ( .A1(n1233), .A2(n1105), .ZN(n1158) );
INV_X1 U888 ( .A(G952), .ZN(n1105) );
XNOR2_X1 U889 ( .A(G953), .B(KEYINPUT15), .ZN(n1233) );
XNOR2_X1 U890 ( .A(G146), .B(n1222), .ZN(G48) );
NAND2_X1 U891 ( .A1(n1212), .A2(n1234), .ZN(n1222) );
XNOR2_X1 U892 ( .A(G143), .B(n1224), .ZN(G45) );
NAND3_X1 U893 ( .A1(n1235), .A2(n1092), .A3(n1236), .ZN(n1224) );
XOR2_X1 U894 ( .A(n1221), .B(n1237), .Z(G42) );
NAND2_X1 U895 ( .A1(KEYINPUT28), .A2(G140), .ZN(n1237) );
NAND3_X1 U896 ( .A1(n1090), .A2(n1212), .A3(n1238), .ZN(n1221) );
AND3_X1 U897 ( .A1(n1082), .A2(n1239), .A3(n1229), .ZN(n1238) );
XOR2_X1 U898 ( .A(G137), .B(n1219), .Z(G39) );
AND4_X1 U899 ( .A1(n1082), .A2(n1236), .A3(n1081), .A4(n1240), .ZN(n1219) );
XOR2_X1 U900 ( .A(n1218), .B(n1241), .Z(G36) );
NOR2_X1 U901 ( .A1(KEYINPUT19), .A2(n1242), .ZN(n1241) );
AND2_X1 U902 ( .A1(n1243), .A2(n1213), .ZN(n1218) );
XOR2_X1 U903 ( .A(G131), .B(n1217), .Z(G33) );
AND2_X1 U904 ( .A1(n1212), .A2(n1243), .ZN(n1217) );
AND3_X1 U905 ( .A1(n1236), .A2(n1102), .A3(n1082), .ZN(n1243) );
AND2_X1 U906 ( .A1(n1078), .A2(n1107), .ZN(n1082) );
XNOR2_X1 U907 ( .A(G128), .B(n1220), .ZN(G30) );
NAND2_X1 U908 ( .A1(n1234), .A2(n1213), .ZN(n1220) );
AND3_X1 U909 ( .A1(n1092), .A2(n1240), .A3(n1236), .ZN(n1234) );
AND3_X1 U910 ( .A1(n1103), .A2(n1239), .A3(n1229), .ZN(n1236) );
NAND2_X1 U911 ( .A1(n1244), .A2(n1245), .ZN(G3) );
NAND2_X1 U912 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XOR2_X1 U913 ( .A(KEYINPUT53), .B(n1248), .Z(n1244) );
NOR2_X1 U914 ( .A1(n1246), .A2(n1247), .ZN(n1248) );
INV_X1 U915 ( .A(n1226), .ZN(n1246) );
NAND3_X1 U916 ( .A1(n1102), .A2(n1103), .A3(n1231), .ZN(n1226) );
XNOR2_X1 U917 ( .A(G125), .B(n1223), .ZN(G27) );
NAND3_X1 U918 ( .A1(n1090), .A2(n1212), .A3(n1249), .ZN(n1223) );
AND3_X1 U919 ( .A1(n1075), .A2(n1239), .A3(n1092), .ZN(n1249) );
NAND2_X1 U920 ( .A1(n1104), .A2(n1250), .ZN(n1239) );
NAND4_X1 U921 ( .A1(n1251), .A2(G902), .A3(n1252), .A4(n1253), .ZN(n1250) );
INV_X1 U922 ( .A(G900), .ZN(n1253) );
XNOR2_X1 U923 ( .A(G953), .B(KEYINPUT5), .ZN(n1251) );
XNOR2_X1 U924 ( .A(G122), .B(n1208), .ZN(G24) );
NAND4_X1 U925 ( .A1(n1235), .A2(n1075), .A3(n1116), .A4(n1228), .ZN(n1208) );
AND3_X1 U926 ( .A1(n1254), .A2(n1255), .A3(n1102), .ZN(n1235) );
XNOR2_X1 U927 ( .A(G119), .B(n1209), .ZN(G21) );
NAND3_X1 U928 ( .A1(n1256), .A2(n1240), .A3(n1081), .ZN(n1209) );
XOR2_X1 U929 ( .A(n1257), .B(n1258), .Z(G18) );
XNOR2_X1 U930 ( .A(G116), .B(KEYINPUT32), .ZN(n1258) );
NAND2_X1 U931 ( .A1(n1259), .A2(n1211), .ZN(n1257) );
XNOR2_X1 U932 ( .A(n1213), .B(KEYINPUT52), .ZN(n1259) );
NOR2_X1 U933 ( .A1(n1255), .A2(n1115), .ZN(n1213) );
XNOR2_X1 U934 ( .A(G113), .B(n1260), .ZN(G15) );
NAND2_X1 U935 ( .A1(n1212), .A2(n1211), .ZN(n1260) );
AND2_X1 U936 ( .A1(n1256), .A2(n1102), .ZN(n1211) );
INV_X1 U937 ( .A(n1230), .ZN(n1102) );
AND3_X1 U938 ( .A1(n1228), .A2(n1103), .A3(n1075), .ZN(n1256) );
AND2_X1 U939 ( .A1(n1096), .A2(n1106), .ZN(n1075) );
AND2_X1 U940 ( .A1(n1115), .A2(n1255), .ZN(n1212) );
INV_X1 U941 ( .A(n1254), .ZN(n1115) );
XNOR2_X1 U942 ( .A(G110), .B(n1261), .ZN(G12) );
NAND2_X1 U943 ( .A1(n1231), .A2(n1090), .ZN(n1261) );
AND2_X1 U944 ( .A1(n1116), .A2(n1240), .ZN(n1090) );
XNOR2_X1 U945 ( .A(n1230), .B(KEYINPUT46), .ZN(n1240) );
NAND3_X1 U946 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1230) );
NAND2_X1 U947 ( .A1(n1265), .A2(n1162), .ZN(n1264) );
NAND2_X1 U948 ( .A1(KEYINPUT18), .A2(n1266), .ZN(n1263) );
NAND2_X1 U949 ( .A1(n1117), .A2(n1267), .ZN(n1266) );
XNOR2_X1 U950 ( .A(KEYINPUT37), .B(n1268), .ZN(n1267) );
NAND2_X1 U951 ( .A1(n1269), .A2(n1270), .ZN(n1262) );
INV_X1 U952 ( .A(KEYINPUT18), .ZN(n1270) );
NAND2_X1 U953 ( .A1(n1271), .A2(n1272), .ZN(n1269) );
NAND3_X1 U954 ( .A1(KEYINPUT37), .A2(n1117), .A3(n1268), .ZN(n1272) );
INV_X1 U955 ( .A(n1162), .ZN(n1117) );
NAND2_X1 U956 ( .A1(G217), .A2(n1273), .ZN(n1162) );
OR2_X1 U957 ( .A1(n1268), .A2(KEYINPUT37), .ZN(n1271) );
INV_X1 U958 ( .A(n1265), .ZN(n1268) );
XOR2_X1 U959 ( .A(n1118), .B(KEYINPUT7), .Z(n1265) );
AND2_X1 U960 ( .A1(n1274), .A2(n1160), .ZN(n1118) );
XNOR2_X1 U961 ( .A(n1275), .B(n1276), .ZN(n1160) );
XOR2_X1 U962 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U963 ( .A(n1279), .B(n1280), .Z(n1278) );
AND3_X1 U964 ( .A1(G221), .A2(n1067), .A3(n1281), .ZN(n1280) );
NAND2_X1 U965 ( .A1(n1282), .A2(KEYINPUT14), .ZN(n1279) );
XNOR2_X1 U966 ( .A(G137), .B(KEYINPUT21), .ZN(n1282) );
NAND2_X1 U967 ( .A1(n1283), .A2(n1284), .ZN(n1277) );
NAND2_X1 U968 ( .A1(n1285), .A2(n1196), .ZN(n1284) );
XOR2_X1 U969 ( .A(n1286), .B(KEYINPUT6), .Z(n1283) );
OR2_X1 U970 ( .A1(n1285), .A2(n1196), .ZN(n1286) );
XOR2_X1 U971 ( .A(G128), .B(n1287), .Z(n1285) );
NOR2_X1 U972 ( .A1(KEYINPUT45), .A2(n1288), .ZN(n1287) );
XOR2_X1 U973 ( .A(n1289), .B(n1290), .Z(n1275) );
NAND2_X1 U974 ( .A1(KEYINPUT48), .A2(n1291), .ZN(n1289) );
INV_X1 U975 ( .A(G146), .ZN(n1291) );
XNOR2_X1 U976 ( .A(G902), .B(KEYINPUT17), .ZN(n1274) );
INV_X1 U977 ( .A(n1103), .ZN(n1116) );
XNOR2_X1 U978 ( .A(n1292), .B(G472), .ZN(n1103) );
NAND2_X1 U979 ( .A1(n1175), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U980 ( .A(n1294), .B(n1295), .ZN(n1175) );
XOR2_X1 U981 ( .A(n1296), .B(n1297), .Z(n1295) );
XNOR2_X1 U982 ( .A(n1298), .B(G113), .ZN(n1297) );
XOR2_X1 U983 ( .A(n1299), .B(n1300), .Z(n1294) );
XNOR2_X1 U984 ( .A(n1301), .B(n1288), .ZN(n1300) );
NAND2_X1 U985 ( .A1(n1302), .A2(G210), .ZN(n1301) );
AND3_X1 U986 ( .A1(n1228), .A2(n1229), .A3(n1081), .ZN(n1231) );
NOR2_X1 U987 ( .A1(n1254), .A2(n1255), .ZN(n1081) );
NAND2_X1 U988 ( .A1(n1303), .A2(n1304), .ZN(n1255) );
NAND2_X1 U989 ( .A1(n1305), .A2(n1119), .ZN(n1304) );
XOR2_X1 U990 ( .A(KEYINPUT41), .B(n1306), .Z(n1303) );
NOR2_X1 U991 ( .A1(n1119), .A2(n1305), .ZN(n1306) );
XNOR2_X1 U992 ( .A(KEYINPUT62), .B(G475), .ZN(n1305) );
AND2_X1 U993 ( .A1(n1172), .A2(n1293), .ZN(n1119) );
XNOR2_X1 U994 ( .A(n1307), .B(n1308), .ZN(n1172) );
XOR2_X1 U995 ( .A(n1309), .B(n1310), .Z(n1308) );
NAND2_X1 U996 ( .A1(KEYINPUT33), .A2(n1311), .ZN(n1310) );
NAND3_X1 U997 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(n1309) );
NAND2_X1 U998 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
INV_X1 U999 ( .A(KEYINPUT13), .ZN(n1316) );
NAND3_X1 U1000 ( .A1(KEYINPUT13), .A2(n1317), .A3(n1318), .ZN(n1313) );
OR2_X1 U1001 ( .A1(n1318), .A2(n1317), .ZN(n1312) );
NOR2_X1 U1002 ( .A1(n1319), .A2(n1315), .ZN(n1317) );
XOR2_X1 U1003 ( .A(G146), .B(n1290), .Z(n1315) );
XNOR2_X1 U1004 ( .A(n1131), .B(KEYINPUT43), .ZN(n1290) );
XNOR2_X1 U1005 ( .A(G125), .B(G140), .ZN(n1131) );
XOR2_X1 U1006 ( .A(KEYINPUT44), .B(KEYINPUT11), .Z(n1319) );
XOR2_X1 U1007 ( .A(n1320), .B(n1321), .Z(n1318) );
XNOR2_X1 U1008 ( .A(G131), .B(n1322), .ZN(n1321) );
NAND2_X1 U1009 ( .A1(n1302), .A2(G214), .ZN(n1322) );
NOR2_X1 U1010 ( .A1(G953), .A2(G237), .ZN(n1302) );
NAND2_X1 U1011 ( .A1(KEYINPUT20), .A2(n1323), .ZN(n1320) );
XNOR2_X1 U1012 ( .A(G104), .B(n1324), .ZN(n1307) );
XNOR2_X1 U1013 ( .A(KEYINPUT3), .B(n1325), .ZN(n1324) );
XNOR2_X1 U1014 ( .A(n1326), .B(G478), .ZN(n1254) );
NAND2_X1 U1015 ( .A1(n1293), .A2(n1167), .ZN(n1326) );
NAND3_X1 U1016 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1167) );
NAND2_X1 U1017 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
NAND2_X1 U1018 ( .A1(KEYINPUT63), .A2(n1332), .ZN(n1331) );
XOR2_X1 U1019 ( .A(KEYINPUT16), .B(n1333), .Z(n1332) );
NAND3_X1 U1020 ( .A1(KEYINPUT63), .A2(n1334), .A3(n1333), .ZN(n1328) );
INV_X1 U1021 ( .A(n1330), .ZN(n1334) );
XNOR2_X1 U1022 ( .A(n1335), .B(n1336), .ZN(n1330) );
XOR2_X1 U1023 ( .A(n1337), .B(n1338), .Z(n1336) );
XNOR2_X1 U1024 ( .A(n1298), .B(G107), .ZN(n1338) );
NOR2_X1 U1025 ( .A1(KEYINPUT8), .A2(n1323), .ZN(n1337) );
XNOR2_X1 U1026 ( .A(G122), .B(n1339), .ZN(n1335) );
XNOR2_X1 U1027 ( .A(n1242), .B(G128), .ZN(n1339) );
INV_X1 U1028 ( .A(G134), .ZN(n1242) );
OR2_X1 U1029 ( .A1(n1333), .A2(KEYINPUT63), .ZN(n1327) );
AND3_X1 U1030 ( .A1(n1281), .A2(n1067), .A3(n1340), .ZN(n1333) );
XNOR2_X1 U1031 ( .A(G217), .B(KEYINPUT60), .ZN(n1340) );
XOR2_X1 U1032 ( .A(G234), .B(KEYINPUT0), .Z(n1281) );
NOR2_X1 U1033 ( .A1(n1096), .A2(n1097), .ZN(n1229) );
INV_X1 U1034 ( .A(n1106), .ZN(n1097) );
NAND2_X1 U1035 ( .A1(G221), .A2(n1273), .ZN(n1106) );
NAND2_X1 U1036 ( .A1(G234), .A2(n1293), .ZN(n1273) );
XNOR2_X1 U1037 ( .A(n1120), .B(n1122), .ZN(n1096) );
INV_X1 U1038 ( .A(G469), .ZN(n1122) );
NAND2_X1 U1039 ( .A1(n1293), .A2(n1341), .ZN(n1120) );
NAND2_X1 U1040 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NAND2_X1 U1041 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
XOR2_X1 U1042 ( .A(n1346), .B(n1347), .Z(n1345) );
NOR2_X1 U1043 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
XOR2_X1 U1044 ( .A(n1195), .B(KEYINPUT56), .Z(n1348) );
XNOR2_X1 U1045 ( .A(G140), .B(n1196), .ZN(n1344) );
INV_X1 U1046 ( .A(G110), .ZN(n1196) );
NAND2_X1 U1047 ( .A1(n1350), .A2(n1351), .ZN(n1342) );
XOR2_X1 U1048 ( .A(n1346), .B(n1352), .Z(n1351) );
NOR2_X1 U1049 ( .A1(n1195), .A2(n1349), .ZN(n1352) );
INV_X1 U1050 ( .A(KEYINPUT1), .ZN(n1349) );
NAND2_X1 U1051 ( .A1(n1353), .A2(n1067), .ZN(n1195) );
XOR2_X1 U1052 ( .A(KEYINPUT24), .B(G227), .Z(n1353) );
XNOR2_X1 U1053 ( .A(n1299), .B(n1189), .ZN(n1346) );
INV_X1 U1054 ( .A(n1197), .ZN(n1189) );
XOR2_X1 U1055 ( .A(G128), .B(n1354), .Z(n1197) );
NOR2_X1 U1056 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
NOR3_X1 U1057 ( .A1(n1357), .A2(G107), .A3(n1358), .ZN(n1356) );
INV_X1 U1058 ( .A(KEYINPUT50), .ZN(n1357) );
NOR2_X1 U1059 ( .A1(KEYINPUT50), .A2(n1359), .ZN(n1355) );
XNOR2_X1 U1060 ( .A(n1199), .B(n1200), .ZN(n1299) );
XNOR2_X1 U1061 ( .A(n1360), .B(n1361), .ZN(n1200) );
NOR2_X1 U1062 ( .A1(KEYINPUT51), .A2(G134), .ZN(n1361) );
XNOR2_X1 U1063 ( .A(G131), .B(G137), .ZN(n1360) );
XOR2_X1 U1064 ( .A(G101), .B(n1132), .Z(n1199) );
XNOR2_X1 U1065 ( .A(G140), .B(G110), .ZN(n1350) );
AND2_X1 U1066 ( .A1(n1092), .A2(n1362), .ZN(n1228) );
NAND2_X1 U1067 ( .A1(n1363), .A2(n1104), .ZN(n1362) );
NAND3_X1 U1068 ( .A1(n1252), .A2(n1067), .A3(G952), .ZN(n1104) );
XOR2_X1 U1069 ( .A(KEYINPUT31), .B(n1364), .Z(n1363) );
AND4_X1 U1070 ( .A1(n1154), .A2(n1252), .A3(G902), .A4(G953), .ZN(n1364) );
NAND2_X1 U1071 ( .A1(G237), .A2(G234), .ZN(n1252) );
INV_X1 U1072 ( .A(G898), .ZN(n1154) );
NOR2_X1 U1073 ( .A1(n1078), .A2(n1079), .ZN(n1092) );
INV_X1 U1074 ( .A(n1107), .ZN(n1079) );
NAND2_X1 U1075 ( .A1(G214), .A2(n1365), .ZN(n1107) );
XNOR2_X1 U1076 ( .A(n1366), .B(n1206), .ZN(n1078) );
NAND2_X1 U1077 ( .A1(G210), .A2(n1365), .ZN(n1206) );
NAND2_X1 U1078 ( .A1(n1367), .A2(n1293), .ZN(n1365) );
INV_X1 U1079 ( .A(G237), .ZN(n1367) );
NAND2_X1 U1080 ( .A1(n1368), .A2(n1293), .ZN(n1366) );
INV_X1 U1081 ( .A(G902), .ZN(n1293) );
XOR2_X1 U1082 ( .A(n1369), .B(n1205), .Z(n1368) );
XOR2_X1 U1083 ( .A(n1155), .B(n1156), .Z(n1205) );
XNOR2_X1 U1084 ( .A(n1370), .B(n1371), .ZN(n1156) );
XNOR2_X1 U1085 ( .A(n1311), .B(G110), .ZN(n1371) );
INV_X1 U1086 ( .A(G122), .ZN(n1311) );
NAND3_X1 U1087 ( .A1(n1372), .A2(n1373), .A3(n1374), .ZN(n1370) );
NAND2_X1 U1088 ( .A1(G113), .A2(n1375), .ZN(n1374) );
NAND2_X1 U1089 ( .A1(n1376), .A2(n1377), .ZN(n1375) );
XNOR2_X1 U1090 ( .A(KEYINPUT30), .B(n1378), .ZN(n1376) );
NAND3_X1 U1091 ( .A1(n1378), .A2(n1379), .A3(n1380), .ZN(n1373) );
INV_X1 U1092 ( .A(KEYINPUT58), .ZN(n1380) );
NAND2_X1 U1093 ( .A1(KEYINPUT30), .A2(n1381), .ZN(n1379) );
INV_X1 U1094 ( .A(n1382), .ZN(n1378) );
NAND3_X1 U1095 ( .A1(n1382), .A2(n1383), .A3(KEYINPUT58), .ZN(n1372) );
NAND2_X1 U1096 ( .A1(n1384), .A2(n1381), .ZN(n1383) );
NAND2_X1 U1097 ( .A1(n1325), .A2(n1377), .ZN(n1381) );
INV_X1 U1098 ( .A(KEYINPUT4), .ZN(n1377) );
INV_X1 U1099 ( .A(G113), .ZN(n1325) );
INV_X1 U1100 ( .A(KEYINPUT30), .ZN(n1384) );
XNOR2_X1 U1101 ( .A(n1385), .B(n1288), .ZN(n1382) );
XOR2_X1 U1102 ( .A(G119), .B(KEYINPUT59), .Z(n1288) );
NAND2_X1 U1103 ( .A1(KEYINPUT47), .A2(n1298), .ZN(n1385) );
INV_X1 U1104 ( .A(G116), .ZN(n1298) );
XNOR2_X1 U1105 ( .A(n1247), .B(n1359), .ZN(n1155) );
XNOR2_X1 U1106 ( .A(n1358), .B(G107), .ZN(n1359) );
INV_X1 U1107 ( .A(G104), .ZN(n1358) );
INV_X1 U1108 ( .A(G101), .ZN(n1247) );
NOR2_X1 U1109 ( .A1(KEYINPUT25), .A2(n1202), .ZN(n1369) );
XOR2_X1 U1110 ( .A(n1386), .B(n1387), .Z(n1202) );
XNOR2_X1 U1111 ( .A(n1388), .B(n1296), .ZN(n1387) );
NOR2_X1 U1112 ( .A1(KEYINPUT23), .A2(G128), .ZN(n1296) );
INV_X1 U1113 ( .A(G125), .ZN(n1388) );
XOR2_X1 U1114 ( .A(n1389), .B(n1132), .Z(n1386) );
XNOR2_X1 U1115 ( .A(n1323), .B(G146), .ZN(n1132) );
INV_X1 U1116 ( .A(G143), .ZN(n1323) );
NAND2_X1 U1117 ( .A1(G224), .A2(n1067), .ZN(n1389) );
INV_X1 U1118 ( .A(G953), .ZN(n1067) );
endmodule


