//Key = 0111010110110110010111111101010111110000011100010100100100111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;

XNOR2_X1 U744 ( .A(G107), .B(n1025), .ZN(G9) );
NOR2_X1 U745 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR3_X1 U746 ( .A1(n1028), .A2(G953), .A3(G952), .ZN(n1027) );
INV_X1 U747 ( .A(n1029), .ZN(n1028) );
NOR3_X1 U748 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1026) );
NOR2_X1 U749 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR3_X1 U750 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1033) );
NOR2_X1 U751 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR2_X1 U752 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U753 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR3_X1 U754 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1036) );
INV_X1 U755 ( .A(n1047), .ZN(n1046) );
NOR2_X1 U756 ( .A1(n1048), .A2(n1049), .ZN(n1045) );
AND2_X1 U757 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
AND3_X1 U758 ( .A1(KEYINPUT41), .A2(n1052), .A3(n1053), .ZN(n1048) );
NOR2_X1 U759 ( .A1(n1054), .A2(KEYINPUT41), .ZN(n1035) );
AND4_X1 U760 ( .A1(n1047), .A2(n1052), .A3(n1053), .A4(n1055), .ZN(n1054) );
NAND3_X1 U761 ( .A1(n1029), .A2(n1056), .A3(n1057), .ZN(n1030) );
NAND2_X1 U762 ( .A1(n1047), .A2(n1058), .ZN(n1057) );
NAND2_X1 U763 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND3_X1 U764 ( .A1(n1061), .A2(n1062), .A3(n1055), .ZN(n1060) );
NAND2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U766 ( .A1(n1065), .A2(n1066), .A3(n1053), .ZN(n1064) );
NAND2_X1 U767 ( .A1(n1067), .A2(n1050), .ZN(n1063) );
NAND2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1059) );
NAND3_X1 U769 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
INV_X1 U770 ( .A(n1073), .ZN(n1072) );
OR2_X1 U771 ( .A1(n1034), .A2(KEYINPUT23), .ZN(n1071) );
NAND3_X1 U772 ( .A1(n1074), .A2(n1075), .A3(KEYINPUT23), .ZN(n1070) );
INV_X1 U773 ( .A(n1039), .ZN(n1068) );
NAND3_X1 U774 ( .A1(n1053), .A2(n1050), .A3(n1055), .ZN(n1039) );
INV_X1 U775 ( .A(n1044), .ZN(n1055) );
NAND2_X1 U776 ( .A1(n1076), .A2(n1077), .ZN(n1029) );
NOR4_X1 U777 ( .A1(n1078), .A2(n1074), .A3(n1079), .A4(n1080), .ZN(n1077) );
XNOR2_X1 U778 ( .A(n1066), .B(KEYINPUT2), .ZN(n1079) );
INV_X1 U779 ( .A(n1042), .ZN(n1078) );
NOR4_X1 U780 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1076) );
XOR2_X1 U781 ( .A(G469), .B(n1085), .Z(n1084) );
NOR2_X1 U782 ( .A1(KEYINPUT46), .A2(n1086), .ZN(n1085) );
AND2_X1 U783 ( .A1(n1087), .A2(KEYINPUT16), .ZN(n1082) );
NOR2_X1 U784 ( .A1(KEYINPUT16), .A2(n1053), .ZN(n1081) );
XOR2_X1 U785 ( .A(n1088), .B(n1089), .Z(G72) );
XOR2_X1 U786 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND2_X1 U787 ( .A1(G953), .A2(n1092), .ZN(n1091) );
NAND2_X1 U788 ( .A1(G900), .A2(G227), .ZN(n1092) );
NAND2_X1 U789 ( .A1(n1093), .A2(n1094), .ZN(n1090) );
NAND2_X1 U790 ( .A1(G953), .A2(n1095), .ZN(n1094) );
XOR2_X1 U791 ( .A(n1096), .B(n1097), .Z(n1093) );
XOR2_X1 U792 ( .A(n1098), .B(n1099), .Z(n1097) );
XOR2_X1 U793 ( .A(G137), .B(G134), .Z(n1096) );
NOR2_X1 U794 ( .A1(n1100), .A2(G953), .ZN(n1088) );
XOR2_X1 U795 ( .A(n1101), .B(n1102), .Z(G69) );
NOR2_X1 U796 ( .A1(n1103), .A2(n1056), .ZN(n1102) );
AND2_X1 U797 ( .A1(G898), .A2(G224), .ZN(n1103) );
NAND2_X1 U798 ( .A1(n1104), .A2(n1105), .ZN(n1101) );
NAND2_X1 U799 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U800 ( .A(KEYINPUT34), .B(n1108), .Z(n1104) );
NOR2_X1 U801 ( .A1(n1106), .A2(n1107), .ZN(n1108) );
NAND2_X1 U802 ( .A1(n1056), .A2(n1109), .ZN(n1107) );
NAND2_X1 U803 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XNOR2_X1 U804 ( .A(n1112), .B(KEYINPUT43), .ZN(n1110) );
AND2_X1 U805 ( .A1(n1113), .A2(n1114), .ZN(n1106) );
XNOR2_X1 U806 ( .A(n1115), .B(n1116), .ZN(n1113) );
XOR2_X1 U807 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U808 ( .A1(n1119), .A2(n1120), .ZN(G66) );
XOR2_X1 U809 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U810 ( .A(n1123), .B(KEYINPUT4), .Z(n1121) );
NAND2_X1 U811 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NOR2_X1 U812 ( .A1(n1119), .A2(n1126), .ZN(G63) );
XOR2_X1 U813 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND2_X1 U814 ( .A1(n1124), .A2(G478), .ZN(n1127) );
NOR2_X1 U815 ( .A1(n1119), .A2(n1129), .ZN(G60) );
XOR2_X1 U816 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U817 ( .A1(n1124), .A2(G475), .ZN(n1130) );
XNOR2_X1 U818 ( .A(G104), .B(n1132), .ZN(G6) );
NOR2_X1 U819 ( .A1(n1119), .A2(n1133), .ZN(G57) );
XOR2_X1 U820 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U821 ( .A(n1136), .B(n1137), .ZN(n1135) );
NAND2_X1 U822 ( .A1(KEYINPUT22), .A2(n1138), .ZN(n1136) );
XOR2_X1 U823 ( .A(n1139), .B(n1140), .Z(n1134) );
NOR2_X1 U824 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XOR2_X1 U825 ( .A(n1143), .B(KEYINPUT11), .Z(n1142) );
NAND2_X1 U826 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NOR2_X1 U827 ( .A1(n1145), .A2(n1144), .ZN(n1141) );
NAND2_X1 U828 ( .A1(n1124), .A2(G472), .ZN(n1139) );
NOR2_X1 U829 ( .A1(n1119), .A2(n1146), .ZN(G54) );
XOR2_X1 U830 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U831 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U832 ( .A1(G110), .A2(KEYINPUT37), .ZN(n1149) );
XOR2_X1 U833 ( .A(n1151), .B(n1152), .Z(n1147) );
XOR2_X1 U834 ( .A(n1153), .B(G140), .Z(n1152) );
NAND2_X1 U835 ( .A1(n1124), .A2(G469), .ZN(n1153) );
NAND2_X1 U836 ( .A1(KEYINPUT59), .A2(n1154), .ZN(n1151) );
NOR2_X1 U837 ( .A1(n1119), .A2(n1155), .ZN(G51) );
XOR2_X1 U838 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U839 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U840 ( .A(KEYINPUT33), .B(G125), .Z(n1159) );
XOR2_X1 U841 ( .A(n1144), .B(n1160), .Z(n1156) );
XOR2_X1 U842 ( .A(n1161), .B(n1162), .Z(n1160) );
NAND2_X1 U843 ( .A1(KEYINPUT42), .A2(n1163), .ZN(n1162) );
NAND2_X1 U844 ( .A1(n1124), .A2(n1164), .ZN(n1161) );
AND2_X1 U845 ( .A1(G902), .A2(n1032), .ZN(n1124) );
NAND3_X1 U846 ( .A1(n1112), .A2(n1111), .A3(n1100), .ZN(n1032) );
AND2_X1 U847 ( .A1(n1165), .A2(n1166), .ZN(n1100) );
NOR4_X1 U848 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
AND4_X1 U849 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1165) );
AND4_X1 U850 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1111) );
NAND3_X1 U851 ( .A1(n1179), .A2(n1050), .A3(n1180), .ZN(n1175) );
AND4_X1 U852 ( .A1(n1132), .A2(n1181), .A3(n1182), .A4(n1025), .ZN(n1112) );
NAND3_X1 U853 ( .A1(n1067), .A2(n1050), .A3(n1183), .ZN(n1025) );
NAND3_X1 U854 ( .A1(n1183), .A2(n1050), .A3(n1051), .ZN(n1132) );
NOR2_X1 U855 ( .A1(n1056), .A2(G952), .ZN(n1119) );
XOR2_X1 U856 ( .A(n1184), .B(n1174), .Z(G48) );
NAND4_X1 U857 ( .A1(n1185), .A2(n1051), .A3(n1073), .A4(n1083), .ZN(n1174) );
XOR2_X1 U858 ( .A(n1173), .B(n1186), .Z(G45) );
NAND2_X1 U859 ( .A1(KEYINPUT14), .A2(G143), .ZN(n1186) );
NAND4_X1 U860 ( .A1(n1179), .A2(n1052), .A3(n1041), .A4(n1187), .ZN(n1173) );
XOR2_X1 U861 ( .A(n1188), .B(n1172), .Z(G42) );
NAND4_X1 U862 ( .A1(n1061), .A2(n1185), .A3(n1065), .A4(n1051), .ZN(n1172) );
XNOR2_X1 U863 ( .A(G137), .B(n1171), .ZN(G39) );
NAND4_X1 U864 ( .A1(n1053), .A2(n1061), .A3(n1185), .A4(n1083), .ZN(n1171) );
XOR2_X1 U865 ( .A(G134), .B(n1170), .Z(G36) );
AND2_X1 U866 ( .A1(n1189), .A2(n1067), .ZN(n1170) );
XOR2_X1 U867 ( .A(n1169), .B(n1190), .Z(G33) );
XOR2_X1 U868 ( .A(KEYINPUT18), .B(G131), .Z(n1190) );
AND2_X1 U869 ( .A1(n1189), .A2(n1051), .ZN(n1169) );
AND4_X1 U870 ( .A1(n1052), .A2(n1061), .A3(n1041), .A4(n1187), .ZN(n1189) );
INV_X1 U871 ( .A(n1034), .ZN(n1061) );
NAND2_X1 U872 ( .A1(n1075), .A2(n1191), .ZN(n1034) );
XOR2_X1 U873 ( .A(n1192), .B(n1193), .Z(G30) );
NOR2_X1 U874 ( .A1(n1168), .A2(KEYINPUT40), .ZN(n1193) );
AND4_X1 U875 ( .A1(n1185), .A2(n1067), .A3(n1073), .A4(n1083), .ZN(n1168) );
AND3_X1 U876 ( .A1(n1066), .A2(n1187), .A3(n1041), .ZN(n1185) );
XNOR2_X1 U877 ( .A(G101), .B(n1181), .ZN(G3) );
NAND3_X1 U878 ( .A1(n1052), .A2(n1183), .A3(n1053), .ZN(n1181) );
XOR2_X1 U879 ( .A(n1194), .B(n1195), .Z(G27) );
NAND2_X1 U880 ( .A1(KEYINPUT3), .A2(n1167), .ZN(n1195) );
AND4_X1 U881 ( .A1(n1065), .A2(n1051), .A3(n1047), .A4(n1196), .ZN(n1167) );
AND3_X1 U882 ( .A1(n1073), .A2(n1187), .A3(n1066), .ZN(n1196) );
NAND2_X1 U883 ( .A1(n1044), .A2(n1197), .ZN(n1187) );
NAND4_X1 U884 ( .A1(G902), .A2(G953), .A3(n1198), .A4(n1095), .ZN(n1197) );
INV_X1 U885 ( .A(G900), .ZN(n1095) );
NAND2_X1 U886 ( .A1(n1199), .A2(n1200), .ZN(G24) );
NAND2_X1 U887 ( .A1(G122), .A2(n1201), .ZN(n1200) );
XOR2_X1 U888 ( .A(KEYINPUT7), .B(n1202), .Z(n1199) );
NOR2_X1 U889 ( .A1(G122), .A2(n1201), .ZN(n1202) );
NAND3_X1 U890 ( .A1(n1180), .A2(n1179), .A3(n1203), .ZN(n1201) );
XNOR2_X1 U891 ( .A(n1050), .B(KEYINPUT20), .ZN(n1203) );
NOR2_X1 U892 ( .A1(n1066), .A2(n1083), .ZN(n1050) );
AND3_X1 U893 ( .A1(n1204), .A2(n1205), .A3(n1073), .ZN(n1179) );
XOR2_X1 U894 ( .A(n1206), .B(n1176), .Z(G21) );
NAND4_X1 U895 ( .A1(n1083), .A2(n1066), .A3(n1073), .A4(n1207), .ZN(n1176) );
AND2_X1 U896 ( .A1(n1053), .A2(n1180), .ZN(n1207) );
INV_X1 U897 ( .A(n1065), .ZN(n1083) );
XNOR2_X1 U898 ( .A(G116), .B(n1178), .ZN(G18) );
NAND4_X1 U899 ( .A1(n1180), .A2(n1052), .A3(n1067), .A4(n1073), .ZN(n1178) );
NOR2_X1 U900 ( .A1(n1204), .A2(n1208), .ZN(n1067) );
XOR2_X1 U901 ( .A(n1209), .B(n1177), .Z(G15) );
NAND4_X1 U902 ( .A1(n1180), .A2(n1052), .A3(n1051), .A4(n1210), .ZN(n1177) );
INV_X1 U903 ( .A(n1087), .ZN(n1051) );
NAND2_X1 U904 ( .A1(n1208), .A2(n1204), .ZN(n1087) );
NOR2_X1 U905 ( .A1(n1066), .A2(n1065), .ZN(n1052) );
AND2_X1 U906 ( .A1(n1047), .A2(n1211), .ZN(n1180) );
NOR2_X1 U907 ( .A1(n1043), .A2(n1212), .ZN(n1047) );
INV_X1 U908 ( .A(n1213), .ZN(n1043) );
NAND2_X1 U909 ( .A1(n1214), .A2(n1215), .ZN(G12) );
NAND2_X1 U910 ( .A1(n1216), .A2(n1182), .ZN(n1215) );
XOR2_X1 U911 ( .A(n1217), .B(KEYINPUT51), .Z(n1214) );
OR2_X1 U912 ( .A1(n1182), .A2(n1216), .ZN(n1217) );
XNOR2_X1 U913 ( .A(G110), .B(KEYINPUT17), .ZN(n1216) );
NAND4_X1 U914 ( .A1(n1053), .A2(n1183), .A3(n1065), .A4(n1066), .ZN(n1182) );
XNOR2_X1 U915 ( .A(n1218), .B(n1125), .ZN(n1066) );
AND2_X1 U916 ( .A1(G217), .A2(n1219), .ZN(n1125) );
NAND2_X1 U917 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
XNOR2_X1 U918 ( .A(n1122), .B(KEYINPUT60), .ZN(n1220) );
XNOR2_X1 U919 ( .A(n1222), .B(n1223), .ZN(n1122) );
XOR2_X1 U920 ( .A(n1224), .B(n1225), .Z(n1223) );
XOR2_X1 U921 ( .A(n1226), .B(n1227), .Z(n1225) );
NOR3_X1 U922 ( .A1(n1228), .A2(KEYINPUT48), .A3(n1229), .ZN(n1227) );
NOR2_X1 U923 ( .A1(G146), .A2(n1230), .ZN(n1229) );
XNOR2_X1 U924 ( .A(KEYINPUT35), .B(n1231), .ZN(n1230) );
XOR2_X1 U925 ( .A(KEYINPUT54), .B(n1232), .Z(n1228) );
NOR2_X1 U926 ( .A1(n1184), .A2(n1233), .ZN(n1232) );
XOR2_X1 U927 ( .A(KEYINPUT35), .B(n1231), .Z(n1233) );
NAND2_X1 U928 ( .A1(n1234), .A2(G221), .ZN(n1226) );
NAND2_X1 U929 ( .A1(KEYINPUT25), .A2(n1206), .ZN(n1224) );
XOR2_X1 U930 ( .A(n1235), .B(n1236), .Z(n1222) );
XOR2_X1 U931 ( .A(KEYINPUT52), .B(G137), .Z(n1236) );
XOR2_X1 U932 ( .A(G110), .B(n1192), .Z(n1235) );
XOR2_X1 U933 ( .A(n1237), .B(G472), .Z(n1065) );
NAND2_X1 U934 ( .A1(n1238), .A2(n1221), .ZN(n1237) );
XOR2_X1 U935 ( .A(n1138), .B(n1239), .Z(n1238) );
NOR2_X1 U936 ( .A1(KEYINPUT63), .A2(n1240), .ZN(n1239) );
XOR2_X1 U937 ( .A(n1241), .B(KEYINPUT10), .Z(n1240) );
NAND2_X1 U938 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND2_X1 U939 ( .A1(n1244), .A2(n1137), .ZN(n1243) );
XOR2_X1 U940 ( .A(KEYINPUT21), .B(n1245), .Z(n1242) );
NOR2_X1 U941 ( .A1(n1244), .A2(n1137), .ZN(n1245) );
XNOR2_X1 U942 ( .A(G113), .B(n1246), .ZN(n1137) );
NOR2_X1 U943 ( .A1(KEYINPUT9), .A2(n1247), .ZN(n1246) );
XNOR2_X1 U944 ( .A(G116), .B(n1248), .ZN(n1247) );
NAND2_X1 U945 ( .A1(KEYINPUT1), .A2(n1206), .ZN(n1248) );
INV_X1 U946 ( .A(G119), .ZN(n1206) );
AND3_X1 U947 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1244) );
OR2_X1 U948 ( .A1(n1145), .A2(KEYINPUT5), .ZN(n1251) );
NAND3_X1 U949 ( .A1(KEYINPUT5), .A2(n1252), .A3(n1253), .ZN(n1250) );
OR2_X1 U950 ( .A1(n1253), .A2(n1252), .ZN(n1249) );
NOR2_X1 U951 ( .A1(KEYINPUT6), .A2(n1254), .ZN(n1252) );
INV_X1 U952 ( .A(n1145), .ZN(n1254) );
XOR2_X1 U953 ( .A(n1255), .B(G101), .Z(n1138) );
NAND2_X1 U954 ( .A1(n1256), .A2(G210), .ZN(n1255) );
AND3_X1 U955 ( .A1(n1210), .A2(n1211), .A3(n1041), .ZN(n1183) );
NOR2_X1 U956 ( .A1(n1212), .A2(n1213), .ZN(n1041) );
XOR2_X1 U957 ( .A(n1086), .B(G469), .Z(n1213) );
NAND2_X1 U958 ( .A1(n1257), .A2(n1221), .ZN(n1086) );
XOR2_X1 U959 ( .A(n1258), .B(n1259), .Z(n1257) );
XNOR2_X1 U960 ( .A(n1154), .B(n1150), .ZN(n1259) );
XOR2_X1 U961 ( .A(n1260), .B(n1145), .Z(n1150) );
XOR2_X1 U962 ( .A(n1261), .B(n1262), .Z(n1145) );
NOR2_X1 U963 ( .A1(G137), .A2(KEYINPUT15), .ZN(n1262) );
XOR2_X1 U964 ( .A(n1263), .B(G134), .Z(n1261) );
INV_X1 U965 ( .A(G131), .ZN(n1263) );
NAND2_X1 U966 ( .A1(n1264), .A2(n1056), .ZN(n1260) );
XOR2_X1 U967 ( .A(KEYINPUT44), .B(G227), .Z(n1264) );
XNOR2_X1 U968 ( .A(n1265), .B(n1266), .ZN(n1154) );
XNOR2_X1 U969 ( .A(n1267), .B(n1099), .ZN(n1266) );
XOR2_X1 U970 ( .A(n1268), .B(n1192), .Z(n1099) );
NAND2_X1 U971 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
XOR2_X1 U972 ( .A(n1271), .B(KEYINPUT45), .Z(n1269) );
XOR2_X1 U973 ( .A(n1272), .B(KEYINPUT27), .Z(n1265) );
XOR2_X1 U974 ( .A(G110), .B(n1188), .Z(n1258) );
INV_X1 U975 ( .A(G140), .ZN(n1188) );
XNOR2_X1 U976 ( .A(n1042), .B(KEYINPUT53), .ZN(n1212) );
NAND2_X1 U977 ( .A1(G221), .A2(n1219), .ZN(n1042) );
NAND2_X1 U978 ( .A1(G234), .A2(n1221), .ZN(n1219) );
NAND2_X1 U979 ( .A1(n1044), .A2(n1273), .ZN(n1211) );
NAND3_X1 U980 ( .A1(n1274), .A2(n1198), .A3(G902), .ZN(n1273) );
INV_X1 U981 ( .A(n1114), .ZN(n1274) );
NAND2_X1 U982 ( .A1(G953), .A2(n1275), .ZN(n1114) );
XOR2_X1 U983 ( .A(KEYINPUT49), .B(G898), .Z(n1275) );
NAND3_X1 U984 ( .A1(n1198), .A2(n1056), .A3(G952), .ZN(n1044) );
NAND2_X1 U985 ( .A1(G237), .A2(G234), .ZN(n1198) );
XOR2_X1 U986 ( .A(n1073), .B(KEYINPUT0), .Z(n1210) );
NOR2_X1 U987 ( .A1(n1075), .A2(n1074), .ZN(n1073) );
INV_X1 U988 ( .A(n1191), .ZN(n1074) );
NAND2_X1 U989 ( .A1(G214), .A2(n1276), .ZN(n1191) );
XOR2_X1 U990 ( .A(n1080), .B(KEYINPUT58), .Z(n1075) );
XNOR2_X1 U991 ( .A(n1277), .B(n1164), .ZN(n1080) );
AND2_X1 U992 ( .A1(G210), .A2(n1276), .ZN(n1164) );
NAND2_X1 U993 ( .A1(n1278), .A2(n1221), .ZN(n1276) );
INV_X1 U994 ( .A(G237), .ZN(n1278) );
NAND2_X1 U995 ( .A1(n1279), .A2(n1221), .ZN(n1277) );
XOR2_X1 U996 ( .A(n1163), .B(n1280), .Z(n1279) );
XNOR2_X1 U997 ( .A(n1158), .B(n1281), .ZN(n1280) );
NAND2_X1 U998 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U999 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U1000 ( .A(KEYINPUT55), .B(n1253), .Z(n1285) );
INV_X1 U1001 ( .A(n1144), .ZN(n1253) );
XOR2_X1 U1002 ( .A(n1194), .B(KEYINPUT32), .Z(n1284) );
INV_X1 U1003 ( .A(G125), .ZN(n1194) );
NAND2_X1 U1004 ( .A1(n1286), .A2(n1287), .ZN(n1282) );
XOR2_X1 U1005 ( .A(KEYINPUT47), .B(G125), .Z(n1287) );
XOR2_X1 U1006 ( .A(KEYINPUT55), .B(n1144), .Z(n1286) );
XOR2_X1 U1007 ( .A(n1288), .B(G128), .Z(n1144) );
NAND3_X1 U1008 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1288) );
XOR2_X1 U1009 ( .A(n1271), .B(KEYINPUT38), .Z(n1291) );
NAND2_X1 U1010 ( .A1(n1292), .A2(n1293), .ZN(n1290) );
OR3_X1 U1011 ( .A1(G143), .A2(G146), .A3(n1293), .ZN(n1289) );
INV_X1 U1012 ( .A(KEYINPUT61), .ZN(n1293) );
AND2_X1 U1013 ( .A1(G224), .A2(n1056), .ZN(n1158) );
XOR2_X1 U1014 ( .A(n1294), .B(n1295), .Z(n1163) );
INV_X1 U1015 ( .A(n1118), .ZN(n1295) );
XOR2_X1 U1016 ( .A(n1272), .B(n1296), .Z(n1118) );
NOR2_X1 U1017 ( .A1(KEYINPUT36), .A2(n1267), .ZN(n1296) );
XNOR2_X1 U1018 ( .A(G101), .B(KEYINPUT24), .ZN(n1267) );
XOR2_X1 U1019 ( .A(n1297), .B(n1298), .Z(n1272) );
XNOR2_X1 U1020 ( .A(n1299), .B(n1300), .ZN(n1294) );
NOR2_X1 U1021 ( .A1(KEYINPUT56), .A2(n1115), .ZN(n1300) );
XOR2_X1 U1022 ( .A(G110), .B(n1301), .Z(n1115) );
NOR2_X1 U1023 ( .A1(KEYINPUT12), .A2(n1117), .ZN(n1299) );
NAND2_X1 U1024 ( .A1(n1302), .A2(n1303), .ZN(n1117) );
NAND2_X1 U1025 ( .A1(n1304), .A2(n1209), .ZN(n1303) );
XOR2_X1 U1026 ( .A(n1305), .B(KEYINPUT57), .Z(n1302) );
OR2_X1 U1027 ( .A1(n1209), .A2(n1304), .ZN(n1305) );
XOR2_X1 U1028 ( .A(G116), .B(n1306), .Z(n1304) );
NOR2_X1 U1029 ( .A1(G119), .A2(KEYINPUT50), .ZN(n1306) );
NOR2_X1 U1030 ( .A1(n1205), .A2(n1204), .ZN(n1053) );
XOR2_X1 U1031 ( .A(G475), .B(n1307), .Z(n1204) );
AND2_X1 U1032 ( .A1(n1221), .A2(n1131), .ZN(n1307) );
XNOR2_X1 U1033 ( .A(n1308), .B(n1309), .ZN(n1131) );
XOR2_X1 U1034 ( .A(n1098), .B(n1310), .Z(n1309) );
INV_X1 U1035 ( .A(n1297), .ZN(n1310) );
XNOR2_X1 U1036 ( .A(G104), .B(KEYINPUT13), .ZN(n1297) );
XOR2_X1 U1037 ( .A(G131), .B(n1231), .Z(n1098) );
XOR2_X1 U1038 ( .A(G125), .B(G140), .Z(n1231) );
NAND2_X1 U1039 ( .A1(n1311), .A2(n1312), .ZN(n1308) );
NAND2_X1 U1040 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
NAND2_X1 U1041 ( .A1(n1271), .A2(n1270), .ZN(n1314) );
INV_X1 U1042 ( .A(n1292), .ZN(n1270) );
NOR2_X1 U1043 ( .A1(n1184), .A2(G143), .ZN(n1292) );
NAND2_X1 U1044 ( .A1(G143), .A2(n1184), .ZN(n1271) );
NAND2_X1 U1045 ( .A1(n1315), .A2(n1316), .ZN(n1311) );
XOR2_X1 U1046 ( .A(G143), .B(n1184), .Z(n1316) );
INV_X1 U1047 ( .A(G146), .ZN(n1184) );
INV_X1 U1048 ( .A(n1313), .ZN(n1315) );
XOR2_X1 U1049 ( .A(n1317), .B(n1318), .Z(n1313) );
NOR3_X1 U1050 ( .A1(KEYINPUT28), .A2(n1319), .A3(n1320), .ZN(n1318) );
NOR2_X1 U1051 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
INV_X1 U1052 ( .A(KEYINPUT26), .ZN(n1322) );
NOR2_X1 U1053 ( .A1(n1323), .A2(n1324), .ZN(n1321) );
NOR2_X1 U1054 ( .A1(n1301), .A2(n1325), .ZN(n1324) );
NOR2_X1 U1055 ( .A1(G122), .A2(n1209), .ZN(n1323) );
NOR2_X1 U1056 ( .A1(KEYINPUT26), .A2(n1326), .ZN(n1319) );
NOR2_X1 U1057 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
NOR2_X1 U1058 ( .A1(n1209), .A2(n1301), .ZN(n1328) );
INV_X1 U1059 ( .A(G122), .ZN(n1301) );
INV_X1 U1060 ( .A(G113), .ZN(n1209) );
NOR2_X1 U1061 ( .A1(G122), .A2(n1325), .ZN(n1327) );
XOR2_X1 U1062 ( .A(n1329), .B(G113), .Z(n1325) );
XNOR2_X1 U1063 ( .A(KEYINPUT39), .B(KEYINPUT29), .ZN(n1329) );
NAND2_X1 U1064 ( .A1(n1256), .A2(G214), .ZN(n1317) );
NOR2_X1 U1065 ( .A1(G953), .A2(G237), .ZN(n1256) );
INV_X1 U1066 ( .A(n1208), .ZN(n1205) );
XOR2_X1 U1067 ( .A(n1330), .B(G478), .Z(n1208) );
NAND2_X1 U1068 ( .A1(n1128), .A2(n1221), .ZN(n1330) );
INV_X1 U1069 ( .A(G902), .ZN(n1221) );
XNOR2_X1 U1070 ( .A(n1331), .B(n1332), .ZN(n1128) );
XOR2_X1 U1071 ( .A(n1333), .B(n1334), .Z(n1332) );
XOR2_X1 U1072 ( .A(KEYINPUT31), .B(G134), .Z(n1334) );
NOR2_X1 U1073 ( .A1(KEYINPUT30), .A2(n1335), .ZN(n1333) );
XOR2_X1 U1074 ( .A(n1192), .B(G143), .Z(n1335) );
INV_X1 U1075 ( .A(G128), .ZN(n1192) );
XOR2_X1 U1076 ( .A(n1336), .B(n1337), .Z(n1331) );
AND2_X1 U1077 ( .A1(n1234), .A2(G217), .ZN(n1337) );
AND2_X1 U1078 ( .A1(G234), .A2(n1056), .ZN(n1234) );
INV_X1 U1079 ( .A(G953), .ZN(n1056) );
NAND3_X1 U1080 ( .A1(n1338), .A2(n1339), .A3(n1340), .ZN(n1336) );
OR2_X1 U1081 ( .A1(n1341), .A2(KEYINPUT8), .ZN(n1340) );
NAND3_X1 U1082 ( .A1(KEYINPUT8), .A2(n1342), .A3(n1298), .ZN(n1339) );
OR2_X1 U1083 ( .A1(n1298), .A2(n1342), .ZN(n1338) );
AND2_X1 U1084 ( .A1(KEYINPUT62), .A2(n1341), .ZN(n1342) );
XOR2_X1 U1085 ( .A(G116), .B(G122), .Z(n1341) );
XOR2_X1 U1086 ( .A(G107), .B(KEYINPUT19), .Z(n1298) );
endmodule


