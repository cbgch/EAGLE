//Key = 0101111001011001000100101111111000011011011110010100001110100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357;

XNOR2_X1 U756 ( .A(G107), .B(n1029), .ZN(G9) );
NOR2_X1 U757 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U758 ( .A1(G953), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1031) );
NOR2_X1 U759 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U760 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U761 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U762 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U763 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U764 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U765 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR3_X1 U766 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1047) );
NOR2_X1 U767 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XOR2_X1 U768 ( .A(KEYINPUT16), .B(n1054), .Z(n1053) );
NOR2_X1 U769 ( .A1(KEYINPUT29), .A2(n1055), .ZN(n1049) );
NOR2_X1 U770 ( .A1(n1056), .A2(n1055), .ZN(n1045) );
NOR2_X1 U771 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
XOR2_X1 U772 ( .A(KEYINPUT50), .B(n1059), .Z(n1058) );
NOR3_X1 U773 ( .A1(n1048), .A2(n1060), .A3(n1055), .ZN(n1041) );
NOR2_X1 U774 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR3_X1 U775 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1061) );
INV_X1 U776 ( .A(KEYINPUT29), .ZN(n1063) );
NOR4_X1 U777 ( .A1(n1066), .A2(n1055), .A3(n1048), .A4(n1044), .ZN(n1037) );
INV_X1 U778 ( .A(n1067), .ZN(n1044) );
INV_X1 U779 ( .A(n1068), .ZN(n1048) );
NOR2_X1 U780 ( .A1(n1069), .A2(n1070), .ZN(n1066) );
NOR3_X1 U781 ( .A1(n1032), .A2(G953), .A3(G952), .ZN(n1030) );
AND4_X1 U782 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1032) );
NOR4_X1 U783 ( .A1(n1065), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1074) );
XOR2_X1 U784 ( .A(KEYINPUT61), .B(n1078), .Z(n1077) );
XNOR2_X1 U785 ( .A(n1079), .B(n1080), .ZN(n1076) );
NOR2_X1 U786 ( .A1(KEYINPUT7), .A2(n1081), .ZN(n1080) );
NOR2_X1 U787 ( .A1(n1082), .A2(n1083), .ZN(n1073) );
XNOR2_X1 U788 ( .A(n1084), .B(KEYINPUT4), .ZN(n1083) );
XOR2_X1 U789 ( .A(n1085), .B(n1086), .Z(n1072) );
NAND2_X1 U790 ( .A1(KEYINPUT54), .A2(n1087), .ZN(n1086) );
XOR2_X1 U791 ( .A(KEYINPUT3), .B(n1088), .Z(n1087) );
XOR2_X1 U792 ( .A(n1089), .B(n1090), .Z(G72) );
XOR2_X1 U793 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U794 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U795 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U796 ( .A1(KEYINPUT48), .A2(n1097), .ZN(n1096) );
XOR2_X1 U797 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND3_X1 U798 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1098) );
NAND2_X1 U799 ( .A1(n1103), .A2(G131), .ZN(n1102) );
NAND2_X1 U800 ( .A1(KEYINPUT0), .A2(n1104), .ZN(n1101) );
NAND2_X1 U801 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XNOR2_X1 U802 ( .A(KEYINPUT18), .B(n1103), .ZN(n1105) );
NAND2_X1 U803 ( .A1(n1107), .A2(n1108), .ZN(n1100) );
INV_X1 U804 ( .A(KEYINPUT0), .ZN(n1108) );
NAND2_X1 U805 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
OR3_X1 U806 ( .A1(n1103), .A2(G131), .A3(KEYINPUT18), .ZN(n1110) );
NAND2_X1 U807 ( .A1(KEYINPUT18), .A2(n1103), .ZN(n1109) );
AND2_X1 U808 ( .A1(n1111), .A2(n1112), .ZN(n1103) );
NAND2_X1 U809 ( .A1(KEYINPUT27), .A2(n1113), .ZN(n1112) );
XOR2_X1 U810 ( .A(G134), .B(n1114), .Z(n1113) );
NAND3_X1 U811 ( .A1(G134), .A2(n1114), .A3(n1115), .ZN(n1111) );
INV_X1 U812 ( .A(KEYINPUT27), .ZN(n1115) );
NAND2_X1 U813 ( .A1(n1116), .A2(n1117), .ZN(n1091) );
NAND2_X1 U814 ( .A1(G900), .A2(G227), .ZN(n1117) );
INV_X1 U815 ( .A(n1118), .ZN(n1116) );
NAND3_X1 U816 ( .A1(n1119), .A2(n1120), .A3(KEYINPUT35), .ZN(n1089) );
XOR2_X1 U817 ( .A(n1121), .B(n1122), .Z(G69) );
NOR2_X1 U818 ( .A1(n1123), .A2(n1118), .ZN(n1122) );
XOR2_X1 U819 ( .A(n1120), .B(KEYINPUT45), .Z(n1118) );
AND2_X1 U820 ( .A1(G224), .A2(G898), .ZN(n1123) );
NAND2_X1 U821 ( .A1(n1124), .A2(n1125), .ZN(n1121) );
NAND2_X1 U822 ( .A1(n1126), .A2(n1120), .ZN(n1125) );
XNOR2_X1 U823 ( .A(n1127), .B(n1128), .ZN(n1126) );
OR3_X1 U824 ( .A1(n1127), .A2(n1129), .A3(n1120), .ZN(n1124) );
NOR2_X1 U825 ( .A1(n1130), .A2(n1131), .ZN(G66) );
XOR2_X1 U826 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U827 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
NOR2_X1 U828 ( .A1(n1130), .A2(n1136), .ZN(G63) );
XOR2_X1 U829 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U830 ( .A1(n1139), .A2(n1135), .ZN(n1138) );
INV_X1 U831 ( .A(G478), .ZN(n1139) );
NOR3_X1 U832 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(G60) );
AND2_X1 U833 ( .A1(KEYINPUT43), .A2(n1130), .ZN(n1142) );
NOR3_X1 U834 ( .A1(KEYINPUT43), .A2(G953), .A3(G952), .ZN(n1141) );
XOR2_X1 U835 ( .A(n1143), .B(n1144), .Z(n1140) );
NOR2_X1 U836 ( .A1(n1085), .A2(n1135), .ZN(n1143) );
INV_X1 U837 ( .A(G475), .ZN(n1085) );
XNOR2_X1 U838 ( .A(G104), .B(n1145), .ZN(G6) );
NOR2_X1 U839 ( .A1(n1130), .A2(n1146), .ZN(G57) );
XOR2_X1 U840 ( .A(n1147), .B(n1148), .Z(n1146) );
NAND3_X1 U841 ( .A1(G472), .A2(n1149), .A3(G902), .ZN(n1147) );
XNOR2_X1 U842 ( .A(KEYINPUT1), .B(n1034), .ZN(n1149) );
NOR2_X1 U843 ( .A1(n1130), .A2(n1150), .ZN(G54) );
XOR2_X1 U844 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U845 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U846 ( .A1(n1155), .A2(n1135), .ZN(n1153) );
INV_X1 U847 ( .A(G469), .ZN(n1155) );
XOR2_X1 U848 ( .A(n1099), .B(n1156), .Z(n1151) );
NOR2_X1 U849 ( .A1(n1130), .A2(n1157), .ZN(G51) );
XOR2_X1 U850 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U851 ( .A1(n1079), .A2(n1135), .ZN(n1159) );
NAND2_X1 U852 ( .A1(G902), .A2(n1034), .ZN(n1135) );
OR2_X1 U853 ( .A1(n1119), .A2(n1128), .ZN(n1034) );
NAND4_X1 U854 ( .A1(n1160), .A2(n1145), .A3(n1161), .A4(n1162), .ZN(n1128) );
AND4_X1 U855 ( .A1(n1029), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1162) );
NAND3_X1 U856 ( .A1(n1068), .A2(n1166), .A3(n1069), .ZN(n1029) );
OR2_X1 U857 ( .A1(n1167), .A2(n1168), .ZN(n1161) );
NAND3_X1 U858 ( .A1(n1068), .A2(n1166), .A3(n1070), .ZN(n1145) );
NAND2_X1 U859 ( .A1(n1169), .A2(n1170), .ZN(n1160) );
NAND2_X1 U860 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND3_X1 U861 ( .A1(n1078), .A2(n1173), .A3(n1068), .ZN(n1172) );
NAND2_X1 U862 ( .A1(n1174), .A2(n1175), .ZN(n1171) );
NAND4_X1 U863 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1119) );
AND4_X1 U864 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1179) );
NOR2_X1 U865 ( .A1(n1184), .A2(n1185), .ZN(n1178) );
NOR2_X1 U866 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NOR2_X1 U867 ( .A1(n1188), .A2(n1189), .ZN(n1186) );
AND2_X1 U868 ( .A1(n1190), .A2(KEYINPUT47), .ZN(n1189) );
NOR3_X1 U869 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1188) );
NOR2_X1 U870 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
INV_X1 U871 ( .A(KEYINPUT17), .ZN(n1195) );
NOR2_X1 U872 ( .A1(n1196), .A2(n1197), .ZN(n1194) );
NOR2_X1 U873 ( .A1(KEYINPUT17), .A2(n1198), .ZN(n1192) );
INV_X1 U874 ( .A(n1057), .ZN(n1191) );
NOR4_X1 U875 ( .A1(KEYINPUT47), .A2(n1070), .A3(n1055), .A4(n1199), .ZN(n1184) );
INV_X1 U876 ( .A(n1200), .ZN(n1055) );
NAND4_X1 U877 ( .A1(n1201), .A2(n1198), .A3(n1069), .A4(n1202), .ZN(n1176) );
XOR2_X1 U878 ( .A(KEYINPUT32), .B(n1175), .Z(n1202) );
XOR2_X1 U879 ( .A(n1168), .B(KEYINPUT41), .Z(n1201) );
NOR2_X1 U880 ( .A1(n1203), .A2(n1204), .ZN(n1158) );
XOR2_X1 U881 ( .A(n1205), .B(KEYINPUT42), .Z(n1204) );
NAND2_X1 U882 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NOR2_X1 U883 ( .A1(n1207), .A2(n1206), .ZN(n1203) );
XNOR2_X1 U884 ( .A(KEYINPUT63), .B(n1208), .ZN(n1206) );
NOR2_X1 U885 ( .A1(n1120), .A2(G952), .ZN(n1130) );
XOR2_X1 U886 ( .A(n1209), .B(n1180), .Z(G48) );
NAND4_X1 U887 ( .A1(n1070), .A2(n1175), .A3(n1198), .A4(n1050), .ZN(n1180) );
XNOR2_X1 U888 ( .A(n1177), .B(n1210), .ZN(G45) );
NOR2_X1 U889 ( .A1(KEYINPUT10), .A2(n1211), .ZN(n1210) );
NAND4_X1 U890 ( .A1(n1190), .A2(n1050), .A3(n1078), .A4(n1173), .ZN(n1177) );
XOR2_X1 U891 ( .A(n1212), .B(n1213), .Z(G42) );
NAND4_X1 U892 ( .A1(n1214), .A2(n1057), .A3(n1215), .A4(n1197), .ZN(n1213) );
XOR2_X1 U893 ( .A(KEYINPUT37), .B(n1062), .Z(n1215) );
INV_X1 U894 ( .A(n1187), .ZN(n1214) );
XOR2_X1 U895 ( .A(n1114), .B(n1183), .Z(G39) );
NAND4_X1 U896 ( .A1(n1174), .A2(n1175), .A3(n1198), .A4(n1200), .ZN(n1183) );
XNOR2_X1 U897 ( .A(G134), .B(n1182), .ZN(G36) );
NAND3_X1 U898 ( .A1(n1069), .A2(n1200), .A3(n1190), .ZN(n1182) );
INV_X1 U899 ( .A(n1199), .ZN(n1190) );
XOR2_X1 U900 ( .A(G131), .B(n1216), .Z(G33) );
NOR2_X1 U901 ( .A1(n1199), .A2(n1187), .ZN(n1216) );
NAND2_X1 U902 ( .A1(n1070), .A2(n1200), .ZN(n1187) );
NAND2_X1 U903 ( .A1(n1217), .A2(n1218), .ZN(n1200) );
OR3_X1 U904 ( .A1(n1054), .A2(n1082), .A3(KEYINPUT16), .ZN(n1218) );
INV_X1 U905 ( .A(n1052), .ZN(n1082) );
NAND2_X1 U906 ( .A1(KEYINPUT16), .A2(n1050), .ZN(n1217) );
NAND2_X1 U907 ( .A1(n1059), .A2(n1198), .ZN(n1199) );
XNOR2_X1 U908 ( .A(G128), .B(n1219), .ZN(G30) );
NAND4_X1 U909 ( .A1(n1175), .A2(n1198), .A3(n1069), .A4(n1050), .ZN(n1219) );
NOR2_X1 U910 ( .A1(n1196), .A2(n1220), .ZN(n1198) );
XOR2_X1 U911 ( .A(n1221), .B(n1165), .Z(G3) );
NAND3_X1 U912 ( .A1(n1059), .A2(n1166), .A3(n1174), .ZN(n1165) );
AND3_X1 U913 ( .A1(n1062), .A2(n1222), .A3(n1050), .ZN(n1166) );
XNOR2_X1 U914 ( .A(G125), .B(n1181), .ZN(G27) );
NAND4_X1 U915 ( .A1(n1057), .A2(n1067), .A3(n1223), .A4(n1070), .ZN(n1181) );
NOR2_X1 U916 ( .A1(n1220), .A2(n1168), .ZN(n1223) );
INV_X1 U917 ( .A(n1197), .ZN(n1220) );
NAND2_X1 U918 ( .A1(n1224), .A2(n1225), .ZN(n1197) );
NAND3_X1 U919 ( .A1(G902), .A2(n1226), .A3(n1093), .ZN(n1225) );
NOR2_X1 U920 ( .A1(n1120), .A2(G900), .ZN(n1093) );
XOR2_X1 U921 ( .A(n1227), .B(n1228), .Z(G24) );
NAND4_X1 U922 ( .A1(KEYINPUT9), .A2(n1169), .A3(n1229), .A4(n1068), .ZN(n1228) );
NOR2_X1 U923 ( .A1(n1075), .A2(n1230), .ZN(n1068) );
NOR2_X1 U924 ( .A1(n1231), .A2(n1232), .ZN(n1229) );
XNOR2_X1 U925 ( .A(G119), .B(n1233), .ZN(G21) );
NAND3_X1 U926 ( .A1(n1174), .A2(n1234), .A3(n1169), .ZN(n1233) );
XOR2_X1 U927 ( .A(KEYINPUT33), .B(n1175), .Z(n1234) );
AND2_X1 U928 ( .A1(n1230), .A2(n1075), .ZN(n1175) );
INV_X1 U929 ( .A(n1235), .ZN(n1230) );
XOR2_X1 U930 ( .A(n1164), .B(n1236), .Z(G18) );
NAND2_X1 U931 ( .A1(KEYINPUT56), .A2(G116), .ZN(n1236) );
NAND3_X1 U932 ( .A1(n1059), .A2(n1069), .A3(n1169), .ZN(n1164) );
NOR2_X1 U933 ( .A1(n1173), .A2(n1232), .ZN(n1069) );
INV_X1 U934 ( .A(n1231), .ZN(n1173) );
XOR2_X1 U935 ( .A(n1237), .B(n1163), .Z(G15) );
NAND3_X1 U936 ( .A1(n1059), .A2(n1070), .A3(n1169), .ZN(n1163) );
AND3_X1 U937 ( .A1(n1050), .A2(n1222), .A3(n1067), .ZN(n1169) );
NOR2_X1 U938 ( .A1(n1065), .A2(n1084), .ZN(n1067) );
INV_X1 U939 ( .A(n1064), .ZN(n1084) );
NOR2_X1 U940 ( .A1(n1078), .A2(n1231), .ZN(n1070) );
INV_X1 U941 ( .A(n1232), .ZN(n1078) );
AND2_X1 U942 ( .A1(n1235), .A2(n1075), .ZN(n1059) );
XOR2_X1 U943 ( .A(n1238), .B(n1239), .Z(G12) );
NAND2_X1 U944 ( .A1(n1240), .A2(n1050), .ZN(n1239) );
INV_X1 U945 ( .A(n1168), .ZN(n1050) );
NAND2_X1 U946 ( .A1(n1054), .A2(n1052), .ZN(n1168) );
NAND2_X1 U947 ( .A1(G214), .A2(n1241), .ZN(n1052) );
XOR2_X1 U948 ( .A(n1081), .B(n1079), .Z(n1054) );
NAND2_X1 U949 ( .A1(G210), .A2(n1241), .ZN(n1079) );
NAND2_X1 U950 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
INV_X1 U951 ( .A(G237), .ZN(n1242) );
NAND2_X1 U952 ( .A1(n1244), .A2(n1243), .ZN(n1081) );
XOR2_X1 U953 ( .A(n1208), .B(n1207), .Z(n1244) );
XOR2_X1 U954 ( .A(n1245), .B(n1127), .Z(n1207) );
XOR2_X1 U955 ( .A(n1246), .B(n1247), .Z(n1127) );
XOR2_X1 U956 ( .A(n1248), .B(n1249), .Z(n1247) );
NAND2_X1 U957 ( .A1(KEYINPUT58), .A2(n1250), .ZN(n1249) );
NAND3_X1 U958 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1248) );
NAND2_X1 U959 ( .A1(n1254), .A2(n1238), .ZN(n1253) );
NAND3_X1 U960 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1254) );
NAND2_X1 U961 ( .A1(KEYINPUT2), .A2(n1258), .ZN(n1257) );
NAND2_X1 U962 ( .A1(KEYINPUT60), .A2(n1227), .ZN(n1256) );
NAND2_X1 U963 ( .A1(n1259), .A2(n1260), .ZN(n1255) );
INV_X1 U964 ( .A(KEYINPUT60), .ZN(n1260) );
NAND2_X1 U965 ( .A1(n1227), .A2(n1261), .ZN(n1259) );
NAND2_X1 U966 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NAND4_X1 U967 ( .A1(n1258), .A2(n1227), .A3(G110), .A4(n1263), .ZN(n1252) );
INV_X1 U968 ( .A(KEYINPUT2), .ZN(n1263) );
INV_X1 U969 ( .A(n1262), .ZN(n1258) );
NAND2_X1 U970 ( .A1(KEYINPUT2), .A2(n1264), .ZN(n1251) );
NAND2_X1 U971 ( .A1(n1227), .A2(n1265), .ZN(n1264) );
NAND2_X1 U972 ( .A1(G110), .A2(n1262), .ZN(n1265) );
XNOR2_X1 U973 ( .A(KEYINPUT53), .B(KEYINPUT30), .ZN(n1262) );
INV_X1 U974 ( .A(G122), .ZN(n1227) );
XOR2_X1 U975 ( .A(n1266), .B(G101), .Z(n1246) );
NAND2_X1 U976 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
XNOR2_X1 U977 ( .A(KEYINPUT6), .B(KEYINPUT36), .ZN(n1245) );
XOR2_X1 U978 ( .A(n1269), .B(n1270), .Z(n1208) );
XOR2_X1 U979 ( .A(KEYINPUT62), .B(G125), .Z(n1270) );
XOR2_X1 U980 ( .A(n1271), .B(n1272), .Z(n1269) );
AND2_X1 U981 ( .A1(n1120), .A2(G224), .ZN(n1272) );
XOR2_X1 U982 ( .A(n1167), .B(KEYINPUT12), .Z(n1240) );
NAND4_X1 U983 ( .A1(n1174), .A2(n1057), .A3(n1062), .A4(n1222), .ZN(n1167) );
NAND2_X1 U984 ( .A1(n1273), .A2(n1224), .ZN(n1222) );
NAND2_X1 U985 ( .A1(n1274), .A2(n1120), .ZN(n1224) );
INV_X1 U986 ( .A(n1036), .ZN(n1274) );
NAND2_X1 U987 ( .A1(G952), .A2(n1226), .ZN(n1036) );
NAND4_X1 U988 ( .A1(n1275), .A2(n1226), .A3(n1129), .A4(G953), .ZN(n1273) );
XOR2_X1 U989 ( .A(G898), .B(KEYINPUT28), .Z(n1129) );
NAND2_X1 U990 ( .A1(G237), .A2(n1276), .ZN(n1226) );
XOR2_X1 U991 ( .A(KEYINPUT59), .B(G902), .Z(n1275) );
INV_X1 U992 ( .A(n1196), .ZN(n1062) );
NAND2_X1 U993 ( .A1(n1065), .A2(n1064), .ZN(n1196) );
NAND2_X1 U994 ( .A1(n1277), .A2(n1278), .ZN(n1064) );
XNOR2_X1 U995 ( .A(G221), .B(KEYINPUT38), .ZN(n1277) );
XNOR2_X1 U996 ( .A(n1279), .B(G469), .ZN(n1065) );
NAND2_X1 U997 ( .A1(n1280), .A2(n1243), .ZN(n1279) );
XNOR2_X1 U998 ( .A(n1281), .B(n1154), .ZN(n1280) );
XNOR2_X1 U999 ( .A(n1282), .B(n1283), .ZN(n1154) );
XOR2_X1 U1000 ( .A(n1284), .B(n1285), .Z(n1283) );
AND2_X1 U1001 ( .A1(n1120), .A2(G227), .ZN(n1284) );
XOR2_X1 U1002 ( .A(n1212), .B(G110), .Z(n1282) );
NAND3_X1 U1003 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1281) );
NAND2_X1 U1004 ( .A1(n1099), .A2(n1289), .ZN(n1288) );
INV_X1 U1005 ( .A(KEYINPUT49), .ZN(n1289) );
NAND3_X1 U1006 ( .A1(KEYINPUT49), .A2(n1290), .A3(n1156), .ZN(n1287) );
OR2_X1 U1007 ( .A1(n1156), .A2(n1290), .ZN(n1286) );
NOR2_X1 U1008 ( .A1(KEYINPUT8), .A2(n1099), .ZN(n1290) );
XOR2_X1 U1009 ( .A(n1291), .B(n1292), .Z(n1099) );
XOR2_X1 U1010 ( .A(n1293), .B(G143), .Z(n1291) );
NAND2_X1 U1011 ( .A1(KEYINPUT24), .A2(n1209), .ZN(n1293) );
INV_X1 U1012 ( .A(G146), .ZN(n1209) );
XOR2_X1 U1013 ( .A(n1221), .B(n1250), .Z(n1156) );
XOR2_X1 U1014 ( .A(G107), .B(G104), .Z(n1250) );
INV_X1 U1015 ( .A(G101), .ZN(n1221) );
NOR2_X1 U1016 ( .A1(n1075), .A2(n1235), .ZN(n1057) );
XOR2_X1 U1017 ( .A(n1071), .B(KEYINPUT14), .Z(n1235) );
XOR2_X1 U1018 ( .A(n1134), .B(n1294), .Z(n1071) );
NOR2_X1 U1019 ( .A1(G902), .A2(n1133), .ZN(n1294) );
XNOR2_X1 U1020 ( .A(n1295), .B(n1296), .ZN(n1133) );
XOR2_X1 U1021 ( .A(n1297), .B(n1298), .Z(n1296) );
AND2_X1 U1022 ( .A1(n1299), .A2(G221), .ZN(n1298) );
NOR2_X1 U1023 ( .A1(KEYINPUT20), .A2(n1300), .ZN(n1297) );
XOR2_X1 U1024 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1025 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U1026 ( .A(n1305), .B(n1306), .ZN(n1304) );
NOR2_X1 U1027 ( .A1(G110), .A2(KEYINPUT21), .ZN(n1306) );
NAND2_X1 U1028 ( .A1(KEYINPUT15), .A2(n1292), .ZN(n1305) );
NOR2_X1 U1029 ( .A1(KEYINPUT57), .A2(n1212), .ZN(n1303) );
XNOR2_X1 U1030 ( .A(G119), .B(n1307), .ZN(n1301) );
XOR2_X1 U1031 ( .A(G146), .B(G125), .Z(n1307) );
NAND2_X1 U1032 ( .A1(KEYINPUT44), .A2(n1114), .ZN(n1295) );
INV_X1 U1033 ( .A(G137), .ZN(n1114) );
NAND2_X1 U1034 ( .A1(G217), .A2(n1278), .ZN(n1134) );
NAND2_X1 U1035 ( .A1(n1276), .A2(n1243), .ZN(n1278) );
XNOR2_X1 U1036 ( .A(G234), .B(KEYINPUT26), .ZN(n1276) );
XNOR2_X1 U1037 ( .A(n1308), .B(G472), .ZN(n1075) );
NAND2_X1 U1038 ( .A1(n1309), .A2(n1243), .ZN(n1308) );
XOR2_X1 U1039 ( .A(KEYINPUT51), .B(n1148), .Z(n1309) );
XNOR2_X1 U1040 ( .A(n1310), .B(n1311), .ZN(n1148) );
AND2_X1 U1041 ( .A1(n1312), .A2(G210), .ZN(n1311) );
XOR2_X1 U1042 ( .A(n1313), .B(G101), .Z(n1310) );
NAND2_X1 U1043 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NAND3_X1 U1044 ( .A1(n1316), .A2(n1268), .A3(n1317), .ZN(n1315) );
XNOR2_X1 U1045 ( .A(KEYINPUT5), .B(n1267), .ZN(n1317) );
XOR2_X1 U1046 ( .A(n1318), .B(n1271), .Z(n1316) );
NAND3_X1 U1047 ( .A1(n1319), .A2(n1320), .A3(n1321), .ZN(n1314) );
XOR2_X1 U1048 ( .A(n1271), .B(n1285), .Z(n1321) );
INV_X1 U1049 ( .A(n1318), .ZN(n1285) );
XOR2_X1 U1050 ( .A(n1106), .B(n1322), .Z(n1318) );
NOR2_X1 U1051 ( .A1(KEYINPUT23), .A2(n1323), .ZN(n1322) );
XOR2_X1 U1052 ( .A(G137), .B(G134), .Z(n1323) );
INV_X1 U1053 ( .A(G131), .ZN(n1106) );
XOR2_X1 U1054 ( .A(n1292), .B(n1324), .Z(n1271) );
XNOR2_X1 U1055 ( .A(n1325), .B(KEYINPUT55), .ZN(n1324) );
NAND2_X1 U1056 ( .A1(KEYINPUT39), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1057 ( .A(G146), .B(n1327), .Z(n1326) );
NOR2_X1 U1058 ( .A1(KEYINPUT13), .A2(n1211), .ZN(n1327) );
INV_X1 U1059 ( .A(G143), .ZN(n1211) );
OR2_X1 U1060 ( .A1(n1267), .A2(KEYINPUT5), .ZN(n1320) );
NAND3_X1 U1061 ( .A1(n1268), .A2(n1267), .A3(KEYINPUT5), .ZN(n1319) );
NAND2_X1 U1062 ( .A1(n1328), .A2(n1237), .ZN(n1267) );
XNOR2_X1 U1063 ( .A(G116), .B(G119), .ZN(n1328) );
NAND2_X1 U1064 ( .A1(G113), .A2(n1329), .ZN(n1268) );
XOR2_X1 U1065 ( .A(G119), .B(G116), .Z(n1329) );
INV_X1 U1066 ( .A(n1040), .ZN(n1174) );
NAND2_X1 U1067 ( .A1(n1232), .A2(n1231), .ZN(n1040) );
XNOR2_X1 U1068 ( .A(n1088), .B(n1330), .ZN(n1231) );
XOR2_X1 U1069 ( .A(KEYINPUT31), .B(G475), .Z(n1330) );
NOR2_X1 U1070 ( .A1(n1144), .A2(G902), .ZN(n1088) );
XNOR2_X1 U1071 ( .A(n1331), .B(n1332), .ZN(n1144) );
NOR2_X1 U1072 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
AND2_X1 U1073 ( .A1(KEYINPUT11), .A2(n1335), .ZN(n1334) );
NOR2_X1 U1074 ( .A1(KEYINPUT25), .A2(n1335), .ZN(n1333) );
XOR2_X1 U1075 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1076 ( .A(G143), .B(G131), .Z(n1337) );
XOR2_X1 U1077 ( .A(n1338), .B(n1339), .Z(n1336) );
NOR2_X1 U1078 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
XOR2_X1 U1079 ( .A(KEYINPUT40), .B(n1342), .Z(n1341) );
NOR2_X1 U1080 ( .A1(G146), .A2(n1343), .ZN(n1342) );
AND2_X1 U1081 ( .A1(n1343), .A2(G146), .ZN(n1340) );
XNOR2_X1 U1082 ( .A(n1095), .B(KEYINPUT52), .ZN(n1343) );
XOR2_X1 U1083 ( .A(G125), .B(n1212), .Z(n1095) );
INV_X1 U1084 ( .A(G140), .ZN(n1212) );
NAND2_X1 U1085 ( .A1(G214), .A2(n1312), .ZN(n1338) );
NOR2_X1 U1086 ( .A1(G953), .A2(G237), .ZN(n1312) );
NAND2_X1 U1087 ( .A1(n1344), .A2(n1345), .ZN(n1331) );
NAND2_X1 U1088 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
XOR2_X1 U1089 ( .A(KEYINPUT46), .B(G104), .Z(n1347) );
XOR2_X1 U1090 ( .A(n1237), .B(G122), .Z(n1346) );
INV_X1 U1091 ( .A(G113), .ZN(n1237) );
NAND2_X1 U1092 ( .A1(n1348), .A2(n1349), .ZN(n1344) );
XOR2_X1 U1093 ( .A(KEYINPUT22), .B(G104), .Z(n1349) );
XOR2_X1 U1094 ( .A(G122), .B(G113), .Z(n1348) );
XOR2_X1 U1095 ( .A(n1350), .B(G478), .Z(n1232) );
NAND2_X1 U1096 ( .A1(n1351), .A2(n1243), .ZN(n1350) );
INV_X1 U1097 ( .A(G902), .ZN(n1243) );
XOR2_X1 U1098 ( .A(n1137), .B(KEYINPUT19), .Z(n1351) );
XOR2_X1 U1099 ( .A(n1352), .B(n1353), .Z(n1137) );
XOR2_X1 U1100 ( .A(n1354), .B(n1355), .Z(n1353) );
XOR2_X1 U1101 ( .A(G122), .B(G116), .Z(n1355) );
XOR2_X1 U1102 ( .A(G143), .B(G134), .Z(n1354) );
XNOR2_X1 U1103 ( .A(n1356), .B(n1292), .ZN(n1352) );
XNOR2_X1 U1104 ( .A(G128), .B(KEYINPUT34), .ZN(n1292) );
XOR2_X1 U1105 ( .A(n1357), .B(G107), .Z(n1356) );
NAND2_X1 U1106 ( .A1(G217), .A2(n1299), .ZN(n1357) );
AND2_X1 U1107 ( .A1(G234), .A2(n1120), .ZN(n1299) );
INV_X1 U1108 ( .A(G953), .ZN(n1120) );
INV_X1 U1109 ( .A(G110), .ZN(n1238) );
endmodule


