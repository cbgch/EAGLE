//Key = 0010010100001111001101111001111011000101111111111001111101010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384;

XNOR2_X1 U748 ( .A(G107), .B(n1050), .ZN(G9) );
NAND4_X1 U749 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1050) );
NOR2_X1 U750 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XOR2_X1 U751 ( .A(KEYINPUT0), .B(n1057), .Z(n1051) );
NOR2_X1 U752 ( .A1(n1058), .A2(n1059), .ZN(G75) );
NOR4_X1 U753 ( .A1(n1060), .A2(n1061), .A3(G953), .A4(n1062), .ZN(n1059) );
NOR3_X1 U754 ( .A1(n1056), .A2(KEYINPUT59), .A3(n1063), .ZN(n1061) );
NOR2_X1 U755 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND3_X1 U756 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1060) );
NAND3_X1 U757 ( .A1(n1069), .A2(n1057), .A3(n1070), .ZN(n1067) );
INV_X1 U758 ( .A(n1065), .ZN(n1070) );
NAND3_X1 U759 ( .A1(n1071), .A2(n1053), .A3(n1072), .ZN(n1065) );
NAND3_X1 U760 ( .A1(n1073), .A2(n1074), .A3(n1072), .ZN(n1066) );
INV_X1 U761 ( .A(n1075), .ZN(n1072) );
NAND2_X1 U762 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NAND4_X1 U763 ( .A1(n1071), .A2(n1053), .A3(n1078), .A4(n1079), .ZN(n1077) );
NAND2_X1 U764 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND4_X1 U765 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1078) );
NAND2_X1 U766 ( .A1(KEYINPUT59), .A2(n1086), .ZN(n1084) );
OR2_X1 U767 ( .A1(n1081), .A2(KEYINPUT2), .ZN(n1083) );
NAND3_X1 U768 ( .A1(n1087), .A2(n1088), .A3(KEYINPUT2), .ZN(n1082) );
NAND3_X1 U769 ( .A1(n1089), .A2(n1090), .A3(n1085), .ZN(n1076) );
NAND2_X1 U770 ( .A1(n1091), .A2(n1081), .ZN(n1090) );
INV_X1 U771 ( .A(n1069), .ZN(n1081) );
NAND3_X1 U772 ( .A1(n1053), .A2(n1092), .A3(n1093), .ZN(n1091) );
INV_X1 U773 ( .A(KEYINPUT46), .ZN(n1092) );
NAND4_X1 U774 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1069), .ZN(n1089) );
NAND2_X1 U775 ( .A1(n1053), .A2(n1097), .ZN(n1096) );
NAND2_X1 U776 ( .A1(n1055), .A2(n1098), .ZN(n1097) );
NAND2_X1 U777 ( .A1(KEYINPUT46), .A2(n1093), .ZN(n1098) );
NAND2_X1 U778 ( .A1(n1071), .A2(n1099), .ZN(n1095) );
NAND2_X1 U779 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U780 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
OR3_X1 U781 ( .A1(n1103), .A2(n1104), .A3(n1071), .ZN(n1094) );
INV_X1 U782 ( .A(KEYINPUT6), .ZN(n1103) );
NOR3_X1 U783 ( .A1(n1062), .A2(G953), .A3(G952), .ZN(n1058) );
AND4_X1 U784 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1062) );
NOR4_X1 U785 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1108) );
XOR2_X1 U786 ( .A(n1113), .B(n1114), .Z(n1112) );
XNOR2_X1 U787 ( .A(KEYINPUT28), .B(n1115), .ZN(n1114) );
NAND2_X1 U788 ( .A1(KEYINPUT39), .A2(n1116), .ZN(n1113) );
XNOR2_X1 U789 ( .A(n1117), .B(KEYINPUT13), .ZN(n1111) );
XOR2_X1 U790 ( .A(n1118), .B(n1119), .Z(n1110) );
NAND3_X1 U791 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1109) );
XNOR2_X1 U792 ( .A(n1123), .B(G472), .ZN(n1122) );
NAND2_X1 U793 ( .A1(n1124), .A2(n1125), .ZN(n1121) );
INV_X1 U794 ( .A(KEYINPUT24), .ZN(n1125) );
NAND2_X1 U795 ( .A1(n1126), .A2(n1127), .ZN(n1124) );
XNOR2_X1 U796 ( .A(n1128), .B(KEYINPUT10), .ZN(n1126) );
NAND2_X1 U797 ( .A1(KEYINPUT24), .A2(n1129), .ZN(n1120) );
NAND2_X1 U798 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
OR3_X1 U799 ( .A1(n1132), .A2(n1128), .A3(KEYINPUT10), .ZN(n1131) );
NAND2_X1 U800 ( .A1(KEYINPUT10), .A2(n1128), .ZN(n1130) );
NOR3_X1 U801 ( .A1(n1080), .A2(n1133), .A3(n1087), .ZN(n1107) );
NAND2_X1 U802 ( .A1(n1128), .A2(n1132), .ZN(n1106) );
INV_X1 U803 ( .A(n1134), .ZN(n1128) );
XOR2_X1 U804 ( .A(G469), .B(n1135), .Z(n1105) );
NOR2_X1 U805 ( .A1(n1136), .A2(KEYINPUT58), .ZN(n1135) );
XOR2_X1 U806 ( .A(n1137), .B(n1138), .Z(G72) );
XOR2_X1 U807 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U808 ( .A1(G953), .A2(n1141), .ZN(n1140) );
NAND2_X1 U809 ( .A1(G900), .A2(G227), .ZN(n1141) );
NAND2_X1 U810 ( .A1(n1142), .A2(n1143), .ZN(n1139) );
NAND2_X1 U811 ( .A1(G953), .A2(n1144), .ZN(n1143) );
XOR2_X1 U812 ( .A(n1145), .B(n1146), .Z(n1142) );
XOR2_X1 U813 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U814 ( .A(G137), .B(n1149), .ZN(n1145) );
NAND2_X1 U815 ( .A1(KEYINPUT18), .A2(n1150), .ZN(n1149) );
NOR2_X1 U816 ( .A1(n1151), .A2(G953), .ZN(n1137) );
XOR2_X1 U817 ( .A(n1152), .B(n1153), .Z(G69) );
NOR2_X1 U818 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NOR2_X1 U819 ( .A1(n1156), .A2(n1157), .ZN(n1154) );
NAND2_X1 U820 ( .A1(n1158), .A2(n1159), .ZN(n1152) );
NAND2_X1 U821 ( .A1(n1160), .A2(n1155), .ZN(n1159) );
XNOR2_X1 U822 ( .A(n1161), .B(n1162), .ZN(n1160) );
NOR2_X1 U823 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NAND3_X1 U824 ( .A1(G898), .A2(n1161), .A3(G953), .ZN(n1158) );
NOR2_X1 U825 ( .A1(n1165), .A2(n1166), .ZN(G66) );
XOR2_X1 U826 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U827 ( .A(n1169), .B(KEYINPUT5), .Z(n1168) );
OR2_X1 U828 ( .A1(n1170), .A2(n1119), .ZN(n1169) );
NAND2_X1 U829 ( .A1(KEYINPUT27), .A2(n1171), .ZN(n1167) );
NOR3_X1 U830 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(G63) );
AND3_X1 U831 ( .A1(KEYINPUT1), .A2(G953), .A3(G952), .ZN(n1174) );
NOR2_X1 U832 ( .A1(KEYINPUT1), .A2(n1175), .ZN(n1173) );
INV_X1 U833 ( .A(n1165), .ZN(n1175) );
NOR3_X1 U834 ( .A1(n1116), .A2(n1176), .A3(n1177), .ZN(n1172) );
NOR3_X1 U835 ( .A1(n1178), .A2(n1115), .A3(n1170), .ZN(n1177) );
NOR2_X1 U836 ( .A1(n1179), .A2(n1180), .ZN(n1176) );
NOR2_X1 U837 ( .A1(n1068), .A2(n1115), .ZN(n1180) );
NOR2_X1 U838 ( .A1(n1165), .A2(n1181), .ZN(G60) );
NOR2_X1 U839 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
XOR2_X1 U840 ( .A(n1184), .B(n1185), .Z(n1183) );
AND2_X1 U841 ( .A1(n1186), .A2(KEYINPUT29), .ZN(n1185) );
AND2_X1 U842 ( .A1(G475), .A2(n1187), .ZN(n1184) );
NOR2_X1 U843 ( .A1(KEYINPUT29), .A2(n1186), .ZN(n1182) );
XNOR2_X1 U844 ( .A(G104), .B(n1188), .ZN(G6) );
NOR2_X1 U845 ( .A1(n1165), .A2(n1189), .ZN(G57) );
XOR2_X1 U846 ( .A(n1190), .B(n1191), .Z(n1189) );
NOR2_X1 U847 ( .A1(KEYINPUT16), .A2(n1192), .ZN(n1191) );
XOR2_X1 U848 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U849 ( .A(n1195), .B(n1196), .Z(n1193) );
AND2_X1 U850 ( .A1(G472), .A2(n1187), .ZN(n1196) );
NAND3_X1 U851 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1190) );
OR2_X1 U852 ( .A1(n1200), .A2(KEYINPUT14), .ZN(n1199) );
OR3_X1 U853 ( .A1(n1201), .A2(n1202), .A3(G101), .ZN(n1198) );
INV_X1 U854 ( .A(KEYINPUT14), .ZN(n1201) );
NAND2_X1 U855 ( .A1(G101), .A2(n1202), .ZN(n1197) );
NAND2_X1 U856 ( .A1(KEYINPUT44), .A2(n1200), .ZN(n1202) );
NOR2_X1 U857 ( .A1(n1165), .A2(n1203), .ZN(G54) );
XOR2_X1 U858 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U859 ( .A(n1206), .B(n1207), .Z(n1205) );
NOR2_X1 U860 ( .A1(n1208), .A2(n1209), .ZN(n1206) );
XOR2_X1 U861 ( .A(n1210), .B(KEYINPUT43), .Z(n1209) );
NAND2_X1 U862 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NOR2_X1 U863 ( .A1(n1212), .A2(n1211), .ZN(n1208) );
XNOR2_X1 U864 ( .A(G140), .B(n1213), .ZN(n1211) );
NOR2_X1 U865 ( .A1(KEYINPUT25), .A2(n1214), .ZN(n1213) );
XOR2_X1 U866 ( .A(KEYINPUT22), .B(n1215), .Z(n1204) );
AND2_X1 U867 ( .A1(G469), .A2(n1187), .ZN(n1215) );
NOR2_X1 U868 ( .A1(n1165), .A2(n1216), .ZN(G51) );
XOR2_X1 U869 ( .A(n1217), .B(n1218), .Z(n1216) );
XOR2_X1 U870 ( .A(n1219), .B(n1220), .Z(n1218) );
NOR2_X1 U871 ( .A1(n1134), .A2(n1170), .ZN(n1220) );
INV_X1 U872 ( .A(n1187), .ZN(n1170) );
NOR2_X1 U873 ( .A1(n1221), .A2(n1068), .ZN(n1187) );
AND3_X1 U874 ( .A1(n1222), .A2(n1223), .A3(n1151), .ZN(n1068) );
AND4_X1 U875 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1151) );
NOR4_X1 U876 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1227) );
INV_X1 U877 ( .A(n1232), .ZN(n1231) );
NAND3_X1 U878 ( .A1(n1233), .A2(n1234), .A3(n1102), .ZN(n1226) );
NAND2_X1 U879 ( .A1(n1055), .A2(n1235), .ZN(n1234) );
XNOR2_X1 U880 ( .A(KEYINPUT20), .B(n1163), .ZN(n1223) );
NAND4_X1 U881 ( .A1(n1236), .A2(n1237), .A3(n1188), .A4(n1238), .ZN(n1163) );
NAND4_X1 U882 ( .A1(n1093), .A2(n1239), .A3(n1053), .A4(n1052), .ZN(n1188) );
NAND4_X1 U883 ( .A1(n1239), .A2(n1240), .A3(n1053), .A4(n1052), .ZN(n1237) );
OR2_X1 U884 ( .A1(n1241), .A2(n1056), .ZN(n1236) );
INV_X1 U885 ( .A(n1164), .ZN(n1222) );
NAND4_X1 U886 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1164) );
NOR2_X1 U887 ( .A1(n1155), .A2(G952), .ZN(n1165) );
XNOR2_X1 U888 ( .A(G146), .B(n1225), .ZN(G48) );
NAND3_X1 U889 ( .A1(n1246), .A2(n1247), .A3(n1093), .ZN(n1225) );
XNOR2_X1 U890 ( .A(G143), .B(n1232), .ZN(G45) );
NAND4_X1 U891 ( .A1(n1102), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1232) );
XNOR2_X1 U892 ( .A(n1250), .B(n1230), .ZN(G42) );
NOR3_X1 U893 ( .A1(n1100), .A2(n1251), .A3(n1235), .ZN(n1230) );
XNOR2_X1 U894 ( .A(n1252), .B(n1229), .ZN(G39) );
AND3_X1 U895 ( .A1(n1233), .A2(n1246), .A3(n1071), .ZN(n1229) );
INV_X1 U896 ( .A(n1251), .ZN(n1233) );
XOR2_X1 U897 ( .A(n1253), .B(n1254), .Z(G36) );
NOR3_X1 U898 ( .A1(n1255), .A2(n1055), .A3(n1251), .ZN(n1254) );
NAND3_X1 U899 ( .A1(n1057), .A2(n1256), .A3(n1069), .ZN(n1251) );
XNOR2_X1 U900 ( .A(KEYINPUT45), .B(n1104), .ZN(n1255) );
XNOR2_X1 U901 ( .A(G134), .B(KEYINPUT15), .ZN(n1253) );
NAND2_X1 U902 ( .A1(n1257), .A2(n1258), .ZN(G33) );
NAND2_X1 U903 ( .A1(G131), .A2(n1259), .ZN(n1258) );
XOR2_X1 U904 ( .A(n1260), .B(KEYINPUT31), .Z(n1257) );
OR2_X1 U905 ( .A1(n1259), .A2(G131), .ZN(n1260) );
NAND4_X1 U906 ( .A1(n1057), .A2(n1261), .A3(n1069), .A4(n1262), .ZN(n1259) );
NOR2_X1 U907 ( .A1(n1235), .A2(n1104), .ZN(n1262) );
NOR2_X1 U908 ( .A1(n1263), .A2(n1087), .ZN(n1069) );
XNOR2_X1 U909 ( .A(KEYINPUT47), .B(n1256), .ZN(n1261) );
XNOR2_X1 U910 ( .A(n1228), .B(n1264), .ZN(G30) );
XNOR2_X1 U911 ( .A(KEYINPUT12), .B(n1265), .ZN(n1264) );
AND3_X1 U912 ( .A1(n1247), .A2(n1240), .A3(n1246), .ZN(n1228) );
AND2_X1 U913 ( .A1(n1239), .A2(n1256), .ZN(n1247) );
XNOR2_X1 U914 ( .A(G101), .B(n1238), .ZN(G3) );
NAND4_X1 U915 ( .A1(n1102), .A2(n1071), .A3(n1239), .A4(n1052), .ZN(n1238) );
AND2_X1 U916 ( .A1(n1086), .A2(n1057), .ZN(n1239) );
XOR2_X1 U917 ( .A(n1266), .B(G125), .Z(G27) );
NAND2_X1 U918 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
OR2_X1 U919 ( .A1(n1224), .A2(KEYINPUT36), .ZN(n1268) );
NAND2_X1 U920 ( .A1(n1269), .A2(n1093), .ZN(n1224) );
NAND3_X1 U921 ( .A1(n1269), .A2(n1235), .A3(KEYINPUT36), .ZN(n1267) );
INV_X1 U922 ( .A(n1093), .ZN(n1235) );
NOR4_X1 U923 ( .A1(n1064), .A2(n1100), .A3(n1056), .A4(n1270), .ZN(n1269) );
INV_X1 U924 ( .A(n1256), .ZN(n1270) );
NAND2_X1 U925 ( .A1(n1075), .A2(n1271), .ZN(n1256) );
NAND4_X1 U926 ( .A1(G953), .A2(G902), .A3(n1272), .A4(n1144), .ZN(n1271) );
INV_X1 U927 ( .A(G900), .ZN(n1144) );
INV_X1 U928 ( .A(n1273), .ZN(n1100) );
XNOR2_X1 U929 ( .A(G122), .B(n1242), .ZN(G24) );
NAND4_X1 U930 ( .A1(n1274), .A2(n1053), .A3(n1248), .A4(n1249), .ZN(n1242) );
NOR2_X1 U931 ( .A1(n1275), .A2(n1276), .ZN(n1053) );
XOR2_X1 U932 ( .A(n1243), .B(n1277), .Z(G21) );
NAND2_X1 U933 ( .A1(KEYINPUT51), .A2(G119), .ZN(n1277) );
NAND3_X1 U934 ( .A1(n1071), .A2(n1246), .A3(n1274), .ZN(n1243) );
NOR2_X1 U935 ( .A1(n1278), .A2(n1279), .ZN(n1246) );
XNOR2_X1 U936 ( .A(n1244), .B(n1280), .ZN(G18) );
XOR2_X1 U937 ( .A(KEYINPUT56), .B(G116), .Z(n1280) );
NAND3_X1 U938 ( .A1(n1102), .A2(n1240), .A3(n1274), .ZN(n1244) );
INV_X1 U939 ( .A(n1055), .ZN(n1240) );
NAND2_X1 U940 ( .A1(n1281), .A2(n1248), .ZN(n1055) );
XNOR2_X1 U941 ( .A(G113), .B(n1245), .ZN(G15) );
NAND3_X1 U942 ( .A1(n1102), .A2(n1093), .A3(n1274), .ZN(n1245) );
NOR3_X1 U943 ( .A1(n1056), .A2(n1282), .A3(n1064), .ZN(n1274) );
NAND2_X1 U944 ( .A1(n1073), .A2(n1085), .ZN(n1064) );
INV_X1 U945 ( .A(n1052), .ZN(n1282) );
INV_X1 U946 ( .A(n1086), .ZN(n1056) );
NOR2_X1 U947 ( .A1(n1248), .A2(n1281), .ZN(n1093) );
INV_X1 U948 ( .A(n1104), .ZN(n1102) );
NAND2_X1 U949 ( .A1(n1275), .A2(n1283), .ZN(n1104) );
XNOR2_X1 U950 ( .A(KEYINPUT34), .B(n1276), .ZN(n1283) );
INV_X1 U951 ( .A(n1278), .ZN(n1276) );
XNOR2_X1 U952 ( .A(G110), .B(n1284), .ZN(G12) );
NAND2_X1 U953 ( .A1(n1285), .A2(n1086), .ZN(n1284) );
NOR2_X1 U954 ( .A1(n1088), .A2(n1087), .ZN(n1086) );
AND2_X1 U955 ( .A1(G214), .A2(n1286), .ZN(n1087) );
INV_X1 U956 ( .A(n1263), .ZN(n1088) );
XNOR2_X1 U957 ( .A(n1127), .B(n1134), .ZN(n1263) );
NAND2_X1 U958 ( .A1(G210), .A2(n1286), .ZN(n1134) );
NAND2_X1 U959 ( .A1(n1287), .A2(n1221), .ZN(n1286) );
XOR2_X1 U960 ( .A(KEYINPUT7), .B(G237), .Z(n1287) );
INV_X1 U961 ( .A(n1132), .ZN(n1127) );
NAND2_X1 U962 ( .A1(n1288), .A2(n1221), .ZN(n1132) );
XOR2_X1 U963 ( .A(n1289), .B(n1217), .Z(n1288) );
XNOR2_X1 U964 ( .A(n1290), .B(n1161), .ZN(n1217) );
XNOR2_X1 U965 ( .A(n1291), .B(n1292), .ZN(n1161) );
XNOR2_X1 U966 ( .A(n1293), .B(n1294), .ZN(n1292) );
XOR2_X1 U967 ( .A(KEYINPUT42), .B(G116), .Z(n1294) );
INV_X1 U968 ( .A(G107), .ZN(n1293) );
XOR2_X1 U969 ( .A(n1295), .B(n1296), .Z(n1291) );
XNOR2_X1 U970 ( .A(G101), .B(n1297), .ZN(n1295) );
XOR2_X1 U971 ( .A(n1298), .B(G125), .Z(n1290) );
NAND2_X1 U972 ( .A1(KEYINPUT40), .A2(n1219), .ZN(n1289) );
NOR2_X1 U973 ( .A1(n1156), .A2(G953), .ZN(n1219) );
INV_X1 U974 ( .A(G224), .ZN(n1156) );
XOR2_X1 U975 ( .A(n1241), .B(KEYINPUT53), .Z(n1285) );
NAND4_X1 U976 ( .A1(n1273), .A2(n1071), .A3(n1057), .A4(n1052), .ZN(n1241) );
NAND2_X1 U977 ( .A1(n1075), .A2(n1299), .ZN(n1052) );
NAND4_X1 U978 ( .A1(G953), .A2(G902), .A3(n1272), .A4(n1157), .ZN(n1299) );
INV_X1 U979 ( .A(G898), .ZN(n1157) );
NAND3_X1 U980 ( .A1(n1272), .A2(n1155), .A3(n1300), .ZN(n1075) );
XOR2_X1 U981 ( .A(KEYINPUT62), .B(G952), .Z(n1300) );
NAND2_X1 U982 ( .A1(G234), .A2(G237), .ZN(n1272) );
NOR2_X1 U983 ( .A1(n1073), .A2(n1080), .ZN(n1057) );
INV_X1 U984 ( .A(n1085), .ZN(n1080) );
NAND2_X1 U985 ( .A1(G221), .A2(n1301), .ZN(n1085) );
XNOR2_X1 U986 ( .A(n1136), .B(G469), .ZN(n1073) );
AND2_X1 U987 ( .A1(n1302), .A2(n1221), .ZN(n1136) );
XOR2_X1 U988 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U989 ( .A(n1214), .B(n1305), .ZN(n1304) );
XNOR2_X1 U990 ( .A(KEYINPUT4), .B(n1250), .ZN(n1305) );
XNOR2_X1 U991 ( .A(n1207), .B(n1212), .ZN(n1303) );
AND2_X1 U992 ( .A1(G227), .A2(n1155), .ZN(n1212) );
XNOR2_X1 U993 ( .A(n1306), .B(n1307), .ZN(n1207) );
XNOR2_X1 U994 ( .A(n1147), .B(n1308), .ZN(n1307) );
XOR2_X1 U995 ( .A(n1309), .B(n1310), .Z(n1147) );
XNOR2_X1 U996 ( .A(G143), .B(G146), .ZN(n1309) );
XOR2_X1 U997 ( .A(n1311), .B(n1312), .Z(n1306) );
XOR2_X1 U998 ( .A(KEYINPUT61), .B(KEYINPUT35), .Z(n1312) );
NAND2_X1 U999 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
NAND2_X1 U1000 ( .A1(G101), .A2(n1315), .ZN(n1314) );
XOR2_X1 U1001 ( .A(KEYINPUT37), .B(n1316), .Z(n1313) );
NOR2_X1 U1002 ( .A1(G101), .A2(n1315), .ZN(n1316) );
NAND2_X1 U1003 ( .A1(n1317), .A2(n1318), .ZN(n1315) );
NAND2_X1 U1004 ( .A1(n1319), .A2(G107), .ZN(n1318) );
XOR2_X1 U1005 ( .A(KEYINPUT55), .B(n1320), .Z(n1317) );
NOR2_X1 U1006 ( .A1(G107), .A2(n1319), .ZN(n1320) );
XNOR2_X1 U1007 ( .A(KEYINPUT3), .B(G104), .ZN(n1319) );
NOR2_X1 U1008 ( .A1(n1248), .A2(n1249), .ZN(n1071) );
INV_X1 U1009 ( .A(n1281), .ZN(n1249) );
NOR2_X1 U1010 ( .A1(n1117), .A2(n1133), .ZN(n1281) );
NOR3_X1 U1011 ( .A1(G475), .A2(G902), .A3(n1321), .ZN(n1133) );
INV_X1 U1012 ( .A(n1186), .ZN(n1321) );
AND2_X1 U1013 ( .A1(G475), .A2(n1322), .ZN(n1117) );
NAND2_X1 U1014 ( .A1(n1186), .A2(n1221), .ZN(n1322) );
XNOR2_X1 U1015 ( .A(n1323), .B(n1324), .ZN(n1186) );
XOR2_X1 U1016 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1017 ( .A(G125), .B(n1327), .Z(n1326) );
NOR3_X1 U1018 ( .A1(n1328), .A2(G953), .A3(G237), .ZN(n1327) );
INV_X1 U1019 ( .A(G214), .ZN(n1328) );
XNOR2_X1 U1020 ( .A(n1329), .B(G131), .ZN(n1325) );
XNOR2_X1 U1021 ( .A(n1296), .B(n1330), .ZN(n1323) );
XNOR2_X1 U1022 ( .A(n1331), .B(n1332), .ZN(n1330) );
NOR2_X1 U1023 ( .A1(G140), .A2(KEYINPUT17), .ZN(n1332) );
NAND2_X1 U1024 ( .A1(KEYINPUT23), .A2(n1333), .ZN(n1331) );
XOR2_X1 U1025 ( .A(G104), .B(n1334), .Z(n1296) );
XNOR2_X1 U1026 ( .A(n1335), .B(G113), .ZN(n1334) );
XNOR2_X1 U1027 ( .A(n1116), .B(n1115), .ZN(n1248) );
INV_X1 U1028 ( .A(G478), .ZN(n1115) );
NOR2_X1 U1029 ( .A1(n1179), .A2(G902), .ZN(n1116) );
INV_X1 U1030 ( .A(n1178), .ZN(n1179) );
NAND2_X1 U1031 ( .A1(n1336), .A2(n1337), .ZN(n1178) );
NAND2_X1 U1032 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
XOR2_X1 U1033 ( .A(n1340), .B(n1341), .Z(n1336) );
NOR2_X1 U1034 ( .A1(n1338), .A2(n1339), .ZN(n1341) );
INV_X1 U1035 ( .A(KEYINPUT33), .ZN(n1339) );
XNOR2_X1 U1036 ( .A(n1342), .B(n1343), .ZN(n1338) );
XNOR2_X1 U1037 ( .A(n1344), .B(n1345), .ZN(n1343) );
NOR2_X1 U1038 ( .A1(KEYINPUT60), .A2(n1346), .ZN(n1345) );
XNOR2_X1 U1039 ( .A(G116), .B(n1347), .ZN(n1346) );
NOR2_X1 U1040 ( .A1(KEYINPUT26), .A2(n1335), .ZN(n1347) );
INV_X1 U1041 ( .A(G122), .ZN(n1335) );
NAND2_X1 U1042 ( .A1(KEYINPUT19), .A2(n1265), .ZN(n1344) );
INV_X1 U1043 ( .A(G128), .ZN(n1265) );
XNOR2_X1 U1044 ( .A(G107), .B(n1348), .ZN(n1342) );
XNOR2_X1 U1045 ( .A(n1333), .B(G134), .ZN(n1348) );
INV_X1 U1046 ( .A(G143), .ZN(n1333) );
NAND2_X1 U1047 ( .A1(G217), .A2(n1349), .ZN(n1340) );
NOR2_X1 U1048 ( .A1(n1278), .A2(n1275), .ZN(n1273) );
INV_X1 U1049 ( .A(n1279), .ZN(n1275) );
XOR2_X1 U1050 ( .A(G472), .B(n1350), .Z(n1279) );
NOR2_X1 U1051 ( .A1(n1123), .A2(KEYINPUT38), .ZN(n1350) );
AND2_X1 U1052 ( .A1(n1351), .A2(n1221), .ZN(n1123) );
XOR2_X1 U1053 ( .A(n1352), .B(n1353), .Z(n1351) );
XOR2_X1 U1054 ( .A(n1354), .B(n1194), .Z(n1353) );
XNOR2_X1 U1055 ( .A(n1355), .B(n1356), .ZN(n1194) );
XOR2_X1 U1056 ( .A(KEYINPUT21), .B(G119), .Z(n1356) );
XNOR2_X1 U1057 ( .A(G113), .B(G116), .ZN(n1355) );
NAND2_X1 U1058 ( .A1(KEYINPUT41), .A2(n1200), .ZN(n1354) );
NOR3_X1 U1059 ( .A1(G237), .A2(G953), .A3(n1357), .ZN(n1200) );
INV_X1 U1060 ( .A(G210), .ZN(n1357) );
XOR2_X1 U1061 ( .A(n1358), .B(G101), .Z(n1352) );
NAND2_X1 U1062 ( .A1(KEYINPUT52), .A2(n1195), .ZN(n1358) );
XNOR2_X1 U1063 ( .A(n1298), .B(n1308), .ZN(n1195) );
NAND2_X1 U1064 ( .A1(n1359), .A2(n1360), .ZN(n1308) );
NAND2_X1 U1065 ( .A1(n1148), .A2(G137), .ZN(n1360) );
NAND2_X1 U1066 ( .A1(n1361), .A2(n1252), .ZN(n1359) );
XNOR2_X1 U1067 ( .A(n1148), .B(KEYINPUT50), .ZN(n1361) );
XOR2_X1 U1068 ( .A(G134), .B(G131), .Z(n1148) );
NAND3_X1 U1069 ( .A1(n1362), .A2(n1363), .A3(n1364), .ZN(n1298) );
OR2_X1 U1070 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
NAND3_X1 U1071 ( .A1(n1366), .A2(n1365), .A3(n1367), .ZN(n1363) );
NAND2_X1 U1072 ( .A1(n1310), .A2(n1368), .ZN(n1362) );
NAND2_X1 U1073 ( .A1(n1369), .A2(n1365), .ZN(n1368) );
INV_X1 U1074 ( .A(KEYINPUT8), .ZN(n1365) );
XNOR2_X1 U1075 ( .A(n1366), .B(KEYINPUT54), .ZN(n1369) );
XOR2_X1 U1076 ( .A(G143), .B(n1370), .Z(n1366) );
NOR2_X1 U1077 ( .A1(KEYINPUT63), .A2(n1329), .ZN(n1370) );
INV_X1 U1078 ( .A(n1367), .ZN(n1310) );
XOR2_X1 U1079 ( .A(G128), .B(KEYINPUT11), .Z(n1367) );
XOR2_X1 U1080 ( .A(n1371), .B(n1118), .Z(n1278) );
NAND2_X1 U1081 ( .A1(n1171), .A2(n1372), .ZN(n1118) );
XNOR2_X1 U1082 ( .A(KEYINPUT48), .B(n1221), .ZN(n1372) );
XOR2_X1 U1083 ( .A(n1373), .B(n1374), .Z(n1171) );
XNOR2_X1 U1084 ( .A(n1297), .B(n1375), .ZN(n1374) );
XOR2_X1 U1085 ( .A(n1376), .B(n1377), .Z(n1375) );
AND2_X1 U1086 ( .A1(n1349), .A2(G221), .ZN(n1377) );
AND2_X1 U1087 ( .A1(G234), .A2(n1155), .ZN(n1349) );
INV_X1 U1088 ( .A(G953), .ZN(n1155) );
NAND2_X1 U1089 ( .A1(n1378), .A2(n1379), .ZN(n1376) );
NAND2_X1 U1090 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
XNOR2_X1 U1091 ( .A(KEYINPUT30), .B(n1329), .ZN(n1381) );
INV_X1 U1092 ( .A(G146), .ZN(n1329) );
XOR2_X1 U1093 ( .A(n1150), .B(KEYINPUT49), .Z(n1380) );
NAND2_X1 U1094 ( .A1(n1382), .A2(n1383), .ZN(n1378) );
XNOR2_X1 U1095 ( .A(KEYINPUT9), .B(n1150), .ZN(n1383) );
XOR2_X1 U1096 ( .A(G125), .B(n1250), .Z(n1150) );
INV_X1 U1097 ( .A(G140), .ZN(n1250) );
XNOR2_X1 U1098 ( .A(KEYINPUT30), .B(G146), .ZN(n1382) );
XNOR2_X1 U1099 ( .A(G119), .B(n1214), .ZN(n1297) );
INV_X1 U1100 ( .A(G110), .ZN(n1214) );
XNOR2_X1 U1101 ( .A(G128), .B(n1384), .ZN(n1373) );
XNOR2_X1 U1102 ( .A(KEYINPUT57), .B(n1252), .ZN(n1384) );
INV_X1 U1103 ( .A(G137), .ZN(n1252) );
NAND2_X1 U1104 ( .A1(KEYINPUT32), .A2(n1119), .ZN(n1371) );
NAND2_X1 U1105 ( .A1(G217), .A2(n1301), .ZN(n1119) );
NAND2_X1 U1106 ( .A1(G234), .A2(n1221), .ZN(n1301) );
INV_X1 U1107 ( .A(G902), .ZN(n1221) );
endmodule


