//Key = 1000111110110100011101111111100110100010011011110111010011110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375;

XNOR2_X1 U750 ( .A(G107), .B(n1043), .ZN(G9) );
NOR2_X1 U751 ( .A1(n1044), .A2(n1045), .ZN(G75) );
NOR3_X1 U752 ( .A1(n1046), .A2(G953), .A3(n1047), .ZN(n1045) );
XOR2_X1 U753 ( .A(n1048), .B(KEYINPUT3), .Z(n1046) );
NAND3_X1 U754 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
INV_X1 U755 ( .A(n1052), .ZN(n1051) );
NAND3_X1 U756 ( .A1(n1053), .A2(n1054), .A3(KEYINPUT33), .ZN(n1050) );
NAND4_X1 U757 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NAND2_X1 U758 ( .A1(n1055), .A2(n1059), .ZN(n1049) );
NAND2_X1 U759 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND3_X1 U760 ( .A1(n1058), .A2(n1062), .A3(n1053), .ZN(n1061) );
NAND2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U762 ( .A1(n1056), .A2(n1065), .ZN(n1064) );
NAND2_X1 U763 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U764 ( .A1(n1057), .A2(n1068), .ZN(n1067) );
INV_X1 U765 ( .A(KEYINPUT33), .ZN(n1068) );
NAND2_X1 U766 ( .A1(n1069), .A2(n1070), .ZN(n1063) );
NAND2_X1 U767 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U768 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
INV_X1 U769 ( .A(n1075), .ZN(n1071) );
NAND3_X1 U770 ( .A1(n1069), .A2(n1076), .A3(n1056), .ZN(n1060) );
NAND2_X1 U771 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U772 ( .A1(n1053), .A2(n1079), .ZN(n1078) );
NAND2_X1 U773 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U774 ( .A1(n1058), .A2(n1082), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
INV_X1 U777 ( .A(n1087), .ZN(n1055) );
NOR3_X1 U778 ( .A1(n1047), .A2(G953), .A3(G952), .ZN(n1044) );
AND4_X1 U779 ( .A1(n1088), .A2(n1053), .A3(n1089), .A4(n1090), .ZN(n1047) );
NOR4_X1 U780 ( .A1(n1073), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1090) );
XNOR2_X1 U781 ( .A(n1094), .B(n1095), .ZN(n1092) );
XNOR2_X1 U782 ( .A(KEYINPUT57), .B(KEYINPUT55), .ZN(n1094) );
XOR2_X1 U783 ( .A(n1096), .B(n1097), .Z(n1091) );
XNOR2_X1 U784 ( .A(KEYINPUT17), .B(n1098), .ZN(n1097) );
XOR2_X1 U785 ( .A(n1099), .B(KEYINPUT6), .Z(n1089) );
NAND2_X1 U786 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U787 ( .A1(G478), .A2(n1102), .ZN(n1101) );
XOR2_X1 U788 ( .A(KEYINPUT38), .B(n1103), .Z(n1100) );
XOR2_X1 U789 ( .A(n1104), .B(n1105), .Z(G72) );
XOR2_X1 U790 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U791 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U792 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NAND3_X1 U793 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1106) );
NAND2_X1 U794 ( .A1(G953), .A2(n1111), .ZN(n1114) );
OR2_X1 U795 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NAND2_X1 U796 ( .A1(n1117), .A2(n1115), .ZN(n1112) );
NAND2_X1 U797 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U798 ( .A1(KEYINPUT34), .A2(n1116), .ZN(n1119) );
NAND2_X1 U799 ( .A1(KEYINPUT13), .A2(n1120), .ZN(n1116) );
NAND2_X1 U800 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
INV_X1 U801 ( .A(KEYINPUT34), .ZN(n1121) );
XNOR2_X1 U802 ( .A(n1122), .B(n1123), .ZN(n1120) );
XNOR2_X1 U803 ( .A(n1124), .B(KEYINPUT63), .ZN(n1123) );
NAND2_X1 U804 ( .A1(KEYINPUT21), .A2(n1125), .ZN(n1124) );
INV_X1 U805 ( .A(G134), .ZN(n1125) );
XOR2_X1 U806 ( .A(n1126), .B(n1127), .Z(n1122) );
NAND2_X1 U807 ( .A1(n1109), .A2(n1128), .ZN(n1104) );
NAND2_X1 U808 ( .A1(n1129), .A2(n1130), .ZN(G69) );
NAND2_X1 U809 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U810 ( .A1(G953), .A2(n1133), .ZN(n1132) );
NAND2_X1 U811 ( .A1(G898), .A2(G224), .ZN(n1133) );
NAND2_X1 U812 ( .A1(n1134), .A2(n1135), .ZN(n1129) );
NAND2_X1 U813 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
OR2_X1 U814 ( .A1(n1109), .A2(G224), .ZN(n1137) );
INV_X1 U815 ( .A(n1138), .ZN(n1136) );
INV_X1 U816 ( .A(n1131), .ZN(n1134) );
XNOR2_X1 U817 ( .A(n1139), .B(n1140), .ZN(n1131) );
NOR3_X1 U818 ( .A1(n1141), .A2(KEYINPUT20), .A3(n1138), .ZN(n1140) );
XNOR2_X1 U819 ( .A(n1142), .B(n1143), .ZN(n1141) );
NAND2_X1 U820 ( .A1(n1144), .A2(n1145), .ZN(n1139) );
NAND2_X1 U821 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XNOR2_X1 U822 ( .A(G953), .B(KEYINPUT60), .ZN(n1144) );
NOR2_X1 U823 ( .A1(n1148), .A2(n1149), .ZN(G66) );
XNOR2_X1 U824 ( .A(n1150), .B(n1151), .ZN(n1149) );
NOR2_X1 U825 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NOR2_X1 U826 ( .A1(n1148), .A2(n1154), .ZN(G63) );
XNOR2_X1 U827 ( .A(n1155), .B(n1156), .ZN(n1154) );
NOR2_X1 U828 ( .A1(n1157), .A2(n1153), .ZN(n1156) );
NOR2_X1 U829 ( .A1(n1148), .A2(n1158), .ZN(G60) );
XNOR2_X1 U830 ( .A(n1159), .B(n1160), .ZN(n1158) );
NOR2_X1 U831 ( .A1(n1161), .A2(n1153), .ZN(n1159) );
XNOR2_X1 U832 ( .A(G104), .B(n1162), .ZN(G6) );
NOR2_X1 U833 ( .A1(n1148), .A2(n1163), .ZN(G57) );
XOR2_X1 U834 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U835 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U836 ( .A1(n1098), .A2(n1153), .ZN(n1166) );
INV_X1 U837 ( .A(G472), .ZN(n1098) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1164) );
XNOR2_X1 U839 ( .A(n1170), .B(n1171), .ZN(n1169) );
NOR3_X1 U840 ( .A1(KEYINPUT39), .A2(n1172), .A3(n1173), .ZN(n1171) );
NOR2_X1 U841 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XNOR2_X1 U842 ( .A(n1176), .B(KEYINPUT46), .ZN(n1175) );
NOR2_X1 U843 ( .A1(n1177), .A2(n1178), .ZN(n1172) );
XNOR2_X1 U844 ( .A(KEYINPUT47), .B(n1179), .ZN(n1178) );
NOR2_X1 U845 ( .A1(n1148), .A2(n1180), .ZN(G54) );
XOR2_X1 U846 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U847 ( .A1(n1183), .A2(n1153), .ZN(n1182) );
NOR2_X1 U848 ( .A1(n1184), .A2(n1185), .ZN(n1181) );
XOR2_X1 U849 ( .A(n1186), .B(KEYINPUT8), .Z(n1185) );
NAND2_X1 U850 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NOR2_X1 U851 ( .A1(n1188), .A2(n1187), .ZN(n1184) );
XOR2_X1 U852 ( .A(n1189), .B(n1190), .Z(n1187) );
XNOR2_X1 U853 ( .A(n1191), .B(n1176), .ZN(n1188) );
NAND2_X1 U854 ( .A1(KEYINPUT45), .A2(n1192), .ZN(n1191) );
XNOR2_X1 U855 ( .A(n1193), .B(n1126), .ZN(n1192) );
NOR2_X1 U856 ( .A1(n1109), .A2(G952), .ZN(n1148) );
NOR2_X1 U857 ( .A1(n1194), .A2(n1195), .ZN(G51) );
XOR2_X1 U858 ( .A(n1196), .B(n1197), .Z(n1195) );
XNOR2_X1 U859 ( .A(n1198), .B(n1199), .ZN(n1197) );
XOR2_X1 U860 ( .A(n1200), .B(n1201), .Z(n1196) );
NOR2_X1 U861 ( .A1(KEYINPUT40), .A2(n1202), .ZN(n1201) );
NOR2_X1 U862 ( .A1(n1203), .A2(n1153), .ZN(n1200) );
NAND2_X1 U863 ( .A1(G902), .A2(n1052), .ZN(n1153) );
NAND3_X1 U864 ( .A1(n1146), .A2(n1204), .A3(n1205), .ZN(n1052) );
INV_X1 U865 ( .A(n1128), .ZN(n1205) );
NAND4_X1 U866 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1128) );
NOR3_X1 U867 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1209) );
NOR2_X1 U868 ( .A1(KEYINPUT52), .A2(n1213), .ZN(n1210) );
NAND2_X1 U869 ( .A1(n1214), .A2(n1215), .ZN(n1208) );
NAND3_X1 U870 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
NAND2_X1 U871 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NAND2_X1 U872 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NAND3_X1 U873 ( .A1(n1223), .A2(n1224), .A3(KEYINPUT52), .ZN(n1222) );
NAND3_X1 U874 ( .A1(n1225), .A2(n1226), .A3(n1056), .ZN(n1221) );
NAND2_X1 U875 ( .A1(n1057), .A2(n1227), .ZN(n1207) );
NAND2_X1 U876 ( .A1(n1228), .A2(n1217), .ZN(n1227) );
NAND2_X1 U877 ( .A1(KEYINPUT4), .A2(n1229), .ZN(n1228) );
OR3_X1 U878 ( .A1(n1216), .A2(KEYINPUT4), .A3(n1057), .ZN(n1206) );
XNOR2_X1 U879 ( .A(KEYINPUT27), .B(n1147), .ZN(n1204) );
AND4_X1 U880 ( .A1(n1162), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1146) );
AND4_X1 U881 ( .A1(n1043), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1232) );
NAND3_X1 U882 ( .A1(n1058), .A2(n1236), .A3(n1057), .ZN(n1043) );
NAND2_X1 U883 ( .A1(n1225), .A2(n1237), .ZN(n1231) );
XNOR2_X1 U884 ( .A(KEYINPUT9), .B(n1238), .ZN(n1237) );
NAND3_X1 U885 ( .A1(n1058), .A2(n1236), .A3(n1214), .ZN(n1162) );
NOR2_X1 U886 ( .A1(G952), .A2(n1239), .ZN(n1194) );
XNOR2_X1 U887 ( .A(KEYINPUT24), .B(n1109), .ZN(n1239) );
XOR2_X1 U888 ( .A(G146), .B(n1240), .Z(G48) );
NOR2_X1 U889 ( .A1(n1066), .A2(n1217), .ZN(n1240) );
INV_X1 U890 ( .A(n1214), .ZN(n1066) );
XNOR2_X1 U891 ( .A(G143), .B(n1241), .ZN(G45) );
NOR2_X1 U892 ( .A1(n1211), .A2(KEYINPUT35), .ZN(n1241) );
AND3_X1 U893 ( .A1(n1223), .A2(n1242), .A3(n1243), .ZN(n1211) );
NOR3_X1 U894 ( .A1(n1083), .A2(n1244), .A3(n1245), .ZN(n1243) );
XNOR2_X1 U895 ( .A(G140), .B(n1213), .ZN(G42) );
NAND3_X1 U896 ( .A1(n1219), .A2(n1246), .A3(n1214), .ZN(n1213) );
XOR2_X1 U897 ( .A(G137), .B(n1212), .Z(G39) );
AND2_X1 U898 ( .A1(n1247), .A2(n1246), .ZN(n1212) );
XNOR2_X1 U899 ( .A(G134), .B(n1248), .ZN(G36) );
NAND2_X1 U900 ( .A1(n1229), .A2(n1057), .ZN(n1248) );
XNOR2_X1 U901 ( .A(G131), .B(n1249), .ZN(G33) );
NAND2_X1 U902 ( .A1(n1229), .A2(n1214), .ZN(n1249) );
INV_X1 U903 ( .A(n1216), .ZN(n1229) );
NAND2_X1 U904 ( .A1(n1246), .A2(n1242), .ZN(n1216) );
AND2_X1 U905 ( .A1(n1223), .A2(n1053), .ZN(n1246) );
INV_X1 U906 ( .A(n1224), .ZN(n1053) );
NAND2_X1 U907 ( .A1(n1086), .A2(n1250), .ZN(n1224) );
XOR2_X1 U908 ( .A(G128), .B(n1251), .Z(G30) );
NOR2_X1 U909 ( .A1(n1217), .A2(n1252), .ZN(n1251) );
XOR2_X1 U910 ( .A(KEYINPUT11), .B(n1057), .Z(n1252) );
NAND4_X1 U911 ( .A1(n1253), .A2(n1223), .A3(n1225), .A4(n1254), .ZN(n1217) );
AND2_X1 U912 ( .A1(n1075), .A2(n1226), .ZN(n1223) );
XNOR2_X1 U913 ( .A(G101), .B(n1147), .ZN(G3) );
NAND3_X1 U914 ( .A1(n1242), .A2(n1236), .A3(n1069), .ZN(n1147) );
AND3_X1 U915 ( .A1(n1075), .A2(n1255), .A3(n1225), .ZN(n1236) );
XNOR2_X1 U916 ( .A(G125), .B(n1256), .ZN(G27) );
NAND4_X1 U917 ( .A1(n1257), .A2(n1056), .A3(n1258), .A4(n1214), .ZN(n1256) );
NOR2_X1 U918 ( .A1(n1083), .A2(n1080), .ZN(n1258) );
XOR2_X1 U919 ( .A(n1226), .B(KEYINPUT12), .Z(n1257) );
NAND2_X1 U920 ( .A1(n1087), .A2(n1259), .ZN(n1226) );
NAND4_X1 U921 ( .A1(G953), .A2(G902), .A3(n1260), .A4(n1111), .ZN(n1259) );
INV_X1 U922 ( .A(G900), .ZN(n1111) );
XNOR2_X1 U923 ( .A(G122), .B(n1230), .ZN(G24) );
NAND4_X1 U924 ( .A1(n1261), .A2(n1058), .A3(n1093), .A4(n1262), .ZN(n1230) );
AND2_X1 U925 ( .A1(n1095), .A2(n1263), .ZN(n1058) );
XOR2_X1 U926 ( .A(G119), .B(n1264), .Z(G21) );
NOR2_X1 U927 ( .A1(KEYINPUT15), .A2(n1235), .ZN(n1264) );
NAND2_X1 U928 ( .A1(n1261), .A2(n1247), .ZN(n1235) );
AND3_X1 U929 ( .A1(n1253), .A2(n1254), .A3(n1069), .ZN(n1247) );
XNOR2_X1 U930 ( .A(n1234), .B(n1265), .ZN(G18) );
NOR2_X1 U931 ( .A1(KEYINPUT43), .A2(n1266), .ZN(n1265) );
INV_X1 U932 ( .A(G116), .ZN(n1266) );
NAND3_X1 U933 ( .A1(n1242), .A2(n1057), .A3(n1261), .ZN(n1234) );
NOR2_X1 U934 ( .A1(n1093), .A2(n1244), .ZN(n1057) );
XNOR2_X1 U935 ( .A(G113), .B(n1233), .ZN(G15) );
NAND3_X1 U936 ( .A1(n1214), .A2(n1242), .A3(n1261), .ZN(n1233) );
AND3_X1 U937 ( .A1(n1225), .A2(n1255), .A3(n1056), .ZN(n1261) );
AND2_X1 U938 ( .A1(n1074), .A2(n1267), .ZN(n1056) );
INV_X1 U939 ( .A(n1081), .ZN(n1242) );
NAND2_X1 U940 ( .A1(n1253), .A2(n1095), .ZN(n1081) );
INV_X1 U941 ( .A(n1254), .ZN(n1095) );
XOR2_X1 U942 ( .A(n1263), .B(KEYINPUT49), .Z(n1253) );
NOR2_X1 U943 ( .A1(n1262), .A2(n1245), .ZN(n1214) );
INV_X1 U944 ( .A(n1093), .ZN(n1245) );
XNOR2_X1 U945 ( .A(n1268), .B(n1269), .ZN(G12) );
NOR2_X1 U946 ( .A1(n1083), .A2(n1238), .ZN(n1269) );
NAND4_X1 U947 ( .A1(n1219), .A2(n1069), .A3(n1075), .A4(n1255), .ZN(n1238) );
NAND2_X1 U948 ( .A1(n1087), .A2(n1270), .ZN(n1255) );
NAND3_X1 U949 ( .A1(G902), .A2(n1260), .A3(n1138), .ZN(n1270) );
NOR2_X1 U950 ( .A1(n1109), .A2(G898), .ZN(n1138) );
NAND3_X1 U951 ( .A1(n1260), .A2(n1109), .A3(G952), .ZN(n1087) );
NAND2_X1 U952 ( .A1(G237), .A2(G234), .ZN(n1260) );
NOR2_X1 U953 ( .A1(n1074), .A2(n1073), .ZN(n1075) );
INV_X1 U954 ( .A(n1267), .ZN(n1073) );
NAND2_X1 U955 ( .A1(G221), .A2(n1271), .ZN(n1267) );
XNOR2_X1 U956 ( .A(n1088), .B(KEYINPUT31), .ZN(n1074) );
XNOR2_X1 U957 ( .A(n1272), .B(n1183), .ZN(n1088) );
INV_X1 U958 ( .A(G469), .ZN(n1183) );
NAND2_X1 U959 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XOR2_X1 U960 ( .A(n1275), .B(n1276), .Z(n1273) );
XNOR2_X1 U961 ( .A(n1189), .B(n1179), .ZN(n1276) );
INV_X1 U962 ( .A(n1176), .ZN(n1179) );
NOR2_X1 U963 ( .A1(n1110), .A2(G953), .ZN(n1189) );
INV_X1 U964 ( .A(G227), .ZN(n1110) );
XOR2_X1 U965 ( .A(n1277), .B(n1278), .Z(n1275) );
XOR2_X1 U966 ( .A(n1279), .B(KEYINPUT10), .Z(n1278) );
NAND3_X1 U967 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1279) );
NAND2_X1 U968 ( .A1(G140), .A2(n1283), .ZN(n1282) );
OR3_X1 U969 ( .A1(n1283), .A2(G140), .A3(n1284), .ZN(n1281) );
NAND2_X1 U970 ( .A1(KEYINPUT50), .A2(n1268), .ZN(n1283) );
NAND2_X1 U971 ( .A1(G110), .A2(n1284), .ZN(n1280) );
INV_X1 U972 ( .A(KEYINPUT58), .ZN(n1284) );
NAND2_X1 U973 ( .A1(n1285), .A2(KEYINPUT5), .ZN(n1277) );
XOR2_X1 U974 ( .A(n1286), .B(n1193), .Z(n1285) );
XNOR2_X1 U975 ( .A(n1287), .B(n1288), .ZN(n1193) );
NAND2_X1 U976 ( .A1(KEYINPUT25), .A2(n1126), .ZN(n1286) );
XOR2_X1 U977 ( .A(n1289), .B(n1290), .Z(n1126) );
XNOR2_X1 U978 ( .A(n1291), .B(KEYINPUT37), .ZN(n1290) );
NAND2_X1 U979 ( .A1(KEYINPUT61), .A2(n1292), .ZN(n1291) );
NOR2_X1 U980 ( .A1(n1262), .A2(n1093), .ZN(n1069) );
XOR2_X1 U981 ( .A(n1293), .B(n1161), .Z(n1093) );
INV_X1 U982 ( .A(G475), .ZN(n1161) );
NAND2_X1 U983 ( .A1(n1160), .A2(n1294), .ZN(n1293) );
XNOR2_X1 U984 ( .A(KEYINPUT59), .B(n1274), .ZN(n1294) );
XOR2_X1 U985 ( .A(n1295), .B(n1296), .Z(n1160) );
XNOR2_X1 U986 ( .A(n1297), .B(n1298), .ZN(n1296) );
XNOR2_X1 U987 ( .A(KEYINPUT62), .B(n1299), .ZN(n1298) );
INV_X1 U988 ( .A(G113), .ZN(n1297) );
XNOR2_X1 U989 ( .A(G104), .B(n1300), .ZN(n1295) );
NOR2_X1 U990 ( .A1(KEYINPUT54), .A2(n1301), .ZN(n1300) );
NOR2_X1 U991 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
XOR2_X1 U992 ( .A(KEYINPUT1), .B(n1304), .Z(n1303) );
AND2_X1 U993 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NOR2_X1 U994 ( .A1(n1306), .A2(n1305), .ZN(n1302) );
NAND2_X1 U995 ( .A1(n1307), .A2(n1308), .ZN(n1305) );
NAND2_X1 U996 ( .A1(G146), .A2(n1309), .ZN(n1308) );
XOR2_X1 U997 ( .A(KEYINPUT18), .B(n1310), .Z(n1307) );
NOR2_X1 U998 ( .A1(G146), .A2(n1309), .ZN(n1310) );
INV_X1 U999 ( .A(n1115), .ZN(n1309) );
XOR2_X1 U1000 ( .A(G140), .B(n1202), .Z(n1115) );
XNOR2_X1 U1001 ( .A(n1311), .B(n1312), .ZN(n1306) );
XNOR2_X1 U1002 ( .A(n1292), .B(G131), .ZN(n1312) );
NAND2_X1 U1003 ( .A1(KEYINPUT56), .A2(n1313), .ZN(n1311) );
NAND3_X1 U1004 ( .A1(n1314), .A2(n1109), .A3(G214), .ZN(n1313) );
INV_X1 U1005 ( .A(n1244), .ZN(n1262) );
NOR2_X1 U1006 ( .A1(n1315), .A2(n1103), .ZN(n1244) );
AND3_X1 U1007 ( .A1(n1157), .A2(n1274), .A3(n1155), .ZN(n1103) );
INV_X1 U1008 ( .A(G478), .ZN(n1157) );
AND2_X1 U1009 ( .A1(G478), .A2(n1102), .ZN(n1315) );
NAND2_X1 U1010 ( .A1(n1274), .A2(n1155), .ZN(n1102) );
NAND2_X1 U1011 ( .A1(n1316), .A2(n1317), .ZN(n1155) );
NAND4_X1 U1012 ( .A1(n1318), .A2(n1109), .A3(n1319), .A4(n1320), .ZN(n1317) );
AND2_X1 U1013 ( .A1(G217), .A2(G234), .ZN(n1320) );
NAND2_X1 U1014 ( .A1(n1321), .A2(n1322), .ZN(n1316) );
NAND3_X1 U1015 ( .A1(G217), .A2(n1109), .A3(G234), .ZN(n1322) );
NAND2_X1 U1016 ( .A1(n1319), .A2(n1318), .ZN(n1321) );
NAND2_X1 U1017 ( .A1(n1323), .A2(n1324), .ZN(n1318) );
XOR2_X1 U1018 ( .A(KEYINPUT51), .B(n1325), .Z(n1323) );
XNOR2_X1 U1019 ( .A(n1326), .B(KEYINPUT0), .ZN(n1319) );
NAND2_X1 U1020 ( .A1(n1327), .A2(n1325), .ZN(n1326) );
XOR2_X1 U1021 ( .A(G107), .B(n1328), .Z(n1325) );
XNOR2_X1 U1022 ( .A(n1299), .B(G116), .ZN(n1328) );
INV_X1 U1023 ( .A(G122), .ZN(n1299) );
INV_X1 U1024 ( .A(n1324), .ZN(n1327) );
XNOR2_X1 U1025 ( .A(n1329), .B(n1330), .ZN(n1324) );
XNOR2_X1 U1026 ( .A(G134), .B(G143), .ZN(n1329) );
INV_X1 U1027 ( .A(n1080), .ZN(n1219) );
NAND2_X1 U1028 ( .A1(n1263), .A2(n1254), .ZN(n1080) );
XOR2_X1 U1029 ( .A(n1331), .B(n1152), .Z(n1254) );
NAND2_X1 U1030 ( .A1(G217), .A2(n1271), .ZN(n1152) );
NAND2_X1 U1031 ( .A1(G234), .A2(n1274), .ZN(n1271) );
NAND2_X1 U1032 ( .A1(n1150), .A2(n1274), .ZN(n1331) );
XNOR2_X1 U1033 ( .A(n1332), .B(n1333), .ZN(n1150) );
XOR2_X1 U1034 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1035 ( .A(G137), .B(G119), .Z(n1335) );
XOR2_X1 U1036 ( .A(KEYINPUT48), .B(KEYINPUT26), .Z(n1334) );
XOR2_X1 U1037 ( .A(n1336), .B(n1337), .Z(n1332) );
XOR2_X1 U1038 ( .A(n1202), .B(n1190), .Z(n1337) );
XNOR2_X1 U1039 ( .A(G140), .B(n1268), .ZN(n1190) );
XOR2_X1 U1040 ( .A(n1289), .B(n1338), .Z(n1336) );
AND3_X1 U1041 ( .A1(G221), .A2(n1109), .A3(G234), .ZN(n1338) );
XNOR2_X1 U1042 ( .A(G146), .B(n1330), .ZN(n1289) );
XNOR2_X1 U1043 ( .A(G472), .B(n1339), .ZN(n1263) );
NOR2_X1 U1044 ( .A1(KEYINPUT36), .A2(n1096), .ZN(n1339) );
NAND2_X1 U1045 ( .A1(n1340), .A2(n1274), .ZN(n1096) );
XOR2_X1 U1046 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1047 ( .A(n1167), .B(n1343), .Z(n1342) );
XNOR2_X1 U1048 ( .A(n1344), .B(n1176), .ZN(n1343) );
XOR2_X1 U1049 ( .A(G134), .B(n1127), .Z(n1176) );
XOR2_X1 U1050 ( .A(G131), .B(G137), .Z(n1127) );
NAND2_X1 U1051 ( .A1(KEYINPUT42), .A2(n1170), .ZN(n1344) );
XOR2_X1 U1052 ( .A(n1345), .B(n1346), .Z(n1341) );
XOR2_X1 U1053 ( .A(KEYINPUT53), .B(KEYINPUT23), .Z(n1346) );
XNOR2_X1 U1054 ( .A(n1347), .B(n1168), .ZN(n1345) );
NAND3_X1 U1055 ( .A1(n1314), .A2(n1109), .A3(G210), .ZN(n1168) );
NAND2_X1 U1056 ( .A1(KEYINPUT7), .A2(n1174), .ZN(n1347) );
INV_X1 U1057 ( .A(n1177), .ZN(n1174) );
XNOR2_X1 U1058 ( .A(n1199), .B(KEYINPUT28), .ZN(n1177) );
INV_X1 U1059 ( .A(n1225), .ZN(n1083) );
NOR2_X1 U1060 ( .A1(n1086), .A2(n1085), .ZN(n1225) );
INV_X1 U1061 ( .A(n1250), .ZN(n1085) );
NAND2_X1 U1062 ( .A1(G214), .A2(n1348), .ZN(n1250) );
XNOR2_X1 U1063 ( .A(n1349), .B(n1203), .ZN(n1086) );
NAND2_X1 U1064 ( .A1(G210), .A2(n1348), .ZN(n1203) );
NAND2_X1 U1065 ( .A1(n1314), .A2(n1274), .ZN(n1348) );
INV_X1 U1066 ( .A(G237), .ZN(n1314) );
NAND2_X1 U1067 ( .A1(n1350), .A2(n1274), .ZN(n1349) );
INV_X1 U1068 ( .A(G902), .ZN(n1274) );
XNOR2_X1 U1069 ( .A(n1351), .B(n1352), .ZN(n1350) );
INV_X1 U1070 ( .A(n1198), .ZN(n1352) );
XOR2_X1 U1071 ( .A(n1353), .B(n1354), .Z(n1198) );
INV_X1 U1072 ( .A(n1142), .ZN(n1354) );
XNOR2_X1 U1073 ( .A(n1355), .B(n1167), .ZN(n1142) );
XNOR2_X1 U1074 ( .A(n1356), .B(n1357), .ZN(n1167) );
XOR2_X1 U1075 ( .A(KEYINPUT32), .B(G119), .Z(n1357) );
XNOR2_X1 U1076 ( .A(G113), .B(G116), .ZN(n1356) );
NAND3_X1 U1077 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1355) );
NAND2_X1 U1078 ( .A1(G122), .A2(n1268), .ZN(n1360) );
NAND2_X1 U1079 ( .A1(KEYINPUT29), .A2(n1361), .ZN(n1359) );
NAND2_X1 U1080 ( .A1(n1362), .A2(G110), .ZN(n1361) );
XNOR2_X1 U1081 ( .A(KEYINPUT2), .B(G122), .ZN(n1362) );
NAND2_X1 U1082 ( .A1(n1363), .A2(n1364), .ZN(n1358) );
INV_X1 U1083 ( .A(KEYINPUT29), .ZN(n1364) );
NAND2_X1 U1084 ( .A1(n1365), .A2(n1366), .ZN(n1363) );
OR3_X1 U1085 ( .A1(n1268), .A2(G122), .A3(KEYINPUT2), .ZN(n1366) );
NAND2_X1 U1086 ( .A1(KEYINPUT2), .A2(G122), .ZN(n1365) );
XOR2_X1 U1087 ( .A(n1367), .B(n1368), .Z(n1353) );
NOR2_X1 U1088 ( .A1(KEYINPUT16), .A2(n1143), .ZN(n1368) );
XNOR2_X1 U1089 ( .A(n1369), .B(n1288), .ZN(n1143) );
XNOR2_X1 U1090 ( .A(G107), .B(n1170), .ZN(n1288) );
INV_X1 U1091 ( .A(G101), .ZN(n1170) );
NAND2_X1 U1092 ( .A1(KEYINPUT41), .A2(n1287), .ZN(n1369) );
INV_X1 U1093 ( .A(G104), .ZN(n1287) );
NAND2_X1 U1094 ( .A1(G224), .A2(n1109), .ZN(n1367) );
INV_X1 U1095 ( .A(G953), .ZN(n1109) );
XNOR2_X1 U1096 ( .A(KEYINPUT19), .B(n1370), .ZN(n1351) );
NOR2_X1 U1097 ( .A1(KEYINPUT14), .A2(n1371), .ZN(n1370) );
XOR2_X1 U1098 ( .A(n1199), .B(n1202), .Z(n1371) );
XOR2_X1 U1099 ( .A(G125), .B(KEYINPUT22), .Z(n1202) );
XOR2_X1 U1100 ( .A(n1372), .B(n1330), .Z(n1199) );
XOR2_X1 U1101 ( .A(G128), .B(KEYINPUT30), .Z(n1330) );
NAND2_X1 U1102 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
NAND2_X1 U1103 ( .A1(G146), .A2(n1292), .ZN(n1374) );
XOR2_X1 U1104 ( .A(KEYINPUT44), .B(n1375), .Z(n1373) );
NOR2_X1 U1105 ( .A1(G146), .A2(n1292), .ZN(n1375) );
INV_X1 U1106 ( .A(G143), .ZN(n1292) );
INV_X1 U1107 ( .A(G110), .ZN(n1268) );
endmodule


