//Key = 1100010111000000011000101110110001001101001101110001001111101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
n1415, n1416, n1417, n1418, n1419, n1420, n1421;

XNOR2_X1 U770 ( .A(n1075), .B(n1076), .ZN(G9) );
NOR2_X1 U771 ( .A1(KEYINPUT63), .A2(n1077), .ZN(n1076) );
NOR2_X1 U772 ( .A1(n1078), .A2(n1079), .ZN(G75) );
XOR2_X1 U773 ( .A(n1080), .B(KEYINPUT58), .Z(n1079) );
NAND4_X1 U774 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1080) );
NOR2_X1 U775 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U776 ( .A(KEYINPUT33), .B(n1087), .Z(n1086) );
NOR2_X1 U777 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR2_X1 U778 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
XOR2_X1 U780 ( .A(n1094), .B(KEYINPUT25), .Z(n1093) );
NAND2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR3_X1 U782 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1092) );
NOR2_X1 U783 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
AND2_X1 U784 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR2_X1 U785 ( .A1(n1104), .A2(n1105), .ZN(n1100) );
XNOR2_X1 U786 ( .A(KEYINPUT0), .B(n1106), .ZN(n1105) );
AND3_X1 U787 ( .A1(n1095), .A2(n1107), .A3(n1108), .ZN(n1088) );
INV_X1 U788 ( .A(n1109), .ZN(n1083) );
NAND3_X1 U789 ( .A1(n1108), .A2(n1110), .A3(n1111), .ZN(n1082) );
INV_X1 U790 ( .A(n1097), .ZN(n1111) );
NAND2_X1 U791 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NAND4_X1 U792 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1113) );
NAND2_X1 U793 ( .A1(n1102), .A2(n1118), .ZN(n1112) );
NAND2_X1 U794 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND3_X1 U795 ( .A1(n1121), .A2(n1117), .A3(n1122), .ZN(n1120) );
NAND2_X1 U796 ( .A1(n1115), .A2(n1123), .ZN(n1119) );
NAND3_X1 U797 ( .A1(n1115), .A2(n1124), .A3(n1095), .ZN(n1081) );
NOR3_X1 U798 ( .A1(n1125), .A2(n1104), .A3(n1097), .ZN(n1095) );
NOR2_X1 U799 ( .A1(G952), .A2(n1109), .ZN(n1078) );
NAND2_X1 U800 ( .A1(n1126), .A2(n1127), .ZN(n1109) );
NAND4_X1 U801 ( .A1(n1128), .A2(n1108), .A3(n1102), .A4(n1129), .ZN(n1127) );
NOR4_X1 U802 ( .A1(n1122), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1129) );
XOR2_X1 U803 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U804 ( .A1(KEYINPUT18), .A2(n1135), .ZN(n1133) );
XOR2_X1 U805 ( .A(n1136), .B(n1137), .Z(G72) );
XOR2_X1 U806 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR3_X1 U807 ( .A1(n1140), .A2(KEYINPUT2), .A3(G953), .ZN(n1139) );
NOR3_X1 U808 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1140) );
INV_X1 U809 ( .A(n1144), .ZN(n1142) );
XNOR2_X1 U810 ( .A(KEYINPUT15), .B(n1145), .ZN(n1141) );
NAND3_X1 U811 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1138) );
XOR2_X1 U812 ( .A(KEYINPUT5), .B(n1149), .Z(n1148) );
NOR2_X1 U813 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XNOR2_X1 U814 ( .A(n1152), .B(n1153), .ZN(n1151) );
AND2_X1 U815 ( .A1(n1154), .A2(KEYINPUT57), .ZN(n1153) );
NAND3_X1 U816 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1147) );
XNOR2_X1 U817 ( .A(KEYINPUT17), .B(n1150), .ZN(n1157) );
XOR2_X1 U818 ( .A(n1158), .B(n1159), .Z(n1150) );
NOR2_X1 U819 ( .A1(G125), .A2(KEYINPUT3), .ZN(n1159) );
NAND2_X1 U820 ( .A1(n1160), .A2(n1154), .ZN(n1156) );
XOR2_X1 U821 ( .A(KEYINPUT57), .B(n1152), .Z(n1160) );
NAND2_X1 U822 ( .A1(n1152), .A2(n1161), .ZN(n1155) );
XNOR2_X1 U823 ( .A(n1162), .B(n1163), .ZN(n1152) );
NOR2_X1 U824 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XOR2_X1 U825 ( .A(KEYINPUT44), .B(n1166), .Z(n1165) );
NOR2_X1 U826 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XNOR2_X1 U827 ( .A(KEYINPUT35), .B(n1169), .ZN(n1168) );
NAND2_X1 U828 ( .A1(KEYINPUT60), .A2(n1170), .ZN(n1162) );
NAND2_X1 U829 ( .A1(G953), .A2(n1171), .ZN(n1146) );
NAND2_X1 U830 ( .A1(n1172), .A2(n1173), .ZN(n1136) );
NAND2_X1 U831 ( .A1(G900), .A2(G227), .ZN(n1173) );
INV_X1 U832 ( .A(n1174), .ZN(n1172) );
XOR2_X1 U833 ( .A(n1175), .B(n1176), .Z(G69) );
NOR2_X1 U834 ( .A1(n1174), .A2(n1177), .ZN(n1176) );
XOR2_X1 U835 ( .A(KEYINPUT52), .B(n1178), .Z(n1177) );
NOR2_X1 U836 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XOR2_X1 U837 ( .A(G953), .B(KEYINPUT54), .Z(n1174) );
NAND2_X1 U838 ( .A1(n1181), .A2(n1182), .ZN(n1175) );
NAND2_X1 U839 ( .A1(n1183), .A2(n1126), .ZN(n1182) );
XNOR2_X1 U840 ( .A(n1184), .B(n1185), .ZN(n1183) );
NAND3_X1 U841 ( .A1(G898), .A2(n1184), .A3(G953), .ZN(n1181) );
XNOR2_X1 U842 ( .A(n1186), .B(n1187), .ZN(n1184) );
NOR2_X1 U843 ( .A1(n1188), .A2(n1189), .ZN(G66) );
NOR3_X1 U844 ( .A1(n1134), .A2(n1190), .A3(n1191), .ZN(n1189) );
NOR3_X1 U845 ( .A1(n1192), .A2(n1135), .A3(n1193), .ZN(n1191) );
INV_X1 U846 ( .A(n1194), .ZN(n1192) );
NOR2_X1 U847 ( .A1(n1195), .A2(n1194), .ZN(n1190) );
NOR2_X1 U848 ( .A1(n1196), .A2(n1135), .ZN(n1195) );
INV_X1 U849 ( .A(n1085), .ZN(n1196) );
NOR2_X1 U850 ( .A1(n1188), .A2(n1197), .ZN(G63) );
XOR2_X1 U851 ( .A(n1198), .B(n1199), .Z(n1197) );
NOR2_X1 U852 ( .A1(n1200), .A2(n1193), .ZN(n1199) );
INV_X1 U853 ( .A(G478), .ZN(n1200) );
NAND2_X1 U854 ( .A1(KEYINPUT42), .A2(n1201), .ZN(n1198) );
INV_X1 U855 ( .A(n1202), .ZN(n1201) );
NOR2_X1 U856 ( .A1(n1188), .A2(n1203), .ZN(G60) );
XNOR2_X1 U857 ( .A(n1204), .B(n1205), .ZN(n1203) );
NOR2_X1 U858 ( .A1(n1206), .A2(n1193), .ZN(n1205) );
XNOR2_X1 U859 ( .A(G104), .B(n1207), .ZN(G6) );
NOR3_X1 U860 ( .A1(n1188), .A2(n1208), .A3(n1209), .ZN(G57) );
NOR3_X1 U861 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1209) );
NOR2_X1 U862 ( .A1(KEYINPUT62), .A2(KEYINPUT9), .ZN(n1211) );
NOR2_X1 U863 ( .A1(n1213), .A2(n1214), .ZN(n1208) );
NOR2_X1 U864 ( .A1(n1215), .A2(n1216), .ZN(n1213) );
XOR2_X1 U865 ( .A(KEYINPUT62), .B(n1212), .Z(n1216) );
XNOR2_X1 U866 ( .A(n1217), .B(n1218), .ZN(n1212) );
XOR2_X1 U867 ( .A(n1219), .B(n1220), .Z(n1218) );
NOR2_X1 U868 ( .A1(n1221), .A2(n1193), .ZN(n1220) );
NOR2_X1 U869 ( .A1(KEYINPUT10), .A2(n1222), .ZN(n1219) );
XNOR2_X1 U870 ( .A(n1223), .B(KEYINPUT23), .ZN(n1222) );
INV_X1 U871 ( .A(KEYINPUT9), .ZN(n1215) );
NOR3_X1 U872 ( .A1(n1188), .A2(n1224), .A3(n1225), .ZN(G54) );
NOR2_X1 U873 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
XOR2_X1 U874 ( .A(n1228), .B(n1229), .Z(n1226) );
NOR2_X1 U875 ( .A1(n1230), .A2(KEYINPUT53), .ZN(n1228) );
INV_X1 U876 ( .A(n1231), .ZN(n1230) );
NOR2_X1 U877 ( .A1(n1232), .A2(n1233), .ZN(n1224) );
XOR2_X1 U878 ( .A(n1234), .B(n1229), .Z(n1233) );
XNOR2_X1 U879 ( .A(n1235), .B(n1236), .ZN(n1229) );
XOR2_X1 U880 ( .A(n1237), .B(n1238), .Z(n1236) );
NOR2_X1 U881 ( .A1(G140), .A2(KEYINPUT31), .ZN(n1238) );
NOR2_X1 U882 ( .A1(n1239), .A2(n1193), .ZN(n1237) );
XNOR2_X1 U883 ( .A(G110), .B(n1240), .ZN(n1235) );
NOR2_X1 U884 ( .A1(KEYINPUT53), .A2(n1231), .ZN(n1234) );
NAND3_X1 U885 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1231) );
NAND2_X1 U886 ( .A1(KEYINPUT30), .A2(n1244), .ZN(n1243) );
NAND3_X1 U887 ( .A1(n1245), .A2(n1246), .A3(n1154), .ZN(n1242) );
INV_X1 U888 ( .A(KEYINPUT30), .ZN(n1246) );
OR2_X1 U889 ( .A1(n1154), .A2(n1245), .ZN(n1241) );
NOR2_X1 U890 ( .A1(KEYINPUT32), .A2(n1244), .ZN(n1245) );
NOR2_X1 U891 ( .A1(n1188), .A2(n1247), .ZN(G51) );
XNOR2_X1 U892 ( .A(n1248), .B(n1249), .ZN(n1247) );
NOR2_X1 U893 ( .A1(n1250), .A2(n1193), .ZN(n1249) );
NAND2_X1 U894 ( .A1(G902), .A2(n1085), .ZN(n1193) );
NAND4_X1 U895 ( .A1(n1185), .A2(n1251), .A3(n1252), .A4(n1145), .ZN(n1085) );
XNOR2_X1 U896 ( .A(KEYINPUT51), .B(n1144), .ZN(n1252) );
INV_X1 U897 ( .A(n1143), .ZN(n1251) );
NAND4_X1 U898 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1143) );
NOR3_X1 U899 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1256) );
NOR2_X1 U900 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND4_X1 U901 ( .A1(n1262), .A2(n1263), .A3(n1264), .A4(n1091), .ZN(n1261) );
INV_X1 U902 ( .A(n1115), .ZN(n1091) );
INV_X1 U903 ( .A(KEYINPUT6), .ZN(n1260) );
NOR2_X1 U904 ( .A1(KEYINPUT6), .A2(n1265), .ZN(n1258) );
NOR2_X1 U905 ( .A1(n1266), .A2(n1267), .ZN(n1257) );
NOR2_X1 U906 ( .A1(n1096), .A2(n1268), .ZN(n1266) );
XOR2_X1 U907 ( .A(KEYINPUT34), .B(n1124), .Z(n1268) );
AND4_X1 U908 ( .A1(n1269), .A2(n1270), .A3(n1271), .A4(n1272), .ZN(n1185) );
AND4_X1 U909 ( .A1(n1273), .A2(n1274), .A3(n1075), .A4(n1207), .ZN(n1272) );
NAND3_X1 U910 ( .A1(n1275), .A2(n1117), .A3(n1096), .ZN(n1207) );
NAND3_X1 U911 ( .A1(n1275), .A2(n1117), .A3(n1124), .ZN(n1075) );
NOR2_X1 U912 ( .A1(n1276), .A2(n1277), .ZN(n1271) );
NOR2_X1 U913 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
XOR2_X1 U914 ( .A(n1280), .B(KEYINPUT41), .Z(n1278) );
AND3_X1 U915 ( .A1(n1123), .A2(n1275), .A3(n1108), .ZN(n1276) );
NOR2_X1 U916 ( .A1(n1126), .A2(G952), .ZN(n1188) );
XOR2_X1 U917 ( .A(n1281), .B(G146), .Z(G48) );
NAND2_X1 U918 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND4_X1 U919 ( .A1(n1096), .A2(n1284), .A3(n1285), .A4(n1286), .ZN(n1283) );
OR2_X1 U920 ( .A1(n1145), .A2(n1286), .ZN(n1282) );
INV_X1 U921 ( .A(KEYINPUT28), .ZN(n1286) );
NAND3_X1 U922 ( .A1(n1287), .A2(n1096), .A3(n1285), .ZN(n1145) );
XNOR2_X1 U923 ( .A(G143), .B(n1255), .ZN(G45) );
NAND4_X1 U924 ( .A1(n1285), .A2(n1103), .A3(n1288), .A4(n1289), .ZN(n1255) );
XNOR2_X1 U925 ( .A(n1158), .B(n1290), .ZN(G42) );
NOR2_X1 U926 ( .A1(KEYINPUT48), .A2(n1144), .ZN(n1290) );
NAND3_X1 U927 ( .A1(n1123), .A2(n1096), .A3(n1291), .ZN(n1144) );
XOR2_X1 U928 ( .A(n1265), .B(n1292), .Z(G39) );
XNOR2_X1 U929 ( .A(KEYINPUT22), .B(n1169), .ZN(n1292) );
NAND2_X1 U930 ( .A1(n1291), .A2(n1262), .ZN(n1265) );
XOR2_X1 U931 ( .A(n1293), .B(n1294), .Z(G36) );
XNOR2_X1 U932 ( .A(G134), .B(KEYINPUT13), .ZN(n1294) );
NAND2_X1 U933 ( .A1(n1295), .A2(n1124), .ZN(n1293) );
INV_X1 U934 ( .A(n1267), .ZN(n1295) );
XOR2_X1 U935 ( .A(G131), .B(n1296), .Z(G33) );
NOR2_X1 U936 ( .A1(n1297), .A2(n1267), .ZN(n1296) );
NAND2_X1 U937 ( .A1(n1291), .A2(n1103), .ZN(n1267) );
AND3_X1 U938 ( .A1(n1263), .A2(n1264), .A3(n1115), .ZN(n1291) );
NOR2_X1 U939 ( .A1(n1298), .A2(n1122), .ZN(n1115) );
XNOR2_X1 U940 ( .A(G128), .B(n1254), .ZN(G30) );
NAND3_X1 U941 ( .A1(n1287), .A2(n1124), .A3(n1285), .ZN(n1254) );
AND3_X1 U942 ( .A1(n1107), .A2(n1264), .A3(n1263), .ZN(n1285) );
XOR2_X1 U943 ( .A(n1269), .B(n1299), .Z(G3) );
XNOR2_X1 U944 ( .A(G101), .B(KEYINPUT40), .ZN(n1299) );
NAND3_X1 U945 ( .A1(n1108), .A2(n1275), .A3(n1103), .ZN(n1269) );
NOR3_X1 U946 ( .A1(n1300), .A2(n1301), .A3(n1106), .ZN(n1275) );
INV_X1 U947 ( .A(n1302), .ZN(n1300) );
XNOR2_X1 U948 ( .A(G125), .B(n1253), .ZN(G27) );
NAND3_X1 U949 ( .A1(n1123), .A2(n1096), .A3(n1303), .ZN(n1253) );
AND3_X1 U950 ( .A1(n1102), .A2(n1264), .A3(n1107), .ZN(n1303) );
NAND2_X1 U951 ( .A1(n1304), .A2(n1097), .ZN(n1264) );
XOR2_X1 U952 ( .A(n1305), .B(KEYINPUT19), .Z(n1304) );
NAND4_X1 U953 ( .A1(G953), .A2(G902), .A3(n1306), .A4(n1171), .ZN(n1305) );
INV_X1 U954 ( .A(G900), .ZN(n1171) );
INV_X1 U955 ( .A(n1125), .ZN(n1102) );
XNOR2_X1 U956 ( .A(G122), .B(n1270), .ZN(G24) );
NAND3_X1 U957 ( .A1(n1307), .A2(n1117), .A3(n1308), .ZN(n1270) );
AND3_X1 U958 ( .A1(n1107), .A2(n1289), .A3(n1288), .ZN(n1308) );
INV_X1 U959 ( .A(n1104), .ZN(n1117) );
NAND2_X1 U960 ( .A1(n1309), .A2(n1128), .ZN(n1104) );
XNOR2_X1 U961 ( .A(G119), .B(n1274), .ZN(G21) );
NAND3_X1 U962 ( .A1(n1307), .A2(n1107), .A3(n1262), .ZN(n1274) );
NOR2_X1 U963 ( .A1(n1284), .A2(n1099), .ZN(n1262) );
INV_X1 U964 ( .A(n1287), .ZN(n1284) );
NOR2_X1 U965 ( .A1(n1128), .A2(n1309), .ZN(n1287) );
INV_X1 U966 ( .A(n1310), .ZN(n1309) );
XOR2_X1 U967 ( .A(G116), .B(n1311), .Z(G18) );
NOR2_X1 U968 ( .A1(n1279), .A2(n1280), .ZN(n1311) );
NAND3_X1 U969 ( .A1(n1307), .A2(n1124), .A3(n1103), .ZN(n1280) );
NOR2_X1 U970 ( .A1(n1288), .A2(n1312), .ZN(n1124) );
INV_X1 U971 ( .A(n1107), .ZN(n1279) );
XNOR2_X1 U972 ( .A(G113), .B(n1273), .ZN(G15) );
NAND4_X1 U973 ( .A1(n1096), .A2(n1103), .A3(n1307), .A4(n1302), .ZN(n1273) );
NOR2_X1 U974 ( .A1(n1125), .A2(n1301), .ZN(n1307) );
NAND2_X1 U975 ( .A1(n1116), .A2(n1313), .ZN(n1125) );
NOR2_X1 U976 ( .A1(n1310), .A2(n1128), .ZN(n1103) );
INV_X1 U977 ( .A(n1297), .ZN(n1096) );
NAND2_X1 U978 ( .A1(n1312), .A2(n1288), .ZN(n1297) );
INV_X1 U979 ( .A(n1289), .ZN(n1312) );
XNOR2_X1 U980 ( .A(G110), .B(n1314), .ZN(G12) );
NAND3_X1 U981 ( .A1(n1315), .A2(n1123), .A3(n1316), .ZN(n1314) );
NOR3_X1 U982 ( .A1(n1099), .A2(n1301), .A3(n1106), .ZN(n1316) );
INV_X1 U983 ( .A(n1263), .ZN(n1106) );
NOR2_X1 U984 ( .A1(n1116), .A2(n1114), .ZN(n1263) );
INV_X1 U985 ( .A(n1313), .ZN(n1114) );
NAND2_X1 U986 ( .A1(G221), .A2(n1317), .ZN(n1313) );
XNOR2_X1 U987 ( .A(n1318), .B(n1239), .ZN(n1116) );
INV_X1 U988 ( .A(G469), .ZN(n1239) );
NAND2_X1 U989 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
XOR2_X1 U990 ( .A(n1321), .B(n1322), .Z(n1319) );
XOR2_X1 U991 ( .A(n1240), .B(n1323), .Z(n1322) );
NOR2_X1 U992 ( .A1(KEYINPUT4), .A2(n1324), .ZN(n1323) );
XNOR2_X1 U993 ( .A(n1325), .B(n1154), .ZN(n1324) );
INV_X1 U994 ( .A(n1161), .ZN(n1154) );
XOR2_X1 U995 ( .A(n1326), .B(n1327), .Z(n1161) );
XNOR2_X1 U996 ( .A(n1232), .B(n1244), .ZN(n1325) );
XNOR2_X1 U997 ( .A(G101), .B(n1328), .ZN(n1244) );
INV_X1 U998 ( .A(n1227), .ZN(n1232) );
AND2_X1 U999 ( .A1(G227), .A2(n1126), .ZN(n1240) );
XNOR2_X1 U1000 ( .A(G110), .B(G140), .ZN(n1321) );
AND2_X1 U1001 ( .A1(n1097), .A2(n1329), .ZN(n1301) );
NAND4_X1 U1002 ( .A1(G953), .A2(G902), .A3(n1306), .A4(n1180), .ZN(n1329) );
INV_X1 U1003 ( .A(G898), .ZN(n1180) );
NAND3_X1 U1004 ( .A1(n1306), .A2(n1126), .A3(G952), .ZN(n1097) );
NAND2_X1 U1005 ( .A1(G237), .A2(G234), .ZN(n1306) );
INV_X1 U1006 ( .A(n1108), .ZN(n1099) );
NOR2_X1 U1007 ( .A1(n1289), .A2(n1288), .ZN(n1108) );
XOR2_X1 U1008 ( .A(n1330), .B(n1206), .Z(n1288) );
INV_X1 U1009 ( .A(G475), .ZN(n1206) );
NAND2_X1 U1010 ( .A1(n1320), .A2(n1204), .ZN(n1330) );
NAND2_X1 U1011 ( .A1(n1331), .A2(n1332), .ZN(n1204) );
NAND2_X1 U1012 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
XOR2_X1 U1013 ( .A(n1335), .B(KEYINPUT11), .Z(n1331) );
OR2_X1 U1014 ( .A1(n1334), .A2(n1333), .ZN(n1335) );
XOR2_X1 U1015 ( .A(G104), .B(n1336), .Z(n1333) );
XNOR2_X1 U1016 ( .A(n1337), .B(G113), .ZN(n1336) );
INV_X1 U1017 ( .A(G122), .ZN(n1337) );
XNOR2_X1 U1018 ( .A(n1338), .B(n1339), .ZN(n1334) );
XOR2_X1 U1019 ( .A(n1340), .B(n1341), .Z(n1339) );
XNOR2_X1 U1020 ( .A(G131), .B(n1342), .ZN(n1341) );
XNOR2_X1 U1021 ( .A(KEYINPUT61), .B(n1158), .ZN(n1340) );
XOR2_X1 U1022 ( .A(n1343), .B(n1344), .Z(n1338) );
XOR2_X1 U1023 ( .A(n1345), .B(n1346), .Z(n1343) );
NOR2_X1 U1024 ( .A1(KEYINPUT20), .A2(G143), .ZN(n1346) );
NAND2_X1 U1025 ( .A1(G214), .A2(n1347), .ZN(n1345) );
XOR2_X1 U1026 ( .A(G478), .B(n1348), .Z(n1289) );
NOR2_X1 U1027 ( .A1(G902), .A2(n1202), .ZN(n1348) );
NAND3_X1 U1028 ( .A1(n1349), .A2(n1350), .A3(n1351), .ZN(n1202) );
NAND2_X1 U1029 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
INV_X1 U1030 ( .A(KEYINPUT37), .ZN(n1353) );
NAND3_X1 U1031 ( .A1(KEYINPUT37), .A2(n1354), .A3(n1355), .ZN(n1350) );
OR2_X1 U1032 ( .A1(n1355), .A2(n1354), .ZN(n1349) );
NOR2_X1 U1033 ( .A1(n1356), .A2(n1352), .ZN(n1354) );
NAND3_X1 U1034 ( .A1(G217), .A2(n1126), .A3(G234), .ZN(n1352) );
INV_X1 U1035 ( .A(KEYINPUT45), .ZN(n1356) );
XNOR2_X1 U1036 ( .A(n1357), .B(n1358), .ZN(n1355) );
XOR2_X1 U1037 ( .A(n1327), .B(n1359), .Z(n1358) );
XNOR2_X1 U1038 ( .A(G107), .B(G134), .ZN(n1357) );
AND2_X1 U1039 ( .A1(n1128), .A2(n1310), .ZN(n1123) );
XNOR2_X1 U1040 ( .A(n1134), .B(n1135), .ZN(n1310) );
NAND2_X1 U1041 ( .A1(G217), .A2(n1317), .ZN(n1135) );
NAND2_X1 U1042 ( .A1(n1360), .A2(n1320), .ZN(n1317) );
XOR2_X1 U1043 ( .A(KEYINPUT21), .B(G234), .Z(n1360) );
NOR2_X1 U1044 ( .A1(n1194), .A2(G902), .ZN(n1134) );
XNOR2_X1 U1045 ( .A(n1361), .B(n1362), .ZN(n1194) );
AND3_X1 U1046 ( .A1(G221), .A2(n1126), .A3(G234), .ZN(n1362) );
INV_X1 U1047 ( .A(G953), .ZN(n1126) );
XNOR2_X1 U1048 ( .A(n1363), .B(n1169), .ZN(n1361) );
NAND2_X1 U1049 ( .A1(n1364), .A2(KEYINPUT55), .ZN(n1363) );
XOR2_X1 U1050 ( .A(n1365), .B(n1344), .Z(n1364) );
XNOR2_X1 U1051 ( .A(n1366), .B(KEYINPUT16), .ZN(n1344) );
XNOR2_X1 U1052 ( .A(n1367), .B(n1368), .ZN(n1365) );
NAND3_X1 U1053 ( .A1(n1369), .A2(n1370), .A3(KEYINPUT56), .ZN(n1368) );
NAND3_X1 U1054 ( .A1(n1371), .A2(n1372), .A3(n1342), .ZN(n1370) );
NAND2_X1 U1055 ( .A1(n1373), .A2(n1158), .ZN(n1372) );
INV_X1 U1056 ( .A(G140), .ZN(n1158) );
NAND2_X1 U1057 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
INV_X1 U1058 ( .A(KEYINPUT14), .ZN(n1375) );
XNOR2_X1 U1059 ( .A(KEYINPUT39), .B(n1376), .ZN(n1374) );
NAND2_X1 U1060 ( .A1(G140), .A2(n1377), .ZN(n1371) );
NAND2_X1 U1061 ( .A1(KEYINPUT39), .A2(KEYINPUT12), .ZN(n1377) );
NAND2_X1 U1062 ( .A1(n1378), .A2(n1376), .ZN(n1369) );
INV_X1 U1063 ( .A(KEYINPUT12), .ZN(n1376) );
NAND2_X1 U1064 ( .A1(n1379), .A2(n1380), .ZN(n1378) );
NAND2_X1 U1065 ( .A1(G140), .A2(n1381), .ZN(n1380) );
NAND2_X1 U1066 ( .A1(KEYINPUT39), .A2(n1342), .ZN(n1381) );
NAND2_X1 U1067 ( .A1(KEYINPUT14), .A2(G125), .ZN(n1379) );
NAND4_X1 U1068 ( .A1(KEYINPUT36), .A2(n1382), .A3(n1383), .A4(n1384), .ZN(n1367) );
OR3_X1 U1069 ( .A1(n1385), .A2(KEYINPUT59), .A3(G110), .ZN(n1384) );
NAND2_X1 U1070 ( .A1(G110), .A2(n1385), .ZN(n1383) );
NAND2_X1 U1071 ( .A1(KEYINPUT8), .A2(n1386), .ZN(n1385) );
INV_X1 U1072 ( .A(n1387), .ZN(n1386) );
NAND2_X1 U1073 ( .A1(KEYINPUT59), .A2(n1387), .ZN(n1382) );
XNOR2_X1 U1074 ( .A(G128), .B(G119), .ZN(n1387) );
XNOR2_X1 U1075 ( .A(n1388), .B(n1221), .ZN(n1128) );
INV_X1 U1076 ( .A(G472), .ZN(n1221) );
NAND2_X1 U1077 ( .A1(n1389), .A2(n1320), .ZN(n1388) );
XNOR2_X1 U1078 ( .A(n1390), .B(n1391), .ZN(n1389) );
INV_X1 U1079 ( .A(n1223), .ZN(n1391) );
XNOR2_X1 U1080 ( .A(n1217), .B(n1210), .ZN(n1390) );
INV_X1 U1081 ( .A(n1214), .ZN(n1210) );
XOR2_X1 U1082 ( .A(n1392), .B(n1393), .Z(n1214) );
INV_X1 U1083 ( .A(G101), .ZN(n1393) );
NAND2_X1 U1084 ( .A1(G210), .A2(n1347), .ZN(n1392) );
NOR2_X1 U1085 ( .A1(G953), .A2(G237), .ZN(n1347) );
XOR2_X1 U1086 ( .A(n1394), .B(n1395), .Z(n1217) );
XNOR2_X1 U1087 ( .A(G113), .B(n1227), .ZN(n1395) );
NAND3_X1 U1088 ( .A1(n1396), .A2(n1397), .A3(n1398), .ZN(n1227) );
NAND2_X1 U1089 ( .A1(n1164), .A2(n1399), .ZN(n1398) );
INV_X1 U1090 ( .A(n1170), .ZN(n1399) );
NOR2_X1 U1091 ( .A1(n1169), .A2(G134), .ZN(n1164) );
NAND3_X1 U1092 ( .A1(G134), .A2(n1170), .A3(G137), .ZN(n1397) );
NAND2_X1 U1093 ( .A1(n1400), .A2(n1169), .ZN(n1396) );
INV_X1 U1094 ( .A(G137), .ZN(n1169) );
XNOR2_X1 U1095 ( .A(n1167), .B(n1170), .ZN(n1400) );
XOR2_X1 U1096 ( .A(G131), .B(KEYINPUT7), .Z(n1170) );
INV_X1 U1097 ( .A(G134), .ZN(n1167) );
NAND2_X1 U1098 ( .A1(KEYINPUT46), .A2(n1401), .ZN(n1394) );
XOR2_X1 U1099 ( .A(G119), .B(G116), .Z(n1401) );
XNOR2_X1 U1100 ( .A(n1302), .B(KEYINPUT43), .ZN(n1315) );
XOR2_X1 U1101 ( .A(n1107), .B(KEYINPUT49), .Z(n1302) );
NOR2_X1 U1102 ( .A1(n1121), .A2(n1122), .ZN(n1107) );
AND2_X1 U1103 ( .A1(G214), .A2(n1402), .ZN(n1122) );
INV_X1 U1104 ( .A(n1298), .ZN(n1121) );
NAND3_X1 U1105 ( .A1(n1403), .A2(n1404), .A3(n1405), .ZN(n1298) );
INV_X1 U1106 ( .A(n1131), .ZN(n1405) );
NOR2_X1 U1107 ( .A1(n1406), .A2(n1407), .ZN(n1131) );
NAND2_X1 U1108 ( .A1(n1130), .A2(KEYINPUT1), .ZN(n1404) );
AND2_X1 U1109 ( .A1(n1407), .A2(n1406), .ZN(n1130) );
NAND2_X1 U1110 ( .A1(n1408), .A2(n1320), .ZN(n1406) );
XNOR2_X1 U1111 ( .A(KEYINPUT27), .B(n1409), .ZN(n1408) );
INV_X1 U1112 ( .A(n1248), .ZN(n1409) );
XNOR2_X1 U1113 ( .A(n1410), .B(n1411), .ZN(n1248) );
XNOR2_X1 U1114 ( .A(n1223), .B(n1186), .ZN(n1411) );
XOR2_X1 U1115 ( .A(n1412), .B(n1413), .Z(n1186) );
XOR2_X1 U1116 ( .A(G113), .B(n1414), .Z(n1413) );
XOR2_X1 U1117 ( .A(KEYINPUT38), .B(G119), .Z(n1414) );
XNOR2_X1 U1118 ( .A(G110), .B(n1359), .ZN(n1412) );
XOR2_X1 U1119 ( .A(G116), .B(G122), .Z(n1359) );
XNOR2_X1 U1120 ( .A(n1415), .B(n1327), .ZN(n1223) );
XOR2_X1 U1121 ( .A(G128), .B(G143), .Z(n1327) );
NAND2_X1 U1122 ( .A1(KEYINPUT26), .A2(n1416), .ZN(n1415) );
XNOR2_X1 U1123 ( .A(KEYINPUT50), .B(n1366), .ZN(n1416) );
INV_X1 U1124 ( .A(n1326), .ZN(n1366) );
XOR2_X1 U1125 ( .A(G146), .B(KEYINPUT47), .Z(n1326) );
XOR2_X1 U1126 ( .A(n1417), .B(n1418), .Z(n1410) );
XNOR2_X1 U1127 ( .A(n1342), .B(n1419), .ZN(n1418) );
NOR2_X1 U1128 ( .A1(G953), .A2(n1179), .ZN(n1419) );
INV_X1 U1129 ( .A(G224), .ZN(n1179) );
INV_X1 U1130 ( .A(G125), .ZN(n1342) );
NAND2_X1 U1131 ( .A1(KEYINPUT24), .A2(n1187), .ZN(n1417) );
XNOR2_X1 U1132 ( .A(n1420), .B(G101), .ZN(n1187) );
NAND2_X1 U1133 ( .A1(KEYINPUT29), .A2(n1328), .ZN(n1420) );
XOR2_X1 U1134 ( .A(G104), .B(n1077), .Z(n1328) );
INV_X1 U1135 ( .A(G107), .ZN(n1077) );
OR2_X1 U1136 ( .A1(n1407), .A2(KEYINPUT1), .ZN(n1403) );
INV_X1 U1137 ( .A(n1250), .ZN(n1407) );
NAND2_X1 U1138 ( .A1(G210), .A2(n1402), .ZN(n1250) );
NAND2_X1 U1139 ( .A1(n1320), .A2(n1421), .ZN(n1402) );
INV_X1 U1140 ( .A(G237), .ZN(n1421) );
INV_X1 U1141 ( .A(G902), .ZN(n1320) );
endmodule


