//Key = 1010011001100111010010110001111100011000110010110011111000111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;

XNOR2_X1 U785 ( .A(G107), .B(n1103), .ZN(G9) );
NOR2_X1 U786 ( .A1(n1104), .A2(n1105), .ZN(G75) );
NOR4_X1 U787 ( .A1(G953), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1105) );
NOR2_X1 U788 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
NOR2_X1 U789 ( .A1(n1111), .A2(n1112), .ZN(n1109) );
NOR3_X1 U790 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1112) );
NOR2_X1 U791 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NOR2_X1 U792 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR3_X1 U793 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1118) );
NOR2_X1 U794 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U795 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NOR3_X1 U796 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1121) );
NOR2_X1 U797 ( .A1(n1130), .A2(n1131), .ZN(n1120) );
XOR2_X1 U798 ( .A(KEYINPUT25), .B(n1128), .Z(n1130) );
NOR3_X1 U799 ( .A1(n1124), .A2(n1132), .A3(n1128), .ZN(n1116) );
NOR2_X1 U800 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U801 ( .A(n1135), .B(KEYINPUT9), .Z(n1134) );
NAND2_X1 U802 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NOR4_X1 U803 ( .A1(n1138), .A2(n1128), .A3(n1119), .A4(n1124), .ZN(n1111) );
NOR2_X1 U804 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR2_X1 U805 ( .A1(n1141), .A2(n1115), .ZN(n1139) );
NOR3_X1 U806 ( .A1(n1106), .A2(G953), .A3(G952), .ZN(n1104) );
AND4_X1 U807 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1106) );
NOR4_X1 U808 ( .A1(n1136), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1145) );
INV_X1 U809 ( .A(n1149), .ZN(n1148) );
XNOR2_X1 U810 ( .A(n1150), .B(n1151), .ZN(n1147) );
NAND2_X1 U811 ( .A1(KEYINPUT15), .A2(n1152), .ZN(n1150) );
XNOR2_X1 U812 ( .A(KEYINPUT23), .B(n1153), .ZN(n1152) );
NOR2_X1 U813 ( .A1(n1113), .A2(n1154), .ZN(n1144) );
XOR2_X1 U814 ( .A(G475), .B(n1155), .Z(n1154) );
NOR2_X1 U815 ( .A1(KEYINPUT4), .A2(n1156), .ZN(n1155) );
XOR2_X1 U816 ( .A(n1157), .B(n1158), .Z(n1143) );
XOR2_X1 U817 ( .A(n1159), .B(n1160), .Z(n1142) );
XOR2_X1 U818 ( .A(n1161), .B(n1162), .Z(G72) );
XOR2_X1 U819 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR3_X1 U820 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1164) );
NOR2_X1 U821 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XOR2_X1 U822 ( .A(KEYINPUT38), .B(n1170), .Z(n1168) );
NOR2_X1 U823 ( .A1(n1171), .A2(n1172), .ZN(n1166) );
XNOR2_X1 U824 ( .A(n1170), .B(KEYINPUT42), .ZN(n1172) );
XNOR2_X1 U825 ( .A(n1173), .B(n1174), .ZN(n1170) );
XOR2_X1 U826 ( .A(n1175), .B(n1176), .Z(n1173) );
NOR2_X1 U827 ( .A1(KEYINPUT49), .A2(n1177), .ZN(n1176) );
INV_X1 U828 ( .A(G131), .ZN(n1177) );
NAND2_X1 U829 ( .A1(n1178), .A2(n1179), .ZN(n1175) );
NAND2_X1 U830 ( .A1(G125), .A2(n1180), .ZN(n1179) );
XOR2_X1 U831 ( .A(n1181), .B(KEYINPUT19), .Z(n1178) );
NAND2_X1 U832 ( .A1(G140), .A2(n1182), .ZN(n1181) );
INV_X1 U833 ( .A(n1169), .ZN(n1171) );
NOR2_X1 U834 ( .A1(G900), .A2(n1183), .ZN(n1165) );
NAND2_X1 U835 ( .A1(n1183), .A2(n1184), .ZN(n1163) );
NAND3_X1 U836 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
INV_X1 U837 ( .A(n1188), .ZN(n1186) );
XNOR2_X1 U838 ( .A(KEYINPUT60), .B(n1189), .ZN(n1185) );
NAND2_X1 U839 ( .A1(G953), .A2(n1190), .ZN(n1161) );
NAND2_X1 U840 ( .A1(G900), .A2(G227), .ZN(n1190) );
NAND2_X1 U841 ( .A1(n1191), .A2(n1192), .ZN(G69) );
NAND2_X1 U842 ( .A1(n1193), .A2(n1183), .ZN(n1192) );
XOR2_X1 U843 ( .A(n1194), .B(n1195), .Z(n1193) );
NAND2_X1 U844 ( .A1(n1196), .A2(G953), .ZN(n1191) );
NAND2_X1 U845 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NAND2_X1 U846 ( .A1(n1194), .A2(n1199), .ZN(n1198) );
NAND2_X1 U847 ( .A1(G224), .A2(n1200), .ZN(n1197) );
NAND2_X1 U848 ( .A1(G898), .A2(n1194), .ZN(n1200) );
NAND2_X1 U849 ( .A1(n1201), .A2(n1202), .ZN(n1194) );
NAND2_X1 U850 ( .A1(G953), .A2(n1203), .ZN(n1202) );
XOR2_X1 U851 ( .A(n1204), .B(n1205), .Z(n1201) );
NOR2_X1 U852 ( .A1(n1206), .A2(KEYINPUT24), .ZN(n1205) );
NAND2_X1 U853 ( .A1(n1207), .A2(n1208), .ZN(n1204) );
NAND2_X1 U854 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND2_X1 U855 ( .A1(KEYINPUT6), .A2(n1211), .ZN(n1210) );
NAND2_X1 U856 ( .A1(KEYINPUT58), .A2(n1212), .ZN(n1211) );
NAND2_X1 U857 ( .A1(n1213), .A2(n1214), .ZN(n1207) );
NAND2_X1 U858 ( .A1(KEYINPUT58), .A2(n1215), .ZN(n1214) );
NAND2_X1 U859 ( .A1(KEYINPUT6), .A2(n1216), .ZN(n1215) );
INV_X1 U860 ( .A(n1212), .ZN(n1213) );
NOR2_X1 U861 ( .A1(n1217), .A2(n1218), .ZN(G66) );
XOR2_X1 U862 ( .A(n1219), .B(n1220), .Z(n1218) );
NOR2_X1 U863 ( .A1(n1151), .A2(n1221), .ZN(n1220) );
NAND2_X1 U864 ( .A1(KEYINPUT31), .A2(n1222), .ZN(n1219) );
NOR2_X1 U865 ( .A1(n1217), .A2(n1223), .ZN(G63) );
XNOR2_X1 U866 ( .A(n1224), .B(n1225), .ZN(n1223) );
NOR2_X1 U867 ( .A1(n1226), .A2(n1221), .ZN(n1225) );
INV_X1 U868 ( .A(G478), .ZN(n1226) );
NOR2_X1 U869 ( .A1(n1217), .A2(n1227), .ZN(G60) );
XNOR2_X1 U870 ( .A(n1228), .B(n1229), .ZN(n1227) );
NOR2_X1 U871 ( .A1(n1230), .A2(n1221), .ZN(n1229) );
INV_X1 U872 ( .A(G475), .ZN(n1230) );
XOR2_X1 U873 ( .A(G104), .B(n1231), .Z(G6) );
NOR2_X1 U874 ( .A1(n1217), .A2(n1232), .ZN(G57) );
XOR2_X1 U875 ( .A(n1233), .B(n1234), .Z(n1232) );
XOR2_X1 U876 ( .A(n1235), .B(n1236), .Z(n1234) );
NOR2_X1 U877 ( .A1(n1237), .A2(n1221), .ZN(n1236) );
INV_X1 U878 ( .A(G472), .ZN(n1237) );
NAND3_X1 U879 ( .A1(n1238), .A2(n1239), .A3(KEYINPUT44), .ZN(n1235) );
NAND3_X1 U880 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1239) );
INV_X1 U881 ( .A(KEYINPUT30), .ZN(n1242) );
NAND2_X1 U882 ( .A1(n1243), .A2(KEYINPUT30), .ZN(n1238) );
NOR2_X1 U883 ( .A1(n1217), .A2(n1244), .ZN(G54) );
XOR2_X1 U884 ( .A(n1245), .B(n1246), .Z(n1244) );
XOR2_X1 U885 ( .A(n1247), .B(n1248), .Z(n1246) );
NOR2_X1 U886 ( .A1(n1160), .A2(n1221), .ZN(n1248) );
NOR2_X1 U887 ( .A1(n1249), .A2(n1250), .ZN(n1247) );
XOR2_X1 U888 ( .A(KEYINPUT61), .B(n1251), .Z(n1250) );
NOR2_X1 U889 ( .A1(n1252), .A2(n1253), .ZN(G51) );
XNOR2_X1 U890 ( .A(n1217), .B(KEYINPUT22), .ZN(n1253) );
NOR2_X1 U891 ( .A1(n1183), .A2(G952), .ZN(n1217) );
XOR2_X1 U892 ( .A(n1254), .B(n1255), .Z(n1252) );
XOR2_X1 U893 ( .A(n1256), .B(n1257), .Z(n1254) );
NOR2_X1 U894 ( .A1(n1158), .A2(n1221), .ZN(n1257) );
NAND2_X1 U895 ( .A1(G902), .A2(n1108), .ZN(n1221) );
NAND4_X1 U896 ( .A1(n1195), .A2(n1187), .A3(n1258), .A4(n1189), .ZN(n1108) );
XOR2_X1 U897 ( .A(KEYINPUT28), .B(n1188), .Z(n1258) );
AND4_X1 U898 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1187) );
NOR2_X1 U899 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
NOR2_X1 U900 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NOR3_X1 U901 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(n1263) );
NOR2_X1 U902 ( .A1(KEYINPUT29), .A2(n1270), .ZN(n1269) );
NOR3_X1 U903 ( .A1(n1271), .A2(n1272), .A3(n1124), .ZN(n1270) );
INV_X1 U904 ( .A(n1273), .ZN(n1124) );
AND2_X1 U905 ( .A1(n1266), .A2(KEYINPUT29), .ZN(n1268) );
NAND3_X1 U906 ( .A1(n1274), .A2(n1271), .A3(n1275), .ZN(n1261) );
NAND2_X1 U907 ( .A1(n1276), .A2(n1277), .ZN(n1274) );
NAND2_X1 U908 ( .A1(n1140), .A2(n1278), .ZN(n1276) );
XOR2_X1 U909 ( .A(KEYINPUT11), .B(n1279), .Z(n1278) );
AND4_X1 U910 ( .A1(n1280), .A2(n1281), .A3(n1282), .A4(n1283), .ZN(n1195) );
NOR4_X1 U911 ( .A1(n1284), .A2(n1285), .A3(n1286), .A4(n1231), .ZN(n1283) );
AND4_X1 U912 ( .A1(n1140), .A2(n1275), .A3(n1287), .A4(n1288), .ZN(n1231) );
NOR3_X1 U913 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1282) );
AND4_X1 U914 ( .A1(KEYINPUT32), .A2(n1292), .A3(n1113), .A4(n1128), .ZN(n1291) );
NOR2_X1 U915 ( .A1(KEYINPUT32), .A2(n1103), .ZN(n1290) );
NAND3_X1 U916 ( .A1(n1287), .A2(n1113), .A3(n1292), .ZN(n1103) );
NOR2_X1 U917 ( .A1(n1293), .A2(n1131), .ZN(n1289) );
XOR2_X1 U918 ( .A(n1294), .B(KEYINPUT16), .Z(n1293) );
INV_X1 U919 ( .A(n1295), .ZN(n1281) );
NAND2_X1 U920 ( .A1(n1296), .A2(n1297), .ZN(n1256) );
NAND4_X1 U921 ( .A1(KEYINPUT27), .A2(n1240), .A3(n1298), .A4(n1299), .ZN(n1297) );
NAND2_X1 U922 ( .A1(n1300), .A2(n1182), .ZN(n1299) );
NAND2_X1 U923 ( .A1(n1301), .A2(G125), .ZN(n1298) );
NAND3_X1 U924 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1296) );
NAND2_X1 U925 ( .A1(KEYINPUT27), .A2(n1240), .ZN(n1304) );
NAND2_X1 U926 ( .A1(n1301), .A2(n1182), .ZN(n1303) );
XOR2_X1 U927 ( .A(KEYINPUT46), .B(n1305), .Z(n1301) );
NAND2_X1 U928 ( .A1(n1300), .A2(G125), .ZN(n1302) );
XNOR2_X1 U929 ( .A(KEYINPUT52), .B(n1305), .ZN(n1300) );
XOR2_X1 U930 ( .A(n1306), .B(n1307), .Z(G48) );
NOR2_X1 U931 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NOR2_X1 U932 ( .A1(KEYINPUT48), .A2(n1310), .ZN(n1306) );
XOR2_X1 U933 ( .A(n1311), .B(n1312), .Z(G45) );
NAND4_X1 U934 ( .A1(n1313), .A2(n1271), .A3(n1314), .A4(n1315), .ZN(n1312) );
OR2_X1 U935 ( .A1(n1316), .A2(n1275), .ZN(n1315) );
NAND2_X1 U936 ( .A1(n1317), .A2(n1316), .ZN(n1314) );
INV_X1 U937 ( .A(KEYINPUT2), .ZN(n1316) );
NAND2_X1 U938 ( .A1(n1133), .A2(n1131), .ZN(n1317) );
INV_X1 U939 ( .A(n1277), .ZN(n1313) );
NAND2_X1 U940 ( .A1(n1318), .A2(n1125), .ZN(n1277) );
INV_X1 U941 ( .A(n1319), .ZN(n1318) );
XOR2_X1 U942 ( .A(n1180), .B(n1259), .Z(G42) );
NAND3_X1 U943 ( .A1(n1140), .A2(n1126), .A3(n1320), .ZN(n1259) );
NAND2_X1 U944 ( .A1(n1321), .A2(n1322), .ZN(G39) );
NAND2_X1 U945 ( .A1(G137), .A2(n1260), .ZN(n1322) );
XOR2_X1 U946 ( .A(n1323), .B(KEYINPUT12), .Z(n1321) );
OR2_X1 U947 ( .A1(n1260), .A2(G137), .ZN(n1323) );
NAND2_X1 U948 ( .A1(n1320), .A2(n1324), .ZN(n1260) );
INV_X1 U949 ( .A(n1266), .ZN(n1320) );
XNOR2_X1 U950 ( .A(G134), .B(n1325), .ZN(G36) );
OR2_X1 U951 ( .A1(n1266), .A2(n1267), .ZN(n1325) );
NAND3_X1 U952 ( .A1(n1133), .A2(n1271), .A3(n1273), .ZN(n1266) );
XOR2_X1 U953 ( .A(n1326), .B(n1327), .Z(G33) );
XOR2_X1 U954 ( .A(KEYINPUT62), .B(G131), .Z(n1327) );
NAND2_X1 U955 ( .A1(n1273), .A2(n1328), .ZN(n1326) );
XOR2_X1 U956 ( .A(KEYINPUT34), .B(n1329), .Z(n1328) );
NOR3_X1 U957 ( .A1(n1265), .A2(n1330), .A3(n1331), .ZN(n1329) );
XOR2_X1 U958 ( .A(n1272), .B(KEYINPUT57), .Z(n1331) );
NOR2_X1 U959 ( .A1(n1129), .A2(n1146), .ZN(n1273) );
INV_X1 U960 ( .A(n1127), .ZN(n1146) );
XOR2_X1 U961 ( .A(G128), .B(n1188), .Z(G30) );
NOR3_X1 U962 ( .A1(n1115), .A2(n1141), .A3(n1309), .ZN(n1188) );
NAND3_X1 U963 ( .A1(n1275), .A2(n1271), .A3(n1279), .ZN(n1309) );
XOR2_X1 U964 ( .A(n1332), .B(n1280), .Z(G3) );
NAND3_X1 U965 ( .A1(n1292), .A2(n1125), .A3(n1141), .ZN(n1280) );
INV_X1 U966 ( .A(n1333), .ZN(n1292) );
XOR2_X1 U967 ( .A(n1189), .B(n1334), .Z(G27) );
XOR2_X1 U968 ( .A(n1182), .B(KEYINPUT21), .Z(n1334) );
NAND3_X1 U969 ( .A1(n1140), .A2(n1335), .A3(n1336), .ZN(n1189) );
NOR3_X1 U970 ( .A1(n1131), .A2(n1330), .A3(n1337), .ZN(n1336) );
INV_X1 U971 ( .A(n1271), .ZN(n1330) );
NAND2_X1 U972 ( .A1(n1110), .A2(n1338), .ZN(n1271) );
NAND4_X1 U973 ( .A1(G953), .A2(G902), .A3(n1339), .A4(n1340), .ZN(n1338) );
INV_X1 U974 ( .A(G900), .ZN(n1340) );
NAND2_X1 U975 ( .A1(n1341), .A2(n1342), .ZN(G24) );
NAND2_X1 U976 ( .A1(n1295), .A2(n1343), .ZN(n1342) );
XOR2_X1 U977 ( .A(KEYINPUT35), .B(n1344), .Z(n1341) );
NOR2_X1 U978 ( .A1(n1295), .A2(n1343), .ZN(n1344) );
NOR3_X1 U979 ( .A1(n1345), .A2(n1128), .A3(n1319), .ZN(n1295) );
NAND2_X1 U980 ( .A1(n1346), .A2(n1115), .ZN(n1319) );
XOR2_X1 U981 ( .A(KEYINPUT55), .B(n1113), .Z(n1346) );
INV_X1 U982 ( .A(n1287), .ZN(n1128) );
NAND2_X1 U983 ( .A1(n1347), .A2(n1348), .ZN(n1287) );
NAND2_X1 U984 ( .A1(n1125), .A2(n1349), .ZN(n1348) );
NAND3_X1 U985 ( .A1(n1350), .A2(n1149), .A3(KEYINPUT36), .ZN(n1347) );
XOR2_X1 U986 ( .A(G119), .B(n1351), .Z(G21) );
NOR2_X1 U987 ( .A1(n1131), .A2(n1294), .ZN(n1351) );
NAND3_X1 U988 ( .A1(n1335), .A2(n1288), .A3(n1324), .ZN(n1294) );
AND3_X1 U989 ( .A1(n1352), .A2(n1141), .A3(n1279), .ZN(n1324) );
XOR2_X1 U990 ( .A(G116), .B(n1286), .Z(G18) );
NOR2_X1 U991 ( .A1(n1267), .A2(n1345), .ZN(n1286) );
NAND3_X1 U992 ( .A1(n1352), .A2(n1113), .A3(n1125), .ZN(n1267) );
XOR2_X1 U993 ( .A(G113), .B(n1285), .Z(G15) );
NOR2_X1 U994 ( .A1(n1345), .A2(n1265), .ZN(n1285) );
NAND2_X1 U995 ( .A1(n1140), .A2(n1125), .ZN(n1265) );
NOR2_X1 U996 ( .A1(n1353), .A2(n1149), .ZN(n1125) );
INV_X1 U997 ( .A(n1308), .ZN(n1140) );
NAND2_X1 U998 ( .A1(n1141), .A2(n1115), .ZN(n1308) );
INV_X1 U999 ( .A(n1352), .ZN(n1115) );
NAND3_X1 U1000 ( .A1(n1354), .A2(n1288), .A3(n1335), .ZN(n1345) );
INV_X1 U1001 ( .A(n1119), .ZN(n1335) );
NAND2_X1 U1002 ( .A1(n1137), .A2(n1355), .ZN(n1119) );
INV_X1 U1003 ( .A(n1131), .ZN(n1354) );
XOR2_X1 U1004 ( .A(G110), .B(n1284), .Z(G12) );
NOR3_X1 U1005 ( .A1(n1333), .A2(n1337), .A3(n1113), .ZN(n1284) );
INV_X1 U1006 ( .A(n1141), .ZN(n1113) );
XOR2_X1 U1007 ( .A(n1356), .B(G478), .Z(n1141) );
NAND2_X1 U1008 ( .A1(n1357), .A2(n1224), .ZN(n1356) );
XNOR2_X1 U1009 ( .A(n1358), .B(n1359), .ZN(n1224) );
XOR2_X1 U1010 ( .A(G107), .B(n1360), .Z(n1359) );
XOR2_X1 U1011 ( .A(KEYINPUT59), .B(G116), .Z(n1360) );
XOR2_X1 U1012 ( .A(n1361), .B(n1362), .Z(n1358) );
XOR2_X1 U1013 ( .A(n1363), .B(n1364), .Z(n1361) );
AND2_X1 U1014 ( .A1(n1365), .A2(G217), .ZN(n1364) );
NAND3_X1 U1015 ( .A1(n1366), .A2(n1367), .A3(n1368), .ZN(n1363) );
NAND2_X1 U1016 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
NAND2_X1 U1017 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
XOR2_X1 U1018 ( .A(n1373), .B(G143), .Z(n1369) );
OR2_X1 U1019 ( .A1(n1371), .A2(KEYINPUT14), .ZN(n1367) );
NAND4_X1 U1020 ( .A1(n1371), .A2(n1372), .A3(n1374), .A4(KEYINPUT14), .ZN(n1366) );
XOR2_X1 U1021 ( .A(G143), .B(G128), .Z(n1374) );
INV_X1 U1022 ( .A(KEYINPUT45), .ZN(n1372) );
XNOR2_X1 U1023 ( .A(G134), .B(KEYINPUT43), .ZN(n1371) );
INV_X1 U1024 ( .A(n1126), .ZN(n1337) );
NAND2_X1 U1025 ( .A1(n1375), .A2(n1376), .ZN(n1126) );
NAND2_X1 U1026 ( .A1(n1279), .A2(n1349), .ZN(n1376) );
INV_X1 U1027 ( .A(KEYINPUT36), .ZN(n1349) );
NOR2_X1 U1028 ( .A1(n1149), .A2(n1350), .ZN(n1279) );
NAND3_X1 U1029 ( .A1(n1353), .A2(n1149), .A3(KEYINPUT36), .ZN(n1375) );
XOR2_X1 U1030 ( .A(n1377), .B(G472), .Z(n1149) );
NAND2_X1 U1031 ( .A1(n1357), .A2(n1378), .ZN(n1377) );
XOR2_X1 U1032 ( .A(n1243), .B(n1379), .Z(n1378) );
INV_X1 U1033 ( .A(n1233), .ZN(n1379) );
XOR2_X1 U1034 ( .A(n1380), .B(n1381), .Z(n1233) );
XOR2_X1 U1035 ( .A(n1332), .B(n1382), .Z(n1381) );
NAND2_X1 U1036 ( .A1(n1383), .A2(G210), .ZN(n1382) );
XOR2_X1 U1037 ( .A(n1384), .B(n1385), .Z(n1380) );
XOR2_X1 U1038 ( .A(G119), .B(G116), .Z(n1385) );
XOR2_X1 U1039 ( .A(n1240), .B(n1241), .Z(n1243) );
INV_X1 U1040 ( .A(n1386), .ZN(n1240) );
INV_X1 U1041 ( .A(n1350), .ZN(n1353) );
XNOR2_X1 U1042 ( .A(n1387), .B(n1151), .ZN(n1350) );
NAND2_X1 U1043 ( .A1(G217), .A2(n1388), .ZN(n1151) );
XOR2_X1 U1044 ( .A(n1153), .B(KEYINPUT3), .Z(n1387) );
NAND2_X1 U1045 ( .A1(n1222), .A2(n1357), .ZN(n1153) );
XOR2_X1 U1046 ( .A(n1389), .B(n1390), .Z(n1222) );
XOR2_X1 U1047 ( .A(n1391), .B(n1392), .Z(n1390) );
XNOR2_X1 U1048 ( .A(n1393), .B(n1394), .ZN(n1392) );
NOR2_X1 U1049 ( .A1(G146), .A2(KEYINPUT8), .ZN(n1394) );
NAND2_X1 U1050 ( .A1(KEYINPUT5), .A2(n1395), .ZN(n1393) );
XNOR2_X1 U1051 ( .A(G137), .B(n1396), .ZN(n1395) );
NAND2_X1 U1052 ( .A1(n1365), .A2(G221), .ZN(n1396) );
AND2_X1 U1053 ( .A1(G234), .A2(n1183), .ZN(n1365) );
XOR2_X1 U1054 ( .A(n1397), .B(n1398), .Z(n1389) );
XOR2_X1 U1055 ( .A(KEYINPUT10), .B(G110), .Z(n1398) );
NAND2_X1 U1056 ( .A1(n1399), .A2(n1400), .ZN(n1397) );
NAND2_X1 U1057 ( .A1(G128), .A2(n1401), .ZN(n1400) );
XOR2_X1 U1058 ( .A(KEYINPUT0), .B(n1402), .Z(n1399) );
NOR2_X1 U1059 ( .A1(G128), .A2(n1401), .ZN(n1402) );
NAND3_X1 U1060 ( .A1(n1352), .A2(n1288), .A3(n1275), .ZN(n1333) );
NOR2_X1 U1061 ( .A1(n1272), .A2(n1131), .ZN(n1275) );
NAND2_X1 U1062 ( .A1(n1129), .A2(n1127), .ZN(n1131) );
NAND2_X1 U1063 ( .A1(G214), .A2(n1403), .ZN(n1127) );
XOR2_X1 U1064 ( .A(n1404), .B(n1158), .Z(n1129) );
NAND2_X1 U1065 ( .A1(G210), .A2(n1403), .ZN(n1158) );
NAND2_X1 U1066 ( .A1(n1405), .A2(n1406), .ZN(n1403) );
INV_X1 U1067 ( .A(G237), .ZN(n1405) );
NAND2_X1 U1068 ( .A1(KEYINPUT13), .A2(n1157), .ZN(n1404) );
AND2_X1 U1069 ( .A1(n1407), .A2(n1357), .ZN(n1157) );
XOR2_X1 U1070 ( .A(n1408), .B(n1409), .Z(n1407) );
XOR2_X1 U1071 ( .A(n1182), .B(n1386), .Z(n1409) );
NAND2_X1 U1072 ( .A1(n1410), .A2(n1411), .ZN(n1386) );
NAND2_X1 U1073 ( .A1(n1412), .A2(n1373), .ZN(n1411) );
XOR2_X1 U1074 ( .A(KEYINPUT54), .B(n1413), .Z(n1410) );
NOR2_X1 U1075 ( .A1(n1373), .A2(n1412), .ZN(n1413) );
NAND3_X1 U1076 ( .A1(n1414), .A2(n1415), .A3(n1416), .ZN(n1412) );
OR2_X1 U1077 ( .A1(n1417), .A2(KEYINPUT26), .ZN(n1415) );
NAND2_X1 U1078 ( .A1(KEYINPUT26), .A2(G146), .ZN(n1414) );
INV_X1 U1079 ( .A(G128), .ZN(n1373) );
INV_X1 U1080 ( .A(G125), .ZN(n1182) );
XNOR2_X1 U1081 ( .A(n1255), .B(n1305), .ZN(n1408) );
NOR2_X1 U1082 ( .A1(n1199), .A2(G953), .ZN(n1305) );
INV_X1 U1083 ( .A(G224), .ZN(n1199) );
XOR2_X1 U1084 ( .A(n1206), .B(n1418), .Z(n1255) );
NOR2_X1 U1085 ( .A1(KEYINPUT18), .A2(n1419), .ZN(n1418) );
XOR2_X1 U1086 ( .A(n1212), .B(n1420), .Z(n1419) );
NOR2_X1 U1087 ( .A1(KEYINPUT7), .A2(n1209), .ZN(n1420) );
INV_X1 U1088 ( .A(n1216), .ZN(n1209) );
XOR2_X1 U1089 ( .A(n1421), .B(n1422), .Z(n1216) );
XOR2_X1 U1090 ( .A(n1423), .B(n1424), .Z(n1422) );
NAND2_X1 U1091 ( .A1(KEYINPUT53), .A2(n1401), .ZN(n1424) );
INV_X1 U1092 ( .A(G119), .ZN(n1401) );
INV_X1 U1093 ( .A(G116), .ZN(n1423) );
NAND2_X1 U1094 ( .A1(KEYINPUT41), .A2(n1384), .ZN(n1421) );
XOR2_X1 U1095 ( .A(n1332), .B(n1425), .Z(n1212) );
INV_X1 U1096 ( .A(G101), .ZN(n1332) );
AND3_X1 U1097 ( .A1(n1426), .A2(n1427), .A3(n1428), .ZN(n1206) );
OR2_X1 U1098 ( .A1(n1362), .A2(KEYINPUT50), .ZN(n1428) );
NAND4_X1 U1099 ( .A1(KEYINPUT20), .A2(n1362), .A3(KEYINPUT50), .A4(G110), .ZN(n1427) );
NAND2_X1 U1100 ( .A1(n1429), .A2(n1430), .ZN(n1426) );
NAND2_X1 U1101 ( .A1(KEYINPUT20), .A2(n1362), .ZN(n1429) );
INV_X1 U1102 ( .A(n1431), .ZN(n1362) );
INV_X1 U1103 ( .A(n1133), .ZN(n1272) );
NOR2_X1 U1104 ( .A1(n1137), .A2(n1136), .ZN(n1133) );
INV_X1 U1105 ( .A(n1355), .ZN(n1136) );
NAND2_X1 U1106 ( .A1(G221), .A2(n1388), .ZN(n1355) );
NAND2_X1 U1107 ( .A1(G234), .A2(n1406), .ZN(n1388) );
XNOR2_X1 U1108 ( .A(n1160), .B(n1432), .ZN(n1137) );
NOR2_X1 U1109 ( .A1(n1159), .A2(KEYINPUT33), .ZN(n1432) );
AND2_X1 U1110 ( .A1(n1433), .A2(n1357), .ZN(n1159) );
XNOR2_X1 U1111 ( .A(n1245), .B(n1434), .ZN(n1433) );
NOR2_X1 U1112 ( .A1(n1249), .A2(n1435), .ZN(n1434) );
XNOR2_X1 U1113 ( .A(n1251), .B(KEYINPUT47), .ZN(n1435) );
NOR2_X1 U1114 ( .A1(n1180), .A2(G110), .ZN(n1251) );
NOR2_X1 U1115 ( .A1(n1430), .A2(G140), .ZN(n1249) );
INV_X1 U1116 ( .A(G110), .ZN(n1430) );
XNOR2_X1 U1117 ( .A(n1436), .B(n1437), .ZN(n1245) );
XNOR2_X1 U1118 ( .A(n1241), .B(n1438), .ZN(n1437) );
XOR2_X1 U1119 ( .A(n1439), .B(n1440), .Z(n1438) );
NOR2_X1 U1120 ( .A1(KEYINPUT37), .A2(n1441), .ZN(n1440) );
XOR2_X1 U1121 ( .A(KEYINPUT63), .B(G101), .Z(n1441) );
NAND2_X1 U1122 ( .A1(G227), .A2(n1183), .ZN(n1439) );
XOR2_X1 U1123 ( .A(n1174), .B(G131), .Z(n1241) );
XOR2_X1 U1124 ( .A(G134), .B(n1442), .Z(n1174) );
XOR2_X1 U1125 ( .A(KEYINPUT39), .B(G137), .Z(n1442) );
XOR2_X1 U1126 ( .A(n1169), .B(n1425), .Z(n1436) );
XOR2_X1 U1127 ( .A(G104), .B(G107), .Z(n1425) );
XOR2_X1 U1128 ( .A(n1443), .B(G128), .Z(n1169) );
NAND3_X1 U1129 ( .A1(n1444), .A2(n1445), .A3(n1446), .ZN(n1443) );
XOR2_X1 U1130 ( .A(n1447), .B(KEYINPUT40), .Z(n1446) );
NAND2_X1 U1131 ( .A1(n1448), .A2(n1449), .ZN(n1447) );
OR2_X1 U1132 ( .A1(n1417), .A2(KEYINPUT51), .ZN(n1449) );
NAND3_X1 U1133 ( .A1(G143), .A2(n1310), .A3(KEYINPUT51), .ZN(n1448) );
OR2_X1 U1134 ( .A1(n1416), .A2(KEYINPUT51), .ZN(n1445) );
NAND3_X1 U1135 ( .A1(G146), .A2(n1311), .A3(KEYINPUT51), .ZN(n1444) );
INV_X1 U1136 ( .A(G469), .ZN(n1160) );
NAND2_X1 U1137 ( .A1(n1110), .A2(n1450), .ZN(n1288) );
NAND4_X1 U1138 ( .A1(G953), .A2(G902), .A3(n1339), .A4(n1203), .ZN(n1450) );
INV_X1 U1139 ( .A(G898), .ZN(n1203) );
NAND3_X1 U1140 ( .A1(n1339), .A2(n1183), .A3(G952), .ZN(n1110) );
INV_X1 U1141 ( .A(G953), .ZN(n1183) );
NAND2_X1 U1142 ( .A1(G237), .A2(G234), .ZN(n1339) );
XOR2_X1 U1143 ( .A(n1156), .B(G475), .Z(n1352) );
NAND2_X1 U1144 ( .A1(n1228), .A2(n1357), .ZN(n1156) );
XOR2_X1 U1145 ( .A(n1406), .B(KEYINPUT56), .Z(n1357) );
INV_X1 U1146 ( .A(G902), .ZN(n1406) );
XNOR2_X1 U1147 ( .A(n1451), .B(n1452), .ZN(n1228) );
XNOR2_X1 U1148 ( .A(n1391), .B(n1453), .ZN(n1452) );
NAND2_X1 U1149 ( .A1(n1454), .A2(n1455), .ZN(n1453) );
NAND2_X1 U1150 ( .A1(n1456), .A2(n1457), .ZN(n1455) );
NAND2_X1 U1151 ( .A1(n1416), .A2(n1417), .ZN(n1457) );
NAND2_X1 U1152 ( .A1(n1311), .A2(n1310), .ZN(n1417) );
INV_X1 U1153 ( .A(G146), .ZN(n1310) );
INV_X1 U1154 ( .A(G143), .ZN(n1311) );
NAND2_X1 U1155 ( .A1(G146), .A2(G143), .ZN(n1416) );
NAND2_X1 U1156 ( .A1(n1458), .A2(n1459), .ZN(n1454) );
INV_X1 U1157 ( .A(n1456), .ZN(n1459) );
XNOR2_X1 U1158 ( .A(n1384), .B(G131), .ZN(n1456) );
INV_X1 U1159 ( .A(G113), .ZN(n1384) );
XOR2_X1 U1160 ( .A(G146), .B(G143), .Z(n1458) );
XNOR2_X1 U1161 ( .A(n1180), .B(G125), .ZN(n1391) );
INV_X1 U1162 ( .A(G140), .ZN(n1180) );
XOR2_X1 U1163 ( .A(n1460), .B(n1461), .Z(n1451) );
AND2_X1 U1164 ( .A1(G214), .A2(n1383), .ZN(n1461) );
NOR2_X1 U1165 ( .A1(G953), .A2(G237), .ZN(n1383) );
XOR2_X1 U1166 ( .A(n1462), .B(G104), .Z(n1460) );
NAND2_X1 U1167 ( .A1(KEYINPUT17), .A2(n1431), .ZN(n1462) );
XOR2_X1 U1168 ( .A(n1343), .B(KEYINPUT1), .Z(n1431) );
INV_X1 U1169 ( .A(G122), .ZN(n1343) );
endmodule


