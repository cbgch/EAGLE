//Key = 0110010010010101010010111000111110101010010110001001110110001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266;

XOR2_X1 U701 ( .A(n966), .B(n967), .Z(G9) );
NAND2_X1 U702 ( .A1(KEYINPUT24), .A2(n968), .ZN(n966) );
NOR2_X1 U703 ( .A1(n969), .A2(n970), .ZN(G75) );
XOR2_X1 U704 ( .A(KEYINPUT7), .B(n971), .Z(n970) );
NOR3_X1 U705 ( .A1(n972), .A2(n973), .A3(n974), .ZN(n971) );
NOR2_X1 U706 ( .A1(n975), .A2(n976), .ZN(n973) );
NOR2_X1 U707 ( .A1(n977), .A2(n978), .ZN(n975) );
NOR3_X1 U708 ( .A1(n979), .A2(n980), .A3(n981), .ZN(n978) );
NOR2_X1 U709 ( .A1(n982), .A2(n983), .ZN(n981) );
NOR2_X1 U710 ( .A1(n984), .A2(n985), .ZN(n983) );
NOR2_X1 U711 ( .A1(n986), .A2(n987), .ZN(n984) );
NOR2_X1 U712 ( .A1(n988), .A2(n989), .ZN(n987) );
NOR2_X1 U713 ( .A1(n990), .A2(n991), .ZN(n988) );
NOR2_X1 U714 ( .A1(n992), .A2(n993), .ZN(n990) );
NOR2_X1 U715 ( .A1(n994), .A2(n995), .ZN(n986) );
NOR2_X1 U716 ( .A1(n996), .A2(n997), .ZN(n994) );
NOR3_X1 U717 ( .A1(n995), .A2(n998), .A3(n989), .ZN(n982) );
NOR2_X1 U718 ( .A1(n999), .A2(n1000), .ZN(n998) );
NOR4_X1 U719 ( .A1(n1001), .A2(n985), .A3(n989), .A4(n995), .ZN(n977) );
NOR2_X1 U720 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NOR2_X1 U721 ( .A1(n979), .A2(n1004), .ZN(n1002) );
NOR2_X1 U722 ( .A1(G952), .A2(n974), .ZN(n969) );
NAND2_X1 U723 ( .A1(n1005), .A2(n1006), .ZN(n974) );
NAND2_X1 U724 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NOR4_X1 U725 ( .A1(n1009), .A2(n980), .A3(n1010), .A4(n1011), .ZN(n1008) );
XOR2_X1 U726 ( .A(n1012), .B(n1013), .Z(n1010) );
XOR2_X1 U727 ( .A(n1014), .B(KEYINPUT40), .Z(n1012) );
NOR4_X1 U728 ( .A1(n979), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1007) );
XNOR2_X1 U729 ( .A(KEYINPUT59), .B(n1018), .ZN(n1017) );
XOR2_X1 U730 ( .A(n1019), .B(n1020), .Z(n1016) );
NAND2_X1 U731 ( .A1(n1021), .A2(n1022), .ZN(G72) );
NAND2_X1 U732 ( .A1(n1023), .A2(n1005), .ZN(n1022) );
NAND2_X1 U733 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND2_X1 U734 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U735 ( .A1(n1028), .A2(n1029), .ZN(n1024) );
INV_X1 U736 ( .A(n1026), .ZN(n1028) );
NAND2_X1 U737 ( .A1(n1030), .A2(n1031), .ZN(n1026) );
NAND2_X1 U738 ( .A1(n1032), .A2(G953), .ZN(n1021) );
XOR2_X1 U739 ( .A(n1033), .B(n1029), .Z(n1032) );
XOR2_X1 U740 ( .A(n1027), .B(KEYINPUT53), .Z(n1029) );
NAND2_X1 U741 ( .A1(n1034), .A2(n1035), .ZN(n1027) );
NAND2_X1 U742 ( .A1(G953), .A2(n1036), .ZN(n1035) );
XOR2_X1 U743 ( .A(n1037), .B(n1038), .Z(n1034) );
XNOR2_X1 U744 ( .A(KEYINPUT47), .B(n1039), .ZN(n1038) );
NOR3_X1 U745 ( .A1(KEYINPUT45), .A2(n1040), .A3(n1041), .ZN(n1039) );
NOR2_X1 U746 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
XNOR2_X1 U747 ( .A(n1044), .B(KEYINPUT11), .ZN(n1043) );
NOR2_X1 U748 ( .A1(G131), .A2(n1045), .ZN(n1040) );
XNOR2_X1 U749 ( .A(KEYINPUT56), .B(n1046), .ZN(n1045) );
INV_X1 U750 ( .A(n1044), .ZN(n1046) );
XNOR2_X1 U751 ( .A(n1047), .B(n1048), .ZN(n1044) );
NAND2_X1 U752 ( .A1(G900), .A2(G227), .ZN(n1033) );
XOR2_X1 U753 ( .A(n1049), .B(n1050), .Z(G69) );
XOR2_X1 U754 ( .A(n1051), .B(n1052), .Z(n1050) );
NOR2_X1 U755 ( .A1(G953), .A2(n1053), .ZN(n1052) );
NOR2_X1 U756 ( .A1(n1054), .A2(n1055), .ZN(n1051) );
XOR2_X1 U757 ( .A(KEYINPUT63), .B(n1056), .Z(n1055) );
NOR2_X1 U758 ( .A1(G898), .A2(n1005), .ZN(n1056) );
XOR2_X1 U759 ( .A(n1057), .B(n1058), .Z(n1054) );
NAND2_X1 U760 ( .A1(n1059), .A2(KEYINPUT55), .ZN(n1057) );
XNOR2_X1 U761 ( .A(G110), .B(G122), .ZN(n1059) );
NOR2_X1 U762 ( .A1(n1060), .A2(n1005), .ZN(n1049) );
NOR2_X1 U763 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U764 ( .A1(n1063), .A2(n1064), .ZN(G66) );
XNOR2_X1 U765 ( .A(n1065), .B(n1066), .ZN(n1064) );
NOR2_X1 U766 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U767 ( .A1(n1063), .A2(n1069), .ZN(G63) );
XNOR2_X1 U768 ( .A(n1070), .B(n1071), .ZN(n1069) );
NOR2_X1 U769 ( .A1(n1072), .A2(n1068), .ZN(n1070) );
NOR2_X1 U770 ( .A1(n1063), .A2(n1073), .ZN(G60) );
XNOR2_X1 U771 ( .A(n1074), .B(n1075), .ZN(n1073) );
NOR2_X1 U772 ( .A1(n1076), .A2(n1068), .ZN(n1075) );
XOR2_X1 U773 ( .A(n1077), .B(n1078), .Z(G6) );
XOR2_X1 U774 ( .A(KEYINPUT58), .B(G104), .Z(n1078) );
NOR4_X1 U775 ( .A1(n1079), .A2(n1080), .A3(n985), .A4(n1081), .ZN(n1077) );
XNOR2_X1 U776 ( .A(n991), .B(KEYINPUT0), .ZN(n1079) );
NOR2_X1 U777 ( .A1(n1063), .A2(n1082), .ZN(G57) );
XOR2_X1 U778 ( .A(n1083), .B(n1084), .Z(n1082) );
XNOR2_X1 U779 ( .A(n1085), .B(n1086), .ZN(n1084) );
XOR2_X1 U780 ( .A(n1087), .B(n1088), .Z(n1086) );
NOR3_X1 U781 ( .A1(n1068), .A2(KEYINPUT10), .A3(n1089), .ZN(n1088) );
XNOR2_X1 U782 ( .A(n1090), .B(n1091), .ZN(n1083) );
NOR2_X1 U783 ( .A1(n1063), .A2(n1092), .ZN(G54) );
XOR2_X1 U784 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U785 ( .A1(n1095), .A2(n1068), .ZN(n1094) );
NAND3_X1 U786 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1093) );
NAND2_X1 U787 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
INV_X1 U788 ( .A(KEYINPUT31), .ZN(n1100) );
NAND3_X1 U789 ( .A1(KEYINPUT31), .A2(n1101), .A3(n1102), .ZN(n1097) );
OR2_X1 U790 ( .A1(n1102), .A2(n1101), .ZN(n1096) );
NOR2_X1 U791 ( .A1(n1103), .A2(n1099), .ZN(n1101) );
XOR2_X1 U792 ( .A(n1104), .B(n1047), .Z(n1099) );
XOR2_X1 U793 ( .A(n1087), .B(n1105), .Z(n1104) );
NOR2_X1 U794 ( .A1(KEYINPUT19), .A2(n1106), .ZN(n1105) );
XOR2_X1 U795 ( .A(n1107), .B(n1108), .Z(n1106) );
INV_X1 U796 ( .A(KEYINPUT61), .ZN(n1103) );
NOR2_X1 U797 ( .A1(n1063), .A2(n1109), .ZN(G51) );
XOR2_X1 U798 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U799 ( .A1(n1112), .A2(n1068), .ZN(n1111) );
NAND2_X1 U800 ( .A1(G902), .A2(n972), .ZN(n1068) );
NAND3_X1 U801 ( .A1(n1053), .A2(n1030), .A3(n1113), .ZN(n972) );
XOR2_X1 U802 ( .A(n1031), .B(KEYINPUT6), .Z(n1113) );
AND4_X1 U803 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1030) );
AND4_X1 U804 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1117) );
OR2_X1 U805 ( .A1(n1122), .A2(n995), .ZN(n1116) );
NAND4_X1 U806 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n991), .ZN(n1114) );
XNOR2_X1 U807 ( .A(n997), .B(KEYINPUT13), .ZN(n1123) );
AND2_X1 U808 ( .A1(n1126), .A2(n1127), .ZN(n1053) );
NOR4_X1 U809 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1127) );
INV_X1 U810 ( .A(n1132), .ZN(n1128) );
NOR4_X1 U811 ( .A1(n967), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1126) );
AND3_X1 U812 ( .A1(n997), .A2(n1136), .A3(n1137), .ZN(n1135) );
AND3_X1 U813 ( .A1(n996), .A2(n1136), .A3(n1137), .ZN(n967) );
INV_X1 U814 ( .A(G210), .ZN(n1112) );
NOR2_X1 U815 ( .A1(n1005), .A2(G952), .ZN(n1063) );
XOR2_X1 U816 ( .A(G146), .B(n1138), .Z(G48) );
NOR2_X1 U817 ( .A1(KEYINPUT42), .A2(n1031), .ZN(n1138) );
NAND3_X1 U818 ( .A1(n997), .A2(n991), .A3(n1139), .ZN(n1031) );
XNOR2_X1 U819 ( .A(G143), .B(n1140), .ZN(G45) );
NOR2_X1 U820 ( .A1(n1141), .A2(KEYINPUT4), .ZN(n1140) );
INV_X1 U821 ( .A(n1115), .ZN(n1141) );
NAND4_X1 U822 ( .A1(n1142), .A2(n991), .A3(n1143), .A4(n1015), .ZN(n1115) );
XNOR2_X1 U823 ( .A(G140), .B(n1121), .ZN(G42) );
NAND4_X1 U824 ( .A1(n1124), .A2(n1144), .A3(n997), .A4(n979), .ZN(n1121) );
INV_X1 U825 ( .A(n1145), .ZN(n1124) );
XNOR2_X1 U826 ( .A(G137), .B(n1120), .ZN(G39) );
NAND3_X1 U827 ( .A1(n1139), .A2(n1146), .A3(n1144), .ZN(n1120) );
XNOR2_X1 U828 ( .A(G134), .B(n1119), .ZN(G36) );
NAND3_X1 U829 ( .A1(n1144), .A2(n996), .A3(n1142), .ZN(n1119) );
XNOR2_X1 U830 ( .A(n1042), .B(n1147), .ZN(G33) );
NOR2_X1 U831 ( .A1(n1148), .A2(n995), .ZN(n1147) );
INV_X1 U832 ( .A(n1144), .ZN(n995) );
NOR2_X1 U833 ( .A1(n992), .A2(n1009), .ZN(n1144) );
XOR2_X1 U834 ( .A(n1122), .B(KEYINPUT12), .Z(n1148) );
NAND2_X1 U835 ( .A1(n1142), .A2(n997), .ZN(n1122) );
AND3_X1 U836 ( .A1(n1000), .A2(n1149), .A3(n1003), .ZN(n1142) );
INV_X1 U837 ( .A(G131), .ZN(n1042) );
XNOR2_X1 U838 ( .A(G128), .B(n1118), .ZN(G30) );
NAND3_X1 U839 ( .A1(n996), .A2(n991), .A3(n1139), .ZN(n1118) );
AND4_X1 U840 ( .A1(n1150), .A2(n1003), .A3(n1151), .A4(n1149), .ZN(n1139) );
XNOR2_X1 U841 ( .A(n1131), .B(n1152), .ZN(G3) );
XNOR2_X1 U842 ( .A(G101), .B(KEYINPUT16), .ZN(n1152) );
AND3_X1 U843 ( .A1(n1136), .A2(n1000), .A3(n1146), .ZN(n1131) );
XOR2_X1 U844 ( .A(n1153), .B(n1154), .Z(G27) );
NOR2_X1 U845 ( .A1(KEYINPUT39), .A2(n1155), .ZN(n1154) );
NOR4_X1 U846 ( .A1(n1156), .A2(n979), .A3(n1081), .A4(n1145), .ZN(n1153) );
NAND3_X1 U847 ( .A1(n1149), .A2(n1004), .A3(n999), .ZN(n1145) );
NAND2_X1 U848 ( .A1(n976), .A2(n1157), .ZN(n1149) );
NAND4_X1 U849 ( .A1(G902), .A2(G953), .A3(n1158), .A4(n1036), .ZN(n1157) );
INV_X1 U850 ( .A(G900), .ZN(n1036) );
INV_X1 U851 ( .A(n997), .ZN(n1081) );
XOR2_X1 U852 ( .A(G122), .B(n1134), .Z(G24) );
AND4_X1 U853 ( .A1(n1159), .A2(n1137), .A3(n1143), .A4(n1015), .ZN(n1134) );
XNOR2_X1 U854 ( .A(n1133), .B(n1160), .ZN(G21) );
NAND2_X1 U855 ( .A1(KEYINPUT2), .A2(G119), .ZN(n1160) );
AND4_X1 U856 ( .A1(n1150), .A2(n1159), .A3(n1146), .A4(n1151), .ZN(n1133) );
XOR2_X1 U857 ( .A(n1161), .B(n1130), .Z(G18) );
AND3_X1 U858 ( .A1(n996), .A2(n1000), .A3(n1159), .ZN(n1130) );
NOR2_X1 U859 ( .A1(n1143), .A2(n1162), .ZN(n996) );
INV_X1 U860 ( .A(n1015), .ZN(n1162) );
XNOR2_X1 U861 ( .A(G116), .B(KEYINPUT51), .ZN(n1161) );
XOR2_X1 U862 ( .A(n1163), .B(n1129), .Z(G15) );
AND3_X1 U863 ( .A1(n997), .A2(n1000), .A3(n1159), .ZN(n1129) );
AND4_X1 U864 ( .A1(n1125), .A2(n991), .A3(n1004), .A4(n1164), .ZN(n1159) );
NAND2_X1 U865 ( .A1(n1165), .A2(n1166), .ZN(n1000) );
OR3_X1 U866 ( .A1(n1151), .A2(n1167), .A3(KEYINPUT37), .ZN(n1166) );
NAND2_X1 U867 ( .A1(KEYINPUT37), .A2(n1137), .ZN(n1165) );
NOR2_X1 U868 ( .A1(n1015), .A2(n1018), .ZN(n997) );
INV_X1 U869 ( .A(n1143), .ZN(n1018) );
NAND2_X1 U870 ( .A1(KEYINPUT20), .A2(n1168), .ZN(n1163) );
XNOR2_X1 U871 ( .A(G110), .B(n1169), .ZN(G12) );
NOR2_X1 U872 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NOR3_X1 U873 ( .A1(n1172), .A2(n1173), .A3(n1156), .ZN(n1171) );
NOR3_X1 U874 ( .A1(n989), .A2(n1174), .A3(n1080), .ZN(n1173) );
INV_X1 U875 ( .A(n999), .ZN(n1174) );
INV_X1 U876 ( .A(n1146), .ZN(n989) );
INV_X1 U877 ( .A(KEYINPUT27), .ZN(n1172) );
NOR2_X1 U878 ( .A1(KEYINPUT27), .A2(n1132), .ZN(n1170) );
NAND3_X1 U879 ( .A1(n1136), .A2(n999), .A3(n1146), .ZN(n1132) );
NOR2_X1 U880 ( .A1(n1015), .A2(n1143), .ZN(n1146) );
XOR2_X1 U881 ( .A(n1175), .B(n1076), .Z(n1143) );
INV_X1 U882 ( .A(G475), .ZN(n1076) );
NAND2_X1 U883 ( .A1(n1074), .A2(n1176), .ZN(n1175) );
XNOR2_X1 U884 ( .A(n1177), .B(n1178), .ZN(n1074) );
XNOR2_X1 U885 ( .A(n1179), .B(n1180), .ZN(n1178) );
NOR2_X1 U886 ( .A1(G104), .A2(KEYINPUT9), .ZN(n1180) );
NAND2_X1 U887 ( .A1(KEYINPUT32), .A2(n1181), .ZN(n1179) );
XOR2_X1 U888 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U889 ( .A(n1037), .B(n1184), .Z(n1183) );
NOR2_X1 U890 ( .A1(KEYINPUT33), .A2(n1185), .ZN(n1184) );
XOR2_X1 U891 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U892 ( .A1(KEYINPUT57), .A2(G143), .ZN(n1187) );
NAND2_X1 U893 ( .A1(G214), .A2(n1188), .ZN(n1186) );
XNOR2_X1 U894 ( .A(G125), .B(G140), .ZN(n1037) );
XNOR2_X1 U895 ( .A(G131), .B(n1189), .ZN(n1182) );
XOR2_X1 U896 ( .A(KEYINPUT21), .B(G146), .Z(n1189) );
XNOR2_X1 U897 ( .A(G113), .B(G122), .ZN(n1177) );
XOR2_X1 U898 ( .A(n1190), .B(n1072), .Z(n1015) );
INV_X1 U899 ( .A(G478), .ZN(n1072) );
NAND2_X1 U900 ( .A1(n1071), .A2(n1191), .ZN(n1190) );
XNOR2_X1 U901 ( .A(KEYINPUT34), .B(n1176), .ZN(n1191) );
XOR2_X1 U902 ( .A(n1192), .B(n1193), .Z(n1071) );
XNOR2_X1 U903 ( .A(n1194), .B(n1195), .ZN(n1193) );
NOR2_X1 U904 ( .A1(KEYINPUT46), .A2(n1196), .ZN(n1195) );
XNOR2_X1 U905 ( .A(G134), .B(n1197), .ZN(n1196) );
NAND2_X1 U906 ( .A1(KEYINPUT1), .A2(n1198), .ZN(n1197) );
XOR2_X1 U907 ( .A(G143), .B(G128), .Z(n1198) );
NAND4_X1 U908 ( .A1(KEYINPUT60), .A2(G217), .A3(n1199), .A4(n1005), .ZN(n1194) );
XNOR2_X1 U909 ( .A(G107), .B(n1200), .ZN(n1192) );
NOR2_X1 U910 ( .A1(KEYINPUT35), .A2(n1201), .ZN(n1200) );
XNOR2_X1 U911 ( .A(G116), .B(G122), .ZN(n1201) );
NAND2_X1 U912 ( .A1(n1202), .A2(n1203), .ZN(n999) );
OR2_X1 U913 ( .A1(n985), .A2(KEYINPUT41), .ZN(n1203) );
INV_X1 U914 ( .A(n1137), .ZN(n985) );
NOR2_X1 U915 ( .A1(n1151), .A2(n1150), .ZN(n1137) );
INV_X1 U916 ( .A(n1167), .ZN(n1150) );
NAND3_X1 U917 ( .A1(n1167), .A2(n1151), .A3(KEYINPUT41), .ZN(n1202) );
XOR2_X1 U918 ( .A(n1011), .B(KEYINPUT25), .Z(n1151) );
XOR2_X1 U919 ( .A(n1204), .B(n1067), .Z(n1011) );
NAND2_X1 U920 ( .A1(G217), .A2(n1205), .ZN(n1067) );
NAND2_X1 U921 ( .A1(n1065), .A2(n1176), .ZN(n1204) );
XNOR2_X1 U922 ( .A(n1206), .B(n1207), .ZN(n1065) );
XNOR2_X1 U923 ( .A(n1208), .B(n1209), .ZN(n1207) );
XOR2_X1 U924 ( .A(G140), .B(G137), .Z(n1209) );
XOR2_X1 U925 ( .A(n1210), .B(n1211), .Z(n1206) );
XOR2_X1 U926 ( .A(n1212), .B(n1213), .Z(n1210) );
NAND3_X1 U927 ( .A1(n1199), .A2(n1214), .A3(G221), .ZN(n1212) );
XNOR2_X1 U928 ( .A(KEYINPUT36), .B(n1005), .ZN(n1214) );
XOR2_X1 U929 ( .A(G234), .B(KEYINPUT26), .Z(n1199) );
XOR2_X1 U930 ( .A(n1215), .B(n1014), .Z(n1167) );
NAND3_X1 U931 ( .A1(n1216), .A2(n1217), .A3(n1176), .ZN(n1014) );
NAND3_X1 U932 ( .A1(n1090), .A2(n1218), .A3(n1219), .ZN(n1217) );
INV_X1 U933 ( .A(KEYINPUT28), .ZN(n1219) );
NAND2_X1 U934 ( .A1(n1220), .A2(KEYINPUT28), .ZN(n1216) );
XNOR2_X1 U935 ( .A(n1218), .B(n1221), .ZN(n1220) );
INV_X1 U936 ( .A(n1090), .ZN(n1221) );
XNOR2_X1 U937 ( .A(n1222), .B(n1108), .ZN(n1090) );
NAND2_X1 U938 ( .A1(G210), .A2(n1188), .ZN(n1222) );
NOR2_X1 U939 ( .A1(G953), .A2(G237), .ZN(n1188) );
XOR2_X1 U940 ( .A(n1091), .B(n1223), .Z(n1218) );
NOR2_X1 U941 ( .A1(KEYINPUT50), .A2(n1224), .ZN(n1223) );
XOR2_X1 U942 ( .A(n1225), .B(n1087), .Z(n1224) );
NAND2_X1 U943 ( .A1(KEYINPUT15), .A2(n1085), .ZN(n1225) );
XNOR2_X1 U944 ( .A(n1226), .B(n1227), .ZN(n1091) );
XNOR2_X1 U945 ( .A(KEYINPUT49), .B(n1208), .ZN(n1227) );
XNOR2_X1 U946 ( .A(G113), .B(G116), .ZN(n1226) );
NAND2_X1 U947 ( .A1(KEYINPUT52), .A2(n1013), .ZN(n1215) );
XNOR2_X1 U948 ( .A(n1089), .B(KEYINPUT29), .ZN(n1013) );
INV_X1 U949 ( .A(G472), .ZN(n1089) );
NOR2_X1 U950 ( .A1(n1156), .A2(n1080), .ZN(n1136) );
NAND2_X1 U951 ( .A1(n1003), .A2(n1164), .ZN(n1080) );
NAND2_X1 U952 ( .A1(n976), .A2(n1228), .ZN(n1164) );
NAND4_X1 U953 ( .A1(G902), .A2(G953), .A3(n1158), .A4(n1062), .ZN(n1228) );
INV_X1 U954 ( .A(G898), .ZN(n1062) );
NAND3_X1 U955 ( .A1(n1158), .A2(n1005), .A3(G952), .ZN(n976) );
NAND2_X1 U956 ( .A1(G237), .A2(G234), .ZN(n1158) );
NOR2_X1 U957 ( .A1(n1125), .A2(n980), .ZN(n1003) );
INV_X1 U958 ( .A(n1004), .ZN(n980) );
NAND2_X1 U959 ( .A1(G221), .A2(n1205), .ZN(n1004) );
NAND2_X1 U960 ( .A1(G234), .A2(n1176), .ZN(n1205) );
INV_X1 U961 ( .A(n979), .ZN(n1125) );
XOR2_X1 U962 ( .A(n1229), .B(n1095), .Z(n979) );
INV_X1 U963 ( .A(G469), .ZN(n1095) );
NAND2_X1 U964 ( .A1(n1230), .A2(n1176), .ZN(n1229) );
XOR2_X1 U965 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U966 ( .A(n1047), .B(n1102), .Z(n1232) );
XOR2_X1 U967 ( .A(n1233), .B(n1234), .Z(n1102) );
XOR2_X1 U968 ( .A(G140), .B(G110), .Z(n1234) );
NAND2_X1 U969 ( .A1(G227), .A2(n1005), .ZN(n1233) );
INV_X1 U970 ( .A(G953), .ZN(n1005) );
XNOR2_X1 U971 ( .A(G143), .B(n1213), .ZN(n1047) );
XOR2_X1 U972 ( .A(G128), .B(G146), .Z(n1213) );
XNOR2_X1 U973 ( .A(n1235), .B(n1236), .ZN(n1231) );
NOR2_X1 U974 ( .A1(KEYINPUT54), .A2(n1087), .ZN(n1236) );
XNOR2_X1 U975 ( .A(G131), .B(n1048), .ZN(n1087) );
XNOR2_X1 U976 ( .A(n1237), .B(G137), .ZN(n1048) );
INV_X1 U977 ( .A(G134), .ZN(n1237) );
NOR2_X1 U978 ( .A1(KEYINPUT3), .A2(n1238), .ZN(n1235) );
XNOR2_X1 U979 ( .A(n1107), .B(n1108), .ZN(n1238) );
INV_X1 U980 ( .A(n991), .ZN(n1156) );
NOR2_X1 U981 ( .A1(n1239), .A2(n1009), .ZN(n991) );
INV_X1 U982 ( .A(n993), .ZN(n1009) );
NAND2_X1 U983 ( .A1(G214), .A2(n1240), .ZN(n993) );
XOR2_X1 U984 ( .A(KEYINPUT44), .B(n1241), .Z(n1240) );
INV_X1 U985 ( .A(n992), .ZN(n1239) );
XOR2_X1 U986 ( .A(n1242), .B(n1020), .Z(n992) );
NAND2_X1 U987 ( .A1(n1243), .A2(n1176), .ZN(n1020) );
INV_X1 U988 ( .A(G902), .ZN(n1176) );
XOR2_X1 U989 ( .A(n1244), .B(n1245), .Z(n1243) );
XOR2_X1 U990 ( .A(KEYINPUT8), .B(KEYINPUT22), .Z(n1245) );
XOR2_X1 U991 ( .A(n1110), .B(KEYINPUT17), .Z(n1244) );
XOR2_X1 U992 ( .A(n1246), .B(n1247), .Z(n1110) );
XOR2_X1 U993 ( .A(n1211), .B(n1248), .Z(n1247) );
XOR2_X1 U994 ( .A(G122), .B(n1249), .Z(n1248) );
NOR2_X1 U995 ( .A1(G953), .A2(n1061), .ZN(n1249) );
INV_X1 U996 ( .A(G224), .ZN(n1061) );
XNOR2_X1 U997 ( .A(n1155), .B(G110), .ZN(n1211) );
INV_X1 U998 ( .A(G125), .ZN(n1155) );
XNOR2_X1 U999 ( .A(n1058), .B(n1250), .ZN(n1246) );
INV_X1 U1000 ( .A(n1085), .ZN(n1250) );
XNOR2_X1 U1001 ( .A(n1251), .B(G128), .ZN(n1085) );
NAND2_X1 U1002 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND2_X1 U1003 ( .A1(G143), .A2(n1254), .ZN(n1253) );
XOR2_X1 U1004 ( .A(KEYINPUT62), .B(n1255), .Z(n1252) );
NOR2_X1 U1005 ( .A1(G143), .A2(n1254), .ZN(n1255) );
XOR2_X1 U1006 ( .A(KEYINPUT38), .B(G146), .Z(n1254) );
XNOR2_X1 U1007 ( .A(n1108), .B(n1256), .ZN(n1058) );
XOR2_X1 U1008 ( .A(n1257), .B(n1258), .Z(n1256) );
NAND2_X1 U1009 ( .A1(KEYINPUT30), .A2(n1107), .ZN(n1258) );
XNOR2_X1 U1010 ( .A(G104), .B(n968), .ZN(n1107) );
INV_X1 U1011 ( .A(G107), .ZN(n968) );
NAND2_X1 U1012 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
OR2_X1 U1013 ( .A1(n1261), .A2(n1168), .ZN(n1260) );
XOR2_X1 U1014 ( .A(n1262), .B(KEYINPUT14), .Z(n1259) );
NAND2_X1 U1015 ( .A1(n1261), .A2(n1168), .ZN(n1262) );
INV_X1 U1016 ( .A(G113), .ZN(n1168) );
XOR2_X1 U1017 ( .A(n1263), .B(n1264), .Z(n1261) );
INV_X1 U1018 ( .A(G116), .ZN(n1264) );
NAND2_X1 U1019 ( .A1(KEYINPUT23), .A2(n1208), .ZN(n1263) );
INV_X1 U1020 ( .A(G119), .ZN(n1208) );
XOR2_X1 U1021 ( .A(G101), .B(KEYINPUT5), .Z(n1108) );
NAND2_X1 U1022 ( .A1(KEYINPUT48), .A2(n1265), .ZN(n1242) );
XNOR2_X1 U1023 ( .A(KEYINPUT18), .B(n1019), .ZN(n1265) );
NAND2_X1 U1024 ( .A1(G210), .A2(n1266), .ZN(n1019) );
XOR2_X1 U1025 ( .A(KEYINPUT43), .B(n1241), .Z(n1266) );
NOR2_X1 U1026 ( .A1(G237), .A2(G902), .ZN(n1241) );
endmodule


