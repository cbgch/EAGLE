//Key = 1111100101110100111011000011110000000001001110101000101010101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362;

XOR2_X1 U760 ( .A(G107), .B(n1052), .Z(G9) );
NOR2_X1 U761 ( .A1(KEYINPUT40), .A2(n1053), .ZN(n1052) );
NOR2_X1 U762 ( .A1(n1054), .A2(n1055), .ZN(G75) );
NOR4_X1 U763 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1055) );
NOR2_X1 U764 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR3_X1 U765 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1058) );
XNOR2_X1 U766 ( .A(n1065), .B(KEYINPUT21), .ZN(n1063) );
XNOR2_X1 U767 ( .A(KEYINPUT44), .B(n1061), .ZN(n1062) );
NAND4_X1 U768 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1061) );
NAND3_X1 U769 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1056) );
NAND4_X1 U770 ( .A1(n1073), .A2(n1066), .A3(n1074), .A4(n1075), .ZN(n1072) );
NAND2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND3_X1 U772 ( .A1(n1069), .A2(n1078), .A3(n1068), .ZN(n1077) );
OR2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U774 ( .A1(n1067), .A2(n1081), .ZN(n1076) );
NAND2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U776 ( .A1(n1069), .A2(n1084), .ZN(n1083) );
XNOR2_X1 U777 ( .A(n1085), .B(n1086), .ZN(n1084) );
NAND2_X1 U778 ( .A1(KEYINPUT1), .A2(n1087), .ZN(n1085) );
NAND2_X1 U779 ( .A1(n1068), .A2(n1088), .ZN(n1082) );
OR2_X1 U780 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
INV_X1 U781 ( .A(n1091), .ZN(n1066) );
NOR3_X1 U782 ( .A1(n1092), .A2(G953), .A3(G952), .ZN(n1054) );
INV_X1 U783 ( .A(n1070), .ZN(n1092) );
NAND4_X1 U784 ( .A1(n1069), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1070) );
NOR4_X1 U785 ( .A1(n1087), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1095) );
XNOR2_X1 U786 ( .A(n1099), .B(n1100), .ZN(n1098) );
NAND2_X1 U787 ( .A1(KEYINPUT16), .A2(n1101), .ZN(n1099) );
XNOR2_X1 U788 ( .A(n1065), .B(KEYINPUT48), .ZN(n1097) );
INV_X1 U789 ( .A(n1064), .ZN(n1096) );
XOR2_X1 U790 ( .A(n1102), .B(n1103), .Z(n1093) );
NOR2_X1 U791 ( .A1(KEYINPUT62), .A2(n1104), .ZN(n1103) );
XNOR2_X1 U792 ( .A(G475), .B(KEYINPUT52), .ZN(n1104) );
NAND3_X1 U793 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(G72) );
NAND2_X1 U794 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
OR3_X1 U795 ( .A1(n1108), .A2(n1110), .A3(KEYINPUT45), .ZN(n1106) );
NOR2_X1 U796 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U797 ( .A1(n1071), .A2(G227), .ZN(n1112) );
NAND2_X1 U798 ( .A1(KEYINPUT45), .A2(n1113), .ZN(n1105) );
OR2_X1 U799 ( .A1(n1109), .A2(n1108), .ZN(n1113) );
XNOR2_X1 U800 ( .A(n1114), .B(n1115), .ZN(n1108) );
NOR3_X1 U801 ( .A1(n1116), .A2(n1111), .A3(n1117), .ZN(n1115) );
NOR2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XOR2_X1 U803 ( .A(KEYINPUT59), .B(n1120), .Z(n1116) );
AND2_X1 U804 ( .A1(n1119), .A2(n1118), .ZN(n1120) );
XNOR2_X1 U805 ( .A(n1121), .B(n1122), .ZN(n1118) );
XNOR2_X1 U806 ( .A(n1123), .B(KEYINPUT18), .ZN(n1121) );
NAND3_X1 U807 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1119) );
NAND2_X1 U808 ( .A1(KEYINPUT15), .A2(G125), .ZN(n1126) );
NAND3_X1 U809 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1125) );
INV_X1 U810 ( .A(KEYINPUT15), .ZN(n1128) );
OR2_X1 U811 ( .A1(n1129), .A2(n1127), .ZN(n1124) );
NOR2_X1 U812 ( .A1(G125), .A2(KEYINPUT55), .ZN(n1127) );
NAND2_X1 U813 ( .A1(n1071), .A2(n1130), .ZN(n1114) );
NAND2_X1 U814 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XNOR2_X1 U815 ( .A(n1133), .B(KEYINPUT26), .ZN(n1131) );
NAND2_X1 U816 ( .A1(G953), .A2(n1134), .ZN(n1109) );
NAND2_X1 U817 ( .A1(G900), .A2(G227), .ZN(n1134) );
NAND2_X1 U818 ( .A1(n1135), .A2(n1136), .ZN(G69) );
NAND3_X1 U819 ( .A1(G953), .A2(n1137), .A3(n1138), .ZN(n1136) );
XOR2_X1 U820 ( .A(KEYINPUT54), .B(n1139), .Z(n1135) );
NOR2_X1 U821 ( .A1(n1140), .A2(n1138), .ZN(n1139) );
XOR2_X1 U822 ( .A(n1141), .B(n1142), .Z(n1138) );
NOR2_X1 U823 ( .A1(n1143), .A2(G953), .ZN(n1142) );
NAND2_X1 U824 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
XOR2_X1 U825 ( .A(KEYINPUT56), .B(n1146), .Z(n1145) );
NOR2_X1 U826 ( .A1(G898), .A2(n1071), .ZN(n1146) );
XOR2_X1 U827 ( .A(n1147), .B(n1148), .Z(n1144) );
NOR2_X1 U828 ( .A1(KEYINPUT57), .A2(n1149), .ZN(n1147) );
XOR2_X1 U829 ( .A(KEYINPUT28), .B(n1150), .Z(n1149) );
AND2_X1 U830 ( .A1(n1137), .A2(G953), .ZN(n1140) );
NAND2_X1 U831 ( .A1(G224), .A2(G898), .ZN(n1137) );
NOR2_X1 U832 ( .A1(n1151), .A2(n1152), .ZN(G66) );
XNOR2_X1 U833 ( .A(n1153), .B(n1154), .ZN(n1152) );
NOR2_X1 U834 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR3_X1 U835 ( .A1(n1151), .A2(n1157), .A3(n1158), .ZN(G63) );
NOR2_X1 U836 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U837 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR3_X1 U838 ( .A1(n1163), .A2(KEYINPUT47), .A3(KEYINPUT30), .ZN(n1162) );
AND2_X1 U839 ( .A1(n1163), .A2(KEYINPUT30), .ZN(n1161) );
NOR2_X1 U840 ( .A1(n1164), .A2(n1165), .ZN(n1157) );
NOR2_X1 U841 ( .A1(KEYINPUT47), .A2(n1163), .ZN(n1164) );
NAND3_X1 U842 ( .A1(G478), .A2(G902), .A3(n1166), .ZN(n1163) );
XOR2_X1 U843 ( .A(n1057), .B(KEYINPUT32), .Z(n1166) );
NOR3_X1 U844 ( .A1(n1151), .A2(n1167), .A3(n1168), .ZN(G60) );
NOR4_X1 U845 ( .A1(n1169), .A2(n1156), .A3(KEYINPUT6), .A4(n1170), .ZN(n1168) );
INV_X1 U846 ( .A(n1171), .ZN(n1169) );
NOR2_X1 U847 ( .A1(n1171), .A2(n1172), .ZN(n1167) );
NOR3_X1 U848 ( .A1(n1156), .A2(n1173), .A3(n1170), .ZN(n1172) );
AND2_X1 U849 ( .A1(n1174), .A2(KEYINPUT6), .ZN(n1173) );
NOR2_X1 U850 ( .A1(KEYINPUT33), .A2(n1174), .ZN(n1171) );
NAND2_X1 U851 ( .A1(n1175), .A2(n1176), .ZN(G6) );
NAND2_X1 U852 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XOR2_X1 U853 ( .A(KEYINPUT9), .B(n1179), .Z(n1175) );
NOR2_X1 U854 ( .A1(n1177), .A2(n1178), .ZN(n1179) );
INV_X1 U855 ( .A(G104), .ZN(n1178) );
NOR2_X1 U856 ( .A1(n1151), .A2(n1180), .ZN(G57) );
XOR2_X1 U857 ( .A(n1181), .B(n1182), .Z(n1180) );
NAND2_X1 U858 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
OR2_X1 U859 ( .A1(n1185), .A2(KEYINPUT0), .ZN(n1184) );
XOR2_X1 U860 ( .A(n1186), .B(n1187), .Z(n1183) );
NOR2_X1 U861 ( .A1(n1188), .A2(n1156), .ZN(n1187) );
NAND2_X1 U862 ( .A1(KEYINPUT0), .A2(n1185), .ZN(n1186) );
XNOR2_X1 U863 ( .A(n1189), .B(n1190), .ZN(n1185) );
XNOR2_X1 U864 ( .A(n1123), .B(n1191), .ZN(n1189) );
NOR2_X1 U865 ( .A1(KEYINPUT12), .A2(n1192), .ZN(n1191) );
NOR2_X1 U866 ( .A1(n1151), .A2(n1193), .ZN(G54) );
XOR2_X1 U867 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U868 ( .A(n1196), .B(n1197), .Z(n1195) );
XOR2_X1 U869 ( .A(n1198), .B(KEYINPUT50), .Z(n1197) );
NAND2_X1 U870 ( .A1(n1199), .A2(KEYINPUT13), .ZN(n1196) );
XNOR2_X1 U871 ( .A(n1200), .B(n1122), .ZN(n1199) );
XOR2_X1 U872 ( .A(n1201), .B(n1202), .Z(n1194) );
NOR2_X1 U873 ( .A1(n1100), .A2(n1156), .ZN(n1202) );
NAND2_X1 U874 ( .A1(n1203), .A2(n1204), .ZN(n1201) );
NAND2_X1 U875 ( .A1(G140), .A2(n1205), .ZN(n1204) );
XNOR2_X1 U876 ( .A(n1206), .B(KEYINPUT22), .ZN(n1203) );
NOR2_X1 U877 ( .A1(n1151), .A2(n1207), .ZN(G51) );
NOR2_X1 U878 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XOR2_X1 U879 ( .A(n1210), .B(KEYINPUT27), .Z(n1209) );
NAND2_X1 U880 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XOR2_X1 U881 ( .A(n1213), .B(KEYINPUT8), .Z(n1212) );
NOR2_X1 U882 ( .A1(n1211), .A2(n1213), .ZN(n1208) );
XOR2_X1 U883 ( .A(n1214), .B(n1215), .Z(n1213) );
XOR2_X1 U884 ( .A(n1216), .B(n1217), .Z(n1214) );
NOR2_X1 U885 ( .A1(KEYINPUT25), .A2(n1218), .ZN(n1217) );
NOR2_X1 U886 ( .A1(n1219), .A2(n1156), .ZN(n1211) );
NAND2_X1 U887 ( .A1(G902), .A2(n1057), .ZN(n1156) );
NAND3_X1 U888 ( .A1(n1143), .A2(n1132), .A3(n1133), .ZN(n1057) );
AND4_X1 U889 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1133) );
NAND4_X1 U890 ( .A1(n1224), .A2(n1225), .A3(n1080), .A4(n1226), .ZN(n1220) );
XNOR2_X1 U891 ( .A(KEYINPUT61), .B(n1227), .ZN(n1226) );
AND4_X1 U892 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1132) );
NAND3_X1 U893 ( .A1(n1232), .A2(n1233), .A3(n1224), .ZN(n1228) );
XOR2_X1 U894 ( .A(KEYINPUT14), .B(n1067), .Z(n1233) );
AND4_X1 U895 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1143) );
NOR4_X1 U896 ( .A1(n1238), .A2(n1239), .A3(n1177), .A4(n1240), .ZN(n1237) );
INV_X1 U897 ( .A(n1053), .ZN(n1240) );
NAND3_X1 U898 ( .A1(n1080), .A2(n1069), .A3(n1241), .ZN(n1053) );
AND3_X1 U899 ( .A1(n1241), .A2(n1069), .A3(n1079), .ZN(n1177) );
NOR2_X1 U900 ( .A1(n1242), .A2(n1243), .ZN(n1236) );
INV_X1 U901 ( .A(n1244), .ZN(n1243) );
XOR2_X1 U902 ( .A(G210), .B(KEYINPUT20), .Z(n1219) );
NOR2_X1 U903 ( .A1(n1071), .A2(G952), .ZN(n1151) );
XNOR2_X1 U904 ( .A(G146), .B(n1230), .ZN(G48) );
NAND4_X1 U905 ( .A1(n1224), .A2(n1225), .A3(n1079), .A4(n1227), .ZN(n1230) );
XOR2_X1 U906 ( .A(n1245), .B(G143), .Z(G45) );
NAND2_X1 U907 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
OR2_X1 U908 ( .A1(n1229), .A2(KEYINPUT34), .ZN(n1247) );
NAND2_X1 U909 ( .A1(n1248), .A2(n1225), .ZN(n1229) );
NAND4_X1 U910 ( .A1(n1249), .A2(n1060), .A3(n1248), .A4(KEYINPUT34), .ZN(n1246) );
AND4_X1 U911 ( .A1(n1089), .A2(n1250), .A3(n1251), .A4(n1227), .ZN(n1248) );
NAND3_X1 U912 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(G42) );
NAND2_X1 U913 ( .A1(G140), .A2(n1231), .ZN(n1254) );
NAND2_X1 U914 ( .A1(KEYINPUT53), .A2(n1255), .ZN(n1253) );
NAND2_X1 U915 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XNOR2_X1 U916 ( .A(KEYINPUT11), .B(n1129), .ZN(n1257) );
NAND2_X1 U917 ( .A1(n1258), .A2(n1259), .ZN(n1252) );
INV_X1 U918 ( .A(KEYINPUT53), .ZN(n1259) );
NAND2_X1 U919 ( .A1(n1260), .A2(n1261), .ZN(n1258) );
OR2_X1 U920 ( .A1(n1129), .A2(KEYINPUT11), .ZN(n1261) );
NAND3_X1 U921 ( .A1(n1256), .A2(n1129), .A3(KEYINPUT11), .ZN(n1260) );
INV_X1 U922 ( .A(n1231), .ZN(n1256) );
NAND3_X1 U923 ( .A1(n1079), .A2(n1090), .A3(n1232), .ZN(n1231) );
NAND2_X1 U924 ( .A1(n1262), .A2(n1263), .ZN(G39) );
NAND4_X1 U925 ( .A1(n1264), .A2(n1067), .A3(n1224), .A4(n1232), .ZN(n1263) );
INV_X1 U926 ( .A(n1265), .ZN(n1264) );
XOR2_X1 U927 ( .A(n1266), .B(KEYINPUT35), .Z(n1262) );
NAND2_X1 U928 ( .A1(n1265), .A2(n1267), .ZN(n1266) );
NAND3_X1 U929 ( .A1(n1224), .A2(n1232), .A3(n1067), .ZN(n1267) );
XOR2_X1 U930 ( .A(G137), .B(KEYINPUT49), .Z(n1265) );
XNOR2_X1 U931 ( .A(G134), .B(n1221), .ZN(G36) );
NAND3_X1 U932 ( .A1(n1232), .A2(n1080), .A3(n1089), .ZN(n1221) );
XNOR2_X1 U933 ( .A(n1222), .B(n1268), .ZN(G33) );
XNOR2_X1 U934 ( .A(KEYINPUT41), .B(n1269), .ZN(n1268) );
NAND3_X1 U935 ( .A1(n1232), .A2(n1079), .A3(n1089), .ZN(n1222) );
AND4_X1 U936 ( .A1(n1073), .A2(n1249), .A3(n1074), .A4(n1227), .ZN(n1232) );
INV_X1 U937 ( .A(n1065), .ZN(n1073) );
XNOR2_X1 U938 ( .A(G128), .B(n1270), .ZN(G30) );
NAND4_X1 U939 ( .A1(n1224), .A2(n1225), .A3(n1080), .A4(n1227), .ZN(n1270) );
AND2_X1 U940 ( .A1(n1271), .A2(n1249), .ZN(n1225) );
XOR2_X1 U941 ( .A(G101), .B(n1239), .Z(G3) );
AND3_X1 U942 ( .A1(n1089), .A2(n1241), .A3(n1067), .ZN(n1239) );
XNOR2_X1 U943 ( .A(G125), .B(n1223), .ZN(G27) );
NAND4_X1 U944 ( .A1(n1271), .A2(n1227), .A3(n1090), .A4(n1272), .ZN(n1223) );
AND2_X1 U945 ( .A1(n1068), .A2(n1079), .ZN(n1272) );
NAND2_X1 U946 ( .A1(n1091), .A2(n1273), .ZN(n1227) );
NAND3_X1 U947 ( .A1(G902), .A2(n1274), .A3(n1111), .ZN(n1273) );
NOR2_X1 U948 ( .A1(n1071), .A2(G900), .ZN(n1111) );
XNOR2_X1 U949 ( .A(n1238), .B(n1275), .ZN(G24) );
NAND2_X1 U950 ( .A1(KEYINPUT17), .A2(G122), .ZN(n1275) );
AND3_X1 U951 ( .A1(n1271), .A2(n1276), .A3(n1277), .ZN(n1238) );
AND3_X1 U952 ( .A1(n1069), .A2(n1251), .A3(n1250), .ZN(n1277) );
NOR2_X1 U953 ( .A1(n1278), .A2(n1279), .ZN(n1069) );
NAND2_X1 U954 ( .A1(n1280), .A2(n1281), .ZN(G21) );
NAND2_X1 U955 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
XOR2_X1 U956 ( .A(KEYINPUT43), .B(n1284), .Z(n1280) );
NOR2_X1 U957 ( .A1(n1283), .A2(n1282), .ZN(n1284) );
NAND2_X1 U958 ( .A1(n1285), .A2(n1286), .ZN(n1282) );
OR2_X1 U959 ( .A1(n1234), .A2(KEYINPUT31), .ZN(n1286) );
OR2_X1 U960 ( .A1(n1287), .A2(n1060), .ZN(n1234) );
NAND3_X1 U961 ( .A1(n1271), .A2(n1287), .A3(KEYINPUT31), .ZN(n1285) );
NAND3_X1 U962 ( .A1(n1276), .A2(n1224), .A3(n1067), .ZN(n1287) );
AND2_X1 U963 ( .A1(n1279), .A2(n1278), .ZN(n1224) );
XNOR2_X1 U964 ( .A(G116), .B(n1235), .ZN(G18) );
NAND4_X1 U965 ( .A1(n1276), .A2(n1089), .A3(n1271), .A4(n1080), .ZN(n1235) );
NOR2_X1 U966 ( .A1(n1250), .A2(n1094), .ZN(n1080) );
INV_X1 U967 ( .A(n1060), .ZN(n1271) );
XOR2_X1 U968 ( .A(n1288), .B(KEYINPUT39), .Z(n1060) );
NAND2_X1 U969 ( .A1(n1289), .A2(n1290), .ZN(G15) );
NAND2_X1 U970 ( .A1(G113), .A2(n1244), .ZN(n1290) );
XOR2_X1 U971 ( .A(KEYINPUT29), .B(n1291), .Z(n1289) );
NOR2_X1 U972 ( .A1(G113), .A2(n1244), .ZN(n1291) );
NAND4_X1 U973 ( .A1(n1276), .A2(n1089), .A3(n1079), .A4(n1288), .ZN(n1244) );
AND2_X1 U974 ( .A1(n1094), .A2(n1250), .ZN(n1079) );
INV_X1 U975 ( .A(n1251), .ZN(n1094) );
NOR2_X1 U976 ( .A1(n1279), .A2(n1292), .ZN(n1089) );
AND2_X1 U977 ( .A1(n1068), .A2(n1293), .ZN(n1276) );
NOR2_X1 U978 ( .A1(n1086), .A2(n1087), .ZN(n1068) );
XNOR2_X1 U979 ( .A(n1205), .B(n1242), .ZN(G12) );
AND3_X1 U980 ( .A1(n1090), .A2(n1241), .A3(n1067), .ZN(n1242) );
NOR2_X1 U981 ( .A1(n1251), .A2(n1250), .ZN(n1067) );
XNOR2_X1 U982 ( .A(n1102), .B(n1170), .ZN(n1250) );
INV_X1 U983 ( .A(G475), .ZN(n1170) );
NOR2_X1 U984 ( .A1(n1174), .A2(G902), .ZN(n1102) );
XOR2_X1 U985 ( .A(n1294), .B(n1295), .Z(n1174) );
XOR2_X1 U986 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U987 ( .A(G122), .B(G113), .Z(n1297) );
XNOR2_X1 U988 ( .A(n1298), .B(G143), .ZN(n1296) );
XOR2_X1 U989 ( .A(n1299), .B(n1300), .Z(n1294) );
XNOR2_X1 U990 ( .A(G104), .B(n1301), .ZN(n1300) );
NAND2_X1 U991 ( .A1(KEYINPUT3), .A2(n1269), .ZN(n1301) );
INV_X1 U992 ( .A(G131), .ZN(n1269) );
XOR2_X1 U993 ( .A(n1302), .B(n1303), .Z(n1299) );
NOR2_X1 U994 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
XOR2_X1 U995 ( .A(KEYINPUT42), .B(G214), .Z(n1305) );
INV_X1 U996 ( .A(n1306), .ZN(n1304) );
NAND2_X1 U997 ( .A1(KEYINPUT58), .A2(n1307), .ZN(n1302) );
XNOR2_X1 U998 ( .A(n1308), .B(G478), .ZN(n1251) );
NAND2_X1 U999 ( .A1(n1165), .A2(n1309), .ZN(n1308) );
INV_X1 U1000 ( .A(n1159), .ZN(n1165) );
XNOR2_X1 U1001 ( .A(n1310), .B(n1311), .ZN(n1159) );
XOR2_X1 U1002 ( .A(G134), .B(n1312), .Z(n1311) );
NOR2_X1 U1003 ( .A1(KEYINPUT51), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1004 ( .A(G107), .B(n1314), .Z(n1313) );
XOR2_X1 U1005 ( .A(G122), .B(G116), .Z(n1314) );
XNOR2_X1 U1006 ( .A(n1315), .B(n1316), .ZN(n1310) );
AND2_X1 U1007 ( .A1(n1317), .A2(G217), .ZN(n1316) );
AND3_X1 U1008 ( .A1(n1288), .A2(n1293), .A3(n1249), .ZN(n1241) );
NOR2_X1 U1009 ( .A1(n1318), .A2(n1087), .ZN(n1249) );
AND2_X1 U1010 ( .A1(G221), .A2(n1319), .ZN(n1087) );
INV_X1 U1011 ( .A(n1086), .ZN(n1318) );
XOR2_X1 U1012 ( .A(n1101), .B(n1100), .Z(n1086) );
INV_X1 U1013 ( .A(G469), .ZN(n1100) );
NAND2_X1 U1014 ( .A1(n1320), .A2(n1309), .ZN(n1101) );
XOR2_X1 U1015 ( .A(n1321), .B(n1322), .Z(n1320) );
XNOR2_X1 U1016 ( .A(n1323), .B(n1198), .ZN(n1322) );
NAND2_X1 U1017 ( .A1(G227), .A2(n1071), .ZN(n1198) );
NOR2_X1 U1018 ( .A1(KEYINPUT37), .A2(n1122), .ZN(n1323) );
XOR2_X1 U1019 ( .A(n1298), .B(n1315), .Z(n1122) );
XOR2_X1 U1020 ( .A(n1200), .B(n1324), .Z(n1321) );
NOR2_X1 U1021 ( .A1(n1325), .A2(n1206), .ZN(n1324) );
NOR2_X1 U1022 ( .A1(n1205), .A2(G140), .ZN(n1206) );
NOR2_X1 U1023 ( .A1(n1129), .A2(n1326), .ZN(n1325) );
XNOR2_X1 U1024 ( .A(KEYINPUT38), .B(n1205), .ZN(n1326) );
XOR2_X1 U1025 ( .A(n1327), .B(n1328), .Z(n1200) );
XNOR2_X1 U1026 ( .A(n1123), .B(KEYINPUT23), .ZN(n1327) );
NAND2_X1 U1027 ( .A1(n1329), .A2(n1091), .ZN(n1293) );
NAND3_X1 U1028 ( .A1(n1274), .A2(n1071), .A3(G952), .ZN(n1091) );
XOR2_X1 U1029 ( .A(n1330), .B(KEYINPUT24), .Z(n1329) );
NAND4_X1 U1030 ( .A1(n1331), .A2(G953), .A3(G902), .A4(n1274), .ZN(n1330) );
NAND2_X1 U1031 ( .A1(G237), .A2(G234), .ZN(n1274) );
XNOR2_X1 U1032 ( .A(G898), .B(KEYINPUT5), .ZN(n1331) );
AND2_X1 U1033 ( .A1(n1065), .A2(n1074), .ZN(n1288) );
XNOR2_X1 U1034 ( .A(n1064), .B(KEYINPUT60), .ZN(n1074) );
NAND2_X1 U1035 ( .A1(G214), .A2(n1332), .ZN(n1064) );
XNOR2_X1 U1036 ( .A(n1333), .B(n1334), .ZN(n1065) );
AND2_X1 U1037 ( .A1(n1332), .A2(G210), .ZN(n1334) );
NAND2_X1 U1038 ( .A1(n1335), .A2(n1309), .ZN(n1332) );
XNOR2_X1 U1039 ( .A(G237), .B(KEYINPUT36), .ZN(n1335) );
NAND2_X1 U1040 ( .A1(n1336), .A2(n1309), .ZN(n1333) );
XNOR2_X1 U1041 ( .A(n1215), .B(n1337), .ZN(n1336) );
XNOR2_X1 U1042 ( .A(n1216), .B(n1218), .ZN(n1337) );
XNOR2_X1 U1043 ( .A(n1192), .B(n1338), .ZN(n1216) );
AND2_X1 U1044 ( .A1(n1071), .A2(G224), .ZN(n1338) );
XOR2_X1 U1045 ( .A(n1150), .B(n1148), .Z(n1215) );
XNOR2_X1 U1046 ( .A(G122), .B(n1205), .ZN(n1148) );
XNOR2_X1 U1047 ( .A(n1339), .B(n1328), .ZN(n1150) );
XNOR2_X1 U1048 ( .A(n1340), .B(n1341), .ZN(n1328) );
XOR2_X1 U1049 ( .A(KEYINPUT19), .B(G107), .Z(n1341) );
XNOR2_X1 U1050 ( .A(G101), .B(G104), .ZN(n1340) );
XOR2_X1 U1051 ( .A(n1342), .B(KEYINPUT7), .Z(n1339) );
AND2_X1 U1052 ( .A1(n1292), .A2(n1279), .ZN(n1090) );
XOR2_X1 U1053 ( .A(n1343), .B(n1155), .Z(n1279) );
NAND2_X1 U1054 ( .A1(G217), .A2(n1319), .ZN(n1155) );
NAND2_X1 U1055 ( .A1(G234), .A2(n1309), .ZN(n1319) );
NAND2_X1 U1056 ( .A1(n1344), .A2(n1153), .ZN(n1343) );
XNOR2_X1 U1057 ( .A(n1345), .B(n1346), .ZN(n1153) );
XOR2_X1 U1058 ( .A(n1347), .B(n1348), .Z(n1346) );
XNOR2_X1 U1059 ( .A(n1283), .B(G110), .ZN(n1348) );
XNOR2_X1 U1060 ( .A(n1298), .B(G137), .ZN(n1347) );
XOR2_X1 U1061 ( .A(n1349), .B(n1350), .Z(n1345) );
XNOR2_X1 U1062 ( .A(n1351), .B(n1307), .ZN(n1349) );
XNOR2_X1 U1063 ( .A(n1218), .B(n1129), .ZN(n1307) );
INV_X1 U1064 ( .A(G140), .ZN(n1129) );
INV_X1 U1065 ( .A(G125), .ZN(n1218) );
NAND2_X1 U1066 ( .A1(n1317), .A2(G221), .ZN(n1351) );
AND2_X1 U1067 ( .A1(G234), .A2(n1071), .ZN(n1317) );
INV_X1 U1068 ( .A(G953), .ZN(n1071) );
XNOR2_X1 U1069 ( .A(KEYINPUT2), .B(n1309), .ZN(n1344) );
INV_X1 U1070 ( .A(n1278), .ZN(n1292) );
XOR2_X1 U1071 ( .A(n1352), .B(n1188), .Z(n1278) );
INV_X1 U1072 ( .A(G472), .ZN(n1188) );
NAND2_X1 U1073 ( .A1(n1353), .A2(n1309), .ZN(n1352) );
INV_X1 U1074 ( .A(G902), .ZN(n1309) );
XOR2_X1 U1075 ( .A(n1354), .B(n1355), .Z(n1353) );
XNOR2_X1 U1076 ( .A(n1192), .B(n1190), .ZN(n1355) );
XNOR2_X1 U1077 ( .A(n1342), .B(KEYINPUT10), .ZN(n1190) );
XNOR2_X1 U1078 ( .A(G113), .B(n1356), .ZN(n1342) );
XNOR2_X1 U1079 ( .A(n1283), .B(G116), .ZN(n1356) );
INV_X1 U1080 ( .A(G119), .ZN(n1283) );
AND2_X1 U1081 ( .A1(n1357), .A2(n1358), .ZN(n1192) );
NAND2_X1 U1082 ( .A1(n1315), .A2(n1298), .ZN(n1358) );
INV_X1 U1083 ( .A(G146), .ZN(n1298) );
NAND2_X1 U1084 ( .A1(n1359), .A2(G146), .ZN(n1357) );
XOR2_X1 U1085 ( .A(KEYINPUT4), .B(n1315), .Z(n1359) );
XOR2_X1 U1086 ( .A(G143), .B(n1350), .Z(n1315) );
XOR2_X1 U1087 ( .A(G128), .B(KEYINPUT63), .Z(n1350) );
XOR2_X1 U1088 ( .A(n1360), .B(n1182), .Z(n1354) );
XNOR2_X1 U1089 ( .A(n1361), .B(G101), .ZN(n1182) );
NAND2_X1 U1090 ( .A1(n1306), .A2(G210), .ZN(n1361) );
NOR2_X1 U1091 ( .A1(G953), .A2(G237), .ZN(n1306) );
NAND2_X1 U1092 ( .A1(KEYINPUT46), .A2(n1123), .ZN(n1360) );
XOR2_X1 U1093 ( .A(G131), .B(n1362), .Z(n1123) );
XOR2_X1 U1094 ( .A(G137), .B(G134), .Z(n1362) );
INV_X1 U1095 ( .A(G110), .ZN(n1205) );
endmodule


