//Key = 0011111111110001101101000001001001010010100011000000111111100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377;

XNOR2_X1 U756 ( .A(G107), .B(n1044), .ZN(G9) );
NOR2_X1 U757 ( .A1(n1045), .A2(n1046), .ZN(G75) );
NOR4_X1 U758 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
NOR3_X1 U759 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1049) );
NAND3_X1 U760 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1051) );
OR2_X1 U761 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NAND3_X1 U762 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1047) );
NAND4_X1 U763 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1061) );
NOR2_X1 U764 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
INV_X1 U765 ( .A(n1053), .ZN(n1064) );
NAND2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1063) );
NAND3_X1 U767 ( .A1(n1056), .A2(n1070), .A3(n1071), .ZN(n1068) );
NAND2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NAND3_X1 U769 ( .A1(n1074), .A2(n1075), .A3(n1054), .ZN(n1062) );
NAND2_X1 U770 ( .A1(n1071), .A2(n1076), .ZN(n1075) );
OR2_X1 U771 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U772 ( .A1(n1079), .A2(n1056), .ZN(n1074) );
XNOR2_X1 U773 ( .A(n1080), .B(n1081), .ZN(n1079) );
NOR2_X1 U774 ( .A1(KEYINPUT46), .A2(n1082), .ZN(n1081) );
AND3_X1 U775 ( .A1(n1059), .A2(n1060), .A3(n1083), .ZN(n1045) );
NAND4_X1 U776 ( .A1(n1084), .A2(n1054), .A3(n1085), .A4(n1086), .ZN(n1059) );
NOR4_X1 U777 ( .A1(n1080), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1086) );
XOR2_X1 U778 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U779 ( .A1(n1092), .A2(KEYINPUT26), .ZN(n1091) );
INV_X1 U780 ( .A(n1093), .ZN(n1092) );
AND2_X1 U781 ( .A1(n1094), .A2(G472), .ZN(n1088) );
NOR2_X1 U782 ( .A1(n1067), .A2(n1095), .ZN(n1085) );
XNOR2_X1 U783 ( .A(n1096), .B(n1097), .ZN(n1084) );
NAND2_X1 U784 ( .A1(KEYINPUT21), .A2(n1098), .ZN(n1096) );
NAND2_X1 U785 ( .A1(n1099), .A2(n1100), .ZN(G72) );
NAND2_X1 U786 ( .A1(n1101), .A2(n1060), .ZN(n1100) );
NAND2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND2_X1 U788 ( .A1(n1104), .A2(n1050), .ZN(n1103) );
NAND2_X1 U789 ( .A1(n1105), .A2(n1106), .ZN(n1102) );
NAND2_X1 U790 ( .A1(n1107), .A2(G953), .ZN(n1099) );
XOR2_X1 U791 ( .A(n1108), .B(n1105), .Z(n1107) );
XOR2_X1 U792 ( .A(n1104), .B(KEYINPUT52), .Z(n1105) );
NAND2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1104) );
NAND2_X1 U794 ( .A1(G953), .A2(n1111), .ZN(n1110) );
XOR2_X1 U795 ( .A(n1112), .B(n1113), .Z(n1109) );
XNOR2_X1 U796 ( .A(n1114), .B(n1115), .ZN(n1113) );
NOR2_X1 U797 ( .A1(G140), .A2(KEYINPUT41), .ZN(n1115) );
NAND2_X1 U798 ( .A1(G900), .A2(G227), .ZN(n1108) );
NAND2_X1 U799 ( .A1(n1116), .A2(n1117), .ZN(G69) );
NAND2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND3_X1 U801 ( .A1(n1120), .A2(n1121), .A3(G953), .ZN(n1119) );
NAND3_X1 U802 ( .A1(n1122), .A2(n1121), .A3(n1123), .ZN(n1116) );
INV_X1 U803 ( .A(n1118), .ZN(n1123) );
XNOR2_X1 U804 ( .A(n1124), .B(n1125), .ZN(n1118) );
NOR2_X1 U805 ( .A1(n1126), .A2(G953), .ZN(n1125) );
NAND2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(n1124) );
XOR2_X1 U807 ( .A(n1129), .B(n1130), .Z(n1127) );
NAND3_X1 U808 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1129) );
NAND2_X1 U809 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND3_X1 U810 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
NAND2_X1 U811 ( .A1(KEYINPUT4), .A2(KEYINPUT0), .ZN(n1138) );
NAND2_X1 U812 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
INV_X1 U813 ( .A(KEYINPUT61), .ZN(n1140) );
NAND2_X1 U814 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
NAND2_X1 U815 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U816 ( .A1(KEYINPUT61), .A2(n1141), .ZN(n1136) );
NAND4_X1 U817 ( .A1(n1145), .A2(n1141), .A3(KEYINPUT4), .A4(n1143), .ZN(n1132) );
INV_X1 U818 ( .A(KEYINPUT0), .ZN(n1143) );
NAND2_X1 U819 ( .A1(KEYINPUT0), .A2(n1146), .ZN(n1131) );
NAND2_X1 U820 ( .A1(n1141), .A2(n1147), .ZN(n1146) );
NAND2_X1 U821 ( .A1(n1145), .A2(n1144), .ZN(n1147) );
INV_X1 U822 ( .A(KEYINPUT4), .ZN(n1144) );
INV_X1 U823 ( .A(KEYINPUT42), .ZN(n1121) );
NAND2_X1 U824 ( .A1(n1128), .A2(n1148), .ZN(n1122) );
NAND2_X1 U825 ( .A1(G953), .A2(n1120), .ZN(n1148) );
INV_X1 U826 ( .A(G224), .ZN(n1120) );
INV_X1 U827 ( .A(n1149), .ZN(n1128) );
NOR2_X1 U828 ( .A1(n1150), .A2(n1151), .ZN(G66) );
NOR3_X1 U829 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
NOR3_X1 U830 ( .A1(n1155), .A2(KEYINPUT25), .A3(n1156), .ZN(n1154) );
NOR3_X1 U831 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1156) );
AND2_X1 U832 ( .A1(n1155), .A2(KEYINPUT25), .ZN(n1153) );
INV_X1 U833 ( .A(n1160), .ZN(n1155) );
NOR3_X1 U834 ( .A1(n1157), .A2(n1161), .A3(n1158), .ZN(n1152) );
NOR2_X1 U835 ( .A1(n1162), .A2(KEYINPUT25), .ZN(n1161) );
NOR2_X1 U836 ( .A1(n1160), .A2(n1159), .ZN(n1162) );
INV_X1 U837 ( .A(KEYINPUT57), .ZN(n1159) );
NOR2_X1 U838 ( .A1(n1150), .A2(n1163), .ZN(G63) );
XNOR2_X1 U839 ( .A(n1164), .B(n1165), .ZN(n1163) );
AND2_X1 U840 ( .A1(G478), .A2(n1166), .ZN(n1165) );
NOR2_X1 U841 ( .A1(n1150), .A2(n1167), .ZN(G60) );
NOR3_X1 U842 ( .A1(n1098), .A2(n1168), .A3(n1169), .ZN(n1167) );
AND3_X1 U843 ( .A1(n1170), .A2(G475), .A3(n1166), .ZN(n1169) );
NOR2_X1 U844 ( .A1(n1171), .A2(n1170), .ZN(n1168) );
NOR2_X1 U845 ( .A1(n1172), .A2(n1097), .ZN(n1171) );
NOR2_X1 U846 ( .A1(n1050), .A2(n1048), .ZN(n1172) );
XNOR2_X1 U847 ( .A(G104), .B(n1173), .ZN(G6) );
NOR3_X1 U848 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(G57) );
NOR3_X1 U849 ( .A1(n1177), .A2(n1060), .A3(n1083), .ZN(n1176) );
INV_X1 U850 ( .A(G952), .ZN(n1083) );
AND2_X1 U851 ( .A1(n1177), .A2(n1150), .ZN(n1175) );
INV_X1 U852 ( .A(KEYINPUT24), .ZN(n1177) );
NOR2_X1 U853 ( .A1(n1178), .A2(n1179), .ZN(n1174) );
XOR2_X1 U854 ( .A(KEYINPUT17), .B(n1180), .Z(n1179) );
NOR2_X1 U855 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
AND2_X1 U856 ( .A1(n1182), .A2(n1181), .ZN(n1178) );
XOR2_X1 U857 ( .A(n1183), .B(n1184), .Z(n1181) );
NOR2_X1 U858 ( .A1(G101), .A2(KEYINPUT28), .ZN(n1184) );
XNOR2_X1 U859 ( .A(n1185), .B(n1186), .ZN(n1182) );
XOR2_X1 U860 ( .A(n1187), .B(n1188), .Z(n1185) );
AND2_X1 U861 ( .A1(G472), .A2(n1166), .ZN(n1188) );
NAND2_X1 U862 ( .A1(KEYINPUT19), .A2(n1189), .ZN(n1187) );
NAND2_X1 U863 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND2_X1 U864 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U865 ( .A(KEYINPUT45), .B(n1194), .Z(n1190) );
NOR2_X1 U866 ( .A1(n1193), .A2(n1192), .ZN(n1194) );
XOR2_X1 U867 ( .A(KEYINPUT32), .B(n1195), .Z(n1192) );
NOR2_X1 U868 ( .A1(n1150), .A2(n1196), .ZN(G54) );
XOR2_X1 U869 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U870 ( .A(n1199), .B(n1200), .Z(n1198) );
XOR2_X1 U871 ( .A(KEYINPUT2), .B(G140), .Z(n1200) );
XOR2_X1 U872 ( .A(KEYINPUT53), .B(KEYINPUT30), .Z(n1199) );
XOR2_X1 U873 ( .A(n1201), .B(n1202), .Z(n1197) );
XNOR2_X1 U874 ( .A(G110), .B(n1203), .ZN(n1202) );
XOR2_X1 U875 ( .A(n1204), .B(n1205), .Z(n1201) );
NAND3_X1 U876 ( .A1(n1166), .A2(G469), .A3(KEYINPUT15), .ZN(n1204) );
INV_X1 U877 ( .A(n1157), .ZN(n1166) );
NOR2_X1 U878 ( .A1(n1150), .A2(n1206), .ZN(G51) );
XOR2_X1 U879 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR2_X1 U880 ( .A1(n1093), .A2(n1157), .ZN(n1208) );
NAND2_X1 U881 ( .A1(G902), .A2(n1209), .ZN(n1157) );
NAND2_X1 U882 ( .A1(n1126), .A2(n1106), .ZN(n1209) );
INV_X1 U883 ( .A(n1050), .ZN(n1106) );
NAND4_X1 U884 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1050) );
AND4_X1 U885 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1213) );
AND2_X1 U886 ( .A1(n1218), .A2(n1219), .ZN(n1212) );
NAND2_X1 U887 ( .A1(n1071), .A2(n1220), .ZN(n1210) );
XNOR2_X1 U888 ( .A(KEYINPUT37), .B(n1221), .ZN(n1220) );
INV_X1 U889 ( .A(n1048), .ZN(n1126) );
NAND4_X1 U890 ( .A1(n1173), .A2(n1044), .A3(n1222), .A4(n1223), .ZN(n1048) );
NOR4_X1 U891 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1223) );
NOR2_X1 U892 ( .A1(n1228), .A2(n1229), .ZN(n1222) );
NOR4_X1 U893 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1229) );
XOR2_X1 U894 ( .A(KEYINPUT62), .B(n1234), .Z(n1233) );
INV_X1 U895 ( .A(n1235), .ZN(n1228) );
NAND2_X1 U896 ( .A1(n1078), .A2(n1236), .ZN(n1044) );
NAND2_X1 U897 ( .A1(n1077), .A2(n1236), .ZN(n1173) );
NOR4_X1 U898 ( .A1(n1230), .A2(n1066), .A3(n1067), .A4(n1234), .ZN(n1236) );
NOR2_X1 U899 ( .A1(n1237), .A2(n1238), .ZN(n1207) );
XOR2_X1 U900 ( .A(n1239), .B(KEYINPUT27), .Z(n1238) );
NAND2_X1 U901 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NOR2_X1 U902 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
XNOR2_X1 U903 ( .A(n1242), .B(n1243), .ZN(n1241) );
NOR2_X1 U904 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XOR2_X1 U905 ( .A(n1246), .B(KEYINPUT3), .Z(n1245) );
NAND2_X1 U906 ( .A1(n1114), .A2(n1193), .ZN(n1246) );
NOR2_X1 U907 ( .A1(n1060), .A2(G952), .ZN(n1150) );
XNOR2_X1 U908 ( .A(G146), .B(n1211), .ZN(G48) );
NAND3_X1 U909 ( .A1(n1077), .A2(n1247), .A3(n1248), .ZN(n1211) );
XOR2_X1 U910 ( .A(n1219), .B(n1249), .Z(G45) );
XNOR2_X1 U911 ( .A(G143), .B(KEYINPUT29), .ZN(n1249) );
NAND4_X1 U912 ( .A1(n1250), .A2(n1251), .A3(n1095), .A4(n1252), .ZN(n1219) );
NOR2_X1 U913 ( .A1(n1230), .A2(n1231), .ZN(n1252) );
NAND2_X1 U914 ( .A1(n1253), .A2(n1254), .ZN(G42) );
NAND2_X1 U915 ( .A1(n1255), .A2(n1218), .ZN(n1254) );
XOR2_X1 U916 ( .A(KEYINPUT54), .B(n1256), .Z(n1253) );
NOR2_X1 U917 ( .A1(n1255), .A2(n1218), .ZN(n1256) );
NAND3_X1 U918 ( .A1(n1058), .A2(n1077), .A3(n1257), .ZN(n1218) );
XNOR2_X1 U919 ( .A(KEYINPUT18), .B(G140), .ZN(n1255) );
XOR2_X1 U920 ( .A(n1258), .B(n1259), .Z(G39) );
NOR2_X1 U921 ( .A1(KEYINPUT34), .A2(n1260), .ZN(n1259) );
NOR2_X1 U922 ( .A1(n1261), .A2(n1052), .ZN(n1258) );
XOR2_X1 U923 ( .A(n1221), .B(KEYINPUT39), .Z(n1261) );
NAND4_X1 U924 ( .A1(n1248), .A2(n1056), .A3(n1073), .A4(n1262), .ZN(n1221) );
XOR2_X1 U925 ( .A(n1263), .B(n1264), .Z(G36) );
XNOR2_X1 U926 ( .A(G134), .B(KEYINPUT9), .ZN(n1264) );
NAND2_X1 U927 ( .A1(KEYINPUT6), .A2(n1217), .ZN(n1263) );
NAND3_X1 U928 ( .A1(n1057), .A2(n1078), .A3(n1257), .ZN(n1217) );
XOR2_X1 U929 ( .A(G131), .B(n1265), .Z(G33) );
NOR2_X1 U930 ( .A1(KEYINPUT49), .A2(n1216), .ZN(n1265) );
NAND3_X1 U931 ( .A1(n1057), .A2(n1077), .A3(n1257), .ZN(n1216) );
NOR4_X1 U932 ( .A1(n1052), .A2(n1266), .A3(n1267), .A4(n1072), .ZN(n1257) );
INV_X1 U933 ( .A(n1071), .ZN(n1052) );
NOR2_X1 U934 ( .A1(n1082), .A2(n1080), .ZN(n1071) );
XNOR2_X1 U935 ( .A(G128), .B(n1215), .ZN(G30) );
NAND3_X1 U936 ( .A1(n1078), .A2(n1247), .A3(n1248), .ZN(n1215) );
NOR3_X1 U937 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(n1248) );
XOR2_X1 U938 ( .A(n1270), .B(n1271), .Z(G3) );
XNOR2_X1 U939 ( .A(G101), .B(KEYINPUT50), .ZN(n1271) );
NAND2_X1 U940 ( .A1(n1272), .A2(n1057), .ZN(n1270) );
XNOR2_X1 U941 ( .A(G125), .B(n1214), .ZN(G27) );
NAND4_X1 U942 ( .A1(n1077), .A2(n1054), .A3(n1058), .A4(n1273), .ZN(n1214) );
NOR3_X1 U943 ( .A1(n1274), .A2(n1080), .A3(n1267), .ZN(n1273) );
INV_X1 U944 ( .A(n1251), .ZN(n1267) );
NAND2_X1 U945 ( .A1(n1053), .A2(n1275), .ZN(n1251) );
NAND3_X1 U946 ( .A1(G953), .A2(n1111), .A3(n1276), .ZN(n1275) );
INV_X1 U947 ( .A(G900), .ZN(n1111) );
INV_X1 U948 ( .A(n1277), .ZN(n1077) );
XOR2_X1 U949 ( .A(G122), .B(n1227), .Z(G24) );
AND4_X1 U950 ( .A1(n1095), .A2(n1250), .A3(n1269), .A4(n1278), .ZN(n1227) );
NOR2_X1 U951 ( .A1(n1066), .A2(n1279), .ZN(n1278) );
XNOR2_X1 U952 ( .A(G119), .B(n1280), .ZN(G21) );
NAND2_X1 U953 ( .A1(KEYINPUT5), .A2(n1226), .ZN(n1280) );
NOR4_X1 U954 ( .A1(n1232), .A2(n1279), .A3(n1269), .A4(n1268), .ZN(n1226) );
XOR2_X1 U955 ( .A(n1225), .B(n1281), .Z(G18) );
NOR2_X1 U956 ( .A1(KEYINPUT23), .A2(n1282), .ZN(n1281) );
INV_X1 U957 ( .A(G116), .ZN(n1282) );
AND3_X1 U958 ( .A1(n1283), .A2(n1078), .A3(n1057), .ZN(n1225) );
NOR2_X1 U959 ( .A1(n1250), .A2(n1284), .ZN(n1078) );
XOR2_X1 U960 ( .A(G113), .B(n1224), .Z(G15) );
NOR3_X1 U961 ( .A1(n1279), .A2(n1277), .A3(n1231), .ZN(n1224) );
INV_X1 U962 ( .A(n1057), .ZN(n1231) );
NOR2_X1 U963 ( .A1(n1067), .A2(n1268), .ZN(n1057) );
NAND2_X1 U964 ( .A1(n1284), .A2(n1250), .ZN(n1277) );
INV_X1 U965 ( .A(n1095), .ZN(n1284) );
INV_X1 U966 ( .A(n1283), .ZN(n1279) );
NOR4_X1 U967 ( .A1(n1069), .A2(n1274), .A3(n1234), .A4(n1080), .ZN(n1283) );
INV_X1 U968 ( .A(n1054), .ZN(n1069) );
NOR2_X1 U969 ( .A1(n1073), .A2(n1072), .ZN(n1054) );
XNOR2_X1 U970 ( .A(G110), .B(n1235), .ZN(G12) );
NAND2_X1 U971 ( .A1(n1272), .A2(n1058), .ZN(n1235) );
NOR2_X1 U972 ( .A1(n1066), .A2(n1269), .ZN(n1058) );
INV_X1 U973 ( .A(n1067), .ZN(n1269) );
XOR2_X1 U974 ( .A(n1285), .B(n1158), .Z(n1067) );
NAND2_X1 U975 ( .A1(G217), .A2(n1286), .ZN(n1158) );
NAND2_X1 U976 ( .A1(n1160), .A2(n1287), .ZN(n1285) );
XNOR2_X1 U977 ( .A(n1288), .B(n1289), .ZN(n1160) );
XOR2_X1 U978 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U979 ( .A(n1292), .B(n1293), .Z(n1291) );
NOR2_X1 U980 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
INV_X1 U981 ( .A(G221), .ZN(n1295) );
NAND2_X1 U982 ( .A1(n1296), .A2(n1297), .ZN(n1292) );
XOR2_X1 U983 ( .A(KEYINPUT11), .B(n1298), .Z(n1296) );
NAND2_X1 U984 ( .A1(KEYINPUT16), .A2(n1299), .ZN(n1290) );
XOR2_X1 U985 ( .A(n1300), .B(n1301), .Z(n1288) );
XNOR2_X1 U986 ( .A(n1302), .B(G110), .ZN(n1301) );
INV_X1 U987 ( .A(G119), .ZN(n1302) );
XNOR2_X1 U988 ( .A(G137), .B(G128), .ZN(n1300) );
INV_X1 U989 ( .A(n1268), .ZN(n1066) );
NOR2_X1 U990 ( .A1(n1303), .A2(n1087), .ZN(n1268) );
NOR2_X1 U991 ( .A1(n1094), .A2(G472), .ZN(n1087) );
AND2_X1 U992 ( .A1(n1304), .A2(G472), .ZN(n1303) );
XOR2_X1 U993 ( .A(n1094), .B(KEYINPUT22), .Z(n1304) );
NAND2_X1 U994 ( .A1(n1305), .A2(n1287), .ZN(n1094) );
XOR2_X1 U995 ( .A(n1306), .B(n1307), .Z(n1305) );
NOR2_X1 U996 ( .A1(KEYINPUT43), .A2(n1308), .ZN(n1307) );
XOR2_X1 U997 ( .A(n1309), .B(n1195), .Z(n1308) );
XOR2_X1 U998 ( .A(n1193), .B(n1186), .Z(n1309) );
XNOR2_X1 U999 ( .A(n1310), .B(G119), .ZN(n1186) );
XOR2_X1 U1000 ( .A(n1183), .B(G101), .Z(n1306) );
NAND3_X1 U1001 ( .A1(n1311), .A2(n1312), .A3(G210), .ZN(n1183) );
NOR3_X1 U1002 ( .A1(n1230), .A2(n1234), .A3(n1232), .ZN(n1272) );
INV_X1 U1003 ( .A(n1056), .ZN(n1232) );
NOR2_X1 U1004 ( .A1(n1095), .A2(n1250), .ZN(n1056) );
XOR2_X1 U1005 ( .A(n1098), .B(n1313), .Z(n1250) );
XNOR2_X1 U1006 ( .A(KEYINPUT13), .B(n1097), .ZN(n1313) );
INV_X1 U1007 ( .A(G475), .ZN(n1097) );
NOR2_X1 U1008 ( .A1(n1170), .A2(G902), .ZN(n1098) );
XOR2_X1 U1009 ( .A(n1314), .B(n1315), .Z(n1170) );
XOR2_X1 U1010 ( .A(n1316), .B(n1317), .Z(n1315) );
XNOR2_X1 U1011 ( .A(n1318), .B(n1319), .ZN(n1317) );
NOR2_X1 U1012 ( .A1(KEYINPUT63), .A2(n1320), .ZN(n1319) );
NOR2_X1 U1013 ( .A1(n1298), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1014 ( .A(n1297), .B(KEYINPUT44), .Z(n1321) );
NAND2_X1 U1015 ( .A1(G140), .A2(n1114), .ZN(n1297) );
NOR2_X1 U1016 ( .A1(G140), .A2(n1114), .ZN(n1298) );
NAND2_X1 U1017 ( .A1(KEYINPUT58), .A2(n1322), .ZN(n1318) );
XOR2_X1 U1018 ( .A(n1323), .B(n1324), .Z(n1322) );
XNOR2_X1 U1019 ( .A(G131), .B(G143), .ZN(n1324) );
NAND3_X1 U1020 ( .A1(n1311), .A2(n1312), .A3(G214), .ZN(n1323) );
XNOR2_X1 U1021 ( .A(G104), .B(n1325), .ZN(n1314) );
XNOR2_X1 U1022 ( .A(n1299), .B(G122), .ZN(n1325) );
INV_X1 U1023 ( .A(G146), .ZN(n1299) );
XNOR2_X1 U1024 ( .A(n1326), .B(G478), .ZN(n1095) );
NAND2_X1 U1025 ( .A1(n1327), .A2(n1164), .ZN(n1326) );
XNOR2_X1 U1026 ( .A(n1328), .B(n1329), .ZN(n1164) );
XOR2_X1 U1027 ( .A(n1330), .B(n1331), .Z(n1329) );
XNOR2_X1 U1028 ( .A(n1332), .B(G122), .ZN(n1331) );
XNOR2_X1 U1029 ( .A(n1333), .B(G134), .ZN(n1330) );
XOR2_X1 U1030 ( .A(n1334), .B(n1335), .Z(n1328) );
NOR2_X1 U1031 ( .A1(n1294), .A2(n1336), .ZN(n1335) );
INV_X1 U1032 ( .A(G217), .ZN(n1336) );
NAND2_X1 U1033 ( .A1(G234), .A2(n1311), .ZN(n1294) );
XNOR2_X1 U1034 ( .A(G107), .B(G116), .ZN(n1334) );
XNOR2_X1 U1035 ( .A(KEYINPUT33), .B(n1287), .ZN(n1327) );
AND2_X1 U1036 ( .A1(n1337), .A2(n1053), .ZN(n1234) );
NAND3_X1 U1037 ( .A1(n1338), .A2(n1060), .A3(G952), .ZN(n1053) );
NAND2_X1 U1038 ( .A1(n1149), .A2(n1276), .ZN(n1337) );
AND2_X1 U1039 ( .A1(n1339), .A2(n1338), .ZN(n1276) );
NAND2_X1 U1040 ( .A1(G237), .A2(G234), .ZN(n1338) );
XNOR2_X1 U1041 ( .A(KEYINPUT51), .B(n1287), .ZN(n1339) );
NOR2_X1 U1042 ( .A1(G898), .A2(n1060), .ZN(n1149) );
INV_X1 U1043 ( .A(n1247), .ZN(n1230) );
NOR4_X1 U1044 ( .A1(n1266), .A2(n1274), .A3(n1072), .A4(n1080), .ZN(n1247) );
AND2_X1 U1045 ( .A1(G214), .A2(n1340), .ZN(n1080) );
INV_X1 U1046 ( .A(n1262), .ZN(n1072) );
NAND2_X1 U1047 ( .A1(G221), .A2(n1286), .ZN(n1262) );
NAND2_X1 U1048 ( .A1(G234), .A2(n1287), .ZN(n1286) );
INV_X1 U1049 ( .A(n1082), .ZN(n1274) );
XOR2_X1 U1050 ( .A(n1090), .B(n1093), .Z(n1082) );
NAND2_X1 U1051 ( .A1(G210), .A2(n1340), .ZN(n1093) );
NAND2_X1 U1052 ( .A1(n1341), .A2(n1287), .ZN(n1340) );
XNOR2_X1 U1053 ( .A(KEYINPUT10), .B(n1312), .ZN(n1341) );
INV_X1 U1054 ( .A(G237), .ZN(n1312) );
NAND2_X1 U1055 ( .A1(n1342), .A2(n1287), .ZN(n1090) );
XOR2_X1 U1056 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1057 ( .A(n1242), .B(n1240), .Z(n1344) );
XOR2_X1 U1058 ( .A(n1345), .B(n1130), .Z(n1240) );
XNOR2_X1 U1059 ( .A(n1346), .B(G122), .ZN(n1130) );
NAND2_X1 U1060 ( .A1(KEYINPUT40), .A2(n1347), .ZN(n1345) );
XOR2_X1 U1061 ( .A(n1348), .B(n1141), .Z(n1347) );
NOR2_X1 U1062 ( .A1(KEYINPUT59), .A2(n1145), .ZN(n1348) );
INV_X1 U1063 ( .A(n1134), .ZN(n1145) );
XNOR2_X1 U1064 ( .A(n1310), .B(n1349), .ZN(n1134) );
NOR2_X1 U1065 ( .A1(G119), .A2(KEYINPUT47), .ZN(n1349) );
XNOR2_X1 U1066 ( .A(G116), .B(n1316), .ZN(n1310) );
XOR2_X1 U1067 ( .A(G113), .B(KEYINPUT36), .Z(n1316) );
NAND2_X1 U1068 ( .A1(G224), .A2(n1311), .ZN(n1242) );
XNOR2_X1 U1069 ( .A(KEYINPUT31), .B(n1350), .ZN(n1343) );
NOR2_X1 U1070 ( .A1(KEYINPUT20), .A2(n1351), .ZN(n1350) );
NOR2_X1 U1071 ( .A1(n1352), .A2(n1244), .ZN(n1351) );
NOR2_X1 U1072 ( .A1(n1193), .A2(n1114), .ZN(n1244) );
AND2_X1 U1073 ( .A1(n1114), .A2(n1193), .ZN(n1352) );
NAND3_X1 U1074 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1193) );
NAND2_X1 U1075 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
INV_X1 U1076 ( .A(KEYINPUT35), .ZN(n1357) );
NAND3_X1 U1077 ( .A1(KEYINPUT35), .A2(n1358), .A3(n1332), .ZN(n1354) );
OR2_X1 U1078 ( .A1(n1332), .A2(n1358), .ZN(n1353) );
NOR2_X1 U1079 ( .A1(KEYINPUT60), .A2(n1356), .ZN(n1358) );
XNOR2_X1 U1080 ( .A(n1359), .B(G143), .ZN(n1356) );
NAND2_X1 U1081 ( .A1(n1360), .A2(KEYINPUT7), .ZN(n1359) );
XNOR2_X1 U1082 ( .A(G146), .B(KEYINPUT1), .ZN(n1360) );
INV_X1 U1083 ( .A(G128), .ZN(n1332) );
INV_X1 U1084 ( .A(G125), .ZN(n1114) );
INV_X1 U1085 ( .A(n1073), .ZN(n1266) );
XNOR2_X1 U1086 ( .A(n1361), .B(G469), .ZN(n1073) );
NAND2_X1 U1087 ( .A1(n1362), .A2(n1287), .ZN(n1361) );
INV_X1 U1088 ( .A(G902), .ZN(n1287) );
NAND2_X1 U1089 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
NAND2_X1 U1090 ( .A1(n1365), .A2(n1205), .ZN(n1364) );
XOR2_X1 U1091 ( .A(n1366), .B(KEYINPUT12), .Z(n1365) );
XOR2_X1 U1092 ( .A(KEYINPUT8), .B(n1367), .Z(n1363) );
NOR2_X1 U1093 ( .A1(n1366), .A2(n1368), .ZN(n1367) );
XNOR2_X1 U1094 ( .A(n1205), .B(KEYINPUT56), .ZN(n1368) );
XNOR2_X1 U1095 ( .A(n1112), .B(n1141), .ZN(n1205) );
XOR2_X1 U1096 ( .A(G101), .B(n1369), .Z(n1141) );
XNOR2_X1 U1097 ( .A(n1370), .B(G104), .ZN(n1369) );
INV_X1 U1098 ( .A(G107), .ZN(n1370) );
XOR2_X1 U1099 ( .A(n1371), .B(n1372), .Z(n1112) );
XNOR2_X1 U1100 ( .A(n1333), .B(G128), .ZN(n1372) );
INV_X1 U1101 ( .A(G143), .ZN(n1333) );
XNOR2_X1 U1102 ( .A(n1195), .B(n1373), .ZN(n1371) );
NOR2_X1 U1103 ( .A1(G146), .A2(KEYINPUT14), .ZN(n1373) );
XOR2_X1 U1104 ( .A(G131), .B(n1374), .Z(n1195) );
XNOR2_X1 U1105 ( .A(n1260), .B(G134), .ZN(n1374) );
INV_X1 U1106 ( .A(G137), .ZN(n1260) );
XOR2_X1 U1107 ( .A(n1375), .B(n1376), .Z(n1366) );
XOR2_X1 U1108 ( .A(G140), .B(n1377), .Z(n1376) );
NOR2_X1 U1109 ( .A1(KEYINPUT48), .A2(n1346), .ZN(n1377) );
INV_X1 U1110 ( .A(G110), .ZN(n1346) );
NAND2_X1 U1111 ( .A1(KEYINPUT55), .A2(n1203), .ZN(n1375) );
NAND2_X1 U1112 ( .A1(G227), .A2(n1311), .ZN(n1203) );
XNOR2_X1 U1113 ( .A(n1060), .B(KEYINPUT38), .ZN(n1311) );
INV_X1 U1114 ( .A(G953), .ZN(n1060) );
endmodule


