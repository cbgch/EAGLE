//Key = 0110011011011110010111110100011101001001101010011100110011110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332;

XOR2_X1 U743 ( .A(G107), .B(n1014), .Z(G9) );
NOR2_X1 U744 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NOR2_X1 U745 ( .A1(n1017), .A2(n1018), .ZN(G75) );
NOR3_X1 U746 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NAND3_X1 U747 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1019) );
NAND2_X1 U748 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U749 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND3_X1 U750 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NAND3_X1 U751 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1030) );
NAND2_X1 U752 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U753 ( .A1(n1037), .A2(n1016), .ZN(n1036) );
INV_X1 U754 ( .A(n1038), .ZN(n1016) );
NAND4_X1 U755 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1032) );
INV_X1 U756 ( .A(KEYINPUT37), .ZN(n1042) );
NAND2_X1 U757 ( .A1(n1040), .A2(n1043), .ZN(n1027) );
NAND2_X1 U758 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND4_X1 U759 ( .A1(KEYINPUT37), .A2(n1039), .A3(n1046), .A4(n1041), .ZN(n1045) );
NOR2_X1 U760 ( .A1(n1031), .A2(n1047), .ZN(n1046) );
NAND2_X1 U761 ( .A1(n1035), .A2(n1048), .ZN(n1044) );
NAND2_X1 U762 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND3_X1 U763 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1050) );
NAND2_X1 U764 ( .A1(n1054), .A2(n1047), .ZN(n1052) );
OR3_X1 U765 ( .A1(n1055), .A2(n1056), .A3(n1054), .ZN(n1051) );
NAND2_X1 U766 ( .A1(n1029), .A2(n1057), .ZN(n1049) );
INV_X1 U767 ( .A(n1058), .ZN(n1025) );
NOR3_X1 U768 ( .A1(n1059), .A2(G953), .A3(n1060), .ZN(n1017) );
INV_X1 U769 ( .A(n1022), .ZN(n1060) );
NAND4_X1 U770 ( .A1(n1035), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1022) );
NOR4_X1 U771 ( .A1(n1064), .A2(n1054), .A3(n1065), .A4(n1066), .ZN(n1063) );
XOR2_X1 U772 ( .A(n1067), .B(n1068), .Z(n1066) );
NOR2_X1 U773 ( .A1(G475), .A2(KEYINPUT3), .ZN(n1068) );
NOR2_X1 U774 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
XOR2_X1 U775 ( .A(KEYINPUT29), .B(G478), .Z(n1070) );
INV_X1 U776 ( .A(n1071), .ZN(n1069) );
NOR2_X1 U777 ( .A1(n1072), .A2(n1073), .ZN(n1062) );
XNOR2_X1 U778 ( .A(n1074), .B(n1075), .ZN(n1073) );
XNOR2_X1 U779 ( .A(G472), .B(n1076), .ZN(n1072) );
XNOR2_X1 U780 ( .A(KEYINPUT9), .B(n1053), .ZN(n1061) );
XNOR2_X1 U781 ( .A(G952), .B(KEYINPUT22), .ZN(n1059) );
XOR2_X1 U782 ( .A(n1077), .B(n1078), .Z(G72) );
NOR3_X1 U783 ( .A1(n1023), .A2(KEYINPUT50), .A3(n1079), .ZN(n1078) );
AND2_X1 U784 ( .A1(G227), .A2(G900), .ZN(n1079) );
NAND2_X1 U785 ( .A1(n1080), .A2(n1081), .ZN(n1077) );
NAND2_X1 U786 ( .A1(n1082), .A2(n1023), .ZN(n1081) );
XOR2_X1 U787 ( .A(n1083), .B(n1084), .Z(n1082) );
NAND3_X1 U788 ( .A1(G900), .A2(n1084), .A3(G953), .ZN(n1080) );
XNOR2_X1 U789 ( .A(n1085), .B(n1086), .ZN(n1084) );
XOR2_X1 U790 ( .A(n1087), .B(n1088), .Z(n1086) );
XOR2_X1 U791 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U792 ( .A1(G131), .A2(KEYINPUT38), .ZN(n1089) );
XOR2_X1 U793 ( .A(KEYINPUT49), .B(KEYINPUT41), .Z(n1087) );
XOR2_X1 U794 ( .A(n1091), .B(n1092), .Z(n1085) );
XOR2_X1 U795 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U796 ( .A(n1095), .B(n1096), .Z(G69) );
NOR2_X1 U797 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR3_X1 U798 ( .A1(n1023), .A2(n1099), .A3(n1100), .ZN(n1098) );
NOR2_X1 U799 ( .A1(G953), .A2(n1101), .ZN(n1097) );
NOR2_X1 U800 ( .A1(n1102), .A2(n1103), .ZN(n1095) );
XOR2_X1 U801 ( .A(n1104), .B(n1105), .Z(n1103) );
XNOR2_X1 U802 ( .A(KEYINPUT46), .B(n1106), .ZN(n1105) );
NOR2_X1 U803 ( .A1(KEYINPUT61), .A2(n1107), .ZN(n1106) );
NOR2_X1 U804 ( .A1(G898), .A2(n1023), .ZN(n1102) );
NOR4_X1 U805 ( .A1(n1108), .A2(n1109), .A3(n1110), .A4(n1111), .ZN(G66) );
NOR3_X1 U806 ( .A1(n1112), .A2(n1023), .A3(n1020), .ZN(n1111) );
INV_X1 U807 ( .A(G952), .ZN(n1020) );
AND2_X1 U808 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
INV_X1 U809 ( .A(KEYINPUT32), .ZN(n1112) );
AND4_X1 U810 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1075), .ZN(n1109) );
NOR2_X1 U811 ( .A1(n1114), .A2(n1117), .ZN(n1108) );
NOR3_X1 U812 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1117) );
NOR2_X1 U813 ( .A1(n1116), .A2(n1121), .ZN(n1119) );
XNOR2_X1 U814 ( .A(n1122), .B(KEYINPUT26), .ZN(n1121) );
INV_X1 U815 ( .A(KEYINPUT54), .ZN(n1116) );
NOR2_X1 U816 ( .A1(KEYINPUT15), .A2(n1123), .ZN(n1114) );
XNOR2_X1 U817 ( .A(KEYINPUT26), .B(n1124), .ZN(n1123) );
NOR2_X1 U818 ( .A1(n1113), .A2(n1125), .ZN(G63) );
XOR2_X1 U819 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND3_X1 U820 ( .A1(G478), .A2(n1128), .A3(G902), .ZN(n1126) );
XNOR2_X1 U821 ( .A(KEYINPUT2), .B(n1021), .ZN(n1128) );
INV_X1 U822 ( .A(n1129), .ZN(n1021) );
NOR2_X1 U823 ( .A1(n1113), .A2(n1130), .ZN(G60) );
XOR2_X1 U824 ( .A(n1131), .B(n1132), .Z(n1130) );
AND2_X1 U825 ( .A1(G475), .A2(n1115), .ZN(n1132) );
NAND2_X1 U826 ( .A1(KEYINPUT53), .A2(n1133), .ZN(n1131) );
XNOR2_X1 U827 ( .A(G104), .B(n1134), .ZN(G6) );
NOR2_X1 U828 ( .A1(n1113), .A2(n1135), .ZN(G57) );
XNOR2_X1 U829 ( .A(n1136), .B(n1137), .ZN(n1135) );
XOR2_X1 U830 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U831 ( .A1(n1115), .A2(G472), .ZN(n1139) );
NAND2_X1 U832 ( .A1(n1140), .A2(KEYINPUT59), .ZN(n1138) );
XNOR2_X1 U833 ( .A(n1141), .B(G101), .ZN(n1140) );
NOR2_X1 U834 ( .A1(n1113), .A2(n1142), .ZN(G54) );
XOR2_X1 U835 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U836 ( .A1(n1115), .A2(G469), .ZN(n1144) );
NAND2_X1 U837 ( .A1(KEYINPUT14), .A2(n1145), .ZN(n1143) );
XOR2_X1 U838 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U839 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U840 ( .A(n1150), .B(n1151), .ZN(n1146) );
NOR2_X1 U841 ( .A1(KEYINPUT16), .A2(n1152), .ZN(n1151) );
NAND2_X1 U842 ( .A1(KEYINPUT20), .A2(n1153), .ZN(n1150) );
NOR3_X1 U843 ( .A1(n1113), .A2(n1154), .A3(n1155), .ZN(G51) );
NOR3_X1 U844 ( .A1(n1156), .A2(n1157), .A3(n1118), .ZN(n1155) );
NOR2_X1 U845 ( .A1(n1158), .A2(n1159), .ZN(n1154) );
XOR2_X1 U846 ( .A(n1160), .B(KEYINPUT25), .Z(n1159) );
OR2_X1 U847 ( .A1(n1118), .A2(n1157), .ZN(n1160) );
INV_X1 U848 ( .A(n1115), .ZN(n1118) );
NOR2_X1 U849 ( .A1(n1161), .A2(n1129), .ZN(n1115) );
NOR2_X1 U850 ( .A1(n1083), .A2(n1101), .ZN(n1129) );
NAND4_X1 U851 ( .A1(n1162), .A2(n1134), .A3(n1163), .A4(n1164), .ZN(n1101) );
AND4_X1 U852 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
NAND2_X1 U853 ( .A1(n1029), .A2(n1169), .ZN(n1163) );
NAND2_X1 U854 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NAND3_X1 U855 ( .A1(n1172), .A2(n1173), .A3(n1038), .ZN(n1171) );
XNOR2_X1 U856 ( .A(KEYINPUT23), .B(n1174), .ZN(n1173) );
NAND4_X1 U857 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1170) );
NAND2_X1 U858 ( .A1(KEYINPUT44), .A2(n1179), .ZN(n1178) );
NAND2_X1 U859 ( .A1(n1180), .A2(n1181), .ZN(n1177) );
INV_X1 U860 ( .A(KEYINPUT44), .ZN(n1181) );
NAND2_X1 U861 ( .A1(n1182), .A2(n1183), .ZN(n1180) );
OR2_X1 U862 ( .A1(n1037), .A2(n1015), .ZN(n1134) );
NAND3_X1 U863 ( .A1(n1029), .A2(n1174), .A3(n1172), .ZN(n1015) );
INV_X1 U864 ( .A(n1184), .ZN(n1037) );
NAND3_X1 U865 ( .A1(n1182), .A2(n1055), .A3(n1185), .ZN(n1162) );
NAND4_X1 U866 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1083) );
AND4_X1 U867 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
NOR2_X1 U868 ( .A1(n1194), .A2(n1195), .ZN(n1188) );
NAND3_X1 U869 ( .A1(n1184), .A2(n1196), .A3(n1055), .ZN(n1187) );
NAND2_X1 U870 ( .A1(n1197), .A2(n1057), .ZN(n1186) );
INV_X1 U871 ( .A(n1156), .ZN(n1158) );
XNOR2_X1 U872 ( .A(n1198), .B(n1199), .ZN(n1156) );
NAND2_X1 U873 ( .A1(KEYINPUT12), .A2(n1200), .ZN(n1198) );
NOR2_X1 U874 ( .A1(n1023), .A2(G952), .ZN(n1113) );
XNOR2_X1 U875 ( .A(n1201), .B(n1195), .ZN(G48) );
AND2_X1 U876 ( .A1(n1184), .A2(n1202), .ZN(n1195) );
XOR2_X1 U877 ( .A(n1203), .B(G143), .Z(G45) );
NAND2_X1 U878 ( .A1(KEYINPUT42), .A2(n1190), .ZN(n1203) );
NAND3_X1 U879 ( .A1(n1056), .A2(n1172), .A3(n1204), .ZN(n1190) );
AND3_X1 U880 ( .A1(n1175), .A2(n1176), .A3(n1205), .ZN(n1204) );
XNOR2_X1 U881 ( .A(G140), .B(n1206), .ZN(G42) );
NAND3_X1 U882 ( .A1(n1184), .A2(n1196), .A3(n1207), .ZN(n1206) );
XNOR2_X1 U883 ( .A(n1055), .B(KEYINPUT6), .ZN(n1207) );
XNOR2_X1 U884 ( .A(n1194), .B(n1208), .ZN(G39) );
NAND2_X1 U885 ( .A1(KEYINPUT52), .A2(G137), .ZN(n1208) );
AND2_X1 U886 ( .A1(n1209), .A2(n1196), .ZN(n1194) );
XNOR2_X1 U887 ( .A(G134), .B(n1193), .ZN(G36) );
NAND3_X1 U888 ( .A1(n1056), .A2(n1038), .A3(n1196), .ZN(n1193) );
XNOR2_X1 U889 ( .A(G131), .B(n1192), .ZN(G33) );
NAND3_X1 U890 ( .A1(n1196), .A2(n1056), .A3(n1184), .ZN(n1192) );
AND3_X1 U891 ( .A1(n1210), .A2(n1205), .A3(n1031), .ZN(n1196) );
NOR2_X1 U892 ( .A1(n1211), .A2(n1054), .ZN(n1031) );
XNOR2_X1 U893 ( .A(G128), .B(n1191), .ZN(G30) );
NAND2_X1 U894 ( .A1(n1202), .A2(n1038), .ZN(n1191) );
AND4_X1 U895 ( .A1(n1212), .A2(n1213), .A3(n1172), .A4(n1205), .ZN(n1202) );
AND2_X1 U896 ( .A1(n1057), .A2(n1210), .ZN(n1172) );
XOR2_X1 U897 ( .A(n1214), .B(n1215), .Z(G3) );
XNOR2_X1 U898 ( .A(G101), .B(KEYINPUT43), .ZN(n1215) );
NAND2_X1 U899 ( .A1(KEYINPUT11), .A2(n1216), .ZN(n1214) );
INV_X1 U900 ( .A(n1168), .ZN(n1216) );
NAND3_X1 U901 ( .A1(n1182), .A2(n1056), .A3(n1185), .ZN(n1168) );
XNOR2_X1 U902 ( .A(G125), .B(n1217), .ZN(G27) );
NAND2_X1 U903 ( .A1(n1218), .A2(n1057), .ZN(n1217) );
XNOR2_X1 U904 ( .A(n1197), .B(KEYINPUT62), .ZN(n1218) );
AND4_X1 U905 ( .A1(n1055), .A2(n1184), .A3(n1035), .A4(n1205), .ZN(n1197) );
NAND2_X1 U906 ( .A1(n1058), .A2(n1219), .ZN(n1205) );
NAND4_X1 U907 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1221), .ZN(n1219) );
INV_X1 U908 ( .A(G900), .ZN(n1221) );
XNOR2_X1 U909 ( .A(G122), .B(n1222), .ZN(G24) );
NAND3_X1 U910 ( .A1(KEYINPUT57), .A2(n1223), .A3(n1224), .ZN(n1222) );
NOR3_X1 U911 ( .A1(n1047), .A2(n1225), .A3(n1226), .ZN(n1224) );
INV_X1 U912 ( .A(n1029), .ZN(n1047) );
NOR2_X1 U913 ( .A1(n1212), .A2(n1213), .ZN(n1029) );
NAND2_X1 U914 ( .A1(n1227), .A2(n1228), .ZN(G21) );
NAND2_X1 U915 ( .A1(G119), .A2(n1167), .ZN(n1228) );
XOR2_X1 U916 ( .A(KEYINPUT39), .B(n1229), .Z(n1227) );
NOR2_X1 U917 ( .A1(G119), .A2(n1167), .ZN(n1229) );
NAND2_X1 U918 ( .A1(n1223), .A2(n1209), .ZN(n1167) );
AND3_X1 U919 ( .A1(n1212), .A2(n1213), .A3(n1040), .ZN(n1209) );
NAND3_X1 U920 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(G18) );
OR2_X1 U921 ( .A1(n1166), .A2(G116), .ZN(n1232) );
NAND2_X1 U922 ( .A1(KEYINPUT60), .A2(n1233), .ZN(n1231) );
NAND2_X1 U923 ( .A1(n1234), .A2(n1166), .ZN(n1233) );
XNOR2_X1 U924 ( .A(KEYINPUT17), .B(G116), .ZN(n1234) );
NAND2_X1 U925 ( .A1(n1235), .A2(n1236), .ZN(n1230) );
INV_X1 U926 ( .A(KEYINPUT60), .ZN(n1236) );
NAND2_X1 U927 ( .A1(n1237), .A2(n1238), .ZN(n1235) );
OR2_X1 U928 ( .A1(G116), .A2(KEYINPUT17), .ZN(n1238) );
NAND3_X1 U929 ( .A1(G116), .A2(n1166), .A3(KEYINPUT17), .ZN(n1237) );
NAND3_X1 U930 ( .A1(n1056), .A2(n1038), .A3(n1223), .ZN(n1166) );
NOR2_X1 U931 ( .A1(n1175), .A2(n1225), .ZN(n1038) );
XNOR2_X1 U932 ( .A(G113), .B(n1165), .ZN(G15) );
NAND3_X1 U933 ( .A1(n1184), .A2(n1056), .A3(n1223), .ZN(n1165) );
INV_X1 U934 ( .A(n1179), .ZN(n1223) );
NAND2_X1 U935 ( .A1(n1182), .A2(n1035), .ZN(n1179) );
INV_X1 U936 ( .A(n1183), .ZN(n1035) );
NAND2_X1 U937 ( .A1(n1041), .A2(n1239), .ZN(n1183) );
AND2_X1 U938 ( .A1(n1057), .A2(n1174), .ZN(n1182) );
NOR2_X1 U939 ( .A1(n1240), .A2(n1212), .ZN(n1056) );
INV_X1 U940 ( .A(n1241), .ZN(n1212) );
NOR2_X1 U941 ( .A1(n1176), .A2(n1226), .ZN(n1184) );
INV_X1 U942 ( .A(n1175), .ZN(n1226) );
XNOR2_X1 U943 ( .A(G110), .B(n1242), .ZN(G12) );
NAND4_X1 U944 ( .A1(n1185), .A2(n1055), .A3(n1243), .A4(n1174), .ZN(n1242) );
NAND2_X1 U945 ( .A1(n1058), .A2(n1244), .ZN(n1174) );
NAND4_X1 U946 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1100), .ZN(n1244) );
INV_X1 U947 ( .A(G898), .ZN(n1100) );
NAND3_X1 U948 ( .A1(n1220), .A2(n1023), .A3(G952), .ZN(n1058) );
NAND2_X1 U949 ( .A1(G237), .A2(G234), .ZN(n1220) );
XOR2_X1 U950 ( .A(KEYINPUT28), .B(n1057), .Z(n1243) );
NOR2_X1 U951 ( .A1(n1053), .A2(n1054), .ZN(n1057) );
AND2_X1 U952 ( .A1(G214), .A2(n1245), .ZN(n1054) );
INV_X1 U953 ( .A(n1211), .ZN(n1053) );
XNOR2_X1 U954 ( .A(n1157), .B(n1246), .ZN(n1211) );
NOR2_X1 U955 ( .A1(G902), .A2(n1247), .ZN(n1246) );
XOR2_X1 U956 ( .A(n1248), .B(KEYINPUT63), .Z(n1247) );
NAND2_X1 U957 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
OR2_X1 U958 ( .A1(n1199), .A2(n1200), .ZN(n1250) );
NAND2_X1 U959 ( .A1(n1251), .A2(n1200), .ZN(n1249) );
XOR2_X1 U960 ( .A(n1104), .B(n1107), .Z(n1200) );
XOR2_X1 U961 ( .A(n1252), .B(n1253), .Z(n1104) );
XOR2_X1 U962 ( .A(G110), .B(n1254), .Z(n1252) );
XOR2_X1 U963 ( .A(KEYINPUT7), .B(n1199), .Z(n1251) );
XNOR2_X1 U964 ( .A(n1255), .B(n1256), .ZN(n1199) );
XNOR2_X1 U965 ( .A(n1257), .B(n1258), .ZN(n1256) );
NOR2_X1 U966 ( .A1(G953), .A2(n1099), .ZN(n1258) );
INV_X1 U967 ( .A(G224), .ZN(n1099) );
NAND2_X1 U968 ( .A1(G210), .A2(n1245), .ZN(n1157) );
NAND2_X1 U969 ( .A1(n1161), .A2(n1259), .ZN(n1245) );
NOR2_X1 U970 ( .A1(n1241), .A2(n1213), .ZN(n1055) );
INV_X1 U971 ( .A(n1240), .ZN(n1213) );
NAND3_X1 U972 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1240) );
NAND2_X1 U973 ( .A1(KEYINPUT35), .A2(n1263), .ZN(n1262) );
INV_X1 U974 ( .A(n1076), .ZN(n1263) );
OR3_X1 U975 ( .A1(n1264), .A2(KEYINPUT35), .A3(G472), .ZN(n1261) );
NAND2_X1 U976 ( .A1(G472), .A2(n1264), .ZN(n1260) );
NAND2_X1 U977 ( .A1(KEYINPUT8), .A2(n1076), .ZN(n1264) );
NAND2_X1 U978 ( .A1(n1265), .A2(n1161), .ZN(n1076) );
XOR2_X1 U979 ( .A(n1266), .B(n1267), .Z(n1265) );
XNOR2_X1 U980 ( .A(G101), .B(n1268), .ZN(n1267) );
NAND2_X1 U981 ( .A1(KEYINPUT58), .A2(n1141), .ZN(n1268) );
AND3_X1 U982 ( .A1(n1259), .A2(n1023), .A3(G210), .ZN(n1141) );
NAND2_X1 U983 ( .A1(KEYINPUT47), .A2(n1136), .ZN(n1266) );
XNOR2_X1 U984 ( .A(n1269), .B(n1270), .ZN(n1136) );
XNOR2_X1 U985 ( .A(n1153), .B(n1255), .ZN(n1270) );
NAND2_X1 U986 ( .A1(n1271), .A2(n1272), .ZN(n1255) );
NAND2_X1 U987 ( .A1(n1273), .A2(n1201), .ZN(n1272) );
XNOR2_X1 U988 ( .A(n1274), .B(KEYINPUT19), .ZN(n1273) );
NAND2_X1 U989 ( .A1(n1275), .A2(G146), .ZN(n1271) );
XNOR2_X1 U990 ( .A(KEYINPUT13), .B(n1276), .ZN(n1275) );
XOR2_X1 U991 ( .A(n1277), .B(G113), .Z(n1269) );
NAND2_X1 U992 ( .A1(KEYINPUT48), .A2(n1254), .ZN(n1277) );
XNOR2_X1 U993 ( .A(G119), .B(G116), .ZN(n1254) );
XNOR2_X1 U994 ( .A(n1074), .B(n1278), .ZN(n1241) );
NOR2_X1 U995 ( .A1(n1075), .A2(KEYINPUT0), .ZN(n1278) );
INV_X1 U996 ( .A(n1120), .ZN(n1075) );
NAND2_X1 U997 ( .A1(G217), .A2(n1279), .ZN(n1120) );
NAND2_X1 U998 ( .A1(n1124), .A2(n1161), .ZN(n1074) );
INV_X1 U999 ( .A(n1122), .ZN(n1124) );
XNOR2_X1 U1000 ( .A(n1280), .B(n1281), .ZN(n1122) );
XOR2_X1 U1001 ( .A(n1282), .B(n1283), .Z(n1281) );
NAND2_X1 U1002 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
OR2_X1 U1003 ( .A1(n1286), .A2(KEYINPUT4), .ZN(n1285) );
NAND3_X1 U1004 ( .A1(n1287), .A2(n1257), .A3(KEYINPUT4), .ZN(n1284) );
XNOR2_X1 U1005 ( .A(KEYINPUT1), .B(G140), .ZN(n1287) );
NAND2_X1 U1006 ( .A1(n1288), .A2(KEYINPUT31), .ZN(n1282) );
XOR2_X1 U1007 ( .A(n1289), .B(n1093), .Z(n1288) );
NAND2_X1 U1008 ( .A1(G221), .A2(n1290), .ZN(n1289) );
XNOR2_X1 U1009 ( .A(G146), .B(n1291), .ZN(n1280) );
NOR2_X1 U1010 ( .A1(KEYINPUT24), .A2(n1292), .ZN(n1291) );
XOR2_X1 U1011 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U1012 ( .A(G119), .B(G110), .Z(n1294) );
XNOR2_X1 U1013 ( .A(G128), .B(KEYINPUT40), .ZN(n1293) );
INV_X1 U1014 ( .A(n1033), .ZN(n1185) );
NAND2_X1 U1015 ( .A1(n1040), .A2(n1210), .ZN(n1033) );
NOR2_X1 U1016 ( .A1(n1041), .A2(n1039), .ZN(n1210) );
INV_X1 U1017 ( .A(n1239), .ZN(n1039) );
NAND2_X1 U1018 ( .A1(G221), .A2(n1279), .ZN(n1239) );
NAND2_X1 U1019 ( .A1(G234), .A2(n1161), .ZN(n1279) );
XOR2_X1 U1020 ( .A(n1295), .B(G469), .Z(n1041) );
NAND3_X1 U1021 ( .A1(n1296), .A2(n1297), .A3(n1161), .ZN(n1295) );
NAND2_X1 U1022 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
INV_X1 U1023 ( .A(KEYINPUT18), .ZN(n1299) );
XOR2_X1 U1024 ( .A(n1300), .B(n1301), .Z(n1298) );
NAND3_X1 U1025 ( .A1(n1301), .A2(n1300), .A3(KEYINPUT18), .ZN(n1296) );
XOR2_X1 U1026 ( .A(n1148), .B(n1302), .Z(n1300) );
XNOR2_X1 U1027 ( .A(n1153), .B(n1107), .ZN(n1302) );
INV_X1 U1028 ( .A(n1152), .ZN(n1107) );
XOR2_X1 U1029 ( .A(G101), .B(n1303), .Z(n1152) );
XOR2_X1 U1030 ( .A(G107), .B(G104), .Z(n1303) );
XNOR2_X1 U1031 ( .A(n1304), .B(G131), .ZN(n1153) );
NAND3_X1 U1032 ( .A1(KEYINPUT21), .A2(n1305), .A3(n1306), .ZN(n1304) );
XOR2_X1 U1033 ( .A(n1307), .B(KEYINPUT10), .Z(n1306) );
NAND2_X1 U1034 ( .A1(n1090), .A2(n1093), .ZN(n1307) );
OR2_X1 U1035 ( .A1(n1093), .A2(n1090), .ZN(n1305) );
XOR2_X1 U1036 ( .A(G134), .B(KEYINPUT55), .Z(n1090) );
XOR2_X1 U1037 ( .A(G137), .B(KEYINPUT33), .Z(n1093) );
XNOR2_X1 U1038 ( .A(n1091), .B(KEYINPUT30), .ZN(n1148) );
XNOR2_X1 U1039 ( .A(G146), .B(n1274), .ZN(n1091) );
XOR2_X1 U1040 ( .A(n1149), .B(KEYINPUT56), .Z(n1301) );
XNOR2_X1 U1041 ( .A(n1308), .B(n1309), .ZN(n1149) );
XNOR2_X1 U1042 ( .A(n1310), .B(G110), .ZN(n1309) );
INV_X1 U1043 ( .A(G140), .ZN(n1310) );
NAND2_X1 U1044 ( .A1(G227), .A2(n1023), .ZN(n1308) );
NOR2_X1 U1045 ( .A1(n1176), .A2(n1175), .ZN(n1040) );
XNOR2_X1 U1046 ( .A(n1067), .B(G475), .ZN(n1175) );
NAND2_X1 U1047 ( .A1(n1133), .A2(n1161), .ZN(n1067) );
XOR2_X1 U1048 ( .A(n1311), .B(n1312), .Z(n1133) );
XOR2_X1 U1049 ( .A(n1313), .B(n1314), .Z(n1312) );
XNOR2_X1 U1050 ( .A(n1315), .B(G104), .ZN(n1314) );
INV_X1 U1051 ( .A(G131), .ZN(n1315) );
XOR2_X1 U1052 ( .A(KEYINPUT34), .B(G143), .Z(n1313) );
XOR2_X1 U1053 ( .A(n1316), .B(n1317), .Z(n1311) );
XOR2_X1 U1054 ( .A(n1318), .B(n1319), .Z(n1317) );
NOR2_X1 U1055 ( .A1(KEYINPUT51), .A2(n1201), .ZN(n1319) );
INV_X1 U1056 ( .A(G146), .ZN(n1201) );
AND3_X1 U1057 ( .A1(G214), .A2(n1023), .A3(n1259), .ZN(n1318) );
INV_X1 U1058 ( .A(G237), .ZN(n1259) );
XOR2_X1 U1059 ( .A(n1286), .B(n1253), .Z(n1316) );
XNOR2_X1 U1060 ( .A(G113), .B(n1320), .ZN(n1253) );
XNOR2_X1 U1061 ( .A(KEYINPUT1), .B(n1094), .ZN(n1286) );
XNOR2_X1 U1062 ( .A(n1257), .B(G140), .ZN(n1094) );
INV_X1 U1063 ( .A(G125), .ZN(n1257) );
INV_X1 U1064 ( .A(n1225), .ZN(n1176) );
NOR2_X1 U1065 ( .A1(n1321), .A2(n1064), .ZN(n1225) );
NOR2_X1 U1066 ( .A1(n1071), .A2(G478), .ZN(n1064) );
AND2_X1 U1067 ( .A1(G478), .A2(n1071), .ZN(n1321) );
NAND2_X1 U1068 ( .A1(n1127), .A2(n1161), .ZN(n1071) );
INV_X1 U1069 ( .A(G902), .ZN(n1161) );
XOR2_X1 U1070 ( .A(n1322), .B(n1323), .Z(n1127) );
XNOR2_X1 U1071 ( .A(n1324), .B(n1325), .ZN(n1323) );
NOR2_X1 U1072 ( .A1(KEYINPUT45), .A2(n1320), .ZN(n1325) );
INV_X1 U1073 ( .A(G122), .ZN(n1320) );
NAND3_X1 U1074 ( .A1(G217), .A2(n1290), .A3(KEYINPUT5), .ZN(n1324) );
AND2_X1 U1075 ( .A1(G234), .A2(n1023), .ZN(n1290) );
INV_X1 U1076 ( .A(G953), .ZN(n1023) );
XOR2_X1 U1077 ( .A(n1326), .B(n1327), .Z(n1322) );
XOR2_X1 U1078 ( .A(G116), .B(G107), .Z(n1327) );
NAND3_X1 U1079 ( .A1(n1328), .A2(n1329), .A3(KEYINPUT36), .ZN(n1326) );
NAND2_X1 U1080 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
INV_X1 U1081 ( .A(KEYINPUT27), .ZN(n1331) );
XNOR2_X1 U1082 ( .A(n1332), .B(n1274), .ZN(n1330) );
NAND3_X1 U1083 ( .A1(n1276), .A2(n1332), .A3(KEYINPUT27), .ZN(n1328) );
INV_X1 U1084 ( .A(G134), .ZN(n1332) );
INV_X1 U1085 ( .A(n1274), .ZN(n1276) );
XOR2_X1 U1086 ( .A(G128), .B(G143), .Z(n1274) );
endmodule


