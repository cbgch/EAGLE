//Key = 1111011000100011100000101110101100010001110010010100001000000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
n1426, n1427;

XNOR2_X1 U776 ( .A(G107), .B(n1076), .ZN(G9) );
NOR2_X1 U777 ( .A1(n1077), .A2(n1078), .ZN(G75) );
NOR3_X1 U778 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
INV_X1 U779 ( .A(n1082), .ZN(n1081) );
INV_X1 U780 ( .A(G952), .ZN(n1080) );
NAND3_X1 U781 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1079) );
NAND2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U784 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
NAND2_X1 U785 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NAND2_X1 U786 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
OR2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1093) );
NAND2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U790 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND3_X1 U791 ( .A1(n1095), .A2(n1105), .A3(n1099), .ZN(n1088) );
NAND2_X1 U792 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U793 ( .A1(n1092), .A2(n1108), .ZN(n1107) );
OR2_X1 U794 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U795 ( .A1(n1090), .A2(n1111), .ZN(n1106) );
NAND2_X1 U796 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U797 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
INV_X1 U798 ( .A(n1116), .ZN(n1086) );
NOR3_X1 U799 ( .A1(n1117), .A2(G953), .A3(n1118), .ZN(n1077) );
INV_X1 U800 ( .A(n1083), .ZN(n1118) );
NAND4_X1 U801 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1083) );
NOR4_X1 U802 ( .A1(n1114), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1122) );
XOR2_X1 U803 ( .A(n1126), .B(KEYINPUT63), .Z(n1124) );
NAND2_X1 U804 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1123) );
INV_X1 U806 ( .A(n1129), .ZN(n1127) );
NOR2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1121) );
XNOR2_X1 U808 ( .A(n1132), .B(G475), .ZN(n1120) );
XNOR2_X1 U809 ( .A(n1133), .B(KEYINPUT4), .ZN(n1119) );
XNOR2_X1 U810 ( .A(G952), .B(KEYINPUT30), .ZN(n1117) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(G72) );
NOR3_X1 U812 ( .A1(n1084), .A2(KEYINPUT36), .A3(n1136), .ZN(n1135) );
AND2_X1 U813 ( .A1(G227), .A2(G900), .ZN(n1136) );
NAND2_X1 U814 ( .A1(n1137), .A2(n1138), .ZN(n1134) );
NAND3_X1 U815 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1138) );
NAND2_X1 U816 ( .A1(KEYINPUT37), .A2(n1142), .ZN(n1140) );
NAND2_X1 U817 ( .A1(G953), .A2(n1143), .ZN(n1142) );
NAND2_X1 U818 ( .A1(G900), .A2(n1144), .ZN(n1143) );
NAND2_X1 U819 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
OR2_X1 U820 ( .A1(n1144), .A2(G953), .ZN(n1145) );
NAND2_X1 U821 ( .A1(n1144), .A2(n1147), .ZN(n1137) );
NAND2_X1 U822 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND2_X1 U823 ( .A1(G900), .A2(n1150), .ZN(n1149) );
NAND2_X1 U824 ( .A1(n1141), .A2(n1151), .ZN(n1150) );
NAND2_X1 U825 ( .A1(G953), .A2(n1146), .ZN(n1151) );
NAND2_X1 U826 ( .A1(n1152), .A2(n1084), .ZN(n1148) );
NAND2_X1 U827 ( .A1(n1146), .A2(n1141), .ZN(n1152) );
INV_X1 U828 ( .A(KEYINPUT37), .ZN(n1146) );
XNOR2_X1 U829 ( .A(n1153), .B(n1154), .ZN(n1144) );
XOR2_X1 U830 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND2_X1 U831 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND2_X1 U832 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U833 ( .A(n1161), .B(KEYINPUT50), .Z(n1157) );
OR2_X1 U834 ( .A1(n1159), .A2(n1160), .ZN(n1161) );
XOR2_X1 U835 ( .A(G137), .B(n1162), .Z(n1159) );
NOR2_X1 U836 ( .A1(KEYINPUT52), .A2(n1163), .ZN(n1162) );
NAND2_X1 U837 ( .A1(n1164), .A2(n1165), .ZN(G69) );
NAND2_X1 U838 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
OR2_X1 U839 ( .A1(n1084), .A2(G224), .ZN(n1167) );
NAND3_X1 U840 ( .A1(G953), .A2(n1168), .A3(n1169), .ZN(n1164) );
INV_X1 U841 ( .A(n1166), .ZN(n1169) );
XNOR2_X1 U842 ( .A(n1170), .B(n1171), .ZN(n1166) );
NOR3_X1 U843 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1171) );
NOR2_X1 U844 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NOR2_X1 U845 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR2_X1 U846 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NOR2_X1 U847 ( .A1(n1181), .A2(n1182), .ZN(n1177) );
NOR2_X1 U848 ( .A1(n1183), .A2(n1184), .ZN(n1173) );
NOR2_X1 U849 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NOR2_X1 U850 ( .A1(n1181), .A2(n1180), .ZN(n1186) );
XNOR2_X1 U851 ( .A(n1182), .B(KEYINPUT7), .ZN(n1180) );
INV_X1 U852 ( .A(n1179), .ZN(n1181) );
NOR2_X1 U853 ( .A1(n1182), .A2(n1179), .ZN(n1185) );
NAND2_X1 U854 ( .A1(n1084), .A2(n1187), .ZN(n1170) );
NAND2_X1 U855 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
INV_X1 U856 ( .A(n1190), .ZN(n1189) );
XOR2_X1 U857 ( .A(n1191), .B(KEYINPUT61), .Z(n1188) );
NAND2_X1 U858 ( .A1(G898), .A2(G224), .ZN(n1168) );
NOR2_X1 U859 ( .A1(n1192), .A2(n1193), .ZN(G66) );
XOR2_X1 U860 ( .A(n1194), .B(n1195), .Z(n1193) );
NOR2_X1 U861 ( .A1(KEYINPUT12), .A2(n1196), .ZN(n1194) );
NOR2_X1 U862 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
XNOR2_X1 U863 ( .A(KEYINPUT2), .B(n1128), .ZN(n1198) );
NOR2_X1 U864 ( .A1(n1192), .A2(n1199), .ZN(G63) );
XOR2_X1 U865 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U866 ( .A(KEYINPUT26), .B(n1202), .Z(n1201) );
AND2_X1 U867 ( .A1(G478), .A2(n1203), .ZN(n1202) );
NOR2_X1 U868 ( .A1(n1192), .A2(n1204), .ZN(G60) );
NOR3_X1 U869 ( .A1(n1132), .A2(n1205), .A3(n1206), .ZN(n1204) );
AND3_X1 U870 ( .A1(n1207), .A2(G475), .A3(n1203), .ZN(n1206) );
NOR2_X1 U871 ( .A1(n1208), .A2(n1207), .ZN(n1205) );
NOR2_X1 U872 ( .A1(n1082), .A2(n1209), .ZN(n1208) );
XNOR2_X1 U873 ( .A(G104), .B(n1210), .ZN(G6) );
NOR2_X1 U874 ( .A1(n1192), .A2(n1211), .ZN(G57) );
XOR2_X1 U875 ( .A(n1212), .B(n1213), .Z(n1211) );
XOR2_X1 U876 ( .A(n1214), .B(n1215), .Z(n1213) );
AND2_X1 U877 ( .A1(G472), .A2(n1203), .ZN(n1215) );
NOR3_X1 U878 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1214) );
NOR2_X1 U879 ( .A1(n1219), .A2(n1183), .ZN(n1218) );
AND3_X1 U880 ( .A1(n1183), .A2(n1219), .A3(KEYINPUT10), .ZN(n1217) );
NOR2_X1 U881 ( .A1(n1220), .A2(KEYINPUT55), .ZN(n1219) );
INV_X1 U882 ( .A(n1221), .ZN(n1220) );
NOR2_X1 U883 ( .A1(KEYINPUT10), .A2(n1221), .ZN(n1216) );
NAND2_X1 U884 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NAND2_X1 U885 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
XOR2_X1 U886 ( .A(KEYINPUT28), .B(n1226), .Z(n1222) );
NOR2_X1 U887 ( .A1(n1225), .A2(n1224), .ZN(n1226) );
XNOR2_X1 U888 ( .A(G101), .B(n1227), .ZN(n1212) );
NOR3_X1 U889 ( .A1(n1228), .A2(n1192), .A3(n1229), .ZN(G54) );
NOR3_X1 U890 ( .A1(n1230), .A2(KEYINPUT38), .A3(n1231), .ZN(n1229) );
XOR2_X1 U891 ( .A(n1232), .B(n1233), .Z(n1230) );
NOR2_X1 U892 ( .A1(KEYINPUT48), .A2(n1234), .ZN(n1233) );
NOR2_X1 U893 ( .A1(n1235), .A2(n1236), .ZN(n1228) );
XOR2_X1 U894 ( .A(n1232), .B(n1237), .Z(n1236) );
NOR2_X1 U895 ( .A1(KEYINPUT48), .A2(n1238), .ZN(n1237) );
AND2_X1 U896 ( .A1(n1203), .A2(G469), .ZN(n1232) );
NOR2_X1 U897 ( .A1(KEYINPUT38), .A2(n1231), .ZN(n1235) );
XNOR2_X1 U898 ( .A(n1239), .B(n1240), .ZN(n1231) );
XNOR2_X1 U899 ( .A(KEYINPUT11), .B(n1241), .ZN(n1240) );
NAND2_X1 U900 ( .A1(n1242), .A2(n1243), .ZN(n1239) );
OR2_X1 U901 ( .A1(n1244), .A2(n1155), .ZN(n1243) );
XOR2_X1 U902 ( .A(n1245), .B(KEYINPUT58), .Z(n1242) );
NAND2_X1 U903 ( .A1(n1244), .A2(n1155), .ZN(n1245) );
XOR2_X1 U904 ( .A(n1246), .B(KEYINPUT59), .Z(n1244) );
NOR2_X1 U905 ( .A1(n1192), .A2(n1247), .ZN(G51) );
XOR2_X1 U906 ( .A(n1248), .B(n1249), .Z(n1247) );
XOR2_X1 U907 ( .A(n1250), .B(n1251), .Z(n1249) );
NOR2_X1 U908 ( .A1(n1252), .A2(n1197), .ZN(n1251) );
INV_X1 U909 ( .A(n1203), .ZN(n1197) );
NOR2_X1 U910 ( .A1(n1253), .A2(n1082), .ZN(n1203) );
NOR3_X1 U911 ( .A1(n1191), .A2(n1141), .A3(n1190), .ZN(n1082) );
NAND4_X1 U912 ( .A1(n1210), .A2(n1254), .A3(n1255), .A4(n1076), .ZN(n1190) );
NAND3_X1 U913 ( .A1(n1098), .A2(n1090), .A3(n1256), .ZN(n1076) );
NAND3_X1 U914 ( .A1(n1256), .A2(n1090), .A3(n1097), .ZN(n1210) );
NAND4_X1 U915 ( .A1(n1257), .A2(n1258), .A3(n1259), .A4(n1260), .ZN(n1141) );
NOR4_X1 U916 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1260) );
NOR2_X1 U917 ( .A1(n1265), .A2(n1266), .ZN(n1259) );
AND3_X1 U918 ( .A1(n1267), .A2(n1098), .A3(n1092), .ZN(n1266) );
INV_X1 U919 ( .A(n1268), .ZN(n1265) );
NAND2_X1 U920 ( .A1(n1269), .A2(n1270), .ZN(n1258) );
XNOR2_X1 U921 ( .A(KEYINPUT17), .B(n1271), .ZN(n1270) );
INV_X1 U922 ( .A(n1272), .ZN(n1269) );
NAND2_X1 U923 ( .A1(n1273), .A2(n1274), .ZN(n1257) );
XOR2_X1 U924 ( .A(n1275), .B(KEYINPUT5), .Z(n1273) );
NAND2_X1 U925 ( .A1(n1276), .A2(n1277), .ZN(n1191) );
NAND2_X1 U926 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NAND3_X1 U927 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1279) );
NAND3_X1 U928 ( .A1(n1110), .A2(n1283), .A3(n1097), .ZN(n1282) );
XOR2_X1 U929 ( .A(n1284), .B(n1285), .Z(n1248) );
NOR2_X1 U930 ( .A1(KEYINPUT18), .A2(n1286), .ZN(n1285) );
NOR2_X1 U931 ( .A1(n1084), .A2(G952), .ZN(n1192) );
XOR2_X1 U932 ( .A(G146), .B(n1264), .Z(G48) );
AND3_X1 U933 ( .A1(n1274), .A2(n1097), .A3(n1287), .ZN(n1264) );
XOR2_X1 U934 ( .A(G143), .B(n1288), .Z(G45) );
NOR2_X1 U935 ( .A1(n1112), .A2(n1275), .ZN(n1288) );
NAND3_X1 U936 ( .A1(n1289), .A2(n1131), .A3(n1267), .ZN(n1275) );
XNOR2_X1 U937 ( .A(G140), .B(n1268), .ZN(G42) );
NAND3_X1 U938 ( .A1(n1092), .A2(n1097), .A3(n1290), .ZN(n1268) );
NOR3_X1 U939 ( .A1(n1271), .A2(n1291), .A3(n1101), .ZN(n1290) );
NAND2_X1 U940 ( .A1(n1292), .A2(n1293), .ZN(G39) );
NAND2_X1 U941 ( .A1(n1263), .A2(n1294), .ZN(n1293) );
XOR2_X1 U942 ( .A(KEYINPUT44), .B(n1295), .Z(n1292) );
NOR2_X1 U943 ( .A1(n1263), .A2(n1294), .ZN(n1295) );
AND3_X1 U944 ( .A1(n1287), .A2(n1099), .A3(n1092), .ZN(n1263) );
XNOR2_X1 U945 ( .A(G134), .B(n1296), .ZN(G36) );
NAND4_X1 U946 ( .A1(n1092), .A2(n1110), .A3(n1297), .A4(n1098), .ZN(n1296) );
NOR2_X1 U947 ( .A1(n1291), .A2(n1298), .ZN(n1297) );
XNOR2_X1 U948 ( .A(n1299), .B(KEYINPUT13), .ZN(n1298) );
INV_X1 U949 ( .A(n1300), .ZN(n1291) );
NAND2_X1 U950 ( .A1(n1301), .A2(n1302), .ZN(G33) );
NAND2_X1 U951 ( .A1(n1303), .A2(n1262), .ZN(n1302) );
XNOR2_X1 U952 ( .A(G131), .B(KEYINPUT9), .ZN(n1303) );
NAND2_X1 U953 ( .A1(n1304), .A2(n1305), .ZN(n1301) );
XOR2_X1 U954 ( .A(KEYINPUT15), .B(n1262), .Z(n1305) );
AND3_X1 U955 ( .A1(n1092), .A2(n1097), .A3(n1267), .ZN(n1262) );
AND3_X1 U956 ( .A1(n1299), .A2(n1300), .A3(n1110), .ZN(n1267) );
NOR2_X1 U957 ( .A1(n1133), .A2(n1114), .ZN(n1092) );
XNOR2_X1 U958 ( .A(G131), .B(KEYINPUT0), .ZN(n1304) );
XNOR2_X1 U959 ( .A(n1261), .B(n1306), .ZN(G30) );
NAND2_X1 U960 ( .A1(KEYINPUT22), .A2(G128), .ZN(n1306) );
AND3_X1 U961 ( .A1(n1274), .A2(n1098), .A3(n1287), .ZN(n1261) );
AND4_X1 U962 ( .A1(n1307), .A2(n1308), .A3(n1299), .A4(n1300), .ZN(n1287) );
XNOR2_X1 U963 ( .A(G101), .B(n1254), .ZN(G3) );
NAND3_X1 U964 ( .A1(n1099), .A2(n1256), .A3(n1110), .ZN(n1254) );
XOR2_X1 U965 ( .A(n1309), .B(n1310), .Z(G27) );
XNOR2_X1 U966 ( .A(KEYINPUT53), .B(n1311), .ZN(n1310) );
NOR2_X1 U967 ( .A1(n1271), .A2(n1272), .ZN(n1309) );
NAND4_X1 U968 ( .A1(n1274), .A2(n1097), .A3(n1095), .A4(n1300), .ZN(n1272) );
NAND2_X1 U969 ( .A1(n1116), .A2(n1312), .ZN(n1300) );
NAND4_X1 U970 ( .A1(G953), .A2(G902), .A3(n1313), .A4(n1314), .ZN(n1312) );
INV_X1 U971 ( .A(G900), .ZN(n1314) );
XNOR2_X1 U972 ( .A(n1315), .B(n1316), .ZN(G24) );
NOR3_X1 U973 ( .A1(n1281), .A2(n1317), .A3(n1318), .ZN(n1316) );
XNOR2_X1 U974 ( .A(n1095), .B(KEYINPUT29), .ZN(n1318) );
INV_X1 U975 ( .A(n1130), .ZN(n1095) );
NAND4_X1 U976 ( .A1(n1274), .A2(n1289), .A3(n1090), .A4(n1131), .ZN(n1281) );
NOR2_X1 U977 ( .A1(n1307), .A2(n1308), .ZN(n1090) );
XNOR2_X1 U978 ( .A(G119), .B(n1276), .ZN(G21) );
NAND4_X1 U979 ( .A1(n1274), .A2(n1278), .A3(n1319), .A4(n1307), .ZN(n1276) );
INV_X1 U980 ( .A(n1320), .ZN(n1307) );
AND2_X1 U981 ( .A1(n1099), .A2(n1308), .ZN(n1319) );
XOR2_X1 U982 ( .A(G116), .B(n1321), .Z(G18) );
NOR3_X1 U983 ( .A1(n1280), .A2(KEYINPUT21), .A3(n1322), .ZN(n1321) );
INV_X1 U984 ( .A(n1278), .ZN(n1322) );
NAND3_X1 U985 ( .A1(n1110), .A2(n1098), .A3(n1274), .ZN(n1280) );
INV_X1 U986 ( .A(n1112), .ZN(n1274) );
XOR2_X1 U987 ( .A(n1283), .B(KEYINPUT24), .Z(n1112) );
NOR2_X1 U988 ( .A1(n1323), .A2(n1289), .ZN(n1098) );
XNOR2_X1 U989 ( .A(G113), .B(n1324), .ZN(G15) );
NAND4_X1 U990 ( .A1(n1325), .A2(n1278), .A3(n1097), .A4(n1110), .ZN(n1324) );
NOR2_X1 U991 ( .A1(n1320), .A2(n1308), .ZN(n1110) );
AND2_X1 U992 ( .A1(n1289), .A2(n1323), .ZN(n1097) );
INV_X1 U993 ( .A(n1131), .ZN(n1323) );
NOR2_X1 U994 ( .A1(n1130), .A2(n1317), .ZN(n1278) );
NAND2_X1 U995 ( .A1(n1104), .A2(n1326), .ZN(n1130) );
XNOR2_X1 U996 ( .A(n1283), .B(KEYINPUT1), .ZN(n1325) );
XNOR2_X1 U997 ( .A(G110), .B(n1255), .ZN(G12) );
NAND3_X1 U998 ( .A1(n1109), .A2(n1256), .A3(n1099), .ZN(n1255) );
NOR2_X1 U999 ( .A1(n1131), .A2(n1289), .ZN(n1099) );
XOR2_X1 U1000 ( .A(n1327), .B(n1328), .Z(n1289) );
XNOR2_X1 U1001 ( .A(KEYINPUT60), .B(n1209), .ZN(n1328) );
INV_X1 U1002 ( .A(G475), .ZN(n1209) );
NAND2_X1 U1003 ( .A1(n1329), .A2(KEYINPUT16), .ZN(n1327) );
XNOR2_X1 U1004 ( .A(n1132), .B(KEYINPUT57), .ZN(n1329) );
NOR2_X1 U1005 ( .A1(n1207), .A2(G902), .ZN(n1132) );
XOR2_X1 U1006 ( .A(n1330), .B(n1331), .Z(n1207) );
XOR2_X1 U1007 ( .A(n1332), .B(n1333), .Z(n1331) );
XOR2_X1 U1008 ( .A(n1334), .B(n1335), .Z(n1333) );
NOR2_X1 U1009 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XOR2_X1 U1010 ( .A(n1338), .B(KEYINPUT39), .Z(n1337) );
NAND2_X1 U1011 ( .A1(G146), .A2(n1339), .ZN(n1338) );
NOR2_X1 U1012 ( .A1(G146), .A2(n1339), .ZN(n1336) );
NAND2_X1 U1013 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
NAND2_X1 U1014 ( .A1(G140), .A2(n1311), .ZN(n1341) );
XOR2_X1 U1015 ( .A(n1342), .B(KEYINPUT8), .Z(n1340) );
NAND2_X1 U1016 ( .A1(G125), .A2(n1343), .ZN(n1342) );
NAND2_X1 U1017 ( .A1(n1344), .A2(G214), .ZN(n1334) );
XNOR2_X1 U1018 ( .A(G104), .B(G113), .ZN(n1332) );
XOR2_X1 U1019 ( .A(n1345), .B(n1346), .Z(n1330) );
XOR2_X1 U1020 ( .A(KEYINPUT23), .B(G143), .Z(n1346) );
XNOR2_X1 U1021 ( .A(G122), .B(G131), .ZN(n1345) );
XNOR2_X1 U1022 ( .A(n1347), .B(G478), .ZN(n1131) );
NAND2_X1 U1023 ( .A1(n1200), .A2(n1253), .ZN(n1347) );
XOR2_X1 U1024 ( .A(n1348), .B(n1349), .Z(n1200) );
XOR2_X1 U1025 ( .A(G128), .B(n1350), .Z(n1349) );
XNOR2_X1 U1026 ( .A(G143), .B(n1163), .ZN(n1350) );
INV_X1 U1027 ( .A(G134), .ZN(n1163) );
XOR2_X1 U1028 ( .A(n1351), .B(n1352), .Z(n1348) );
NOR2_X1 U1029 ( .A1(KEYINPUT43), .A2(n1353), .ZN(n1352) );
NOR2_X1 U1030 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
XOR2_X1 U1031 ( .A(n1356), .B(KEYINPUT62), .Z(n1355) );
NAND2_X1 U1032 ( .A1(n1357), .A2(G107), .ZN(n1356) );
NOR2_X1 U1033 ( .A1(G107), .A2(n1357), .ZN(n1354) );
XNOR2_X1 U1034 ( .A(G116), .B(n1358), .ZN(n1357) );
XNOR2_X1 U1035 ( .A(KEYINPUT25), .B(n1315), .ZN(n1358) );
NAND2_X1 U1036 ( .A1(n1359), .A2(n1360), .ZN(n1351) );
XOR2_X1 U1037 ( .A(KEYINPUT32), .B(G217), .Z(n1360) );
NOR3_X1 U1038 ( .A1(n1361), .A2(n1317), .A3(n1101), .ZN(n1256) );
INV_X1 U1039 ( .A(n1299), .ZN(n1101) );
NOR2_X1 U1040 ( .A1(n1104), .A2(n1103), .ZN(n1299) );
INV_X1 U1041 ( .A(n1326), .ZN(n1103) );
NAND2_X1 U1042 ( .A1(G221), .A2(n1362), .ZN(n1326) );
XOR2_X1 U1043 ( .A(n1363), .B(G469), .Z(n1104) );
NAND2_X1 U1044 ( .A1(n1364), .A2(n1365), .ZN(n1363) );
XNOR2_X1 U1045 ( .A(KEYINPUT31), .B(n1253), .ZN(n1365) );
XOR2_X1 U1046 ( .A(n1366), .B(n1367), .Z(n1364) );
XNOR2_X1 U1047 ( .A(n1368), .B(n1369), .ZN(n1367) );
INV_X1 U1048 ( .A(n1246), .ZN(n1369) );
XNOR2_X1 U1049 ( .A(n1370), .B(n1371), .ZN(n1246) );
XNOR2_X1 U1050 ( .A(KEYINPUT47), .B(n1372), .ZN(n1370) );
NOR2_X1 U1051 ( .A1(KEYINPUT33), .A2(n1373), .ZN(n1372) );
NOR2_X1 U1052 ( .A1(KEYINPUT51), .A2(n1234), .ZN(n1368) );
INV_X1 U1053 ( .A(n1238), .ZN(n1234) );
XNOR2_X1 U1054 ( .A(n1374), .B(n1375), .ZN(n1238) );
XNOR2_X1 U1055 ( .A(n1343), .B(G110), .ZN(n1375) );
NAND2_X1 U1056 ( .A1(G227), .A2(n1084), .ZN(n1374) );
XNOR2_X1 U1057 ( .A(n1241), .B(n1155), .ZN(n1366) );
NAND2_X1 U1058 ( .A1(n1376), .A2(n1377), .ZN(n1155) );
NAND2_X1 U1059 ( .A1(G128), .A2(n1378), .ZN(n1377) );
XOR2_X1 U1060 ( .A(n1379), .B(KEYINPUT19), .Z(n1376) );
OR2_X1 U1061 ( .A1(n1378), .A2(G128), .ZN(n1379) );
AND2_X1 U1062 ( .A1(n1116), .A2(n1380), .ZN(n1317) );
NAND3_X1 U1063 ( .A1(G902), .A2(n1313), .A3(n1172), .ZN(n1380) );
NOR2_X1 U1064 ( .A1(n1084), .A2(G898), .ZN(n1172) );
NAND3_X1 U1065 ( .A1(n1313), .A2(n1084), .A3(G952), .ZN(n1116) );
NAND2_X1 U1066 ( .A1(G237), .A2(G234), .ZN(n1313) );
INV_X1 U1067 ( .A(n1283), .ZN(n1361) );
NOR2_X1 U1068 ( .A1(n1115), .A2(n1114), .ZN(n1283) );
AND2_X1 U1069 ( .A1(G214), .A2(n1381), .ZN(n1114) );
INV_X1 U1070 ( .A(n1133), .ZN(n1115) );
XOR2_X1 U1071 ( .A(n1382), .B(n1252), .Z(n1133) );
NAND2_X1 U1072 ( .A1(G210), .A2(n1381), .ZN(n1252) );
NAND2_X1 U1073 ( .A1(n1383), .A2(n1253), .ZN(n1381) );
INV_X1 U1074 ( .A(G237), .ZN(n1383) );
NAND2_X1 U1075 ( .A1(n1384), .A2(n1253), .ZN(n1382) );
XOR2_X1 U1076 ( .A(n1250), .B(n1385), .Z(n1384) );
XOR2_X1 U1077 ( .A(n1284), .B(n1386), .Z(n1385) );
NAND2_X1 U1078 ( .A1(KEYINPUT40), .A2(n1387), .ZN(n1386) );
INV_X1 U1079 ( .A(n1286), .ZN(n1387) );
NAND2_X1 U1080 ( .A1(G224), .A2(n1084), .ZN(n1286) );
NAND2_X1 U1081 ( .A1(n1388), .A2(n1389), .ZN(n1284) );
OR2_X1 U1082 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
XOR2_X1 U1083 ( .A(n1392), .B(KEYINPUT20), .Z(n1388) );
NAND2_X1 U1084 ( .A1(n1391), .A2(n1390), .ZN(n1392) );
NAND2_X1 U1085 ( .A1(n1393), .A2(n1394), .ZN(n1390) );
NAND2_X1 U1086 ( .A1(n1179), .A2(n1183), .ZN(n1394) );
XOR2_X1 U1087 ( .A(KEYINPUT41), .B(n1395), .Z(n1393) );
NOR2_X1 U1088 ( .A1(n1179), .A2(n1183), .ZN(n1395) );
XOR2_X1 U1089 ( .A(G101), .B(n1371), .Z(n1179) );
XOR2_X1 U1090 ( .A(G104), .B(G107), .Z(n1371) );
INV_X1 U1091 ( .A(n1182), .ZN(n1391) );
XOR2_X1 U1092 ( .A(G110), .B(n1315), .Z(n1182) );
INV_X1 U1093 ( .A(G122), .ZN(n1315) );
XNOR2_X1 U1094 ( .A(n1396), .B(n1311), .ZN(n1250) );
INV_X1 U1095 ( .A(G125), .ZN(n1311) );
INV_X1 U1096 ( .A(n1271), .ZN(n1109) );
NAND2_X1 U1097 ( .A1(n1308), .A2(n1320), .ZN(n1271) );
XOR2_X1 U1098 ( .A(n1125), .B(KEYINPUT3), .Z(n1320) );
XNOR2_X1 U1099 ( .A(n1397), .B(G472), .ZN(n1125) );
NAND2_X1 U1100 ( .A1(n1398), .A2(n1253), .ZN(n1397) );
XOR2_X1 U1101 ( .A(n1399), .B(n1400), .Z(n1398) );
XNOR2_X1 U1102 ( .A(n1401), .B(n1224), .ZN(n1400) );
XOR2_X1 U1103 ( .A(n1396), .B(KEYINPUT35), .Z(n1224) );
XNOR2_X1 U1104 ( .A(G128), .B(n1378), .ZN(n1396) );
XOR2_X1 U1105 ( .A(G143), .B(G146), .Z(n1378) );
NOR2_X1 U1106 ( .A1(KEYINPUT46), .A2(n1175), .ZN(n1401) );
INV_X1 U1107 ( .A(n1183), .ZN(n1175) );
XOR2_X1 U1108 ( .A(G113), .B(n1402), .Z(n1183) );
XOR2_X1 U1109 ( .A(G119), .B(G116), .Z(n1402) );
XNOR2_X1 U1110 ( .A(n1225), .B(n1403), .ZN(n1399) );
NOR2_X1 U1111 ( .A1(n1404), .A2(n1405), .ZN(n1403) );
XOR2_X1 U1112 ( .A(KEYINPUT27), .B(n1406), .Z(n1405) );
NOR2_X1 U1113 ( .A1(n1373), .A2(n1227), .ZN(n1406) );
AND2_X1 U1114 ( .A1(n1373), .A2(n1227), .ZN(n1404) );
NAND2_X1 U1115 ( .A1(n1344), .A2(G210), .ZN(n1227) );
NOR2_X1 U1116 ( .A1(G953), .A2(G237), .ZN(n1344) );
INV_X1 U1117 ( .A(G101), .ZN(n1373) );
INV_X1 U1118 ( .A(n1241), .ZN(n1225) );
NAND3_X1 U1119 ( .A1(n1407), .A2(n1408), .A3(n1409), .ZN(n1241) );
OR2_X1 U1120 ( .A1(n1410), .A2(n1160), .ZN(n1409) );
NAND2_X1 U1121 ( .A1(KEYINPUT34), .A2(n1411), .ZN(n1408) );
NAND2_X1 U1122 ( .A1(n1412), .A2(n1410), .ZN(n1411) );
XNOR2_X1 U1123 ( .A(KEYINPUT49), .B(n1160), .ZN(n1412) );
NAND2_X1 U1124 ( .A1(n1413), .A2(n1414), .ZN(n1407) );
INV_X1 U1125 ( .A(KEYINPUT34), .ZN(n1414) );
NAND2_X1 U1126 ( .A1(n1415), .A2(n1416), .ZN(n1413) );
OR2_X1 U1127 ( .A1(n1160), .A2(KEYINPUT49), .ZN(n1416) );
NAND3_X1 U1128 ( .A1(n1160), .A2(n1410), .A3(KEYINPUT49), .ZN(n1415) );
XNOR2_X1 U1129 ( .A(G134), .B(n1294), .ZN(n1410) );
XOR2_X1 U1130 ( .A(G131), .B(KEYINPUT42), .Z(n1160) );
XNOR2_X1 U1131 ( .A(n1417), .B(n1128), .ZN(n1308) );
NAND2_X1 U1132 ( .A1(G217), .A2(n1362), .ZN(n1128) );
NAND2_X1 U1133 ( .A1(G234), .A2(n1253), .ZN(n1362) );
INV_X1 U1134 ( .A(G902), .ZN(n1253) );
NAND2_X1 U1135 ( .A1(KEYINPUT6), .A2(n1129), .ZN(n1417) );
NAND2_X1 U1136 ( .A1(n1418), .A2(n1195), .ZN(n1129) );
XNOR2_X1 U1137 ( .A(n1419), .B(n1420), .ZN(n1195) );
AND2_X1 U1138 ( .A1(G221), .A2(n1359), .ZN(n1420) );
AND2_X1 U1139 ( .A1(G234), .A2(n1084), .ZN(n1359) );
INV_X1 U1140 ( .A(G953), .ZN(n1084) );
XNOR2_X1 U1141 ( .A(n1421), .B(n1294), .ZN(n1419) );
INV_X1 U1142 ( .A(G137), .ZN(n1294) );
NAND2_X1 U1143 ( .A1(n1422), .A2(KEYINPUT54), .ZN(n1421) );
XOR2_X1 U1144 ( .A(n1423), .B(n1424), .Z(n1422) );
XOR2_X1 U1145 ( .A(G110), .B(n1425), .Z(n1424) );
NOR2_X1 U1146 ( .A1(KEYINPUT56), .A2(n1426), .ZN(n1425) );
XNOR2_X1 U1147 ( .A(G146), .B(n1427), .ZN(n1426) );
NAND2_X1 U1148 ( .A1(KEYINPUT14), .A2(n1153), .ZN(n1427) );
XNOR2_X1 U1149 ( .A(G125), .B(n1343), .ZN(n1153) );
INV_X1 U1150 ( .A(G140), .ZN(n1343) );
XNOR2_X1 U1151 ( .A(G119), .B(G128), .ZN(n1423) );
XNOR2_X1 U1152 ( .A(G902), .B(KEYINPUT45), .ZN(n1418) );
endmodule


