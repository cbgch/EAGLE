//Key = 0100011111011111111000100101101110111100000110011101110111010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311;

XNOR2_X1 U720 ( .A(G107), .B(n994), .ZN(G9) );
NOR2_X1 U721 ( .A1(n995), .A2(n996), .ZN(G75) );
NOR3_X1 U722 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n996) );
NOR3_X1 U723 ( .A1(n1000), .A2(n1001), .A3(n1002), .ZN(n998) );
NOR2_X1 U724 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
XOR2_X1 U725 ( .A(KEYINPUT26), .B(n1005), .Z(n1004) );
NOR3_X1 U726 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n1005) );
XOR2_X1 U727 ( .A(n1009), .B(KEYINPUT10), .Z(n1007) );
NOR2_X1 U728 ( .A1(n1010), .A2(n1009), .ZN(n1003) );
NOR2_X1 U729 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NOR2_X1 U730 ( .A1(n1013), .A2(n1006), .ZN(n1012) );
NOR2_X1 U731 ( .A1(n1014), .A2(n1015), .ZN(n1011) );
NOR2_X1 U732 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR2_X1 U733 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NOR2_X1 U734 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR3_X1 U735 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1016) );
NOR2_X1 U736 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NOR2_X1 U737 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NAND3_X1 U738 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n997) );
NAND3_X1 U739 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NAND2_X1 U740 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
OR3_X1 U741 ( .A1(n1000), .A2(n1009), .A3(n1037), .ZN(n1036) );
NAND2_X1 U742 ( .A1(n1038), .A2(n1039), .ZN(n1035) );
XNOR2_X1 U743 ( .A(KEYINPUT58), .B(n1009), .ZN(n1039) );
AND3_X1 U744 ( .A1(n1029), .A2(n1030), .A3(n1040), .ZN(n995) );
NAND4_X1 U745 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1029) );
NOR4_X1 U746 ( .A1(n1001), .A2(n1045), .A3(n1046), .A4(n1019), .ZN(n1044) );
XOR2_X1 U747 ( .A(n1047), .B(n1048), .Z(n1046) );
NAND2_X1 U748 ( .A1(KEYINPUT15), .A2(n1049), .ZN(n1047) );
XNOR2_X1 U749 ( .A(n1050), .B(n1051), .ZN(n1045) );
NAND2_X1 U750 ( .A1(KEYINPUT49), .A2(n1052), .ZN(n1050) );
INV_X1 U751 ( .A(n1037), .ZN(n1001) );
XOR2_X1 U752 ( .A(n1053), .B(n1054), .Z(n1043) );
NOR2_X1 U753 ( .A1(KEYINPUT19), .A2(n1055), .ZN(n1054) );
XOR2_X1 U754 ( .A(n1056), .B(KEYINPUT60), .Z(n1042) );
XOR2_X1 U755 ( .A(n1057), .B(n1058), .Z(n1041) );
XNOR2_X1 U756 ( .A(KEYINPUT17), .B(n1059), .ZN(n1058) );
NAND2_X1 U757 ( .A1(KEYINPUT22), .A2(n1060), .ZN(n1057) );
XOR2_X1 U758 ( .A(n1061), .B(n1062), .Z(G72) );
XOR2_X1 U759 ( .A(n1063), .B(n1064), .Z(n1062) );
NAND2_X1 U760 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
INV_X1 U761 ( .A(n1067), .ZN(n1066) );
XOR2_X1 U762 ( .A(n1068), .B(n1069), .Z(n1065) );
XOR2_X1 U763 ( .A(n1070), .B(G125), .Z(n1069) );
NAND2_X1 U764 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U765 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XOR2_X1 U766 ( .A(KEYINPUT32), .B(n1075), .Z(n1071) );
NOR2_X1 U767 ( .A1(n1073), .A2(n1074), .ZN(n1075) );
XNOR2_X1 U768 ( .A(KEYINPUT6), .B(n1076), .ZN(n1074) );
XNOR2_X1 U769 ( .A(G140), .B(KEYINPUT31), .ZN(n1068) );
NAND2_X1 U770 ( .A1(n1077), .A2(n1078), .ZN(n1063) );
XOR2_X1 U771 ( .A(n1030), .B(KEYINPUT33), .Z(n1077) );
NOR2_X1 U772 ( .A1(n1079), .A2(n1030), .ZN(n1061) );
AND2_X1 U773 ( .A1(G227), .A2(G900), .ZN(n1079) );
XOR2_X1 U774 ( .A(n1080), .B(n1081), .Z(G69) );
XOR2_X1 U775 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U776 ( .A1(n1084), .A2(G953), .ZN(n1083) );
NOR3_X1 U777 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
NOR2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(n1082) );
XOR2_X1 U779 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U780 ( .A1(KEYINPUT3), .A2(n1092), .ZN(n1090) );
NOR2_X1 U781 ( .A1(G898), .A2(n1030), .ZN(n1088) );
NOR2_X1 U782 ( .A1(n1093), .A2(n1030), .ZN(n1080) );
NOR2_X1 U783 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NOR3_X1 U784 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(G66) );
NOR3_X1 U785 ( .A1(n1099), .A2(n1030), .A3(n1040), .ZN(n1098) );
INV_X1 U786 ( .A(G952), .ZN(n1040) );
AND2_X1 U787 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
INV_X1 U788 ( .A(KEYINPUT41), .ZN(n1099) );
XNOR2_X1 U789 ( .A(n1101), .B(n1102), .ZN(n1096) );
NOR2_X1 U790 ( .A1(n1059), .A2(n1103), .ZN(n1102) );
NOR2_X1 U791 ( .A1(n1100), .A2(n1104), .ZN(G63) );
XOR2_X1 U792 ( .A(n1105), .B(n1106), .Z(n1104) );
OR2_X1 U793 ( .A1(n1103), .A2(n1049), .ZN(n1106) );
INV_X1 U794 ( .A(G478), .ZN(n1049) );
NAND2_X1 U795 ( .A1(KEYINPUT62), .A2(n1107), .ZN(n1105) );
NOR2_X1 U796 ( .A1(n1100), .A2(n1108), .ZN(G60) );
XOR2_X1 U797 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U798 ( .A1(n1052), .A2(n1103), .ZN(n1109) );
INV_X1 U799 ( .A(G475), .ZN(n1052) );
XNOR2_X1 U800 ( .A(G104), .B(n1111), .ZN(G6) );
NAND2_X1 U801 ( .A1(KEYINPUT12), .A2(n1112), .ZN(n1111) );
NOR2_X1 U802 ( .A1(n1100), .A2(n1113), .ZN(G57) );
XOR2_X1 U803 ( .A(n1114), .B(n1115), .Z(n1113) );
XNOR2_X1 U804 ( .A(n1116), .B(n1117), .ZN(n1115) );
NOR2_X1 U805 ( .A1(n1053), .A2(n1103), .ZN(n1117) );
INV_X1 U806 ( .A(G472), .ZN(n1053) );
XOR2_X1 U807 ( .A(n1118), .B(n1119), .Z(n1114) );
XNOR2_X1 U808 ( .A(n1120), .B(KEYINPUT55), .ZN(n1119) );
NAND2_X1 U809 ( .A1(n1121), .A2(KEYINPUT25), .ZN(n1120) );
XOR2_X1 U810 ( .A(n1122), .B(G101), .Z(n1121) );
NAND2_X1 U811 ( .A1(KEYINPUT14), .A2(n1123), .ZN(n1118) );
NOR2_X1 U812 ( .A1(n1100), .A2(n1124), .ZN(G54) );
XOR2_X1 U813 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U814 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U815 ( .A(n1129), .B(n1130), .Z(n1127) );
XOR2_X1 U816 ( .A(n1131), .B(n1132), .Z(n1125) );
NOR3_X1 U817 ( .A1(n1103), .A2(KEYINPUT21), .A3(n1133), .ZN(n1132) );
INV_X1 U818 ( .A(G469), .ZN(n1133) );
XNOR2_X1 U819 ( .A(KEYINPUT56), .B(KEYINPUT20), .ZN(n1131) );
NOR2_X1 U820 ( .A1(n1100), .A2(n1134), .ZN(G51) );
XOR2_X1 U821 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U822 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U823 ( .A1(n1139), .A2(n1103), .ZN(n1138) );
NAND2_X1 U824 ( .A1(G902), .A2(n999), .ZN(n1103) );
NAND4_X1 U825 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n999) );
XOR2_X1 U826 ( .A(KEYINPUT57), .B(n1087), .Z(n1143) );
AND2_X1 U827 ( .A1(n1144), .A2(n1145), .ZN(n1087) );
INV_X1 U828 ( .A(n1085), .ZN(n1142) );
NAND4_X1 U829 ( .A1(n1146), .A2(n994), .A3(n1147), .A4(n1148), .ZN(n1085) );
NOR3_X1 U830 ( .A1(n1112), .A2(n1149), .A3(n1150), .ZN(n1148) );
INV_X1 U831 ( .A(n1151), .ZN(n1149) );
AND2_X1 U832 ( .A1(n1152), .A2(n1153), .ZN(n1112) );
NAND2_X1 U833 ( .A1(n1154), .A2(n1153), .ZN(n994) );
AND4_X1 U834 ( .A1(n1145), .A2(n1026), .A3(n1155), .A4(n1156), .ZN(n1153) );
INV_X1 U835 ( .A(n1078), .ZN(n1141) );
NAND4_X1 U836 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1078) );
NOR4_X1 U837 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1160) );
INV_X1 U838 ( .A(n1165), .ZN(n1161) );
NAND2_X1 U839 ( .A1(n1166), .A2(n1167), .ZN(n1159) );
NAND2_X1 U840 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U841 ( .A1(n1032), .A2(n1170), .ZN(n1169) );
NAND2_X1 U842 ( .A1(n1152), .A2(n1021), .ZN(n1168) );
XOR2_X1 U843 ( .A(n1171), .B(KEYINPUT2), .Z(n1140) );
XOR2_X1 U844 ( .A(n1172), .B(n1173), .Z(n1135) );
NOR2_X1 U845 ( .A1(n1174), .A2(KEYINPUT29), .ZN(n1173) );
NOR2_X1 U846 ( .A1(n1030), .A2(G952), .ZN(n1100) );
XOR2_X1 U847 ( .A(n1175), .B(n1157), .Z(G48) );
NAND2_X1 U848 ( .A1(n1176), .A2(n1152), .ZN(n1157) );
XOR2_X1 U849 ( .A(n1177), .B(G143), .Z(G45) );
NAND2_X1 U850 ( .A1(KEYINPUT35), .A2(n1158), .ZN(n1177) );
NAND3_X1 U851 ( .A1(n1178), .A2(n1026), .A3(n1179), .ZN(n1158) );
AND3_X1 U852 ( .A1(n1021), .A2(n1180), .A3(n1181), .ZN(n1179) );
XOR2_X1 U853 ( .A(G140), .B(n1164), .Z(G42) );
AND3_X1 U854 ( .A1(n1152), .A2(n1020), .A3(n1166), .ZN(n1164) );
XOR2_X1 U855 ( .A(G137), .B(n1182), .Z(G39) );
NOR3_X1 U856 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1182) );
XOR2_X1 U857 ( .A(KEYINPUT13), .B(n1032), .Z(n1183) );
XOR2_X1 U858 ( .A(G134), .B(n1163), .Z(G36) );
NOR3_X1 U859 ( .A1(n1013), .A2(n1186), .A3(n1185), .ZN(n1163) );
XNOR2_X1 U860 ( .A(G131), .B(n1187), .ZN(G33) );
NAND4_X1 U861 ( .A1(n1188), .A2(n1189), .A3(KEYINPUT47), .A4(n1190), .ZN(n1187) );
NOR2_X1 U862 ( .A1(n1186), .A2(n1008), .ZN(n1190) );
INV_X1 U863 ( .A(n1021), .ZN(n1186) );
OR2_X1 U864 ( .A1(n1166), .A2(KEYINPUT4), .ZN(n1189) );
INV_X1 U865 ( .A(n1185), .ZN(n1166) );
NAND4_X1 U866 ( .A1(n1056), .A2(n1026), .A3(n1191), .A4(n1037), .ZN(n1185) );
NAND2_X1 U867 ( .A1(KEYINPUT4), .A2(n1192), .ZN(n1188) );
NAND4_X1 U868 ( .A1(n1056), .A2(n1193), .A3(n1026), .A4(n1037), .ZN(n1192) );
XOR2_X1 U869 ( .A(G128), .B(n1162), .Z(G30) );
AND2_X1 U870 ( .A1(n1176), .A2(n1154), .ZN(n1162) );
AND3_X1 U871 ( .A1(n1178), .A2(n1026), .A3(n1170), .ZN(n1176) );
XOR2_X1 U872 ( .A(n1194), .B(n1195), .Z(G3) );
NOR2_X1 U873 ( .A1(n1150), .A2(KEYINPUT45), .ZN(n1195) );
AND3_X1 U874 ( .A1(n1032), .A2(n1026), .A3(n1196), .ZN(n1150) );
XOR2_X1 U875 ( .A(n1172), .B(n1165), .Z(G27) );
NAND4_X1 U876 ( .A1(n1152), .A2(n1020), .A3(n1178), .A4(n1197), .ZN(n1165) );
NOR2_X1 U877 ( .A1(n1198), .A2(n1193), .ZN(n1178) );
INV_X1 U878 ( .A(n1191), .ZN(n1193) );
NAND2_X1 U879 ( .A1(n1009), .A2(n1199), .ZN(n1191) );
NAND3_X1 U880 ( .A1(G902), .A2(n1200), .A3(n1067), .ZN(n1199) );
NOR2_X1 U881 ( .A1(n1030), .A2(G900), .ZN(n1067) );
XOR2_X1 U882 ( .A(n1086), .B(n1201), .Z(G24) );
NOR2_X1 U883 ( .A1(KEYINPUT50), .A2(n1202), .ZN(n1201) );
INV_X1 U884 ( .A(n1171), .ZN(n1086) );
NAND4_X1 U885 ( .A1(n1034), .A2(n1145), .A3(n1181), .A4(n1180), .ZN(n1171) );
INV_X1 U886 ( .A(n1006), .ZN(n1034) );
NAND3_X1 U887 ( .A1(n1155), .A2(n1156), .A3(n1197), .ZN(n1006) );
XOR2_X1 U888 ( .A(n1203), .B(n1151), .Z(G21) );
NAND4_X1 U889 ( .A1(n1032), .A2(n1170), .A3(n1197), .A4(n1145), .ZN(n1151) );
INV_X1 U890 ( .A(n1184), .ZN(n1170) );
XNOR2_X1 U891 ( .A(G116), .B(n1147), .ZN(G18) );
NAND3_X1 U892 ( .A1(n1197), .A2(n1154), .A3(n1196), .ZN(n1147) );
INV_X1 U893 ( .A(n1013), .ZN(n1154) );
NAND2_X1 U894 ( .A1(n1181), .A2(n1204), .ZN(n1013) );
XNOR2_X1 U895 ( .A(G113), .B(n1146), .ZN(G15) );
NAND3_X1 U896 ( .A1(n1152), .A2(n1197), .A3(n1196), .ZN(n1146) );
AND2_X1 U897 ( .A1(n1145), .A2(n1021), .ZN(n1196) );
NAND2_X1 U898 ( .A1(n1205), .A2(n1206), .ZN(n1021) );
OR2_X1 U899 ( .A1(n1184), .A2(KEYINPUT61), .ZN(n1206) );
NAND2_X1 U900 ( .A1(n1023), .A2(n1022), .ZN(n1184) );
INV_X1 U901 ( .A(n1155), .ZN(n1022) );
NAND3_X1 U902 ( .A1(n1023), .A2(n1155), .A3(KEYINPUT61), .ZN(n1205) );
AND2_X1 U903 ( .A1(n1038), .A2(n1207), .ZN(n1145) );
INV_X1 U904 ( .A(n1198), .ZN(n1038) );
INV_X1 U905 ( .A(n1019), .ZN(n1197) );
NAND2_X1 U906 ( .A1(n1208), .A2(n1028), .ZN(n1019) );
INV_X1 U907 ( .A(n1027), .ZN(n1208) );
INV_X1 U908 ( .A(n1008), .ZN(n1152) );
NAND2_X1 U909 ( .A1(n1209), .A2(n1180), .ZN(n1008) );
XNOR2_X1 U910 ( .A(G110), .B(n1210), .ZN(G12) );
NAND3_X1 U911 ( .A1(n1144), .A2(n1207), .A3(n1211), .ZN(n1210) );
XOR2_X1 U912 ( .A(n1198), .B(KEYINPUT5), .Z(n1211) );
NAND2_X1 U913 ( .A1(n1000), .A2(n1037), .ZN(n1198) );
NAND2_X1 U914 ( .A1(G214), .A2(n1212), .ZN(n1037) );
INV_X1 U915 ( .A(n1056), .ZN(n1000) );
XNOR2_X1 U916 ( .A(n1213), .B(n1139), .ZN(n1056) );
NAND2_X1 U917 ( .A1(G210), .A2(n1212), .ZN(n1139) );
NAND2_X1 U918 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
INV_X1 U919 ( .A(G237), .ZN(n1214) );
NAND2_X1 U920 ( .A1(n1216), .A2(n1215), .ZN(n1213) );
XOR2_X1 U921 ( .A(n1217), .B(n1218), .Z(n1216) );
XOR2_X1 U922 ( .A(n1219), .B(n1137), .Z(n1218) );
XOR2_X1 U923 ( .A(n1220), .B(n1091), .Z(n1137) );
XOR2_X1 U924 ( .A(G110), .B(n1221), .Z(n1091) );
XOR2_X1 U925 ( .A(KEYINPUT39), .B(G122), .Z(n1221) );
XOR2_X1 U926 ( .A(n1092), .B(n1222), .Z(n1220) );
NOR2_X1 U927 ( .A1(G953), .A2(n1094), .ZN(n1222) );
INV_X1 U928 ( .A(G224), .ZN(n1094) );
XOR2_X1 U929 ( .A(n1223), .B(n1224), .Z(n1092) );
INV_X1 U930 ( .A(n1123), .ZN(n1224) );
XOR2_X1 U931 ( .A(n1225), .B(G101), .Z(n1223) );
NAND2_X1 U932 ( .A1(n1226), .A2(KEYINPUT28), .ZN(n1225) );
XOR2_X1 U933 ( .A(n1227), .B(G107), .Z(n1226) );
NAND2_X1 U934 ( .A1(KEYINPUT7), .A2(n1228), .ZN(n1227) );
NAND2_X1 U935 ( .A1(KEYINPUT16), .A2(n1172), .ZN(n1219) );
XOR2_X1 U936 ( .A(KEYINPUT37), .B(n1174), .Z(n1217) );
INV_X1 U937 ( .A(n1229), .ZN(n1174) );
NAND2_X1 U938 ( .A1(n1230), .A2(n1009), .ZN(n1207) );
NAND3_X1 U939 ( .A1(n1200), .A2(n1030), .A3(G952), .ZN(n1009) );
NAND4_X1 U940 ( .A1(G902), .A2(G953), .A3(n1200), .A4(n1095), .ZN(n1230) );
INV_X1 U941 ( .A(G898), .ZN(n1095) );
NAND2_X1 U942 ( .A1(G237), .A2(G234), .ZN(n1200) );
AND3_X1 U943 ( .A1(n1020), .A2(n1026), .A3(n1032), .ZN(n1144) );
INV_X1 U944 ( .A(n1015), .ZN(n1032) );
NAND2_X1 U945 ( .A1(n1209), .A2(n1204), .ZN(n1015) );
XOR2_X1 U946 ( .A(n1180), .B(KEYINPUT44), .Z(n1204) );
XNOR2_X1 U947 ( .A(n1051), .B(G475), .ZN(n1180) );
NAND2_X1 U948 ( .A1(n1231), .A2(n1215), .ZN(n1051) );
XOR2_X1 U949 ( .A(KEYINPUT27), .B(n1110), .Z(n1231) );
XNOR2_X1 U950 ( .A(n1232), .B(n1233), .ZN(n1110) );
XOR2_X1 U951 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U952 ( .A(G131), .B(n1236), .Z(n1235) );
NAND2_X1 U953 ( .A1(G214), .A2(n1237), .ZN(n1234) );
XOR2_X1 U954 ( .A(n1238), .B(n1128), .Z(n1232) );
XOR2_X1 U955 ( .A(G104), .B(G140), .Z(n1128) );
XOR2_X1 U956 ( .A(n1239), .B(n1240), .Z(n1238) );
NAND2_X1 U957 ( .A1(n1241), .A2(KEYINPUT53), .ZN(n1239) );
XOR2_X1 U958 ( .A(G113), .B(n1202), .Z(n1241) );
INV_X1 U959 ( .A(G122), .ZN(n1202) );
INV_X1 U960 ( .A(n1181), .ZN(n1209) );
XOR2_X1 U961 ( .A(n1048), .B(G478), .Z(n1181) );
NOR2_X1 U962 ( .A1(n1107), .A2(G902), .ZN(n1048) );
XNOR2_X1 U963 ( .A(n1242), .B(n1243), .ZN(n1107) );
XOR2_X1 U964 ( .A(n1244), .B(n1245), .Z(n1243) );
XOR2_X1 U965 ( .A(n1246), .B(G107), .Z(n1245) );
NAND2_X1 U966 ( .A1(KEYINPUT51), .A2(n1247), .ZN(n1246) );
XOR2_X1 U967 ( .A(G122), .B(G116), .Z(n1247) );
NAND3_X1 U968 ( .A1(n1248), .A2(n1249), .A3(G217), .ZN(n1244) );
XOR2_X1 U969 ( .A(KEYINPUT30), .B(G953), .Z(n1249) );
XOR2_X1 U970 ( .A(n1250), .B(n1251), .Z(n1242) );
XOR2_X1 U971 ( .A(KEYINPUT48), .B(G143), .Z(n1251) );
XOR2_X1 U972 ( .A(G134), .B(n1252), .Z(n1250) );
AND2_X1 U973 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U974 ( .A1(n1253), .A2(G221), .ZN(n1028) );
XOR2_X1 U975 ( .A(n1254), .B(KEYINPUT38), .Z(n1253) );
XNOR2_X1 U976 ( .A(n1255), .B(G469), .ZN(n1027) );
NAND3_X1 U977 ( .A1(n1256), .A2(n1257), .A3(n1215), .ZN(n1255) );
NAND2_X1 U978 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
INV_X1 U979 ( .A(KEYINPUT0), .ZN(n1259) );
XOR2_X1 U980 ( .A(n1260), .B(n1261), .Z(n1258) );
NAND3_X1 U981 ( .A1(n1261), .A2(n1260), .A3(KEYINPUT0), .ZN(n1256) );
XOR2_X1 U982 ( .A(G140), .B(n1262), .Z(n1260) );
INV_X1 U983 ( .A(n1129), .ZN(n1262) );
XNOR2_X1 U984 ( .A(G110), .B(n1263), .ZN(n1129) );
AND2_X1 U985 ( .A1(n1030), .A2(G227), .ZN(n1263) );
XOR2_X1 U986 ( .A(n1228), .B(n1130), .Z(n1261) );
XNOR2_X1 U987 ( .A(n1264), .B(n1265), .ZN(n1130) );
XNOR2_X1 U988 ( .A(n1073), .B(n1076), .ZN(n1265) );
XNOR2_X1 U989 ( .A(n1266), .B(n1267), .ZN(n1076) );
XOR2_X1 U990 ( .A(KEYINPUT24), .B(n1268), .Z(n1267) );
NOR2_X1 U991 ( .A1(G128), .A2(KEYINPUT42), .ZN(n1268) );
NAND2_X1 U992 ( .A1(n1269), .A2(n1270), .ZN(n1266) );
NAND2_X1 U993 ( .A1(n1271), .A2(n1175), .ZN(n1270) );
XOR2_X1 U994 ( .A(KEYINPUT34), .B(G143), .Z(n1271) );
NAND2_X1 U995 ( .A1(G146), .A2(n1272), .ZN(n1269) );
XOR2_X1 U996 ( .A(n1236), .B(KEYINPUT52), .Z(n1272) );
XOR2_X1 U997 ( .A(n1194), .B(n1273), .Z(n1264) );
XOR2_X1 U998 ( .A(KEYINPUT59), .B(G107), .Z(n1273) );
XOR2_X1 U999 ( .A(G104), .B(KEYINPUT56), .Z(n1228) );
NOR2_X1 U1000 ( .A1(n1155), .A2(n1023), .ZN(n1020) );
INV_X1 U1001 ( .A(n1156), .ZN(n1023) );
NAND3_X1 U1002 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1156) );
NAND2_X1 U1003 ( .A1(G472), .A2(n1277), .ZN(n1276) );
NAND2_X1 U1004 ( .A1(n1278), .A2(n1055), .ZN(n1277) );
NAND3_X1 U1005 ( .A1(n1279), .A2(n1055), .A3(n1280), .ZN(n1275) );
INV_X1 U1006 ( .A(n1278), .ZN(n1279) );
XOR2_X1 U1007 ( .A(n1281), .B(G472), .Z(n1278) );
XNOR2_X1 U1008 ( .A(KEYINPUT46), .B(KEYINPUT1), .ZN(n1281) );
OR2_X1 U1009 ( .A1(n1280), .A2(n1055), .ZN(n1274) );
NAND2_X1 U1010 ( .A1(n1282), .A2(n1215), .ZN(n1055) );
XOR2_X1 U1011 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U1012 ( .A(n1194), .B(n1285), .Z(n1284) );
NAND2_X1 U1013 ( .A1(KEYINPUT8), .A2(n1122), .ZN(n1285) );
NAND2_X1 U1014 ( .A1(G210), .A2(n1237), .ZN(n1122) );
NOR2_X1 U1015 ( .A1(G953), .A2(G237), .ZN(n1237) );
INV_X1 U1016 ( .A(G101), .ZN(n1194) );
XOR2_X1 U1017 ( .A(n1123), .B(n1116), .Z(n1283) );
XOR2_X1 U1018 ( .A(n1229), .B(n1073), .Z(n1116) );
XNOR2_X1 U1019 ( .A(G131), .B(n1286), .ZN(n1073) );
XOR2_X1 U1020 ( .A(G137), .B(G134), .Z(n1286) );
NAND2_X1 U1021 ( .A1(n1287), .A2(n1288), .ZN(n1229) );
NAND4_X1 U1022 ( .A1(KEYINPUT11), .A2(n1175), .A3(n1289), .A4(n1290), .ZN(n1288) );
NAND2_X1 U1023 ( .A1(n1291), .A2(n1236), .ZN(n1290) );
NAND2_X1 U1024 ( .A1(G143), .A2(n1292), .ZN(n1289) );
NAND3_X1 U1025 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(n1287) );
NAND2_X1 U1026 ( .A1(KEYINPUT11), .A2(n1175), .ZN(n1295) );
INV_X1 U1027 ( .A(G146), .ZN(n1175) );
NAND2_X1 U1028 ( .A1(n1292), .A2(n1236), .ZN(n1294) );
INV_X1 U1029 ( .A(G143), .ZN(n1236) );
XOR2_X1 U1030 ( .A(KEYINPUT40), .B(n1252), .Z(n1292) );
NAND2_X1 U1031 ( .A1(G143), .A2(n1291), .ZN(n1293) );
XOR2_X1 U1032 ( .A(KEYINPUT43), .B(n1252), .Z(n1291) );
XNOR2_X1 U1033 ( .A(G113), .B(n1296), .ZN(n1123) );
XOR2_X1 U1034 ( .A(G119), .B(G116), .Z(n1296) );
INV_X1 U1035 ( .A(KEYINPUT23), .ZN(n1280) );
XNOR2_X1 U1036 ( .A(n1060), .B(n1059), .ZN(n1155) );
NAND2_X1 U1037 ( .A1(G217), .A2(n1254), .ZN(n1059) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1215), .ZN(n1254) );
NAND2_X1 U1039 ( .A1(n1101), .A2(n1215), .ZN(n1060) );
INV_X1 U1040 ( .A(G902), .ZN(n1215) );
XNOR2_X1 U1041 ( .A(n1297), .B(n1298), .ZN(n1101) );
XNOR2_X1 U1042 ( .A(n1299), .B(n1240), .ZN(n1298) );
XNOR2_X1 U1043 ( .A(n1172), .B(G146), .ZN(n1240) );
INV_X1 U1044 ( .A(G125), .ZN(n1172) );
NAND2_X1 U1045 ( .A1(KEYINPUT18), .A2(G140), .ZN(n1299) );
XOR2_X1 U1046 ( .A(n1300), .B(n1301), .Z(n1297) );
NOR2_X1 U1047 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
XOR2_X1 U1048 ( .A(n1304), .B(KEYINPUT63), .Z(n1303) );
NAND2_X1 U1049 ( .A1(G110), .A2(n1305), .ZN(n1304) );
NOR2_X1 U1050 ( .A1(G110), .A2(n1305), .ZN(n1302) );
NAND3_X1 U1051 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1305) );
OR2_X1 U1052 ( .A1(n1203), .A2(KEYINPUT9), .ZN(n1308) );
NAND3_X1 U1053 ( .A1(KEYINPUT9), .A2(n1203), .A3(G128), .ZN(n1307) );
INV_X1 U1054 ( .A(G119), .ZN(n1203) );
NAND2_X1 U1055 ( .A1(n1309), .A2(n1252), .ZN(n1306) );
INV_X1 U1056 ( .A(G128), .ZN(n1252) );
NAND2_X1 U1057 ( .A1(KEYINPUT9), .A2(n1310), .ZN(n1309) );
XOR2_X1 U1058 ( .A(KEYINPUT36), .B(G119), .Z(n1310) );
XOR2_X1 U1059 ( .A(n1311), .B(G137), .Z(n1300) );
NAND3_X1 U1060 ( .A1(n1248), .A2(n1030), .A3(G221), .ZN(n1311) );
INV_X1 U1061 ( .A(G953), .ZN(n1030) );
XOR2_X1 U1062 ( .A(G234), .B(KEYINPUT54), .Z(n1248) );
endmodule


