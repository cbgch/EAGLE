//Key = 1111101111100011111101011111100100100011001111000100101011001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359;

NAND2_X1 U747 ( .A1(n1030), .A2(n1031), .ZN(G9) );
NAND2_X1 U748 ( .A1(G107), .A2(n1032), .ZN(n1031) );
XOR2_X1 U749 ( .A(KEYINPUT3), .B(n1033), .Z(n1030) );
NOR2_X1 U750 ( .A1(G107), .A2(n1032), .ZN(n1033) );
NAND3_X1 U751 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1032) );
XOR2_X1 U752 ( .A(n1037), .B(KEYINPUT23), .Z(n1036) );
NOR2_X1 U753 ( .A1(n1038), .A2(n1039), .ZN(G75) );
NOR3_X1 U754 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
NAND3_X1 U755 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1040) );
NAND2_X1 U756 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U757 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND4_X1 U758 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1049) );
NAND2_X1 U759 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NAND2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U761 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U762 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1054) );
OR2_X1 U764 ( .A1(n1064), .A2(n1034), .ZN(n1063) );
NAND3_X1 U765 ( .A1(n1056), .A2(n1065), .A3(n1062), .ZN(n1048) );
NAND2_X1 U766 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND3_X1 U767 ( .A1(n1068), .A2(n1069), .A3(n1050), .ZN(n1067) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
OR3_X1 U769 ( .A1(n1072), .A2(n1073), .A3(n1070), .ZN(n1068) );
NAND2_X1 U770 ( .A1(n1074), .A2(n1051), .ZN(n1066) );
INV_X1 U771 ( .A(n1075), .ZN(n1046) );
NOR3_X1 U772 ( .A1(n1076), .A2(G953), .A3(n1077), .ZN(n1038) );
INV_X1 U773 ( .A(n1043), .ZN(n1077) );
NAND4_X1 U774 ( .A1(n1078), .A2(n1050), .A3(n1079), .A4(n1080), .ZN(n1043) );
NOR4_X1 U775 ( .A1(n1060), .A2(n1081), .A3(n1082), .A4(n1070), .ZN(n1080) );
INV_X1 U776 ( .A(n1083), .ZN(n1082) );
NOR2_X1 U777 ( .A1(n1084), .A2(n1071), .ZN(n1079) );
XOR2_X1 U778 ( .A(n1085), .B(KEYINPUT14), .Z(n1084) );
XOR2_X1 U779 ( .A(n1041), .B(KEYINPUT4), .Z(n1076) );
INV_X1 U780 ( .A(G952), .ZN(n1041) );
XOR2_X1 U781 ( .A(n1086), .B(n1087), .Z(G72) );
NOR2_X1 U782 ( .A1(n1088), .A2(n1044), .ZN(n1087) );
AND2_X1 U783 ( .A1(G227), .A2(G900), .ZN(n1088) );
NAND2_X1 U784 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NAND2_X1 U785 ( .A1(n1091), .A2(n1044), .ZN(n1090) );
XNOR2_X1 U786 ( .A(n1092), .B(n1093), .ZN(n1091) );
NOR3_X1 U787 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
XOR2_X1 U788 ( .A(n1097), .B(KEYINPUT52), .Z(n1095) );
NAND3_X1 U789 ( .A1(G900), .A2(n1092), .A3(G953), .ZN(n1089) );
XNOR2_X1 U790 ( .A(n1098), .B(n1099), .ZN(n1092) );
XOR2_X1 U791 ( .A(n1100), .B(n1101), .Z(n1098) );
NOR2_X1 U792 ( .A1(KEYINPUT48), .A2(n1102), .ZN(n1101) );
XOR2_X1 U793 ( .A(KEYINPUT9), .B(n1103), .Z(n1102) );
NAND2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(G69) );
NAND2_X1 U795 ( .A1(n1106), .A2(n1044), .ZN(n1105) );
XNOR2_X1 U796 ( .A(n1107), .B(n1108), .ZN(n1106) );
NAND2_X1 U797 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
XOR2_X1 U798 ( .A(n1111), .B(KEYINPUT61), .Z(n1109) );
NAND2_X1 U799 ( .A1(n1112), .A2(G953), .ZN(n1104) );
NAND2_X1 U800 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND2_X1 U801 ( .A1(n1108), .A2(n1115), .ZN(n1114) );
INV_X1 U802 ( .A(G224), .ZN(n1115) );
NAND2_X1 U803 ( .A1(G224), .A2(n1116), .ZN(n1113) );
NAND2_X1 U804 ( .A1(G898), .A2(n1108), .ZN(n1116) );
NAND2_X1 U805 ( .A1(n1117), .A2(n1118), .ZN(n1108) );
NAND2_X1 U806 ( .A1(G953), .A2(n1119), .ZN(n1118) );
XNOR2_X1 U807 ( .A(n1120), .B(n1121), .ZN(n1117) );
XNOR2_X1 U808 ( .A(n1122), .B(n1123), .ZN(n1121) );
NAND2_X1 U809 ( .A1(KEYINPUT42), .A2(n1124), .ZN(n1123) );
NAND2_X1 U810 ( .A1(KEYINPUT27), .A2(n1125), .ZN(n1122) );
NOR2_X1 U811 ( .A1(n1126), .A2(n1127), .ZN(G66) );
XNOR2_X1 U812 ( .A(n1128), .B(n1129), .ZN(n1127) );
NAND3_X1 U813 ( .A1(n1130), .A2(G217), .A3(KEYINPUT44), .ZN(n1128) );
NOR2_X1 U814 ( .A1(n1126), .A2(n1131), .ZN(G63) );
XOR2_X1 U815 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND3_X1 U816 ( .A1(n1130), .A2(G478), .A3(KEYINPUT28), .ZN(n1132) );
NOR2_X1 U817 ( .A1(n1126), .A2(n1134), .ZN(G60) );
NOR2_X1 U818 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U819 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U820 ( .A1(KEYINPUT30), .A2(n1139), .ZN(n1138) );
AND2_X1 U821 ( .A1(G475), .A2(n1130), .ZN(n1137) );
AND2_X1 U822 ( .A1(n1139), .A2(KEYINPUT30), .ZN(n1135) );
XOR2_X1 U823 ( .A(n1140), .B(n1141), .Z(G6) );
NOR2_X1 U824 ( .A1(n1126), .A2(n1142), .ZN(G57) );
XOR2_X1 U825 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U826 ( .A1(KEYINPUT20), .A2(n1145), .ZN(n1143) );
XOR2_X1 U827 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U828 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U829 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XOR2_X1 U830 ( .A(KEYINPUT21), .B(G472), .Z(n1151) );
NAND2_X1 U831 ( .A1(n1152), .A2(n1153), .ZN(n1148) );
NAND2_X1 U832 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XOR2_X1 U833 ( .A(n1156), .B(KEYINPUT32), .Z(n1152) );
NAND2_X1 U834 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NOR2_X1 U835 ( .A1(n1126), .A2(n1159), .ZN(G54) );
XOR2_X1 U836 ( .A(n1160), .B(KEYINPUT2), .Z(n1159) );
NAND2_X1 U837 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U838 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U839 ( .A(KEYINPUT17), .B(n1165), .Z(n1161) );
NOR2_X1 U840 ( .A1(n1163), .A2(n1164), .ZN(n1165) );
NAND2_X1 U841 ( .A1(n1130), .A2(G469), .ZN(n1164) );
INV_X1 U842 ( .A(n1150), .ZN(n1130) );
XOR2_X1 U843 ( .A(n1166), .B(n1167), .Z(n1163) );
XOR2_X1 U844 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND2_X1 U845 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NAND2_X1 U846 ( .A1(G140), .A2(n1172), .ZN(n1171) );
XOR2_X1 U847 ( .A(KEYINPUT16), .B(n1173), .Z(n1170) );
NOR2_X1 U848 ( .A1(G140), .A2(n1172), .ZN(n1173) );
NAND2_X1 U849 ( .A1(n1174), .A2(n1175), .ZN(n1166) );
OR2_X1 U850 ( .A1(n1176), .A2(n1157), .ZN(n1175) );
XOR2_X1 U851 ( .A(n1177), .B(KEYINPUT62), .Z(n1174) );
NAND2_X1 U852 ( .A1(n1176), .A2(n1157), .ZN(n1177) );
XNOR2_X1 U853 ( .A(n1178), .B(n1179), .ZN(n1176) );
NOR2_X1 U854 ( .A1(KEYINPUT51), .A2(n1180), .ZN(n1179) );
NOR2_X1 U855 ( .A1(n1126), .A2(n1181), .ZN(G51) );
XOR2_X1 U856 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U857 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U858 ( .A1(n1186), .A2(n1150), .ZN(n1185) );
NAND2_X1 U859 ( .A1(G902), .A2(n1042), .ZN(n1150) );
NAND4_X1 U860 ( .A1(n1187), .A2(n1110), .A3(n1188), .A4(n1111), .ZN(n1042) );
XOR2_X1 U861 ( .A(KEYINPUT5), .B(n1189), .Z(n1188) );
NOR2_X1 U862 ( .A1(n1190), .A2(n1096), .ZN(n1189) );
NAND3_X1 U863 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1096) );
NAND3_X1 U864 ( .A1(n1034), .A2(n1194), .A3(n1195), .ZN(n1193) );
AND3_X1 U865 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1110) );
AND3_X1 U866 ( .A1(n1141), .A2(n1199), .A3(n1200), .ZN(n1198) );
NAND3_X1 U867 ( .A1(n1035), .A2(n1074), .A3(n1064), .ZN(n1141) );
NAND2_X1 U868 ( .A1(n1074), .A2(n1201), .ZN(n1197) );
NAND2_X1 U869 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NAND2_X1 U870 ( .A1(n1034), .A2(n1035), .ZN(n1203) );
AND3_X1 U871 ( .A1(n1051), .A2(n1204), .A3(n1194), .ZN(n1035) );
NAND2_X1 U872 ( .A1(n1205), .A2(n1206), .ZN(n1196) );
NAND2_X1 U873 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U874 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XOR2_X1 U875 ( .A(KEYINPUT37), .B(n1062), .Z(n1210) );
NAND2_X1 U876 ( .A1(n1194), .A2(n1072), .ZN(n1207) );
INV_X1 U877 ( .A(n1094), .ZN(n1187) );
NAND4_X1 U878 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1094) );
NAND2_X1 U879 ( .A1(n1215), .A2(n1216), .ZN(n1211) );
XOR2_X1 U880 ( .A(KEYINPUT22), .B(n1074), .Z(n1216) );
INV_X1 U881 ( .A(n1217), .ZN(n1215) );
NOR2_X1 U882 ( .A1(n1218), .A2(n1219), .ZN(n1184) );
AND2_X1 U883 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
NOR2_X1 U884 ( .A1(n1044), .A2(G952), .ZN(n1126) );
XNOR2_X1 U885 ( .A(G146), .B(n1212), .ZN(G48) );
NAND3_X1 U886 ( .A1(n1064), .A2(n1194), .A3(n1195), .ZN(n1212) );
XOR2_X1 U887 ( .A(G143), .B(n1222), .Z(G45) );
NOR2_X1 U888 ( .A1(n1217), .A2(n1223), .ZN(n1222) );
XOR2_X1 U889 ( .A(KEYINPUT10), .B(n1074), .Z(n1223) );
NAND4_X1 U890 ( .A1(n1194), .A2(n1072), .A3(n1224), .A4(n1225), .ZN(n1217) );
NOR2_X1 U891 ( .A1(n1226), .A2(n1227), .ZN(n1224) );
XNOR2_X1 U892 ( .A(n1213), .B(n1228), .ZN(G42) );
XOR2_X1 U893 ( .A(KEYINPUT29), .B(G140), .Z(n1228) );
NAND3_X1 U894 ( .A1(n1229), .A2(n1073), .A3(n1064), .ZN(n1213) );
XNOR2_X1 U895 ( .A(G137), .B(n1214), .ZN(G39) );
NAND3_X1 U896 ( .A1(n1209), .A2(n1056), .A3(n1229), .ZN(n1214) );
INV_X1 U897 ( .A(n1230), .ZN(n1209) );
XOR2_X1 U898 ( .A(n1191), .B(n1231), .Z(G36) );
NAND2_X1 U899 ( .A1(KEYINPUT45), .A2(G134), .ZN(n1231) );
NAND3_X1 U900 ( .A1(n1034), .A2(n1072), .A3(n1229), .ZN(n1191) );
NAND3_X1 U901 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(G33) );
NAND2_X1 U902 ( .A1(n1235), .A2(n1192), .ZN(n1234) );
NAND2_X1 U903 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
INV_X1 U904 ( .A(KEYINPUT35), .ZN(n1237) );
XOR2_X1 U905 ( .A(KEYINPUT25), .B(G131), .Z(n1236) );
OR3_X1 U906 ( .A1(n1192), .A2(G131), .A3(KEYINPUT35), .ZN(n1233) );
NAND3_X1 U907 ( .A1(n1229), .A2(n1072), .A3(n1064), .ZN(n1192) );
NOR4_X1 U908 ( .A1(n1238), .A2(n1058), .A3(n1227), .A4(n1070), .ZN(n1229) );
INV_X1 U909 ( .A(n1053), .ZN(n1070) );
NAND2_X1 U910 ( .A1(KEYINPUT35), .A2(G131), .ZN(n1232) );
XOR2_X1 U911 ( .A(G128), .B(n1239), .Z(G30) );
AND3_X1 U912 ( .A1(n1240), .A2(n1034), .A3(n1195), .ZN(n1239) );
NOR3_X1 U913 ( .A1(n1037), .A2(n1227), .A3(n1230), .ZN(n1195) );
XOR2_X1 U914 ( .A(KEYINPUT18), .B(n1058), .Z(n1240) );
XOR2_X1 U915 ( .A(n1241), .B(n1242), .Z(G3) );
NAND3_X1 U916 ( .A1(n1205), .A2(n1072), .A3(n1243), .ZN(n1242) );
XOR2_X1 U917 ( .A(n1058), .B(KEYINPUT43), .Z(n1243) );
INV_X1 U918 ( .A(n1194), .ZN(n1058) );
XOR2_X1 U919 ( .A(G125), .B(n1190), .Z(G27) );
INV_X1 U920 ( .A(n1097), .ZN(n1190) );
NAND3_X1 U921 ( .A1(n1062), .A2(n1064), .A3(n1244), .ZN(n1097) );
NOR3_X1 U922 ( .A1(n1245), .A2(n1227), .A3(n1037), .ZN(n1244) );
AND2_X1 U923 ( .A1(n1075), .A2(n1246), .ZN(n1227) );
NAND4_X1 U924 ( .A1(G953), .A2(G902), .A3(n1247), .A4(n1248), .ZN(n1246) );
INV_X1 U925 ( .A(G900), .ZN(n1248) );
XOR2_X1 U926 ( .A(n1249), .B(n1250), .Z(G24) );
NOR2_X1 U927 ( .A1(n1251), .A2(n1037), .ZN(n1250) );
XOR2_X1 U928 ( .A(n1202), .B(KEYINPUT41), .Z(n1251) );
NAND4_X1 U929 ( .A1(n1204), .A2(n1252), .A3(n1225), .A4(n1253), .ZN(n1202) );
NOR2_X1 U930 ( .A1(n1071), .A2(n1254), .ZN(n1253) );
INV_X1 U931 ( .A(n1051), .ZN(n1071) );
NAND2_X1 U932 ( .A1(KEYINPUT24), .A2(n1255), .ZN(n1249) );
XOR2_X1 U933 ( .A(G119), .B(n1256), .Z(G21) );
NOR3_X1 U934 ( .A1(n1254), .A2(n1257), .A3(n1230), .ZN(n1256) );
NAND2_X1 U935 ( .A1(n1258), .A2(n1259), .ZN(n1230) );
XNOR2_X1 U936 ( .A(G116), .B(n1200), .ZN(G18) );
NAND2_X1 U937 ( .A1(n1260), .A2(n1034), .ZN(n1200) );
NOR2_X1 U938 ( .A1(n1252), .A2(n1078), .ZN(n1034) );
XOR2_X1 U939 ( .A(n1199), .B(n1261), .Z(G15) );
NOR2_X1 U940 ( .A1(KEYINPUT11), .A2(n1262), .ZN(n1261) );
XOR2_X1 U941 ( .A(n1263), .B(KEYINPUT56), .Z(n1262) );
NAND2_X1 U942 ( .A1(n1260), .A2(n1064), .ZN(n1199) );
NOR2_X1 U943 ( .A1(n1225), .A2(n1226), .ZN(n1064) );
INV_X1 U944 ( .A(n1252), .ZN(n1226) );
AND4_X1 U945 ( .A1(n1062), .A2(n1074), .A3(n1072), .A4(n1204), .ZN(n1260) );
NAND2_X1 U946 ( .A1(n1264), .A2(n1265), .ZN(n1072) );
OR3_X1 U947 ( .A1(n1259), .A2(n1266), .A3(KEYINPUT58), .ZN(n1265) );
NAND2_X1 U948 ( .A1(KEYINPUT58), .A2(n1051), .ZN(n1264) );
NOR2_X1 U949 ( .A1(n1259), .A2(n1258), .ZN(n1051) );
INV_X1 U950 ( .A(n1266), .ZN(n1258) );
INV_X1 U951 ( .A(n1254), .ZN(n1062) );
NAND2_X1 U952 ( .A1(n1061), .A2(n1267), .ZN(n1254) );
XOR2_X1 U953 ( .A(n1172), .B(n1111), .Z(G12) );
NAND3_X1 U954 ( .A1(n1073), .A2(n1194), .A3(n1205), .ZN(n1111) );
INV_X1 U955 ( .A(n1257), .ZN(n1205) );
NAND3_X1 U956 ( .A1(n1074), .A2(n1204), .A3(n1056), .ZN(n1257) );
NOR2_X1 U957 ( .A1(n1225), .A2(n1252), .ZN(n1056) );
NAND2_X1 U958 ( .A1(n1268), .A2(n1083), .ZN(n1252) );
NAND2_X1 U959 ( .A1(n1269), .A2(n1270), .ZN(n1083) );
XOR2_X1 U960 ( .A(KEYINPUT26), .B(n1081), .Z(n1268) );
NOR2_X1 U961 ( .A1(n1270), .A2(n1269), .ZN(n1081) );
NOR2_X1 U962 ( .A1(n1139), .A2(G902), .ZN(n1269) );
XNOR2_X1 U963 ( .A(n1271), .B(n1272), .ZN(n1139) );
XOR2_X1 U964 ( .A(n1273), .B(n1274), .Z(n1272) );
XOR2_X1 U965 ( .A(G104), .B(n1275), .Z(n1274) );
NOR2_X1 U966 ( .A1(KEYINPUT36), .A2(n1276), .ZN(n1275) );
XOR2_X1 U967 ( .A(n1277), .B(n1278), .Z(n1276) );
NOR2_X1 U968 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NOR2_X1 U969 ( .A1(n1281), .A2(G143), .ZN(n1280) );
NOR2_X1 U970 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NOR3_X1 U971 ( .A1(n1283), .A2(n1284), .A3(n1282), .ZN(n1279) );
XOR2_X1 U972 ( .A(n1285), .B(KEYINPUT50), .Z(n1284) );
INV_X1 U973 ( .A(G214), .ZN(n1283) );
NAND2_X1 U974 ( .A1(KEYINPUT49), .A2(G131), .ZN(n1277) );
INV_X1 U975 ( .A(n1286), .ZN(n1273) );
XOR2_X1 U976 ( .A(n1263), .B(n1287), .Z(n1271) );
XOR2_X1 U977 ( .A(KEYINPUT34), .B(G122), .Z(n1287) );
XNOR2_X1 U978 ( .A(G475), .B(KEYINPUT59), .ZN(n1270) );
INV_X1 U979 ( .A(n1078), .ZN(n1225) );
XOR2_X1 U980 ( .A(n1288), .B(G478), .Z(n1078) );
NAND2_X1 U981 ( .A1(n1133), .A2(n1289), .ZN(n1288) );
XOR2_X1 U982 ( .A(n1290), .B(n1291), .Z(n1133) );
XOR2_X1 U983 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U984 ( .A(G107), .B(n1294), .Z(n1293) );
NOR2_X1 U985 ( .A1(KEYINPUT40), .A2(n1295), .ZN(n1294) );
XOR2_X1 U986 ( .A(G122), .B(G116), .Z(n1295) );
AND3_X1 U987 ( .A1(G234), .A2(n1044), .A3(G217), .ZN(n1292) );
XOR2_X1 U988 ( .A(n1296), .B(n1297), .Z(n1290) );
XOR2_X1 U989 ( .A(G143), .B(G134), .Z(n1297) );
NAND2_X1 U990 ( .A1(n1075), .A2(n1298), .ZN(n1204) );
NAND4_X1 U991 ( .A1(G953), .A2(G902), .A3(n1247), .A4(n1119), .ZN(n1298) );
INV_X1 U992 ( .A(G898), .ZN(n1119) );
NAND3_X1 U993 ( .A1(n1247), .A2(n1044), .A3(G952), .ZN(n1075) );
NAND2_X1 U994 ( .A1(G237), .A2(G234), .ZN(n1247) );
INV_X1 U995 ( .A(n1037), .ZN(n1074) );
NAND2_X1 U996 ( .A1(n1238), .A2(n1053), .ZN(n1037) );
NAND2_X1 U997 ( .A1(G214), .A2(n1299), .ZN(n1053) );
INV_X1 U998 ( .A(n1050), .ZN(n1238) );
XNOR2_X1 U999 ( .A(n1300), .B(n1186), .ZN(n1050) );
NAND2_X1 U1000 ( .A1(G210), .A2(n1299), .ZN(n1186) );
NAND2_X1 U1001 ( .A1(n1301), .A2(n1289), .ZN(n1299) );
NAND2_X1 U1002 ( .A1(n1302), .A2(n1289), .ZN(n1300) );
XOR2_X1 U1003 ( .A(n1303), .B(n1182), .Z(n1302) );
XNOR2_X1 U1004 ( .A(n1304), .B(n1120), .ZN(n1182) );
XNOR2_X1 U1005 ( .A(n1305), .B(G113), .ZN(n1120) );
NAND2_X1 U1006 ( .A1(KEYINPUT54), .A2(n1306), .ZN(n1305) );
XOR2_X1 U1007 ( .A(n1124), .B(n1125), .Z(n1304) );
XOR2_X1 U1008 ( .A(n1307), .B(n1172), .Z(n1125) );
NAND2_X1 U1009 ( .A1(KEYINPUT15), .A2(n1255), .ZN(n1307) );
INV_X1 U1010 ( .A(G122), .ZN(n1255) );
XOR2_X1 U1011 ( .A(n1308), .B(n1309), .Z(n1124) );
NAND2_X1 U1012 ( .A1(KEYINPUT19), .A2(n1140), .ZN(n1308) );
XOR2_X1 U1013 ( .A(n1310), .B(KEYINPUT46), .Z(n1303) );
NAND3_X1 U1014 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1310) );
INV_X1 U1015 ( .A(n1219), .ZN(n1313) );
NOR2_X1 U1016 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NAND3_X1 U1017 ( .A1(KEYINPUT6), .A2(n1220), .A3(n1221), .ZN(n1312) );
NAND2_X1 U1018 ( .A1(G224), .A2(n1044), .ZN(n1220) );
OR2_X1 U1019 ( .A1(n1221), .A2(KEYINPUT6), .ZN(n1311) );
XNOR2_X1 U1020 ( .A(G125), .B(n1158), .ZN(n1221) );
INV_X1 U1021 ( .A(n1154), .ZN(n1158) );
NOR2_X1 U1022 ( .A1(n1061), .A2(n1060), .ZN(n1194) );
INV_X1 U1023 ( .A(n1267), .ZN(n1060) );
NAND2_X1 U1024 ( .A1(G221), .A2(n1314), .ZN(n1267) );
NAND2_X1 U1025 ( .A1(G234), .A2(n1289), .ZN(n1314) );
XOR2_X1 U1026 ( .A(n1085), .B(KEYINPUT55), .Z(n1061) );
XOR2_X1 U1027 ( .A(n1315), .B(G469), .Z(n1085) );
NAND2_X1 U1028 ( .A1(n1316), .A2(n1289), .ZN(n1315) );
XOR2_X1 U1029 ( .A(n1317), .B(n1318), .Z(n1316) );
XOR2_X1 U1030 ( .A(n1157), .B(n1103), .Z(n1318) );
INV_X1 U1031 ( .A(n1178), .ZN(n1103) );
XOR2_X1 U1032 ( .A(n1285), .B(n1319), .Z(n1178) );
INV_X1 U1033 ( .A(G143), .ZN(n1285) );
XNOR2_X1 U1034 ( .A(n1320), .B(n1321), .ZN(n1317) );
NOR2_X1 U1035 ( .A1(KEYINPUT53), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1036 ( .A(n1168), .B(n1323), .Z(n1322) );
NAND2_X1 U1037 ( .A1(n1324), .A2(KEYINPUT57), .ZN(n1323) );
XOR2_X1 U1038 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1039 ( .A(KEYINPUT12), .B(G140), .Z(n1326) );
NAND2_X1 U1040 ( .A1(KEYINPUT1), .A2(G110), .ZN(n1325) );
NAND2_X1 U1041 ( .A1(G227), .A2(n1044), .ZN(n1168) );
NAND2_X1 U1042 ( .A1(KEYINPUT8), .A2(n1327), .ZN(n1320) );
INV_X1 U1043 ( .A(n1180), .ZN(n1327) );
XNOR2_X1 U1044 ( .A(n1309), .B(n1328), .ZN(n1180) );
XNOR2_X1 U1045 ( .A(n1329), .B(KEYINPUT63), .ZN(n1328) );
NAND2_X1 U1046 ( .A1(KEYINPUT39), .A2(n1140), .ZN(n1329) );
INV_X1 U1047 ( .A(G104), .ZN(n1140) );
XNOR2_X1 U1048 ( .A(n1241), .B(G107), .ZN(n1309) );
INV_X1 U1049 ( .A(n1245), .ZN(n1073) );
NAND2_X1 U1050 ( .A1(n1266), .A2(n1259), .ZN(n1245) );
NAND3_X1 U1051 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n1259) );
NAND2_X1 U1052 ( .A1(n1333), .A2(n1129), .ZN(n1332) );
OR3_X1 U1053 ( .A1(n1129), .A2(n1333), .A3(G902), .ZN(n1331) );
NOR2_X1 U1054 ( .A1(n1334), .A2(G234), .ZN(n1333) );
INV_X1 U1055 ( .A(G217), .ZN(n1334) );
XOR2_X1 U1056 ( .A(n1335), .B(n1336), .Z(n1129) );
XOR2_X1 U1057 ( .A(n1337), .B(n1286), .Z(n1336) );
XNOR2_X1 U1058 ( .A(G146), .B(n1099), .ZN(n1286) );
XOR2_X1 U1059 ( .A(G125), .B(G140), .Z(n1099) );
NAND2_X1 U1060 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
NAND4_X1 U1061 ( .A1(G221), .A2(G234), .A3(n1340), .A4(n1044), .ZN(n1339) );
INV_X1 U1062 ( .A(n1341), .ZN(n1340) );
XOR2_X1 U1063 ( .A(n1342), .B(KEYINPUT33), .Z(n1338) );
NAND2_X1 U1064 ( .A1(n1341), .A2(n1343), .ZN(n1342) );
NAND3_X1 U1065 ( .A1(G234), .A2(n1044), .A3(G221), .ZN(n1343) );
XNOR2_X1 U1066 ( .A(n1344), .B(KEYINPUT38), .ZN(n1341) );
XOR2_X1 U1067 ( .A(n1345), .B(n1346), .Z(n1335) );
XNOR2_X1 U1068 ( .A(G119), .B(n1347), .ZN(n1346) );
NAND2_X1 U1069 ( .A1(KEYINPUT7), .A2(n1172), .ZN(n1347) );
NAND2_X1 U1070 ( .A1(KEYINPUT31), .A2(n1296), .ZN(n1345) );
INV_X1 U1071 ( .A(G128), .ZN(n1296) );
NAND2_X1 U1072 ( .A1(G902), .A2(G217), .ZN(n1330) );
XOR2_X1 U1073 ( .A(n1348), .B(G472), .Z(n1266) );
NAND2_X1 U1074 ( .A1(n1349), .A2(n1289), .ZN(n1348) );
INV_X1 U1075 ( .A(G902), .ZN(n1289) );
XOR2_X1 U1076 ( .A(n1350), .B(n1144), .Z(n1349) );
AND2_X1 U1077 ( .A1(n1351), .A2(n1352), .ZN(n1144) );
NAND2_X1 U1078 ( .A1(n1353), .A2(n1241), .ZN(n1352) );
INV_X1 U1079 ( .A(G101), .ZN(n1241) );
NAND2_X1 U1080 ( .A1(G210), .A2(n1354), .ZN(n1353) );
NAND3_X1 U1081 ( .A1(G210), .A2(n1354), .A3(G101), .ZN(n1351) );
INV_X1 U1082 ( .A(n1282), .ZN(n1354) );
NAND2_X1 U1083 ( .A1(n1301), .A2(n1044), .ZN(n1282) );
INV_X1 U1084 ( .A(G953), .ZN(n1044) );
INV_X1 U1085 ( .A(G237), .ZN(n1301) );
XOR2_X1 U1086 ( .A(n1355), .B(n1356), .Z(n1350) );
INV_X1 U1087 ( .A(n1146), .ZN(n1356) );
XOR2_X1 U1088 ( .A(n1263), .B(n1306), .Z(n1146) );
XOR2_X1 U1089 ( .A(G116), .B(G119), .Z(n1306) );
INV_X1 U1090 ( .A(G113), .ZN(n1263) );
NAND2_X1 U1091 ( .A1(n1357), .A2(KEYINPUT60), .ZN(n1355) );
XOR2_X1 U1092 ( .A(n1154), .B(n1157), .Z(n1357) );
INV_X1 U1093 ( .A(n1155), .ZN(n1157) );
XOR2_X1 U1094 ( .A(n1100), .B(KEYINPUT47), .Z(n1155) );
XOR2_X1 U1095 ( .A(n1358), .B(n1344), .Z(n1100) );
XOR2_X1 U1096 ( .A(G137), .B(KEYINPUT0), .Z(n1344) );
XNOR2_X1 U1097 ( .A(G134), .B(G131), .ZN(n1358) );
XNOR2_X1 U1098 ( .A(n1319), .B(n1359), .ZN(n1154) );
NOR2_X1 U1099 ( .A1(G143), .A2(KEYINPUT13), .ZN(n1359) );
XOR2_X1 U1100 ( .A(G146), .B(G128), .Z(n1319) );
INV_X1 U1101 ( .A(G110), .ZN(n1172) );
endmodule


