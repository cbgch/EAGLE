//Key = 1001110100011100100011111111100001000011111011111101011100100101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310;

XNOR2_X1 U716 ( .A(G107), .B(n986), .ZN(G9) );
NOR2_X1 U717 ( .A1(n987), .A2(n988), .ZN(G75) );
NOR3_X1 U718 ( .A1(n989), .A2(n990), .A3(n991), .ZN(n988) );
XNOR2_X1 U719 ( .A(KEYINPUT40), .B(n992), .ZN(n991) );
NAND3_X1 U720 ( .A1(n993), .A2(n994), .A3(n995), .ZN(n989) );
NAND2_X1 U721 ( .A1(n996), .A2(n997), .ZN(n995) );
NAND2_X1 U722 ( .A1(n998), .A2(n999), .ZN(n997) );
NAND4_X1 U723 ( .A1(n1000), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(n999) );
NAND3_X1 U724 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1002) );
NAND2_X1 U725 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
OR2_X1 U726 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND2_X1 U727 ( .A1(n1011), .A2(n1012), .ZN(n1005) );
NAND2_X1 U728 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U729 ( .A1(KEYINPUT21), .A2(n1015), .ZN(n1014) );
OR3_X1 U730 ( .A1(n1016), .A2(KEYINPUT21), .A3(n1011), .ZN(n1004) );
INV_X1 U731 ( .A(n1015), .ZN(n1016) );
NAND3_X1 U732 ( .A1(n1007), .A2(n1017), .A3(n1011), .ZN(n998) );
NAND2_X1 U733 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND3_X1 U734 ( .A1(n1020), .A2(n1021), .A3(n1000), .ZN(n1019) );
OR2_X1 U735 ( .A1(n1003), .A2(n1001), .ZN(n1021) );
NAND3_X1 U736 ( .A1(n1022), .A2(n1023), .A3(n1003), .ZN(n1020) );
INV_X1 U737 ( .A(n1024), .ZN(n1023) );
NAND2_X1 U738 ( .A1(n1025), .A2(n1026), .ZN(n1022) );
NAND2_X1 U739 ( .A1(n1001), .A2(n1027), .ZN(n1018) );
INV_X1 U740 ( .A(n1028), .ZN(n996) );
NOR3_X1 U741 ( .A1(n1029), .A2(G953), .A3(G952), .ZN(n987) );
INV_X1 U742 ( .A(n993), .ZN(n1029) );
NAND4_X1 U743 ( .A1(n1030), .A2(n1003), .A3(n1031), .A4(n1032), .ZN(n993) );
NOR4_X1 U744 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1032) );
XNOR2_X1 U745 ( .A(KEYINPUT29), .B(n1026), .ZN(n1036) );
NOR2_X1 U746 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR3_X1 U747 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NOR2_X1 U748 ( .A1(KEYINPUT50), .A2(n1042), .ZN(n1041) );
NOR2_X1 U749 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U750 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
AND2_X1 U751 ( .A1(n1047), .A2(KEYINPUT50), .ZN(n1040) );
NOR2_X1 U752 ( .A1(KEYINPUT61), .A2(KEYINPUT19), .ZN(n1039) );
NOR2_X1 U753 ( .A1(KEYINPUT61), .A2(n1048), .ZN(n1034) );
NOR2_X1 U754 ( .A1(n1049), .A2(n1044), .ZN(n1048) );
NOR2_X1 U755 ( .A1(n1050), .A2(n1045), .ZN(n1049) );
INV_X1 U756 ( .A(KEYINPUT19), .ZN(n1045) );
NOR4_X1 U757 ( .A1(n1046), .A2(n1050), .A3(KEYINPUT19), .A4(n1044), .ZN(n1033) );
INV_X1 U758 ( .A(KEYINPUT61), .ZN(n1046) );
XOR2_X1 U759 ( .A(KEYINPUT17), .B(n1051), .Z(n1031) );
NOR4_X1 U760 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1051) );
XNOR2_X1 U761 ( .A(KEYINPUT6), .B(n1056), .ZN(n1055) );
XNOR2_X1 U762 ( .A(n1057), .B(n1058), .ZN(n1054) );
XOR2_X1 U763 ( .A(n1059), .B(n1060), .Z(n1052) );
XNOR2_X1 U764 ( .A(KEYINPUT30), .B(n1061), .ZN(n1060) );
NAND2_X1 U765 ( .A1(KEYINPUT41), .A2(n1062), .ZN(n1059) );
XOR2_X1 U766 ( .A(n1063), .B(n1064), .Z(G72) );
XOR2_X1 U767 ( .A(n1065), .B(n1066), .Z(n1064) );
NOR2_X1 U768 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
AND2_X1 U769 ( .A1(G227), .A2(G900), .ZN(n1067) );
NAND3_X1 U770 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1065) );
XOR2_X1 U771 ( .A(KEYINPUT5), .B(n1072), .Z(n1071) );
NOR2_X1 U772 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U773 ( .A1(n1073), .A2(n1074), .ZN(n1070) );
XNOR2_X1 U774 ( .A(n1075), .B(G125), .ZN(n1074) );
NAND2_X1 U775 ( .A1(KEYINPUT45), .A2(n1076), .ZN(n1075) );
AND2_X1 U776 ( .A1(n1077), .A2(n1078), .ZN(n1073) );
NAND2_X1 U777 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U778 ( .A(KEYINPUT44), .B(n1081), .Z(n1077) );
NOR2_X1 U779 ( .A1(n1079), .A2(n1082), .ZN(n1081) );
XNOR2_X1 U780 ( .A(KEYINPUT0), .B(n1080), .ZN(n1082) );
XNOR2_X1 U781 ( .A(KEYINPUT56), .B(n1083), .ZN(n1079) );
INV_X1 U782 ( .A(n1084), .ZN(n1069) );
NAND2_X1 U783 ( .A1(n1085), .A2(n994), .ZN(n1063) );
XOR2_X1 U784 ( .A(KEYINPUT16), .B(n1086), .Z(n1085) );
NAND3_X1 U785 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(G69) );
NAND2_X1 U786 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U787 ( .A1(n1092), .A2(KEYINPUT11), .ZN(n1091) );
XNOR2_X1 U788 ( .A(n1093), .B(KEYINPUT28), .ZN(n1092) );
NAND2_X1 U789 ( .A1(n1094), .A2(n1095), .ZN(n1090) );
OR2_X1 U790 ( .A1(n1093), .A2(KEYINPUT11), .ZN(n1088) );
NAND4_X1 U791 ( .A1(n1094), .A2(n1095), .A3(n1093), .A4(KEYINPUT11), .ZN(n1087) );
NOR2_X1 U792 ( .A1(n1068), .A2(n1096), .ZN(n1093) );
AND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1096) );
XNOR2_X1 U794 ( .A(G953), .B(KEYINPUT18), .ZN(n1068) );
NAND3_X1 U795 ( .A1(n1097), .A2(n994), .A3(n1098), .ZN(n1095) );
NAND2_X1 U796 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
XOR2_X1 U797 ( .A(n1101), .B(KEYINPUT43), .Z(n1094) );
NAND4_X1 U798 ( .A1(n1102), .A2(n1099), .A3(n1100), .A4(n1103), .ZN(n1101) );
NAND2_X1 U799 ( .A1(G953), .A2(n1104), .ZN(n1103) );
INV_X1 U800 ( .A(n1098), .ZN(n1102) );
XNOR2_X1 U801 ( .A(n1105), .B(n1106), .ZN(n1098) );
XNOR2_X1 U802 ( .A(n1107), .B(n1108), .ZN(n1106) );
NAND2_X1 U803 ( .A1(n1109), .A2(KEYINPUT24), .ZN(n1107) );
XNOR2_X1 U804 ( .A(G113), .B(n1110), .ZN(n1109) );
NOR2_X1 U805 ( .A1(n1111), .A2(n1112), .ZN(G66) );
XNOR2_X1 U806 ( .A(n1113), .B(n1114), .ZN(n1112) );
XNOR2_X1 U807 ( .A(KEYINPUT12), .B(n1115), .ZN(n1114) );
NOR3_X1 U808 ( .A1(n1116), .A2(KEYINPUT35), .A3(n1117), .ZN(n1115) );
NOR2_X1 U809 ( .A1(n1111), .A2(n1118), .ZN(G63) );
XOR2_X1 U810 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U811 ( .A(KEYINPUT47), .B(n1121), .Z(n1120) );
NOR2_X1 U812 ( .A1(n1122), .A2(n1116), .ZN(n1121) );
NOR2_X1 U813 ( .A1(n1111), .A2(n1123), .ZN(G60) );
XNOR2_X1 U814 ( .A(n1124), .B(n1125), .ZN(n1123) );
XOR2_X1 U815 ( .A(KEYINPUT31), .B(n1126), .Z(n1125) );
NOR2_X1 U816 ( .A1(n1061), .A2(n1116), .ZN(n1126) );
INV_X1 U817 ( .A(G475), .ZN(n1061) );
XNOR2_X1 U818 ( .A(n1127), .B(n1128), .ZN(G6) );
NOR2_X1 U819 ( .A1(KEYINPUT10), .A2(n1129), .ZN(n1128) );
NOR2_X1 U820 ( .A1(n1111), .A2(n1130), .ZN(G57) );
XOR2_X1 U821 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U822 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U823 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U824 ( .A1(n1057), .A2(n1116), .ZN(n1136) );
NAND2_X1 U825 ( .A1(KEYINPUT7), .A2(n1137), .ZN(n1135) );
NAND2_X1 U826 ( .A1(KEYINPUT48), .A2(n1138), .ZN(n1133) );
XNOR2_X1 U827 ( .A(n1139), .B(n1140), .ZN(n1131) );
NOR2_X1 U828 ( .A1(n1111), .A2(n1141), .ZN(G54) );
NOR2_X1 U829 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XOR2_X1 U830 ( .A(n1144), .B(n1145), .Z(n1143) );
NOR2_X1 U831 ( .A1(KEYINPUT52), .A2(n1146), .ZN(n1145) );
NOR2_X1 U832 ( .A1(n1147), .A2(n1116), .ZN(n1144) );
AND2_X1 U833 ( .A1(n1146), .A2(KEYINPUT52), .ZN(n1142) );
XOR2_X1 U834 ( .A(n1148), .B(n1149), .Z(n1146) );
XNOR2_X1 U835 ( .A(n1150), .B(n1076), .ZN(n1149) );
NOR2_X1 U836 ( .A1(KEYINPUT59), .A2(n1080), .ZN(n1150) );
INV_X1 U837 ( .A(n1139), .ZN(n1080) );
XNOR2_X1 U838 ( .A(n1151), .B(n1152), .ZN(n1148) );
NOR2_X1 U839 ( .A1(n1111), .A2(n1153), .ZN(G51) );
XOR2_X1 U840 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U841 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR2_X1 U842 ( .A1(n1047), .A2(n1116), .ZN(n1156) );
NAND2_X1 U843 ( .A1(G902), .A2(n1158), .ZN(n1116) );
NAND2_X1 U844 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
INV_X1 U845 ( .A(n990), .ZN(n1160) );
NAND2_X1 U846 ( .A1(n1086), .A2(n1100), .ZN(n990) );
AND4_X1 U847 ( .A1(n1127), .A2(n986), .A3(n1161), .A4(n1162), .ZN(n1100) );
NAND3_X1 U848 ( .A1(n1010), .A2(n1007), .A3(n1163), .ZN(n986) );
NAND3_X1 U849 ( .A1(n1163), .A2(n1007), .A3(n1009), .ZN(n1127) );
AND2_X1 U850 ( .A1(n1164), .A2(n1165), .ZN(n1086) );
NOR4_X1 U851 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
INV_X1 U852 ( .A(n1170), .ZN(n1169) );
INV_X1 U853 ( .A(n1171), .ZN(n1168) );
NOR4_X1 U854 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1164) );
NOR3_X1 U855 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1174) );
INV_X1 U856 ( .A(n1010), .ZN(n1177) );
XNOR2_X1 U857 ( .A(KEYINPUT39), .B(n1013), .ZN(n1176) );
XNOR2_X1 U858 ( .A(n1099), .B(KEYINPUT40), .ZN(n1159) );
INV_X1 U859 ( .A(n992), .ZN(n1099) );
NAND4_X1 U860 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n992) );
NOR2_X1 U861 ( .A1(n1183), .A2(n1184), .ZN(n1179) );
AND2_X1 U862 ( .A1(KEYINPUT46), .A2(n1185), .ZN(n1184) );
NOR4_X1 U863 ( .A1(KEYINPUT46), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1183) );
NOR2_X1 U864 ( .A1(n1189), .A2(n1190), .ZN(n1187) );
NOR2_X1 U865 ( .A1(n994), .A2(G952), .ZN(n1111) );
XNOR2_X1 U866 ( .A(n1191), .B(n1192), .ZN(G48) );
NAND2_X1 U867 ( .A1(n1193), .A2(n1194), .ZN(n1191) );
NAND3_X1 U868 ( .A1(n1027), .A2(n1195), .A3(n1196), .ZN(n1194) );
INV_X1 U869 ( .A(KEYINPUT38), .ZN(n1196) );
NAND2_X1 U870 ( .A1(n1175), .A2(KEYINPUT38), .ZN(n1193) );
NOR2_X1 U871 ( .A1(n1195), .A2(n1197), .ZN(n1175) );
NAND4_X1 U872 ( .A1(n1198), .A2(n1009), .A3(n1199), .A4(n1024), .ZN(n1195) );
AND2_X1 U873 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U874 ( .A(G143), .B(n1173), .Z(G45) );
AND4_X1 U875 ( .A1(n1202), .A2(n1203), .A3(n1053), .A4(n1204), .ZN(n1173) );
XOR2_X1 U876 ( .A(G140), .B(n1167), .Z(G42) );
AND3_X1 U877 ( .A1(n1009), .A2(n1205), .A3(n1015), .ZN(n1167) );
XOR2_X1 U878 ( .A(G137), .B(n1166), .Z(G39) );
AND2_X1 U879 ( .A1(n1205), .A2(n1206), .ZN(n1166) );
XOR2_X1 U880 ( .A(G134), .B(n1207), .Z(G36) );
NOR2_X1 U881 ( .A1(n1178), .A2(n1208), .ZN(n1207) );
XOR2_X1 U882 ( .A(G131), .B(n1172), .Z(G33) );
AND3_X1 U883 ( .A1(n1009), .A2(n1205), .A3(n1202), .ZN(n1172) );
INV_X1 U884 ( .A(n1178), .ZN(n1205) );
NAND4_X1 U885 ( .A1(n1000), .A2(n1024), .A3(n1200), .A4(n1003), .ZN(n1178) );
XNOR2_X1 U886 ( .A(G128), .B(n1170), .ZN(G30) );
NAND4_X1 U887 ( .A1(n1198), .A2(n1203), .A3(n1010), .A4(n1201), .ZN(n1170) );
AND3_X1 U888 ( .A1(n1027), .A2(n1200), .A3(n1024), .ZN(n1203) );
XNOR2_X1 U889 ( .A(G101), .B(n1161), .ZN(G3) );
NAND3_X1 U890 ( .A1(n1011), .A2(n1163), .A3(n1202), .ZN(n1161) );
XNOR2_X1 U891 ( .A(G125), .B(n1171), .ZN(G27) );
NAND4_X1 U892 ( .A1(n1027), .A2(n1200), .A3(n1009), .A4(n1209), .ZN(n1171) );
AND2_X1 U893 ( .A1(n1015), .A2(n1001), .ZN(n1209) );
NAND2_X1 U894 ( .A1(n1028), .A2(n1210), .ZN(n1200) );
NAND3_X1 U895 ( .A1(G902), .A2(n1211), .A3(n1084), .ZN(n1210) );
NOR2_X1 U896 ( .A1(n994), .A2(G900), .ZN(n1084) );
XNOR2_X1 U897 ( .A(G122), .B(n1212), .ZN(G24) );
NOR2_X1 U898 ( .A1(KEYINPUT34), .A2(n1185), .ZN(n1212) );
NOR4_X1 U899 ( .A1(n1186), .A2(n1188), .A3(n1190), .A4(n1189), .ZN(n1185) );
INV_X1 U900 ( .A(n1007), .ZN(n1188) );
NOR2_X1 U901 ( .A1(n1201), .A2(n1213), .ZN(n1007) );
XNOR2_X1 U902 ( .A(G119), .B(n1182), .ZN(G21) );
NAND2_X1 U903 ( .A1(n1214), .A2(n1206), .ZN(n1182) );
AND3_X1 U904 ( .A1(n1198), .A2(n1201), .A3(n1011), .ZN(n1206) );
XNOR2_X1 U905 ( .A(G116), .B(n1180), .ZN(G18) );
OR2_X1 U906 ( .A1(n1208), .A2(n1186), .ZN(n1180) );
NAND2_X1 U907 ( .A1(n1202), .A2(n1010), .ZN(n1208) );
NOR2_X1 U908 ( .A1(n1204), .A2(n1190), .ZN(n1010) );
INV_X1 U909 ( .A(n1053), .ZN(n1190) );
NAND2_X1 U910 ( .A1(n1215), .A2(n1216), .ZN(G15) );
NAND2_X1 U911 ( .A1(G113), .A2(n1181), .ZN(n1216) );
XOR2_X1 U912 ( .A(KEYINPUT26), .B(n1217), .Z(n1215) );
NOR2_X1 U913 ( .A1(G113), .A2(n1181), .ZN(n1217) );
NAND3_X1 U914 ( .A1(n1202), .A2(n1009), .A3(n1214), .ZN(n1181) );
INV_X1 U915 ( .A(n1186), .ZN(n1214) );
NAND2_X1 U916 ( .A1(n1001), .A2(n1218), .ZN(n1186) );
NOR2_X1 U917 ( .A1(n1219), .A2(n1025), .ZN(n1001) );
NOR2_X1 U918 ( .A1(n1053), .A2(n1189), .ZN(n1009) );
INV_X1 U919 ( .A(n1204), .ZN(n1189) );
INV_X1 U920 ( .A(n1013), .ZN(n1202) );
NAND2_X1 U921 ( .A1(n1198), .A2(n1056), .ZN(n1013) );
XNOR2_X1 U922 ( .A(n1220), .B(KEYINPUT1), .ZN(n1198) );
XNOR2_X1 U923 ( .A(G110), .B(n1162), .ZN(G12) );
NAND3_X1 U924 ( .A1(n1011), .A2(n1163), .A3(n1015), .ZN(n1162) );
NOR2_X1 U925 ( .A1(n1056), .A2(n1213), .ZN(n1015) );
INV_X1 U926 ( .A(n1220), .ZN(n1213) );
XNOR2_X1 U927 ( .A(n1221), .B(n1222), .ZN(n1220) );
XOR2_X1 U928 ( .A(KEYINPUT37), .B(n1058), .Z(n1222) );
AND2_X1 U929 ( .A1(n1223), .A2(n1224), .ZN(n1058) );
XOR2_X1 U930 ( .A(n1225), .B(n1226), .Z(n1223) );
NOR2_X1 U931 ( .A1(KEYINPUT62), .A2(n1227), .ZN(n1226) );
XOR2_X1 U932 ( .A(n1137), .B(n1228), .Z(n1227) );
XNOR2_X1 U933 ( .A(n1083), .B(n1229), .ZN(n1228) );
NOR2_X1 U934 ( .A1(KEYINPUT8), .A2(n1139), .ZN(n1229) );
XOR2_X1 U935 ( .A(n1230), .B(n1110), .Z(n1137) );
NAND2_X1 U936 ( .A1(KEYINPUT23), .A2(n1231), .ZN(n1230) );
XNOR2_X1 U937 ( .A(n1138), .B(G101), .ZN(n1225) );
AND3_X1 U938 ( .A1(n1232), .A2(n994), .A3(G210), .ZN(n1138) );
NAND2_X1 U939 ( .A1(KEYINPUT13), .A2(n1057), .ZN(n1221) );
INV_X1 U940 ( .A(G472), .ZN(n1057) );
INV_X1 U941 ( .A(n1201), .ZN(n1056) );
XOR2_X1 U942 ( .A(n1233), .B(n1117), .Z(n1201) );
NAND2_X1 U943 ( .A1(G217), .A2(n1234), .ZN(n1117) );
NAND2_X1 U944 ( .A1(n1113), .A2(n1224), .ZN(n1233) );
XNOR2_X1 U945 ( .A(n1235), .B(n1236), .ZN(n1113) );
XOR2_X1 U946 ( .A(n1237), .B(n1238), .Z(n1236) );
XNOR2_X1 U947 ( .A(n1152), .B(n1239), .ZN(n1238) );
NOR2_X1 U948 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
NOR2_X1 U949 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U950 ( .A(KEYINPUT25), .B(G119), .Z(n1242) );
NOR2_X1 U951 ( .A1(G128), .A2(n1244), .ZN(n1240) );
XOR2_X1 U952 ( .A(KEYINPUT14), .B(G119), .Z(n1244) );
XOR2_X1 U953 ( .A(n1245), .B(n1246), .Z(n1235) );
NOR2_X1 U954 ( .A1(KEYINPUT15), .A2(n1247), .ZN(n1246) );
XOR2_X1 U955 ( .A(n1248), .B(G137), .Z(n1245) );
NAND2_X1 U956 ( .A1(n1249), .A2(G221), .ZN(n1248) );
AND2_X1 U957 ( .A1(n1218), .A2(n1024), .ZN(n1163) );
NOR2_X1 U958 ( .A1(n1026), .A2(n1025), .ZN(n1024) );
INV_X1 U959 ( .A(n1030), .ZN(n1025) );
NAND2_X1 U960 ( .A1(G221), .A2(n1234), .ZN(n1030) );
NAND2_X1 U961 ( .A1(G234), .A2(n1250), .ZN(n1234) );
INV_X1 U962 ( .A(n1219), .ZN(n1026) );
XOR2_X1 U963 ( .A(n1251), .B(n1147), .Z(n1219) );
INV_X1 U964 ( .A(G469), .ZN(n1147) );
NAND2_X1 U965 ( .A1(n1252), .A2(n1224), .ZN(n1251) );
XOR2_X1 U966 ( .A(n1253), .B(n1254), .Z(n1252) );
XNOR2_X1 U967 ( .A(n1151), .B(n1076), .ZN(n1254) );
XOR2_X1 U968 ( .A(n1255), .B(n1256), .Z(n1151) );
XOR2_X1 U969 ( .A(n1257), .B(n1140), .Z(n1256) );
XNOR2_X1 U970 ( .A(n1258), .B(n1083), .ZN(n1140) );
XOR2_X1 U971 ( .A(n1259), .B(n1260), .Z(n1255) );
XOR2_X1 U972 ( .A(KEYINPUT56), .B(KEYINPUT42), .Z(n1260) );
NAND2_X1 U973 ( .A1(G227), .A2(n994), .ZN(n1259) );
XNOR2_X1 U974 ( .A(n1139), .B(n1261), .ZN(n1253) );
NOR2_X1 U975 ( .A1(KEYINPUT32), .A2(n1152), .ZN(n1261) );
XOR2_X1 U976 ( .A(G131), .B(n1262), .Z(n1139) );
XOR2_X1 U977 ( .A(G137), .B(G134), .Z(n1262) );
AND2_X1 U978 ( .A1(n1027), .A2(n1263), .ZN(n1218) );
NAND2_X1 U979 ( .A1(n1028), .A2(n1264), .ZN(n1263) );
NAND4_X1 U980 ( .A1(G953), .A2(G902), .A3(n1211), .A4(n1104), .ZN(n1264) );
INV_X1 U981 ( .A(G898), .ZN(n1104) );
NAND3_X1 U982 ( .A1(n1211), .A2(n994), .A3(G952), .ZN(n1028) );
NAND2_X1 U983 ( .A1(G237), .A2(G234), .ZN(n1211) );
INV_X1 U984 ( .A(n1197), .ZN(n1027) );
NAND2_X1 U985 ( .A1(n1265), .A2(n1003), .ZN(n1197) );
NAND2_X1 U986 ( .A1(G214), .A2(n1266), .ZN(n1003) );
XOR2_X1 U987 ( .A(n1000), .B(KEYINPUT55), .Z(n1265) );
XNOR2_X1 U988 ( .A(n1037), .B(n1044), .ZN(n1000) );
INV_X1 U989 ( .A(n1047), .ZN(n1044) );
NAND2_X1 U990 ( .A1(G210), .A2(n1266), .ZN(n1047) );
NAND2_X1 U991 ( .A1(n1250), .A2(n1232), .ZN(n1266) );
XNOR2_X1 U992 ( .A(n1224), .B(KEYINPUT20), .ZN(n1250) );
INV_X1 U993 ( .A(n1050), .ZN(n1037) );
NAND2_X1 U994 ( .A1(n1267), .A2(n1224), .ZN(n1050) );
XOR2_X1 U995 ( .A(n1268), .B(n1269), .Z(n1267) );
XNOR2_X1 U996 ( .A(n1154), .B(KEYINPUT54), .ZN(n1269) );
XOR2_X1 U997 ( .A(n1270), .B(n1271), .Z(n1154) );
INV_X1 U998 ( .A(n1108), .ZN(n1271) );
XNOR2_X1 U999 ( .A(G122), .B(n1152), .ZN(n1108) );
XNOR2_X1 U1000 ( .A(G110), .B(KEYINPUT27), .ZN(n1152) );
XOR2_X1 U1001 ( .A(n1272), .B(n1273), .Z(n1270) );
AND2_X1 U1002 ( .A1(n994), .A2(G224), .ZN(n1273) );
NAND2_X1 U1003 ( .A1(n1274), .A2(KEYINPUT4), .ZN(n1272) );
XOR2_X1 U1004 ( .A(n1105), .B(n1275), .Z(n1274) );
NOR2_X1 U1005 ( .A1(KEYINPUT2), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U1006 ( .A(n1231), .B(n1110), .ZN(n1276) );
XOR2_X1 U1007 ( .A(G116), .B(G119), .Z(n1110) );
XNOR2_X1 U1008 ( .A(n1277), .B(n1258), .ZN(n1105) );
INV_X1 U1009 ( .A(G101), .ZN(n1258) );
NAND2_X1 U1010 ( .A1(KEYINPUT33), .A2(n1257), .ZN(n1277) );
XNOR2_X1 U1011 ( .A(n1278), .B(G104), .ZN(n1257) );
INV_X1 U1012 ( .A(G107), .ZN(n1278) );
NAND2_X1 U1013 ( .A1(n1279), .A2(n1280), .ZN(n1268) );
OR2_X1 U1014 ( .A1(n1281), .A2(n1157), .ZN(n1280) );
XOR2_X1 U1015 ( .A(G125), .B(n1083), .Z(n1157) );
NAND3_X1 U1016 ( .A1(n1083), .A2(n1282), .A3(n1281), .ZN(n1279) );
INV_X1 U1017 ( .A(KEYINPUT51), .ZN(n1281) );
XOR2_X1 U1018 ( .A(G146), .B(n1283), .Z(n1083) );
NOR2_X1 U1019 ( .A1(n1053), .A2(n1204), .ZN(n1011) );
XOR2_X1 U1020 ( .A(n1284), .B(n1062), .Z(n1204) );
NAND2_X1 U1021 ( .A1(n1124), .A2(n1224), .ZN(n1062) );
XNOR2_X1 U1022 ( .A(n1285), .B(n1286), .ZN(n1124) );
XNOR2_X1 U1023 ( .A(n1247), .B(n1239), .ZN(n1286) );
XNOR2_X1 U1024 ( .A(n1192), .B(KEYINPUT58), .ZN(n1239) );
INV_X1 U1025 ( .A(G146), .ZN(n1192) );
XNOR2_X1 U1026 ( .A(n1282), .B(n1076), .ZN(n1247) );
XNOR2_X1 U1027 ( .A(G140), .B(KEYINPUT36), .ZN(n1076) );
INV_X1 U1028 ( .A(G125), .ZN(n1282) );
XOR2_X1 U1029 ( .A(n1287), .B(n1288), .Z(n1285) );
NOR2_X1 U1030 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XOR2_X1 U1031 ( .A(n1291), .B(KEYINPUT22), .Z(n1290) );
NAND3_X1 U1032 ( .A1(n1292), .A2(n1129), .A3(n1293), .ZN(n1291) );
NOR2_X1 U1033 ( .A1(n1294), .A2(n1129), .ZN(n1289) );
INV_X1 U1034 ( .A(G104), .ZN(n1129) );
AND2_X1 U1035 ( .A1(n1292), .A2(n1293), .ZN(n1294) );
XNOR2_X1 U1036 ( .A(n1295), .B(KEYINPUT63), .ZN(n1293) );
NAND2_X1 U1037 ( .A1(G122), .A2(n1231), .ZN(n1295) );
OR2_X1 U1038 ( .A1(n1231), .A2(G122), .ZN(n1292) );
INV_X1 U1039 ( .A(G113), .ZN(n1231) );
NAND2_X1 U1040 ( .A1(n1296), .A2(KEYINPUT49), .ZN(n1287) );
XOR2_X1 U1041 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U1042 ( .A(G143), .B(G131), .Z(n1298) );
NAND3_X1 U1043 ( .A1(n1232), .A2(n994), .A3(G214), .ZN(n1297) );
INV_X1 U1044 ( .A(G237), .ZN(n1232) );
XOR2_X1 U1045 ( .A(n1299), .B(KEYINPUT53), .Z(n1284) );
NAND2_X1 U1046 ( .A1(n1300), .A2(KEYINPUT3), .ZN(n1299) );
XNOR2_X1 U1047 ( .A(G475), .B(KEYINPUT60), .ZN(n1300) );
XOR2_X1 U1048 ( .A(n1301), .B(n1122), .Z(n1053) );
INV_X1 U1049 ( .A(G478), .ZN(n1122) );
NAND2_X1 U1050 ( .A1(n1119), .A2(n1224), .ZN(n1301) );
INV_X1 U1051 ( .A(G902), .ZN(n1224) );
XNOR2_X1 U1052 ( .A(n1302), .B(n1303), .ZN(n1119) );
NOR2_X1 U1053 ( .A1(KEYINPUT9), .A2(n1304), .ZN(n1303) );
XOR2_X1 U1054 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1055 ( .A(G107), .B(n1307), .ZN(n1306) );
NAND2_X1 U1056 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND2_X1 U1057 ( .A1(G134), .A2(n1283), .ZN(n1309) );
XOR2_X1 U1058 ( .A(n1310), .B(KEYINPUT57), .Z(n1308) );
OR2_X1 U1059 ( .A1(n1283), .A2(G134), .ZN(n1310) );
XNOR2_X1 U1060 ( .A(G143), .B(n1243), .ZN(n1283) );
INV_X1 U1061 ( .A(G128), .ZN(n1243) );
XNOR2_X1 U1062 ( .A(G116), .B(G122), .ZN(n1305) );
NAND2_X1 U1063 ( .A1(G217), .A2(n1249), .ZN(n1302) );
AND2_X1 U1064 ( .A1(G234), .A2(n994), .ZN(n1249) );
INV_X1 U1065 ( .A(G953), .ZN(n994) );
endmodule


