//Key = 0000011001011011000010010001100010100110000001110100101101000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383;

XNOR2_X1 U772 ( .A(G107), .B(n1055), .ZN(G9) );
NOR2_X1 U773 ( .A1(n1056), .A2(n1057), .ZN(G75) );
NOR4_X1 U774 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1057) );
XOR2_X1 U775 ( .A(KEYINPUT50), .B(n1062), .Z(n1059) );
NOR4_X1 U776 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1062) );
NAND4_X1 U777 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1058) );
NAND4_X1 U778 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1068) );
NAND2_X1 U779 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U780 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
OR2_X1 U781 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U782 ( .A1(n1081), .A2(n1082), .ZN(n1075) );
NAND2_X1 U783 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U784 ( .A(KEYINPUT49), .B(n1085), .Z(n1083) );
NOR2_X1 U785 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U786 ( .A1(n1088), .A2(n1089), .ZN(n1067) );
NAND3_X1 U787 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
NAND2_X1 U788 ( .A1(n1073), .A2(n1093), .ZN(n1092) );
NAND2_X1 U789 ( .A1(n1094), .A2(n1072), .ZN(n1090) );
INV_X1 U790 ( .A(n1065), .ZN(n1088) );
NAND3_X1 U791 ( .A1(n1081), .A2(n1077), .A3(n1071), .ZN(n1065) );
INV_X1 U792 ( .A(n1095), .ZN(n1071) );
NOR3_X1 U793 ( .A1(n1096), .A2(G953), .A3(G952), .ZN(n1056) );
INV_X1 U794 ( .A(n1069), .ZN(n1096) );
NAND4_X1 U795 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1069) );
NOR4_X1 U796 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1100) );
XNOR2_X1 U797 ( .A(n1105), .B(n1106), .ZN(n1104) );
XOR2_X1 U798 ( .A(KEYINPUT63), .B(KEYINPUT4), .Z(n1106) );
XNOR2_X1 U799 ( .A(G478), .B(n1107), .ZN(n1102) );
NOR2_X1 U800 ( .A1(n1108), .A2(KEYINPUT29), .ZN(n1107) );
XNOR2_X1 U801 ( .A(n1109), .B(G472), .ZN(n1099) );
XNOR2_X1 U802 ( .A(n1110), .B(KEYINPUT2), .ZN(n1098) );
XOR2_X1 U803 ( .A(n1111), .B(G469), .Z(n1097) );
XOR2_X1 U804 ( .A(n1112), .B(n1113), .Z(G72) );
XOR2_X1 U805 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U806 ( .A1(G953), .A2(n1116), .ZN(n1115) );
NAND2_X1 U807 ( .A1(G900), .A2(G227), .ZN(n1116) );
NAND2_X1 U808 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
NAND2_X1 U809 ( .A1(G953), .A2(n1119), .ZN(n1118) );
XOR2_X1 U810 ( .A(n1120), .B(n1121), .Z(n1117) );
XNOR2_X1 U811 ( .A(n1122), .B(n1123), .ZN(n1121) );
NAND2_X1 U812 ( .A1(KEYINPUT57), .A2(n1124), .ZN(n1122) );
XNOR2_X1 U813 ( .A(n1125), .B(n1126), .ZN(n1124) );
XOR2_X1 U814 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U815 ( .A1(KEYINPUT41), .A2(n1129), .ZN(n1128) );
XOR2_X1 U816 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U817 ( .A1(G137), .A2(KEYINPUT60), .ZN(n1130) );
XNOR2_X1 U818 ( .A(G140), .B(KEYINPUT58), .ZN(n1120) );
AND2_X1 U819 ( .A1(n1061), .A2(n1070), .ZN(n1112) );
XOR2_X1 U820 ( .A(n1132), .B(n1133), .Z(G69) );
NOR2_X1 U821 ( .A1(n1134), .A2(n1070), .ZN(n1133) );
NOR2_X1 U822 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U823 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
NAND2_X1 U824 ( .A1(n1139), .A2(n1070), .ZN(n1138) );
XOR2_X1 U825 ( .A(n1060), .B(n1140), .Z(n1139) );
NAND3_X1 U826 ( .A1(G898), .A2(n1140), .A3(G953), .ZN(n1137) );
XOR2_X1 U827 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U828 ( .A(KEYINPUT48), .B(n1143), .Z(n1142) );
XNOR2_X1 U829 ( .A(n1144), .B(n1145), .ZN(n1141) );
NOR2_X1 U830 ( .A1(n1146), .A2(n1147), .ZN(G66) );
XOR2_X1 U831 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U832 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
NOR2_X1 U833 ( .A1(n1146), .A2(n1152), .ZN(G63) );
XOR2_X1 U834 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U835 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND2_X1 U836 ( .A1(KEYINPUT38), .A2(n1157), .ZN(n1153) );
NOR2_X1 U837 ( .A1(n1146), .A2(n1158), .ZN(G60) );
XOR2_X1 U838 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND2_X1 U839 ( .A1(n1150), .A2(G475), .ZN(n1159) );
XNOR2_X1 U840 ( .A(G104), .B(n1161), .ZN(G6) );
NOR2_X1 U841 ( .A1(n1146), .A2(n1162), .ZN(G57) );
XNOR2_X1 U842 ( .A(n1163), .B(n1164), .ZN(n1162) );
XNOR2_X1 U843 ( .A(n1165), .B(n1166), .ZN(n1164) );
NOR2_X1 U844 ( .A1(KEYINPUT44), .A2(n1167), .ZN(n1166) );
NOR2_X1 U845 ( .A1(KEYINPUT18), .A2(n1168), .ZN(n1165) );
XOR2_X1 U846 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U847 ( .A1(n1171), .A2(n1156), .ZN(n1170) );
NOR4_X1 U848 ( .A1(n1172), .A2(n1173), .A3(KEYINPUT26), .A4(n1174), .ZN(n1169) );
NOR2_X1 U849 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XNOR2_X1 U850 ( .A(n1177), .B(n1178), .ZN(n1176) );
NOR3_X1 U851 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1173) );
NOR3_X1 U852 ( .A1(n1177), .A2(n1181), .A3(n1178), .ZN(n1172) );
NOR3_X1 U853 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(G54) );
AND2_X1 U854 ( .A1(KEYINPUT46), .A2(n1146), .ZN(n1184) );
NOR3_X1 U855 ( .A1(KEYINPUT46), .A2(G953), .A3(G952), .ZN(n1183) );
XOR2_X1 U856 ( .A(n1185), .B(n1186), .Z(n1182) );
XNOR2_X1 U857 ( .A(n1187), .B(n1188), .ZN(n1185) );
NAND2_X1 U858 ( .A1(KEYINPUT37), .A2(n1189), .ZN(n1188) );
NAND3_X1 U859 ( .A1(n1150), .A2(G469), .A3(KEYINPUT54), .ZN(n1187) );
NOR2_X1 U860 ( .A1(n1146), .A2(n1190), .ZN(G51) );
XOR2_X1 U861 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U862 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U863 ( .A1(KEYINPUT21), .A2(n1195), .ZN(n1194) );
XNOR2_X1 U864 ( .A(n1181), .B(n1196), .ZN(n1195) );
XNOR2_X1 U865 ( .A(G125), .B(n1197), .ZN(n1196) );
NAND2_X1 U866 ( .A1(n1150), .A2(n1198), .ZN(n1193) );
INV_X1 U867 ( .A(n1156), .ZN(n1150) );
NAND2_X1 U868 ( .A1(n1199), .A2(n1200), .ZN(n1156) );
OR2_X1 U869 ( .A1(n1061), .A2(n1060), .ZN(n1200) );
NAND4_X1 U870 ( .A1(n1201), .A2(n1161), .A3(n1202), .A4(n1203), .ZN(n1060) );
AND4_X1 U871 ( .A1(n1204), .A2(n1055), .A3(n1205), .A4(n1206), .ZN(n1203) );
NAND3_X1 U872 ( .A1(n1080), .A2(n1073), .A3(n1207), .ZN(n1055) );
NOR2_X1 U873 ( .A1(n1208), .A2(n1209), .ZN(n1202) );
NOR2_X1 U874 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
AND2_X1 U875 ( .A1(n1094), .A2(n1212), .ZN(n1208) );
NAND3_X1 U876 ( .A1(n1207), .A2(n1073), .A3(n1079), .ZN(n1161) );
NAND2_X1 U877 ( .A1(n1213), .A2(n1093), .ZN(n1201) );
XOR2_X1 U878 ( .A(n1214), .B(KEYINPUT11), .Z(n1213) );
NAND4_X1 U879 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1061) );
AND4_X1 U880 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1218) );
NOR3_X1 U881 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1217) );
NOR3_X1 U882 ( .A1(n1226), .A2(n1093), .A3(n1227), .ZN(n1225) );
AND2_X1 U883 ( .A1(n1226), .A2(n1228), .ZN(n1224) );
INV_X1 U884 ( .A(KEYINPUT17), .ZN(n1226) );
INV_X1 U885 ( .A(n1229), .ZN(n1223) );
XNOR2_X1 U886 ( .A(G902), .B(KEYINPUT6), .ZN(n1199) );
NOR2_X1 U887 ( .A1(n1070), .A2(G952), .ZN(n1146) );
XNOR2_X1 U888 ( .A(G146), .B(n1229), .ZN(G48) );
NAND3_X1 U889 ( .A1(n1079), .A2(n1093), .A3(n1230), .ZN(n1229) );
NAND2_X1 U890 ( .A1(n1231), .A2(n1232), .ZN(G45) );
NAND2_X1 U891 ( .A1(KEYINPUT13), .A2(n1233), .ZN(n1232) );
XOR2_X1 U892 ( .A(n1234), .B(n1228), .Z(n1231) );
NOR2_X1 U893 ( .A1(n1227), .A2(n1235), .ZN(n1228) );
NAND3_X1 U894 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1227) );
OR2_X1 U895 ( .A1(n1233), .A2(KEYINPUT13), .ZN(n1234) );
XNOR2_X1 U896 ( .A(G140), .B(n1215), .ZN(G42) );
NAND4_X1 U897 ( .A1(n1236), .A2(n1094), .A3(n1079), .A4(n1072), .ZN(n1215) );
XNOR2_X1 U898 ( .A(G137), .B(n1216), .ZN(G39) );
NAND3_X1 U899 ( .A1(n1230), .A2(n1072), .A3(n1081), .ZN(n1216) );
XNOR2_X1 U900 ( .A(G134), .B(n1222), .ZN(G36) );
NAND3_X1 U901 ( .A1(n1236), .A2(n1080), .A3(n1239), .ZN(n1222) );
XNOR2_X1 U902 ( .A(G131), .B(n1221), .ZN(G33) );
NAND3_X1 U903 ( .A1(n1236), .A2(n1079), .A3(n1239), .ZN(n1221) );
INV_X1 U904 ( .A(n1091), .ZN(n1239) );
NAND2_X1 U905 ( .A1(n1238), .A2(n1072), .ZN(n1091) );
INV_X1 U906 ( .A(n1103), .ZN(n1072) );
NAND2_X1 U907 ( .A1(n1240), .A2(n1066), .ZN(n1103) );
INV_X1 U908 ( .A(n1064), .ZN(n1240) );
XNOR2_X1 U909 ( .A(n1220), .B(n1241), .ZN(G30) );
NOR2_X1 U910 ( .A1(KEYINPUT7), .A2(n1242), .ZN(n1241) );
INV_X1 U911 ( .A(G128), .ZN(n1242) );
NAND3_X1 U912 ( .A1(n1080), .A2(n1093), .A3(n1230), .ZN(n1220) );
AND3_X1 U913 ( .A1(n1243), .A2(n1244), .A3(n1236), .ZN(n1230) );
NOR2_X1 U914 ( .A1(n1084), .A2(n1245), .ZN(n1236) );
XNOR2_X1 U915 ( .A(G101), .B(n1204), .ZN(G3) );
NAND2_X1 U916 ( .A1(n1212), .A2(n1238), .ZN(n1204) );
XOR2_X1 U917 ( .A(n1219), .B(n1246), .Z(G27) );
NAND2_X1 U918 ( .A1(G125), .A2(n1247), .ZN(n1246) );
XOR2_X1 U919 ( .A(KEYINPUT5), .B(KEYINPUT3), .Z(n1247) );
NAND3_X1 U920 ( .A1(n1077), .A2(n1094), .A3(n1248), .ZN(n1219) );
NOR3_X1 U921 ( .A1(n1249), .A2(n1245), .A3(n1235), .ZN(n1248) );
AND2_X1 U922 ( .A1(n1250), .A2(n1095), .ZN(n1245) );
NAND4_X1 U923 ( .A1(G953), .A2(G902), .A3(n1251), .A4(n1119), .ZN(n1250) );
INV_X1 U924 ( .A(G900), .ZN(n1119) );
XNOR2_X1 U925 ( .A(G122), .B(n1252), .ZN(G24) );
NOR2_X1 U926 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NOR3_X1 U927 ( .A1(n1255), .A2(n1235), .A3(n1214), .ZN(n1254) );
NAND4_X1 U928 ( .A1(n1077), .A2(n1073), .A3(n1237), .A4(n1256), .ZN(n1214) );
INV_X1 U929 ( .A(KEYINPUT55), .ZN(n1255) );
NOR4_X1 U930 ( .A1(KEYINPUT55), .A2(n1210), .A3(n1063), .A4(n1237), .ZN(n1253) );
NAND2_X1 U931 ( .A1(n1257), .A2(n1258), .ZN(n1237) );
NAND3_X1 U932 ( .A1(n1259), .A2(n1110), .A3(n1260), .ZN(n1258) );
INV_X1 U933 ( .A(KEYINPUT8), .ZN(n1260) );
NAND2_X1 U934 ( .A1(KEYINPUT8), .A2(n1080), .ZN(n1257) );
INV_X1 U935 ( .A(n1073), .ZN(n1063) );
NOR2_X1 U936 ( .A1(n1244), .A2(n1243), .ZN(n1073) );
XOR2_X1 U937 ( .A(n1261), .B(n1262), .Z(G21) );
NOR2_X1 U938 ( .A1(KEYINPUT33), .A2(n1263), .ZN(n1262) );
NOR3_X1 U939 ( .A1(n1211), .A2(n1264), .A3(n1265), .ZN(n1261) );
NOR2_X1 U940 ( .A1(KEYINPUT12), .A2(n1266), .ZN(n1265) );
NOR3_X1 U941 ( .A1(n1235), .A2(n1077), .A3(n1267), .ZN(n1266) );
AND2_X1 U942 ( .A1(n1210), .A2(KEYINPUT12), .ZN(n1264) );
NAND3_X1 U943 ( .A1(n1243), .A2(n1244), .A3(n1081), .ZN(n1211) );
XNOR2_X1 U944 ( .A(G116), .B(n1206), .ZN(G18) );
NAND3_X1 U945 ( .A1(n1238), .A2(n1080), .A3(n1268), .ZN(n1206) );
NOR2_X1 U946 ( .A1(n1110), .A2(n1269), .ZN(n1080) );
XNOR2_X1 U947 ( .A(G113), .B(n1205), .ZN(G15) );
NAND3_X1 U948 ( .A1(n1238), .A2(n1079), .A3(n1268), .ZN(n1205) );
INV_X1 U949 ( .A(n1210), .ZN(n1268) );
NAND3_X1 U950 ( .A1(n1093), .A2(n1256), .A3(n1077), .ZN(n1210) );
NOR2_X1 U951 ( .A1(n1086), .A2(n1101), .ZN(n1077) );
INV_X1 U952 ( .A(n1087), .ZN(n1101) );
XNOR2_X1 U953 ( .A(n1270), .B(KEYINPUT45), .ZN(n1086) );
INV_X1 U954 ( .A(n1235), .ZN(n1093) );
INV_X1 U955 ( .A(n1249), .ZN(n1079) );
NAND2_X1 U956 ( .A1(n1269), .A2(n1110), .ZN(n1249) );
AND2_X1 U957 ( .A1(n1105), .A2(n1243), .ZN(n1238) );
XNOR2_X1 U958 ( .A(G110), .B(n1271), .ZN(G12) );
NAND2_X1 U959 ( .A1(n1212), .A2(n1272), .ZN(n1271) );
XOR2_X1 U960 ( .A(KEYINPUT59), .B(n1094), .Z(n1272) );
NOR2_X1 U961 ( .A1(n1243), .A2(n1105), .ZN(n1094) );
INV_X1 U962 ( .A(n1244), .ZN(n1105) );
XNOR2_X1 U963 ( .A(n1273), .B(n1151), .ZN(n1244) );
AND2_X1 U964 ( .A1(G217), .A2(n1274), .ZN(n1151) );
NAND2_X1 U965 ( .A1(n1149), .A2(n1275), .ZN(n1273) );
XOR2_X1 U966 ( .A(n1276), .B(n1277), .Z(n1149) );
NOR2_X1 U967 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
INV_X1 U968 ( .A(G221), .ZN(n1278) );
XNOR2_X1 U969 ( .A(n1280), .B(n1281), .ZN(n1276) );
NAND3_X1 U970 ( .A1(KEYINPUT32), .A2(n1282), .A3(n1283), .ZN(n1280) );
XOR2_X1 U971 ( .A(n1284), .B(KEYINPUT30), .Z(n1283) );
NAND2_X1 U972 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
OR2_X1 U973 ( .A1(n1286), .A2(n1285), .ZN(n1282) );
XNOR2_X1 U974 ( .A(n1287), .B(G110), .ZN(n1285) );
NAND2_X1 U975 ( .A1(KEYINPUT34), .A2(n1288), .ZN(n1287) );
XNOR2_X1 U976 ( .A(n1263), .B(n1289), .ZN(n1288) );
NAND3_X1 U977 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1286) );
NAND2_X1 U978 ( .A1(G146), .A2(n1293), .ZN(n1292) );
OR3_X1 U979 ( .A1(n1293), .A2(G146), .A3(KEYINPUT1), .ZN(n1291) );
NAND2_X1 U980 ( .A1(KEYINPUT9), .A2(n1294), .ZN(n1293) );
INV_X1 U981 ( .A(n1295), .ZN(n1294) );
NAND2_X1 U982 ( .A1(n1295), .A2(KEYINPUT1), .ZN(n1290) );
XOR2_X1 U983 ( .A(G125), .B(n1296), .Z(n1295) );
NOR2_X1 U984 ( .A1(G140), .A2(KEYINPUT43), .ZN(n1296) );
XOR2_X1 U985 ( .A(n1297), .B(n1171), .Z(n1243) );
INV_X1 U986 ( .A(G472), .ZN(n1171) );
NAND2_X1 U987 ( .A1(KEYINPUT20), .A2(n1109), .ZN(n1297) );
AND2_X1 U988 ( .A1(n1298), .A2(n1275), .ZN(n1109) );
XOR2_X1 U989 ( .A(n1299), .B(n1300), .Z(n1298) );
XNOR2_X1 U990 ( .A(n1167), .B(n1163), .ZN(n1300) );
NAND3_X1 U991 ( .A1(n1301), .A2(n1070), .A3(G210), .ZN(n1167) );
INV_X1 U992 ( .A(G237), .ZN(n1301) );
XNOR2_X1 U993 ( .A(n1177), .B(n1302), .ZN(n1299) );
XOR2_X1 U994 ( .A(n1303), .B(KEYINPUT10), .Z(n1302) );
NAND3_X1 U995 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n1303) );
NAND2_X1 U996 ( .A1(n1180), .A2(n1175), .ZN(n1306) );
NAND2_X1 U997 ( .A1(KEYINPUT39), .A2(n1307), .ZN(n1305) );
NAND2_X1 U998 ( .A1(n1178), .A2(n1308), .ZN(n1307) );
XNOR2_X1 U999 ( .A(n1181), .B(KEYINPUT28), .ZN(n1308) );
NAND2_X1 U1000 ( .A1(n1309), .A2(n1310), .ZN(n1304) );
INV_X1 U1001 ( .A(KEYINPUT39), .ZN(n1310) );
NAND2_X1 U1002 ( .A1(n1311), .A2(n1312), .ZN(n1309) );
NAND3_X1 U1003 ( .A1(KEYINPUT28), .A2(n1178), .A3(n1181), .ZN(n1312) );
INV_X1 U1004 ( .A(n1180), .ZN(n1178) );
XOR2_X1 U1005 ( .A(n1313), .B(n1314), .Z(n1180) );
INV_X1 U1006 ( .A(G131), .ZN(n1314) );
OR2_X1 U1007 ( .A1(n1181), .A2(KEYINPUT28), .ZN(n1311) );
INV_X1 U1008 ( .A(n1179), .ZN(n1177) );
NAND2_X1 U1009 ( .A1(n1315), .A2(n1316), .ZN(n1179) );
NAND2_X1 U1010 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
XOR2_X1 U1011 ( .A(n1319), .B(KEYINPUT25), .Z(n1315) );
NAND2_X1 U1012 ( .A1(G113), .A2(n1320), .ZN(n1319) );
INV_X1 U1013 ( .A(n1317), .ZN(n1320) );
AND2_X1 U1014 ( .A1(n1081), .A2(n1207), .ZN(n1212) );
NOR3_X1 U1015 ( .A1(n1235), .A2(n1267), .A3(n1084), .ZN(n1207) );
NAND2_X1 U1016 ( .A1(n1087), .A2(n1270), .ZN(n1084) );
NAND2_X1 U1017 ( .A1(n1321), .A2(n1322), .ZN(n1270) );
NAND2_X1 U1018 ( .A1(G469), .A2(n1111), .ZN(n1322) );
XOR2_X1 U1019 ( .A(n1323), .B(KEYINPUT22), .Z(n1321) );
OR2_X1 U1020 ( .A1(n1111), .A2(G469), .ZN(n1323) );
NAND2_X1 U1021 ( .A1(n1324), .A2(n1275), .ZN(n1111) );
XOR2_X1 U1022 ( .A(n1186), .B(n1325), .Z(n1324) );
XOR2_X1 U1023 ( .A(KEYINPUT0), .B(n1189), .Z(n1325) );
AND2_X1 U1024 ( .A1(G227), .A2(n1070), .ZN(n1189) );
XNOR2_X1 U1025 ( .A(n1326), .B(n1327), .ZN(n1186) );
XOR2_X1 U1026 ( .A(n1127), .B(n1328), .Z(n1327) );
NAND3_X1 U1027 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1127) );
OR2_X1 U1028 ( .A1(n1332), .A2(KEYINPUT19), .ZN(n1330) );
NAND2_X1 U1029 ( .A1(KEYINPUT19), .A2(n1289), .ZN(n1329) );
XOR2_X1 U1030 ( .A(n1333), .B(n1334), .Z(n1326) );
XNOR2_X1 U1031 ( .A(G110), .B(n1313), .ZN(n1334) );
NAND2_X1 U1032 ( .A1(n1335), .A2(n1336), .ZN(n1313) );
NAND2_X1 U1033 ( .A1(n1131), .A2(n1281), .ZN(n1336) );
XOR2_X1 U1034 ( .A(KEYINPUT27), .B(n1337), .Z(n1335) );
NOR2_X1 U1035 ( .A1(n1131), .A2(n1281), .ZN(n1337) );
INV_X1 U1036 ( .A(G137), .ZN(n1281) );
XOR2_X1 U1037 ( .A(G134), .B(KEYINPUT36), .Z(n1131) );
NAND2_X1 U1038 ( .A1(n1338), .A2(n1339), .ZN(n1333) );
OR2_X1 U1039 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
XOR2_X1 U1040 ( .A(n1342), .B(KEYINPUT56), .Z(n1338) );
NAND2_X1 U1041 ( .A1(n1341), .A2(n1340), .ZN(n1342) );
XNOR2_X1 U1042 ( .A(n1343), .B(KEYINPUT15), .ZN(n1340) );
NAND2_X1 U1043 ( .A1(G221), .A2(n1274), .ZN(n1087) );
NAND2_X1 U1044 ( .A1(G234), .A2(n1275), .ZN(n1274) );
INV_X1 U1045 ( .A(n1256), .ZN(n1267) );
NAND2_X1 U1046 ( .A1(n1095), .A2(n1344), .ZN(n1256) );
NAND4_X1 U1047 ( .A1(G953), .A2(G902), .A3(n1251), .A4(n1136), .ZN(n1344) );
INV_X1 U1048 ( .A(G898), .ZN(n1136) );
NAND3_X1 U1049 ( .A1(n1251), .A2(n1070), .A3(G952), .ZN(n1095) );
NAND2_X1 U1050 ( .A1(G237), .A2(G234), .ZN(n1251) );
NAND2_X1 U1051 ( .A1(n1064), .A2(n1066), .ZN(n1235) );
NAND2_X1 U1052 ( .A1(G214), .A2(n1345), .ZN(n1066) );
XNOR2_X1 U1053 ( .A(n1346), .B(n1198), .ZN(n1064) );
AND2_X1 U1054 ( .A1(G210), .A2(n1345), .ZN(n1198) );
NAND2_X1 U1055 ( .A1(n1347), .A2(n1275), .ZN(n1345) );
XOR2_X1 U1056 ( .A(KEYINPUT52), .B(G237), .Z(n1347) );
NAND2_X1 U1057 ( .A1(n1348), .A2(n1349), .ZN(n1346) );
XOR2_X1 U1058 ( .A(n1350), .B(n1351), .Z(n1349) );
XOR2_X1 U1059 ( .A(n1197), .B(n1352), .Z(n1351) );
XNOR2_X1 U1060 ( .A(KEYINPUT31), .B(n1123), .ZN(n1352) );
INV_X1 U1061 ( .A(G125), .ZN(n1123) );
NOR2_X1 U1062 ( .A1(n1135), .A2(G953), .ZN(n1197) );
INV_X1 U1063 ( .A(G224), .ZN(n1135) );
XOR2_X1 U1064 ( .A(n1191), .B(n1353), .Z(n1350) );
NOR2_X1 U1065 ( .A1(KEYINPUT35), .A2(n1181), .ZN(n1353) );
INV_X1 U1066 ( .A(n1175), .ZN(n1181) );
NAND2_X1 U1067 ( .A1(n1354), .A2(n1355), .ZN(n1175) );
NAND2_X1 U1068 ( .A1(G146), .A2(n1356), .ZN(n1355) );
NAND2_X1 U1069 ( .A1(n1331), .A2(n1332), .ZN(n1356) );
NAND2_X1 U1070 ( .A1(n1357), .A2(n1358), .ZN(n1354) );
XNOR2_X1 U1071 ( .A(n1233), .B(n1289), .ZN(n1357) );
XOR2_X1 U1072 ( .A(n1359), .B(n1143), .Z(n1191) );
XOR2_X1 U1073 ( .A(G110), .B(G122), .Z(n1143) );
NAND2_X1 U1074 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NAND2_X1 U1075 ( .A1(n1144), .A2(n1145), .ZN(n1361) );
XOR2_X1 U1076 ( .A(KEYINPUT62), .B(n1362), .Z(n1360) );
NOR2_X1 U1077 ( .A1(n1144), .A2(n1145), .ZN(n1362) );
XNOR2_X1 U1078 ( .A(n1317), .B(n1363), .ZN(n1145) );
NOR2_X1 U1079 ( .A1(KEYINPUT24), .A2(n1318), .ZN(n1363) );
XOR2_X1 U1080 ( .A(G116), .B(n1263), .Z(n1317) );
INV_X1 U1081 ( .A(G119), .ZN(n1263) );
XOR2_X1 U1082 ( .A(n1343), .B(n1341), .Z(n1144) );
INV_X1 U1083 ( .A(n1163), .ZN(n1341) );
XOR2_X1 U1084 ( .A(G101), .B(KEYINPUT40), .Z(n1163) );
XNOR2_X1 U1085 ( .A(G107), .B(n1364), .ZN(n1343) );
XNOR2_X1 U1086 ( .A(G902), .B(KEYINPUT51), .ZN(n1348) );
NOR2_X1 U1087 ( .A1(n1259), .A2(n1110), .ZN(n1081) );
XNOR2_X1 U1088 ( .A(n1365), .B(G475), .ZN(n1110) );
NAND2_X1 U1089 ( .A1(n1160), .A2(n1275), .ZN(n1365) );
XNOR2_X1 U1090 ( .A(n1366), .B(n1367), .ZN(n1160) );
XOR2_X1 U1091 ( .A(n1328), .B(n1368), .Z(n1367) );
XNOR2_X1 U1092 ( .A(n1369), .B(n1370), .ZN(n1368) );
NOR4_X1 U1093 ( .A1(KEYINPUT42), .A2(G953), .A3(G237), .A4(n1371), .ZN(n1370) );
INV_X1 U1094 ( .A(G214), .ZN(n1371) );
NOR2_X1 U1095 ( .A1(KEYINPUT53), .A2(n1372), .ZN(n1369) );
XOR2_X1 U1096 ( .A(n1364), .B(n1373), .Z(n1372) );
XNOR2_X1 U1097 ( .A(G122), .B(n1318), .ZN(n1373) );
INV_X1 U1098 ( .A(G113), .ZN(n1318) );
XOR2_X1 U1099 ( .A(G104), .B(KEYINPUT16), .Z(n1364) );
XNOR2_X1 U1100 ( .A(G140), .B(n1125), .ZN(n1328) );
XNOR2_X1 U1101 ( .A(G131), .B(n1358), .ZN(n1125) );
INV_X1 U1102 ( .A(G146), .ZN(n1358) );
XNOR2_X1 U1103 ( .A(G125), .B(n1374), .ZN(n1366) );
XNOR2_X1 U1104 ( .A(KEYINPUT23), .B(n1233), .ZN(n1374) );
INV_X1 U1105 ( .A(G143), .ZN(n1233) );
INV_X1 U1106 ( .A(n1269), .ZN(n1259) );
XOR2_X1 U1107 ( .A(n1108), .B(n1155), .Z(n1269) );
INV_X1 U1108 ( .A(G478), .ZN(n1155) );
AND2_X1 U1109 ( .A1(n1157), .A2(n1275), .ZN(n1108) );
INV_X1 U1110 ( .A(G902), .ZN(n1275) );
XOR2_X1 U1111 ( .A(n1375), .B(n1376), .Z(n1157) );
XOR2_X1 U1112 ( .A(n1377), .B(n1378), .Z(n1376) );
XOR2_X1 U1113 ( .A(n1379), .B(n1380), .Z(n1378) );
NOR2_X1 U1114 ( .A1(n1279), .A2(n1381), .ZN(n1380) );
INV_X1 U1115 ( .A(G217), .ZN(n1381) );
NAND2_X1 U1116 ( .A1(G234), .A2(n1070), .ZN(n1279) );
INV_X1 U1117 ( .A(G953), .ZN(n1070) );
NAND2_X1 U1118 ( .A1(n1382), .A2(n1331), .ZN(n1379) );
NAND2_X1 U1119 ( .A1(G143), .A2(n1289), .ZN(n1331) );
XOR2_X1 U1120 ( .A(n1332), .B(KEYINPUT61), .Z(n1382) );
OR2_X1 U1121 ( .A1(n1289), .A2(G143), .ZN(n1332) );
XOR2_X1 U1122 ( .A(G128), .B(KEYINPUT14), .Z(n1289) );
NAND2_X1 U1123 ( .A1(KEYINPUT47), .A2(G116), .ZN(n1377) );
XNOR2_X1 U1124 ( .A(G107), .B(n1383), .ZN(n1375) );
XOR2_X1 U1125 ( .A(G134), .B(G122), .Z(n1383) );
endmodule


