//Key = 0011100100111011010010000011111111110000011100110100110101110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437;

XNOR2_X1 U785 ( .A(G107), .B(n1100), .ZN(G9) );
NAND4_X1 U786 ( .A1(KEYINPUT20), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1100) );
NOR2_X1 U787 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NOR2_X1 U788 ( .A1(n1106), .A2(n1107), .ZN(G75) );
XOR2_X1 U789 ( .A(n1108), .B(KEYINPUT12), .Z(n1107) );
NAND3_X1 U790 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1108) );
NOR3_X1 U791 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
NOR2_X1 U792 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U793 ( .A1(n1117), .A2(n1118), .ZN(n1115) );
NOR3_X1 U794 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1118) );
NOR3_X1 U795 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1121) );
AND2_X1 U796 ( .A1(n1125), .A2(KEYINPUT14), .ZN(n1124) );
AND2_X1 U797 ( .A1(n1103), .A2(n1101), .ZN(n1123) );
NOR2_X1 U798 ( .A1(n1126), .A2(n1127), .ZN(n1120) );
NOR2_X1 U799 ( .A1(KEYINPUT14), .A2(n1128), .ZN(n1127) );
NOR4_X1 U800 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1117) );
NOR4_X1 U801 ( .A1(n1119), .A2(n1133), .A3(n1131), .A4(n1134), .ZN(n1113) );
XOR2_X1 U802 ( .A(n1135), .B(KEYINPUT5), .Z(n1112) );
NAND2_X1 U803 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND3_X1 U804 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1137) );
NAND2_X1 U805 ( .A1(n1141), .A2(n1142), .ZN(n1136) );
NAND2_X1 U806 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND3_X1 U807 ( .A1(n1139), .A2(n1145), .A3(n1126), .ZN(n1144) );
NAND2_X1 U808 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND2_X1 U809 ( .A1(n1148), .A2(n1103), .ZN(n1147) );
NAND2_X1 U810 ( .A1(n1140), .A2(n1149), .ZN(n1143) );
INV_X1 U811 ( .A(n1131), .ZN(n1140) );
NAND3_X1 U812 ( .A1(n1150), .A2(n1103), .A3(n1126), .ZN(n1131) );
INV_X1 U813 ( .A(n1122), .ZN(n1126) );
INV_X1 U814 ( .A(n1151), .ZN(n1110) );
NOR2_X1 U815 ( .A1(G952), .A2(n1151), .ZN(n1106) );
NAND2_X1 U816 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND4_X1 U817 ( .A1(n1154), .A2(n1132), .A3(n1155), .A4(n1156), .ZN(n1153) );
NOR4_X1 U818 ( .A1(n1157), .A2(n1116), .A3(n1158), .A4(n1159), .ZN(n1156) );
XNOR2_X1 U819 ( .A(n1130), .B(KEYINPUT3), .ZN(n1159) );
NOR2_X1 U820 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
NAND3_X1 U821 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1157) );
XNOR2_X1 U822 ( .A(G478), .B(n1165), .ZN(n1164) );
NAND2_X1 U823 ( .A1(n1166), .A2(n1167), .ZN(n1163) );
NAND2_X1 U824 ( .A1(n1168), .A2(G472), .ZN(n1162) );
NAND2_X1 U825 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND2_X1 U826 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
OR2_X1 U827 ( .A1(n1172), .A2(n1166), .ZN(n1169) );
NOR2_X1 U828 ( .A1(KEYINPUT9), .A2(n1173), .ZN(n1166) );
INV_X1 U829 ( .A(KEYINPUT52), .ZN(n1172) );
NOR3_X1 U830 ( .A1(n1174), .A2(n1129), .A3(n1175), .ZN(n1155) );
INV_X1 U831 ( .A(n1176), .ZN(n1129) );
INV_X1 U832 ( .A(n1177), .ZN(n1174) );
NAND2_X1 U833 ( .A1(n1178), .A2(n1179), .ZN(n1154) );
XNOR2_X1 U834 ( .A(G475), .B(KEYINPUT29), .ZN(n1178) );
XOR2_X1 U835 ( .A(n1180), .B(n1181), .Z(G72) );
XOR2_X1 U836 ( .A(n1182), .B(n1183), .Z(n1181) );
NAND2_X1 U837 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
INV_X1 U838 ( .A(n1186), .ZN(n1185) );
XOR2_X1 U839 ( .A(n1187), .B(n1188), .Z(n1184) );
XOR2_X1 U840 ( .A(n1189), .B(n1190), .Z(n1188) );
XNOR2_X1 U841 ( .A(G131), .B(n1191), .ZN(n1187) );
NOR2_X1 U842 ( .A1(KEYINPUT50), .A2(n1192), .ZN(n1191) );
XNOR2_X1 U843 ( .A(n1193), .B(G125), .ZN(n1192) );
NAND2_X1 U844 ( .A1(n1194), .A2(n1195), .ZN(n1182) );
XNOR2_X1 U845 ( .A(KEYINPUT42), .B(n1152), .ZN(n1194) );
NOR2_X1 U846 ( .A1(n1196), .A2(n1152), .ZN(n1180) );
AND2_X1 U847 ( .A1(G227), .A2(G900), .ZN(n1196) );
NAND2_X1 U848 ( .A1(n1197), .A2(n1198), .ZN(G69) );
NAND2_X1 U849 ( .A1(n1199), .A2(n1152), .ZN(n1198) );
XNOR2_X1 U850 ( .A(n1200), .B(n1201), .ZN(n1199) );
NAND2_X1 U851 ( .A1(n1202), .A2(G953), .ZN(n1197) );
NAND2_X1 U852 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NAND2_X1 U853 ( .A1(n1201), .A2(n1205), .ZN(n1204) );
NAND2_X1 U854 ( .A1(G224), .A2(n1206), .ZN(n1203) );
NAND2_X1 U855 ( .A1(G898), .A2(n1201), .ZN(n1206) );
NAND2_X1 U856 ( .A1(n1207), .A2(n1208), .ZN(n1201) );
NAND2_X1 U857 ( .A1(G953), .A2(n1209), .ZN(n1208) );
XOR2_X1 U858 ( .A(n1210), .B(n1211), .Z(n1207) );
XOR2_X1 U859 ( .A(n1212), .B(n1213), .Z(n1211) );
NOR2_X1 U860 ( .A1(KEYINPUT22), .A2(n1214), .ZN(n1213) );
NOR3_X1 U861 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(G66) );
AND2_X1 U862 ( .A1(KEYINPUT58), .A2(n1218), .ZN(n1217) );
NOR3_X1 U863 ( .A1(KEYINPUT58), .A2(n1152), .A3(n1219), .ZN(n1216) );
INV_X1 U864 ( .A(G952), .ZN(n1219) );
XOR2_X1 U865 ( .A(n1220), .B(n1221), .Z(n1215) );
NOR2_X1 U866 ( .A1(n1161), .A2(n1222), .ZN(n1220) );
NOR2_X1 U867 ( .A1(n1218), .A2(n1223), .ZN(G63) );
XOR2_X1 U868 ( .A(n1224), .B(n1225), .Z(n1223) );
NAND2_X1 U869 ( .A1(n1226), .A2(G478), .ZN(n1224) );
NOR2_X1 U870 ( .A1(n1218), .A2(n1227), .ZN(G60) );
XOR2_X1 U871 ( .A(n1228), .B(n1229), .Z(n1227) );
NAND3_X1 U872 ( .A1(n1226), .A2(G475), .A3(KEYINPUT33), .ZN(n1228) );
XOR2_X1 U873 ( .A(G104), .B(n1230), .Z(G6) );
NOR2_X1 U874 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NOR2_X1 U875 ( .A1(n1233), .A2(n1234), .ZN(G57) );
XOR2_X1 U876 ( .A(n1235), .B(n1236), .Z(n1234) );
NOR2_X1 U877 ( .A1(n1167), .A2(n1222), .ZN(n1235) );
INV_X1 U878 ( .A(n1226), .ZN(n1222) );
XNOR2_X1 U879 ( .A(n1218), .B(KEYINPUT10), .ZN(n1233) );
NOR2_X1 U880 ( .A1(n1218), .A2(n1237), .ZN(G54) );
XOR2_X1 U881 ( .A(n1238), .B(n1239), .Z(n1237) );
XNOR2_X1 U882 ( .A(n1240), .B(n1241), .ZN(n1239) );
XOR2_X1 U883 ( .A(n1242), .B(n1243), .Z(n1238) );
NOR2_X1 U884 ( .A1(KEYINPUT36), .A2(n1244), .ZN(n1243) );
XOR2_X1 U885 ( .A(n1245), .B(n1246), .Z(n1244) );
NOR2_X1 U886 ( .A1(KEYINPUT39), .A2(n1247), .ZN(n1245) );
NOR3_X1 U887 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1247) );
NOR2_X1 U888 ( .A1(G140), .A2(n1251), .ZN(n1250) );
NOR2_X1 U889 ( .A1(KEYINPUT40), .A2(n1252), .ZN(n1251) );
XOR2_X1 U890 ( .A(KEYINPUT54), .B(G110), .Z(n1252) );
NOR3_X1 U891 ( .A1(n1193), .A2(KEYINPUT40), .A3(G110), .ZN(n1249) );
AND2_X1 U892 ( .A1(G110), .A2(KEYINPUT40), .ZN(n1248) );
NAND2_X1 U893 ( .A1(n1226), .A2(G469), .ZN(n1242) );
NOR2_X1 U894 ( .A1(n1218), .A2(n1253), .ZN(G51) );
XOR2_X1 U895 ( .A(n1254), .B(n1255), .Z(n1253) );
XNOR2_X1 U896 ( .A(n1256), .B(n1257), .ZN(n1255) );
AND2_X1 U897 ( .A1(G210), .A2(n1226), .ZN(n1256) );
NOR2_X1 U898 ( .A1(n1258), .A2(n1109), .ZN(n1226) );
NOR2_X1 U899 ( .A1(n1195), .A2(n1200), .ZN(n1109) );
NAND4_X1 U900 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1200) );
AND2_X1 U901 ( .A1(n1263), .A2(n1264), .ZN(n1261) );
NAND3_X1 U902 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1260) );
NAND4_X1 U903 ( .A1(n1149), .A2(n1268), .A3(n1269), .A4(n1128), .ZN(n1266) );
NAND2_X1 U904 ( .A1(KEYINPUT49), .A2(n1270), .ZN(n1269) );
NAND2_X1 U905 ( .A1(n1101), .A2(n1103), .ZN(n1268) );
NAND2_X1 U906 ( .A1(n1104), .A2(n1271), .ZN(n1265) );
NAND3_X1 U907 ( .A1(n1272), .A2(n1273), .A3(n1270), .ZN(n1271) );
INV_X1 U908 ( .A(KEYINPUT49), .ZN(n1273) );
NAND2_X1 U909 ( .A1(n1149), .A2(n1274), .ZN(n1259) );
NAND2_X1 U910 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
XNOR2_X1 U911 ( .A(KEYINPUT63), .B(n1232), .ZN(n1276) );
NAND4_X1 U912 ( .A1(n1148), .A2(n1103), .A3(n1267), .A4(n1272), .ZN(n1232) );
XOR2_X1 U913 ( .A(n1277), .B(KEYINPUT38), .Z(n1275) );
NAND4_X1 U914 ( .A1(n1278), .A2(n1279), .A3(n1280), .A4(n1281), .ZN(n1195) );
NOR4_X1 U915 ( .A1(n1282), .A2(n1283), .A3(n1284), .A4(n1285), .ZN(n1281) );
INV_X1 U916 ( .A(n1286), .ZN(n1284) );
AND2_X1 U917 ( .A1(n1287), .A2(n1288), .ZN(n1280) );
NOR2_X1 U918 ( .A1(n1289), .A2(n1290), .ZN(n1254) );
NOR2_X1 U919 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XNOR2_X1 U920 ( .A(n1293), .B(KEYINPUT7), .ZN(n1292) );
AND2_X1 U921 ( .A1(n1293), .A2(n1291), .ZN(n1289) );
XOR2_X1 U922 ( .A(n1294), .B(n1295), .Z(n1291) );
NAND2_X1 U923 ( .A1(KEYINPUT2), .A2(n1296), .ZN(n1294) );
NOR2_X1 U924 ( .A1(n1152), .A2(G952), .ZN(n1218) );
XNOR2_X1 U925 ( .A(G146), .B(n1288), .ZN(G48) );
NAND4_X1 U926 ( .A1(n1297), .A2(n1148), .A3(n1138), .A4(n1298), .ZN(n1288) );
XNOR2_X1 U927 ( .A(G143), .B(n1287), .ZN(G45) );
NAND4_X1 U928 ( .A1(n1138), .A2(n1149), .A3(n1299), .A4(n1300), .ZN(n1287) );
AND3_X1 U929 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1300) );
XOR2_X1 U930 ( .A(n1278), .B(n1304), .Z(G42) );
XNOR2_X1 U931 ( .A(G140), .B(KEYINPUT18), .ZN(n1304) );
NAND4_X1 U932 ( .A1(n1148), .A2(n1305), .A3(n1306), .A4(n1307), .ZN(n1278) );
NAND3_X1 U933 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(G39) );
NAND2_X1 U934 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
OR3_X1 U935 ( .A1(n1312), .A2(n1311), .A3(KEYINPUT45), .ZN(n1309) );
NOR2_X1 U936 ( .A1(KEYINPUT0), .A2(n1279), .ZN(n1311) );
NAND2_X1 U937 ( .A1(KEYINPUT45), .A2(n1313), .ZN(n1308) );
NAND2_X1 U938 ( .A1(G137), .A2(n1279), .ZN(n1313) );
NAND3_X1 U939 ( .A1(n1298), .A2(n1305), .A3(n1314), .ZN(n1279) );
XNOR2_X1 U940 ( .A(n1315), .B(n1283), .ZN(G36) );
AND3_X1 U941 ( .A1(n1305), .A2(n1101), .A3(n1299), .ZN(n1283) );
XNOR2_X1 U942 ( .A(n1316), .B(n1282), .ZN(G33) );
AND3_X1 U943 ( .A1(n1299), .A2(n1305), .A3(n1148), .ZN(n1282) );
AND3_X1 U944 ( .A1(n1138), .A2(n1303), .A3(n1139), .ZN(n1305) );
INV_X1 U945 ( .A(n1119), .ZN(n1139) );
NAND3_X1 U946 ( .A1(n1132), .A2(n1176), .A3(n1317), .ZN(n1119) );
XNOR2_X1 U947 ( .A(n1267), .B(KEYINPUT59), .ZN(n1138) );
XOR2_X1 U948 ( .A(G128), .B(n1285), .Z(G30) );
AND4_X1 U949 ( .A1(n1298), .A2(n1297), .A3(n1101), .A4(n1267), .ZN(n1285) );
XNOR2_X1 U950 ( .A(G101), .B(n1318), .ZN(G3) );
NAND4_X1 U951 ( .A1(KEYINPUT43), .A2(n1270), .A3(n1267), .A4(n1319), .ZN(n1318) );
INV_X1 U952 ( .A(n1146), .ZN(n1270) );
NAND2_X1 U953 ( .A1(n1150), .A2(n1299), .ZN(n1146) );
XNOR2_X1 U954 ( .A(G125), .B(n1286), .ZN(G27) );
NAND4_X1 U955 ( .A1(n1297), .A2(n1148), .A3(n1141), .A4(n1306), .ZN(n1286) );
AND3_X1 U956 ( .A1(n1303), .A2(n1307), .A3(n1149), .ZN(n1297) );
NAND2_X1 U957 ( .A1(n1122), .A2(n1320), .ZN(n1303) );
NAND3_X1 U958 ( .A1(G902), .A2(n1321), .A3(n1186), .ZN(n1320) );
NOR2_X1 U959 ( .A1(n1152), .A2(G900), .ZN(n1186) );
XNOR2_X1 U960 ( .A(G122), .B(n1262), .ZN(G24) );
NAND4_X1 U961 ( .A1(n1322), .A2(n1103), .A3(n1301), .A4(n1302), .ZN(n1262) );
NOR2_X1 U962 ( .A1(n1307), .A2(n1298), .ZN(n1103) );
XNOR2_X1 U963 ( .A(G119), .B(n1264), .ZN(G21) );
NAND3_X1 U964 ( .A1(n1298), .A2(n1314), .A3(n1322), .ZN(n1264) );
INV_X1 U965 ( .A(n1306), .ZN(n1298) );
XNOR2_X1 U966 ( .A(G116), .B(n1263), .ZN(G18) );
NAND3_X1 U967 ( .A1(n1299), .A2(n1101), .A3(n1322), .ZN(n1263) );
NOR2_X1 U968 ( .A1(n1116), .A2(n1104), .ZN(n1322) );
AND2_X1 U969 ( .A1(n1323), .A2(n1301), .ZN(n1101) );
XOR2_X1 U970 ( .A(G113), .B(n1324), .Z(G15) );
NOR2_X1 U971 ( .A1(n1231), .A2(n1277), .ZN(n1324) );
NAND4_X1 U972 ( .A1(n1148), .A2(n1299), .A3(n1141), .A4(n1272), .ZN(n1277) );
INV_X1 U973 ( .A(n1116), .ZN(n1141) );
NAND2_X1 U974 ( .A1(n1325), .A2(n1134), .ZN(n1116) );
INV_X1 U975 ( .A(n1133), .ZN(n1325) );
NOR2_X1 U976 ( .A1(n1306), .A2(n1307), .ZN(n1299) );
NOR2_X1 U977 ( .A1(n1301), .A2(n1323), .ZN(n1148) );
XOR2_X1 U978 ( .A(n1326), .B(G110), .Z(G12) );
NAND2_X1 U979 ( .A1(KEYINPUT61), .A2(n1327), .ZN(n1326) );
NAND3_X1 U980 ( .A1(n1267), .A2(n1319), .A3(n1125), .ZN(n1327) );
INV_X1 U981 ( .A(n1128), .ZN(n1125) );
NAND2_X1 U982 ( .A1(n1314), .A2(n1306), .ZN(n1128) );
XOR2_X1 U983 ( .A(n1328), .B(n1173), .Z(n1306) );
INV_X1 U984 ( .A(n1171), .ZN(n1173) );
NOR2_X1 U985 ( .A1(n1236), .A2(G902), .ZN(n1171) );
XNOR2_X1 U986 ( .A(n1329), .B(n1330), .ZN(n1236) );
XOR2_X1 U987 ( .A(n1331), .B(n1332), .Z(n1330) );
XNOR2_X1 U988 ( .A(G101), .B(G113), .ZN(n1332) );
NAND2_X1 U989 ( .A1(KEYINPUT26), .A2(n1333), .ZN(n1331) );
XNOR2_X1 U990 ( .A(n1334), .B(G116), .ZN(n1333) );
XNOR2_X1 U991 ( .A(n1335), .B(n1241), .ZN(n1329) );
XOR2_X1 U992 ( .A(n1336), .B(n1295), .Z(n1335) );
NAND3_X1 U993 ( .A1(n1337), .A2(n1152), .A3(G210), .ZN(n1336) );
NAND2_X1 U994 ( .A1(KEYINPUT57), .A2(n1167), .ZN(n1328) );
INV_X1 U995 ( .A(G472), .ZN(n1167) );
AND2_X1 U996 ( .A1(n1150), .A2(n1307), .ZN(n1314) );
NAND3_X1 U997 ( .A1(n1338), .A2(n1339), .A3(n1177), .ZN(n1307) );
NAND2_X1 U998 ( .A1(n1160), .A2(n1161), .ZN(n1177) );
NAND2_X1 U999 ( .A1(n1161), .A2(n1340), .ZN(n1339) );
OR3_X1 U1000 ( .A1(n1161), .A2(n1160), .A3(n1340), .ZN(n1338) );
INV_X1 U1001 ( .A(KEYINPUT31), .ZN(n1340) );
NOR2_X1 U1002 ( .A1(n1221), .A2(G902), .ZN(n1160) );
XOR2_X1 U1003 ( .A(G119), .B(n1341), .Z(n1221) );
XOR2_X1 U1004 ( .A(n1342), .B(n1343), .Z(n1341) );
XOR2_X1 U1005 ( .A(n1344), .B(n1345), .Z(n1343) );
XOR2_X1 U1006 ( .A(G110), .B(n1346), .Z(n1345) );
AND2_X1 U1007 ( .A1(n1347), .A2(G221), .ZN(n1346) );
XOR2_X1 U1008 ( .A(n1348), .B(n1349), .Z(n1344) );
NOR2_X1 U1009 ( .A1(G128), .A2(KEYINPUT51), .ZN(n1349) );
NAND2_X1 U1010 ( .A1(KEYINPUT17), .A2(G140), .ZN(n1348) );
XOR2_X1 U1011 ( .A(n1350), .B(n1351), .Z(n1342) );
XOR2_X1 U1012 ( .A(KEYINPUT21), .B(G146), .Z(n1351) );
XNOR2_X1 U1013 ( .A(G137), .B(G125), .ZN(n1350) );
NAND2_X1 U1014 ( .A1(G217), .A2(n1352), .ZN(n1161) );
NOR2_X1 U1015 ( .A1(n1301), .A2(n1302), .ZN(n1150) );
INV_X1 U1016 ( .A(n1323), .ZN(n1302) );
NOR2_X1 U1017 ( .A1(n1353), .A2(n1175), .ZN(n1323) );
NOR2_X1 U1018 ( .A1(n1179), .A2(G475), .ZN(n1175) );
AND2_X1 U1019 ( .A1(G475), .A2(n1179), .ZN(n1353) );
NAND2_X1 U1020 ( .A1(n1229), .A2(n1258), .ZN(n1179) );
XOR2_X1 U1021 ( .A(n1354), .B(n1355), .Z(n1229) );
XOR2_X1 U1022 ( .A(n1356), .B(n1357), .Z(n1355) );
XOR2_X1 U1023 ( .A(n1358), .B(n1359), .Z(n1357) );
XNOR2_X1 U1024 ( .A(n1360), .B(n1361), .ZN(n1359) );
NOR2_X1 U1025 ( .A1(G140), .A2(KEYINPUT6), .ZN(n1361) );
NOR4_X1 U1026 ( .A1(KEYINPUT23), .A2(G953), .A3(G237), .A4(n1362), .ZN(n1360) );
INV_X1 U1027 ( .A(G214), .ZN(n1362) );
XNOR2_X1 U1028 ( .A(G104), .B(G113), .ZN(n1358) );
XOR2_X1 U1029 ( .A(n1363), .B(n1364), .Z(n1356) );
XNOR2_X1 U1030 ( .A(n1296), .B(G122), .ZN(n1364) );
XNOR2_X1 U1031 ( .A(G146), .B(n1316), .ZN(n1363) );
XNOR2_X1 U1032 ( .A(G143), .B(KEYINPUT44), .ZN(n1354) );
XOR2_X1 U1033 ( .A(n1165), .B(n1365), .Z(n1301) );
NOR2_X1 U1034 ( .A1(KEYINPUT1), .A2(n1366), .ZN(n1365) );
INV_X1 U1035 ( .A(G478), .ZN(n1366) );
AND2_X1 U1036 ( .A1(n1367), .A2(n1225), .ZN(n1165) );
XNOR2_X1 U1037 ( .A(n1368), .B(n1369), .ZN(n1225) );
NOR2_X1 U1038 ( .A1(KEYINPUT13), .A2(n1370), .ZN(n1369) );
XOR2_X1 U1039 ( .A(n1371), .B(n1372), .Z(n1370) );
XOR2_X1 U1040 ( .A(n1373), .B(n1374), .Z(n1372) );
NAND2_X1 U1041 ( .A1(n1375), .A2(n1376), .ZN(n1373) );
NAND2_X1 U1042 ( .A1(G116), .A2(n1377), .ZN(n1376) );
XOR2_X1 U1043 ( .A(KEYINPUT28), .B(n1378), .Z(n1375) );
NOR2_X1 U1044 ( .A1(G116), .A2(n1377), .ZN(n1378) );
XNOR2_X1 U1045 ( .A(n1315), .B(G107), .ZN(n1371) );
INV_X1 U1046 ( .A(G134), .ZN(n1315) );
NAND2_X1 U1047 ( .A1(G217), .A2(n1347), .ZN(n1368) );
AND2_X1 U1048 ( .A1(n1379), .A2(n1152), .ZN(n1347) );
XNOR2_X1 U1049 ( .A(G234), .B(KEYINPUT27), .ZN(n1379) );
XNOR2_X1 U1050 ( .A(KEYINPUT55), .B(n1258), .ZN(n1367) );
INV_X1 U1051 ( .A(n1104), .ZN(n1319) );
NAND2_X1 U1052 ( .A1(n1149), .A2(n1272), .ZN(n1104) );
NAND2_X1 U1053 ( .A1(n1122), .A2(n1380), .ZN(n1272) );
NAND4_X1 U1054 ( .A1(G953), .A2(G902), .A3(n1321), .A4(n1209), .ZN(n1380) );
INV_X1 U1055 ( .A(G898), .ZN(n1209) );
NAND3_X1 U1056 ( .A1(n1321), .A2(n1152), .A3(G952), .ZN(n1122) );
NAND2_X1 U1057 ( .A1(G237), .A2(n1381), .ZN(n1321) );
INV_X1 U1058 ( .A(n1231), .ZN(n1149) );
NAND2_X1 U1059 ( .A1(n1132), .A2(n1382), .ZN(n1231) );
NAND2_X1 U1060 ( .A1(n1317), .A2(n1176), .ZN(n1382) );
NAND2_X1 U1061 ( .A1(n1383), .A2(n1384), .ZN(n1176) );
INV_X1 U1062 ( .A(n1130), .ZN(n1317) );
NOR2_X1 U1063 ( .A1(n1384), .A2(n1383), .ZN(n1130) );
AND2_X1 U1064 ( .A1(n1385), .A2(n1258), .ZN(n1383) );
XOR2_X1 U1065 ( .A(n1386), .B(n1387), .Z(n1385) );
XNOR2_X1 U1066 ( .A(n1388), .B(n1295), .ZN(n1387) );
XNOR2_X1 U1067 ( .A(n1374), .B(n1389), .ZN(n1295) );
NOR2_X1 U1068 ( .A1(G146), .A2(KEYINPUT60), .ZN(n1389) );
XNOR2_X1 U1069 ( .A(G128), .B(G143), .ZN(n1374) );
NAND2_X1 U1070 ( .A1(KEYINPUT62), .A2(n1296), .ZN(n1388) );
INV_X1 U1071 ( .A(G125), .ZN(n1296) );
XNOR2_X1 U1072 ( .A(n1390), .B(n1391), .ZN(n1386) );
NOR2_X1 U1073 ( .A1(KEYINPUT25), .A2(n1257), .ZN(n1391) );
XOR2_X1 U1074 ( .A(n1392), .B(n1393), .Z(n1257) );
XNOR2_X1 U1075 ( .A(n1214), .B(n1210), .ZN(n1393) );
NAND2_X1 U1076 ( .A1(n1394), .A2(n1395), .ZN(n1210) );
NAND2_X1 U1077 ( .A1(G101), .A2(n1396), .ZN(n1395) );
NAND2_X1 U1078 ( .A1(n1397), .A2(n1398), .ZN(n1396) );
XNOR2_X1 U1079 ( .A(KEYINPUT41), .B(n1399), .ZN(n1397) );
NAND2_X1 U1080 ( .A1(n1400), .A2(n1401), .ZN(n1394) );
INV_X1 U1081 ( .A(G101), .ZN(n1401) );
NAND2_X1 U1082 ( .A1(n1402), .A2(n1403), .ZN(n1400) );
NAND2_X1 U1083 ( .A1(n1404), .A2(n1405), .ZN(n1403) );
OR2_X1 U1084 ( .A1(n1406), .A2(n1405), .ZN(n1402) );
INV_X1 U1085 ( .A(KEYINPUT41), .ZN(n1405) );
XOR2_X1 U1086 ( .A(G110), .B(n1407), .Z(n1214) );
XNOR2_X1 U1087 ( .A(KEYINPUT37), .B(n1377), .ZN(n1407) );
INV_X1 U1088 ( .A(G122), .ZN(n1377) );
XOR2_X1 U1089 ( .A(n1408), .B(KEYINPUT35), .Z(n1392) );
NAND2_X1 U1090 ( .A1(KEYINPUT34), .A2(n1212), .ZN(n1408) );
XOR2_X1 U1091 ( .A(n1409), .B(n1410), .Z(n1212) );
XNOR2_X1 U1092 ( .A(n1334), .B(G113), .ZN(n1410) );
INV_X1 U1093 ( .A(G119), .ZN(n1334) );
NAND2_X1 U1094 ( .A1(KEYINPUT30), .A2(G116), .ZN(n1409) );
NAND2_X1 U1095 ( .A1(KEYINPUT15), .A2(n1293), .ZN(n1390) );
NOR2_X1 U1096 ( .A1(n1205), .A2(G953), .ZN(n1293) );
INV_X1 U1097 ( .A(G224), .ZN(n1205) );
NAND2_X1 U1098 ( .A1(n1411), .A2(n1412), .ZN(n1384) );
XOR2_X1 U1099 ( .A(KEYINPUT8), .B(G210), .Z(n1411) );
NAND2_X1 U1100 ( .A1(G214), .A2(n1412), .ZN(n1132) );
NAND2_X1 U1101 ( .A1(n1337), .A2(n1258), .ZN(n1412) );
INV_X1 U1102 ( .A(G237), .ZN(n1337) );
INV_X1 U1103 ( .A(n1105), .ZN(n1267) );
NAND2_X1 U1104 ( .A1(n1133), .A2(n1134), .ZN(n1105) );
NAND2_X1 U1105 ( .A1(n1413), .A2(n1352), .ZN(n1134) );
NAND2_X1 U1106 ( .A1(n1381), .A2(n1258), .ZN(n1352) );
XOR2_X1 U1107 ( .A(G234), .B(KEYINPUT56), .Z(n1381) );
XOR2_X1 U1108 ( .A(KEYINPUT19), .B(G221), .Z(n1413) );
XNOR2_X1 U1109 ( .A(n1414), .B(G469), .ZN(n1133) );
NAND2_X1 U1110 ( .A1(n1415), .A2(n1258), .ZN(n1414) );
INV_X1 U1111 ( .A(G902), .ZN(n1258) );
XOR2_X1 U1112 ( .A(KEYINPUT32), .B(n1416), .Z(n1415) );
NOR2_X1 U1113 ( .A1(n1417), .A2(n1418), .ZN(n1416) );
XOR2_X1 U1114 ( .A(n1419), .B(KEYINPUT46), .Z(n1418) );
NAND2_X1 U1115 ( .A1(n1420), .A2(n1421), .ZN(n1419) );
NOR2_X1 U1116 ( .A1(n1420), .A2(n1421), .ZN(n1417) );
XNOR2_X1 U1117 ( .A(KEYINPUT16), .B(n1422), .ZN(n1421) );
NAND2_X1 U1118 ( .A1(n1423), .A2(n1424), .ZN(n1422) );
NAND2_X1 U1119 ( .A1(n1241), .A2(n1240), .ZN(n1424) );
XOR2_X1 U1120 ( .A(KEYINPUT47), .B(n1425), .Z(n1423) );
NOR2_X1 U1121 ( .A1(n1241), .A2(n1240), .ZN(n1425) );
XNOR2_X1 U1122 ( .A(n1189), .B(n1426), .ZN(n1240) );
XNOR2_X1 U1123 ( .A(G101), .B(n1406), .ZN(n1426) );
NAND2_X1 U1124 ( .A1(n1399), .A2(n1398), .ZN(n1406) );
NAND2_X1 U1125 ( .A1(G104), .A2(n1427), .ZN(n1398) );
INV_X1 U1126 ( .A(n1404), .ZN(n1399) );
NOR2_X1 U1127 ( .A1(n1427), .A2(G104), .ZN(n1404) );
INV_X1 U1128 ( .A(G107), .ZN(n1427) );
XOR2_X1 U1129 ( .A(n1428), .B(n1429), .Z(n1189) );
NOR2_X1 U1130 ( .A1(n1430), .A2(n1431), .ZN(n1429) );
XOR2_X1 U1131 ( .A(n1432), .B(KEYINPUT4), .Z(n1431) );
NAND2_X1 U1132 ( .A1(n1433), .A2(n1434), .ZN(n1432) );
XOR2_X1 U1133 ( .A(KEYINPUT24), .B(G146), .Z(n1433) );
NOR2_X1 U1134 ( .A1(G146), .A2(n1434), .ZN(n1430) );
XNOR2_X1 U1135 ( .A(KEYINPUT53), .B(n1435), .ZN(n1434) );
INV_X1 U1136 ( .A(G143), .ZN(n1435) );
XNOR2_X1 U1137 ( .A(G128), .B(KEYINPUT11), .ZN(n1428) );
XNOR2_X1 U1138 ( .A(n1190), .B(n1436), .ZN(n1241) );
NOR2_X1 U1139 ( .A1(KEYINPUT48), .A2(n1316), .ZN(n1436) );
INV_X1 U1140 ( .A(G131), .ZN(n1316) );
XNOR2_X1 U1141 ( .A(G134), .B(n1312), .ZN(n1190) );
INV_X1 U1142 ( .A(G137), .ZN(n1312) );
XNOR2_X1 U1143 ( .A(n1246), .B(n1437), .ZN(n1420) );
XNOR2_X1 U1144 ( .A(n1193), .B(G110), .ZN(n1437) );
INV_X1 U1145 ( .A(G140), .ZN(n1193) );
AND2_X1 U1146 ( .A1(G227), .A2(n1152), .ZN(n1246) );
INV_X1 U1147 ( .A(G953), .ZN(n1152) );
endmodule


