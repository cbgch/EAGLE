//Key = 0110010110001010100000101001011110001111001111101110010011001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360;

XOR2_X1 U746 ( .A(G107), .B(n1029), .Z(G9) );
NOR2_X1 U747 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U748 ( .A1(G953), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1031) );
NOR2_X1 U749 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR4_X1 U751 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1038) );
NOR3_X1 U752 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1040) );
NOR2_X1 U753 ( .A1(n1046), .A2(n1047), .ZN(n1039) );
NOR2_X1 U754 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U755 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR3_X1 U756 ( .A1(n1043), .A2(n1052), .A3(n1049), .ZN(n1037) );
INV_X1 U757 ( .A(n1053), .ZN(n1049) );
NOR2_X1 U758 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U759 ( .A1(n1056), .A2(n1042), .ZN(n1055) );
NOR3_X1 U760 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
NOR3_X1 U761 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
INV_X1 U762 ( .A(KEYINPUT8), .ZN(n1060) );
NOR2_X1 U763 ( .A1(KEYINPUT8), .A2(n1041), .ZN(n1058) );
NOR2_X1 U764 ( .A1(n1063), .A2(n1041), .ZN(n1054) );
NOR2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR3_X1 U766 ( .A1(n1032), .A2(G953), .A3(G952), .ZN(n1030) );
AND4_X1 U767 ( .A1(n1066), .A2(n1051), .A3(n1067), .A4(n1068), .ZN(n1032) );
NOR3_X1 U768 ( .A1(n1069), .A2(n1041), .A3(n1042), .ZN(n1068) );
XOR2_X1 U769 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND2_X1 U770 ( .A1(KEYINPUT49), .A2(G472), .ZN(n1071) );
XOR2_X1 U771 ( .A(KEYINPUT17), .B(n1072), .Z(n1066) );
NOR2_X1 U772 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XOR2_X1 U773 ( .A(n1075), .B(KEYINPUT38), .Z(n1074) );
XOR2_X1 U774 ( .A(n1076), .B(n1077), .Z(G72) );
NOR2_X1 U775 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XOR2_X1 U776 ( .A(n1080), .B(KEYINPUT33), .Z(n1079) );
AND2_X1 U777 ( .A1(G227), .A2(G900), .ZN(n1078) );
NAND2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1076) );
NAND2_X1 U779 ( .A1(n1083), .A2(n1080), .ZN(n1082) );
XOR2_X1 U780 ( .A(n1084), .B(n1085), .Z(n1083) );
NAND3_X1 U781 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1084) );
XOR2_X1 U782 ( .A(n1089), .B(KEYINPUT61), .Z(n1088) );
NAND3_X1 U783 ( .A1(G900), .A2(n1085), .A3(G953), .ZN(n1081) );
XNOR2_X1 U784 ( .A(n1090), .B(n1091), .ZN(n1085) );
NOR2_X1 U785 ( .A1(KEYINPUT20), .A2(n1092), .ZN(n1091) );
XOR2_X1 U786 ( .A(n1093), .B(n1094), .Z(n1092) );
XNOR2_X1 U787 ( .A(n1095), .B(n1096), .ZN(n1094) );
NAND2_X1 U788 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U789 ( .A1(n1099), .A2(G134), .ZN(n1098) );
XOR2_X1 U790 ( .A(n1100), .B(KEYINPUT18), .Z(n1097) );
NAND2_X1 U791 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U792 ( .A(n1103), .B(n1104), .Z(G69) );
XOR2_X1 U793 ( .A(n1105), .B(n1106), .Z(n1104) );
NAND2_X1 U794 ( .A1(G953), .A2(n1107), .ZN(n1106) );
NAND2_X1 U795 ( .A1(G898), .A2(G224), .ZN(n1107) );
NAND2_X1 U796 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
NAND2_X1 U797 ( .A1(G953), .A2(n1110), .ZN(n1109) );
XOR2_X1 U798 ( .A(n1111), .B(n1112), .Z(n1108) );
XNOR2_X1 U799 ( .A(n1113), .B(KEYINPUT2), .ZN(n1112) );
NAND2_X1 U800 ( .A1(n1114), .A2(KEYINPUT39), .ZN(n1113) );
XOR2_X1 U801 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U802 ( .A(n1117), .B(n1118), .Z(n1111) );
NOR2_X1 U803 ( .A1(n1119), .A2(G953), .ZN(n1103) );
NOR2_X1 U804 ( .A1(n1120), .A2(n1121), .ZN(G66) );
XNOR2_X1 U805 ( .A(n1122), .B(n1123), .ZN(n1121) );
NOR2_X1 U806 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NOR2_X1 U807 ( .A1(n1120), .A2(n1126), .ZN(G63) );
XOR2_X1 U808 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U809 ( .A1(n1129), .A2(n1125), .ZN(n1127) );
INV_X1 U810 ( .A(G478), .ZN(n1129) );
NOR2_X1 U811 ( .A1(n1120), .A2(n1130), .ZN(G60) );
XOR2_X1 U812 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U813 ( .A(KEYINPUT16), .B(n1133), .Z(n1132) );
NOR2_X1 U814 ( .A1(n1134), .A2(n1125), .ZN(n1133) );
INV_X1 U815 ( .A(G475), .ZN(n1134) );
XNOR2_X1 U816 ( .A(G104), .B(n1135), .ZN(G6) );
NOR2_X1 U817 ( .A1(n1120), .A2(n1136), .ZN(G57) );
NOR3_X1 U818 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
NOR2_X1 U819 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR2_X1 U820 ( .A1(KEYINPUT23), .A2(n1142), .ZN(n1140) );
XNOR2_X1 U821 ( .A(n1143), .B(KEYINPUT60), .ZN(n1142) );
NOR3_X1 U822 ( .A1(n1144), .A2(KEYINPUT23), .A3(n1143), .ZN(n1138) );
INV_X1 U823 ( .A(n1141), .ZN(n1144) );
XOR2_X1 U824 ( .A(n1145), .B(KEYINPUT43), .Z(n1141) );
AND2_X1 U825 ( .A1(n1143), .A2(KEYINPUT23), .ZN(n1137) );
XNOR2_X1 U826 ( .A(n1146), .B(n1147), .ZN(n1143) );
NOR2_X1 U827 ( .A1(n1148), .A2(n1125), .ZN(n1147) );
INV_X1 U828 ( .A(G472), .ZN(n1148) );
NAND2_X1 U829 ( .A1(KEYINPUT53), .A2(n1149), .ZN(n1146) );
XOR2_X1 U830 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U831 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U832 ( .A1(n1120), .A2(n1154), .ZN(G54) );
XOR2_X1 U833 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U834 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U835 ( .A(n1152), .B(n1159), .Z(n1158) );
NOR2_X1 U836 ( .A1(KEYINPUT58), .A2(n1160), .ZN(n1159) );
XOR2_X1 U837 ( .A(n1161), .B(n1162), .Z(n1155) );
XNOR2_X1 U838 ( .A(n1095), .B(n1163), .ZN(n1162) );
NAND2_X1 U839 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U840 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U841 ( .A(KEYINPUT45), .B(n1168), .Z(n1164) );
NOR2_X1 U842 ( .A1(n1166), .A2(n1167), .ZN(n1168) );
XNOR2_X1 U843 ( .A(KEYINPUT62), .B(G110), .ZN(n1166) );
NOR2_X1 U844 ( .A1(n1169), .A2(n1125), .ZN(n1161) );
NOR2_X1 U845 ( .A1(n1120), .A2(n1170), .ZN(G51) );
XOR2_X1 U846 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U847 ( .A(n1173), .B(n1174), .Z(n1171) );
NOR2_X1 U848 ( .A1(n1175), .A2(n1125), .ZN(n1174) );
NAND2_X1 U849 ( .A1(G902), .A2(n1034), .ZN(n1125) );
NAND4_X1 U850 ( .A1(n1119), .A2(n1086), .A3(n1176), .A4(n1177), .ZN(n1034) );
XNOR2_X1 U851 ( .A(KEYINPUT11), .B(n1089), .ZN(n1177) );
NAND3_X1 U852 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1089) );
NAND3_X1 U853 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
NAND2_X1 U854 ( .A1(n1184), .A2(n1185), .ZN(n1182) );
NAND2_X1 U855 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NAND2_X1 U856 ( .A1(KEYINPUT35), .A2(n1188), .ZN(n1184) );
NAND2_X1 U857 ( .A1(n1189), .A2(n1190), .ZN(n1181) );
INV_X1 U858 ( .A(n1187), .ZN(n1189) );
NAND2_X1 U859 ( .A1(n1191), .A2(n1192), .ZN(n1187) );
OR3_X1 U860 ( .A1(n1193), .A2(KEYINPUT35), .A3(n1042), .ZN(n1192) );
NAND2_X1 U861 ( .A1(n1194), .A2(n1195), .ZN(n1191) );
XOR2_X1 U862 ( .A(n1196), .B(KEYINPUT7), .Z(n1194) );
XNOR2_X1 U863 ( .A(KEYINPUT42), .B(n1087), .ZN(n1176) );
AND3_X1 U864 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1086) );
NAND2_X1 U865 ( .A1(n1057), .A2(n1200), .ZN(n1199) );
XOR2_X1 U866 ( .A(KEYINPUT26), .B(n1201), .Z(n1200) );
NAND3_X1 U867 ( .A1(n1044), .A2(n1064), .A3(n1183), .ZN(n1197) );
AND4_X1 U868 ( .A1(n1135), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1119) );
NOR4_X1 U869 ( .A1(n1205), .A2(n1206), .A3(n1029), .A4(n1207), .ZN(n1204) );
AND3_X1 U870 ( .A1(n1053), .A2(n1208), .A3(n1064), .ZN(n1029) );
NAND2_X1 U871 ( .A1(n1044), .A2(n1209), .ZN(n1203) );
NAND2_X1 U872 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND3_X1 U873 ( .A1(n1212), .A2(n1213), .A3(n1065), .ZN(n1211) );
XOR2_X1 U874 ( .A(KEYINPUT54), .B(n1046), .Z(n1213) );
NAND2_X1 U875 ( .A1(n1188), .A2(n1208), .ZN(n1210) );
NAND3_X1 U876 ( .A1(n1053), .A2(n1208), .A3(n1065), .ZN(n1135) );
INV_X1 U877 ( .A(n1214), .ZN(n1208) );
NOR2_X1 U878 ( .A1(n1080), .A2(G952), .ZN(n1120) );
XOR2_X1 U879 ( .A(n1215), .B(n1178), .Z(G48) );
NAND3_X1 U880 ( .A1(n1065), .A2(n1190), .A3(n1216), .ZN(n1178) );
XNOR2_X1 U881 ( .A(G143), .B(n1179), .ZN(G45) );
NAND4_X1 U882 ( .A1(n1216), .A2(n1044), .A3(n1217), .A4(n1218), .ZN(n1179) );
XOR2_X1 U883 ( .A(G140), .B(n1219), .Z(G42) );
NOR3_X1 U884 ( .A1(n1220), .A2(n1221), .A3(n1196), .ZN(n1219) );
XOR2_X1 U885 ( .A(G137), .B(n1222), .Z(G39) );
NOR2_X1 U886 ( .A1(n1223), .A2(n1220), .ZN(n1222) );
XOR2_X1 U887 ( .A(n1102), .B(n1224), .Z(G36) );
NAND4_X1 U888 ( .A1(KEYINPUT1), .A2(n1183), .A3(n1044), .A4(n1064), .ZN(n1224) );
XNOR2_X1 U889 ( .A(G131), .B(n1087), .ZN(G33) );
NAND3_X1 U890 ( .A1(n1065), .A2(n1044), .A3(n1183), .ZN(n1087) );
INV_X1 U891 ( .A(n1220), .ZN(n1183) );
NAND4_X1 U892 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1051), .ZN(n1220) );
INV_X1 U893 ( .A(n1041), .ZN(n1226) );
NAND2_X1 U894 ( .A1(n1228), .A2(n1062), .ZN(n1041) );
XOR2_X1 U895 ( .A(n1229), .B(n1198), .Z(G30) );
NAND3_X1 U896 ( .A1(n1190), .A2(n1064), .A3(n1216), .ZN(n1198) );
AND4_X1 U897 ( .A1(n1225), .A2(n1057), .A3(n1227), .A4(n1051), .ZN(n1216) );
XOR2_X1 U898 ( .A(G101), .B(n1230), .Z(G3) );
NOR3_X1 U899 ( .A1(n1231), .A2(n1232), .A3(n1214), .ZN(n1230) );
XOR2_X1 U900 ( .A(n1042), .B(KEYINPUT28), .Z(n1232) );
XOR2_X1 U901 ( .A(n1173), .B(n1233), .Z(G27) );
NAND2_X1 U902 ( .A1(n1201), .A2(n1057), .ZN(n1233) );
AND4_X1 U903 ( .A1(n1065), .A2(n1046), .A3(n1045), .A4(n1227), .ZN(n1201) );
NAND2_X1 U904 ( .A1(n1036), .A2(n1234), .ZN(n1227) );
NAND4_X1 U905 ( .A1(G902), .A2(G953), .A3(n1235), .A4(n1236), .ZN(n1234) );
INV_X1 U906 ( .A(G900), .ZN(n1236) );
INV_X1 U907 ( .A(n1221), .ZN(n1045) );
INV_X1 U908 ( .A(n1196), .ZN(n1065) );
XNOR2_X1 U909 ( .A(G122), .B(n1202), .ZN(G24) );
NAND4_X1 U910 ( .A1(n1237), .A2(n1053), .A3(n1217), .A4(n1218), .ZN(n1202) );
NOR2_X1 U911 ( .A1(n1238), .A2(n1239), .ZN(n1053) );
XOR2_X1 U912 ( .A(G119), .B(n1207), .Z(G21) );
NOR2_X1 U913 ( .A1(n1223), .A2(n1240), .ZN(n1207) );
NAND2_X1 U914 ( .A1(n1190), .A2(n1188), .ZN(n1223) );
AND2_X1 U915 ( .A1(n1186), .A2(n1239), .ZN(n1190) );
INV_X1 U916 ( .A(n1193), .ZN(n1239) );
XOR2_X1 U917 ( .A(G116), .B(n1206), .Z(G18) );
AND3_X1 U918 ( .A1(n1237), .A2(n1064), .A3(n1044), .ZN(n1206) );
NOR2_X1 U919 ( .A1(n1218), .A2(n1241), .ZN(n1064) );
INV_X1 U920 ( .A(n1240), .ZN(n1237) );
XNOR2_X1 U921 ( .A(G113), .B(n1242), .ZN(G15) );
NOR2_X1 U922 ( .A1(KEYINPUT15), .A2(n1243), .ZN(n1242) );
NOR3_X1 U923 ( .A1(n1196), .A2(n1240), .A3(n1231), .ZN(n1243) );
INV_X1 U924 ( .A(n1044), .ZN(n1231) );
NOR2_X1 U925 ( .A1(n1238), .A2(n1193), .ZN(n1044) );
NAND2_X1 U926 ( .A1(n1046), .A2(n1212), .ZN(n1240) );
INV_X1 U927 ( .A(n1043), .ZN(n1046) );
NAND2_X1 U928 ( .A1(n1050), .A2(n1051), .ZN(n1043) );
INV_X1 U929 ( .A(n1225), .ZN(n1050) );
NAND2_X1 U930 ( .A1(n1241), .A2(n1218), .ZN(n1196) );
XOR2_X1 U931 ( .A(G110), .B(n1205), .Z(G12) );
NOR3_X1 U932 ( .A1(n1042), .A2(n1214), .A3(n1221), .ZN(n1205) );
NAND2_X1 U933 ( .A1(n1195), .A2(n1186), .ZN(n1221) );
XNOR2_X1 U934 ( .A(n1238), .B(KEYINPUT56), .ZN(n1186) );
NAND2_X1 U935 ( .A1(n1244), .A2(n1075), .ZN(n1238) );
NAND2_X1 U936 ( .A1(n1245), .A2(n1246), .ZN(n1075) );
NAND2_X1 U937 ( .A1(n1122), .A2(n1247), .ZN(n1246) );
INV_X1 U938 ( .A(n1124), .ZN(n1245) );
XOR2_X1 U939 ( .A(KEYINPUT30), .B(n1073), .Z(n1244) );
AND3_X1 U940 ( .A1(n1122), .A2(n1247), .A3(n1124), .ZN(n1073) );
NAND2_X1 U941 ( .A1(G217), .A2(n1248), .ZN(n1124) );
NAND2_X1 U942 ( .A1(n1249), .A2(n1250), .ZN(n1122) );
NAND2_X1 U943 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XOR2_X1 U944 ( .A(KEYINPUT10), .B(n1253), .Z(n1251) );
NAND2_X1 U945 ( .A1(n1254), .A2(n1255), .ZN(n1249) );
XOR2_X1 U946 ( .A(KEYINPUT29), .B(n1252), .Z(n1255) );
XNOR2_X1 U947 ( .A(n1256), .B(n1257), .ZN(n1252) );
XOR2_X1 U948 ( .A(n1258), .B(n1259), .Z(n1257) );
NAND2_X1 U949 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND2_X1 U950 ( .A1(n1099), .A2(n1262), .ZN(n1261) );
XOR2_X1 U951 ( .A(KEYINPUT31), .B(n1263), .Z(n1260) );
NOR2_X1 U952 ( .A1(n1099), .A2(n1262), .ZN(n1263) );
NAND3_X1 U953 ( .A1(G221), .A2(G234), .A3(n1264), .ZN(n1262) );
XOR2_X1 U954 ( .A(n1080), .B(KEYINPUT9), .Z(n1264) );
NAND2_X1 U955 ( .A1(n1265), .A2(n1266), .ZN(n1258) );
OR2_X1 U956 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
XOR2_X1 U957 ( .A(n1269), .B(KEYINPUT52), .Z(n1265) );
NAND2_X1 U958 ( .A1(n1268), .A2(n1267), .ZN(n1269) );
INV_X1 U959 ( .A(G119), .ZN(n1267) );
XNOR2_X1 U960 ( .A(n1229), .B(KEYINPUT51), .ZN(n1268) );
NAND2_X1 U961 ( .A1(KEYINPUT37), .A2(G110), .ZN(n1256) );
XNOR2_X1 U962 ( .A(n1253), .B(KEYINPUT10), .ZN(n1254) );
XOR2_X1 U963 ( .A(n1193), .B(KEYINPUT40), .Z(n1195) );
XOR2_X1 U964 ( .A(n1070), .B(G472), .Z(n1193) );
NAND2_X1 U965 ( .A1(n1270), .A2(n1247), .ZN(n1070) );
XOR2_X1 U966 ( .A(n1271), .B(n1145), .Z(n1270) );
XOR2_X1 U967 ( .A(n1272), .B(G101), .Z(n1145) );
NAND2_X1 U968 ( .A1(G210), .A2(n1273), .ZN(n1272) );
NAND2_X1 U969 ( .A1(n1274), .A2(n1275), .ZN(n1271) );
NAND2_X1 U970 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XOR2_X1 U971 ( .A(KEYINPUT34), .B(n1278), .Z(n1277) );
XOR2_X1 U972 ( .A(KEYINPUT41), .B(n1279), .Z(n1276) );
XOR2_X1 U973 ( .A(KEYINPUT5), .B(n1280), .Z(n1274) );
NOR2_X1 U974 ( .A1(n1278), .A2(n1279), .ZN(n1280) );
XNOR2_X1 U975 ( .A(n1152), .B(n1281), .ZN(n1279) );
XOR2_X1 U976 ( .A(n1153), .B(n1116), .Z(n1278) );
NAND3_X1 U977 ( .A1(n1225), .A2(n1051), .A3(n1212), .ZN(n1214) );
AND2_X1 U978 ( .A1(n1057), .A2(n1282), .ZN(n1212) );
NAND2_X1 U979 ( .A1(n1036), .A2(n1283), .ZN(n1282) );
NAND4_X1 U980 ( .A1(G902), .A2(G953), .A3(n1235), .A4(n1110), .ZN(n1283) );
INV_X1 U981 ( .A(G898), .ZN(n1110) );
NAND3_X1 U982 ( .A1(n1235), .A2(n1080), .A3(G952), .ZN(n1036) );
NAND2_X1 U983 ( .A1(G237), .A2(G234), .ZN(n1235) );
AND2_X1 U984 ( .A1(n1061), .A2(n1062), .ZN(n1057) );
NAND2_X1 U985 ( .A1(G214), .A2(n1284), .ZN(n1062) );
INV_X1 U986 ( .A(n1228), .ZN(n1061) );
XNOR2_X1 U987 ( .A(n1285), .B(n1175), .ZN(n1228) );
NAND2_X1 U988 ( .A1(G210), .A2(n1284), .ZN(n1175) );
NAND2_X1 U989 ( .A1(n1286), .A2(n1247), .ZN(n1284) );
INV_X1 U990 ( .A(G237), .ZN(n1286) );
NAND2_X1 U991 ( .A1(n1287), .A2(n1247), .ZN(n1285) );
XOR2_X1 U992 ( .A(n1288), .B(n1172), .Z(n1287) );
XNOR2_X1 U993 ( .A(n1289), .B(n1290), .ZN(n1172) );
XOR2_X1 U994 ( .A(n1118), .B(n1291), .Z(n1290) );
INV_X1 U995 ( .A(n1150), .ZN(n1291) );
XNOR2_X1 U996 ( .A(n1281), .B(n1116), .ZN(n1150) );
XNOR2_X1 U997 ( .A(n1292), .B(n1293), .ZN(n1281) );
NOR2_X1 U998 ( .A1(KEYINPUT6), .A2(n1294), .ZN(n1293) );
XOR2_X1 U999 ( .A(KEYINPUT25), .B(G128), .Z(n1294) );
XOR2_X1 U1000 ( .A(n1215), .B(G143), .Z(n1292) );
XOR2_X1 U1001 ( .A(n1295), .B(n1296), .Z(n1118) );
INV_X1 U1002 ( .A(G101), .ZN(n1296) );
NAND2_X1 U1003 ( .A1(n1297), .A2(n1298), .ZN(n1295) );
OR2_X1 U1004 ( .A1(n1299), .A2(G104), .ZN(n1298) );
XOR2_X1 U1005 ( .A(n1300), .B(KEYINPUT4), .Z(n1297) );
NAND2_X1 U1006 ( .A1(G104), .A2(n1299), .ZN(n1300) );
XOR2_X1 U1007 ( .A(n1301), .B(n1302), .Z(n1289) );
XOR2_X1 U1008 ( .A(n1115), .B(n1303), .Z(n1302) );
NAND2_X1 U1009 ( .A1(G224), .A2(n1080), .ZN(n1303) );
NAND2_X1 U1010 ( .A1(KEYINPUT22), .A2(n1153), .ZN(n1115) );
XOR2_X1 U1011 ( .A(G116), .B(G119), .Z(n1153) );
NAND2_X1 U1012 ( .A1(KEYINPUT27), .A2(n1117), .ZN(n1301) );
XNOR2_X1 U1013 ( .A(G110), .B(n1304), .ZN(n1117) );
XOR2_X1 U1014 ( .A(KEYINPUT63), .B(G122), .Z(n1304) );
NAND2_X1 U1015 ( .A1(KEYINPUT36), .A2(n1173), .ZN(n1288) );
INV_X1 U1016 ( .A(G125), .ZN(n1173) );
NAND2_X1 U1017 ( .A1(n1305), .A2(n1248), .ZN(n1051) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1247), .ZN(n1248) );
XNOR2_X1 U1019 ( .A(G221), .B(KEYINPUT44), .ZN(n1305) );
XOR2_X1 U1020 ( .A(n1067), .B(KEYINPUT14), .Z(n1225) );
XOR2_X1 U1021 ( .A(n1169), .B(n1306), .Z(n1067) );
NOR2_X1 U1022 ( .A1(G902), .A2(n1307), .ZN(n1306) );
XOR2_X1 U1023 ( .A(n1308), .B(n1309), .Z(n1307) );
XNOR2_X1 U1024 ( .A(n1152), .B(n1160), .ZN(n1309) );
NAND2_X1 U1025 ( .A1(G227), .A2(n1080), .ZN(n1160) );
XNOR2_X1 U1026 ( .A(n1093), .B(n1310), .ZN(n1152) );
NOR2_X1 U1027 ( .A1(KEYINPUT3), .A2(n1311), .ZN(n1310) );
XOR2_X1 U1028 ( .A(n1102), .B(n1101), .Z(n1311) );
INV_X1 U1029 ( .A(n1099), .ZN(n1101) );
XNOR2_X1 U1030 ( .A(G137), .B(KEYINPUT13), .ZN(n1099) );
INV_X1 U1031 ( .A(G134), .ZN(n1102) );
XOR2_X1 U1032 ( .A(n1312), .B(n1313), .Z(n1308) );
NOR2_X1 U1033 ( .A1(KEYINPUT55), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1034 ( .A(n1315), .B(n1157), .Z(n1314) );
NAND2_X1 U1035 ( .A1(n1316), .A2(n1317), .ZN(n1157) );
NAND2_X1 U1036 ( .A1(n1318), .A2(n1299), .ZN(n1317) );
INV_X1 U1037 ( .A(G107), .ZN(n1299) );
NAND2_X1 U1038 ( .A1(n1319), .A2(G107), .ZN(n1316) );
XOR2_X1 U1039 ( .A(KEYINPUT57), .B(n1318), .Z(n1319) );
XOR2_X1 U1040 ( .A(G101), .B(G104), .Z(n1318) );
NAND2_X1 U1041 ( .A1(KEYINPUT48), .A2(n1095), .ZN(n1315) );
AND2_X1 U1042 ( .A1(n1320), .A2(n1321), .ZN(n1095) );
NAND2_X1 U1043 ( .A1(n1322), .A2(n1229), .ZN(n1321) );
XOR2_X1 U1044 ( .A(KEYINPUT50), .B(n1323), .Z(n1320) );
NOR2_X1 U1045 ( .A1(n1322), .A2(n1229), .ZN(n1323) );
INV_X1 U1046 ( .A(G128), .ZN(n1229) );
AND2_X1 U1047 ( .A1(n1324), .A2(n1325), .ZN(n1322) );
NAND2_X1 U1048 ( .A1(G143), .A2(n1215), .ZN(n1325) );
NAND2_X1 U1049 ( .A1(G146), .A2(n1326), .ZN(n1324) );
XNOR2_X1 U1050 ( .A(G143), .B(KEYINPUT0), .ZN(n1326) );
XOR2_X1 U1051 ( .A(n1167), .B(G110), .Z(n1312) );
INV_X1 U1052 ( .A(G469), .ZN(n1169) );
INV_X1 U1053 ( .A(n1188), .ZN(n1042) );
NOR2_X1 U1054 ( .A1(n1217), .A2(n1218), .ZN(n1188) );
XNOR2_X1 U1055 ( .A(n1327), .B(G475), .ZN(n1218) );
NAND2_X1 U1056 ( .A1(n1247), .A2(n1131), .ZN(n1327) );
NAND3_X1 U1057 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1131) );
NAND2_X1 U1058 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NAND2_X1 U1059 ( .A1(n1333), .A2(n1334), .ZN(n1329) );
INV_X1 U1060 ( .A(KEYINPUT32), .ZN(n1334) );
NAND2_X1 U1061 ( .A1(n1335), .A2(n1336), .ZN(n1333) );
INV_X1 U1062 ( .A(n1331), .ZN(n1336) );
XNOR2_X1 U1063 ( .A(KEYINPUT59), .B(n1332), .ZN(n1335) );
NAND2_X1 U1064 ( .A1(KEYINPUT32), .A2(n1337), .ZN(n1328) );
NAND2_X1 U1065 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
OR3_X1 U1066 ( .A1(n1331), .A2(n1332), .A3(KEYINPUT59), .ZN(n1339) );
XOR2_X1 U1067 ( .A(n1340), .B(n1253), .Z(n1331) );
XOR2_X1 U1068 ( .A(n1215), .B(n1090), .Z(n1253) );
XOR2_X1 U1069 ( .A(G125), .B(n1167), .Z(n1090) );
INV_X1 U1070 ( .A(G140), .ZN(n1167) );
INV_X1 U1071 ( .A(G146), .ZN(n1215) );
NAND3_X1 U1072 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1340) );
NAND2_X1 U1073 ( .A1(KEYINPUT21), .A2(n1344), .ZN(n1343) );
NAND3_X1 U1074 ( .A1(n1345), .A2(n1346), .A3(n1093), .ZN(n1342) );
INV_X1 U1075 ( .A(KEYINPUT21), .ZN(n1346) );
OR2_X1 U1076 ( .A1(n1093), .A2(n1345), .ZN(n1341) );
NOR2_X1 U1077 ( .A1(n1347), .A2(n1344), .ZN(n1345) );
XNOR2_X1 U1078 ( .A(n1348), .B(G143), .ZN(n1344) );
NAND2_X1 U1079 ( .A1(G214), .A2(n1273), .ZN(n1348) );
NOR2_X1 U1080 ( .A1(G953), .A2(G237), .ZN(n1273) );
INV_X1 U1081 ( .A(KEYINPUT12), .ZN(n1347) );
XOR2_X1 U1082 ( .A(G131), .B(KEYINPUT24), .Z(n1093) );
NAND2_X1 U1083 ( .A1(KEYINPUT59), .A2(n1332), .ZN(n1338) );
XNOR2_X1 U1084 ( .A(n1349), .B(n1116), .ZN(n1332) );
XOR2_X1 U1085 ( .A(G113), .B(KEYINPUT19), .Z(n1116) );
XNOR2_X1 U1086 ( .A(G104), .B(G122), .ZN(n1349) );
INV_X1 U1087 ( .A(G902), .ZN(n1247) );
INV_X1 U1088 ( .A(n1241), .ZN(n1217) );
XOR2_X1 U1089 ( .A(n1350), .B(G478), .Z(n1241) );
OR2_X1 U1090 ( .A1(n1128), .A2(G902), .ZN(n1350) );
XNOR2_X1 U1091 ( .A(n1351), .B(n1352), .ZN(n1128) );
XOR2_X1 U1092 ( .A(G107), .B(n1353), .Z(n1352) );
XOR2_X1 U1093 ( .A(G122), .B(G116), .Z(n1353) );
XOR2_X1 U1094 ( .A(n1354), .B(n1355), .Z(n1351) );
NOR2_X1 U1095 ( .A1(n1356), .A2(KEYINPUT47), .ZN(n1355) );
AND3_X1 U1096 ( .A1(G234), .A2(n1080), .A3(G217), .ZN(n1356) );
INV_X1 U1097 ( .A(G953), .ZN(n1080) );
NAND2_X1 U1098 ( .A1(n1357), .A2(n1358), .ZN(n1354) );
NAND2_X1 U1099 ( .A1(G134), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1100 ( .A(KEYINPUT46), .B(n1360), .Z(n1357) );
NOR2_X1 U1101 ( .A1(G134), .A2(n1359), .ZN(n1360) );
XOR2_X1 U1102 ( .A(G143), .B(G128), .Z(n1359) );
endmodule


