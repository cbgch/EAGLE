//Key = 1110011001000000010000100101000101010001000001011001000011000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337;

XNOR2_X1 U743 ( .A(n1018), .B(n1019), .ZN(G9) );
NOR3_X1 U744 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1019) );
XOR2_X1 U745 ( .A(KEYINPUT51), .B(n1023), .Z(n1020) );
NOR2_X1 U746 ( .A1(n1024), .A2(n1025), .ZN(G75) );
NOR3_X1 U747 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NAND3_X1 U748 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1026) );
NAND2_X1 U749 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U750 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND4_X1 U751 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
NAND4_X1 U752 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NAND2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U754 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
OR2_X1 U755 ( .A1(n1048), .A2(KEYINPUT49), .ZN(n1047) );
NAND3_X1 U756 ( .A1(KEYINPUT49), .A2(n1049), .A3(n1050), .ZN(n1042) );
NAND2_X1 U757 ( .A1(n1051), .A2(n1023), .ZN(n1040) );
NAND3_X1 U758 ( .A1(n1023), .A2(n1052), .A3(n1044), .ZN(n1034) );
NAND2_X1 U759 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U760 ( .A1(n1037), .A2(n1055), .ZN(n1054) );
XNOR2_X1 U761 ( .A(KEYINPUT4), .B(n1056), .ZN(n1055) );
NAND2_X1 U762 ( .A1(n1036), .A2(n1057), .ZN(n1053) );
NAND2_X1 U763 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U764 ( .A1(n1038), .A2(n1060), .ZN(n1059) );
NAND2_X1 U765 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U766 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U767 ( .A1(n1065), .A2(n1037), .ZN(n1058) );
INV_X1 U768 ( .A(n1066), .ZN(n1032) );
NOR3_X1 U769 ( .A1(n1067), .A2(G953), .A3(n1068), .ZN(n1024) );
INV_X1 U770 ( .A(n1029), .ZN(n1068) );
NAND2_X1 U771 ( .A1(n1069), .A2(n1070), .ZN(n1029) );
NOR4_X1 U772 ( .A1(n1065), .A2(n1063), .A3(n1071), .A4(n1072), .ZN(n1070) );
XOR2_X1 U773 ( .A(n1064), .B(KEYINPUT45), .Z(n1072) );
INV_X1 U774 ( .A(n1073), .ZN(n1071) );
INV_X1 U775 ( .A(n1074), .ZN(n1063) );
NOR4_X1 U776 ( .A1(n1075), .A2(n1076), .A3(n1050), .A4(n1077), .ZN(n1069) );
XNOR2_X1 U777 ( .A(KEYINPUT59), .B(n1078), .ZN(n1077) );
XNOR2_X1 U778 ( .A(KEYINPUT41), .B(n1027), .ZN(n1067) );
INV_X1 U779 ( .A(G952), .ZN(n1027) );
XOR2_X1 U780 ( .A(n1079), .B(n1080), .Z(G72) );
XOR2_X1 U781 ( .A(n1081), .B(n1082), .Z(n1080) );
NOR2_X1 U782 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U783 ( .A(n1085), .B(n1086), .Z(n1084) );
XOR2_X1 U784 ( .A(n1087), .B(n1088), .Z(n1086) );
XNOR2_X1 U785 ( .A(n1089), .B(n1090), .ZN(n1085) );
NOR2_X1 U786 ( .A1(G900), .A2(n1030), .ZN(n1083) );
NAND2_X1 U787 ( .A1(n1030), .A2(n1091), .ZN(n1081) );
NAND2_X1 U788 ( .A1(G953), .A2(n1092), .ZN(n1079) );
NAND2_X1 U789 ( .A1(G900), .A2(G227), .ZN(n1092) );
XOR2_X1 U790 ( .A(n1093), .B(n1094), .Z(G69) );
NOR2_X1 U791 ( .A1(n1095), .A2(n1030), .ZN(n1094) );
AND2_X1 U792 ( .A1(G224), .A2(G898), .ZN(n1095) );
NAND2_X1 U793 ( .A1(n1096), .A2(n1097), .ZN(n1093) );
NAND2_X1 U794 ( .A1(n1098), .A2(n1030), .ZN(n1097) );
XNOR2_X1 U795 ( .A(n1099), .B(n1100), .ZN(n1098) );
NAND3_X1 U796 ( .A1(G898), .A2(n1099), .A3(G953), .ZN(n1096) );
XNOR2_X1 U797 ( .A(n1101), .B(KEYINPUT30), .ZN(n1099) );
NOR2_X1 U798 ( .A1(n1102), .A2(n1103), .ZN(G66) );
XOR2_X1 U799 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U800 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NOR2_X1 U801 ( .A1(n1102), .A2(n1108), .ZN(G63) );
XOR2_X1 U802 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U803 ( .A1(n1111), .A2(KEYINPUT55), .ZN(n1110) );
NOR2_X1 U804 ( .A1(n1112), .A2(n1107), .ZN(n1111) );
NOR2_X1 U805 ( .A1(n1102), .A2(n1113), .ZN(G60) );
XOR2_X1 U806 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U807 ( .A(KEYINPUT0), .B(n1116), .Z(n1115) );
NOR2_X1 U808 ( .A1(n1117), .A2(n1107), .ZN(n1116) );
XNOR2_X1 U809 ( .A(n1118), .B(n1119), .ZN(G6) );
NOR2_X1 U810 ( .A1(n1022), .A2(n1041), .ZN(n1119) );
NOR2_X1 U811 ( .A1(n1102), .A2(n1120), .ZN(G57) );
XOR2_X1 U812 ( .A(n1121), .B(n1122), .Z(n1120) );
XNOR2_X1 U813 ( .A(n1123), .B(n1124), .ZN(n1122) );
XNOR2_X1 U814 ( .A(KEYINPUT19), .B(n1125), .ZN(n1121) );
NOR3_X1 U815 ( .A1(n1107), .A2(KEYINPUT11), .A3(n1126), .ZN(n1125) );
NOR2_X1 U816 ( .A1(n1102), .A2(n1127), .ZN(G54) );
XOR2_X1 U817 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U818 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U819 ( .A1(n1132), .A2(n1107), .ZN(n1131) );
NAND2_X1 U820 ( .A1(G902), .A2(n1028), .ZN(n1107) );
NOR2_X1 U821 ( .A1(KEYINPUT8), .A2(n1133), .ZN(n1130) );
XOR2_X1 U822 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U823 ( .A1(KEYINPUT14), .A2(n1136), .ZN(n1134) );
XNOR2_X1 U824 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR2_X1 U825 ( .A1(n1102), .A2(n1139), .ZN(G51) );
XOR2_X1 U826 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U827 ( .A(n1142), .B(n1101), .Z(n1141) );
NAND3_X1 U828 ( .A1(G902), .A2(G210), .A3(n1143), .ZN(n1142) );
XOR2_X1 U829 ( .A(n1028), .B(KEYINPUT36), .Z(n1143) );
NAND2_X1 U830 ( .A1(n1100), .A2(n1144), .ZN(n1028) );
INV_X1 U831 ( .A(n1091), .ZN(n1144) );
NAND4_X1 U832 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1091) );
NOR4_X1 U833 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1148) );
NOR2_X1 U834 ( .A1(n1153), .A2(n1154), .ZN(n1147) );
NOR2_X1 U835 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XNOR2_X1 U836 ( .A(n1157), .B(KEYINPUT48), .ZN(n1155) );
NOR3_X1 U837 ( .A1(n1158), .A2(n1050), .A3(n1159), .ZN(n1153) );
AND4_X1 U838 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1100) );
AND4_X1 U839 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1163) );
NOR2_X1 U840 ( .A1(n1168), .A2(n1169), .ZN(n1162) );
NOR3_X1 U841 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1169) );
XNOR2_X1 U842 ( .A(KEYINPUT22), .B(n1048), .ZN(n1170) );
NOR2_X1 U843 ( .A1(n1056), .A2(n1173), .ZN(n1168) );
NAND3_X1 U844 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1161) );
INV_X1 U845 ( .A(n1041), .ZN(n1176) );
NAND2_X1 U846 ( .A1(n1177), .A2(n1023), .ZN(n1041) );
NAND2_X1 U847 ( .A1(KEYINPUT5), .A2(n1022), .ZN(n1175) );
NAND2_X1 U848 ( .A1(n1178), .A2(n1179), .ZN(n1174) );
INV_X1 U849 ( .A(KEYINPUT5), .ZN(n1179) );
NAND2_X1 U850 ( .A1(n1180), .A2(n1181), .ZN(n1178) );
INV_X1 U851 ( .A(n1182), .ZN(n1180) );
NAND3_X1 U852 ( .A1(n1051), .A2(n1023), .A3(n1183), .ZN(n1160) );
XOR2_X1 U853 ( .A(n1184), .B(KEYINPUT15), .Z(n1140) );
NAND2_X1 U854 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND2_X1 U855 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U856 ( .A(n1189), .B(KEYINPUT26), .Z(n1187) );
XOR2_X1 U857 ( .A(n1190), .B(KEYINPUT29), .Z(n1185) );
OR2_X1 U858 ( .A1(n1188), .A2(n1189), .ZN(n1190) );
XOR2_X1 U859 ( .A(n1191), .B(n1192), .Z(n1188) );
NOR2_X1 U860 ( .A1(G125), .A2(KEYINPUT58), .ZN(n1192) );
NOR2_X1 U861 ( .A1(n1030), .A2(G952), .ZN(n1102) );
XNOR2_X1 U862 ( .A(G146), .B(n1145), .ZN(G48) );
NAND3_X1 U863 ( .A1(n1177), .A2(n1193), .A3(n1194), .ZN(n1145) );
XNOR2_X1 U864 ( .A(G143), .B(n1146), .ZN(G45) );
NAND4_X1 U865 ( .A1(n1194), .A2(n1049), .A3(n1195), .A4(n1196), .ZN(n1146) );
NOR3_X1 U866 ( .A1(n1056), .A2(n1157), .A3(n1061), .ZN(n1194) );
XOR2_X1 U867 ( .A(G140), .B(n1152), .Z(G42) );
NOR3_X1 U868 ( .A1(n1172), .A2(n1046), .A3(n1158), .ZN(n1152) );
NAND2_X1 U869 ( .A1(n1197), .A2(n1198), .ZN(G39) );
NAND2_X1 U870 ( .A1(G137), .A2(n1199), .ZN(n1198) );
XOR2_X1 U871 ( .A(KEYINPUT6), .B(n1200), .Z(n1197) );
NOR2_X1 U872 ( .A1(G137), .A2(n1199), .ZN(n1200) );
NAND3_X1 U873 ( .A1(n1193), .A2(n1201), .A3(n1202), .ZN(n1199) );
INV_X1 U874 ( .A(n1158), .ZN(n1202) );
XNOR2_X1 U875 ( .A(KEYINPUT60), .B(n1050), .ZN(n1201) );
XOR2_X1 U876 ( .A(G134), .B(n1151), .Z(G36) );
NOR3_X1 U877 ( .A1(n1048), .A2(n1021), .A3(n1158), .ZN(n1151) );
XNOR2_X1 U878 ( .A(n1203), .B(n1150), .ZN(G33) );
NOR3_X1 U879 ( .A1(n1172), .A2(n1048), .A3(n1158), .ZN(n1150) );
NAND4_X1 U880 ( .A1(n1036), .A2(n1204), .A3(n1038), .A4(n1205), .ZN(n1158) );
XOR2_X1 U881 ( .A(n1065), .B(KEYINPUT35), .Z(n1038) );
XOR2_X1 U882 ( .A(G128), .B(n1206), .Z(G30) );
NOR2_X1 U883 ( .A1(n1157), .A2(n1156), .ZN(n1206) );
NAND4_X1 U884 ( .A1(n1193), .A2(n1051), .A3(n1207), .A4(n1182), .ZN(n1156) );
INV_X1 U885 ( .A(n1159), .ZN(n1193) );
NAND2_X1 U886 ( .A1(n1208), .A2(n1209), .ZN(G3) );
NAND2_X1 U887 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
INV_X1 U888 ( .A(G101), .ZN(n1211) );
NAND2_X1 U889 ( .A1(n1212), .A2(G101), .ZN(n1208) );
NAND2_X1 U890 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND2_X1 U891 ( .A1(KEYINPUT44), .A2(n1215), .ZN(n1214) );
OR2_X1 U892 ( .A1(n1210), .A2(KEYINPUT44), .ZN(n1213) );
NOR2_X1 U893 ( .A1(KEYINPUT46), .A2(n1167), .ZN(n1210) );
INV_X1 U894 ( .A(n1215), .ZN(n1167) );
NOR3_X1 U895 ( .A1(n1050), .A2(n1022), .A3(n1048), .ZN(n1215) );
XNOR2_X1 U896 ( .A(n1149), .B(n1216), .ZN(G27) );
XOR2_X1 U897 ( .A(KEYINPUT61), .B(G125), .Z(n1216) );
AND4_X1 U898 ( .A1(n1177), .A2(n1037), .A3(n1217), .A4(n1218), .ZN(n1149) );
NOR2_X1 U899 ( .A1(n1157), .A2(n1056), .ZN(n1217) );
INV_X1 U900 ( .A(n1207), .ZN(n1056) );
INV_X1 U901 ( .A(n1205), .ZN(n1157) );
NAND2_X1 U902 ( .A1(n1066), .A2(n1219), .ZN(n1205) );
NAND4_X1 U903 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1221), .ZN(n1219) );
INV_X1 U904 ( .A(G900), .ZN(n1221) );
INV_X1 U905 ( .A(n1172), .ZN(n1177) );
XOR2_X1 U906 ( .A(n1166), .B(n1222), .Z(G24) );
XNOR2_X1 U907 ( .A(G122), .B(KEYINPUT3), .ZN(n1222) );
NAND4_X1 U908 ( .A1(n1223), .A2(n1023), .A3(n1195), .A4(n1196), .ZN(n1166) );
AND2_X1 U909 ( .A1(n1224), .A2(n1225), .ZN(n1023) );
INV_X1 U910 ( .A(n1171), .ZN(n1223) );
NAND3_X1 U911 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(G21) );
NAND2_X1 U912 ( .A1(G119), .A2(n1165), .ZN(n1228) );
NAND2_X1 U913 ( .A1(KEYINPUT28), .A2(n1229), .ZN(n1227) );
NAND2_X1 U914 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XNOR2_X1 U915 ( .A(KEYINPUT32), .B(G119), .ZN(n1230) );
NAND2_X1 U916 ( .A1(n1232), .A2(n1233), .ZN(n1226) );
INV_X1 U917 ( .A(KEYINPUT28), .ZN(n1233) );
NAND2_X1 U918 ( .A1(n1234), .A2(n1235), .ZN(n1232) );
OR3_X1 U919 ( .A1(n1165), .A2(G119), .A3(KEYINPUT32), .ZN(n1235) );
INV_X1 U920 ( .A(n1231), .ZN(n1165) );
NOR3_X1 U921 ( .A1(n1159), .A2(n1050), .A3(n1171), .ZN(n1231) );
NAND2_X1 U922 ( .A1(n1236), .A2(n1075), .ZN(n1159) );
XNOR2_X1 U923 ( .A(KEYINPUT43), .B(n1224), .ZN(n1236) );
NAND2_X1 U924 ( .A1(KEYINPUT32), .A2(G119), .ZN(n1234) );
XNOR2_X1 U925 ( .A(G116), .B(n1237), .ZN(G18) );
NAND3_X1 U926 ( .A1(n1238), .A2(n1239), .A3(n1207), .ZN(n1237) );
XOR2_X1 U927 ( .A(KEYINPUT16), .B(KEYINPUT1), .Z(n1239) );
XNOR2_X1 U928 ( .A(KEYINPUT42), .B(n1173), .ZN(n1238) );
NAND4_X1 U929 ( .A1(n1049), .A2(n1037), .A3(n1051), .A4(n1240), .ZN(n1173) );
INV_X1 U930 ( .A(n1021), .ZN(n1051) );
NAND2_X1 U931 ( .A1(n1241), .A2(n1242), .ZN(n1021) );
XNOR2_X1 U932 ( .A(n1195), .B(KEYINPUT47), .ZN(n1241) );
XNOR2_X1 U933 ( .A(n1243), .B(KEYINPUT38), .ZN(n1195) );
INV_X1 U934 ( .A(n1048), .ZN(n1049) );
XNOR2_X1 U935 ( .A(G113), .B(n1244), .ZN(G15) );
NOR2_X1 U936 ( .A1(n1245), .A2(KEYINPUT21), .ZN(n1244) );
NOR3_X1 U937 ( .A1(n1172), .A2(n1171), .A3(n1048), .ZN(n1245) );
NAND2_X1 U938 ( .A1(n1224), .A2(n1075), .ZN(n1048) );
INV_X1 U939 ( .A(n1076), .ZN(n1224) );
NAND2_X1 U940 ( .A1(n1037), .A2(n1181), .ZN(n1171) );
AND2_X1 U941 ( .A1(n1064), .A2(n1074), .ZN(n1037) );
NAND2_X1 U942 ( .A1(n1243), .A2(n1196), .ZN(n1172) );
XOR2_X1 U943 ( .A(n1164), .B(n1246), .Z(G12) );
NOR2_X1 U944 ( .A1(G110), .A2(KEYINPUT7), .ZN(n1246) );
NAND3_X1 U945 ( .A1(n1044), .A2(n1183), .A3(n1218), .ZN(n1164) );
INV_X1 U946 ( .A(n1046), .ZN(n1218) );
NAND2_X1 U947 ( .A1(n1076), .A2(n1225), .ZN(n1046) );
XOR2_X1 U948 ( .A(n1075), .B(KEYINPUT39), .Z(n1225) );
XOR2_X1 U949 ( .A(n1247), .B(n1126), .Z(n1075) );
INV_X1 U950 ( .A(G472), .ZN(n1126) );
NAND2_X1 U951 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
XOR2_X1 U952 ( .A(n1250), .B(n1123), .Z(n1248) );
XNOR2_X1 U953 ( .A(n1251), .B(G101), .ZN(n1123) );
NAND3_X1 U954 ( .A1(n1252), .A2(n1030), .A3(G210), .ZN(n1251) );
NOR2_X1 U955 ( .A1(KEYINPUT54), .A2(n1124), .ZN(n1250) );
XOR2_X1 U956 ( .A(n1253), .B(n1254), .Z(n1124) );
XNOR2_X1 U957 ( .A(n1135), .B(n1255), .ZN(n1254) );
NAND2_X1 U958 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND2_X1 U959 ( .A1(KEYINPUT33), .A2(n1258), .ZN(n1257) );
XNOR2_X1 U960 ( .A(G116), .B(G119), .ZN(n1258) );
NAND3_X1 U961 ( .A1(G116), .A2(n1259), .A3(n1260), .ZN(n1256) );
INV_X1 U962 ( .A(KEYINPUT33), .ZN(n1260) );
XNOR2_X1 U963 ( .A(n1191), .B(G113), .ZN(n1253) );
INV_X1 U964 ( .A(n1261), .ZN(n1191) );
XOR2_X1 U965 ( .A(n1262), .B(n1106), .Z(n1076) );
NAND2_X1 U966 ( .A1(G217), .A2(n1263), .ZN(n1106) );
OR2_X1 U967 ( .A1(n1105), .A2(G902), .ZN(n1262) );
XNOR2_X1 U968 ( .A(n1264), .B(n1265), .ZN(n1105) );
XNOR2_X1 U969 ( .A(n1266), .B(n1267), .ZN(n1265) );
XOR2_X1 U970 ( .A(n1268), .B(n1269), .Z(n1264) );
XNOR2_X1 U971 ( .A(G110), .B(n1270), .ZN(n1269) );
NAND2_X1 U972 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND2_X1 U973 ( .A1(KEYINPUT23), .A2(G137), .ZN(n1272) );
XOR2_X1 U974 ( .A(n1273), .B(n1274), .Z(n1271) );
NOR2_X1 U975 ( .A1(G137), .A2(KEYINPUT23), .ZN(n1274) );
NAND2_X1 U976 ( .A1(n1275), .A2(G221), .ZN(n1273) );
NAND2_X1 U977 ( .A1(KEYINPUT57), .A2(G119), .ZN(n1268) );
INV_X1 U978 ( .A(n1022), .ZN(n1183) );
NAND2_X1 U979 ( .A1(n1181), .A2(n1182), .ZN(n1022) );
XOR2_X1 U980 ( .A(n1204), .B(KEYINPUT34), .Z(n1182) );
INV_X1 U981 ( .A(n1061), .ZN(n1204) );
NAND2_X1 U982 ( .A1(n1276), .A2(n1074), .ZN(n1061) );
NAND2_X1 U983 ( .A1(G221), .A2(n1263), .ZN(n1074) );
NAND2_X1 U984 ( .A1(G234), .A2(n1249), .ZN(n1263) );
XOR2_X1 U985 ( .A(n1064), .B(KEYINPUT31), .Z(n1276) );
XNOR2_X1 U986 ( .A(n1277), .B(n1132), .ZN(n1064) );
INV_X1 U987 ( .A(G469), .ZN(n1132) );
NAND2_X1 U988 ( .A1(n1278), .A2(n1249), .ZN(n1277) );
XOR2_X1 U989 ( .A(n1279), .B(n1128), .Z(n1278) );
XNOR2_X1 U990 ( .A(n1280), .B(n1281), .ZN(n1128) );
XOR2_X1 U991 ( .A(G140), .B(G110), .Z(n1281) );
NAND2_X1 U992 ( .A1(G227), .A2(n1030), .ZN(n1280) );
XNOR2_X1 U993 ( .A(n1135), .B(n1282), .ZN(n1279) );
NOR2_X1 U994 ( .A1(KEYINPUT13), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U995 ( .A(n1137), .B(n1284), .ZN(n1283) );
NOR2_X1 U996 ( .A1(KEYINPUT62), .A2(n1138), .ZN(n1284) );
XNOR2_X1 U997 ( .A(n1285), .B(n1286), .ZN(n1138) );
NOR2_X1 U998 ( .A1(G101), .A2(KEYINPUT40), .ZN(n1286) );
XNOR2_X1 U999 ( .A(G146), .B(n1287), .ZN(n1137) );
INV_X1 U1000 ( .A(n1089), .ZN(n1287) );
XOR2_X1 U1001 ( .A(n1087), .B(n1288), .Z(n1135) );
NOR2_X1 U1002 ( .A1(KEYINPUT24), .A2(n1088), .ZN(n1288) );
XNOR2_X1 U1003 ( .A(n1203), .B(KEYINPUT18), .ZN(n1088) );
XOR2_X1 U1004 ( .A(G134), .B(G137), .Z(n1087) );
AND2_X1 U1005 ( .A1(n1207), .A2(n1240), .ZN(n1181) );
NAND2_X1 U1006 ( .A1(n1066), .A2(n1289), .ZN(n1240) );
NAND4_X1 U1007 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1290), .ZN(n1289) );
INV_X1 U1008 ( .A(G898), .ZN(n1290) );
NAND3_X1 U1009 ( .A1(n1220), .A2(n1030), .A3(G952), .ZN(n1066) );
NAND2_X1 U1010 ( .A1(G234), .A2(G237), .ZN(n1220) );
NOR2_X1 U1011 ( .A1(n1065), .A2(n1036), .ZN(n1207) );
AND2_X1 U1012 ( .A1(n1291), .A2(n1073), .ZN(n1036) );
NAND2_X1 U1013 ( .A1(G210), .A2(n1292), .ZN(n1073) );
NAND2_X1 U1014 ( .A1(n1293), .A2(n1249), .ZN(n1292) );
OR2_X1 U1015 ( .A1(n1252), .A2(n1294), .ZN(n1293) );
XOR2_X1 U1016 ( .A(n1078), .B(KEYINPUT63), .Z(n1291) );
NAND3_X1 U1017 ( .A1(n1295), .A2(n1249), .A3(n1294), .ZN(n1078) );
XNOR2_X1 U1018 ( .A(n1296), .B(n1297), .ZN(n1294) );
XNOR2_X1 U1019 ( .A(G125), .B(n1189), .ZN(n1297) );
NAND2_X1 U1020 ( .A1(G224), .A2(n1030), .ZN(n1189) );
XNOR2_X1 U1021 ( .A(n1101), .B(n1261), .ZN(n1296) );
NAND3_X1 U1022 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1261) );
NAND2_X1 U1023 ( .A1(KEYINPUT52), .A2(n1301), .ZN(n1300) );
NAND3_X1 U1024 ( .A1(n1302), .A2(n1303), .A3(n1266), .ZN(n1299) );
INV_X1 U1025 ( .A(KEYINPUT52), .ZN(n1303) );
OR2_X1 U1026 ( .A1(n1266), .A2(n1302), .ZN(n1298) );
NOR2_X1 U1027 ( .A1(KEYINPUT12), .A2(n1301), .ZN(n1302) );
XOR2_X1 U1028 ( .A(G146), .B(n1304), .Z(n1301) );
NOR2_X1 U1029 ( .A1(G143), .A2(KEYINPUT10), .ZN(n1304) );
XOR2_X1 U1030 ( .A(n1305), .B(n1306), .Z(n1101) );
XNOR2_X1 U1031 ( .A(n1307), .B(n1308), .ZN(n1306) );
XNOR2_X1 U1032 ( .A(KEYINPUT25), .B(n1259), .ZN(n1308) );
INV_X1 U1033 ( .A(G119), .ZN(n1259) );
INV_X1 U1034 ( .A(G113), .ZN(n1307) );
XNOR2_X1 U1035 ( .A(n1309), .B(n1310), .ZN(n1305) );
XNOR2_X1 U1036 ( .A(G110), .B(n1311), .ZN(n1310) );
NAND2_X1 U1037 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NAND2_X1 U1038 ( .A1(G101), .A2(n1285), .ZN(n1313) );
XOR2_X1 U1039 ( .A(n1314), .B(KEYINPUT20), .Z(n1312) );
OR2_X1 U1040 ( .A1(n1285), .A2(G101), .ZN(n1314) );
XOR2_X1 U1041 ( .A(G107), .B(G104), .Z(n1285) );
NAND2_X1 U1042 ( .A1(G210), .A2(G237), .ZN(n1295) );
AND2_X1 U1043 ( .A1(G214), .A2(n1315), .ZN(n1065) );
NAND2_X1 U1044 ( .A1(n1249), .A2(n1252), .ZN(n1315) );
INV_X1 U1045 ( .A(n1050), .ZN(n1044) );
NAND2_X1 U1046 ( .A1(n1242), .A2(n1243), .ZN(n1050) );
XNOR2_X1 U1047 ( .A(n1316), .B(n1112), .ZN(n1243) );
INV_X1 U1048 ( .A(G478), .ZN(n1112) );
NAND2_X1 U1049 ( .A1(n1109), .A2(n1249), .ZN(n1316) );
XOR2_X1 U1050 ( .A(n1317), .B(n1318), .Z(n1109) );
XNOR2_X1 U1051 ( .A(n1018), .B(n1319), .ZN(n1318) );
XOR2_X1 U1052 ( .A(KEYINPUT53), .B(G134), .Z(n1319) );
INV_X1 U1053 ( .A(G107), .ZN(n1018) );
XOR2_X1 U1054 ( .A(n1320), .B(n1309), .Z(n1317) );
XOR2_X1 U1055 ( .A(G116), .B(G122), .Z(n1309) );
XNOR2_X1 U1056 ( .A(n1089), .B(n1321), .ZN(n1320) );
AND2_X1 U1057 ( .A1(n1275), .A2(G217), .ZN(n1321) );
AND2_X1 U1058 ( .A1(n1322), .A2(n1030), .ZN(n1275) );
XNOR2_X1 U1059 ( .A(G234), .B(KEYINPUT9), .ZN(n1322) );
XOR2_X1 U1060 ( .A(G143), .B(n1266), .Z(n1089) );
XOR2_X1 U1061 ( .A(G128), .B(KEYINPUT2), .Z(n1266) );
INV_X1 U1062 ( .A(n1196), .ZN(n1242) );
XOR2_X1 U1063 ( .A(n1323), .B(n1117), .Z(n1196) );
INV_X1 U1064 ( .A(G475), .ZN(n1117) );
NAND2_X1 U1065 ( .A1(n1114), .A2(n1249), .ZN(n1323) );
INV_X1 U1066 ( .A(G902), .ZN(n1249) );
XOR2_X1 U1067 ( .A(n1324), .B(n1325), .Z(n1114) );
XOR2_X1 U1068 ( .A(n1326), .B(n1327), .Z(n1325) );
XNOR2_X1 U1069 ( .A(n1328), .B(n1329), .ZN(n1327) );
INV_X1 U1070 ( .A(G143), .ZN(n1329) );
NAND2_X1 U1071 ( .A1(KEYINPUT27), .A2(n1203), .ZN(n1328) );
INV_X1 U1072 ( .A(G131), .ZN(n1203) );
NAND2_X1 U1073 ( .A1(KEYINPUT56), .A2(n1267), .ZN(n1326) );
XNOR2_X1 U1074 ( .A(n1090), .B(KEYINPUT50), .ZN(n1267) );
XOR2_X1 U1075 ( .A(G125), .B(n1330), .Z(n1090) );
XOR2_X1 U1076 ( .A(G146), .B(G140), .Z(n1330) );
XOR2_X1 U1077 ( .A(n1331), .B(n1332), .Z(n1324) );
NOR2_X1 U1078 ( .A1(KEYINPUT37), .A2(n1333), .ZN(n1332) );
AND3_X1 U1079 ( .A1(G214), .A2(n1030), .A3(n1252), .ZN(n1333) );
INV_X1 U1080 ( .A(G237), .ZN(n1252) );
INV_X1 U1081 ( .A(G953), .ZN(n1030) );
NAND2_X1 U1082 ( .A1(n1334), .A2(n1335), .ZN(n1331) );
NAND2_X1 U1083 ( .A1(n1336), .A2(n1118), .ZN(n1335) );
XOR2_X1 U1084 ( .A(KEYINPUT17), .B(n1337), .Z(n1334) );
NOR2_X1 U1085 ( .A1(n1336), .A2(n1118), .ZN(n1337) );
INV_X1 U1086 ( .A(G104), .ZN(n1118) );
XNOR2_X1 U1087 ( .A(G113), .B(G122), .ZN(n1336) );
endmodule


