//Key = 0110101000101111010010010010111110111110101001111110001000100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352;

XNOR2_X1 U760 ( .A(G107), .B(n1048), .ZN(G9) );
NOR2_X1 U761 ( .A1(n1049), .A2(n1050), .ZN(G75) );
NOR4_X1 U762 ( .A1(G953), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1050) );
NOR2_X1 U763 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U764 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR3_X1 U765 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
NOR2_X1 U766 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR2_X1 U767 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U768 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NOR2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U770 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
NOR2_X1 U771 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR2_X1 U772 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U773 ( .A1(n1075), .A2(n1070), .ZN(n1061) );
NOR2_X1 U774 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR3_X1 U775 ( .A1(n1068), .A2(n1078), .A3(n1079), .ZN(n1076) );
NOR4_X1 U776 ( .A1(n1080), .A2(n1070), .A3(n1068), .A4(n1064), .ZN(n1056) );
INV_X1 U777 ( .A(n1081), .ZN(n1070) );
NOR2_X1 U778 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NOR3_X1 U779 ( .A1(n1051), .A2(G953), .A3(G952), .ZN(n1049) );
AND4_X1 U780 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1051) );
NOR4_X1 U781 ( .A1(n1058), .A2(n1079), .A3(n1068), .A4(n1088), .ZN(n1087) );
XOR2_X1 U782 ( .A(KEYINPUT55), .B(n1089), .Z(n1088) );
NOR2_X1 U783 ( .A1(G472), .A2(n1090), .ZN(n1089) );
AND3_X1 U784 ( .A1(n1091), .A2(n1078), .A3(n1092), .ZN(n1086) );
OR2_X1 U785 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NAND2_X1 U786 ( .A1(G472), .A2(n1090), .ZN(n1085) );
XOR2_X1 U787 ( .A(G478), .B(n1095), .Z(n1084) );
NOR2_X1 U788 ( .A1(n1096), .A2(KEYINPUT8), .ZN(n1095) );
XOR2_X1 U789 ( .A(n1097), .B(n1098), .Z(G72) );
NOR2_X1 U790 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U791 ( .A(n1101), .B(n1102), .Z(n1100) );
XOR2_X1 U792 ( .A(n1103), .B(n1104), .Z(n1102) );
XOR2_X1 U793 ( .A(n1105), .B(n1106), .Z(n1101) );
NAND2_X1 U794 ( .A1(KEYINPUT30), .A2(n1107), .ZN(n1106) );
NOR2_X1 U795 ( .A1(G900), .A2(n1108), .ZN(n1099) );
NAND3_X1 U796 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1097) );
NAND2_X1 U797 ( .A1(G953), .A2(n1112), .ZN(n1109) );
NAND2_X1 U798 ( .A1(G900), .A2(G227), .ZN(n1112) );
XOR2_X1 U799 ( .A(n1113), .B(n1114), .Z(G69) );
NOR2_X1 U800 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U801 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U802 ( .A(n1119), .B(KEYINPUT11), .Z(n1118) );
NAND2_X1 U803 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U804 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XNOR2_X1 U805 ( .A(n1124), .B(KEYINPUT19), .ZN(n1120) );
NOR2_X1 U806 ( .A1(G898), .A2(n1108), .ZN(n1115) );
NAND2_X1 U807 ( .A1(n1125), .A2(n1126), .ZN(n1113) );
NAND2_X1 U808 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND3_X1 U809 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1127) );
XOR2_X1 U810 ( .A(KEYINPUT62), .B(n1132), .Z(n1130) );
XOR2_X1 U811 ( .A(KEYINPUT15), .B(n1133), .Z(n1129) );
NAND3_X1 U812 ( .A1(KEYINPUT48), .A2(n1134), .A3(G953), .ZN(n1125) );
NAND2_X1 U813 ( .A1(G898), .A2(G224), .ZN(n1134) );
NOR2_X1 U814 ( .A1(n1135), .A2(n1136), .ZN(G66) );
XOR2_X1 U815 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U816 ( .A1(n1094), .A2(n1139), .ZN(n1138) );
NOR2_X1 U817 ( .A1(n1135), .A2(n1140), .ZN(G63) );
NOR3_X1 U818 ( .A1(n1096), .A2(n1141), .A3(n1142), .ZN(n1140) );
NOR3_X1 U819 ( .A1(n1143), .A2(n1144), .A3(n1139), .ZN(n1142) );
INV_X1 U820 ( .A(n1145), .ZN(n1143) );
NOR2_X1 U821 ( .A1(n1146), .A2(n1145), .ZN(n1141) );
AND2_X1 U822 ( .A1(n1053), .A2(G478), .ZN(n1146) );
NOR2_X1 U823 ( .A1(n1135), .A2(n1147), .ZN(G60) );
XOR2_X1 U824 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U825 ( .A(KEYINPUT26), .B(n1150), .Z(n1149) );
NOR2_X1 U826 ( .A1(n1151), .A2(n1139), .ZN(n1150) );
XNOR2_X1 U827 ( .A(G475), .B(KEYINPUT24), .ZN(n1151) );
XOR2_X1 U828 ( .A(n1133), .B(n1152), .Z(G6) );
NOR2_X1 U829 ( .A1(KEYINPUT16), .A2(n1153), .ZN(n1152) );
NOR2_X1 U830 ( .A1(n1135), .A2(n1154), .ZN(G57) );
XOR2_X1 U831 ( .A(n1155), .B(n1156), .Z(n1154) );
XNOR2_X1 U832 ( .A(n1157), .B(n1158), .ZN(n1156) );
XOR2_X1 U833 ( .A(n1159), .B(n1160), .Z(n1155) );
NOR2_X1 U834 ( .A1(n1161), .A2(n1139), .ZN(n1160) );
INV_X1 U835 ( .A(G472), .ZN(n1161) );
NAND2_X1 U836 ( .A1(KEYINPUT4), .A2(n1162), .ZN(n1159) );
NOR2_X1 U837 ( .A1(n1135), .A2(n1163), .ZN(G54) );
XOR2_X1 U838 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U839 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U840 ( .A1(KEYINPUT0), .A2(n1105), .ZN(n1166) );
XOR2_X1 U841 ( .A(n1168), .B(n1169), .Z(n1164) );
XOR2_X1 U842 ( .A(G110), .B(n1170), .Z(n1169) );
NOR2_X1 U843 ( .A1(n1171), .A2(n1139), .ZN(n1170) );
INV_X1 U844 ( .A(G469), .ZN(n1171) );
NAND2_X1 U845 ( .A1(KEYINPUT54), .A2(n1172), .ZN(n1168) );
NOR2_X1 U846 ( .A1(n1135), .A2(n1173), .ZN(G51) );
XOR2_X1 U847 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U848 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U849 ( .A1(KEYINPUT34), .A2(n1178), .ZN(n1176) );
XOR2_X1 U850 ( .A(n1179), .B(n1180), .Z(n1174) );
NOR2_X1 U851 ( .A1(n1181), .A2(n1139), .ZN(n1180) );
NAND2_X1 U852 ( .A1(G902), .A2(n1053), .ZN(n1139) );
NAND4_X1 U853 ( .A1(n1182), .A2(n1111), .A3(n1183), .A4(n1131), .ZN(n1053) );
AND4_X1 U854 ( .A1(n1048), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1131) );
NOR2_X1 U855 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NOR2_X1 U856 ( .A1(n1067), .A2(n1189), .ZN(n1188) );
NOR2_X1 U857 ( .A1(n1190), .A2(n1191), .ZN(n1067) );
NOR3_X1 U858 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1187) );
INV_X1 U859 ( .A(n1077), .ZN(n1194) );
XOR2_X1 U860 ( .A(n1195), .B(KEYINPUT10), .Z(n1193) );
NAND3_X1 U861 ( .A1(n1082), .A2(n1081), .A3(n1196), .ZN(n1048) );
NOR2_X1 U862 ( .A1(n1132), .A2(n1133), .ZN(n1183) );
AND3_X1 U863 ( .A1(n1196), .A2(n1081), .A3(n1083), .ZN(n1133) );
AND3_X1 U864 ( .A1(n1197), .A2(n1082), .A3(n1190), .ZN(n1132) );
AND4_X1 U865 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1111) );
NOR4_X1 U866 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
INV_X1 U867 ( .A(n1206), .ZN(n1204) );
NAND3_X1 U868 ( .A1(n1082), .A2(n1072), .A3(n1207), .ZN(n1200) );
XOR2_X1 U869 ( .A(n1110), .B(KEYINPUT21), .Z(n1182) );
NOR2_X1 U870 ( .A1(n1208), .A2(n1209), .ZN(n1179) );
XOR2_X1 U871 ( .A(KEYINPUT41), .B(n1210), .Z(n1209) );
NOR2_X1 U872 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NOR2_X1 U873 ( .A1(G125), .A2(n1213), .ZN(n1208) );
XOR2_X1 U874 ( .A(n1211), .B(KEYINPUT2), .Z(n1213) );
NOR2_X1 U875 ( .A1(n1214), .A2(G952), .ZN(n1135) );
XOR2_X1 U876 ( .A(KEYINPUT51), .B(n1128), .Z(n1214) );
XNOR2_X1 U877 ( .A(G146), .B(n1215), .ZN(G48) );
NAND2_X1 U878 ( .A1(KEYINPUT28), .A2(n1203), .ZN(n1215) );
AND3_X1 U879 ( .A1(n1083), .A2(n1072), .A3(n1207), .ZN(n1203) );
XOR2_X1 U880 ( .A(n1216), .B(n1199), .Z(G45) );
NAND4_X1 U881 ( .A1(n1217), .A2(n1072), .A3(n1190), .A4(n1218), .ZN(n1199) );
NOR3_X1 U882 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1218) );
XOR2_X1 U883 ( .A(G140), .B(n1202), .Z(G42) );
AND3_X1 U884 ( .A1(n1222), .A2(n1083), .A3(n1191), .ZN(n1202) );
XOR2_X1 U885 ( .A(n1223), .B(G137), .Z(G39) );
NAND2_X1 U886 ( .A1(KEYINPUT29), .A2(n1198), .ZN(n1223) );
NAND2_X1 U887 ( .A1(n1224), .A2(n1222), .ZN(n1198) );
INV_X1 U888 ( .A(n1192), .ZN(n1224) );
XOR2_X1 U889 ( .A(n1107), .B(n1225), .Z(G36) );
NAND2_X1 U890 ( .A1(KEYINPUT63), .A2(n1226), .ZN(n1225) );
INV_X1 U891 ( .A(n1110), .ZN(n1226) );
NAND3_X1 U892 ( .A1(n1190), .A2(n1082), .A3(n1222), .ZN(n1110) );
XOR2_X1 U893 ( .A(G131), .B(n1205), .Z(G33) );
AND3_X1 U894 ( .A1(n1083), .A2(n1190), .A3(n1222), .ZN(n1205) );
NOR3_X1 U895 ( .A1(n1227), .A2(n1220), .A3(n1064), .ZN(n1222) );
NAND2_X1 U896 ( .A1(n1228), .A2(n1229), .ZN(n1064) );
XOR2_X1 U897 ( .A(KEYINPUT42), .B(n1079), .Z(n1229) );
INV_X1 U898 ( .A(n1230), .ZN(n1220) );
XNOR2_X1 U899 ( .A(G128), .B(n1231), .ZN(G30) );
NAND3_X1 U900 ( .A1(n1082), .A2(n1232), .A3(n1207), .ZN(n1231) );
AND4_X1 U901 ( .A1(n1233), .A2(n1234), .A3(n1230), .A4(n1235), .ZN(n1207) );
XOR2_X1 U902 ( .A(KEYINPUT59), .B(n1072), .Z(n1232) );
XOR2_X1 U903 ( .A(G101), .B(n1236), .Z(G3) );
NOR2_X1 U904 ( .A1(n1237), .A2(n1189), .ZN(n1236) );
INV_X1 U905 ( .A(n1190), .ZN(n1237) );
XOR2_X1 U906 ( .A(n1212), .B(n1206), .Z(G27) );
NAND4_X1 U907 ( .A1(n1191), .A2(n1083), .A3(n1077), .A4(n1230), .ZN(n1206) );
NAND2_X1 U908 ( .A1(n1055), .A2(n1238), .ZN(n1230) );
NAND2_X1 U909 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
INV_X1 U910 ( .A(G900), .ZN(n1240) );
XNOR2_X1 U911 ( .A(n1184), .B(n1241), .ZN(G24) );
NOR2_X1 U912 ( .A1(KEYINPUT39), .A2(n1242), .ZN(n1241) );
NAND4_X1 U913 ( .A1(n1197), .A2(n1081), .A3(n1217), .A4(n1058), .ZN(n1184) );
INV_X1 U914 ( .A(n1221), .ZN(n1058) );
NOR2_X1 U915 ( .A1(n1235), .A2(n1234), .ZN(n1081) );
XOR2_X1 U916 ( .A(n1243), .B(n1244), .Z(G21) );
NOR2_X1 U917 ( .A1(n1245), .A2(n1192), .ZN(n1244) );
NAND4_X1 U918 ( .A1(n1221), .A2(n1234), .A3(n1246), .A4(n1235), .ZN(n1192) );
INV_X1 U919 ( .A(n1247), .ZN(n1234) );
XNOR2_X1 U920 ( .A(G119), .B(KEYINPUT13), .ZN(n1243) );
NAND2_X1 U921 ( .A1(n1248), .A2(n1249), .ZN(G18) );
NAND2_X1 U922 ( .A1(G116), .A2(n1250), .ZN(n1249) );
XOR2_X1 U923 ( .A(KEYINPUT36), .B(n1251), .Z(n1248) );
NOR2_X1 U924 ( .A1(G116), .A2(n1250), .ZN(n1251) );
NAND4_X1 U925 ( .A1(n1252), .A2(n1190), .A3(n1077), .A4(n1082), .ZN(n1250) );
AND2_X1 U926 ( .A1(n1221), .A2(n1217), .ZN(n1082) );
XOR2_X1 U927 ( .A(n1060), .B(KEYINPUT25), .Z(n1217) );
XOR2_X1 U928 ( .A(n1195), .B(KEYINPUT52), .Z(n1252) );
NAND2_X1 U929 ( .A1(n1253), .A2(n1254), .ZN(G15) );
NAND2_X1 U930 ( .A1(G113), .A2(n1185), .ZN(n1254) );
XOR2_X1 U931 ( .A(KEYINPUT1), .B(n1255), .Z(n1253) );
NOR2_X1 U932 ( .A1(G113), .A2(n1185), .ZN(n1255) );
NAND3_X1 U933 ( .A1(n1190), .A2(n1197), .A3(n1083), .ZN(n1185) );
NOR2_X1 U934 ( .A1(n1060), .A2(n1221), .ZN(n1083) );
INV_X1 U935 ( .A(n1245), .ZN(n1197) );
NAND2_X1 U936 ( .A1(n1077), .A2(n1195), .ZN(n1245) );
NOR2_X1 U937 ( .A1(n1068), .A2(n1219), .ZN(n1077) );
NAND2_X1 U938 ( .A1(n1256), .A2(n1074), .ZN(n1068) );
NOR2_X1 U939 ( .A1(n1235), .A2(n1247), .ZN(n1190) );
XOR2_X1 U940 ( .A(G110), .B(n1257), .Z(G12) );
NOR2_X1 U941 ( .A1(n1258), .A2(n1189), .ZN(n1257) );
NAND3_X1 U942 ( .A1(n1221), .A2(n1246), .A3(n1196), .ZN(n1189) );
AND3_X1 U943 ( .A1(n1233), .A2(n1195), .A3(n1072), .ZN(n1196) );
INV_X1 U944 ( .A(n1227), .ZN(n1072) );
NAND2_X1 U945 ( .A1(n1073), .A2(n1074), .ZN(n1227) );
NAND2_X1 U946 ( .A1(G221), .A2(n1259), .ZN(n1074) );
INV_X1 U947 ( .A(n1256), .ZN(n1073) );
XOR2_X1 U948 ( .A(n1260), .B(G469), .Z(n1256) );
NAND2_X1 U949 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U950 ( .A(n1263), .B(n1264), .Z(n1261) );
XNOR2_X1 U951 ( .A(n1265), .B(n1167), .ZN(n1264) );
XNOR2_X1 U952 ( .A(n1266), .B(n1267), .ZN(n1167) );
XOR2_X1 U953 ( .A(G104), .B(n1268), .Z(n1267) );
AND2_X1 U954 ( .A1(n1128), .A2(G227), .ZN(n1268) );
XNOR2_X1 U955 ( .A(n1158), .B(n1269), .ZN(n1266) );
NAND2_X1 U956 ( .A1(KEYINPUT23), .A2(n1270), .ZN(n1265) );
XOR2_X1 U957 ( .A(n1105), .B(n1271), .Z(n1263) );
XOR2_X1 U958 ( .A(n1172), .B(KEYINPUT7), .Z(n1271) );
NAND2_X1 U959 ( .A1(n1272), .A2(n1273), .ZN(n1105) );
OR2_X1 U960 ( .A1(n1274), .A2(G128), .ZN(n1273) );
XOR2_X1 U961 ( .A(n1275), .B(KEYINPUT18), .Z(n1272) );
NAND2_X1 U962 ( .A1(G128), .A2(n1274), .ZN(n1275) );
XNOR2_X1 U963 ( .A(n1216), .B(n1276), .ZN(n1274) );
XOR2_X1 U964 ( .A(KEYINPUT44), .B(G146), .Z(n1276) );
NAND2_X1 U965 ( .A1(n1055), .A2(n1277), .ZN(n1195) );
NAND2_X1 U966 ( .A1(n1239), .A2(n1278), .ZN(n1277) );
INV_X1 U967 ( .A(G898), .ZN(n1278) );
NOR3_X1 U968 ( .A1(n1108), .A2(n1279), .A3(n1262), .ZN(n1239) );
INV_X1 U969 ( .A(n1280), .ZN(n1279) );
XNOR2_X1 U970 ( .A(n1128), .B(KEYINPUT38), .ZN(n1108) );
NAND3_X1 U971 ( .A1(n1280), .A2(n1128), .A3(G952), .ZN(n1055) );
NAND2_X1 U972 ( .A1(G237), .A2(G234), .ZN(n1280) );
INV_X1 U973 ( .A(n1219), .ZN(n1233) );
NAND2_X1 U974 ( .A1(n1228), .A2(n1079), .ZN(n1219) );
XOR2_X1 U975 ( .A(n1281), .B(n1181), .Z(n1079) );
NAND2_X1 U976 ( .A1(G210), .A2(n1282), .ZN(n1181) );
NAND2_X1 U977 ( .A1(n1283), .A2(n1262), .ZN(n1281) );
XOR2_X1 U978 ( .A(n1177), .B(n1284), .Z(n1283) );
XNOR2_X1 U979 ( .A(n1285), .B(KEYINPUT46), .ZN(n1284) );
NAND2_X1 U980 ( .A1(n1286), .A2(KEYINPUT61), .ZN(n1285) );
XOR2_X1 U981 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U982 ( .A(KEYINPUT17), .B(G125), .Z(n1288) );
XOR2_X1 U983 ( .A(n1162), .B(n1178), .Z(n1287) );
NAND2_X1 U984 ( .A1(G224), .A2(n1128), .ZN(n1178) );
INV_X1 U985 ( .A(n1211), .ZN(n1162) );
XOR2_X1 U986 ( .A(n1289), .B(n1290), .Z(n1177) );
NOR2_X1 U987 ( .A1(n1124), .A2(n1291), .ZN(n1290) );
AND2_X1 U988 ( .A1(n1123), .A2(n1122), .ZN(n1291) );
NOR2_X1 U989 ( .A1(n1123), .A2(n1122), .ZN(n1124) );
AND2_X1 U990 ( .A1(n1292), .A2(n1293), .ZN(n1122) );
OR2_X1 U991 ( .A1(n1294), .A2(G119), .ZN(n1293) );
NAND2_X1 U992 ( .A1(G119), .A2(n1295), .ZN(n1292) );
XNOR2_X1 U993 ( .A(n1294), .B(KEYINPUT37), .ZN(n1295) );
XOR2_X1 U994 ( .A(n1269), .B(n1296), .Z(n1123) );
NOR2_X1 U995 ( .A1(KEYINPUT9), .A2(n1153), .ZN(n1296) );
INV_X1 U996 ( .A(G104), .ZN(n1153) );
XOR2_X1 U997 ( .A(G101), .B(G107), .Z(n1269) );
NAND2_X1 U998 ( .A1(KEYINPUT14), .A2(n1117), .ZN(n1289) );
XOR2_X1 U999 ( .A(n1270), .B(G122), .Z(n1117) );
XOR2_X1 U1000 ( .A(n1078), .B(KEYINPUT56), .Z(n1228) );
NAND2_X1 U1001 ( .A1(G214), .A2(n1282), .ZN(n1078) );
NAND2_X1 U1002 ( .A1(n1297), .A2(n1262), .ZN(n1282) );
INV_X1 U1003 ( .A(G237), .ZN(n1297) );
INV_X1 U1004 ( .A(n1060), .ZN(n1246) );
XOR2_X1 U1005 ( .A(n1298), .B(n1096), .Z(n1060) );
NOR2_X1 U1006 ( .A1(n1145), .A2(G902), .ZN(n1096) );
XOR2_X1 U1007 ( .A(n1299), .B(n1300), .Z(n1145) );
NOR2_X1 U1008 ( .A1(KEYINPUT22), .A2(n1301), .ZN(n1300) );
XOR2_X1 U1009 ( .A(n1302), .B(n1303), .Z(n1301) );
NAND2_X1 U1010 ( .A1(KEYINPUT20), .A2(n1304), .ZN(n1303) );
NAND2_X1 U1011 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND2_X1 U1012 ( .A1(n1307), .A2(n1107), .ZN(n1306) );
XOR2_X1 U1013 ( .A(n1308), .B(KEYINPUT3), .Z(n1305) );
OR2_X1 U1014 ( .A1(n1307), .A2(n1107), .ZN(n1308) );
INV_X1 U1015 ( .A(G134), .ZN(n1107) );
XNOR2_X1 U1016 ( .A(n1309), .B(G128), .ZN(n1307) );
NAND2_X1 U1017 ( .A1(KEYINPUT47), .A2(n1216), .ZN(n1309) );
NAND2_X1 U1018 ( .A1(n1310), .A2(n1311), .ZN(n1302) );
NAND3_X1 U1019 ( .A1(KEYINPUT50), .A2(n1312), .A3(n1313), .ZN(n1311) );
XOR2_X1 U1020 ( .A(n1314), .B(G107), .Z(n1313) );
NAND2_X1 U1021 ( .A1(KEYINPUT35), .A2(G122), .ZN(n1314) );
NAND2_X1 U1022 ( .A1(n1315), .A2(n1316), .ZN(n1310) );
NAND2_X1 U1023 ( .A1(KEYINPUT50), .A2(n1312), .ZN(n1316) );
INV_X1 U1024 ( .A(G116), .ZN(n1312) );
XOR2_X1 U1025 ( .A(n1317), .B(G107), .Z(n1315) );
NAND2_X1 U1026 ( .A1(KEYINPUT35), .A2(n1242), .ZN(n1317) );
INV_X1 U1027 ( .A(G122), .ZN(n1242) );
NAND2_X1 U1028 ( .A1(G217), .A2(n1318), .ZN(n1299) );
NAND2_X1 U1029 ( .A1(KEYINPUT12), .A2(n1144), .ZN(n1298) );
INV_X1 U1030 ( .A(G478), .ZN(n1144) );
XOR2_X1 U1031 ( .A(n1319), .B(G475), .Z(n1221) );
NAND2_X1 U1032 ( .A1(n1148), .A2(n1262), .ZN(n1319) );
XOR2_X1 U1033 ( .A(n1320), .B(n1321), .Z(n1148) );
XOR2_X1 U1034 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U1035 ( .A(G122), .B(G113), .Z(n1323) );
XOR2_X1 U1036 ( .A(G146), .B(G143), .Z(n1322) );
XOR2_X1 U1037 ( .A(n1324), .B(n1325), .Z(n1320) );
XOR2_X1 U1038 ( .A(G104), .B(n1326), .Z(n1325) );
NOR2_X1 U1039 ( .A1(KEYINPUT5), .A2(n1327), .ZN(n1326) );
XOR2_X1 U1040 ( .A(n1212), .B(n1328), .Z(n1327) );
NAND2_X1 U1041 ( .A1(KEYINPUT40), .A2(n1172), .ZN(n1328) );
INV_X1 U1042 ( .A(G140), .ZN(n1172) );
INV_X1 U1043 ( .A(G125), .ZN(n1212) );
XOR2_X1 U1044 ( .A(n1329), .B(n1330), .Z(n1324) );
NOR2_X1 U1045 ( .A1(KEYINPUT43), .A2(G131), .ZN(n1330) );
NAND2_X1 U1046 ( .A1(n1331), .A2(G214), .ZN(n1329) );
XNOR2_X1 U1047 ( .A(n1191), .B(KEYINPUT27), .ZN(n1258) );
AND2_X1 U1048 ( .A1(n1247), .A2(n1235), .ZN(n1191) );
NAND3_X1 U1049 ( .A1(n1332), .A2(n1333), .A3(n1092), .ZN(n1235) );
NAND2_X1 U1050 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U1051 ( .A1(KEYINPUT53), .A2(n1094), .ZN(n1333) );
OR3_X1 U1052 ( .A1(n1093), .A2(KEYINPUT53), .A3(n1094), .ZN(n1332) );
NAND2_X1 U1053 ( .A1(G217), .A2(n1259), .ZN(n1094) );
NAND2_X1 U1054 ( .A1(G234), .A2(n1262), .ZN(n1259) );
NOR2_X1 U1055 ( .A1(n1137), .A2(G902), .ZN(n1093) );
XOR2_X1 U1056 ( .A(n1334), .B(n1335), .Z(n1137) );
XOR2_X1 U1057 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1058 ( .A(G137), .B(G119), .Z(n1337) );
XOR2_X1 U1059 ( .A(KEYINPUT57), .B(KEYINPUT32), .Z(n1336) );
XOR2_X1 U1060 ( .A(n1338), .B(n1339), .Z(n1334) );
XOR2_X1 U1061 ( .A(n1340), .B(n1104), .Z(n1339) );
XOR2_X1 U1062 ( .A(G140), .B(G125), .Z(n1104) );
XNOR2_X1 U1063 ( .A(n1341), .B(n1342), .ZN(n1338) );
NAND3_X1 U1064 ( .A1(n1318), .A2(G221), .A3(KEYINPUT6), .ZN(n1342) );
AND2_X1 U1065 ( .A1(G234), .A2(n1128), .ZN(n1318) );
INV_X1 U1066 ( .A(G953), .ZN(n1128) );
NAND2_X1 U1067 ( .A1(KEYINPUT45), .A2(n1270), .ZN(n1341) );
INV_X1 U1068 ( .A(G110), .ZN(n1270) );
XOR2_X1 U1069 ( .A(n1090), .B(G472), .Z(n1247) );
NAND2_X1 U1070 ( .A1(n1343), .A2(n1262), .ZN(n1090) );
INV_X1 U1071 ( .A(G902), .ZN(n1262) );
XOR2_X1 U1072 ( .A(n1344), .B(n1157), .Z(n1343) );
XOR2_X1 U1073 ( .A(n1345), .B(n1346), .Z(n1157) );
XOR2_X1 U1074 ( .A(G119), .B(G101), .Z(n1346) );
XOR2_X1 U1075 ( .A(n1347), .B(n1294), .Z(n1345) );
XOR2_X1 U1076 ( .A(G113), .B(G116), .Z(n1294) );
NAND2_X1 U1077 ( .A1(n1331), .A2(G210), .ZN(n1347) );
NOR2_X1 U1078 ( .A1(G953), .A2(G237), .ZN(n1331) );
NAND2_X1 U1079 ( .A1(n1348), .A2(KEYINPUT58), .ZN(n1344) );
XOR2_X1 U1080 ( .A(n1211), .B(n1349), .Z(n1348) );
NOR2_X1 U1081 ( .A1(KEYINPUT60), .A2(n1350), .ZN(n1349) );
XOR2_X1 U1082 ( .A(KEYINPUT33), .B(n1158), .Z(n1350) );
XOR2_X1 U1083 ( .A(n1103), .B(G134), .Z(n1158) );
XOR2_X1 U1084 ( .A(G131), .B(n1351), .Z(n1103) );
XOR2_X1 U1085 ( .A(KEYINPUT31), .B(G137), .Z(n1351) );
XOR2_X1 U1086 ( .A(n1352), .B(n1340), .Z(n1211) );
XOR2_X1 U1087 ( .A(G128), .B(G146), .Z(n1340) );
NAND2_X1 U1088 ( .A1(KEYINPUT49), .A2(n1216), .ZN(n1352) );
INV_X1 U1089 ( .A(G143), .ZN(n1216) );
endmodule


