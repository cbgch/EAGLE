//Key = 0001101010011010011111101111100100010001010001111110000000101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376;

XOR2_X1 U745 ( .A(G107), .B(n1038), .Z(G9) );
NOR2_X1 U746 ( .A1(n1039), .A2(n1040), .ZN(G75) );
AND3_X1 U747 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NOR4_X1 U748 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1039) );
NOR2_X1 U749 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR3_X1 U750 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1048) );
NAND4_X1 U751 ( .A1(n1041), .A2(n1053), .A3(n1054), .A4(n1042), .ZN(n1044) );
NAND4_X1 U752 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NAND2_X1 U753 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U754 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
OR2_X1 U755 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U756 ( .A1(n1065), .A2(n1066), .ZN(n1059) );
XOR2_X1 U757 ( .A(n1067), .B(n1068), .Z(n1065) );
NAND2_X1 U758 ( .A1(n1069), .A2(n1070), .ZN(n1053) );
NAND2_X1 U759 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U760 ( .A1(n1056), .A2(n1073), .ZN(n1072) );
NAND2_X1 U761 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U762 ( .A1(n1076), .A2(n1049), .ZN(n1075) );
INV_X1 U763 ( .A(KEYINPUT13), .ZN(n1049) );
INV_X1 U764 ( .A(n1052), .ZN(n1056) );
NAND2_X1 U765 ( .A1(n1057), .A2(n1077), .ZN(n1071) );
NAND2_X1 U766 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U767 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U768 ( .A(n1082), .B(KEYINPUT17), .Z(n1080) );
INV_X1 U769 ( .A(n1050), .ZN(n1069) );
NAND3_X1 U770 ( .A1(n1066), .A2(n1061), .A3(n1055), .ZN(n1050) );
INV_X1 U771 ( .A(n1083), .ZN(n1055) );
NAND4_X1 U772 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1041) );
NOR4_X1 U773 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1087) );
XNOR2_X1 U774 ( .A(KEYINPUT42), .B(n1092), .ZN(n1091) );
XOR2_X1 U775 ( .A(n1093), .B(n1094), .Z(n1090) );
XNOR2_X1 U776 ( .A(G472), .B(n1095), .ZN(n1089) );
NAND3_X1 U777 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1088) );
XOR2_X1 U778 ( .A(n1099), .B(G478), .Z(n1098) );
OR3_X1 U779 ( .A1(n1100), .A2(n1101), .A3(KEYINPUT32), .ZN(n1097) );
NAND2_X1 U780 ( .A1(KEYINPUT32), .A2(n1100), .ZN(n1096) );
NOR3_X1 U781 ( .A1(n1067), .A2(n1102), .A3(n1103), .ZN(n1086) );
XOR2_X1 U782 ( .A(KEYINPUT48), .B(n1104), .Z(n1084) );
XOR2_X1 U783 ( .A(n1105), .B(n1106), .Z(G72) );
XOR2_X1 U784 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U785 ( .A1(n1109), .A2(n1042), .ZN(n1108) );
NOR2_X1 U786 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U787 ( .A1(n1112), .A2(n1113), .ZN(n1107) );
NAND2_X1 U788 ( .A1(G953), .A2(n1111), .ZN(n1113) );
XOR2_X1 U789 ( .A(n1114), .B(n1115), .Z(n1112) );
XOR2_X1 U790 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U791 ( .A(G131), .B(n1118), .Z(n1117) );
XOR2_X1 U792 ( .A(n1119), .B(n1120), .Z(n1114) );
XOR2_X1 U793 ( .A(G137), .B(G134), .Z(n1120) );
XNOR2_X1 U794 ( .A(KEYINPUT6), .B(KEYINPUT47), .ZN(n1119) );
NAND2_X1 U795 ( .A1(n1042), .A2(n1047), .ZN(n1105) );
NAND2_X1 U796 ( .A1(n1121), .A2(n1122), .ZN(G69) );
NAND2_X1 U797 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U798 ( .A(n1125), .B(KEYINPUT40), .Z(n1123) );
XOR2_X1 U799 ( .A(KEYINPUT21), .B(n1126), .Z(n1121) );
NOR2_X1 U800 ( .A1(n1124), .A2(n1125), .ZN(n1126) );
XOR2_X1 U801 ( .A(n1127), .B(n1128), .Z(n1125) );
NOR2_X1 U802 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XOR2_X1 U803 ( .A(n1042), .B(KEYINPUT22), .Z(n1130) );
INV_X1 U804 ( .A(n1045), .ZN(n1129) );
NAND2_X1 U805 ( .A1(n1131), .A2(n1132), .ZN(n1127) );
NAND2_X1 U806 ( .A1(G953), .A2(n1133), .ZN(n1132) );
XOR2_X1 U807 ( .A(n1134), .B(G101), .Z(n1131) );
AND2_X1 U808 ( .A1(G953), .A2(n1135), .ZN(n1124) );
NAND2_X1 U809 ( .A1(G898), .A2(G224), .ZN(n1135) );
NOR3_X1 U810 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(G66) );
AND2_X1 U811 ( .A1(KEYINPUT18), .A2(n1139), .ZN(n1138) );
NOR3_X1 U812 ( .A1(KEYINPUT18), .A2(G953), .A3(G952), .ZN(n1137) );
XOR2_X1 U813 ( .A(n1140), .B(n1141), .Z(n1136) );
NOR2_X1 U814 ( .A1(KEYINPUT16), .A2(n1142), .ZN(n1141) );
INV_X1 U815 ( .A(n1143), .ZN(n1142) );
NAND2_X1 U816 ( .A1(n1144), .A2(n1145), .ZN(n1140) );
NOR2_X1 U817 ( .A1(n1139), .A2(n1146), .ZN(G63) );
XOR2_X1 U818 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U819 ( .A(KEYINPUT63), .B(n1149), .Z(n1148) );
AND2_X1 U820 ( .A1(G478), .A2(n1144), .ZN(n1149) );
NOR3_X1 U821 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(G60) );
AND2_X1 U822 ( .A1(n1139), .A2(KEYINPUT31), .ZN(n1152) );
NOR3_X1 U823 ( .A1(KEYINPUT31), .A2(n1042), .A3(n1043), .ZN(n1151) );
INV_X1 U824 ( .A(G952), .ZN(n1043) );
NOR2_X1 U825 ( .A1(n1153), .A2(n1154), .ZN(n1150) );
XOR2_X1 U826 ( .A(KEYINPUT38), .B(n1155), .Z(n1154) );
NOR2_X1 U827 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
AND2_X1 U828 ( .A1(n1157), .A2(n1156), .ZN(n1153) );
NAND2_X1 U829 ( .A1(n1144), .A2(G475), .ZN(n1156) );
XOR2_X1 U830 ( .A(n1158), .B(n1159), .Z(G6) );
XNOR2_X1 U831 ( .A(G104), .B(KEYINPUT11), .ZN(n1159) );
NAND2_X1 U832 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
NAND2_X1 U833 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
INV_X1 U834 ( .A(KEYINPUT56), .ZN(n1163) );
NAND3_X1 U835 ( .A1(n1164), .A2(n1165), .A3(KEYINPUT56), .ZN(n1160) );
NOR2_X1 U836 ( .A1(n1166), .A2(n1167), .ZN(G57) );
XOR2_X1 U837 ( .A(KEYINPUT51), .B(n1139), .Z(n1167) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1166) );
XOR2_X1 U839 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U840 ( .A(n1172), .B(n1173), .Z(n1168) );
AND2_X1 U841 ( .A1(G472), .A2(n1144), .ZN(n1173) );
INV_X1 U842 ( .A(n1174), .ZN(n1144) );
XOR2_X1 U843 ( .A(n1175), .B(KEYINPUT36), .Z(n1172) );
NOR2_X1 U844 ( .A1(n1139), .A2(n1176), .ZN(G54) );
XOR2_X1 U845 ( .A(n1177), .B(n1178), .Z(n1176) );
XNOR2_X1 U846 ( .A(n1179), .B(n1180), .ZN(n1178) );
XOR2_X1 U847 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U848 ( .A1(n1093), .A2(n1174), .ZN(n1182) );
NAND2_X1 U849 ( .A1(KEYINPUT28), .A2(n1116), .ZN(n1181) );
XNOR2_X1 U850 ( .A(n1183), .B(n1184), .ZN(n1116) );
XOR2_X1 U851 ( .A(n1185), .B(n1186), .Z(n1177) );
XNOR2_X1 U852 ( .A(n1187), .B(n1188), .ZN(n1186) );
NOR2_X1 U853 ( .A1(KEYINPUT53), .A2(n1189), .ZN(n1188) );
XOR2_X1 U854 ( .A(n1190), .B(n1191), .Z(n1185) );
NOR2_X1 U855 ( .A1(n1139), .A2(n1192), .ZN(G51) );
NOR2_X1 U856 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XOR2_X1 U857 ( .A(n1195), .B(n1196), .Z(n1194) );
NOR2_X1 U858 ( .A1(n1100), .A2(n1174), .ZN(n1196) );
NAND2_X1 U859 ( .A1(G902), .A2(n1197), .ZN(n1174) );
OR2_X1 U860 ( .A1(n1045), .A2(n1047), .ZN(n1197) );
NAND2_X1 U861 ( .A1(n1198), .A2(n1199), .ZN(n1047) );
AND4_X1 U862 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
NOR4_X1 U863 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1198) );
INV_X1 U864 ( .A(n1208), .ZN(n1207) );
INV_X1 U865 ( .A(n1209), .ZN(n1206) );
NAND4_X1 U866 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1045) );
NOR4_X1 U867 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1213) );
AND3_X1 U868 ( .A1(n1218), .A2(n1219), .A3(n1066), .ZN(n1217) );
INV_X1 U869 ( .A(n1220), .ZN(n1216) );
INV_X1 U870 ( .A(n1221), .ZN(n1214) );
NOR2_X1 U871 ( .A1(n1162), .A2(n1038), .ZN(n1212) );
AND4_X1 U872 ( .A1(n1064), .A2(n1222), .A3(n1057), .A4(n1223), .ZN(n1038) );
AND2_X1 U873 ( .A1(n1165), .A2(n1223), .ZN(n1162) );
AND3_X1 U874 ( .A1(n1222), .A2(n1057), .A3(n1063), .ZN(n1165) );
NOR2_X1 U875 ( .A1(KEYINPUT29), .A2(n1224), .ZN(n1195) );
AND2_X1 U876 ( .A1(n1224), .A2(KEYINPUT29), .ZN(n1193) );
NOR2_X1 U877 ( .A1(n1042), .A2(G952), .ZN(n1139) );
NAND2_X1 U878 ( .A1(n1225), .A2(n1226), .ZN(G48) );
NAND2_X1 U879 ( .A1(G146), .A2(n1208), .ZN(n1226) );
XOR2_X1 U880 ( .A(KEYINPUT25), .B(n1227), .Z(n1225) );
NOR2_X1 U881 ( .A1(G146), .A2(n1208), .ZN(n1227) );
NAND4_X1 U882 ( .A1(n1218), .A2(n1063), .A3(n1222), .A4(n1228), .ZN(n1208) );
XOR2_X1 U883 ( .A(n1229), .B(n1209), .Z(G45) );
NAND3_X1 U884 ( .A1(n1230), .A2(n1222), .A3(n1231), .ZN(n1209) );
NOR3_X1 U885 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1231) );
XOR2_X1 U886 ( .A(G140), .B(n1205), .Z(G42) );
AND3_X1 U887 ( .A1(n1076), .A2(n1063), .A3(n1235), .ZN(n1205) );
XOR2_X1 U888 ( .A(G137), .B(n1204), .Z(G39) );
AND3_X1 U889 ( .A1(n1218), .A2(n1066), .A3(n1235), .ZN(n1204) );
XNOR2_X1 U890 ( .A(n1203), .B(n1236), .ZN(G36) );
XOR2_X1 U891 ( .A(KEYINPUT61), .B(G134), .Z(n1236) );
NAND3_X1 U892 ( .A1(n1230), .A2(n1064), .A3(n1235), .ZN(n1203) );
XOR2_X1 U893 ( .A(n1202), .B(n1237), .Z(G33) );
NOR2_X1 U894 ( .A1(G131), .A2(KEYINPUT55), .ZN(n1237) );
NAND3_X1 U895 ( .A1(n1063), .A2(n1230), .A3(n1235), .ZN(n1202) );
NOR4_X1 U896 ( .A1(n1238), .A2(n1052), .A3(n1233), .A4(n1067), .ZN(n1235) );
NAND2_X1 U897 ( .A1(n1239), .A2(n1082), .ZN(n1052) );
XNOR2_X1 U898 ( .A(n1081), .B(KEYINPUT35), .ZN(n1239) );
XNOR2_X1 U899 ( .A(G128), .B(n1201), .ZN(G30) );
NAND4_X1 U900 ( .A1(n1218), .A2(n1064), .A3(n1222), .A4(n1228), .ZN(n1201) );
XOR2_X1 U901 ( .A(n1190), .B(n1210), .Z(G3) );
NAND4_X1 U902 ( .A1(n1230), .A2(n1066), .A3(n1222), .A4(n1223), .ZN(n1210) );
XOR2_X1 U903 ( .A(n1240), .B(n1200), .Z(G27) );
NAND4_X1 U904 ( .A1(n1076), .A2(n1063), .A3(n1241), .A4(n1061), .ZN(n1200) );
NOR2_X1 U905 ( .A1(n1233), .A2(n1078), .ZN(n1241) );
INV_X1 U906 ( .A(n1228), .ZN(n1233) );
NAND2_X1 U907 ( .A1(n1083), .A2(n1242), .ZN(n1228) );
NAND4_X1 U908 ( .A1(G953), .A2(G902), .A3(n1243), .A4(n1111), .ZN(n1242) );
INV_X1 U909 ( .A(G900), .ZN(n1111) );
INV_X1 U910 ( .A(n1244), .ZN(n1063) );
XNOR2_X1 U911 ( .A(G122), .B(n1211), .ZN(G24) );
NAND4_X1 U912 ( .A1(n1219), .A2(n1057), .A3(n1245), .A4(n1104), .ZN(n1211) );
NOR2_X1 U913 ( .A1(n1246), .A2(n1247), .ZN(n1057) );
XOR2_X1 U914 ( .A(n1248), .B(n1249), .Z(G21) );
NAND2_X1 U915 ( .A1(KEYINPUT4), .A2(G119), .ZN(n1249) );
NAND4_X1 U916 ( .A1(n1218), .A2(n1066), .A3(n1250), .A4(n1061), .ZN(n1248) );
NOR2_X1 U917 ( .A1(n1164), .A2(n1251), .ZN(n1250) );
XOR2_X1 U918 ( .A(n1078), .B(KEYINPUT34), .Z(n1251) );
INV_X1 U919 ( .A(n1223), .ZN(n1164) );
AND2_X1 U920 ( .A1(n1247), .A2(n1246), .ZN(n1218) );
INV_X1 U921 ( .A(n1252), .ZN(n1247) );
XOR2_X1 U922 ( .A(G116), .B(n1253), .Z(G18) );
NOR2_X1 U923 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
AND2_X1 U924 ( .A1(KEYINPUT46), .A2(n1220), .ZN(n1255) );
NOR2_X1 U925 ( .A1(KEYINPUT8), .A2(n1220), .ZN(n1254) );
NAND3_X1 U926 ( .A1(n1219), .A2(n1064), .A3(n1230), .ZN(n1220) );
NOR2_X1 U927 ( .A1(n1104), .A2(n1232), .ZN(n1064) );
INV_X1 U928 ( .A(n1256), .ZN(n1219) );
XOR2_X1 U929 ( .A(G113), .B(n1215), .Z(G15) );
NOR3_X1 U930 ( .A1(n1074), .A2(n1256), .A3(n1244), .ZN(n1215) );
NAND2_X1 U931 ( .A1(n1257), .A2(n1232), .ZN(n1244) );
INV_X1 U932 ( .A(n1245), .ZN(n1232) );
XOR2_X1 U933 ( .A(n1234), .B(KEYINPUT58), .Z(n1257) );
NAND3_X1 U934 ( .A1(n1258), .A2(n1223), .A3(n1061), .ZN(n1256) );
NOR2_X1 U935 ( .A1(n1068), .A2(n1067), .ZN(n1061) );
INV_X1 U936 ( .A(n1230), .ZN(n1074) );
NOR2_X1 U937 ( .A1(n1246), .A2(n1252), .ZN(n1230) );
XOR2_X1 U938 ( .A(n1259), .B(n1221), .Z(G12) );
NAND4_X1 U939 ( .A1(n1076), .A2(n1066), .A3(n1222), .A4(n1223), .ZN(n1221) );
NAND2_X1 U940 ( .A1(n1083), .A2(n1260), .ZN(n1223) );
NAND4_X1 U941 ( .A1(G953), .A2(G902), .A3(n1243), .A4(n1133), .ZN(n1260) );
INV_X1 U942 ( .A(G898), .ZN(n1133) );
NAND3_X1 U943 ( .A1(n1243), .A2(n1042), .A3(G952), .ZN(n1083) );
NAND2_X1 U944 ( .A1(G234), .A2(G237), .ZN(n1243) );
NOR3_X1 U945 ( .A1(n1238), .A2(n1067), .A3(n1078), .ZN(n1222) );
INV_X1 U946 ( .A(n1258), .ZN(n1078) );
NOR2_X1 U947 ( .A1(n1081), .A2(n1103), .ZN(n1258) );
INV_X1 U948 ( .A(n1082), .ZN(n1103) );
NAND2_X1 U949 ( .A1(G214), .A2(n1261), .ZN(n1082) );
NOR2_X1 U950 ( .A1(n1102), .A2(n1262), .ZN(n1081) );
NOR2_X1 U951 ( .A1(n1100), .A2(n1101), .ZN(n1262) );
AND2_X1 U952 ( .A1(n1101), .A2(n1100), .ZN(n1102) );
NAND2_X1 U953 ( .A1(G210), .A2(n1261), .ZN(n1100) );
NAND2_X1 U954 ( .A1(n1263), .A2(n1264), .ZN(n1261) );
NOR2_X1 U955 ( .A1(n1224), .A2(G902), .ZN(n1101) );
XOR2_X1 U956 ( .A(n1265), .B(n1266), .Z(n1224) );
XOR2_X1 U957 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U958 ( .A(G143), .B(G125), .Z(n1268) );
AND2_X1 U959 ( .A1(n1042), .A2(G224), .ZN(n1267) );
XOR2_X1 U960 ( .A(n1134), .B(n1269), .Z(n1265) );
INV_X1 U961 ( .A(n1171), .ZN(n1269) );
XOR2_X1 U962 ( .A(n1270), .B(n1271), .Z(n1134) );
XOR2_X1 U963 ( .A(G110), .B(G107), .Z(n1271) );
XOR2_X1 U964 ( .A(n1272), .B(n1273), .Z(n1270) );
NAND2_X1 U965 ( .A1(n1274), .A2(n1275), .ZN(n1272) );
OR2_X1 U966 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XOR2_X1 U967 ( .A(n1278), .B(KEYINPUT44), .Z(n1274) );
NAND2_X1 U968 ( .A1(n1276), .A2(n1277), .ZN(n1278) );
INV_X1 U969 ( .A(G113), .ZN(n1277) );
XNOR2_X1 U970 ( .A(n1279), .B(G119), .ZN(n1276) );
NAND2_X1 U971 ( .A1(KEYINPUT50), .A2(n1280), .ZN(n1279) );
AND2_X1 U972 ( .A1(G221), .A2(n1281), .ZN(n1067) );
INV_X1 U973 ( .A(n1068), .ZN(n1238) );
XNOR2_X1 U974 ( .A(n1282), .B(n1094), .ZN(n1068) );
NAND2_X1 U975 ( .A1(n1283), .A2(n1284), .ZN(n1094) );
XOR2_X1 U976 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U977 ( .A(n1191), .B(n1287), .ZN(n1286) );
NAND2_X1 U978 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U979 ( .A1(n1290), .A2(n1189), .ZN(n1289) );
XOR2_X1 U980 ( .A(KEYINPUT45), .B(n1291), .Z(n1288) );
NOR2_X1 U981 ( .A1(n1290), .A2(n1189), .ZN(n1291) );
XOR2_X1 U982 ( .A(n1171), .B(n1292), .Z(n1290) );
XOR2_X1 U983 ( .A(n1187), .B(n1183), .Z(n1292) );
XNOR2_X1 U984 ( .A(KEYINPUT54), .B(n1293), .ZN(n1183) );
NOR2_X1 U985 ( .A1(KEYINPUT1), .A2(n1294), .ZN(n1293) );
XOR2_X1 U986 ( .A(n1229), .B(KEYINPUT9), .Z(n1294) );
NAND3_X1 U987 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1187) );
OR2_X1 U988 ( .A1(n1298), .A2(G107), .ZN(n1297) );
NAND2_X1 U989 ( .A1(n1299), .A2(n1300), .ZN(n1296) );
INV_X1 U990 ( .A(KEYINPUT14), .ZN(n1300) );
NAND2_X1 U991 ( .A1(n1301), .A2(n1298), .ZN(n1299) );
XNOR2_X1 U992 ( .A(KEYINPUT39), .B(G107), .ZN(n1301) );
NAND2_X1 U993 ( .A1(KEYINPUT14), .A2(n1302), .ZN(n1295) );
NAND2_X1 U994 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
OR2_X1 U995 ( .A1(G107), .A2(KEYINPUT39), .ZN(n1304) );
NAND3_X1 U996 ( .A1(G107), .A2(n1298), .A3(KEYINPUT39), .ZN(n1303) );
XNOR2_X1 U997 ( .A(G104), .B(KEYINPUT2), .ZN(n1298) );
XOR2_X1 U998 ( .A(n1190), .B(n1184), .Z(n1171) );
INV_X1 U999 ( .A(G101), .ZN(n1190) );
NOR2_X1 U1000 ( .A1(n1110), .A2(G953), .ZN(n1191) );
INV_X1 U1001 ( .A(G227), .ZN(n1110) );
NOR3_X1 U1002 ( .A1(KEYINPUT43), .A2(n1305), .A3(n1306), .ZN(n1285) );
NOR3_X1 U1003 ( .A1(KEYINPUT60), .A2(G110), .A3(n1307), .ZN(n1306) );
NOR2_X1 U1004 ( .A1(n1179), .A2(n1308), .ZN(n1305) );
INV_X1 U1005 ( .A(KEYINPUT60), .ZN(n1308) );
XNOR2_X1 U1006 ( .A(n1259), .B(G140), .ZN(n1179) );
XOR2_X1 U1007 ( .A(KEYINPUT24), .B(G902), .Z(n1283) );
NAND2_X1 U1008 ( .A1(KEYINPUT20), .A2(n1093), .ZN(n1282) );
INV_X1 U1009 ( .A(G469), .ZN(n1093) );
NOR2_X1 U1010 ( .A1(n1104), .A2(n1245), .ZN(n1066) );
XOR2_X1 U1011 ( .A(n1099), .B(n1309), .Z(n1245) );
NOR2_X1 U1012 ( .A1(G478), .A2(KEYINPUT30), .ZN(n1309) );
OR2_X1 U1013 ( .A1(n1147), .A2(G902), .ZN(n1099) );
XNOR2_X1 U1014 ( .A(n1310), .B(n1311), .ZN(n1147) );
XNOR2_X1 U1015 ( .A(n1312), .B(n1313), .ZN(n1311) );
XOR2_X1 U1016 ( .A(n1314), .B(n1315), .Z(n1313) );
NOR2_X1 U1017 ( .A1(KEYINPUT15), .A2(n1316), .ZN(n1315) );
XOR2_X1 U1018 ( .A(KEYINPUT57), .B(G128), .Z(n1316) );
NAND2_X1 U1019 ( .A1(G217), .A2(n1317), .ZN(n1314) );
XNOR2_X1 U1020 ( .A(G107), .B(n1318), .ZN(n1310) );
XOR2_X1 U1021 ( .A(G134), .B(G122), .Z(n1318) );
INV_X1 U1022 ( .A(n1234), .ZN(n1104) );
XOR2_X1 U1023 ( .A(n1319), .B(G475), .Z(n1234) );
NAND2_X1 U1024 ( .A1(n1264), .A2(n1157), .ZN(n1319) );
NAND2_X1 U1025 ( .A1(n1320), .A2(n1321), .ZN(n1157) );
NAND2_X1 U1026 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XOR2_X1 U1027 ( .A(KEYINPUT3), .B(n1324), .Z(n1320) );
NOR2_X1 U1028 ( .A1(n1323), .A2(n1322), .ZN(n1324) );
XOR2_X1 U1029 ( .A(G113), .B(n1273), .Z(n1322) );
XOR2_X1 U1030 ( .A(G104), .B(G122), .Z(n1273) );
XOR2_X1 U1031 ( .A(n1325), .B(n1326), .Z(n1323) );
XOR2_X1 U1032 ( .A(n1327), .B(n1328), .Z(n1326) );
NOR2_X1 U1033 ( .A1(G131), .A2(KEYINPUT10), .ZN(n1328) );
AND2_X1 U1034 ( .A1(n1329), .A2(G214), .ZN(n1327) );
NAND2_X1 U1035 ( .A1(n1330), .A2(n1331), .ZN(n1325) );
NAND2_X1 U1036 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
INV_X1 U1037 ( .A(KEYINPUT33), .ZN(n1333) );
XOR2_X1 U1038 ( .A(n1334), .B(n1118), .Z(n1332) );
XOR2_X1 U1039 ( .A(G125), .B(G140), .Z(n1118) );
NAND2_X1 U1040 ( .A1(KEYINPUT33), .A2(n1335), .ZN(n1330) );
XOR2_X1 U1041 ( .A(n1240), .B(n1334), .Z(n1335) );
XOR2_X1 U1042 ( .A(G143), .B(G146), .Z(n1334) );
INV_X1 U1043 ( .A(G125), .ZN(n1240) );
INV_X1 U1044 ( .A(n1051), .ZN(n1076) );
NAND2_X1 U1045 ( .A1(n1252), .A2(n1246), .ZN(n1051) );
NAND2_X1 U1046 ( .A1(n1092), .A2(n1085), .ZN(n1246) );
NAND3_X1 U1047 ( .A1(n1336), .A2(n1264), .A3(n1143), .ZN(n1085) );
NAND2_X1 U1048 ( .A1(G217), .A2(n1337), .ZN(n1336) );
NAND2_X1 U1049 ( .A1(n1145), .A2(n1338), .ZN(n1092) );
NAND2_X1 U1050 ( .A1(n1143), .A2(n1264), .ZN(n1338) );
XOR2_X1 U1051 ( .A(n1339), .B(n1340), .Z(n1143) );
XOR2_X1 U1052 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1053 ( .A(G146), .B(G110), .Z(n1342) );
NOR2_X1 U1054 ( .A1(KEYINPUT37), .A2(n1343), .ZN(n1341) );
XOR2_X1 U1055 ( .A(n1344), .B(G128), .Z(n1343) );
INV_X1 U1056 ( .A(G119), .ZN(n1344) );
XOR2_X1 U1057 ( .A(n1345), .B(n1346), .Z(n1339) );
NOR2_X1 U1058 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
NOR3_X1 U1059 ( .A1(G140), .A2(G125), .A3(n1349), .ZN(n1348) );
NOR2_X1 U1060 ( .A1(n1350), .A2(n1307), .ZN(n1347) );
INV_X1 U1061 ( .A(G140), .ZN(n1307) );
NOR2_X1 U1062 ( .A1(G125), .A2(n1349), .ZN(n1350) );
INV_X1 U1063 ( .A(KEYINPUT41), .ZN(n1349) );
NAND4_X1 U1064 ( .A1(n1351), .A2(n1352), .A3(n1353), .A4(n1354), .ZN(n1345) );
NAND3_X1 U1065 ( .A1(KEYINPUT49), .A2(n1355), .A3(n1356), .ZN(n1354) );
XOR2_X1 U1066 ( .A(n1357), .B(KEYINPUT27), .Z(n1355) );
OR2_X1 U1067 ( .A1(n1356), .A2(KEYINPUT49), .ZN(n1353) );
OR3_X1 U1068 ( .A1(n1357), .A2(n1358), .A3(KEYINPUT62), .ZN(n1352) );
NOR2_X1 U1069 ( .A1(KEYINPUT27), .A2(G137), .ZN(n1358) );
NAND3_X1 U1070 ( .A1(n1359), .A2(n1357), .A3(KEYINPUT62), .ZN(n1351) );
NAND2_X1 U1071 ( .A1(G221), .A2(n1317), .ZN(n1357) );
NOR2_X1 U1072 ( .A1(n1337), .A2(G953), .ZN(n1317) );
INV_X1 U1073 ( .A(G234), .ZN(n1337) );
NAND2_X1 U1074 ( .A1(KEYINPUT27), .A2(n1356), .ZN(n1359) );
INV_X1 U1075 ( .A(G137), .ZN(n1356) );
AND2_X1 U1076 ( .A1(G217), .A2(n1281), .ZN(n1145) );
NAND2_X1 U1077 ( .A1(G234), .A2(n1264), .ZN(n1281) );
XNOR2_X1 U1078 ( .A(G472), .B(n1360), .ZN(n1252) );
NOR2_X1 U1079 ( .A1(KEYINPUT5), .A2(n1095), .ZN(n1360) );
NAND2_X1 U1080 ( .A1(n1361), .A2(n1264), .ZN(n1095) );
INV_X1 U1081 ( .A(G902), .ZN(n1264) );
XOR2_X1 U1082 ( .A(n1362), .B(n1363), .Z(n1361) );
XOR2_X1 U1083 ( .A(KEYINPUT26), .B(n1364), .Z(n1363) );
NOR2_X1 U1084 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
XOR2_X1 U1085 ( .A(KEYINPUT7), .B(KEYINPUT0), .Z(n1366) );
XOR2_X1 U1086 ( .A(n1175), .B(n1367), .Z(n1365) );
XOR2_X1 U1087 ( .A(KEYINPUT23), .B(G101), .Z(n1367) );
NAND2_X1 U1088 ( .A1(G210), .A2(n1329), .ZN(n1175) );
AND2_X1 U1089 ( .A1(n1368), .A2(n1042), .ZN(n1329) );
INV_X1 U1090 ( .A(G953), .ZN(n1042) );
XOR2_X1 U1091 ( .A(n1263), .B(KEYINPUT52), .Z(n1368) );
INV_X1 U1092 ( .A(G237), .ZN(n1263) );
XOR2_X1 U1093 ( .A(n1170), .B(n1184), .Z(n1362) );
XOR2_X1 U1094 ( .A(G128), .B(G146), .Z(n1184) );
XOR2_X1 U1095 ( .A(n1369), .B(n1370), .Z(n1170) );
XOR2_X1 U1096 ( .A(G119), .B(G113), .Z(n1370) );
XNOR2_X1 U1097 ( .A(n1189), .B(n1312), .ZN(n1369) );
XOR2_X1 U1098 ( .A(n1280), .B(n1229), .Z(n1312) );
INV_X1 U1099 ( .A(G143), .ZN(n1229) );
INV_X1 U1100 ( .A(G116), .ZN(n1280) );
XOR2_X1 U1101 ( .A(G131), .B(n1371), .Z(n1189) );
NOR2_X1 U1102 ( .A1(KEYINPUT59), .A2(n1372), .ZN(n1371) );
NOR2_X1 U1103 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
XOR2_X1 U1104 ( .A(n1375), .B(KEYINPUT19), .Z(n1374) );
NAND2_X1 U1105 ( .A1(G134), .A2(n1376), .ZN(n1375) );
NOR2_X1 U1106 ( .A1(G134), .A2(n1376), .ZN(n1373) );
XOR2_X1 U1107 ( .A(G137), .B(KEYINPUT12), .Z(n1376) );
INV_X1 U1108 ( .A(G110), .ZN(n1259) );
endmodule


