//Key = 1110000110010011111100010100110111010110001110110000011000000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315;

NAND2_X1 U726 ( .A1(n1003), .A2(n1004), .ZN(G9) );
NAND2_X1 U727 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
XOR2_X1 U728 ( .A(KEYINPUT2), .B(n1007), .Z(n1003) );
NOR2_X1 U729 ( .A1(n1005), .A2(n1006), .ZN(n1007) );
INV_X1 U730 ( .A(n1008), .ZN(n1005) );
NOR2_X1 U731 ( .A1(n1009), .A2(n1010), .ZN(G75) );
NOR4_X1 U732 ( .A1(G953), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1010) );
NOR2_X1 U733 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR2_X1 U734 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR3_X1 U735 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1017) );
NOR2_X1 U736 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
AND2_X1 U737 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR3_X1 U738 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1021) );
NOR3_X1 U739 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
NOR2_X1 U740 ( .A1(n1023), .A2(n1031), .ZN(n1026) );
NOR4_X1 U741 ( .A1(n1028), .A2(n1032), .A3(n1033), .A4(n1025), .ZN(n1016) );
INV_X1 U742 ( .A(n1023), .ZN(n1033) );
NOR4_X1 U743 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1032) );
AND2_X1 U744 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR3_X1 U745 ( .A1(n1040), .A2(KEYINPUT54), .A3(n1041), .ZN(n1035) );
NOR2_X1 U746 ( .A1(n1042), .A2(n1020), .ZN(n1034) );
INV_X1 U747 ( .A(n1040), .ZN(n1020) );
NOR2_X1 U748 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
XOR2_X1 U749 ( .A(KEYINPUT30), .B(n1045), .Z(n1044) );
NOR2_X1 U750 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
AND2_X1 U751 ( .A1(n1048), .A2(KEYINPUT54), .ZN(n1043) );
NOR3_X1 U752 ( .A1(n1011), .A2(G953), .A3(G952), .ZN(n1009) );
AND4_X1 U753 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1011) );
NOR3_X1 U754 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
INV_X1 U755 ( .A(n1056), .ZN(n1055) );
NAND3_X1 U756 ( .A1(n1057), .A2(n1058), .A3(n1031), .ZN(n1053) );
NOR3_X1 U757 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1051) );
XNOR2_X1 U758 ( .A(n1062), .B(KEYINPUT18), .ZN(n1061) );
INV_X1 U759 ( .A(n1046), .ZN(n1060) );
XOR2_X1 U760 ( .A(n1063), .B(n1064), .Z(n1049) );
XOR2_X1 U761 ( .A(KEYINPUT19), .B(n1065), .Z(n1064) );
NOR2_X1 U762 ( .A1(KEYINPUT20), .A2(G478), .ZN(n1065) );
XOR2_X1 U763 ( .A(n1066), .B(n1067), .Z(G72) );
NOR2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NAND2_X1 U766 ( .A1(n1072), .A2(n1073), .ZN(n1066) );
NAND3_X1 U767 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
NAND2_X1 U768 ( .A1(G953), .A2(n1071), .ZN(n1075) );
OR2_X1 U769 ( .A1(n1076), .A2(n1074), .ZN(n1072) );
XNOR2_X1 U770 ( .A(n1077), .B(n1078), .ZN(n1074) );
XNOR2_X1 U771 ( .A(G131), .B(n1079), .ZN(n1078) );
XNOR2_X1 U772 ( .A(KEYINPUT57), .B(KEYINPUT55), .ZN(n1079) );
XOR2_X1 U773 ( .A(n1080), .B(n1081), .Z(n1077) );
XOR2_X1 U774 ( .A(n1082), .B(n1083), .Z(n1080) );
NAND2_X1 U775 ( .A1(n1069), .A2(n1084), .ZN(n1076) );
NAND4_X1 U776 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1084) );
NOR2_X1 U777 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XOR2_X1 U778 ( .A(n1091), .B(KEYINPUT46), .Z(n1089) );
XOR2_X1 U779 ( .A(n1092), .B(n1093), .Z(G69) );
XOR2_X1 U780 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U781 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XNOR2_X1 U782 ( .A(n1098), .B(n1099), .ZN(n1097) );
NOR2_X1 U783 ( .A1(n1069), .A2(n1100), .ZN(n1096) );
XNOR2_X1 U784 ( .A(KEYINPUT12), .B(n1101), .ZN(n1100) );
NAND2_X1 U785 ( .A1(n1069), .A2(n1102), .ZN(n1094) );
NAND2_X1 U786 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U787 ( .A(KEYINPUT28), .B(n1008), .ZN(n1104) );
NAND3_X1 U788 ( .A1(G953), .A2(n1105), .A3(KEYINPUT47), .ZN(n1092) );
XOR2_X1 U789 ( .A(KEYINPUT43), .B(n1106), .Z(n1105) );
AND2_X1 U790 ( .A1(G224), .A2(G898), .ZN(n1106) );
NOR2_X1 U791 ( .A1(n1107), .A2(n1108), .ZN(G66) );
NOR2_X1 U792 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U793 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U794 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U795 ( .A1(KEYINPUT26), .A2(n1115), .ZN(n1111) );
AND2_X1 U796 ( .A1(n1115), .A2(KEYINPUT26), .ZN(n1109) );
NOR2_X1 U797 ( .A1(n1107), .A2(n1116), .ZN(G63) );
XOR2_X1 U798 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND3_X1 U799 ( .A1(n1119), .A2(n1013), .A3(G478), .ZN(n1118) );
XNOR2_X1 U800 ( .A(KEYINPUT50), .B(n1120), .ZN(n1119) );
NOR2_X1 U801 ( .A1(n1107), .A2(n1121), .ZN(G60) );
XOR2_X1 U802 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U803 ( .A1(KEYINPUT56), .A2(n1124), .ZN(n1123) );
NAND2_X1 U804 ( .A1(n1125), .A2(G475), .ZN(n1122) );
XNOR2_X1 U805 ( .A(G104), .B(n1126), .ZN(G6) );
NOR2_X1 U806 ( .A1(n1107), .A2(n1127), .ZN(G57) );
XOR2_X1 U807 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U808 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U809 ( .A1(KEYINPUT13), .A2(n1132), .ZN(n1131) );
XNOR2_X1 U810 ( .A(KEYINPUT31), .B(n1133), .ZN(n1132) );
NOR2_X1 U811 ( .A1(KEYINPUT58), .A2(n1134), .ZN(n1130) );
XNOR2_X1 U812 ( .A(n1135), .B(n1136), .ZN(n1134) );
XOR2_X1 U813 ( .A(n1137), .B(n1138), .Z(n1128) );
AND2_X1 U814 ( .A1(G472), .A2(n1125), .ZN(n1138) );
NOR2_X1 U815 ( .A1(n1107), .A2(n1139), .ZN(G54) );
XOR2_X1 U816 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U817 ( .A(n1142), .B(n1143), .ZN(n1141) );
AND2_X1 U818 ( .A1(G469), .A2(n1125), .ZN(n1142) );
INV_X1 U819 ( .A(n1114), .ZN(n1125) );
XOR2_X1 U820 ( .A(n1144), .B(n1145), .Z(n1140) );
NOR2_X1 U821 ( .A1(KEYINPUT5), .A2(n1146), .ZN(n1144) );
NOR2_X1 U822 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U823 ( .A(n1149), .B(KEYINPUT15), .Z(n1148) );
NAND2_X1 U824 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NOR2_X1 U825 ( .A1(n1151), .A2(n1150), .ZN(n1147) );
XOR2_X1 U826 ( .A(n1152), .B(KEYINPUT40), .Z(n1150) );
NOR2_X1 U827 ( .A1(n1107), .A2(n1153), .ZN(G51) );
XOR2_X1 U828 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U829 ( .A1(n1156), .A2(n1114), .ZN(n1155) );
NAND2_X1 U830 ( .A1(G902), .A2(n1013), .ZN(n1114) );
NAND4_X1 U831 ( .A1(n1157), .A2(n1091), .A3(n1103), .A4(n1158), .ZN(n1013) );
AND4_X1 U832 ( .A1(n1086), .A2(n1085), .A3(n1008), .A4(n1087), .ZN(n1158) );
NAND3_X1 U833 ( .A1(n1040), .A2(n1159), .A3(n1029), .ZN(n1008) );
AND4_X1 U834 ( .A1(n1160), .A2(n1161), .A3(n1126), .A4(n1162), .ZN(n1103) );
AND4_X1 U835 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1162) );
NAND3_X1 U836 ( .A1(n1040), .A2(n1159), .A3(n1030), .ZN(n1126) );
NAND2_X1 U837 ( .A1(n1048), .A2(n1167), .ZN(n1091) );
XOR2_X1 U838 ( .A(KEYINPUT27), .B(n1168), .Z(n1167) );
XNOR2_X1 U839 ( .A(KEYINPUT59), .B(n1090), .ZN(n1157) );
NAND4_X1 U840 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1090) );
NOR3_X1 U841 ( .A1(n1173), .A2(KEYINPUT52), .A3(n1174), .ZN(n1154) );
NOR2_X1 U842 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XOR2_X1 U843 ( .A(KEYINPUT51), .B(n1177), .Z(n1173) );
NOR2_X1 U844 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XNOR2_X1 U845 ( .A(n1180), .B(KEYINPUT61), .ZN(n1179) );
INV_X1 U846 ( .A(n1176), .ZN(n1178) );
NAND2_X1 U847 ( .A1(n1181), .A2(n1182), .ZN(n1176) );
XOR2_X1 U848 ( .A(n1183), .B(KEYINPUT45), .Z(n1181) );
NOR2_X1 U849 ( .A1(n1069), .A2(G952), .ZN(n1107) );
XNOR2_X1 U850 ( .A(G146), .B(n1184), .ZN(G48) );
NAND2_X1 U851 ( .A1(n1168), .A2(n1048), .ZN(n1184) );
AND2_X1 U852 ( .A1(n1030), .A2(n1185), .ZN(n1168) );
XNOR2_X1 U853 ( .A(G143), .B(n1087), .ZN(G45) );
NAND3_X1 U854 ( .A1(n1186), .A2(n1048), .A3(n1187), .ZN(n1087) );
XOR2_X1 U855 ( .A(n1085), .B(n1188), .Z(G42) );
XOR2_X1 U856 ( .A(KEYINPUT38), .B(G140), .Z(n1188) );
NAND4_X1 U857 ( .A1(n1030), .A2(n1036), .A3(n1024), .A4(n1189), .ZN(n1085) );
NOR3_X1 U858 ( .A1(n1062), .A2(n1190), .A3(n1018), .ZN(n1036) );
INV_X1 U859 ( .A(n1038), .ZN(n1018) );
XNOR2_X1 U860 ( .A(G137), .B(n1086), .ZN(G39) );
NAND3_X1 U861 ( .A1(n1038), .A2(n1023), .A3(n1185), .ZN(n1086) );
XNOR2_X1 U862 ( .A(G134), .B(n1191), .ZN(G36) );
NOR2_X1 U863 ( .A1(n1192), .A2(KEYINPUT62), .ZN(n1191) );
INV_X1 U864 ( .A(n1169), .ZN(n1192) );
NAND3_X1 U865 ( .A1(n1038), .A2(n1029), .A3(n1187), .ZN(n1169) );
XNOR2_X1 U866 ( .A(n1170), .B(n1193), .ZN(G33) );
NOR2_X1 U867 ( .A1(KEYINPUT22), .A2(n1194), .ZN(n1193) );
NAND3_X1 U868 ( .A1(n1030), .A2(n1038), .A3(n1187), .ZN(n1170) );
AND3_X1 U869 ( .A1(n1024), .A2(n1189), .A3(n1039), .ZN(n1187) );
NOR2_X1 U870 ( .A1(n1047), .A2(n1195), .ZN(n1038) );
INV_X1 U871 ( .A(n1196), .ZN(n1195) );
XNOR2_X1 U872 ( .A(G128), .B(n1171), .ZN(G30) );
NAND3_X1 U873 ( .A1(n1029), .A2(n1048), .A3(n1185), .ZN(n1171) );
AND4_X1 U874 ( .A1(n1197), .A2(n1024), .A3(n1062), .A4(n1189), .ZN(n1185) );
XNOR2_X1 U875 ( .A(G101), .B(n1160), .ZN(G3) );
NAND3_X1 U876 ( .A1(n1159), .A2(n1023), .A3(n1039), .ZN(n1160) );
XNOR2_X1 U877 ( .A(G125), .B(n1172), .ZN(G27) );
NAND4_X1 U878 ( .A1(n1197), .A2(n1030), .A3(n1198), .A4(n1199), .ZN(n1172) );
AND4_X1 U879 ( .A1(n1031), .A2(n1189), .A3(n1048), .A4(n1200), .ZN(n1199) );
NAND2_X1 U880 ( .A1(n1015), .A2(n1201), .ZN(n1189) );
NAND4_X1 U881 ( .A1(G953), .A2(G902), .A3(n1202), .A4(n1071), .ZN(n1201) );
INV_X1 U882 ( .A(G900), .ZN(n1071) );
XNOR2_X1 U883 ( .A(G122), .B(n1161), .ZN(G24) );
NAND3_X1 U884 ( .A1(n1203), .A2(n1040), .A3(n1186), .ZN(n1161) );
AND2_X1 U885 ( .A1(n1204), .A2(n1205), .ZN(n1186) );
XOR2_X1 U886 ( .A(KEYINPUT4), .B(n1059), .Z(n1204) );
NOR2_X1 U887 ( .A1(n1062), .A2(n1197), .ZN(n1040) );
XOR2_X1 U888 ( .A(n1165), .B(n1206), .Z(G21) );
NOR2_X1 U889 ( .A1(G119), .A2(KEYINPUT36), .ZN(n1206) );
NAND4_X1 U890 ( .A1(n1197), .A2(n1203), .A3(n1023), .A4(n1062), .ZN(n1165) );
XNOR2_X1 U891 ( .A(G116), .B(n1207), .ZN(G18) );
NAND2_X1 U892 ( .A1(KEYINPUT16), .A2(n1208), .ZN(n1207) );
INV_X1 U893 ( .A(n1164), .ZN(n1208) );
NAND3_X1 U894 ( .A1(n1203), .A2(n1029), .A3(n1039), .ZN(n1164) );
XNOR2_X1 U895 ( .A(G113), .B(n1163), .ZN(G15) );
NAND3_X1 U896 ( .A1(n1203), .A2(n1030), .A3(n1039), .ZN(n1163) );
NOR2_X1 U897 ( .A1(n1197), .A2(n1200), .ZN(n1039) );
AND2_X1 U898 ( .A1(n1209), .A2(n1059), .ZN(n1030) );
XNOR2_X1 U899 ( .A(KEYINPUT0), .B(n1210), .ZN(n1209) );
AND3_X1 U900 ( .A1(n1211), .A2(n1031), .A3(n1198), .ZN(n1203) );
XNOR2_X1 U901 ( .A(G110), .B(n1166), .ZN(G12) );
NAND4_X1 U902 ( .A1(n1197), .A2(n1159), .A3(n1200), .A4(n1023), .ZN(n1166) );
NAND2_X1 U903 ( .A1(n1212), .A2(n1213), .ZN(n1023) );
NAND2_X1 U904 ( .A1(n1029), .A2(n1214), .ZN(n1213) );
NOR2_X1 U905 ( .A1(n1059), .A2(n1210), .ZN(n1029) );
INV_X1 U906 ( .A(n1205), .ZN(n1210) );
OR3_X1 U907 ( .A1(n1059), .A2(n1205), .A3(n1214), .ZN(n1212) );
INV_X1 U908 ( .A(KEYINPUT0), .ZN(n1214) );
XNOR2_X1 U909 ( .A(n1063), .B(G478), .ZN(n1205) );
NAND2_X1 U910 ( .A1(n1120), .A2(n1117), .ZN(n1063) );
NAND2_X1 U911 ( .A1(n1215), .A2(n1216), .ZN(n1117) );
NAND4_X1 U912 ( .A1(G217), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1216) );
NAND2_X1 U913 ( .A1(n1220), .A2(n1221), .ZN(n1215) );
NAND2_X1 U914 ( .A1(G217), .A2(n1217), .ZN(n1221) );
NAND2_X1 U915 ( .A1(n1218), .A2(n1219), .ZN(n1220) );
NAND2_X1 U916 ( .A1(n1222), .A2(n1223), .ZN(n1219) );
XNOR2_X1 U917 ( .A(n1224), .B(KEYINPUT23), .ZN(n1218) );
OR2_X1 U918 ( .A1(n1223), .A2(n1222), .ZN(n1224) );
XOR2_X1 U919 ( .A(n1006), .B(n1225), .Z(n1222) );
XNOR2_X1 U920 ( .A(n1226), .B(G116), .ZN(n1225) );
XOR2_X1 U921 ( .A(G128), .B(n1227), .Z(n1223) );
XOR2_X1 U922 ( .A(G143), .B(G134), .Z(n1227) );
XNOR2_X1 U923 ( .A(n1228), .B(G475), .ZN(n1059) );
OR2_X1 U924 ( .A1(n1124), .A2(G902), .ZN(n1228) );
XNOR2_X1 U925 ( .A(n1229), .B(n1230), .ZN(n1124) );
XOR2_X1 U926 ( .A(n1231), .B(n1232), .Z(n1230) );
XNOR2_X1 U927 ( .A(n1233), .B(n1234), .ZN(n1232) );
NAND2_X1 U928 ( .A1(G214), .A2(n1235), .ZN(n1233) );
XNOR2_X1 U929 ( .A(G113), .B(G131), .ZN(n1231) );
XOR2_X1 U930 ( .A(n1236), .B(n1081), .Z(n1229) );
XNOR2_X1 U931 ( .A(n1237), .B(n1238), .ZN(n1236) );
NAND2_X1 U932 ( .A1(KEYINPUT7), .A2(n1226), .ZN(n1237) );
INV_X1 U933 ( .A(n1062), .ZN(n1200) );
XNOR2_X1 U934 ( .A(n1239), .B(G472), .ZN(n1062) );
NAND2_X1 U935 ( .A1(n1240), .A2(n1120), .ZN(n1239) );
XOR2_X1 U936 ( .A(n1241), .B(n1242), .Z(n1240) );
NOR2_X1 U937 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XOR2_X1 U938 ( .A(n1245), .B(KEYINPUT37), .Z(n1244) );
NAND2_X1 U939 ( .A1(n1246), .A2(n1136), .ZN(n1245) );
XOR2_X1 U940 ( .A(KEYINPUT49), .B(n1135), .Z(n1246) );
NOR2_X1 U941 ( .A1(n1247), .A2(n1135), .ZN(n1243) );
XNOR2_X1 U942 ( .A(n1248), .B(n1151), .ZN(n1135) );
INV_X1 U943 ( .A(n1249), .ZN(n1151) );
XNOR2_X1 U944 ( .A(n1136), .B(KEYINPUT14), .ZN(n1247) );
XNOR2_X1 U945 ( .A(n1250), .B(n1251), .ZN(n1136) );
NOR2_X1 U946 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
XOR2_X1 U947 ( .A(KEYINPUT6), .B(n1254), .Z(n1253) );
NOR2_X1 U948 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XNOR2_X1 U949 ( .A(KEYINPUT29), .B(n1257), .ZN(n1256) );
INV_X1 U950 ( .A(G116), .ZN(n1257) );
NOR2_X1 U951 ( .A1(KEYINPUT3), .A2(n1258), .ZN(n1241) );
XOR2_X1 U952 ( .A(n1137), .B(n1259), .Z(n1258) );
XNOR2_X1 U953 ( .A(KEYINPUT39), .B(n1133), .ZN(n1259) );
NAND2_X1 U954 ( .A1(G210), .A2(n1235), .ZN(n1137) );
NOR2_X1 U955 ( .A1(G953), .A2(G237), .ZN(n1235) );
AND2_X1 U956 ( .A1(n1024), .A2(n1211), .ZN(n1159) );
AND2_X1 U957 ( .A1(n1048), .A2(n1260), .ZN(n1211) );
NAND2_X1 U958 ( .A1(n1015), .A2(n1261), .ZN(n1260) );
NAND4_X1 U959 ( .A1(G953), .A2(G902), .A3(n1202), .A4(n1101), .ZN(n1261) );
INV_X1 U960 ( .A(G898), .ZN(n1101) );
NAND3_X1 U961 ( .A1(n1202), .A2(n1069), .A3(G952), .ZN(n1015) );
NAND2_X1 U962 ( .A1(G237), .A2(G234), .ZN(n1202) );
INV_X1 U963 ( .A(n1041), .ZN(n1048) );
NAND2_X1 U964 ( .A1(n1196), .A2(n1047), .ZN(n1041) );
NAND3_X1 U965 ( .A1(n1262), .A2(n1263), .A3(n1056), .ZN(n1047) );
NAND3_X1 U966 ( .A1(n1156), .A2(n1120), .A3(n1264), .ZN(n1056) );
NAND2_X1 U967 ( .A1(n1156), .A2(n1265), .ZN(n1263) );
INV_X1 U968 ( .A(KEYINPUT1), .ZN(n1265) );
NAND2_X1 U969 ( .A1(n1054), .A2(KEYINPUT1), .ZN(n1262) );
NOR2_X1 U970 ( .A1(n1156), .A2(n1266), .ZN(n1054) );
AND2_X1 U971 ( .A1(n1264), .A2(n1120), .ZN(n1266) );
XNOR2_X1 U972 ( .A(n1267), .B(n1175), .ZN(n1264) );
INV_X1 U973 ( .A(n1180), .ZN(n1175) );
XOR2_X1 U974 ( .A(n1099), .B(n1268), .Z(n1180) );
NOR2_X1 U975 ( .A1(KEYINPUT48), .A2(n1098), .ZN(n1268) );
XNOR2_X1 U976 ( .A(n1269), .B(n1270), .ZN(n1098) );
XNOR2_X1 U977 ( .A(G107), .B(n1271), .ZN(n1270) );
NAND2_X1 U978 ( .A1(KEYINPUT8), .A2(n1234), .ZN(n1271) );
INV_X1 U979 ( .A(G104), .ZN(n1234) );
NAND2_X1 U980 ( .A1(KEYINPUT25), .A2(n1133), .ZN(n1269) );
INV_X1 U981 ( .A(G101), .ZN(n1133) );
XNOR2_X1 U982 ( .A(n1272), .B(n1273), .ZN(n1099) );
XOR2_X1 U983 ( .A(n1274), .B(n1250), .Z(n1273) );
XNOR2_X1 U984 ( .A(G113), .B(KEYINPUT11), .ZN(n1250) );
NAND2_X1 U985 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
INV_X1 U986 ( .A(n1252), .ZN(n1276) );
NOR2_X1 U987 ( .A1(n1277), .A2(G116), .ZN(n1252) );
XOR2_X1 U988 ( .A(n1278), .B(KEYINPUT34), .Z(n1275) );
NAND2_X1 U989 ( .A1(n1277), .A2(G116), .ZN(n1278) );
INV_X1 U990 ( .A(n1255), .ZN(n1277) );
XNOR2_X1 U991 ( .A(G110), .B(n1279), .ZN(n1272) );
XNOR2_X1 U992 ( .A(KEYINPUT42), .B(n1226), .ZN(n1279) );
INV_X1 U993 ( .A(G122), .ZN(n1226) );
NAND2_X1 U994 ( .A1(n1183), .A2(n1182), .ZN(n1267) );
NAND2_X1 U995 ( .A1(n1280), .A2(n1281), .ZN(n1182) );
NAND2_X1 U996 ( .A1(G224), .A2(n1069), .ZN(n1281) );
XOR2_X1 U997 ( .A(G125), .B(n1248), .Z(n1280) );
NAND3_X1 U998 ( .A1(G224), .A2(n1069), .A3(n1282), .ZN(n1183) );
XNOR2_X1 U999 ( .A(n1248), .B(G125), .ZN(n1282) );
XNOR2_X1 U1000 ( .A(G128), .B(n1238), .ZN(n1248) );
NAND2_X1 U1001 ( .A1(G210), .A2(n1283), .ZN(n1156) );
XNOR2_X1 U1002 ( .A(n1046), .B(KEYINPUT44), .ZN(n1196) );
NAND2_X1 U1003 ( .A1(G214), .A2(n1283), .ZN(n1046) );
NAND2_X1 U1004 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
INV_X1 U1005 ( .A(G237), .ZN(n1285) );
NOR2_X1 U1006 ( .A1(n1028), .A2(n1198), .ZN(n1024) );
INV_X1 U1007 ( .A(n1025), .ZN(n1198) );
NAND2_X1 U1008 ( .A1(n1286), .A2(n1057), .ZN(n1025) );
NAND2_X1 U1009 ( .A1(G469), .A2(n1287), .ZN(n1057) );
XNOR2_X1 U1010 ( .A(KEYINPUT17), .B(n1058), .ZN(n1286) );
OR2_X1 U1011 ( .A1(n1287), .A2(G469), .ZN(n1058) );
NAND2_X1 U1012 ( .A1(n1288), .A2(n1120), .ZN(n1287) );
XOR2_X1 U1013 ( .A(n1145), .B(n1289), .Z(n1288) );
XNOR2_X1 U1014 ( .A(n1290), .B(n1291), .ZN(n1289) );
NOR2_X1 U1015 ( .A1(KEYINPUT60), .A2(n1143), .ZN(n1291) );
XNOR2_X1 U1016 ( .A(G140), .B(KEYINPUT21), .ZN(n1143) );
NAND2_X1 U1017 ( .A1(KEYINPUT32), .A2(n1292), .ZN(n1290) );
XNOR2_X1 U1018 ( .A(n1249), .B(n1152), .ZN(n1292) );
XOR2_X1 U1019 ( .A(n1293), .B(n1294), .Z(n1152) );
XNOR2_X1 U1020 ( .A(n1006), .B(G104), .ZN(n1294) );
INV_X1 U1021 ( .A(G107), .ZN(n1006) );
XNOR2_X1 U1022 ( .A(G101), .B(n1083), .ZN(n1293) );
XNOR2_X1 U1023 ( .A(n1295), .B(n1296), .ZN(n1083) );
NOR2_X1 U1024 ( .A1(KEYINPUT9), .A2(n1238), .ZN(n1296) );
XNOR2_X1 U1025 ( .A(G143), .B(G146), .ZN(n1238) );
XOR2_X1 U1026 ( .A(n1297), .B(n1194), .Z(n1249) );
INV_X1 U1027 ( .A(G131), .ZN(n1194) );
NAND2_X1 U1028 ( .A1(KEYINPUT63), .A2(n1082), .ZN(n1297) );
XNOR2_X1 U1029 ( .A(G134), .B(n1298), .ZN(n1082) );
XNOR2_X1 U1030 ( .A(n1299), .B(n1300), .ZN(n1145) );
NOR2_X1 U1031 ( .A1(n1070), .A2(G953), .ZN(n1300) );
INV_X1 U1032 ( .A(G227), .ZN(n1070) );
INV_X1 U1033 ( .A(G110), .ZN(n1299) );
INV_X1 U1034 ( .A(n1031), .ZN(n1028) );
NAND2_X1 U1035 ( .A1(G221), .A2(n1301), .ZN(n1031) );
INV_X1 U1036 ( .A(n1190), .ZN(n1197) );
XNOR2_X1 U1037 ( .A(n1050), .B(KEYINPUT53), .ZN(n1190) );
XNOR2_X1 U1038 ( .A(n1302), .B(n1113), .ZN(n1050) );
NAND2_X1 U1039 ( .A1(G217), .A2(n1301), .ZN(n1113) );
NAND2_X1 U1040 ( .A1(G234), .A2(n1284), .ZN(n1301) );
XNOR2_X1 U1041 ( .A(n1120), .B(KEYINPUT35), .ZN(n1284) );
INV_X1 U1042 ( .A(G902), .ZN(n1120) );
OR2_X1 U1043 ( .A1(n1115), .A2(G902), .ZN(n1302) );
XOR2_X1 U1044 ( .A(n1303), .B(n1304), .Z(n1115) );
XNOR2_X1 U1045 ( .A(n1305), .B(n1255), .ZN(n1304) );
XOR2_X1 U1046 ( .A(G119), .B(KEYINPUT41), .Z(n1255) );
NAND2_X1 U1047 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U1048 ( .A1(G146), .A2(n1081), .ZN(n1307) );
XOR2_X1 U1049 ( .A(n1308), .B(KEYINPUT10), .Z(n1306) );
OR2_X1 U1050 ( .A1(n1081), .A2(G146), .ZN(n1308) );
XOR2_X1 U1051 ( .A(G140), .B(G125), .Z(n1081) );
XOR2_X1 U1052 ( .A(n1309), .B(n1310), .Z(n1303) );
XNOR2_X1 U1053 ( .A(n1295), .B(G110), .ZN(n1310) );
INV_X1 U1054 ( .A(G128), .ZN(n1295) );
NAND2_X1 U1055 ( .A1(n1311), .A2(n1312), .ZN(n1309) );
NAND3_X1 U1056 ( .A1(n1313), .A2(n1217), .A3(G221), .ZN(n1312) );
INV_X1 U1057 ( .A(n1298), .ZN(n1313) );
XOR2_X1 U1058 ( .A(n1314), .B(KEYINPUT24), .Z(n1311) );
NAND2_X1 U1059 ( .A1(n1298), .A2(n1315), .ZN(n1314) );
NAND2_X1 U1060 ( .A1(G221), .A2(n1217), .ZN(n1315) );
AND2_X1 U1061 ( .A1(G234), .A2(n1069), .ZN(n1217) );
INV_X1 U1062 ( .A(G953), .ZN(n1069) );
XOR2_X1 U1063 ( .A(G137), .B(KEYINPUT33), .Z(n1298) );
endmodule


