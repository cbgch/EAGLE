//Key = 1101001010000011100001011101001011000101111101111110011000000101
module c3540 ( G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107,
G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270,
G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
G1698, G2897, G353, G355, G361, G358, G351, G372, G369, G399, G364,
G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405,
G402, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63 );

input G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330,
G343, G1698, G2897, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3,
KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9,
KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39,
KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63;

output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;

wire   n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347;

NOR3_X2 U1727 ( .A1(n3011), .A2(n3005), .A3(n3003), .ZN(n2615) );
NOR3_X2 U1728 ( .A1(n3003), .A2(n3011), .A3(n3004), .ZN(n2601) );
NOR3_X2 U1729 ( .A1(n2787), .A2(G1), .A3(n3031), .ZN(n3079) );
NOR3_X2 U1730 ( .A1(n3005), .A2(G200), .A3(n3003), .ZN(n2602) );
NAND3_X1 U1731 ( .A1(n2518), .A2(n2519), .A3(G213), .ZN(G409) );
NAND2_X1 U1732 ( .A1(n2520), .A2(n2521), .ZN(n2519) );
NAND3_X1 U1733 ( .A1(n2522), .A2(n2523), .A3(n2524), .ZN(n2518) );
NAND2_X1 U1734 ( .A1(n2521), .A2(n2525), .ZN(G407) );
XOR2_X1 U1735 ( .A(KEYINPUT13), .B(n2520), .Z(n2525) );
NOR4_X1 U1736 ( .A1(G384), .A2(G375), .A3(G378), .A4(G381), .ZN(n2520) );
NOR4_X1 U1737 ( .A1(n2526), .A2(n2527), .A3(G396), .A4(G393), .ZN(n2521) );
INV_X1 U1738 ( .A(n2528), .ZN(n2527) );
XNOR2_X1 U1739 ( .A(n2529), .B(n2530), .ZN(G405) );
INV_X1 U1740 ( .A(n2531), .ZN(n2530) );
NAND3_X1 U1741 ( .A1(n2532), .A2(n2533), .A3(n2534), .ZN(n2529) );
NAND4_X1 U1742 ( .A1(G2897), .A2(n2535), .A3(n2536), .A4(n2537), .ZN(n2534) );
OR2_X1 U1743 ( .A1(n2538), .A2(n2539), .ZN(n2535) );
NAND3_X1 U1744 ( .A1(n2540), .A2(n2538), .A3(n2541), .ZN(n2533) );
NAND2_X1 U1745 ( .A1(n2542), .A2(n2536), .ZN(n2538) );
XNOR2_X1 U1746 ( .A(n2522), .B(n2543), .ZN(n2542) );
NOR2_X1 U1747 ( .A1(n2523), .A2(KEYINPUT28), .ZN(n2543) );
NAND2_X1 U1748 ( .A1(n2544), .A2(n2545), .ZN(n2532) );
NAND2_X1 U1749 ( .A1(n2546), .A2(n2547), .ZN(n2545) );
OR2_X1 U1750 ( .A1(n2537), .A2(n2540), .ZN(n2547) );
NAND2_X1 U1751 ( .A1(G2897), .A2(n2524), .ZN(n2540) );
INV_X1 U1752 ( .A(KEYINPUT46), .ZN(n2537) );
NAND2_X1 U1753 ( .A1(n2539), .A2(n2536), .ZN(n2546) );
INV_X1 U1754 ( .A(n2524), .ZN(n2536) );
NOR2_X1 U1755 ( .A1(n2548), .A2(G343), .ZN(n2524) );
XOR2_X1 U1756 ( .A(G213), .B(KEYINPUT33), .Z(n2548) );
XNOR2_X1 U1757 ( .A(n2522), .B(G378), .ZN(n2539) );
XNOR2_X1 U1758 ( .A(n2549), .B(n2544), .ZN(G402) );
INV_X1 U1759 ( .A(n2541), .ZN(n2544) );
XOR2_X1 U1760 ( .A(G381), .B(G384), .Z(n2541) );
XNOR2_X1 U1761 ( .A(n2531), .B(n2550), .ZN(n2549) );
NOR2_X1 U1762 ( .A1(n2551), .A2(n2552), .ZN(n2550) );
XOR2_X1 U1763 ( .A(KEYINPUT2), .B(n2553), .Z(n2552) );
NOR2_X1 U1764 ( .A1(n2523), .A2(G375), .ZN(n2553) );
INV_X1 U1765 ( .A(G378), .ZN(n2523) );
NOR2_X1 U1766 ( .A1(G378), .A2(n2522), .ZN(n2551) );
INV_X1 U1767 ( .A(G375), .ZN(n2522) );
XNOR2_X1 U1768 ( .A(n2554), .B(n2555), .ZN(n2531) );
XNOR2_X1 U1769 ( .A(n2556), .B(G393), .ZN(n2555) );
XNOR2_X1 U1770 ( .A(G396), .B(n2557), .ZN(n2554) );
NAND2_X1 U1771 ( .A1(n2558), .A2(n2559), .ZN(G396) );
NAND3_X1 U1772 ( .A1(n2560), .A2(n2561), .A3(n2562), .ZN(n2559) );
NAND2_X1 U1773 ( .A1(n2563), .A2(n2564), .ZN(n2560) );
XNOR2_X1 U1774 ( .A(n2565), .B(n2566), .ZN(n2563) );
NAND2_X1 U1775 ( .A1(n2567), .A2(n2568), .ZN(n2558) );
NOR4_X1 U1776 ( .A1(n2569), .A2(n2570), .A3(n2571), .A4(n2572), .ZN(n2567) );
NOR2_X1 U1777 ( .A1(n2573), .A2(n2574), .ZN(n2572) );
NOR3_X1 U1778 ( .A1(n2575), .A2(n2576), .A3(n2577), .ZN(n2573) );
NOR2_X1 U1779 ( .A1(n2578), .A2(n2579), .ZN(n2577) );
NOR2_X1 U1780 ( .A1(n2580), .A2(n2581), .ZN(n2579) );
AND2_X1 U1781 ( .A1(n2582), .A2(G45), .ZN(n2581) );
NOR2_X1 U1782 ( .A1(G45), .A2(n2583), .ZN(n2580) );
NOR3_X1 U1783 ( .A1(n2584), .A2(n2585), .A3(n2586), .ZN(n2576) );
XNOR2_X1 U1784 ( .A(KEYINPUT52), .B(n2587), .ZN(n2586) );
AND2_X1 U1785 ( .A1(G355), .A2(n2585), .ZN(n2575) );
NOR3_X1 U1786 ( .A1(n2588), .A2(KEYINPUT20), .A3(n2565), .ZN(n2571) );
INV_X1 U1787 ( .A(n2589), .ZN(n2565) );
NOR4_X1 U1788 ( .A1(n2590), .A2(n2591), .A3(n2592), .A4(n2593), .ZN(n2570) );
NOR2_X1 U1789 ( .A1(n2594), .A2(n2595), .ZN(n2593) );
NOR2_X1 U1790 ( .A1(n2596), .A2(n2597), .ZN(n2592) );
NAND3_X1 U1791 ( .A1(n2598), .A2(n2599), .A3(n2600), .ZN(n2591) );
NAND2_X1 U1792 ( .A1(G68), .A2(n2601), .ZN(n2600) );
NAND2_X1 U1793 ( .A1(G58), .A2(n2602), .ZN(n2598) );
NAND4_X1 U1794 ( .A1(n2603), .A2(n2604), .A3(n2605), .A4(n2606), .ZN(n2590) );
NAND2_X1 U1795 ( .A1(n2607), .A2(G107), .ZN(n2606) );
NAND2_X1 U1796 ( .A1(G159), .A2(n2608), .ZN(n2605) );
NAND2_X1 U1797 ( .A1(G87), .A2(n2609), .ZN(n2604) );
NOR4_X1 U1798 ( .A1(n2610), .A2(n2611), .A3(n2612), .A4(n2613), .ZN(n2569) );
NOR2_X1 U1799 ( .A1(n2595), .A2(n2614), .ZN(n2613) );
AND2_X1 U1800 ( .A1(n2615), .A2(G326), .ZN(n2612) );
NAND3_X1 U1801 ( .A1(n2616), .A2(n2617), .A3(n2618), .ZN(n2611) );
NAND2_X1 U1802 ( .A1(G317), .A2(n2601), .ZN(n2618) );
NAND2_X1 U1803 ( .A1(G303), .A2(n2619), .ZN(n2617) );
NAND2_X1 U1804 ( .A1(G322), .A2(n2602), .ZN(n2616) );
NAND4_X1 U1805 ( .A1(n2620), .A2(n2621), .A3(n2622), .A4(n2623), .ZN(n2610) );
NAND2_X1 U1806 ( .A1(G283), .A2(n2607), .ZN(n2623) );
NAND2_X1 U1807 ( .A1(G329), .A2(n2608), .ZN(n2622) );
NAND2_X1 U1808 ( .A1(G294), .A2(n2624), .ZN(n2621) );
NAND3_X1 U1809 ( .A1(n2625), .A2(n2626), .A3(n2627), .ZN(G393) );
NAND2_X1 U1810 ( .A1(n2628), .A2(n2629), .ZN(n2627) );
XOR2_X1 U1811 ( .A(n2630), .B(n2631), .Z(n2628) );
XOR2_X1 U1812 ( .A(KEYINPUT11), .B(n2632), .Z(n2631) );
XNOR2_X1 U1813 ( .A(n2561), .B(n2633), .ZN(n2630) );
NAND4_X1 U1814 ( .A1(n2568), .A2(n2634), .A3(n2635), .A4(n2636), .ZN(n2626) );
NAND2_X1 U1815 ( .A1(n2637), .A2(n2638), .ZN(n2636) );
NAND3_X1 U1816 ( .A1(n2639), .A2(n2640), .A3(n2641), .ZN(n2638) );
NAND2_X1 U1817 ( .A1(n2585), .A2(n2642), .ZN(n2641) );
NAND3_X1 U1818 ( .A1(n2643), .A2(n2644), .A3(n2578), .ZN(n2640) );
NAND2_X1 U1819 ( .A1(n2645), .A2(n2584), .ZN(n2639) );
NAND2_X1 U1820 ( .A1(n2646), .A2(n2647), .ZN(n2645) );
NAND2_X1 U1821 ( .A1(n2648), .A2(n2649), .ZN(n2647) );
NAND4_X1 U1822 ( .A1(n2650), .A2(G58), .A3(n2651), .A4(n2597), .ZN(n2648) );
NAND2_X1 U1823 ( .A1(n2652), .A2(G77), .ZN(n2651) );
NAND2_X1 U1824 ( .A1(n2653), .A2(G45), .ZN(n2646) );
XOR2_X1 U1825 ( .A(n2654), .B(n2655), .Z(n2653) );
XOR2_X1 U1826 ( .A(KEYINPUT25), .B(n2656), .Z(n2655) );
NOR2_X1 U1827 ( .A1(n2657), .A2(n2658), .ZN(n2635) );
NOR4_X1 U1828 ( .A1(n2659), .A2(n2660), .A3(n2661), .A4(n2662), .ZN(n2658) );
NOR2_X1 U1829 ( .A1(n2595), .A2(n2663), .ZN(n2662) );
NOR2_X1 U1830 ( .A1(n2596), .A2(n2664), .ZN(n2661) );
NAND3_X1 U1831 ( .A1(n2665), .A2(n2666), .A3(n2667), .ZN(n2660) );
NAND2_X1 U1832 ( .A1(G58), .A2(n2601), .ZN(n2667) );
NAND2_X1 U1833 ( .A1(G50), .A2(n2602), .ZN(n2665) );
NAND4_X1 U1834 ( .A1(n2603), .A2(n2668), .A3(n2669), .A4(n2670), .ZN(n2659) );
NAND2_X1 U1835 ( .A1(G150), .A2(n2608), .ZN(n2669) );
NAND2_X1 U1836 ( .A1(G77), .A2(n2609), .ZN(n2668) );
NOR4_X1 U1837 ( .A1(n2671), .A2(n2672), .A3(n2673), .A4(n2674), .ZN(n2657) );
NOR2_X1 U1838 ( .A1(n2595), .A2(n2675), .ZN(n2674) );
NOR2_X1 U1839 ( .A1(n2596), .A2(n2676), .ZN(n2673) );
NAND3_X1 U1840 ( .A1(n2677), .A2(n2678), .A3(n2679), .ZN(n2672) );
NAND2_X1 U1841 ( .A1(G311), .A2(n2601), .ZN(n2679) );
NAND2_X1 U1842 ( .A1(n2680), .A2(n2619), .ZN(n2678) );
XNOR2_X1 U1843 ( .A(G294), .B(KEYINPUT47), .ZN(n2680) );
NAND2_X1 U1844 ( .A1(G317), .A2(n2602), .ZN(n2677) );
NAND4_X1 U1845 ( .A1(n2620), .A2(n2681), .A3(n2682), .A4(n2683), .ZN(n2671) );
NAND2_X1 U1846 ( .A1(n2607), .A2(G116), .ZN(n2683) );
NAND2_X1 U1847 ( .A1(G326), .A2(n2608), .ZN(n2682) );
NAND2_X1 U1848 ( .A1(G283), .A2(n2624), .ZN(n2681) );
NAND2_X1 U1849 ( .A1(n2684), .A2(n2685), .ZN(n2634) );
NAND2_X1 U1850 ( .A1(n2686), .A2(n2687), .ZN(n2625) );
XNOR2_X1 U1851 ( .A(KEYINPUT43), .B(n2688), .ZN(n2686) );
NOR2_X1 U1852 ( .A1(n2689), .A2(n2557), .ZN(G390) );
NAND2_X1 U1853 ( .A1(n2690), .A2(n2691), .ZN(n2557) );
OR2_X1 U1854 ( .A1(n2526), .A2(KEYINPUT22), .ZN(n2691) );
NAND3_X1 U1855 ( .A1(n2692), .A2(n2688), .A3(KEYINPUT22), .ZN(n2690) );
INV_X1 U1856 ( .A(n2526), .ZN(n2689) );
NAND3_X1 U1857 ( .A1(n2693), .A2(n2694), .A3(n2695), .ZN(n2526) );
NAND2_X1 U1858 ( .A1(n2692), .A2(n2688), .ZN(n2695) );
NAND4_X1 U1859 ( .A1(n2568), .A2(n2696), .A3(n2697), .A4(n2698), .ZN(n2694) );
NAND3_X1 U1860 ( .A1(n2699), .A2(n2700), .A3(n2701), .ZN(n2698) );
XNOR2_X1 U1861 ( .A(KEYINPUT26), .B(n2702), .ZN(n2701) );
NAND2_X1 U1862 ( .A1(G33), .A2(n2703), .ZN(n2700) );
NAND2_X1 U1863 ( .A1(n2704), .A2(n2705), .ZN(n2703) );
NOR4_X1 U1864 ( .A1(n2706), .A2(n2707), .A3(n2708), .A4(n2709), .ZN(n2705) );
NOR2_X1 U1865 ( .A1(n2710), .A2(n2711), .ZN(n2709) );
NOR2_X1 U1866 ( .A1(n2712), .A2(n2675), .ZN(n2708) );
NOR2_X1 U1867 ( .A1(n2713), .A2(n2614), .ZN(n2707) );
INV_X1 U1868 ( .A(G311), .ZN(n2614) );
NOR2_X1 U1869 ( .A1(n2714), .A2(n2715), .ZN(n2706) );
XNOR2_X1 U1870 ( .A(G107), .B(KEYINPUT19), .ZN(n2714) );
NOR4_X1 U1871 ( .A1(n2716), .A2(n2717), .A3(n2718), .A4(n2719), .ZN(n2704) );
NOR2_X1 U1872 ( .A1(n2720), .A2(n2587), .ZN(n2719) );
NOR2_X1 U1873 ( .A1(n2721), .A2(n2676), .ZN(n2718) );
INV_X1 U1874 ( .A(G322), .ZN(n2676) );
AND2_X1 U1875 ( .A1(n2722), .A2(G294), .ZN(n2717) );
AND2_X1 U1876 ( .A1(n2615), .A2(G317), .ZN(n2716) );
NAND2_X1 U1877 ( .A1(n2723), .A2(n2724), .ZN(n2699) );
NAND4_X1 U1878 ( .A1(n2725), .A2(n2726), .A3(n2727), .A4(n2728), .ZN(n2723) );
NOR4_X1 U1879 ( .A1(n2729), .A2(n2730), .A3(n2731), .A4(n2732), .ZN(n2728) );
NOR2_X1 U1880 ( .A1(n2721), .A2(n2733), .ZN(n2732) );
NOR2_X1 U1881 ( .A1(n2734), .A2(n2715), .ZN(n2731) );
NOR2_X1 U1882 ( .A1(n2595), .A2(n2735), .ZN(n2730) );
NOR2_X1 U1883 ( .A1(n2596), .A2(n2736), .ZN(n2729) );
NOR2_X1 U1884 ( .A1(n2737), .A2(n2738), .ZN(n2727) );
NOR2_X1 U1885 ( .A1(n2739), .A2(n2663), .ZN(n2738) );
NAND2_X1 U1886 ( .A1(G159), .A2(n2602), .ZN(n2726) );
NAND2_X1 U1887 ( .A1(G50), .A2(n2601), .ZN(n2725) );
NAND2_X1 U1888 ( .A1(n2637), .A2(n2740), .ZN(n2697) );
NAND3_X1 U1889 ( .A1(n2741), .A2(n2742), .A3(n2643), .ZN(n2740) );
INV_X1 U1890 ( .A(n2585), .ZN(n2643) );
NAND2_X1 U1891 ( .A1(n2578), .A2(n2743), .ZN(n2742) );
NAND2_X1 U1892 ( .A1(n2744), .A2(n2584), .ZN(n2741) );
INV_X1 U1893 ( .A(n2574), .ZN(n2637) );
NAND2_X1 U1894 ( .A1(n2745), .A2(n2684), .ZN(n2696) );
NAND2_X1 U1895 ( .A1(n2629), .A2(n2746), .ZN(n2693) );
XNOR2_X1 U1896 ( .A(n2747), .B(n2692), .ZN(n2746) );
NAND2_X1 U1897 ( .A1(n2632), .A2(n2687), .ZN(n2747) );
NOR2_X1 U1898 ( .A1(n2556), .A2(n2528), .ZN(G387) );
NAND2_X1 U1899 ( .A1(n2748), .A2(n2749), .ZN(n2528) );
OR2_X1 U1900 ( .A1(n2750), .A2(KEYINPUT3), .ZN(n2749) );
NAND2_X1 U1901 ( .A1(n2556), .A2(KEYINPUT3), .ZN(n2748) );
AND3_X1 U1902 ( .A1(n2751), .A2(n2750), .A3(n2752), .ZN(n2556) );
NAND2_X1 U1903 ( .A1(n2753), .A2(n2688), .ZN(n2752) );
NAND3_X1 U1904 ( .A1(n2568), .A2(n2754), .A3(n2755), .ZN(n2750) );
NOR3_X1 U1905 ( .A1(n2756), .A2(n2757), .A3(n2758), .ZN(n2755) );
NOR4_X1 U1906 ( .A1(n2759), .A2(n2760), .A3(n2761), .A4(n2762), .ZN(n2758) );
NOR2_X1 U1907 ( .A1(n2587), .A2(n2710), .ZN(n2762) );
NOR2_X1 U1908 ( .A1(n2595), .A2(n2711), .ZN(n2761) );
NAND3_X1 U1909 ( .A1(n2763), .A2(n2764), .A3(n2765), .ZN(n2760) );
NAND2_X1 U1910 ( .A1(G294), .A2(n2601), .ZN(n2765) );
NAND2_X1 U1911 ( .A1(G311), .A2(n2615), .ZN(n2764) );
NAND2_X1 U1912 ( .A1(G303), .A2(n2602), .ZN(n2763) );
NAND4_X1 U1913 ( .A1(n2620), .A2(n2766), .A3(n2767), .A4(n2670), .ZN(n2759) );
NAND2_X1 U1914 ( .A1(n2607), .A2(G97), .ZN(n2670) );
NAND2_X1 U1915 ( .A1(G317), .A2(n2608), .ZN(n2767) );
NAND2_X1 U1916 ( .A1(G107), .A2(n2624), .ZN(n2766) );
NOR2_X1 U1917 ( .A1(n2724), .A2(n2702), .ZN(n2620) );
NOR4_X1 U1918 ( .A1(n2768), .A2(n2769), .A3(n2770), .A4(n2771), .ZN(n2757) );
NOR2_X1 U1919 ( .A1(n2596), .A2(n2733), .ZN(n2771) );
NOR2_X1 U1920 ( .A1(n2712), .A2(n2664), .ZN(n2770) );
NAND3_X1 U1921 ( .A1(n2772), .A2(n2773), .A3(n2774), .ZN(n2769) );
NAND2_X1 U1922 ( .A1(G150), .A2(n2602), .ZN(n2774) );
NAND2_X1 U1923 ( .A1(n2775), .A2(G50), .ZN(n2773) );
XNOR2_X1 U1924 ( .A(n2722), .B(KEYINPUT32), .ZN(n2775) );
NAND4_X1 U1925 ( .A1(n2603), .A2(n2776), .A3(n2777), .A4(n2778), .ZN(n2768) );
NAND2_X1 U1926 ( .A1(G58), .A2(n2609), .ZN(n2778) );
NAND2_X1 U1927 ( .A1(G137), .A2(n2608), .ZN(n2776) );
NOR2_X1 U1928 ( .A1(n2702), .A2(G33), .ZN(n2603) );
NOR2_X1 U1929 ( .A1(n2779), .A2(n2574), .ZN(n2756) );
NAND2_X1 U1930 ( .A1(n2702), .A2(n2588), .ZN(n2574) );
NOR3_X1 U1931 ( .A1(n2780), .A2(n2585), .A3(n2781), .ZN(n2779) );
NOR2_X1 U1932 ( .A1(n2782), .A2(n2578), .ZN(n2781) );
NOR2_X1 U1933 ( .A1(n2783), .A2(G33), .ZN(n2585) );
XOR2_X1 U1934 ( .A(n2784), .B(KEYINPUT39), .Z(n2780) );
NAND2_X1 U1935 ( .A1(n2734), .A2(n2578), .ZN(n2784) );
INV_X1 U1936 ( .A(n2584), .ZN(n2578) );
NOR2_X1 U1937 ( .A1(n2724), .A2(n2783), .ZN(n2584) );
NAND2_X1 U1938 ( .A1(n2785), .A2(n2684), .ZN(n2754) );
INV_X1 U1939 ( .A(n2588), .ZN(n2684) );
NAND2_X1 U1940 ( .A1(n2786), .A2(n2787), .ZN(n2588) );
NAND3_X1 U1941 ( .A1(n2629), .A2(n2788), .A3(n2753), .ZN(n2751) );
XNOR2_X1 U1942 ( .A(n2789), .B(n2785), .ZN(n2753) );
XOR2_X1 U1943 ( .A(n2790), .B(n2791), .Z(n2785) );
NOR2_X1 U1944 ( .A1(n2792), .A2(n2793), .ZN(n2791) );
XOR2_X1 U1945 ( .A(n2794), .B(n2795), .Z(n2789) );
NOR3_X1 U1946 ( .A1(n2561), .A2(n2745), .A3(n2796), .ZN(n2795) );
NAND2_X1 U1947 ( .A1(n2797), .A2(n2798), .ZN(n2794) );
NAND2_X1 U1948 ( .A1(n2799), .A2(n2800), .ZN(n2798) );
OR2_X1 U1949 ( .A1(n2801), .A2(n2802), .ZN(n2797) );
NAND2_X1 U1950 ( .A1(n2632), .A2(n2803), .ZN(n2788) );
NAND2_X1 U1951 ( .A1(n2692), .A2(n2687), .ZN(n2803) );
XNOR2_X1 U1952 ( .A(n2804), .B(n2805), .ZN(n2687) );
NAND2_X1 U1953 ( .A1(KEYINPUT24), .A2(n2633), .ZN(n2804) );
XNOR2_X1 U1954 ( .A(n2806), .B(n2807), .ZN(n2633) );
NAND2_X1 U1955 ( .A1(n2808), .A2(n2793), .ZN(n2806) );
XOR2_X1 U1956 ( .A(n2809), .B(n2745), .Z(n2692) );
INV_X1 U1957 ( .A(n2800), .ZN(n2745) );
XOR2_X1 U1958 ( .A(n2810), .B(n2811), .Z(n2800) );
NOR2_X1 U1959 ( .A1(n2812), .A2(n2793), .ZN(n2811) );
NAND2_X1 U1960 ( .A1(G399), .A2(n2813), .ZN(n2809) );
NAND3_X1 U1961 ( .A1(n2807), .A2(n2805), .A3(n2799), .ZN(n2813) );
INV_X1 U1962 ( .A(n2814), .ZN(n2799) );
NAND2_X1 U1963 ( .A1(n2814), .A2(n2815), .ZN(G399) );
NAND2_X1 U1964 ( .A1(n2805), .A2(n2807), .ZN(n2815) );
INV_X1 U1965 ( .A(n2561), .ZN(n2805) );
NAND2_X1 U1966 ( .A1(G330), .A2(n2816), .ZN(n2561) );
XNOR2_X1 U1967 ( .A(n2589), .B(n2566), .ZN(n2816) );
NOR2_X1 U1968 ( .A1(n2793), .A2(n2817), .ZN(n2566) );
NAND2_X1 U1969 ( .A1(n2793), .A2(n2818), .ZN(n2814) );
NAND2_X1 U1970 ( .A1(n2819), .A2(n2820), .ZN(n2818) );
NAND2_X1 U1971 ( .A1(n2807), .A2(n2808), .ZN(n2819) );
INV_X1 U1972 ( .A(n2821), .ZN(n2808) );
INV_X1 U1973 ( .A(n2796), .ZN(n2807) );
XOR2_X1 U1974 ( .A(n2822), .B(n2685), .Z(n2796) );
NAND2_X1 U1975 ( .A1(KEYINPUT30), .A2(n2823), .ZN(n2822) );
NAND2_X1 U1976 ( .A1(n2802), .A2(n2824), .ZN(n2823) );
NAND2_X1 U1977 ( .A1(n2825), .A2(n2826), .ZN(G384) );
NAND4_X1 U1978 ( .A1(n2827), .A2(n2828), .A3(n2829), .A4(n2562), .ZN(n2826) );
NAND2_X1 U1979 ( .A1(n2830), .A2(n2632), .ZN(n2828) );
NAND2_X1 U1980 ( .A1(n2831), .A2(n2832), .ZN(n2827) );
NAND4_X1 U1981 ( .A1(n2833), .A2(n2834), .A3(n2835), .A4(n2568), .ZN(n2825) );
NOR2_X1 U1982 ( .A1(n2836), .A2(n2837), .ZN(n2835) );
NOR4_X1 U1983 ( .A1(n2838), .A2(n2839), .A3(n2840), .A4(n2841), .ZN(n2837) );
NOR2_X1 U1984 ( .A1(n2712), .A2(n2736), .ZN(n2841) );
NOR2_X1 U1985 ( .A1(n2720), .A2(n2735), .ZN(n2840) );
NAND3_X1 U1986 ( .A1(n2842), .A2(n2843), .A3(n2844), .ZN(n2839) );
NAND2_X1 U1987 ( .A1(G132), .A2(n2608), .ZN(n2844) );
NAND2_X1 U1988 ( .A1(G50), .A2(n2609), .ZN(n2843) );
NAND2_X1 U1989 ( .A1(G137), .A2(n2615), .ZN(n2842) );
NAND3_X1 U1990 ( .A1(n2845), .A2(n2846), .A3(n2847), .ZN(n2838) );
NOR3_X1 U1991 ( .A1(n2848), .A2(n2849), .A3(n2850), .ZN(n2847) );
NOR2_X1 U1992 ( .A1(n2715), .A2(n2663), .ZN(n2850) );
NOR2_X1 U1993 ( .A1(n2595), .A2(n2664), .ZN(n2849) );
NOR2_X1 U1994 ( .A1(n2713), .A2(n2733), .ZN(n2848) );
XNOR2_X1 U1995 ( .A(KEYINPUT0), .B(n2724), .ZN(n2846) );
NOR4_X1 U1996 ( .A1(n2851), .A2(n2852), .A3(n2853), .A4(n2854), .ZN(n2836) );
NOR2_X1 U1997 ( .A1(n2587), .A2(n2595), .ZN(n2854) );
NOR2_X1 U1998 ( .A1(n2596), .A2(n2675), .ZN(n2853) );
INV_X1 U1999 ( .A(G303), .ZN(n2675) );
NAND3_X1 U2000 ( .A1(n2855), .A2(n2599), .A3(n2856), .ZN(n2852) );
NAND2_X1 U2001 ( .A1(n2619), .A2(G107), .ZN(n2856) );
NAND2_X1 U2002 ( .A1(G97), .A2(n2624), .ZN(n2599) );
NAND2_X1 U2003 ( .A1(G294), .A2(n2602), .ZN(n2855) );
NAND4_X1 U2004 ( .A1(n2857), .A2(n2858), .A3(n2859), .A4(n2860), .ZN(n2851) );
NAND2_X1 U2005 ( .A1(n2607), .A2(G87), .ZN(n2860) );
NAND2_X1 U2006 ( .A1(G311), .A2(n2608), .ZN(n2859) );
NAND2_X1 U2007 ( .A1(G283), .A2(n2861), .ZN(n2858) );
XNOR2_X1 U2008 ( .A(KEYINPUT51), .B(n2712), .ZN(n2861) );
NAND2_X1 U2009 ( .A1(n2862), .A2(n2594), .ZN(n2834) );
NAND2_X1 U2010 ( .A1(n2786), .A2(n2863), .ZN(n2833) );
NAND3_X1 U2011 ( .A1(n2864), .A2(n2865), .A3(n2866), .ZN(G381) );
NAND2_X1 U2012 ( .A1(n2867), .A2(n2629), .ZN(n2866) );
XOR2_X1 U2013 ( .A(n2868), .B(n2869), .Z(n2867) );
XNOR2_X1 U2014 ( .A(n2870), .B(n2871), .ZN(n2869) );
XNOR2_X1 U2015 ( .A(KEYINPUT53), .B(KEYINPUT21), .ZN(n2868) );
NAND3_X1 U2016 ( .A1(n2568), .A2(n2872), .A3(n2873), .ZN(n2865) );
NOR3_X1 U2017 ( .A1(n2874), .A2(n2875), .A3(n2876), .ZN(n2873) );
NOR4_X1 U2018 ( .A1(n2877), .A2(n2878), .A3(n2879), .A4(n2880), .ZN(n2876) );
NOR2_X1 U2019 ( .A1(n2713), .A2(n2881), .ZN(n2880) );
INV_X1 U2020 ( .A(n2602), .ZN(n2713) );
NOR2_X1 U2021 ( .A1(n2739), .A2(n2664), .ZN(n2879) );
INV_X1 U2022 ( .A(n2609), .ZN(n2739) );
NAND3_X1 U2023 ( .A1(n2882), .A2(n2724), .A3(n2883), .ZN(n2878) );
NAND2_X1 U2024 ( .A1(G58), .A2(n2884), .ZN(n2883) );
XNOR2_X1 U2025 ( .A(KEYINPUT18), .B(n2715), .ZN(n2884) );
NAND2_X1 U2026 ( .A1(G143), .A2(n2601), .ZN(n2882) );
NAND4_X1 U2027 ( .A1(n2885), .A2(n2886), .A3(n2887), .A4(n2888), .ZN(n2877) );
NOR2_X1 U2028 ( .A1(n2889), .A2(n2890), .ZN(n2888) );
NOR2_X1 U2029 ( .A1(n2596), .A2(n2891), .ZN(n2889) );
NAND2_X1 U2030 ( .A1(G50), .A2(n2624), .ZN(n2887) );
NAND2_X1 U2031 ( .A1(G128), .A2(n2608), .ZN(n2886) );
NAND2_X1 U2032 ( .A1(G150), .A2(n2722), .ZN(n2885) );
NOR4_X1 U2033 ( .A1(n2892), .A2(n2893), .A3(n2894), .A4(n2895), .ZN(n2875) );
NOR2_X1 U2034 ( .A1(n2710), .A2(n2896), .ZN(n2895) );
XNOR2_X1 U2035 ( .A(KEYINPUT42), .B(n2743), .ZN(n2896) );
NOR2_X1 U2036 ( .A1(n2644), .A2(n2595), .ZN(n2894) );
NAND3_X1 U2037 ( .A1(n2897), .A2(n2666), .A3(n2898), .ZN(n2893) );
NAND2_X1 U2038 ( .A1(n2601), .A2(G116), .ZN(n2898) );
NAND2_X1 U2039 ( .A1(G87), .A2(n2624), .ZN(n2666) );
NAND2_X1 U2040 ( .A1(G283), .A2(n2602), .ZN(n2897) );
NAND4_X1 U2041 ( .A1(n2857), .A2(n2899), .A3(n2900), .A4(n2777), .ZN(n2892) );
NAND2_X1 U2042 ( .A1(n2607), .A2(G77), .ZN(n2777) );
NAND2_X1 U2043 ( .A1(G303), .A2(n2608), .ZN(n2900) );
NAND2_X1 U2044 ( .A1(n2615), .A2(G294), .ZN(n2899) );
NOR2_X1 U2045 ( .A1(G68), .A2(n2901), .ZN(n2874) );
NAND2_X1 U2046 ( .A1(n2902), .A2(n2786), .ZN(n2872) );
NAND2_X1 U2047 ( .A1(n2903), .A2(n2871), .ZN(n2864) );
XNOR2_X1 U2048 ( .A(n2904), .B(KEYINPUT62), .ZN(n2903) );
NAND3_X1 U2049 ( .A1(n2905), .A2(n2906), .A3(n2907), .ZN(G378) );
NAND2_X1 U2050 ( .A1(n2908), .A2(n2688), .ZN(n2907) );
NAND3_X1 U2051 ( .A1(n2568), .A2(n2909), .A3(n2910), .ZN(n2906) );
NOR3_X1 U2052 ( .A1(n2911), .A2(n2912), .A3(n2913), .ZN(n2910) );
NOR4_X1 U2053 ( .A1(n2914), .A2(n2915), .A3(n2916), .A4(n2917), .ZN(n2913) );
NOR2_X1 U2054 ( .A1(n2720), .A2(n2664), .ZN(n2917) );
NOR2_X1 U2055 ( .A1(n2721), .A2(n2918), .ZN(n2916) );
NAND3_X1 U2056 ( .A1(n2919), .A2(n2724), .A3(n2920), .ZN(n2915) );
NAND2_X1 U2057 ( .A1(G150), .A2(n2609), .ZN(n2920) );
NAND2_X1 U2058 ( .A1(G132), .A2(n2602), .ZN(n2919) );
NAND4_X1 U2059 ( .A1(n2921), .A2(n2922), .A3(n2923), .A4(n2924), .ZN(n2914) );
NOR2_X1 U2060 ( .A1(n2890), .A2(n2925), .ZN(n2924) );
XOR2_X1 U2061 ( .A(KEYINPUT9), .B(n2926), .Z(n2925) );
NOR2_X1 U2062 ( .A1(n2595), .A2(n2733), .ZN(n2926) );
INV_X1 U2063 ( .A(G143), .ZN(n2733) );
NAND2_X1 U2064 ( .A1(G137), .A2(n2601), .ZN(n2923) );
NAND2_X1 U2065 ( .A1(G128), .A2(n2615), .ZN(n2922) );
NAND2_X1 U2066 ( .A1(G50), .A2(n2607), .ZN(n2921) );
NOR4_X1 U2067 ( .A1(n2927), .A2(n2928), .A3(n2929), .A4(n2930), .ZN(n2912) );
NOR2_X1 U2068 ( .A1(n2710), .A2(n2734), .ZN(n2930) );
NOR2_X1 U2069 ( .A1(n2595), .A2(n2743), .ZN(n2929) );
NAND3_X1 U2070 ( .A1(n2931), .A2(n2932), .A3(n2933), .ZN(n2928) );
NAND2_X1 U2071 ( .A1(G107), .A2(n2601), .ZN(n2933) );
INV_X1 U2072 ( .A(n2737), .ZN(n2932) );
NOR2_X1 U2073 ( .A1(n2594), .A2(n2720), .ZN(n2737) );
NAND2_X1 U2074 ( .A1(G116), .A2(n2602), .ZN(n2931) );
NAND4_X1 U2075 ( .A1(n2857), .A2(n2934), .A3(n2935), .A4(n2936), .ZN(n2927) );
NAND2_X1 U2076 ( .A1(G68), .A2(n2607), .ZN(n2936) );
NAND2_X1 U2077 ( .A1(G294), .A2(n2608), .ZN(n2935) );
NAND2_X1 U2078 ( .A1(G283), .A2(n2615), .ZN(n2934) );
NOR2_X1 U2079 ( .A1(n2724), .A2(n2890), .ZN(n2857) );
NOR2_X1 U2080 ( .A1(G58), .A2(n2901), .ZN(n2911) );
NAND2_X1 U2081 ( .A1(n2786), .A2(n2937), .ZN(n2909) );
NAND2_X1 U2082 ( .A1(n2629), .A2(n2938), .ZN(n2905) );
XOR2_X1 U2083 ( .A(n2939), .B(n2908), .Z(n2938) );
AND2_X1 U2084 ( .A1(n2871), .A2(n2870), .ZN(n2939) );
NAND2_X1 U2085 ( .A1(n2940), .A2(n2941), .ZN(G375) );
NAND3_X1 U2086 ( .A1(n2942), .A2(n2943), .A3(n2562), .ZN(n2941) );
INV_X1 U2087 ( .A(n2568), .ZN(n2562) );
NAND3_X1 U2088 ( .A1(n2944), .A2(n2945), .A3(n2904), .ZN(n2943) );
INV_X1 U2089 ( .A(n2688), .ZN(n2904) );
OR2_X1 U2090 ( .A1(n2946), .A2(KEYINPUT8), .ZN(n2945) );
NAND2_X1 U2091 ( .A1(KEYINPUT8), .A2(n2947), .ZN(n2944) );
NAND2_X1 U2092 ( .A1(n2870), .A2(n2948), .ZN(n2947) );
NAND2_X1 U2093 ( .A1(n2871), .A2(n2908), .ZN(n2948) );
XOR2_X1 U2094 ( .A(n2949), .B(n2950), .Z(n2908) );
XOR2_X1 U2095 ( .A(n2951), .B(n2952), .Z(n2949) );
NOR2_X1 U2096 ( .A1(n2902), .A2(n2829), .ZN(n2952) );
INV_X1 U2097 ( .A(n2953), .ZN(n2902) );
XOR2_X1 U2098 ( .A(n2954), .B(n2955), .Z(n2871) );
XNOR2_X1 U2099 ( .A(n2956), .B(n2953), .ZN(n2955) );
NAND2_X1 U2100 ( .A1(n2957), .A2(n2958), .ZN(n2956) );
NAND2_X1 U2101 ( .A1(n2831), .A2(n2959), .ZN(n2958) );
XNOR2_X1 U2102 ( .A(KEYINPUT60), .B(n2830), .ZN(n2959) );
INV_X1 U2103 ( .A(n2832), .ZN(n2830) );
NAND2_X1 U2104 ( .A1(n2960), .A2(n2793), .ZN(n2957) );
XOR2_X1 U2105 ( .A(n2829), .B(KEYINPUT36), .Z(n2954) );
NAND2_X1 U2106 ( .A1(n2961), .A2(n2832), .ZN(n2829) );
INV_X1 U2107 ( .A(n2946), .ZN(n2870) );
NAND2_X1 U2108 ( .A1(n2962), .A2(n2963), .ZN(n2946) );
NAND2_X1 U2109 ( .A1(n2961), .A2(n2964), .ZN(n2963) );
XOR2_X1 U2110 ( .A(n2965), .B(n2966), .Z(n2942) );
XOR2_X1 U2111 ( .A(n2967), .B(n2968), .Z(n2966) );
NAND2_X1 U2112 ( .A1(n2969), .A2(n2970), .ZN(n2968) );
NAND2_X1 U2113 ( .A1(KEYINPUT63), .A2(n2971), .ZN(n2967) );
XOR2_X1 U2114 ( .A(n2972), .B(n2973), .Z(n2965) );
NOR2_X1 U2115 ( .A1(n2564), .A2(n2974), .ZN(n2973) );
INV_X1 U2116 ( .A(G330), .ZN(n2564) );
XNOR2_X1 U2117 ( .A(n2975), .B(KEYINPUT16), .ZN(n2972) );
NAND4_X1 U2118 ( .A1(n2976), .A2(n2977), .A3(n2978), .A4(n2568), .ZN(n2940) );
NOR2_X1 U2119 ( .A1(n2688), .A2(n2629), .ZN(n2568) );
NAND2_X1 U2120 ( .A1(G1), .A2(n2979), .ZN(n2688) );
NAND3_X1 U2121 ( .A1(G13), .A2(n2787), .A3(G45), .ZN(n2979) );
NAND2_X1 U2122 ( .A1(n2786), .A2(n2980), .ZN(n2978) );
NAND4_X1 U2123 ( .A1(n2845), .A2(n2981), .A3(n2982), .A4(n2983), .ZN(n2977) );
NAND2_X1 U2124 ( .A1(n2984), .A2(n2724), .ZN(n2983) );
XOR2_X1 U2125 ( .A(n2985), .B(KEYINPUT7), .Z(n2984) );
NAND4_X1 U2126 ( .A1(n2986), .A2(n2987), .A3(n2988), .A4(n2989), .ZN(n2985) );
NOR4_X1 U2127 ( .A1(n2990), .A2(n2991), .A3(n2992), .A4(n2993), .ZN(n2989) );
NOR2_X1 U2128 ( .A1(n2596), .A2(n2918), .ZN(n2993) );
INV_X1 U2129 ( .A(G125), .ZN(n2918) );
INV_X1 U2130 ( .A(n2615), .ZN(n2596) );
NOR2_X1 U2131 ( .A1(n2712), .A2(n2891), .ZN(n2992) );
INV_X1 U2132 ( .A(G132), .ZN(n2891) );
INV_X1 U2133 ( .A(n2601), .ZN(n2712) );
AND2_X1 U2134 ( .A1(n2602), .A2(G128), .ZN(n2991) );
NOR2_X1 U2135 ( .A1(n2595), .A2(n2881), .ZN(n2990) );
INV_X1 U2136 ( .A(G137), .ZN(n2881) );
NOR2_X1 U2137 ( .A1(n2994), .A2(n2995), .ZN(n2988) );
NOR2_X1 U2138 ( .A1(n2715), .A2(n2664), .ZN(n2995) );
INV_X1 U2139 ( .A(G159), .ZN(n2664) );
NOR2_X1 U2140 ( .A1(n2720), .A2(n2736), .ZN(n2994) );
INV_X1 U2141 ( .A(G150), .ZN(n2736) );
NAND2_X1 U2142 ( .A1(G124), .A2(n2608), .ZN(n2987) );
INV_X1 U2143 ( .A(n2721), .ZN(n2608) );
NAND2_X1 U2144 ( .A1(G143), .A2(n2609), .ZN(n2986) );
XOR2_X1 U2145 ( .A(n2619), .B(KEYINPUT5), .Z(n2609) );
NAND2_X1 U2146 ( .A1(n2996), .A2(G33), .ZN(n2982) );
XOR2_X1 U2147 ( .A(KEYINPUT48), .B(n2997), .Z(n2996) );
NOR4_X1 U2148 ( .A1(n2998), .A2(n2999), .A3(n3000), .A4(n3001), .ZN(n2997) );
XOR2_X1 U2149 ( .A(KEYINPUT55), .B(n3002), .Z(n3001) );
NOR2_X1 U2150 ( .A1(n2595), .A2(n2734), .ZN(n3002) );
INV_X1 U2151 ( .A(n2722), .ZN(n2595) );
NOR3_X1 U2152 ( .A1(n3003), .A2(G200), .A3(n3004), .ZN(n2722) );
NOR2_X1 U2153 ( .A1(n2721), .A2(n2711), .ZN(n3000) );
INV_X1 U2154 ( .A(G283), .ZN(n2711) );
NAND2_X1 U2155 ( .A1(n3005), .A2(n3006), .ZN(n2721) );
NAND2_X1 U2156 ( .A1(n3007), .A2(n3008), .ZN(n2999) );
NAND2_X1 U2157 ( .A1(n2619), .A2(G77), .ZN(n3008) );
INV_X1 U2158 ( .A(n2710), .ZN(n2619) );
NAND3_X1 U2159 ( .A1(G20), .A2(n3004), .A3(n3009), .ZN(n2710) );
NAND2_X1 U2160 ( .A1(G58), .A2(n2607), .ZN(n3007) );
INV_X1 U2161 ( .A(n2715), .ZN(n2607) );
NAND2_X1 U2162 ( .A1(n3009), .A2(n3005), .ZN(n2715) );
AND2_X1 U2163 ( .A1(n3010), .A2(n3003), .ZN(n3009) );
XNOR2_X1 U2164 ( .A(KEYINPUT35), .B(n3011), .ZN(n3010) );
NAND4_X1 U2165 ( .A1(n3012), .A2(n3013), .A3(n3014), .A4(n2772), .ZN(n2998) );
NAND2_X1 U2166 ( .A1(G68), .A2(n2624), .ZN(n2772) );
INV_X1 U2167 ( .A(n2720), .ZN(n2624) );
NAND2_X1 U2168 ( .A1(n3006), .A2(n3004), .ZN(n2720) );
AND2_X1 U2169 ( .A1(n3003), .A2(n3015), .ZN(n3006) );
NAND2_X1 U2170 ( .A1(G200), .A2(G20), .ZN(n3015) );
NAND2_X1 U2171 ( .A1(n2615), .A2(n3016), .ZN(n3014) );
XNOR2_X1 U2172 ( .A(KEYINPUT58), .B(n2587), .ZN(n3016) );
NAND2_X1 U2173 ( .A1(G107), .A2(n2602), .ZN(n3013) );
NAND2_X1 U2174 ( .A1(G97), .A2(n2601), .ZN(n3012) );
INV_X1 U2175 ( .A(n3005), .ZN(n3004) );
NOR2_X1 U2176 ( .A1(n2787), .A2(G190), .ZN(n3005) );
NAND2_X1 U2177 ( .A1(G179), .A2(G20), .ZN(n3003) );
NAND2_X1 U2178 ( .A1(n3017), .A2(n2597), .ZN(n2976) );
NAND2_X1 U2179 ( .A1(n2901), .A2(n3018), .ZN(n3017) );
NAND2_X1 U2180 ( .A1(G41), .A2(n2845), .ZN(n3018) );
INV_X1 U2181 ( .A(n2862), .ZN(n2901) );
NOR2_X1 U2182 ( .A1(n2845), .A2(n2786), .ZN(n2862) );
NOR2_X1 U2183 ( .A1(G13), .A2(G33), .ZN(n2786) );
INV_X1 U2184 ( .A(n2890), .ZN(n2845) );
XNOR2_X1 U2185 ( .A(n2702), .B(KEYINPUT14), .ZN(n2890) );
NAND2_X1 U2186 ( .A1(G13), .A2(n3019), .ZN(n2702) );
NAND2_X1 U2187 ( .A1(G20), .A2(n3020), .ZN(n3019) );
AND2_X1 U2188 ( .A1(n2964), .A2(n3021), .ZN(G372) );
NAND4_X1 U2189 ( .A1(n3022), .A2(n3023), .A3(n3024), .A4(n3025), .ZN(G369) );
NAND2_X1 U2190 ( .A1(n2964), .A2(n3026), .ZN(n3022) );
NAND3_X1 U2191 ( .A1(n3027), .A2(n3028), .A3(n3029), .ZN(G367) );
NAND3_X1 U2192 ( .A1(n3030), .A2(n3031), .A3(G1), .ZN(n3029) );
NAND2_X1 U2193 ( .A1(n3032), .A2(n3033), .ZN(n3030) );
NAND2_X1 U2194 ( .A1(n2652), .A2(n2597), .ZN(n3033) );
XNOR2_X1 U2195 ( .A(G68), .B(KEYINPUT23), .ZN(n2652) );
NAND3_X1 U2196 ( .A1(n3034), .A2(n3035), .A3(n3036), .ZN(n3028) );
NAND2_X1 U2197 ( .A1(G1), .A2(n3031), .ZN(n3035) );
XOR2_X1 U2198 ( .A(n2971), .B(n3037), .Z(n3034) );
XOR2_X1 U2199 ( .A(n3038), .B(n2962), .Z(n3037) );
AND4_X1 U2200 ( .A1(n3023), .A2(n3039), .A3(n3024), .A4(n3025), .ZN(n2962) );
NAND3_X1 U2201 ( .A1(n3040), .A2(n3041), .A3(n3042), .ZN(n3024) );
NAND2_X1 U2202 ( .A1(n3043), .A2(n2980), .ZN(n3041) );
NAND2_X1 U2203 ( .A1(n3044), .A2(n3045), .ZN(n3043) );
NAND2_X1 U2204 ( .A1(n3046), .A2(n3047), .ZN(n3040) );
NAND2_X1 U2205 ( .A1(n3044), .A2(n3048), .ZN(n3046) );
NAND2_X1 U2206 ( .A1(n2975), .A2(n3045), .ZN(n3048) );
INV_X1 U2207 ( .A(KEYINPUT1), .ZN(n3045) );
NOR2_X1 U2208 ( .A1(n3049), .A2(n3050), .ZN(n3044) );
NAND2_X1 U2209 ( .A1(n2964), .A2(n2831), .ZN(n3039) );
NAND2_X1 U2210 ( .A1(n3051), .A2(n2975), .ZN(n3023) );
INV_X1 U2211 ( .A(n2980), .ZN(n2975) );
NAND2_X1 U2212 ( .A1(n3052), .A2(n3053), .ZN(n3038) );
XOR2_X1 U2213 ( .A(n2974), .B(n3054), .Z(n3053) );
NAND2_X1 U2214 ( .A1(n2964), .A2(n3055), .ZN(n3054) );
NOR4_X1 U2215 ( .A1(n2863), .A2(n2937), .A3(n2980), .A4(n3049), .ZN(n2964) );
NAND2_X1 U2216 ( .A1(n3025), .A2(n3056), .ZN(n2980) );
NAND2_X1 U2217 ( .A1(n3057), .A2(n3058), .ZN(n3056) );
NAND3_X1 U2218 ( .A1(n3059), .A2(n3060), .A3(n3061), .ZN(n3058) );
NAND2_X1 U2219 ( .A1(n3062), .A2(n3011), .ZN(n3061) );
INV_X1 U2220 ( .A(G200), .ZN(n3011) );
NAND2_X1 U2221 ( .A1(n3063), .A2(G190), .ZN(n3062) );
NAND2_X1 U2222 ( .A1(KEYINPUT10), .A2(n3064), .ZN(n3060) );
OR3_X1 U2223 ( .A1(G190), .A2(KEYINPUT10), .A3(n3064), .ZN(n3059) );
INV_X1 U2224 ( .A(n2970), .ZN(n3057) );
NAND3_X1 U2225 ( .A1(n3065), .A2(n3066), .A3(n2970), .ZN(n3025) );
NAND3_X1 U2226 ( .A1(n3067), .A2(n3068), .A3(n3069), .ZN(n2970) );
NAND2_X1 U2227 ( .A1(n3070), .A2(n3071), .ZN(n3069) );
NAND3_X1 U2228 ( .A1(n3072), .A2(n3073), .A3(n3074), .ZN(n3071) );
NAND2_X1 U2229 ( .A1(G20), .A2(n3075), .ZN(n3074) );
NAND2_X1 U2230 ( .A1(n2597), .A2(n2663), .ZN(n3075) );
NAND2_X1 U2231 ( .A1(G58), .A2(n3076), .ZN(n3073) );
NAND2_X1 U2232 ( .A1(n3077), .A2(G150), .ZN(n3072) );
XNOR2_X1 U2233 ( .A(KEYINPUT31), .B(n3078), .ZN(n3070) );
NAND2_X1 U2234 ( .A1(n3079), .A2(n2597), .ZN(n3068) );
NAND2_X1 U2235 ( .A1(n3080), .A2(G50), .ZN(n3067) );
NAND2_X1 U2236 ( .A1(n3063), .A2(n3081), .ZN(n3066) );
INV_X1 U2237 ( .A(n3064), .ZN(n3063) );
NAND2_X1 U2238 ( .A1(n3064), .A2(n3020), .ZN(n3065) );
NAND3_X1 U2239 ( .A1(n3082), .A2(n3083), .A3(n3084), .ZN(n3064) );
NAND2_X1 U2240 ( .A1(n3085), .A2(G226), .ZN(n3084) );
NAND2_X1 U2241 ( .A1(n3086), .A2(n3087), .ZN(n3082) );
NAND3_X1 U2242 ( .A1(n3088), .A2(n3089), .A3(n3090), .ZN(n3087) );
NAND2_X1 U2243 ( .A1(G33), .A2(G77), .ZN(n3090) );
NAND2_X1 U2244 ( .A1(G223), .A2(n3091), .ZN(n3089) );
NAND2_X1 U2245 ( .A1(G222), .A2(n3092), .ZN(n3088) );
NAND4_X1 U2246 ( .A1(n2950), .A2(n2953), .A3(n2832), .A4(n3055), .ZN(n2974) );
XNOR2_X1 U2247 ( .A(G330), .B(KEYINPUT27), .ZN(n3052) );
NAND2_X1 U2248 ( .A1(n3093), .A2(n3094), .ZN(n2971) );
NAND2_X1 U2249 ( .A1(n2950), .A2(n2951), .ZN(n3094) );
NAND2_X1 U2250 ( .A1(n3095), .A2(n3096), .ZN(n2951) );
NAND3_X1 U2251 ( .A1(n2953), .A2(n2832), .A3(n2831), .ZN(n3096) );
XNOR2_X1 U2252 ( .A(n3097), .B(n3098), .ZN(n2832) );
NOR2_X1 U2253 ( .A1(n3099), .A2(n2793), .ZN(n3098) );
NAND2_X1 U2254 ( .A1(KEYINPUT45), .A2(n3100), .ZN(n3097) );
INV_X1 U2255 ( .A(n2863), .ZN(n3100) );
NAND2_X1 U2256 ( .A1(n3050), .A2(n3101), .ZN(n2863) );
NAND3_X1 U2257 ( .A1(n3102), .A2(n3103), .A3(n3099), .ZN(n3101) );
INV_X1 U2258 ( .A(n3104), .ZN(n3099) );
NAND2_X1 U2259 ( .A1(G200), .A2(n3105), .ZN(n3103) );
NAND2_X1 U2260 ( .A1(n3106), .A2(G190), .ZN(n3102) );
NAND2_X1 U2261 ( .A1(n3107), .A2(n2793), .ZN(n3095) );
NAND2_X1 U2262 ( .A1(n3047), .A2(n3108), .ZN(n3107) );
NAND2_X1 U2263 ( .A1(n2960), .A2(n2953), .ZN(n3108) );
XNOR2_X1 U2264 ( .A(n3049), .B(n3109), .ZN(n2953) );
NOR2_X1 U2265 ( .A1(n3110), .A2(n2793), .ZN(n3109) );
NAND2_X1 U2266 ( .A1(n3111), .A2(n3112), .ZN(n3049) );
NAND3_X1 U2267 ( .A1(n3113), .A2(n3114), .A3(n3110), .ZN(n3112) );
INV_X1 U2268 ( .A(n3115), .ZN(n3110) );
NAND2_X1 U2269 ( .A1(G200), .A2(n3116), .ZN(n3114) );
NAND2_X1 U2270 ( .A1(n3117), .A2(G190), .ZN(n3113) );
XNOR2_X1 U2271 ( .A(KEYINPUT37), .B(n3047), .ZN(n3111) );
INV_X1 U2272 ( .A(n3050), .ZN(n2960) );
NAND3_X1 U2273 ( .A1(n3118), .A2(n3119), .A3(n3104), .ZN(n3050) );
NAND3_X1 U2274 ( .A1(n3120), .A2(n3121), .A3(n3122), .ZN(n3104) );
NAND2_X1 U2275 ( .A1(n3123), .A2(n3124), .ZN(n3122) );
NAND3_X1 U2276 ( .A1(n3125), .A2(n3126), .A3(n3127), .ZN(n3124) );
NAND2_X1 U2277 ( .A1(G77), .A2(G20), .ZN(n3127) );
NAND2_X1 U2278 ( .A1(G58), .A2(n3077), .ZN(n3126) );
NAND2_X1 U2279 ( .A1(n3128), .A2(G87), .ZN(n3125) );
NAND2_X1 U2280 ( .A1(n3079), .A2(n2594), .ZN(n3121) );
NAND2_X1 U2281 ( .A1(n3080), .A2(G77), .ZN(n3120) );
NAND2_X1 U2282 ( .A1(n3106), .A2(n3081), .ZN(n3119) );
INV_X1 U2283 ( .A(n3105), .ZN(n3106) );
NAND2_X1 U2284 ( .A1(n3105), .A2(n3020), .ZN(n3118) );
NAND3_X1 U2285 ( .A1(n3129), .A2(n3083), .A3(n3130), .ZN(n3105) );
NAND2_X1 U2286 ( .A1(G244), .A2(n3085), .ZN(n3130) );
NAND2_X1 U2287 ( .A1(n3086), .A2(n3131), .ZN(n3129) );
NAND3_X1 U2288 ( .A1(n3132), .A2(n3133), .A3(n3134), .ZN(n3131) );
NAND2_X1 U2289 ( .A1(G107), .A2(G33), .ZN(n3134) );
NAND2_X1 U2290 ( .A1(G238), .A2(n3091), .ZN(n3133) );
NAND2_X1 U2291 ( .A1(G232), .A2(n3092), .ZN(n3132) );
NAND3_X1 U2292 ( .A1(n3135), .A2(n3136), .A3(n3115), .ZN(n3047) );
NAND3_X1 U2293 ( .A1(n3137), .A2(n3138), .A3(n3139), .ZN(n3115) );
NAND2_X1 U2294 ( .A1(n3140), .A2(n3141), .ZN(n3139) );
NAND3_X1 U2295 ( .A1(n3142), .A2(n3143), .A3(n3144), .ZN(n3141) );
NAND2_X1 U2296 ( .A1(G20), .A2(n2663), .ZN(n3144) );
NAND2_X1 U2297 ( .A1(n3077), .A2(G50), .ZN(n3143) );
NAND2_X1 U2298 ( .A1(n3128), .A2(G77), .ZN(n3142) );
XNOR2_X1 U2299 ( .A(n3123), .B(KEYINPUT54), .ZN(n3140) );
NAND2_X1 U2300 ( .A1(n3079), .A2(n2663), .ZN(n3138) );
NAND2_X1 U2301 ( .A1(n3080), .A2(G68), .ZN(n3137) );
NAND2_X1 U2302 ( .A1(n3117), .A2(n3081), .ZN(n3136) );
INV_X1 U2303 ( .A(n3116), .ZN(n3117) );
NAND2_X1 U2304 ( .A1(n3116), .A2(n3020), .ZN(n3135) );
NAND3_X1 U2305 ( .A1(n3145), .A2(n3083), .A3(n3146), .ZN(n3116) );
NAND2_X1 U2306 ( .A1(G238), .A2(n3085), .ZN(n3146) );
NAND2_X1 U2307 ( .A1(n3086), .A2(n3147), .ZN(n3145) );
NAND3_X1 U2308 ( .A1(n3148), .A2(n3149), .A3(n3150), .ZN(n3147) );
NAND2_X1 U2309 ( .A1(G97), .A2(G33), .ZN(n3150) );
NAND2_X1 U2310 ( .A1(G232), .A2(n3091), .ZN(n3149) );
NAND2_X1 U2311 ( .A1(n3092), .A2(G226), .ZN(n3148) );
XOR2_X1 U2312 ( .A(n3151), .B(n3152), .Z(n2950) );
NOR2_X1 U2313 ( .A1(n3153), .A2(n3154), .ZN(n3152) );
XNOR2_X1 U2314 ( .A(n3042), .B(KEYINPUT49), .ZN(n3151) );
INV_X1 U2315 ( .A(n2937), .ZN(n3042) );
NAND2_X1 U2316 ( .A1(n3155), .A2(n3156), .ZN(n2937) );
XOR2_X1 U2317 ( .A(n3157), .B(KEYINPUT59), .Z(n3155) );
NAND3_X1 U2318 ( .A1(n3158), .A2(n3159), .A3(n3153), .ZN(n3157) );
INV_X1 U2319 ( .A(n3160), .ZN(n3153) );
NAND2_X1 U2320 ( .A1(G200), .A2(n3161), .ZN(n3159) );
NAND2_X1 U2321 ( .A1(n3162), .A2(G190), .ZN(n3158) );
NAND2_X1 U2322 ( .A1(n3051), .A2(n3154), .ZN(n3093) );
INV_X1 U2323 ( .A(n3156), .ZN(n3051) );
NAND3_X1 U2324 ( .A1(n3163), .A2(n3164), .A3(n3160), .ZN(n3156) );
NAND3_X1 U2325 ( .A1(n3165), .A2(n3166), .A3(n3167), .ZN(n3160) );
NAND2_X1 U2326 ( .A1(n3123), .A2(n3168), .ZN(n3167) );
NAND3_X1 U2327 ( .A1(n3169), .A2(n3170), .A3(n3171), .ZN(n3168) );
NAND2_X1 U2328 ( .A1(n3077), .A2(G159), .ZN(n3171) );
NAND3_X1 U2329 ( .A1(n3172), .A2(G20), .A3(KEYINPUT6), .ZN(n3170) );
NAND2_X1 U2330 ( .A1(G68), .A2(n3173), .ZN(n3169) );
NAND2_X1 U2331 ( .A1(n3174), .A2(n3175), .ZN(n3173) );
NAND2_X1 U2332 ( .A1(G20), .A2(n3176), .ZN(n3175) );
NAND2_X1 U2333 ( .A1(KEYINPUT6), .A2(n2735), .ZN(n3176) );
INV_X1 U2334 ( .A(n3128), .ZN(n3174) );
NAND2_X1 U2335 ( .A1(n3079), .A2(n2735), .ZN(n3166) );
INV_X1 U2336 ( .A(G58), .ZN(n2735) );
NAND2_X1 U2337 ( .A1(n3080), .A2(G58), .ZN(n3165) );
AND3_X1 U2338 ( .A1(n3177), .A2(n3078), .A3(n3178), .ZN(n3080) );
NAND2_X1 U2339 ( .A1(n3179), .A2(n3180), .ZN(n3178) );
XNOR2_X1 U2340 ( .A(KEYINPUT44), .B(n2787), .ZN(n3179) );
NAND2_X1 U2341 ( .A1(n3162), .A2(n3081), .ZN(n3164) );
INV_X1 U2342 ( .A(n3161), .ZN(n3162) );
NAND2_X1 U2343 ( .A1(n3161), .A2(n3020), .ZN(n3163) );
NAND3_X1 U2344 ( .A1(n3181), .A2(n3083), .A3(n3182), .ZN(n3161) );
NAND2_X1 U2345 ( .A1(G232), .A2(n3085), .ZN(n3182) );
NOR2_X1 U2346 ( .A1(n3183), .A2(n3086), .ZN(n3085) );
NAND2_X1 U2347 ( .A1(G274), .A2(n3183), .ZN(n3083) );
AND2_X1 U2348 ( .A1(n3180), .A2(n3184), .ZN(n3183) );
NAND2_X1 U2349 ( .A1(n2981), .A2(n2649), .ZN(n3184) );
INV_X1 U2350 ( .A(G41), .ZN(n2981) );
NAND2_X1 U2351 ( .A1(n3086), .A2(n3185), .ZN(n3181) );
NAND3_X1 U2352 ( .A1(n3186), .A2(n3187), .A3(n3188), .ZN(n3185) );
NAND2_X1 U2353 ( .A1(G87), .A2(G33), .ZN(n3188) );
NAND2_X1 U2354 ( .A1(G226), .A2(n3091), .ZN(n3187) );
NAND2_X1 U2355 ( .A1(G223), .A2(n3092), .ZN(n3186) );
NAND3_X1 U2356 ( .A1(G116), .A2(n3189), .A3(n3190), .ZN(n3027) );
XOR2_X1 U2357 ( .A(KEYINPUT29), .B(n3191), .Z(n3189) );
NOR2_X1 U2358 ( .A1(n3192), .A2(n3193), .ZN(G364) );
NOR3_X1 U2359 ( .A1(n3194), .A2(n3195), .A3(n3196), .ZN(n3193) );
NOR3_X1 U2360 ( .A1(n2642), .A2(n2629), .A3(n3180), .ZN(n3194) );
INV_X1 U2361 ( .A(n2650), .ZN(n2642) );
NOR2_X1 U2362 ( .A1(n3197), .A2(G116), .ZN(n2650) );
NOR3_X1 U2363 ( .A1(n3196), .A2(KEYINPUT40), .A3(n3195), .ZN(n3192) );
NOR2_X1 U2364 ( .A1(n2632), .A2(G1), .ZN(n3195) );
NOR2_X1 U2365 ( .A1(n2961), .A2(n2831), .ZN(n2632) );
AND2_X1 U2366 ( .A1(n2793), .A2(n3026), .ZN(n2831) );
NAND2_X1 U2367 ( .A1(n3198), .A2(n3199), .ZN(n3026) );
NAND2_X1 U2368 ( .A1(n3200), .A2(n3201), .ZN(n3199) );
NAND2_X1 U2369 ( .A1(n2801), .A2(n3202), .ZN(n3201) );
NAND2_X1 U2370 ( .A1(n2810), .A2(n3203), .ZN(n3202) );
NAND2_X1 U2371 ( .A1(n2820), .A2(n3204), .ZN(n3203) );
OR2_X1 U2372 ( .A1(n2821), .A2(n2685), .ZN(n3204) );
INV_X1 U2373 ( .A(n3205), .ZN(n2810) );
INV_X1 U2374 ( .A(n2790), .ZN(n3200) );
AND2_X1 U2375 ( .A1(G330), .A2(n3055), .ZN(n2961) );
NAND2_X1 U2376 ( .A1(n3206), .A2(n3207), .ZN(n3055) );
NAND2_X1 U2377 ( .A1(n3021), .A2(n2793), .ZN(n3207) );
NOR4_X1 U2378 ( .A1(n2589), .A2(n2790), .A3(n3205), .A4(n2685), .ZN(n3021) );
NAND2_X1 U2379 ( .A1(n2820), .A2(n3208), .ZN(n2685) );
NAND3_X1 U2380 ( .A1(n3209), .A2(n3210), .A3(n3211), .ZN(n3208) );
INV_X1 U2381 ( .A(n2824), .ZN(n3211) );
NAND2_X1 U2382 ( .A1(G200), .A2(n3212), .ZN(n3210) );
NAND2_X1 U2383 ( .A1(n3213), .A2(G190), .ZN(n3209) );
NAND3_X1 U2384 ( .A1(n3214), .A2(n3215), .A3(n2824), .ZN(n2820) );
NAND3_X1 U2385 ( .A1(n3216), .A2(n3217), .A3(n3218), .ZN(n2824) );
NAND2_X1 U2386 ( .A1(n3123), .A2(n3219), .ZN(n3218) );
NAND3_X1 U2387 ( .A1(n3220), .A2(n3221), .A3(n3222), .ZN(n3219) );
NAND2_X1 U2388 ( .A1(n3128), .A2(G116), .ZN(n3222) );
NAND2_X1 U2389 ( .A1(n3223), .A2(G20), .ZN(n3221) );
NAND2_X1 U2390 ( .A1(n3077), .A2(G87), .ZN(n3220) );
NAND2_X1 U2391 ( .A1(n3079), .A2(n2644), .ZN(n3217) );
NAND2_X1 U2392 ( .A1(n3224), .A2(G107), .ZN(n3216) );
NAND2_X1 U2393 ( .A1(n3213), .A2(n3081), .ZN(n3215) );
NAND2_X1 U2394 ( .A1(n3212), .A2(n3020), .ZN(n3214) );
NAND2_X1 U2395 ( .A1(n2801), .A2(n3225), .ZN(n3205) );
NAND3_X1 U2396 ( .A1(n3226), .A2(n3227), .A3(n2812), .ZN(n3225) );
INV_X1 U2397 ( .A(n3228), .ZN(n2812) );
NAND2_X1 U2398 ( .A1(G200), .A2(n3229), .ZN(n3227) );
NAND2_X1 U2399 ( .A1(n3230), .A2(G190), .ZN(n3226) );
NAND3_X1 U2400 ( .A1(n3231), .A2(n3232), .A3(n3228), .ZN(n2801) );
NAND3_X1 U2401 ( .A1(n3233), .A2(n3234), .A3(n3235), .ZN(n3228) );
NAND2_X1 U2402 ( .A1(n3123), .A2(n3236), .ZN(n3235) );
NAND3_X1 U2403 ( .A1(n3237), .A2(n3238), .A3(n3239), .ZN(n3236) );
OR2_X1 U2404 ( .A1(n3191), .A2(n2787), .ZN(n3239) );
NAND3_X1 U2405 ( .A1(n3240), .A2(n3241), .A3(G77), .ZN(n3238) );
OR2_X1 U2406 ( .A1(G20), .A2(KEYINPUT15), .ZN(n3241) );
NAND2_X1 U2407 ( .A1(KEYINPUT15), .A2(n3076), .ZN(n3240) );
INV_X1 U2408 ( .A(n3077), .ZN(n3076) );
NAND2_X1 U2409 ( .A1(n3128), .A2(G107), .ZN(n3237) );
NAND2_X1 U2410 ( .A1(n3079), .A2(n2743), .ZN(n3234) );
NAND2_X1 U2411 ( .A1(n3224), .A2(G97), .ZN(n3233) );
NAND2_X1 U2412 ( .A1(n3230), .A2(n3081), .ZN(n3232) );
NAND2_X1 U2413 ( .A1(n3229), .A2(n3020), .ZN(n3231) );
NAND2_X1 U2414 ( .A1(n3198), .A2(n3242), .ZN(n2790) );
NAND3_X1 U2415 ( .A1(n3243), .A2(n3244), .A3(n2792), .ZN(n3242) );
INV_X1 U2416 ( .A(n3245), .ZN(n2792) );
NAND2_X1 U2417 ( .A1(G200), .A2(n3246), .ZN(n3244) );
NAND2_X1 U2418 ( .A1(n3247), .A2(G190), .ZN(n3243) );
NAND3_X1 U2419 ( .A1(n3248), .A2(n3249), .A3(n3245), .ZN(n3198) );
NAND3_X1 U2420 ( .A1(n3250), .A2(n3251), .A3(n3252), .ZN(n3245) );
NAND2_X1 U2421 ( .A1(n3123), .A2(n3253), .ZN(n3252) );
NAND3_X1 U2422 ( .A1(n3254), .A2(n3255), .A3(n3256), .ZN(n3253) );
NAND2_X1 U2423 ( .A1(n3128), .A2(G97), .ZN(n3256) );
NAND2_X1 U2424 ( .A1(G20), .A2(n3197), .ZN(n3255) );
NAND3_X1 U2425 ( .A1(n3257), .A2(n2734), .A3(n3223), .ZN(n3197) );
XNOR2_X1 U2426 ( .A(KEYINPUT34), .B(G107), .ZN(n3223) );
XNOR2_X1 U2427 ( .A(G97), .B(KEYINPUT57), .ZN(n3257) );
NAND2_X1 U2428 ( .A1(n3077), .A2(G68), .ZN(n3254) );
NAND2_X1 U2429 ( .A1(n3079), .A2(n2734), .ZN(n3251) );
INV_X1 U2430 ( .A(G87), .ZN(n2734) );
NAND2_X1 U2431 ( .A1(n3224), .A2(G87), .ZN(n3250) );
NAND2_X1 U2432 ( .A1(n3247), .A2(n3081), .ZN(n3249) );
INV_X1 U2433 ( .A(n3246), .ZN(n3247) );
NAND2_X1 U2434 ( .A1(n3246), .A2(n3020), .ZN(n3248) );
NAND2_X1 U2435 ( .A1(n3258), .A2(n2821), .ZN(n2589) );
NAND3_X1 U2436 ( .A1(n3259), .A2(n3260), .A3(n3261), .ZN(n2821) );
NAND2_X1 U2437 ( .A1(n3262), .A2(n3081), .ZN(n3260) );
NAND2_X1 U2438 ( .A1(n3263), .A2(n3020), .ZN(n3259) );
INV_X1 U2439 ( .A(G169), .ZN(n3020) );
NAND3_X1 U2440 ( .A1(n3264), .A2(n3265), .A3(n2817), .ZN(n3258) );
INV_X1 U2441 ( .A(n3261), .ZN(n2817) );
NAND3_X1 U2442 ( .A1(n3266), .A2(n3267), .A3(n3268), .ZN(n3261) );
NAND2_X1 U2443 ( .A1(n3123), .A2(n3269), .ZN(n3268) );
NAND3_X1 U2444 ( .A1(n3270), .A2(n3271), .A3(n3272), .ZN(n3269) );
NAND2_X1 U2445 ( .A1(n3128), .A2(G283), .ZN(n3272) );
NAND2_X1 U2446 ( .A1(G116), .A2(n3273), .ZN(n3271) );
XNOR2_X1 U2447 ( .A(KEYINPUT4), .B(n2787), .ZN(n3273) );
NAND2_X1 U2448 ( .A1(n3077), .A2(G97), .ZN(n3270) );
NOR2_X1 U2449 ( .A1(n3128), .A2(G20), .ZN(n3077) );
NOR2_X1 U2450 ( .A1(n2724), .A2(G20), .ZN(n3128) );
INV_X1 U2451 ( .A(n3078), .ZN(n3123) );
NAND2_X1 U2452 ( .A1(n3079), .A2(n2587), .ZN(n3267) );
NAND2_X1 U2453 ( .A1(n3224), .A2(G116), .ZN(n3266) );
AND3_X1 U2454 ( .A1(n3177), .A2(n3078), .A3(n3274), .ZN(n3224) );
NAND2_X1 U2455 ( .A1(G33), .A2(n3180), .ZN(n3274) );
NAND2_X1 U2456 ( .A1(G1), .A2(n3275), .ZN(n3078) );
NAND2_X1 U2457 ( .A1(n3031), .A2(n3276), .ZN(n3275) );
NAND2_X1 U2458 ( .A1(G20), .A2(n3277), .ZN(n3276) );
XNOR2_X1 U2459 ( .A(KEYINPUT17), .B(n2724), .ZN(n3277) );
INV_X1 U2460 ( .A(n3079), .ZN(n3177) );
NAND2_X1 U2461 ( .A1(G200), .A2(n3263), .ZN(n3265) );
NAND2_X1 U2462 ( .A1(n3262), .A2(G190), .ZN(n3264) );
NAND2_X1 U2463 ( .A1(n3278), .A2(n2802), .ZN(n3206) );
INV_X1 U2464 ( .A(n2793), .ZN(n2802) );
NAND2_X1 U2465 ( .A1(G343), .A2(n2969), .ZN(n2793) );
INV_X1 U2466 ( .A(n3154), .ZN(n2969) );
NAND4_X1 U2467 ( .A1(G213), .A2(G13), .A3(n3180), .A4(n2787), .ZN(n3154) );
NAND2_X1 U2468 ( .A1(n3279), .A2(n3280), .ZN(n3278) );
NAND4_X1 U2469 ( .A1(n3246), .A2(n3263), .A3(n3281), .A4(n3081), .ZN(n3280) );
INV_X1 U2470 ( .A(G179), .ZN(n3081) );
NOR2_X1 U2471 ( .A1(n3230), .A2(n3282), .ZN(n3281) );
XNOR2_X1 U2472 ( .A(KEYINPUT12), .B(n3212), .ZN(n3282) );
INV_X1 U2473 ( .A(n3229), .ZN(n3230) );
NAND4_X1 U2474 ( .A1(n3213), .A2(n3262), .A3(n3283), .A4(G179), .ZN(n3279) );
NOR2_X1 U2475 ( .A1(n3246), .A2(n3229), .ZN(n3283) );
NAND3_X1 U2476 ( .A1(n3284), .A2(n3285), .A3(n3286), .ZN(n3229) );
NAND2_X1 U2477 ( .A1(n3086), .A2(n3287), .ZN(n3286) );
NAND3_X1 U2478 ( .A1(n3288), .A2(n3289), .A3(n3290), .ZN(n3287) );
NAND2_X1 U2479 ( .A1(G283), .A2(G33), .ZN(n3290) );
NAND2_X1 U2480 ( .A1(n3291), .A2(n3092), .ZN(n3289) );
XNOR2_X1 U2481 ( .A(G244), .B(KEYINPUT61), .ZN(n3291) );
NAND2_X1 U2482 ( .A1(G250), .A2(n3091), .ZN(n3288) );
NAND2_X1 U2483 ( .A1(G257), .A2(n3292), .ZN(n3284) );
NAND3_X1 U2484 ( .A1(n3293), .A2(n3294), .A3(n3295), .ZN(n3246) );
NAND2_X1 U2485 ( .A1(n3086), .A2(n3296), .ZN(n3295) );
NAND3_X1 U2486 ( .A1(n3297), .A2(n3298), .A3(n3299), .ZN(n3296) );
XOR2_X1 U2487 ( .A(KEYINPUT41), .B(n3300), .Z(n3299) );
NOR2_X1 U2488 ( .A1(n2724), .A2(n2587), .ZN(n3300) );
INV_X1 U2489 ( .A(G116), .ZN(n2587) );
INV_X1 U2490 ( .A(G33), .ZN(n2724) );
NAND2_X1 U2491 ( .A1(G244), .A2(n3091), .ZN(n3298) );
NAND2_X1 U2492 ( .A1(G238), .A2(n3092), .ZN(n3297) );
NAND3_X1 U2493 ( .A1(G250), .A2(n3301), .A3(n3302), .ZN(n3294) );
NAND2_X1 U2494 ( .A1(n3303), .A2(G274), .ZN(n3293) );
INV_X1 U2495 ( .A(n3263), .ZN(n3262) );
NAND3_X1 U2496 ( .A1(n3304), .A2(n3285), .A3(n3305), .ZN(n3263) );
NAND2_X1 U2497 ( .A1(n3086), .A2(n3306), .ZN(n3305) );
NAND3_X1 U2498 ( .A1(n3307), .A2(n3308), .A3(n3309), .ZN(n3306) );
NAND2_X1 U2499 ( .A1(G303), .A2(G33), .ZN(n3309) );
NAND2_X1 U2500 ( .A1(G264), .A2(n3091), .ZN(n3308) );
NAND2_X1 U2501 ( .A1(G257), .A2(n3092), .ZN(n3307) );
NAND2_X1 U2502 ( .A1(G270), .A2(n3292), .ZN(n3304) );
INV_X1 U2503 ( .A(n3212), .ZN(n3213) );
NAND3_X1 U2504 ( .A1(n3310), .A2(n3285), .A3(n3311), .ZN(n3212) );
NAND2_X1 U2505 ( .A1(n3086), .A2(n3312), .ZN(n3311) );
NAND3_X1 U2506 ( .A1(n3313), .A2(n3314), .A3(n3315), .ZN(n3312) );
NAND2_X1 U2507 ( .A1(G294), .A2(G33), .ZN(n3315) );
NAND2_X1 U2508 ( .A1(G257), .A2(n3091), .ZN(n3314) );
NOR2_X1 U2509 ( .A1(n3092), .A2(G33), .ZN(n3091) );
NAND2_X1 U2510 ( .A1(G250), .A2(n3092), .ZN(n3313) );
NOR2_X1 U2511 ( .A1(G33), .A2(G1698), .ZN(n3092) );
NAND2_X1 U2512 ( .A1(n3316), .A2(G274), .ZN(n3285) );
NAND2_X1 U2513 ( .A1(G264), .A2(n3292), .ZN(n3310) );
NOR2_X1 U2514 ( .A1(n3316), .A2(n3086), .ZN(n3292) );
INV_X1 U2515 ( .A(n3301), .ZN(n3086) );
NAND3_X1 U2516 ( .A1(G1), .A2(n3317), .A3(G13), .ZN(n3301) );
NAND2_X1 U2517 ( .A1(G41), .A2(G33), .ZN(n3317) );
NOR2_X1 U2518 ( .A1(n3302), .A2(G41), .ZN(n3316) );
INV_X1 U2519 ( .A(n3303), .ZN(n3302) );
NOR2_X1 U2520 ( .A1(n2649), .A2(G1), .ZN(n3303) );
INV_X1 U2521 ( .A(G45), .ZN(n2649) );
AND2_X1 U2522 ( .A1(n2583), .A2(n2629), .ZN(n3196) );
NOR2_X1 U2523 ( .A1(n2783), .A2(G41), .ZN(n2629) );
NOR3_X1 U2524 ( .A1(n3318), .A2(n3319), .A3(n3320), .ZN(G361) );
NOR3_X1 U2525 ( .A1(n2783), .A2(n3321), .A3(n3322), .ZN(n3320) );
NOR2_X1 U2526 ( .A1(G264), .A2(n3323), .ZN(n3321) );
XOR2_X1 U2527 ( .A(KEYINPUT38), .B(G257), .Z(n3323) );
INV_X1 U2528 ( .A(n3324), .ZN(n2783) );
NOR3_X1 U2529 ( .A1(n3324), .A2(n3190), .A3(n3325), .ZN(n3319) );
NOR2_X1 U2530 ( .A1(n3326), .A2(n3327), .ZN(n3325) );
NAND4_X1 U2531 ( .A1(n3328), .A2(n3329), .A3(n3330), .A4(n3331), .ZN(n3327) );
NAND2_X1 U2532 ( .A1(G238), .A2(G68), .ZN(n3331) );
NAND2_X1 U2533 ( .A1(G244), .A2(G77), .ZN(n3330) );
NAND2_X1 U2534 ( .A1(G250), .A2(G87), .ZN(n3329) );
NAND2_X1 U2535 ( .A1(G257), .A2(G97), .ZN(n3328) );
NAND4_X1 U2536 ( .A1(n3332), .A2(n3333), .A3(n3334), .A4(n3335), .ZN(n3326) );
NAND2_X1 U2537 ( .A1(G264), .A2(G107), .ZN(n3335) );
NAND2_X1 U2538 ( .A1(G270), .A2(G116), .ZN(n3334) );
NAND2_X1 U2539 ( .A1(G226), .A2(G50), .ZN(n3333) );
NAND2_X1 U2540 ( .A1(G232), .A2(G58), .ZN(n3332) );
NOR3_X1 U2541 ( .A1(n3180), .A2(G13), .A3(n2787), .ZN(n3324) );
NOR2_X1 U2542 ( .A1(n3336), .A2(n3337), .ZN(n3318) );
XNOR2_X1 U2543 ( .A(KEYINPUT50), .B(n3036), .ZN(n3337) );
INV_X1 U2544 ( .A(n3190), .ZN(n3036) );
NOR3_X1 U2545 ( .A1(n2787), .A2(n3180), .A3(n3031), .ZN(n3190) );
INV_X1 U2546 ( .A(G13), .ZN(n3031) );
INV_X1 U2547 ( .A(G1), .ZN(n3180) );
INV_X1 U2548 ( .A(G20), .ZN(n2787) );
INV_X1 U2549 ( .A(n2583), .ZN(n3336) );
NOR2_X1 U2550 ( .A1(n2597), .A2(n3172), .ZN(n2583) );
XOR2_X1 U2551 ( .A(n2782), .B(n3338), .Z(G358) );
XOR2_X1 U2552 ( .A(n3339), .B(n2656), .Z(n3338) );
XOR2_X1 U2553 ( .A(G238), .B(G244), .Z(n2656) );
NOR2_X1 U2554 ( .A1(KEYINPUT56), .A2(n2654), .ZN(n3339) );
XNOR2_X1 U2555 ( .A(G226), .B(G232), .ZN(n2654) );
XOR2_X1 U2556 ( .A(n3340), .B(n3341), .Z(n2782) );
XNOR2_X1 U2557 ( .A(G257), .B(n3322), .ZN(n3341) );
INV_X1 U2558 ( .A(G250), .ZN(n3322) );
XNOR2_X1 U2559 ( .A(G270), .B(G264), .ZN(n3340) );
NAND2_X1 U2560 ( .A1(G87), .A2(n3342), .ZN(G355) );
NAND2_X1 U2561 ( .A1(n2644), .A2(n2743), .ZN(n3342) );
INV_X1 U2562 ( .A(G107), .ZN(n2644) );
AND3_X1 U2563 ( .A1(n3172), .A2(n2594), .A3(n2597), .ZN(G353) );
NOR2_X1 U2564 ( .A1(G58), .A2(G68), .ZN(n3172) );
XNOR2_X1 U2565 ( .A(n2582), .B(n2744), .ZN(G351) );
XNOR2_X1 U2566 ( .A(n3343), .B(n3191), .ZN(n2744) );
XNOR2_X1 U2567 ( .A(G107), .B(n2743), .ZN(n3191) );
INV_X1 U2568 ( .A(G97), .ZN(n2743) );
XNOR2_X1 U2569 ( .A(G116), .B(G87), .ZN(n3343) );
NAND3_X1 U2570 ( .A1(n3344), .A2(n3345), .A3(n3032), .ZN(n2582) );
NAND3_X1 U2571 ( .A1(G77), .A2(n3346), .A3(G50), .ZN(n3032) );
NAND2_X1 U2572 ( .A1(n3347), .A2(n2594), .ZN(n3345) );
XNOR2_X1 U2573 ( .A(n2597), .B(n3346), .ZN(n3347) );
INV_X1 U2574 ( .A(G50), .ZN(n2597) );
OR3_X1 U2575 ( .A1(n3346), .A2(G50), .A3(n2594), .ZN(n3344) );
INV_X1 U2576 ( .A(G77), .ZN(n2594) );
XNOR2_X1 U2577 ( .A(G58), .B(n2663), .ZN(n3346) );
INV_X1 U2578 ( .A(G68), .ZN(n2663) );
endmodule


