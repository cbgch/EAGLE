//Key = 1110011000110100100001101001010100100111100110101101100101010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341;

XNOR2_X1 U741 ( .A(G107), .B(n1023), .ZN(G9) );
NOR2_X1 U742 ( .A1(n1024), .A2(n1025), .ZN(G75) );
NOR2_X1 U743 ( .A1(G952), .A2(n1026), .ZN(n1025) );
NOR4_X1 U744 ( .A1(n1027), .A2(n1028), .A3(n1026), .A4(n1029), .ZN(n1024) );
NAND2_X1 U745 ( .A1(n1030), .A2(n1031), .ZN(n1026) );
NAND4_X1 U746 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
NOR4_X1 U747 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
XNOR2_X1 U748 ( .A(KEYINPUT20), .B(n1040), .ZN(n1039) );
XOR2_X1 U749 ( .A(KEYINPUT8), .B(n1041), .Z(n1038) );
NOR3_X1 U750 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1034) );
INV_X1 U751 ( .A(n1045), .ZN(n1044) );
NAND2_X1 U752 ( .A1(n1046), .A2(n1047), .ZN(n1033) );
XOR2_X1 U753 ( .A(KEYINPUT25), .B(G475), .Z(n1046) );
NOR3_X1 U754 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1028) );
AND2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U756 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1049) );
NOR2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR3_X1 U758 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1056) );
AND2_X1 U759 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U760 ( .A1(n1063), .A2(n1064), .ZN(n1059) );
XNOR2_X1 U761 ( .A(KEYINPUT2), .B(n1065), .ZN(n1064) );
INV_X1 U762 ( .A(n1066), .ZN(n1063) );
NOR2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1058) );
NOR3_X1 U764 ( .A1(n1068), .A2(n1069), .A3(n1065), .ZN(n1054) );
NOR2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR2_X1 U766 ( .A1(n1045), .A2(n1037), .ZN(n1071) );
NOR2_X1 U767 ( .A1(KEYINPUT7), .A2(n1072), .ZN(n1070) );
NOR2_X1 U768 ( .A1(n1073), .A2(n1051), .ZN(n1053) );
INV_X1 U769 ( .A(KEYINPUT7), .ZN(n1051) );
NOR4_X1 U770 ( .A1(n1072), .A2(n1065), .A3(n1068), .A4(n1052), .ZN(n1073) );
NOR4_X1 U771 ( .A1(n1074), .A2(n1057), .A3(n1068), .A4(n1052), .ZN(n1027) );
INV_X1 U772 ( .A(n1075), .ZN(n1068) );
NOR2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XNOR2_X1 U775 ( .A(KEYINPUT38), .B(n1048), .ZN(n1079) );
INV_X1 U776 ( .A(n1080), .ZN(n1048) );
NOR2_X1 U777 ( .A1(n1081), .A2(n1065), .ZN(n1076) );
NOR2_X1 U778 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U779 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
XOR2_X1 U780 ( .A(n1086), .B(n1087), .Z(G72) );
XOR2_X1 U781 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U782 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U783 ( .A1(G953), .A2(n1092), .ZN(n1091) );
XNOR2_X1 U784 ( .A(KEYINPUT37), .B(n1093), .ZN(n1092) );
XOR2_X1 U785 ( .A(n1094), .B(n1095), .Z(n1090) );
XNOR2_X1 U786 ( .A(n1096), .B(n1097), .ZN(n1095) );
INV_X1 U787 ( .A(n1098), .ZN(n1097) );
NAND2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1096) );
NAND3_X1 U789 ( .A1(G134), .A2(n1101), .A3(KEYINPUT31), .ZN(n1100) );
NAND3_X1 U790 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
NAND2_X1 U791 ( .A1(G131), .A2(n1105), .ZN(n1103) );
OR2_X1 U792 ( .A1(n1106), .A2(n1105), .ZN(n1102) );
NAND4_X1 U793 ( .A1(n1107), .A2(n1106), .A3(n1108), .A4(n1109), .ZN(n1099) );
NAND2_X1 U794 ( .A1(n1110), .A2(n1105), .ZN(n1109) );
OR2_X1 U795 ( .A1(n1104), .A2(n1105), .ZN(n1108) );
INV_X1 U796 ( .A(KEYINPUT62), .ZN(n1105) );
NAND2_X1 U797 ( .A1(KEYINPUT31), .A2(G134), .ZN(n1107) );
NAND2_X1 U798 ( .A1(n1111), .A2(n1112), .ZN(n1088) );
XNOR2_X1 U799 ( .A(G953), .B(KEYINPUT17), .ZN(n1111) );
NOR2_X1 U800 ( .A1(n1113), .A2(n1030), .ZN(n1086) );
AND2_X1 U801 ( .A1(G227), .A2(G900), .ZN(n1113) );
XOR2_X1 U802 ( .A(n1114), .B(n1115), .Z(G69) );
XOR2_X1 U803 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U805 ( .A1(G953), .A2(n1120), .ZN(n1119) );
XOR2_X1 U806 ( .A(KEYINPUT44), .B(n1121), .Z(n1118) );
NAND2_X1 U807 ( .A1(n1122), .A2(n1030), .ZN(n1116) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1030), .ZN(n1114) );
AND2_X1 U809 ( .A1(G224), .A2(G898), .ZN(n1123) );
NOR2_X1 U810 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XOR2_X1 U811 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U812 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U813 ( .A1(KEYINPUT21), .A2(n1130), .ZN(n1126) );
NOR2_X1 U814 ( .A1(n1124), .A2(n1131), .ZN(G63) );
XOR2_X1 U815 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND3_X1 U816 ( .A1(n1134), .A2(n1029), .A3(G478), .ZN(n1132) );
XOR2_X1 U817 ( .A(KEYINPUT19), .B(n1135), .Z(n1134) );
NOR2_X1 U818 ( .A1(n1124), .A2(n1136), .ZN(G60) );
XOR2_X1 U819 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U820 ( .A1(n1139), .A2(G475), .ZN(n1137) );
XNOR2_X1 U821 ( .A(G104), .B(n1140), .ZN(G6) );
NAND3_X1 U822 ( .A1(n1141), .A2(n1062), .A3(n1142), .ZN(n1140) );
NOR3_X1 U823 ( .A1(n1065), .A2(n1143), .A3(n1144), .ZN(n1142) );
INV_X1 U824 ( .A(n1061), .ZN(n1065) );
XNOR2_X1 U825 ( .A(n1145), .B(KEYINPUT61), .ZN(n1141) );
NOR2_X1 U826 ( .A1(n1146), .A2(n1147), .ZN(G57) );
XOR2_X1 U827 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U828 ( .A(n1150), .B(n1151), .ZN(n1149) );
XOR2_X1 U829 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U830 ( .A1(KEYINPUT40), .A2(n1154), .ZN(n1152) );
XOR2_X1 U831 ( .A(n1155), .B(n1156), .Z(n1148) );
NOR2_X1 U832 ( .A1(G101), .A2(n1157), .ZN(n1156) );
XOR2_X1 U833 ( .A(KEYINPUT29), .B(KEYINPUT0), .Z(n1157) );
XOR2_X1 U834 ( .A(n1158), .B(KEYINPUT3), .Z(n1155) );
NAND2_X1 U835 ( .A1(n1139), .A2(G472), .ZN(n1158) );
NOR2_X1 U836 ( .A1(n1159), .A2(n1030), .ZN(n1146) );
XNOR2_X1 U837 ( .A(G952), .B(KEYINPUT57), .ZN(n1159) );
NOR2_X1 U838 ( .A1(n1124), .A2(n1160), .ZN(G54) );
XOR2_X1 U839 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U840 ( .A(n1150), .B(n1163), .ZN(n1162) );
XOR2_X1 U841 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U842 ( .A1(n1139), .A2(G469), .ZN(n1165) );
NAND2_X1 U843 ( .A1(KEYINPUT6), .A2(n1166), .ZN(n1164) );
XNOR2_X1 U844 ( .A(n1098), .B(n1167), .ZN(n1166) );
XNOR2_X1 U845 ( .A(KEYINPUT41), .B(n1168), .ZN(n1167) );
NOR2_X1 U846 ( .A1(KEYINPUT9), .A2(n1169), .ZN(n1168) );
XOR2_X1 U847 ( .A(n1170), .B(n1171), .Z(n1161) );
XOR2_X1 U848 ( .A(G110), .B(n1172), .Z(n1171) );
XNOR2_X1 U849 ( .A(G140), .B(KEYINPUT58), .ZN(n1170) );
NOR2_X1 U850 ( .A1(n1030), .A2(G952), .ZN(n1124) );
NOR2_X1 U851 ( .A1(n1173), .A2(n1174), .ZN(G51) );
XOR2_X1 U852 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U853 ( .A(n1177), .B(n1178), .ZN(n1176) );
NAND2_X1 U854 ( .A1(KEYINPUT13), .A2(n1154), .ZN(n1177) );
XNOR2_X1 U855 ( .A(n1179), .B(n1180), .ZN(n1175) );
NAND2_X1 U856 ( .A1(n1139), .A2(n1181), .ZN(n1179) );
INV_X1 U857 ( .A(n1129), .ZN(n1139) );
NAND2_X1 U858 ( .A1(n1135), .A2(n1029), .ZN(n1129) );
OR2_X1 U859 ( .A1(n1112), .A2(n1122), .ZN(n1029) );
NAND4_X1 U860 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1122) );
AND4_X1 U861 ( .A1(n1186), .A2(n1187), .A3(n1023), .A4(n1188), .ZN(n1185) );
NAND3_X1 U862 ( .A1(n1061), .A2(n1189), .A3(n1066), .ZN(n1023) );
NAND2_X1 U863 ( .A1(n1062), .A2(n1190), .ZN(n1184) );
NAND2_X1 U864 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NAND2_X1 U865 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XNOR2_X1 U866 ( .A(KEYINPUT12), .B(n1078), .ZN(n1194) );
NAND2_X1 U867 ( .A1(n1061), .A2(n1189), .ZN(n1191) );
NAND4_X1 U868 ( .A1(n1193), .A2(n1061), .A3(n1195), .A4(n1196), .ZN(n1182) );
NAND4_X1 U869 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1112) );
NOR4_X1 U870 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
NAND2_X1 U871 ( .A1(n1205), .A2(n1206), .ZN(n1199) );
NAND2_X1 U872 ( .A1(n1207), .A2(n1078), .ZN(n1206) );
XNOR2_X1 U873 ( .A(KEYINPUT24), .B(n1067), .ZN(n1207) );
INV_X1 U874 ( .A(n1208), .ZN(n1205) );
XNOR2_X1 U875 ( .A(n1209), .B(KEYINPUT32), .ZN(n1135) );
NOR2_X1 U876 ( .A1(n1210), .A2(n1030), .ZN(n1173) );
XNOR2_X1 U877 ( .A(G952), .B(KEYINPUT1), .ZN(n1210) );
XNOR2_X1 U878 ( .A(G146), .B(n1197), .ZN(G48) );
NAND3_X1 U879 ( .A1(n1062), .A2(n1083), .A3(n1211), .ZN(n1197) );
XNOR2_X1 U880 ( .A(G143), .B(n1198), .ZN(G45) );
NAND4_X1 U881 ( .A1(n1212), .A2(n1083), .A3(n1195), .A4(n1196), .ZN(n1198) );
XOR2_X1 U882 ( .A(G140), .B(n1213), .Z(G42) );
NOR2_X1 U883 ( .A1(n1067), .A2(n1208), .ZN(n1213) );
XOR2_X1 U884 ( .A(G137), .B(n1204), .Z(G39) );
AND3_X1 U885 ( .A1(n1080), .A2(n1211), .A3(n1075), .ZN(n1204) );
XNOR2_X1 U886 ( .A(n1214), .B(n1203), .ZN(G36) );
AND3_X1 U887 ( .A1(n1080), .A2(n1066), .A3(n1212), .ZN(n1203) );
NOR3_X1 U888 ( .A1(n1072), .A2(n1215), .A3(n1078), .ZN(n1212) );
XNOR2_X1 U889 ( .A(n1110), .B(n1216), .ZN(G33) );
NOR2_X1 U890 ( .A1(n1078), .A2(n1208), .ZN(n1216) );
NAND4_X1 U891 ( .A1(n1080), .A2(n1062), .A3(n1145), .A4(n1217), .ZN(n1208) );
NOR2_X1 U892 ( .A1(n1084), .A2(n1042), .ZN(n1080) );
INV_X1 U893 ( .A(n1085), .ZN(n1042) );
INV_X1 U894 ( .A(n1218), .ZN(n1078) );
XOR2_X1 U895 ( .A(G128), .B(n1202), .Z(G30) );
AND3_X1 U896 ( .A1(n1066), .A2(n1083), .A3(n1211), .ZN(n1202) );
AND4_X1 U897 ( .A1(n1145), .A2(n1041), .A3(n1219), .A4(n1217), .ZN(n1211) );
INV_X1 U898 ( .A(n1072), .ZN(n1145) );
XNOR2_X1 U899 ( .A(G101), .B(n1187), .ZN(G3) );
NAND3_X1 U900 ( .A1(n1218), .A2(n1189), .A3(n1075), .ZN(n1187) );
NAND2_X1 U901 ( .A1(n1220), .A2(n1221), .ZN(G27) );
NAND2_X1 U902 ( .A1(n1222), .A2(n1180), .ZN(n1221) );
INV_X1 U903 ( .A(G125), .ZN(n1180) );
NAND2_X1 U904 ( .A1(G125), .A2(n1223), .ZN(n1220) );
NAND2_X1 U905 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NAND2_X1 U906 ( .A1(KEYINPUT18), .A2(n1201), .ZN(n1225) );
OR2_X1 U907 ( .A1(n1222), .A2(KEYINPUT18), .ZN(n1224) );
AND2_X1 U908 ( .A1(KEYINPUT11), .A2(n1201), .ZN(n1222) );
AND4_X1 U909 ( .A1(n1226), .A2(n1062), .A3(n1227), .A4(n1228), .ZN(n1201) );
NOR2_X1 U910 ( .A1(n1215), .A2(n1144), .ZN(n1227) );
INV_X1 U911 ( .A(n1217), .ZN(n1215) );
NAND2_X1 U912 ( .A1(n1052), .A2(n1229), .ZN(n1217) );
NAND4_X1 U913 ( .A1(G902), .A2(G953), .A3(n1230), .A4(n1093), .ZN(n1229) );
INV_X1 U914 ( .A(G900), .ZN(n1093) );
XNOR2_X1 U915 ( .A(G122), .B(n1231), .ZN(G24) );
NAND4_X1 U916 ( .A1(n1228), .A2(n1061), .A3(n1232), .A4(n1233), .ZN(n1231) );
NOR3_X1 U917 ( .A1(n1040), .A2(n1234), .A3(n1143), .ZN(n1233) );
XNOR2_X1 U918 ( .A(n1083), .B(KEYINPUT49), .ZN(n1232) );
INV_X1 U919 ( .A(n1144), .ZN(n1083) );
NOR2_X1 U920 ( .A1(n1219), .A2(n1041), .ZN(n1061) );
INV_X1 U921 ( .A(n1057), .ZN(n1228) );
XNOR2_X1 U922 ( .A(G119), .B(n1183), .ZN(G21) );
NAND4_X1 U923 ( .A1(n1193), .A2(n1075), .A3(n1041), .A4(n1219), .ZN(n1183) );
XNOR2_X1 U924 ( .A(G116), .B(n1188), .ZN(G18) );
NAND2_X1 U925 ( .A1(n1235), .A2(n1066), .ZN(n1188) );
NOR2_X1 U926 ( .A1(n1196), .A2(n1040), .ZN(n1066) );
INV_X1 U927 ( .A(n1195), .ZN(n1040) );
XNOR2_X1 U928 ( .A(G113), .B(n1236), .ZN(G15) );
NAND2_X1 U929 ( .A1(n1235), .A2(n1062), .ZN(n1236) );
NOR2_X1 U930 ( .A1(n1195), .A2(n1234), .ZN(n1062) );
AND2_X1 U931 ( .A1(n1193), .A2(n1218), .ZN(n1235) );
NOR2_X1 U932 ( .A1(n1041), .A2(n1032), .ZN(n1218) );
NOR3_X1 U933 ( .A1(n1144), .A2(n1143), .A3(n1057), .ZN(n1193) );
NAND2_X1 U934 ( .A1(n1237), .A2(n1238), .ZN(n1057) );
INV_X1 U935 ( .A(n1037), .ZN(n1237) );
XOR2_X1 U936 ( .A(n1186), .B(n1239), .Z(G12) );
NOR2_X1 U937 ( .A1(G110), .A2(KEYINPUT14), .ZN(n1239) );
NAND3_X1 U938 ( .A1(n1226), .A2(n1189), .A3(n1075), .ZN(n1186) );
NOR2_X1 U939 ( .A1(n1195), .A2(n1196), .ZN(n1075) );
INV_X1 U940 ( .A(n1234), .ZN(n1196) );
NOR2_X1 U941 ( .A1(n1240), .A2(n1043), .ZN(n1234) );
NOR2_X1 U942 ( .A1(n1047), .A2(G475), .ZN(n1043) );
AND2_X1 U943 ( .A1(G475), .A2(n1047), .ZN(n1240) );
NAND2_X1 U944 ( .A1(n1138), .A2(n1209), .ZN(n1047) );
XOR2_X1 U945 ( .A(n1241), .B(n1242), .Z(n1138) );
XOR2_X1 U946 ( .A(G113), .B(n1243), .Z(n1242) );
XNOR2_X1 U947 ( .A(KEYINPUT43), .B(n1244), .ZN(n1243) );
XNOR2_X1 U948 ( .A(n1245), .B(n1246), .ZN(n1241) );
INV_X1 U949 ( .A(G104), .ZN(n1246) );
NAND2_X1 U950 ( .A1(n1247), .A2(n1248), .ZN(n1245) );
NAND2_X1 U951 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
XOR2_X1 U952 ( .A(n1251), .B(KEYINPUT53), .Z(n1247) );
OR2_X1 U953 ( .A1(n1250), .A2(n1249), .ZN(n1251) );
XOR2_X1 U954 ( .A(n1094), .B(n1252), .Z(n1249) );
NOR2_X1 U955 ( .A1(G146), .A2(KEYINPUT23), .ZN(n1252) );
XNOR2_X1 U956 ( .A(n1253), .B(n1254), .ZN(n1250) );
XNOR2_X1 U957 ( .A(n1255), .B(G131), .ZN(n1254) );
INV_X1 U958 ( .A(G143), .ZN(n1255) );
NAND2_X1 U959 ( .A1(G214), .A2(n1256), .ZN(n1253) );
XNOR2_X1 U960 ( .A(n1257), .B(G478), .ZN(n1195) );
NAND2_X1 U961 ( .A1(n1133), .A2(n1209), .ZN(n1257) );
XOR2_X1 U962 ( .A(n1258), .B(n1259), .Z(n1133) );
NOR2_X1 U963 ( .A1(KEYINPUT35), .A2(n1260), .ZN(n1259) );
XOR2_X1 U964 ( .A(n1261), .B(n1262), .Z(n1260) );
XNOR2_X1 U965 ( .A(n1263), .B(n1264), .ZN(n1262) );
NOR2_X1 U966 ( .A1(G134), .A2(KEYINPUT45), .ZN(n1264) );
NAND2_X1 U967 ( .A1(KEYINPUT48), .A2(n1265), .ZN(n1263) );
NAND2_X1 U968 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NAND2_X1 U969 ( .A1(G107), .A2(n1268), .ZN(n1267) );
XOR2_X1 U970 ( .A(KEYINPUT63), .B(n1269), .Z(n1266) );
NOR2_X1 U971 ( .A1(G107), .A2(n1268), .ZN(n1269) );
XNOR2_X1 U972 ( .A(n1244), .B(G116), .ZN(n1268) );
INV_X1 U973 ( .A(G122), .ZN(n1244) );
NAND2_X1 U974 ( .A1(G217), .A2(n1270), .ZN(n1258) );
NOR3_X1 U975 ( .A1(n1144), .A2(n1143), .A3(n1072), .ZN(n1189) );
NAND2_X1 U976 ( .A1(n1238), .A2(n1037), .ZN(n1072) );
XNOR2_X1 U977 ( .A(n1271), .B(G469), .ZN(n1037) );
NAND2_X1 U978 ( .A1(n1272), .A2(n1209), .ZN(n1271) );
XOR2_X1 U979 ( .A(n1273), .B(n1274), .Z(n1272) );
NOR3_X1 U980 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1274) );
NOR2_X1 U981 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
INV_X1 U982 ( .A(KEYINPUT33), .ZN(n1279) );
NOR2_X1 U983 ( .A1(n1172), .A2(n1280), .ZN(n1278) );
NOR3_X1 U984 ( .A1(KEYINPUT33), .A2(n1281), .A3(n1280), .ZN(n1276) );
AND2_X1 U985 ( .A1(n1172), .A2(KEYINPUT46), .ZN(n1281) );
AND3_X1 U986 ( .A1(KEYINPUT46), .A2(n1280), .A3(n1172), .ZN(n1275) );
AND2_X1 U987 ( .A1(G227), .A2(n1282), .ZN(n1172) );
XOR2_X1 U988 ( .A(G140), .B(n1283), .Z(n1280) );
NOR2_X1 U989 ( .A1(G110), .A2(KEYINPUT42), .ZN(n1283) );
NAND2_X1 U990 ( .A1(n1284), .A2(n1285), .ZN(n1273) );
NAND2_X1 U991 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XNOR2_X1 U992 ( .A(n1150), .B(KEYINPUT39), .ZN(n1287) );
XOR2_X1 U993 ( .A(KEYINPUT27), .B(n1288), .Z(n1284) );
NOR2_X1 U994 ( .A1(n1150), .A2(n1286), .ZN(n1288) );
XOR2_X1 U995 ( .A(n1289), .B(n1169), .Z(n1286) );
NOR2_X1 U996 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NOR2_X1 U997 ( .A1(KEYINPUT59), .A2(n1292), .ZN(n1291) );
NOR2_X1 U998 ( .A1(KEYINPUT28), .A2(n1293), .ZN(n1290) );
INV_X1 U999 ( .A(n1292), .ZN(n1293) );
XOR2_X1 U1000 ( .A(n1098), .B(KEYINPUT51), .Z(n1292) );
XNOR2_X1 U1001 ( .A(n1294), .B(n1154), .ZN(n1098) );
XNOR2_X1 U1002 ( .A(KEYINPUT60), .B(KEYINPUT56), .ZN(n1294) );
INV_X1 U1003 ( .A(n1295), .ZN(n1150) );
XOR2_X1 U1004 ( .A(n1045), .B(KEYINPUT50), .Z(n1238) );
NAND2_X1 U1005 ( .A1(G221), .A2(n1296), .ZN(n1045) );
AND2_X1 U1006 ( .A1(n1297), .A2(n1052), .ZN(n1143) );
NAND3_X1 U1007 ( .A1(n1230), .A2(n1030), .A3(G952), .ZN(n1052) );
INV_X1 U1008 ( .A(G953), .ZN(n1030) );
NAND4_X1 U1009 ( .A1(G902), .A2(G953), .A3(n1230), .A4(n1120), .ZN(n1297) );
INV_X1 U1010 ( .A(G898), .ZN(n1120) );
NAND2_X1 U1011 ( .A1(G237), .A2(G234), .ZN(n1230) );
NAND2_X1 U1012 ( .A1(n1084), .A2(n1085), .ZN(n1144) );
NAND2_X1 U1013 ( .A1(G214), .A2(n1298), .ZN(n1085) );
XOR2_X1 U1014 ( .A(n1036), .B(KEYINPUT15), .Z(n1084) );
XNOR2_X1 U1015 ( .A(n1299), .B(n1181), .ZN(n1036) );
AND2_X1 U1016 ( .A1(G210), .A2(n1298), .ZN(n1181) );
NAND2_X1 U1017 ( .A1(n1300), .A2(n1209), .ZN(n1298) );
NAND2_X1 U1018 ( .A1(n1301), .A2(n1209), .ZN(n1299) );
XNOR2_X1 U1019 ( .A(n1302), .B(n1303), .ZN(n1301) );
XNOR2_X1 U1020 ( .A(n1304), .B(KEYINPUT34), .ZN(n1303) );
NAND2_X1 U1021 ( .A1(n1305), .A2(KEYINPUT10), .ZN(n1304) );
XNOR2_X1 U1022 ( .A(G125), .B(n1154), .ZN(n1305) );
INV_X1 U1023 ( .A(n1178), .ZN(n1302) );
XNOR2_X1 U1024 ( .A(n1306), .B(n1121), .ZN(n1178) );
XNOR2_X1 U1025 ( .A(n1307), .B(n1308), .ZN(n1121) );
XOR2_X1 U1026 ( .A(n1169), .B(n1309), .Z(n1308) );
XNOR2_X1 U1027 ( .A(n1310), .B(n1311), .ZN(n1169) );
XOR2_X1 U1028 ( .A(KEYINPUT36), .B(G107), .Z(n1311) );
XNOR2_X1 U1029 ( .A(G104), .B(G101), .ZN(n1310) );
XOR2_X1 U1030 ( .A(n1312), .B(n1313), .Z(n1307) );
XNOR2_X1 U1031 ( .A(G122), .B(n1314), .ZN(n1313) );
NAND2_X1 U1032 ( .A1(n1315), .A2(KEYINPUT55), .ZN(n1314) );
XNOR2_X1 U1033 ( .A(G110), .B(KEYINPUT30), .ZN(n1315) );
NAND2_X1 U1034 ( .A1(KEYINPUT5), .A2(n1316), .ZN(n1312) );
XOR2_X1 U1035 ( .A(n1317), .B(KEYINPUT16), .Z(n1306) );
NAND2_X1 U1036 ( .A1(G224), .A2(n1282), .ZN(n1317) );
INV_X1 U1037 ( .A(n1067), .ZN(n1226) );
NAND2_X1 U1038 ( .A1(n1032), .A2(n1041), .ZN(n1067) );
XOR2_X1 U1039 ( .A(n1318), .B(n1128), .Z(n1041) );
NAND2_X1 U1040 ( .A1(G217), .A2(n1296), .ZN(n1128) );
NAND2_X1 U1041 ( .A1(G234), .A2(n1319), .ZN(n1296) );
XNOR2_X1 U1042 ( .A(KEYINPUT52), .B(n1209), .ZN(n1319) );
NAND2_X1 U1043 ( .A1(n1130), .A2(n1209), .ZN(n1318) );
XNOR2_X1 U1044 ( .A(n1320), .B(n1321), .ZN(n1130) );
XOR2_X1 U1045 ( .A(G137), .B(n1322), .Z(n1321) );
XOR2_X1 U1046 ( .A(KEYINPUT26), .B(G146), .Z(n1322) );
XOR2_X1 U1047 ( .A(n1094), .B(n1323), .Z(n1320) );
XOR2_X1 U1048 ( .A(n1324), .B(n1325), .Z(n1323) );
NAND2_X1 U1049 ( .A1(G221), .A2(n1270), .ZN(n1325) );
AND2_X1 U1050 ( .A1(G234), .A2(n1282), .ZN(n1270) );
NAND2_X1 U1051 ( .A1(n1326), .A2(n1327), .ZN(n1324) );
OR2_X1 U1052 ( .A1(n1328), .A2(G110), .ZN(n1327) );
XOR2_X1 U1053 ( .A(n1329), .B(KEYINPUT4), .Z(n1326) );
NAND2_X1 U1054 ( .A1(G110), .A2(n1328), .ZN(n1329) );
XOR2_X1 U1055 ( .A(G119), .B(G128), .Z(n1328) );
XNOR2_X1 U1056 ( .A(G125), .B(G140), .ZN(n1094) );
INV_X1 U1057 ( .A(n1219), .ZN(n1032) );
XNOR2_X1 U1058 ( .A(n1330), .B(G472), .ZN(n1219) );
NAND2_X1 U1059 ( .A1(n1331), .A2(n1209), .ZN(n1330) );
INV_X1 U1060 ( .A(G902), .ZN(n1209) );
XOR2_X1 U1061 ( .A(n1153), .B(n1332), .Z(n1331) );
XOR2_X1 U1062 ( .A(G101), .B(n1333), .Z(n1332) );
NOR2_X1 U1063 ( .A1(KEYINPUT47), .A2(n1334), .ZN(n1333) );
XNOR2_X1 U1064 ( .A(n1295), .B(n1154), .ZN(n1334) );
XNOR2_X1 U1065 ( .A(n1335), .B(n1261), .ZN(n1154) );
XOR2_X1 U1066 ( .A(G128), .B(G143), .Z(n1261) );
XNOR2_X1 U1067 ( .A(G146), .B(KEYINPUT22), .ZN(n1335) );
NAND2_X1 U1068 ( .A1(n1336), .A2(n1337), .ZN(n1295) );
NAND2_X1 U1069 ( .A1(n1338), .A2(n1214), .ZN(n1337) );
INV_X1 U1070 ( .A(G134), .ZN(n1214) );
NAND2_X1 U1071 ( .A1(n1106), .A2(n1104), .ZN(n1338) );
OR2_X1 U1072 ( .A1(n1110), .A2(G137), .ZN(n1104) );
NAND2_X1 U1073 ( .A1(G137), .A2(n1110), .ZN(n1106) );
INV_X1 U1074 ( .A(G131), .ZN(n1110) );
NAND2_X1 U1075 ( .A1(n1339), .A2(G134), .ZN(n1336) );
XNOR2_X1 U1076 ( .A(G137), .B(G131), .ZN(n1339) );
XOR2_X1 U1077 ( .A(n1340), .B(n1309), .Z(n1153) );
XOR2_X1 U1078 ( .A(G113), .B(G119), .Z(n1309) );
XNOR2_X1 U1079 ( .A(n1341), .B(n1316), .ZN(n1340) );
INV_X1 U1080 ( .A(G116), .ZN(n1316) );
NAND2_X1 U1081 ( .A1(G210), .A2(n1256), .ZN(n1341) );
AND2_X1 U1082 ( .A1(n1282), .A2(n1300), .ZN(n1256) );
INV_X1 U1083 ( .A(G237), .ZN(n1300) );
XNOR2_X1 U1084 ( .A(G953), .B(KEYINPUT54), .ZN(n1282) );
endmodule


