//Key = 1111111110001110101100011000110000110000111010001100100101101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380;

XNOR2_X1 U758 ( .A(G107), .B(n1047), .ZN(G9) );
NAND2_X1 U759 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U760 ( .A1(n1050), .A2(n1051), .ZN(G75) );
NOR4_X1 U761 ( .A1(G953), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1051) );
NOR2_X1 U762 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U763 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR3_X1 U764 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
NOR2_X1 U765 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR3_X1 U767 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1062) );
NOR3_X1 U768 ( .A1(n1069), .A2(n1048), .A3(n1070), .ZN(n1068) );
AND2_X1 U769 ( .A1(n1065), .A2(n1069), .ZN(n1067) );
NOR3_X1 U770 ( .A1(n1071), .A2(n1072), .A3(n1065), .ZN(n1057) );
NOR2_X1 U771 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U772 ( .A1(n1075), .A2(n1059), .ZN(n1074) );
NOR2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR2_X1 U774 ( .A1(n1078), .A2(n1061), .ZN(n1073) );
NOR2_X1 U775 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U776 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NOR3_X1 U777 ( .A1(n1052), .A2(G953), .A3(G952), .ZN(n1050) );
AND4_X1 U778 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1052) );
NOR4_X1 U779 ( .A1(n1069), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1086) );
XOR2_X1 U780 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U781 ( .A1(n1092), .A2(KEYINPUT10), .ZN(n1091) );
XNOR2_X1 U782 ( .A(n1093), .B(n1094), .ZN(n1088) );
NAND2_X1 U783 ( .A1(KEYINPUT13), .A2(n1095), .ZN(n1093) );
NOR3_X1 U784 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1087) );
XNOR2_X1 U785 ( .A(G475), .B(KEYINPUT42), .ZN(n1098) );
NOR2_X1 U786 ( .A1(n1099), .A2(n1100), .ZN(n1085) );
XOR2_X1 U787 ( .A(n1101), .B(KEYINPUT3), .Z(n1099) );
XOR2_X1 U788 ( .A(n1102), .B(n1103), .Z(n1083) );
NOR2_X1 U789 ( .A1(KEYINPUT39), .A2(n1104), .ZN(n1103) );
XOR2_X1 U790 ( .A(n1105), .B(n1106), .Z(G72) );
NOR2_X1 U791 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U792 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
NAND2_X1 U793 ( .A1(n1111), .A2(n1112), .ZN(n1105) );
NAND2_X1 U794 ( .A1(n1113), .A2(n1108), .ZN(n1112) );
XNOR2_X1 U795 ( .A(n1114), .B(n1115), .ZN(n1113) );
NOR2_X1 U796 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U797 ( .A(KEYINPUT7), .B(n1118), .Z(n1117) );
NOR2_X1 U798 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND3_X1 U799 ( .A1(G900), .A2(n1114), .A3(G953), .ZN(n1111) );
XNOR2_X1 U800 ( .A(n1121), .B(n1122), .ZN(n1114) );
XNOR2_X1 U801 ( .A(KEYINPUT15), .B(n1123), .ZN(n1122) );
XNOR2_X1 U802 ( .A(n1124), .B(n1125), .ZN(n1121) );
NOR2_X1 U803 ( .A1(G140), .A2(n1126), .ZN(n1125) );
XOR2_X1 U804 ( .A(KEYINPUT63), .B(KEYINPUT0), .Z(n1126) );
XOR2_X1 U805 ( .A(n1127), .B(n1128), .Z(G69) );
XOR2_X1 U806 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U807 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U808 ( .A(KEYINPUT47), .B(n1133), .Z(n1132) );
XOR2_X1 U809 ( .A(n1134), .B(n1135), .Z(n1131) );
XNOR2_X1 U810 ( .A(G110), .B(G122), .ZN(n1135) );
NAND2_X1 U811 ( .A1(KEYINPUT23), .A2(n1136), .ZN(n1134) );
XOR2_X1 U812 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U813 ( .A1(n1139), .A2(n1140), .ZN(n1129) );
XNOR2_X1 U814 ( .A(KEYINPUT49), .B(n1108), .ZN(n1139) );
NAND2_X1 U815 ( .A1(G953), .A2(n1141), .ZN(n1127) );
NAND2_X1 U816 ( .A1(G224), .A2(G898), .ZN(n1141) );
NOR2_X1 U817 ( .A1(n1142), .A2(n1143), .ZN(G66) );
XOR2_X1 U818 ( .A(n1144), .B(n1145), .Z(n1143) );
NAND2_X1 U819 ( .A1(KEYINPUT6), .A2(n1146), .ZN(n1144) );
OR2_X1 U820 ( .A1(n1147), .A2(n1102), .ZN(n1146) );
NOR2_X1 U821 ( .A1(n1142), .A2(n1148), .ZN(G63) );
XNOR2_X1 U822 ( .A(n1149), .B(n1150), .ZN(n1148) );
XOR2_X1 U823 ( .A(KEYINPUT46), .B(n1151), .Z(n1150) );
NOR2_X1 U824 ( .A1(n1095), .A2(n1147), .ZN(n1151) );
NOR2_X1 U825 ( .A1(n1142), .A2(n1152), .ZN(G60) );
XOR2_X1 U826 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U827 ( .A1(KEYINPUT20), .A2(n1155), .ZN(n1154) );
XOR2_X1 U828 ( .A(KEYINPUT59), .B(n1096), .Z(n1155) );
NAND2_X1 U829 ( .A1(n1156), .A2(G475), .ZN(n1153) );
XOR2_X1 U830 ( .A(G104), .B(n1157), .Z(G6) );
NOR2_X1 U831 ( .A1(n1142), .A2(n1158), .ZN(G57) );
XNOR2_X1 U832 ( .A(n1159), .B(n1160), .ZN(n1158) );
XOR2_X1 U833 ( .A(n1161), .B(n1162), .Z(n1160) );
AND2_X1 U834 ( .A1(G472), .A2(n1156), .ZN(n1162) );
NAND2_X1 U835 ( .A1(n1163), .A2(n1164), .ZN(n1161) );
NOR2_X1 U836 ( .A1(n1142), .A2(n1165), .ZN(G54) );
XOR2_X1 U837 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U839 ( .A1(KEYINPUT26), .A2(n1170), .ZN(n1168) );
XOR2_X1 U840 ( .A(n1171), .B(n1172), .Z(n1166) );
AND2_X1 U841 ( .A1(G469), .A2(n1156), .ZN(n1172) );
NAND2_X1 U842 ( .A1(KEYINPUT62), .A2(n1173), .ZN(n1171) );
NOR3_X1 U843 ( .A1(n1142), .A2(n1174), .A3(n1175), .ZN(G51) );
NOR2_X1 U844 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
INV_X1 U845 ( .A(n1178), .ZN(n1177) );
NOR2_X1 U846 ( .A1(n1179), .A2(n1180), .ZN(n1176) );
NOR2_X1 U847 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NOR2_X1 U848 ( .A1(n1183), .A2(n1184), .ZN(n1179) );
NOR2_X1 U849 ( .A1(n1178), .A2(n1185), .ZN(n1174) );
NOR2_X1 U850 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NOR2_X1 U851 ( .A1(n1182), .A2(n1184), .ZN(n1187) );
XNOR2_X1 U852 ( .A(KEYINPUT56), .B(n1188), .ZN(n1184) );
INV_X1 U853 ( .A(n1183), .ZN(n1182) );
NOR2_X1 U854 ( .A1(n1183), .A2(n1181), .ZN(n1186) );
XOR2_X1 U855 ( .A(KEYINPUT30), .B(n1188), .Z(n1181) );
AND2_X1 U856 ( .A1(n1156), .A2(n1092), .ZN(n1188) );
INV_X1 U857 ( .A(n1147), .ZN(n1156) );
NAND2_X1 U858 ( .A1(G902), .A2(n1054), .ZN(n1147) );
OR4_X1 U859 ( .A1(n1140), .A2(n1116), .A3(n1120), .A4(n1189), .ZN(n1054) );
XNOR2_X1 U860 ( .A(KEYINPUT41), .B(n1119), .ZN(n1189) );
NAND3_X1 U861 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1120) );
NAND4_X1 U862 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1116) );
NAND3_X1 U863 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1195) );
OR2_X1 U864 ( .A1(n1200), .A2(KEYINPUT61), .ZN(n1198) );
NAND2_X1 U865 ( .A1(KEYINPUT61), .A2(n1201), .ZN(n1197) );
NAND3_X1 U866 ( .A1(n1202), .A2(n1080), .A3(n1203), .ZN(n1201) );
NAND2_X1 U867 ( .A1(n1204), .A2(n1077), .ZN(n1194) );
OR2_X1 U868 ( .A1(n1205), .A2(n1206), .ZN(n1193) );
NAND4_X1 U869 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1140) );
AND4_X1 U870 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1210) );
NOR2_X1 U871 ( .A1(n1157), .A2(n1215), .ZN(n1209) );
NOR2_X1 U872 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NOR2_X1 U873 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
NOR2_X1 U874 ( .A1(n1065), .A2(n1220), .ZN(n1219) );
XOR2_X1 U875 ( .A(KEYINPUT52), .B(n1077), .Z(n1220) );
NOR3_X1 U876 ( .A1(n1221), .A2(n1061), .A3(n1222), .ZN(n1218) );
AND2_X1 U877 ( .A1(n1070), .A2(n1049), .ZN(n1157) );
NOR2_X1 U878 ( .A1(n1061), .A2(n1217), .ZN(n1049) );
INV_X1 U879 ( .A(n1223), .ZN(n1061) );
NAND4_X1 U880 ( .A1(n1048), .A2(n1223), .A3(n1224), .A4(n1064), .ZN(n1208) );
AND3_X1 U881 ( .A1(n1080), .A2(n1221), .A3(n1225), .ZN(n1224) );
INV_X1 U882 ( .A(KEYINPUT55), .ZN(n1221) );
INV_X1 U883 ( .A(n1226), .ZN(n1080) );
NAND2_X1 U884 ( .A1(n1227), .A2(n1228), .ZN(n1207) );
XNOR2_X1 U885 ( .A(KEYINPUT25), .B(n1229), .ZN(n1227) );
XNOR2_X1 U886 ( .A(n1230), .B(n1231), .ZN(n1183) );
NAND2_X1 U887 ( .A1(n1232), .A2(KEYINPUT5), .ZN(n1230) );
XNOR2_X1 U888 ( .A(n1233), .B(n1170), .ZN(n1232) );
NAND2_X1 U889 ( .A1(KEYINPUT16), .A2(n1123), .ZN(n1233) );
NOR2_X1 U890 ( .A1(n1108), .A2(G952), .ZN(n1142) );
XNOR2_X1 U891 ( .A(n1234), .B(n1235), .ZN(G48) );
NOR2_X1 U892 ( .A1(n1206), .A2(n1205), .ZN(n1235) );
INV_X1 U893 ( .A(n1070), .ZN(n1206) );
NAND2_X1 U894 ( .A1(n1236), .A2(n1237), .ZN(G45) );
OR2_X1 U895 ( .A1(n1238), .A2(G143), .ZN(n1237) );
NAND2_X1 U896 ( .A1(G143), .A2(n1239), .ZN(n1236) );
NAND2_X1 U897 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
OR2_X1 U898 ( .A1(n1196), .A2(KEYINPUT48), .ZN(n1241) );
NAND2_X1 U899 ( .A1(KEYINPUT48), .A2(n1238), .ZN(n1240) );
OR2_X1 U900 ( .A1(KEYINPUT37), .A2(n1196), .ZN(n1238) );
NAND3_X1 U901 ( .A1(n1076), .A2(n1242), .A3(n1243), .ZN(n1196) );
NOR3_X1 U902 ( .A1(n1203), .A2(n1244), .A3(n1245), .ZN(n1243) );
XNOR2_X1 U903 ( .A(G140), .B(n1246), .ZN(G42) );
NOR2_X1 U904 ( .A1(KEYINPUT43), .A2(n1247), .ZN(n1246) );
NOR2_X1 U905 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
XOR2_X1 U906 ( .A(KEYINPUT8), .B(n1077), .Z(n1249) );
XOR2_X1 U907 ( .A(n1250), .B(n1251), .Z(G39) );
XNOR2_X1 U908 ( .A(KEYINPUT27), .B(n1252), .ZN(n1251) );
AND2_X1 U909 ( .A1(n1199), .A2(n1200), .ZN(n1250) );
XNOR2_X1 U910 ( .A(G134), .B(n1190), .ZN(G36) );
NAND3_X1 U911 ( .A1(n1076), .A2(n1048), .A3(n1200), .ZN(n1190) );
XNOR2_X1 U912 ( .A(G131), .B(n1192), .ZN(G33) );
NAND2_X1 U913 ( .A1(n1204), .A2(n1076), .ZN(n1192) );
INV_X1 U914 ( .A(n1248), .ZN(n1204) );
NAND2_X1 U915 ( .A1(n1200), .A2(n1070), .ZN(n1248) );
NOR3_X1 U916 ( .A1(n1226), .A2(n1203), .A3(n1071), .ZN(n1200) );
INV_X1 U917 ( .A(n1202), .ZN(n1071) );
NOR2_X1 U918 ( .A1(n1066), .A2(n1069), .ZN(n1202) );
INV_X1 U919 ( .A(n1253), .ZN(n1069) );
XNOR2_X1 U920 ( .A(n1254), .B(n1255), .ZN(G30) );
NAND2_X1 U921 ( .A1(n1256), .A2(n1257), .ZN(n1254) );
OR3_X1 U922 ( .A1(n1205), .A2(n1048), .A3(KEYINPUT2), .ZN(n1257) );
NAND2_X1 U923 ( .A1(n1119), .A2(KEYINPUT2), .ZN(n1256) );
NOR2_X1 U924 ( .A1(n1205), .A2(n1222), .ZN(n1119) );
INV_X1 U925 ( .A(n1048), .ZN(n1222) );
NAND4_X1 U926 ( .A1(n1258), .A2(n1242), .A3(n1100), .A4(n1259), .ZN(n1205) );
NAND2_X1 U927 ( .A1(n1260), .A2(n1261), .ZN(G3) );
NAND2_X1 U928 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XOR2_X1 U929 ( .A(KEYINPUT60), .B(n1264), .Z(n1260) );
NOR2_X1 U930 ( .A1(n1262), .A2(n1263), .ZN(n1264) );
INV_X1 U931 ( .A(G101), .ZN(n1263) );
INV_X1 U932 ( .A(n1214), .ZN(n1262) );
NAND2_X1 U933 ( .A1(n1265), .A2(n1076), .ZN(n1214) );
NAND2_X1 U934 ( .A1(n1266), .A2(n1267), .ZN(G27) );
NAND2_X1 U935 ( .A1(G125), .A2(n1191), .ZN(n1267) );
XOR2_X1 U936 ( .A(n1268), .B(KEYINPUT33), .Z(n1266) );
OR2_X1 U937 ( .A1(n1191), .A2(G125), .ZN(n1268) );
NAND3_X1 U938 ( .A1(n1077), .A2(n1070), .A3(n1269), .ZN(n1191) );
NOR3_X1 U939 ( .A1(n1059), .A2(n1203), .A3(n1064), .ZN(n1269) );
INV_X1 U940 ( .A(n1259), .ZN(n1203) );
NAND2_X1 U941 ( .A1(n1056), .A2(n1270), .ZN(n1259) );
NAND4_X1 U942 ( .A1(G953), .A2(G902), .A3(n1271), .A4(n1110), .ZN(n1270) );
INV_X1 U943 ( .A(G900), .ZN(n1110) );
INV_X1 U944 ( .A(n1084), .ZN(n1059) );
XNOR2_X1 U945 ( .A(G122), .B(n1213), .ZN(G24) );
NAND4_X1 U946 ( .A1(n1272), .A2(n1223), .A3(n1273), .A4(n1274), .ZN(n1213) );
NOR2_X1 U947 ( .A1(n1100), .A2(n1258), .ZN(n1223) );
XNOR2_X1 U948 ( .A(n1275), .B(n1276), .ZN(G21) );
NAND2_X1 U949 ( .A1(KEYINPUT34), .A2(n1212), .ZN(n1275) );
NAND2_X1 U950 ( .A1(n1199), .A2(n1272), .ZN(n1212) );
NOR3_X1 U951 ( .A1(n1277), .A2(n1278), .A3(n1065), .ZN(n1199) );
XNOR2_X1 U952 ( .A(G116), .B(n1211), .ZN(G18) );
NAND3_X1 U953 ( .A1(n1272), .A2(n1048), .A3(n1076), .ZN(n1211) );
NOR2_X1 U954 ( .A1(n1273), .A2(n1244), .ZN(n1048) );
AND3_X1 U955 ( .A1(n1228), .A2(n1225), .A3(n1084), .ZN(n1272) );
INV_X1 U956 ( .A(n1064), .ZN(n1228) );
XOR2_X1 U957 ( .A(G113), .B(n1279), .Z(G15) );
NOR2_X1 U958 ( .A1(n1064), .A2(n1229), .ZN(n1279) );
NAND4_X1 U959 ( .A1(n1070), .A2(n1076), .A3(n1084), .A4(n1225), .ZN(n1229) );
NOR2_X1 U960 ( .A1(n1081), .A2(n1280), .ZN(n1084) );
INV_X1 U961 ( .A(n1082), .ZN(n1280) );
NOR2_X1 U962 ( .A1(n1278), .A2(n1258), .ZN(n1076) );
INV_X1 U963 ( .A(n1277), .ZN(n1258) );
INV_X1 U964 ( .A(n1100), .ZN(n1278) );
NOR2_X1 U965 ( .A1(n1274), .A2(n1245), .ZN(n1070) );
XNOR2_X1 U966 ( .A(G110), .B(n1281), .ZN(G12) );
NAND2_X1 U967 ( .A1(n1077), .A2(n1265), .ZN(n1281) );
NOR2_X1 U968 ( .A1(n1065), .A2(n1217), .ZN(n1265) );
NAND2_X1 U969 ( .A1(n1242), .A2(n1225), .ZN(n1217) );
NAND2_X1 U970 ( .A1(n1056), .A2(n1282), .ZN(n1225) );
NAND3_X1 U971 ( .A1(G902), .A2(n1271), .A3(n1133), .ZN(n1282) );
AND2_X1 U972 ( .A1(G953), .A2(n1283), .ZN(n1133) );
XOR2_X1 U973 ( .A(KEYINPUT18), .B(G898), .Z(n1283) );
NAND3_X1 U974 ( .A1(n1271), .A2(n1108), .A3(G952), .ZN(n1056) );
NAND2_X1 U975 ( .A1(G237), .A2(G234), .ZN(n1271) );
NOR2_X1 U976 ( .A1(n1064), .A2(n1226), .ZN(n1242) );
NAND2_X1 U977 ( .A1(n1081), .A2(n1082), .ZN(n1226) );
NAND2_X1 U978 ( .A1(G221), .A2(n1284), .ZN(n1082) );
XOR2_X1 U979 ( .A(n1285), .B(n1286), .Z(n1081) );
XOR2_X1 U980 ( .A(KEYINPUT24), .B(G469), .Z(n1286) );
NAND2_X1 U981 ( .A1(n1287), .A2(n1288), .ZN(n1285) );
XNOR2_X1 U982 ( .A(n1169), .B(n1124), .ZN(n1287) );
XNOR2_X1 U983 ( .A(n1289), .B(n1290), .ZN(n1169) );
XNOR2_X1 U984 ( .A(n1291), .B(n1292), .ZN(n1290) );
NOR2_X1 U985 ( .A1(G953), .A2(n1109), .ZN(n1292) );
INV_X1 U986 ( .A(G227), .ZN(n1109) );
NAND2_X1 U987 ( .A1(n1066), .A2(n1253), .ZN(n1064) );
NAND2_X1 U988 ( .A1(G214), .A2(n1293), .ZN(n1253) );
XOR2_X1 U989 ( .A(n1090), .B(n1294), .Z(n1066) );
XOR2_X1 U990 ( .A(KEYINPUT29), .B(n1092), .Z(n1294) );
AND2_X1 U991 ( .A1(G210), .A2(n1293), .ZN(n1092) );
NAND2_X1 U992 ( .A1(n1295), .A2(n1288), .ZN(n1293) );
INV_X1 U993 ( .A(G237), .ZN(n1295) );
NAND2_X1 U994 ( .A1(n1296), .A2(n1288), .ZN(n1090) );
XOR2_X1 U995 ( .A(n1297), .B(n1298), .Z(n1296) );
XNOR2_X1 U996 ( .A(n1178), .B(n1299), .ZN(n1298) );
XNOR2_X1 U997 ( .A(n1300), .B(n1138), .ZN(n1178) );
XNOR2_X1 U998 ( .A(n1301), .B(G113), .ZN(n1138) );
NAND2_X1 U999 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
OR2_X1 U1000 ( .A1(n1276), .A2(G116), .ZN(n1303) );
XOR2_X1 U1001 ( .A(n1304), .B(KEYINPUT9), .Z(n1302) );
NAND2_X1 U1002 ( .A1(G116), .A2(n1276), .ZN(n1304) );
XNOR2_X1 U1003 ( .A(n1289), .B(n1305), .ZN(n1300) );
XNOR2_X1 U1004 ( .A(G110), .B(n1137), .ZN(n1289) );
XNOR2_X1 U1005 ( .A(n1306), .B(n1307), .ZN(n1137) );
XNOR2_X1 U1006 ( .A(G104), .B(G107), .ZN(n1306) );
XNOR2_X1 U1007 ( .A(G125), .B(n1308), .ZN(n1297) );
NOR2_X1 U1008 ( .A1(KEYINPUT17), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1009 ( .A(KEYINPUT28), .B(n1231), .Z(n1309) );
AND2_X1 U1010 ( .A1(G224), .A2(n1108), .ZN(n1231) );
NAND2_X1 U1011 ( .A1(n1244), .A2(n1245), .ZN(n1065) );
INV_X1 U1012 ( .A(n1273), .ZN(n1245) );
NAND2_X1 U1013 ( .A1(n1310), .A2(n1101), .ZN(n1273) );
NAND2_X1 U1014 ( .A1(G475), .A2(n1311), .ZN(n1101) );
OR2_X1 U1015 ( .A1(n1096), .A2(n1097), .ZN(n1311) );
XOR2_X1 U1016 ( .A(KEYINPUT44), .B(n1312), .Z(n1310) );
NOR3_X1 U1017 ( .A1(n1096), .A2(G475), .A3(n1097), .ZN(n1312) );
XOR2_X1 U1018 ( .A(n1288), .B(KEYINPUT14), .Z(n1097) );
XNOR2_X1 U1019 ( .A(n1313), .B(n1314), .ZN(n1096) );
XOR2_X1 U1020 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1021 ( .A(n1317), .B(n1318), .Z(n1316) );
NAND2_X1 U1022 ( .A1(G214), .A2(n1319), .ZN(n1318) );
NAND4_X1 U1023 ( .A1(KEYINPUT19), .A2(n1320), .A3(n1321), .A4(n1322), .ZN(n1317) );
NAND3_X1 U1024 ( .A1(n1323), .A2(n1324), .A3(G146), .ZN(n1322) );
NAND2_X1 U1025 ( .A1(n1325), .A2(n1234), .ZN(n1321) );
NAND2_X1 U1026 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
NAND2_X1 U1027 ( .A1(G140), .A2(n1123), .ZN(n1327) );
XNOR2_X1 U1028 ( .A(n1328), .B(n1324), .ZN(n1326) );
NAND2_X1 U1029 ( .A1(G125), .A2(n1291), .ZN(n1328) );
OR2_X1 U1030 ( .A1(n1329), .A2(n1324), .ZN(n1320) );
INV_X1 U1031 ( .A(KEYINPUT45), .ZN(n1324) );
NOR2_X1 U1032 ( .A1(G143), .A2(KEYINPUT22), .ZN(n1315) );
XOR2_X1 U1033 ( .A(n1330), .B(n1331), .Z(n1313) );
XOR2_X1 U1034 ( .A(G104), .B(n1332), .Z(n1331) );
NOR2_X1 U1035 ( .A1(G113), .A2(KEYINPUT31), .ZN(n1332) );
XNOR2_X1 U1036 ( .A(G131), .B(G122), .ZN(n1330) );
INV_X1 U1037 ( .A(n1274), .ZN(n1244) );
NAND2_X1 U1038 ( .A1(n1333), .A2(n1334), .ZN(n1274) );
OR2_X1 U1039 ( .A1(n1094), .A2(G478), .ZN(n1334) );
XOR2_X1 U1040 ( .A(n1335), .B(KEYINPUT36), .Z(n1333) );
NAND2_X1 U1041 ( .A1(n1336), .A2(n1094), .ZN(n1335) );
NAND2_X1 U1042 ( .A1(n1149), .A2(n1288), .ZN(n1094) );
XNOR2_X1 U1043 ( .A(n1337), .B(n1338), .ZN(n1149) );
XNOR2_X1 U1044 ( .A(G134), .B(n1339), .ZN(n1338) );
NAND2_X1 U1045 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
XNOR2_X1 U1046 ( .A(KEYINPUT57), .B(KEYINPUT40), .ZN(n1340) );
XOR2_X1 U1047 ( .A(n1342), .B(n1343), .Z(n1337) );
AND3_X1 U1048 ( .A1(G234), .A2(n1108), .A3(G217), .ZN(n1343) );
NAND2_X1 U1049 ( .A1(n1344), .A2(n1345), .ZN(n1342) );
NAND2_X1 U1050 ( .A1(G107), .A2(n1346), .ZN(n1345) );
XOR2_X1 U1051 ( .A(KEYINPUT12), .B(n1347), .Z(n1344) );
NOR2_X1 U1052 ( .A1(G107), .A2(n1346), .ZN(n1347) );
XNOR2_X1 U1053 ( .A(n1305), .B(G116), .ZN(n1346) );
INV_X1 U1054 ( .A(G122), .ZN(n1305) );
XNOR2_X1 U1055 ( .A(KEYINPUT51), .B(n1095), .ZN(n1336) );
INV_X1 U1056 ( .A(G478), .ZN(n1095) );
NOR2_X1 U1057 ( .A1(n1277), .A2(n1100), .ZN(n1077) );
XNOR2_X1 U1058 ( .A(n1348), .B(n1349), .ZN(n1100) );
XOR2_X1 U1059 ( .A(KEYINPUT11), .B(G472), .Z(n1349) );
NAND2_X1 U1060 ( .A1(n1350), .A2(n1288), .ZN(n1348) );
XOR2_X1 U1061 ( .A(n1351), .B(n1352), .Z(n1350) );
NOR2_X1 U1062 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
XOR2_X1 U1063 ( .A(n1163), .B(KEYINPUT35), .Z(n1354) );
NAND2_X1 U1064 ( .A1(n1307), .A2(n1355), .ZN(n1163) );
NAND2_X1 U1065 ( .A1(G210), .A2(n1319), .ZN(n1355) );
INV_X1 U1066 ( .A(n1164), .ZN(n1353) );
NAND3_X1 U1067 ( .A1(n1356), .A2(n1319), .A3(G210), .ZN(n1164) );
AND2_X1 U1068 ( .A1(n1357), .A2(n1108), .ZN(n1319) );
XNOR2_X1 U1069 ( .A(G237), .B(KEYINPUT54), .ZN(n1357) );
INV_X1 U1070 ( .A(n1307), .ZN(n1356) );
XOR2_X1 U1071 ( .A(G101), .B(KEYINPUT1), .Z(n1307) );
NOR2_X1 U1072 ( .A1(KEYINPUT38), .A2(n1358), .ZN(n1351) );
XNOR2_X1 U1073 ( .A(KEYINPUT53), .B(n1359), .ZN(n1358) );
INV_X1 U1074 ( .A(n1159), .ZN(n1359) );
XNOR2_X1 U1075 ( .A(n1360), .B(n1361), .ZN(n1159) );
XOR2_X1 U1076 ( .A(G116), .B(G113), .Z(n1361) );
XNOR2_X1 U1077 ( .A(n1124), .B(n1362), .ZN(n1360) );
NOR2_X1 U1078 ( .A1(G119), .A2(KEYINPUT32), .ZN(n1362) );
XOR2_X1 U1079 ( .A(n1173), .B(n1170), .Z(n1124) );
INV_X1 U1080 ( .A(n1299), .ZN(n1170) );
XOR2_X1 U1081 ( .A(G146), .B(n1341), .Z(n1299) );
XNOR2_X1 U1082 ( .A(n1255), .B(G143), .ZN(n1341) );
INV_X1 U1083 ( .A(G128), .ZN(n1255) );
XNOR2_X1 U1084 ( .A(G131), .B(n1363), .ZN(n1173) );
XNOR2_X1 U1085 ( .A(n1252), .B(G134), .ZN(n1363) );
XOR2_X1 U1086 ( .A(n1364), .B(n1104), .Z(n1277) );
OR2_X1 U1087 ( .A1(n1145), .A2(G902), .ZN(n1104) );
XNOR2_X1 U1088 ( .A(n1365), .B(n1366), .ZN(n1145) );
NOR2_X1 U1089 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
XOR2_X1 U1090 ( .A(KEYINPUT50), .B(n1369), .Z(n1368) );
NOR2_X1 U1091 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
AND2_X1 U1092 ( .A1(n1371), .A2(n1370), .ZN(n1367) );
XOR2_X1 U1093 ( .A(n1372), .B(n1373), .Z(n1370) );
XNOR2_X1 U1094 ( .A(n1276), .B(G110), .ZN(n1373) );
INV_X1 U1095 ( .A(G119), .ZN(n1276) );
XNOR2_X1 U1096 ( .A(G128), .B(KEYINPUT58), .ZN(n1372) );
NAND3_X1 U1097 ( .A1(n1374), .A2(n1375), .A3(n1329), .ZN(n1371) );
NAND3_X1 U1098 ( .A1(G125), .A2(n1291), .A3(G146), .ZN(n1329) );
INV_X1 U1099 ( .A(G140), .ZN(n1291) );
NAND2_X1 U1100 ( .A1(n1323), .A2(n1234), .ZN(n1375) );
INV_X1 U1101 ( .A(G146), .ZN(n1234) );
XNOR2_X1 U1102 ( .A(G140), .B(G125), .ZN(n1323) );
NAND3_X1 U1103 ( .A1(G140), .A2(n1123), .A3(G146), .ZN(n1374) );
INV_X1 U1104 ( .A(G125), .ZN(n1123) );
NAND2_X1 U1105 ( .A1(n1376), .A2(n1377), .ZN(n1365) );
NAND2_X1 U1106 ( .A1(n1378), .A2(n1252), .ZN(n1377) );
NAND2_X1 U1107 ( .A1(n1379), .A2(n1380), .ZN(n1376) );
INV_X1 U1108 ( .A(n1378), .ZN(n1380) );
NAND3_X1 U1109 ( .A1(G234), .A2(n1108), .A3(G221), .ZN(n1378) );
INV_X1 U1110 ( .A(G953), .ZN(n1108) );
XNOR2_X1 U1111 ( .A(KEYINPUT21), .B(n1252), .ZN(n1379) );
INV_X1 U1112 ( .A(G137), .ZN(n1252) );
NAND2_X1 U1113 ( .A1(KEYINPUT4), .A2(n1102), .ZN(n1364) );
NAND2_X1 U1114 ( .A1(G217), .A2(n1284), .ZN(n1102) );
NAND2_X1 U1115 ( .A1(G234), .A2(n1288), .ZN(n1284) );
INV_X1 U1116 ( .A(G902), .ZN(n1288) );
endmodule


