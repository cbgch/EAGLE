//Key = 1101000110100001110110100001010000100001110011001111100111100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399;

XNOR2_X1 U770 ( .A(G107), .B(n1058), .ZN(G9) );
NOR2_X1 U771 ( .A1(n1059), .A2(n1060), .ZN(G75) );
NOR4_X1 U772 ( .A1(n1061), .A2(n1062), .A3(G953), .A4(n1063), .ZN(n1060) );
NOR3_X1 U773 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1062) );
NOR4_X1 U774 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1065) );
NAND3_X1 U775 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1061) );
NAND2_X1 U776 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NAND2_X1 U777 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND4_X1 U778 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1077) );
NAND2_X1 U779 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U780 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U781 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
OR2_X1 U782 ( .A1(n1088), .A2(KEYINPUT17), .ZN(n1087) );
NAND3_X1 U783 ( .A1(n1089), .A2(n1090), .A3(n1088), .ZN(n1082) );
NAND2_X1 U784 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U785 ( .A1(KEYINPUT17), .A2(n1084), .ZN(n1092) );
INV_X1 U786 ( .A(n1093), .ZN(n1091) );
NAND3_X1 U787 ( .A1(n1094), .A2(n1095), .A3(n1093), .ZN(n1089) );
NAND2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NAND3_X1 U789 ( .A1(n1084), .A2(n1098), .A3(n1099), .ZN(n1076) );
NAND2_X1 U790 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NAND3_X1 U791 ( .A1(n1080), .A2(n1102), .A3(n1079), .ZN(n1101) );
NAND2_X1 U792 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND2_X1 U793 ( .A1(n1078), .A2(n1105), .ZN(n1100) );
NAND2_X1 U794 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U795 ( .A1(n1108), .A2(n1064), .ZN(n1107) );
INV_X1 U796 ( .A(KEYINPUT5), .ZN(n1064) );
NAND2_X1 U797 ( .A1(n1080), .A2(n1109), .ZN(n1106) );
INV_X1 U798 ( .A(n1070), .ZN(n1074) );
XOR2_X1 U799 ( .A(KEYINPUT6), .B(n1110), .Z(n1071) );
NOR3_X1 U800 ( .A1(n1063), .A2(G953), .A3(G952), .ZN(n1059) );
AND4_X1 U801 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1063) );
NOR4_X1 U802 ( .A1(n1115), .A2(n1116), .A3(n1067), .A4(n1066), .ZN(n1114) );
AND2_X1 U803 ( .A1(KEYINPUT8), .A2(n1117), .ZN(n1116) );
NOR2_X1 U804 ( .A1(KEYINPUT8), .A2(n1118), .ZN(n1115) );
NOR2_X1 U805 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XOR2_X1 U806 ( .A(KEYINPUT39), .B(n1121), .Z(n1112) );
XOR2_X1 U807 ( .A(KEYINPUT9), .B(n1122), .Z(n1111) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
INV_X1 U809 ( .A(n1125), .ZN(n1123) );
XOR2_X1 U810 ( .A(n1126), .B(n1127), .Z(G72) );
XOR2_X1 U811 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U812 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U813 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U814 ( .A1(KEYINPUT34), .A2(n1134), .ZN(n1133) );
NAND3_X1 U815 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1132) );
NAND2_X1 U816 ( .A1(KEYINPUT53), .A2(n1138), .ZN(n1137) );
NAND3_X1 U817 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1136) );
INV_X1 U818 ( .A(KEYINPUT53), .ZN(n1140) );
OR2_X1 U819 ( .A1(n1141), .A2(n1139), .ZN(n1135) );
NOR2_X1 U820 ( .A1(KEYINPUT47), .A2(n1138), .ZN(n1139) );
NAND2_X1 U821 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U822 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U823 ( .A(KEYINPUT49), .B(n1146), .Z(n1144) );
XOR2_X1 U824 ( .A(n1147), .B(KEYINPUT4), .Z(n1142) );
NAND2_X1 U825 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XNOR2_X1 U826 ( .A(KEYINPUT49), .B(n1146), .ZN(n1149) );
XOR2_X1 U827 ( .A(n1145), .B(KEYINPUT45), .Z(n1148) );
NOR2_X1 U828 ( .A1(n1150), .A2(n1151), .ZN(n1128) );
NOR2_X1 U829 ( .A1(n1152), .A2(n1153), .ZN(n1150) );
INV_X1 U830 ( .A(G900), .ZN(n1153) );
XNOR2_X1 U831 ( .A(G227), .B(KEYINPUT43), .ZN(n1152) );
NOR2_X1 U832 ( .A1(n1073), .A2(G953), .ZN(n1126) );
XOR2_X1 U833 ( .A(n1154), .B(n1155), .Z(G69) );
XOR2_X1 U834 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND3_X1 U835 ( .A1(n1158), .A2(n1159), .A3(n1151), .ZN(n1157) );
OR3_X1 U836 ( .A1(n1160), .A2(n1161), .A3(KEYINPUT1), .ZN(n1159) );
NAND2_X1 U837 ( .A1(KEYINPUT1), .A2(n1110), .ZN(n1158) );
NAND4_X1 U838 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1156) );
OR2_X1 U839 ( .A1(n1166), .A2(KEYINPUT26), .ZN(n1165) );
NAND2_X1 U840 ( .A1(n1167), .A2(KEYINPUT26), .ZN(n1164) );
XOR2_X1 U841 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U842 ( .A1(n1170), .A2(n1151), .ZN(n1154) );
AND2_X1 U843 ( .A1(G224), .A2(G898), .ZN(n1170) );
NOR3_X1 U844 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(G66) );
AND2_X1 U845 ( .A1(KEYINPUT16), .A2(n1174), .ZN(n1173) );
NOR3_X1 U846 ( .A1(KEYINPUT16), .A2(G953), .A3(G952), .ZN(n1172) );
XNOR2_X1 U847 ( .A(n1175), .B(n1176), .ZN(n1171) );
NOR2_X1 U848 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR2_X1 U849 ( .A1(n1174), .A2(n1179), .ZN(G63) );
XOR2_X1 U850 ( .A(n1180), .B(n1181), .Z(n1179) );
NAND3_X1 U851 ( .A1(G478), .A2(n1182), .A3(n1183), .ZN(n1180) );
XOR2_X1 U852 ( .A(n1184), .B(KEYINPUT27), .Z(n1183) );
NOR2_X1 U853 ( .A1(n1174), .A2(n1185), .ZN(G60) );
XNOR2_X1 U854 ( .A(n1186), .B(n1187), .ZN(n1185) );
NOR2_X1 U855 ( .A1(n1188), .A2(n1178), .ZN(n1187) );
INV_X1 U856 ( .A(G475), .ZN(n1188) );
XOR2_X1 U857 ( .A(n1189), .B(n1190), .Z(G6) );
NOR2_X1 U858 ( .A1(n1174), .A2(n1191), .ZN(G57) );
XOR2_X1 U859 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U860 ( .A(n1194), .B(n1195), .Z(n1193) );
NOR2_X1 U861 ( .A1(n1120), .A2(n1178), .ZN(n1195) );
INV_X1 U862 ( .A(G472), .ZN(n1120) );
NAND2_X1 U863 ( .A1(n1196), .A2(KEYINPUT51), .ZN(n1194) );
XOR2_X1 U864 ( .A(n1197), .B(n1198), .Z(n1196) );
NAND3_X1 U865 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1197) );
OR2_X1 U866 ( .A1(n1202), .A2(KEYINPUT48), .ZN(n1201) );
NAND3_X1 U867 ( .A1(KEYINPUT48), .A2(n1202), .A3(n1203), .ZN(n1200) );
NAND2_X1 U868 ( .A1(n1204), .A2(n1205), .ZN(n1199) );
NAND2_X1 U869 ( .A1(KEYINPUT48), .A2(n1206), .ZN(n1205) );
XNOR2_X1 U870 ( .A(KEYINPUT56), .B(n1202), .ZN(n1206) );
XOR2_X1 U871 ( .A(n1207), .B(G101), .Z(n1192) );
NOR2_X1 U872 ( .A1(n1174), .A2(n1208), .ZN(G54) );
XOR2_X1 U873 ( .A(n1209), .B(n1210), .Z(n1208) );
XOR2_X1 U874 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U875 ( .A(n1213), .B(n1214), .Z(n1212) );
XOR2_X1 U876 ( .A(n1215), .B(n1216), .Z(n1209) );
XNOR2_X1 U877 ( .A(n1217), .B(n1218), .ZN(n1216) );
NOR2_X1 U878 ( .A1(KEYINPUT60), .A2(n1203), .ZN(n1218) );
NAND2_X1 U879 ( .A1(KEYINPUT22), .A2(G110), .ZN(n1217) );
XNOR2_X1 U880 ( .A(n1219), .B(n1220), .ZN(n1215) );
NOR2_X1 U881 ( .A1(n1221), .A2(n1178), .ZN(n1220) );
INV_X1 U882 ( .A(G469), .ZN(n1221) );
NOR2_X1 U883 ( .A1(n1174), .A2(n1222), .ZN(G51) );
XOR2_X1 U884 ( .A(n1223), .B(n1224), .Z(n1222) );
NOR2_X1 U885 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U886 ( .A(KEYINPUT11), .B(n1227), .Z(n1226) );
AND2_X1 U887 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NOR2_X1 U888 ( .A1(n1230), .A2(n1178), .ZN(n1223) );
NAND2_X1 U889 ( .A1(G902), .A2(n1182), .ZN(n1178) );
NAND2_X1 U890 ( .A1(n1073), .A2(n1110), .ZN(n1182) );
NOR2_X1 U891 ( .A1(n1161), .A2(n1231), .ZN(n1110) );
INV_X1 U892 ( .A(n1160), .ZN(n1231) );
NAND2_X1 U893 ( .A1(n1232), .A2(n1233), .ZN(n1160) );
NAND4_X1 U894 ( .A1(n1190), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1161) );
AND3_X1 U895 ( .A1(n1237), .A2(n1058), .A3(n1238), .ZN(n1236) );
NAND3_X1 U896 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(n1058) );
NAND2_X1 U897 ( .A1(n1242), .A2(n1243), .ZN(n1235) );
NAND2_X1 U898 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XNOR2_X1 U899 ( .A(KEYINPUT41), .B(n1246), .ZN(n1245) );
XOR2_X1 U900 ( .A(n1247), .B(KEYINPUT31), .Z(n1244) );
NAND3_X1 U901 ( .A1(n1239), .A2(n1240), .A3(n1233), .ZN(n1190) );
AND4_X1 U902 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1073) );
AND4_X1 U903 ( .A1(n1252), .A2(n1253), .A3(n1254), .A4(n1255), .ZN(n1251) );
NOR4_X1 U904 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1250) );
AND2_X1 U905 ( .A1(KEYINPUT10), .A2(n1260), .ZN(n1259) );
NOR3_X1 U906 ( .A1(KEYINPUT10), .A2(n1084), .A3(n1261), .ZN(n1258) );
NOR4_X1 U907 ( .A1(n1262), .A2(n1263), .A3(n1104), .A4(n1264), .ZN(n1257) );
INV_X1 U908 ( .A(KEYINPUT14), .ZN(n1262) );
NOR2_X1 U909 ( .A1(KEYINPUT14), .A2(n1265), .ZN(n1256) );
NOR2_X1 U910 ( .A1(n1151), .A2(G952), .ZN(n1174) );
XOR2_X1 U911 ( .A(n1266), .B(n1254), .Z(G48) );
NAND3_X1 U912 ( .A1(n1267), .A2(n1263), .A3(n1233), .ZN(n1254) );
NAND2_X1 U913 ( .A1(n1268), .A2(n1269), .ZN(G45) );
NAND2_X1 U914 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U915 ( .A1(G143), .A2(n1272), .ZN(n1268) );
NAND2_X1 U916 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U917 ( .A1(KEYINPUT32), .A2(n1275), .ZN(n1274) );
INV_X1 U918 ( .A(n1248), .ZN(n1275) );
OR2_X1 U919 ( .A1(n1270), .A2(KEYINPUT32), .ZN(n1273) );
NOR2_X1 U920 ( .A1(KEYINPUT35), .A2(n1248), .ZN(n1270) );
NAND3_X1 U921 ( .A1(n1108), .A2(n1239), .A3(n1276), .ZN(n1248) );
AND3_X1 U922 ( .A1(n1277), .A2(n1263), .A3(n1121), .ZN(n1276) );
XNOR2_X1 U923 ( .A(G140), .B(n1249), .ZN(G42) );
NAND4_X1 U924 ( .A1(n1233), .A2(n1278), .A3(n1080), .A4(n1109), .ZN(n1249) );
XNOR2_X1 U925 ( .A(G137), .B(n1253), .ZN(G39) );
NAND4_X1 U926 ( .A1(n1078), .A2(n1278), .A3(n1279), .A4(n1109), .ZN(n1253) );
XNOR2_X1 U927 ( .A(G134), .B(n1252), .ZN(G36) );
NAND3_X1 U928 ( .A1(n1108), .A2(n1241), .A3(n1278), .ZN(n1252) );
NAND3_X1 U929 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(G33) );
NAND2_X1 U930 ( .A1(G131), .A2(n1255), .ZN(n1282) );
NAND2_X1 U931 ( .A1(n1283), .A2(n1284), .ZN(n1281) );
INV_X1 U932 ( .A(KEYINPUT15), .ZN(n1284) );
NAND2_X1 U933 ( .A1(n1285), .A2(n1145), .ZN(n1283) );
XNOR2_X1 U934 ( .A(KEYINPUT63), .B(n1255), .ZN(n1285) );
NAND2_X1 U935 ( .A1(KEYINPUT15), .A2(n1286), .ZN(n1280) );
NAND2_X1 U936 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
NAND2_X1 U937 ( .A1(KEYINPUT63), .A2(n1255), .ZN(n1288) );
OR3_X1 U938 ( .A1(G131), .A2(KEYINPUT63), .A3(n1255), .ZN(n1287) );
NAND3_X1 U939 ( .A1(n1278), .A2(n1108), .A3(n1233), .ZN(n1255) );
AND3_X1 U940 ( .A1(n1289), .A2(n1263), .A3(n1099), .ZN(n1278) );
INV_X1 U941 ( .A(n1066), .ZN(n1099) );
NAND2_X1 U942 ( .A1(n1088), .A2(n1093), .ZN(n1066) );
XNOR2_X1 U943 ( .A(G128), .B(n1265), .ZN(G30) );
NAND3_X1 U944 ( .A1(n1241), .A2(n1263), .A3(n1267), .ZN(n1265) );
INV_X1 U945 ( .A(n1264), .ZN(n1267) );
NAND3_X1 U946 ( .A1(n1279), .A2(n1109), .A3(n1239), .ZN(n1264) );
XOR2_X1 U947 ( .A(n1290), .B(n1234), .Z(G3) );
NAND4_X1 U948 ( .A1(n1078), .A2(n1108), .A3(n1239), .A4(n1291), .ZN(n1234) );
NOR2_X1 U949 ( .A1(n1095), .A2(n1086), .ZN(n1239) );
INV_X1 U950 ( .A(n1289), .ZN(n1095) );
XOR2_X1 U951 ( .A(G125), .B(n1260), .Z(G27) );
NOR2_X1 U952 ( .A1(n1261), .A2(n1067), .ZN(n1260) );
NAND4_X1 U953 ( .A1(n1263), .A2(n1109), .A3(n1242), .A4(n1292), .ZN(n1261) );
NOR2_X1 U954 ( .A1(n1103), .A2(n1117), .ZN(n1292) );
NAND2_X1 U955 ( .A1(n1070), .A2(n1293), .ZN(n1263) );
NAND3_X1 U956 ( .A1(G902), .A2(n1294), .A3(n1130), .ZN(n1293) );
NOR2_X1 U957 ( .A1(n1151), .A2(G900), .ZN(n1130) );
XOR2_X1 U958 ( .A(n1237), .B(n1295), .Z(G24) );
XOR2_X1 U959 ( .A(n1296), .B(KEYINPUT36), .Z(n1295) );
NAND4_X1 U960 ( .A1(n1084), .A2(n1240), .A3(n1297), .A4(n1242), .ZN(n1237) );
NOR2_X1 U961 ( .A1(n1298), .A2(n1113), .ZN(n1297) );
AND3_X1 U962 ( .A1(n1080), .A2(n1291), .A3(n1079), .ZN(n1240) );
XOR2_X1 U963 ( .A(G119), .B(n1299), .Z(G21) );
NOR2_X1 U964 ( .A1(n1300), .A2(n1246), .ZN(n1299) );
NAND3_X1 U965 ( .A1(n1084), .A2(n1279), .A3(n1301), .ZN(n1246) );
XOR2_X1 U966 ( .A(n1086), .B(KEYINPUT54), .Z(n1300) );
XNOR2_X1 U967 ( .A(G116), .B(n1238), .ZN(G18) );
NAND2_X1 U968 ( .A1(n1232), .A2(n1241), .ZN(n1238) );
INV_X1 U969 ( .A(n1104), .ZN(n1241) );
NAND2_X1 U970 ( .A1(n1113), .A2(n1121), .ZN(n1104) );
INV_X1 U971 ( .A(n1298), .ZN(n1121) );
AND4_X1 U972 ( .A1(n1108), .A2(n1084), .A3(n1242), .A4(n1291), .ZN(n1232) );
INV_X1 U973 ( .A(n1086), .ZN(n1242) );
INV_X1 U974 ( .A(n1067), .ZN(n1084) );
XOR2_X1 U975 ( .A(G113), .B(n1302), .Z(G15) );
NOR2_X1 U976 ( .A1(n1303), .A2(n1086), .ZN(n1302) );
XOR2_X1 U977 ( .A(n1304), .B(KEYINPUT23), .Z(n1303) );
NAND4_X1 U978 ( .A1(n1305), .A2(n1233), .A3(n1108), .A4(n1291), .ZN(n1304) );
INV_X1 U979 ( .A(n1068), .ZN(n1108) );
NAND2_X1 U980 ( .A1(n1306), .A2(n1079), .ZN(n1068) );
INV_X1 U981 ( .A(n1109), .ZN(n1079) );
XNOR2_X1 U982 ( .A(n1279), .B(KEYINPUT50), .ZN(n1306) );
XNOR2_X1 U983 ( .A(n1080), .B(KEYINPUT21), .ZN(n1279) );
INV_X1 U984 ( .A(n1103), .ZN(n1233) );
NAND2_X1 U985 ( .A1(n1307), .A2(n1277), .ZN(n1103) );
INV_X1 U986 ( .A(n1113), .ZN(n1277) );
XOR2_X1 U987 ( .A(n1067), .B(KEYINPUT44), .Z(n1305) );
NAND2_X1 U988 ( .A1(n1097), .A2(n1308), .ZN(n1067) );
XOR2_X1 U989 ( .A(n1309), .B(n1310), .Z(G12) );
NOR2_X1 U990 ( .A1(KEYINPUT37), .A2(n1311), .ZN(n1310) );
NOR2_X1 U991 ( .A1(n1086), .A2(n1312), .ZN(n1309) );
XNOR2_X1 U992 ( .A(KEYINPUT20), .B(n1247), .ZN(n1312) );
NAND3_X1 U993 ( .A1(n1080), .A2(n1289), .A3(n1301), .ZN(n1247) );
AND3_X1 U994 ( .A1(n1291), .A2(n1109), .A3(n1078), .ZN(n1301) );
INV_X1 U995 ( .A(n1069), .ZN(n1078) );
NAND2_X1 U996 ( .A1(n1307), .A2(n1113), .ZN(n1069) );
XOR2_X1 U997 ( .A(n1313), .B(G475), .Z(n1113) );
NAND2_X1 U998 ( .A1(n1186), .A2(n1184), .ZN(n1313) );
XNOR2_X1 U999 ( .A(n1314), .B(n1315), .ZN(n1186) );
XOR2_X1 U1000 ( .A(G113), .B(n1316), .Z(n1315) );
XOR2_X1 U1001 ( .A(G146), .B(G122), .Z(n1316) );
XOR2_X1 U1002 ( .A(n1317), .B(n1211), .Z(n1314) );
XOR2_X1 U1003 ( .A(G104), .B(G140), .Z(n1211) );
XNOR2_X1 U1004 ( .A(n1318), .B(n1319), .ZN(n1317) );
NOR2_X1 U1005 ( .A1(G125), .A2(KEYINPUT25), .ZN(n1319) );
NOR2_X1 U1006 ( .A1(KEYINPUT38), .A2(n1320), .ZN(n1318) );
XNOR2_X1 U1007 ( .A(n1321), .B(n1322), .ZN(n1320) );
XOR2_X1 U1008 ( .A(G131), .B(n1323), .Z(n1322) );
AND3_X1 U1009 ( .A1(G214), .A2(n1151), .A3(n1324), .ZN(n1323) );
XOR2_X1 U1010 ( .A(KEYINPUT24), .B(n1298), .Z(n1307) );
XOR2_X1 U1011 ( .A(n1325), .B(G478), .Z(n1298) );
NAND2_X1 U1012 ( .A1(n1181), .A2(n1184), .ZN(n1325) );
XOR2_X1 U1013 ( .A(n1326), .B(n1327), .Z(n1181) );
XOR2_X1 U1014 ( .A(n1328), .B(n1329), .Z(n1327) );
XNOR2_X1 U1015 ( .A(G107), .B(n1330), .ZN(n1329) );
NAND2_X1 U1016 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
OR2_X1 U1017 ( .A1(n1321), .A2(n1333), .ZN(n1332) );
XOR2_X1 U1018 ( .A(n1334), .B(KEYINPUT62), .Z(n1331) );
NAND2_X1 U1019 ( .A1(n1333), .A2(n1321), .ZN(n1334) );
AND3_X1 U1020 ( .A1(G234), .A2(n1151), .A3(G217), .ZN(n1328) );
XOR2_X1 U1021 ( .A(n1335), .B(n1336), .Z(n1326) );
XOR2_X1 U1022 ( .A(G122), .B(G116), .Z(n1336) );
XNOR2_X1 U1023 ( .A(G134), .B(KEYINPUT59), .ZN(n1335) );
NAND2_X1 U1024 ( .A1(n1337), .A2(n1125), .ZN(n1109) );
NAND3_X1 U1025 ( .A1(n1338), .A2(n1184), .A3(n1175), .ZN(n1125) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1339), .ZN(n1338) );
INV_X1 U1027 ( .A(G234), .ZN(n1339) );
XNOR2_X1 U1028 ( .A(n1124), .B(KEYINPUT42), .ZN(n1337) );
NOR2_X1 U1029 ( .A1(n1177), .A2(n1340), .ZN(n1124) );
AND2_X1 U1030 ( .A1(n1175), .A2(n1184), .ZN(n1340) );
XNOR2_X1 U1031 ( .A(n1341), .B(n1342), .ZN(n1175) );
XOR2_X1 U1032 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1033 ( .A(G110), .B(n1345), .Z(n1344) );
AND3_X1 U1034 ( .A1(G221), .A2(n1151), .A3(G234), .ZN(n1345) );
XOR2_X1 U1035 ( .A(G137), .B(G119), .Z(n1343) );
XOR2_X1 U1036 ( .A(n1134), .B(n1346), .Z(n1341) );
XNOR2_X1 U1037 ( .A(n1347), .B(n1348), .ZN(n1346) );
NOR2_X1 U1038 ( .A1(KEYINPUT28), .A2(n1333), .ZN(n1348) );
NAND2_X1 U1039 ( .A1(KEYINPUT58), .A2(n1266), .ZN(n1347) );
INV_X1 U1040 ( .A(G146), .ZN(n1266) );
XNOR2_X1 U1041 ( .A(G125), .B(G140), .ZN(n1134) );
NAND2_X1 U1042 ( .A1(G217), .A2(n1349), .ZN(n1177) );
NAND2_X1 U1043 ( .A1(n1070), .A2(n1350), .ZN(n1291) );
NAND3_X1 U1044 ( .A1(n1351), .A2(n1294), .A3(G902), .ZN(n1350) );
INV_X1 U1045 ( .A(n1163), .ZN(n1351) );
NAND2_X1 U1046 ( .A1(n1352), .A2(G953), .ZN(n1163) );
XNOR2_X1 U1047 ( .A(G898), .B(KEYINPUT13), .ZN(n1352) );
NAND3_X1 U1048 ( .A1(n1294), .A2(n1151), .A3(n1353), .ZN(n1070) );
XNOR2_X1 U1049 ( .A(G952), .B(KEYINPUT29), .ZN(n1353) );
NAND2_X1 U1050 ( .A1(G237), .A2(G234), .ZN(n1294) );
NOR2_X1 U1051 ( .A1(n1097), .A2(n1096), .ZN(n1289) );
INV_X1 U1052 ( .A(n1308), .ZN(n1096) );
NAND2_X1 U1053 ( .A1(G221), .A2(n1349), .ZN(n1308) );
NAND2_X1 U1054 ( .A1(G234), .A2(n1184), .ZN(n1349) );
XOR2_X1 U1055 ( .A(n1354), .B(G469), .Z(n1097) );
NAND2_X1 U1056 ( .A1(n1355), .A2(n1184), .ZN(n1354) );
XOR2_X1 U1057 ( .A(n1356), .B(n1357), .Z(n1355) );
XOR2_X1 U1058 ( .A(n1204), .B(n1214), .Z(n1357) );
XOR2_X1 U1059 ( .A(G107), .B(n1358), .Z(n1214) );
NOR2_X1 U1060 ( .A1(G101), .A2(KEYINPUT46), .ZN(n1358) );
INV_X1 U1061 ( .A(n1203), .ZN(n1204) );
XOR2_X1 U1062 ( .A(n1359), .B(n1360), .Z(n1356) );
XOR2_X1 U1063 ( .A(n1361), .B(G104), .Z(n1360) );
NAND3_X1 U1064 ( .A1(n1362), .A2(n1363), .A3(KEYINPUT3), .ZN(n1361) );
NAND2_X1 U1065 ( .A1(n1364), .A2(n1219), .ZN(n1363) );
XOR2_X1 U1066 ( .A(KEYINPUT7), .B(n1365), .Z(n1362) );
NOR2_X1 U1067 ( .A1(n1219), .A2(n1364), .ZN(n1365) );
XOR2_X1 U1068 ( .A(G140), .B(G110), .Z(n1364) );
NAND2_X1 U1069 ( .A1(G227), .A2(n1151), .ZN(n1219) );
NAND2_X1 U1070 ( .A1(KEYINPUT40), .A2(n1213), .ZN(n1359) );
INV_X1 U1071 ( .A(n1138), .ZN(n1213) );
XOR2_X1 U1072 ( .A(n1333), .B(n1366), .Z(n1138) );
INV_X1 U1073 ( .A(n1117), .ZN(n1080) );
XOR2_X1 U1074 ( .A(n1119), .B(G472), .Z(n1117) );
AND2_X1 U1075 ( .A1(n1367), .A2(n1184), .ZN(n1119) );
XOR2_X1 U1076 ( .A(n1368), .B(n1369), .Z(n1367) );
XOR2_X1 U1077 ( .A(n1202), .B(n1203), .Z(n1369) );
XOR2_X1 U1078 ( .A(n1370), .B(n1146), .Z(n1203) );
XOR2_X1 U1079 ( .A(G134), .B(G137), .Z(n1146) );
XOR2_X1 U1080 ( .A(n1145), .B(KEYINPUT33), .Z(n1370) );
INV_X1 U1081 ( .A(G131), .ZN(n1145) );
XNOR2_X1 U1082 ( .A(n1198), .B(n1371), .ZN(n1368) );
XOR2_X1 U1083 ( .A(n1207), .B(n1372), .Z(n1371) );
NAND2_X1 U1084 ( .A1(KEYINPUT55), .A2(n1290), .ZN(n1372) );
NAND3_X1 U1085 ( .A1(G210), .A2(n1151), .A3(n1373), .ZN(n1207) );
XOR2_X1 U1086 ( .A(n1324), .B(KEYINPUT30), .Z(n1373) );
XNOR2_X1 U1087 ( .A(n1374), .B(G113), .ZN(n1198) );
NAND2_X1 U1088 ( .A1(n1375), .A2(KEYINPUT0), .ZN(n1374) );
XNOR2_X1 U1089 ( .A(G116), .B(n1376), .ZN(n1375) );
NOR2_X1 U1090 ( .A1(G119), .A2(KEYINPUT12), .ZN(n1376) );
NAND2_X1 U1091 ( .A1(n1377), .A2(n1093), .ZN(n1086) );
NAND2_X1 U1092 ( .A1(G214), .A2(n1378), .ZN(n1093) );
INV_X1 U1093 ( .A(n1088), .ZN(n1377) );
XNOR2_X1 U1094 ( .A(n1379), .B(n1230), .ZN(n1088) );
NAND2_X1 U1095 ( .A1(G210), .A2(n1378), .ZN(n1230) );
NAND2_X1 U1096 ( .A1(n1324), .A2(n1184), .ZN(n1378) );
INV_X1 U1097 ( .A(G237), .ZN(n1324) );
NAND3_X1 U1098 ( .A1(n1380), .A2(n1381), .A3(n1184), .ZN(n1379) );
INV_X1 U1099 ( .A(G902), .ZN(n1184) );
NAND2_X1 U1100 ( .A1(KEYINPUT18), .A2(n1382), .ZN(n1381) );
NAND2_X1 U1101 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
NAND2_X1 U1102 ( .A1(n1229), .A2(n1228), .ZN(n1384) );
INV_X1 U1103 ( .A(n1225), .ZN(n1383) );
NOR2_X1 U1104 ( .A1(n1228), .A2(n1229), .ZN(n1225) );
NAND2_X1 U1105 ( .A1(n1385), .A2(n1386), .ZN(n1380) );
INV_X1 U1106 ( .A(KEYINPUT18), .ZN(n1386) );
XOR2_X1 U1107 ( .A(n1229), .B(n1228), .Z(n1385) );
NAND2_X1 U1108 ( .A1(n1166), .A2(n1162), .ZN(n1228) );
NAND2_X1 U1109 ( .A1(n1387), .A2(n1168), .ZN(n1162) );
AND2_X1 U1110 ( .A1(n1388), .A2(n1389), .ZN(n1166) );
OR3_X1 U1111 ( .A1(n1390), .A2(n1387), .A3(n1168), .ZN(n1389) );
NOR2_X1 U1112 ( .A1(n1391), .A2(n1169), .ZN(n1387) );
AND2_X1 U1113 ( .A1(n1169), .A2(n1391), .ZN(n1390) );
NAND3_X1 U1114 ( .A1(n1169), .A2(n1391), .A3(n1168), .ZN(n1388) );
XOR2_X1 U1115 ( .A(n1296), .B(n1311), .Z(n1168) );
INV_X1 U1116 ( .A(G110), .ZN(n1311) );
INV_X1 U1117 ( .A(G122), .ZN(n1296) );
XNOR2_X1 U1118 ( .A(n1290), .B(n1392), .ZN(n1391) );
NOR2_X1 U1119 ( .A1(KEYINPUT2), .A2(n1393), .ZN(n1392) );
XOR2_X1 U1120 ( .A(n1189), .B(G107), .Z(n1393) );
INV_X1 U1121 ( .A(G104), .ZN(n1189) );
INV_X1 U1122 ( .A(G101), .ZN(n1290) );
XOR2_X1 U1123 ( .A(G113), .B(n1394), .Z(n1169) );
XOR2_X1 U1124 ( .A(G119), .B(G116), .Z(n1394) );
XNOR2_X1 U1125 ( .A(n1395), .B(n1396), .ZN(n1229) );
XNOR2_X1 U1126 ( .A(n1397), .B(n1202), .ZN(n1396) );
XOR2_X1 U1127 ( .A(n1398), .B(n1366), .Z(n1202) );
XOR2_X1 U1128 ( .A(G146), .B(n1321), .Z(n1366) );
XNOR2_X1 U1129 ( .A(n1271), .B(KEYINPUT57), .ZN(n1321) );
INV_X1 U1130 ( .A(G143), .ZN(n1271) );
NAND2_X1 U1131 ( .A1(KEYINPUT19), .A2(n1399), .ZN(n1398) );
INV_X1 U1132 ( .A(n1333), .ZN(n1399) );
XNOR2_X1 U1133 ( .A(G128), .B(KEYINPUT52), .ZN(n1333) );
AND2_X1 U1134 ( .A1(n1151), .A2(G224), .ZN(n1397) );
INV_X1 U1135 ( .A(G953), .ZN(n1151) );
XNOR2_X1 U1136 ( .A(G125), .B(KEYINPUT61), .ZN(n1395) );
endmodule


