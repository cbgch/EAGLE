//Key = 0100011011101111000000100100001001010001101111011101111110000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354;

XNOR2_X1 U735 ( .A(G107), .B(n1031), .ZN(G9) );
NAND2_X1 U736 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U737 ( .A1(n1034), .A2(n1035), .ZN(G75) );
NOR3_X1 U738 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NAND3_X1 U739 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1036) );
NAND2_X1 U740 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U741 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND4_X1 U742 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1045) );
NAND2_X1 U743 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U744 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U745 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U746 ( .A1(n1056), .A2(n1057), .ZN(n1050) );
NAND2_X1 U747 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U748 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND3_X1 U749 ( .A1(n1052), .A2(n1062), .A3(n1056), .ZN(n1044) );
NAND2_X1 U750 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U751 ( .A1(n1065), .A2(n1066), .A3(n1048), .ZN(n1064) );
OR2_X1 U752 ( .A1(n1046), .A2(n1047), .ZN(n1066) );
NAND3_X1 U753 ( .A1(n1067), .A2(n1068), .A3(n1046), .ZN(n1065) );
OR2_X1 U754 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
INV_X1 U755 ( .A(n1071), .ZN(n1042) );
NOR3_X1 U756 ( .A1(n1072), .A2(G953), .A3(n1073), .ZN(n1034) );
INV_X1 U757 ( .A(n1039), .ZN(n1073) );
NAND4_X1 U758 ( .A1(n1061), .A2(n1046), .A3(n1074), .A4(n1075), .ZN(n1039) );
NOR3_X1 U759 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NAND3_X1 U760 ( .A1(n1079), .A2(n1069), .A3(n1080), .ZN(n1076) );
NAND2_X1 U761 ( .A1(KEYINPUT27), .A2(n1081), .ZN(n1080) );
NOR3_X1 U762 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1074) );
NOR2_X1 U763 ( .A1(G475), .A2(n1085), .ZN(n1084) );
NOR2_X1 U764 ( .A1(KEYINPUT27), .A2(n1086), .ZN(n1085) );
XNOR2_X1 U765 ( .A(n1081), .B(KEYINPUT14), .ZN(n1086) );
NOR3_X1 U766 ( .A1(n1087), .A2(KEYINPUT27), .A3(n1081), .ZN(n1083) );
XNOR2_X1 U767 ( .A(KEYINPUT50), .B(n1088), .ZN(n1082) );
XNOR2_X1 U768 ( .A(KEYINPUT59), .B(n1037), .ZN(n1072) );
INV_X1 U769 ( .A(G952), .ZN(n1037) );
XOR2_X1 U770 ( .A(n1089), .B(n1090), .Z(G72) );
NOR2_X1 U771 ( .A1(n1091), .A2(n1040), .ZN(n1090) );
AND2_X1 U772 ( .A1(G227), .A2(G900), .ZN(n1091) );
NAND3_X1 U773 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1089) );
OR2_X1 U774 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND3_X1 U775 ( .A1(n1096), .A2(n1095), .A3(KEYINPUT51), .ZN(n1093) );
NAND2_X1 U776 ( .A1(KEYINPUT22), .A2(n1097), .ZN(n1096) );
NAND2_X1 U777 ( .A1(n1098), .A2(n1099), .ZN(n1092) );
INV_X1 U778 ( .A(KEYINPUT51), .ZN(n1099) );
NAND2_X1 U779 ( .A1(n1100), .A2(n1095), .ZN(n1098) );
NAND2_X1 U780 ( .A1(n1101), .A2(n1102), .ZN(n1095) );
NAND2_X1 U781 ( .A1(G953), .A2(n1103), .ZN(n1102) );
XOR2_X1 U782 ( .A(n1104), .B(n1105), .Z(n1101) );
XNOR2_X1 U783 ( .A(n1106), .B(n1107), .ZN(n1105) );
NAND2_X1 U784 ( .A1(KEYINPUT40), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U785 ( .A(n1109), .B(n1110), .ZN(n1104) );
NOR3_X1 U786 ( .A1(KEYINPUT60), .A2(n1111), .A3(n1112), .ZN(n1110) );
NOR2_X1 U787 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XNOR2_X1 U788 ( .A(n1115), .B(KEYINPUT63), .ZN(n1114) );
NOR2_X1 U789 ( .A1(G137), .A2(n1116), .ZN(n1111) );
XOR2_X1 U790 ( .A(KEYINPUT43), .B(n1115), .Z(n1116) );
XOR2_X1 U791 ( .A(G131), .B(n1117), .Z(n1115) );
INV_X1 U792 ( .A(n1097), .ZN(n1100) );
NAND2_X1 U793 ( .A1(n1040), .A2(n1118), .ZN(n1097) );
OR4_X1 U794 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1118) );
AND2_X1 U795 ( .A1(n1123), .A2(n1124), .ZN(n1120) );
NAND2_X1 U796 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XOR2_X1 U797 ( .A(n1127), .B(n1128), .Z(G69) );
XOR2_X1 U798 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U799 ( .A1(n1040), .A2(n1131), .ZN(n1130) );
NAND3_X1 U800 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
XNOR2_X1 U801 ( .A(n1135), .B(KEYINPUT52), .ZN(n1134) );
INV_X1 U802 ( .A(n1136), .ZN(n1133) );
XNOR2_X1 U803 ( .A(n1137), .B(KEYINPUT62), .ZN(n1132) );
NAND4_X1 U804 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1129) );
NAND3_X1 U805 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1141) );
NAND3_X1 U806 ( .A1(KEYINPUT13), .A2(n1145), .A3(n1146), .ZN(n1140) );
NAND2_X1 U807 ( .A1(G953), .A2(n1147), .ZN(n1139) );
XNOR2_X1 U808 ( .A(KEYINPUT49), .B(n1148), .ZN(n1147) );
NAND3_X1 U809 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1138) );
NAND2_X1 U810 ( .A1(n1146), .A2(KEYINPUT13), .ZN(n1150) );
NAND2_X1 U811 ( .A1(n1144), .A2(n1143), .ZN(n1149) );
NAND2_X1 U812 ( .A1(KEYINPUT13), .A2(n1152), .ZN(n1143) );
NOR2_X1 U813 ( .A1(n1153), .A2(n1040), .ZN(n1127) );
NOR2_X1 U814 ( .A1(n1154), .A2(n1148), .ZN(n1153) );
NOR2_X1 U815 ( .A1(n1155), .A2(n1156), .ZN(G66) );
XOR2_X1 U816 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U817 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NOR2_X1 U818 ( .A1(n1155), .A2(n1161), .ZN(G63) );
XOR2_X1 U819 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR3_X1 U820 ( .A1(n1160), .A2(KEYINPUT41), .A3(n1164), .ZN(n1162) );
NOR2_X1 U821 ( .A1(n1155), .A2(n1165), .ZN(G60) );
XOR2_X1 U822 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U823 ( .A1(KEYINPUT3), .A2(n1168), .ZN(n1167) );
NOR2_X1 U824 ( .A1(n1087), .A2(n1160), .ZN(n1166) );
XNOR2_X1 U825 ( .A(G104), .B(n1169), .ZN(G6) );
NAND2_X1 U826 ( .A1(n1123), .A2(n1033), .ZN(n1169) );
NOR2_X1 U827 ( .A1(n1155), .A2(n1170), .ZN(G57) );
XOR2_X1 U828 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U829 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U830 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U831 ( .A1(n1177), .A2(n1160), .ZN(n1176) );
NOR2_X1 U832 ( .A1(n1178), .A2(n1179), .ZN(n1175) );
NOR2_X1 U833 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NOR2_X1 U834 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NOR2_X1 U835 ( .A1(G101), .A2(n1184), .ZN(n1180) );
AND2_X1 U836 ( .A1(n1182), .A2(KEYINPUT7), .ZN(n1184) );
NOR4_X1 U837 ( .A1(KEYINPUT7), .A2(G101), .A3(n1182), .A4(n1183), .ZN(n1178) );
INV_X1 U838 ( .A(KEYINPUT44), .ZN(n1183) );
NOR2_X1 U839 ( .A1(KEYINPUT34), .A2(n1142), .ZN(n1173) );
XNOR2_X1 U840 ( .A(n1117), .B(n1185), .ZN(n1171) );
NOR2_X1 U841 ( .A1(n1155), .A2(n1186), .ZN(G54) );
XOR2_X1 U842 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U843 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U844 ( .A(n1191), .B(n1192), .Z(n1190) );
NOR2_X1 U845 ( .A1(n1193), .A2(n1160), .ZN(n1192) );
NAND2_X1 U846 ( .A1(KEYINPUT6), .A2(n1194), .ZN(n1191) );
NAND2_X1 U847 ( .A1(KEYINPUT48), .A2(n1195), .ZN(n1189) );
XNOR2_X1 U848 ( .A(n1107), .B(n1196), .ZN(n1187) );
NOR2_X1 U849 ( .A1(n1040), .A2(G952), .ZN(n1155) );
NOR2_X1 U850 ( .A1(n1197), .A2(n1198), .ZN(G51) );
XNOR2_X1 U851 ( .A(n1199), .B(n1200), .ZN(n1198) );
XOR2_X1 U852 ( .A(n1201), .B(n1202), .Z(n1200) );
NOR2_X1 U853 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
INV_X1 U854 ( .A(n1205), .ZN(n1203) );
NOR4_X1 U855 ( .A1(KEYINPUT37), .A2(n1206), .A3(n1207), .A4(n1160), .ZN(n1201) );
NAND2_X1 U856 ( .A1(G902), .A2(n1038), .ZN(n1160) );
NAND4_X1 U857 ( .A1(n1208), .A2(n1135), .A3(n1209), .A4(n1210), .ZN(n1038) );
NOR4_X1 U858 ( .A1(n1137), .A2(n1122), .A3(n1121), .A4(n1211), .ZN(n1210) );
NOR2_X1 U859 ( .A1(n1054), .A2(n1125), .ZN(n1211) );
NOR2_X1 U860 ( .A1(n1136), .A2(n1119), .ZN(n1209) );
NAND4_X1 U861 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1119) );
OR2_X1 U862 ( .A1(n1125), .A2(n1055), .ZN(n1212) );
NAND3_X1 U863 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1136) );
NAND4_X1 U864 ( .A1(n1219), .A2(n1032), .A3(n1220), .A4(n1221), .ZN(n1218) );
XOR2_X1 U865 ( .A(KEYINPUT18), .B(n1047), .Z(n1221) );
INV_X1 U866 ( .A(n1055), .ZN(n1032) );
AND3_X1 U867 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1135) );
NAND2_X1 U868 ( .A1(n1033), .A2(n1225), .ZN(n1224) );
NAND2_X1 U869 ( .A1(n1226), .A2(n1054), .ZN(n1225) );
XNOR2_X1 U870 ( .A(KEYINPUT12), .B(n1055), .ZN(n1226) );
AND2_X1 U871 ( .A1(n1227), .A2(n1046), .ZN(n1033) );
XOR2_X1 U872 ( .A(n1228), .B(KEYINPUT4), .Z(n1208) );
OR2_X1 U873 ( .A1(n1126), .A2(n1054), .ZN(n1228) );
NOR2_X1 U874 ( .A1(n1229), .A2(n1040), .ZN(n1197) );
XNOR2_X1 U875 ( .A(G952), .B(KEYINPUT1), .ZN(n1229) );
XOR2_X1 U876 ( .A(n1230), .B(n1231), .Z(G48) );
NOR2_X1 U877 ( .A1(n1126), .A2(n1232), .ZN(n1231) );
XNOR2_X1 U878 ( .A(KEYINPUT56), .B(n1054), .ZN(n1232) );
XNOR2_X1 U879 ( .A(G146), .B(KEYINPUT53), .ZN(n1230) );
XOR2_X1 U880 ( .A(G143), .B(n1121), .Z(G45) );
AND3_X1 U881 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(n1121) );
NOR3_X1 U882 ( .A1(n1088), .A2(n1236), .A3(n1237), .ZN(n1235) );
XNOR2_X1 U883 ( .A(G140), .B(n1213), .ZN(G42) );
NAND4_X1 U884 ( .A1(n1238), .A2(n1123), .A3(n1052), .A4(n1048), .ZN(n1213) );
XNOR2_X1 U885 ( .A(G137), .B(n1214), .ZN(G39) );
NAND4_X1 U886 ( .A1(n1056), .A2(n1238), .A3(n1052), .A4(n1077), .ZN(n1214) );
XOR2_X1 U887 ( .A(G134), .B(n1239), .Z(G36) );
NOR2_X1 U888 ( .A1(n1055), .A2(n1125), .ZN(n1239) );
NAND3_X1 U889 ( .A1(n1052), .A2(n1240), .A3(n1233), .ZN(n1125) );
XNOR2_X1 U890 ( .A(G131), .B(n1241), .ZN(G33) );
NAND4_X1 U891 ( .A1(n1242), .A2(n1233), .A3(n1123), .A4(n1052), .ZN(n1241) );
NAND2_X1 U892 ( .A1(n1243), .A2(n1244), .ZN(n1052) );
OR2_X1 U893 ( .A1(n1058), .A2(KEYINPUT10), .ZN(n1244) );
INV_X1 U894 ( .A(n1234), .ZN(n1058) );
NAND3_X1 U895 ( .A1(n1061), .A2(n1079), .A3(KEYINPUT10), .ZN(n1243) );
INV_X1 U896 ( .A(n1060), .ZN(n1079) );
XNOR2_X1 U897 ( .A(n1236), .B(KEYINPUT23), .ZN(n1242) );
XOR2_X1 U898 ( .A(G128), .B(n1122), .Z(G30) );
NOR2_X1 U899 ( .A1(n1126), .A2(n1055), .ZN(n1122) );
NAND3_X1 U900 ( .A1(n1234), .A2(n1077), .A3(n1238), .ZN(n1126) );
NOR3_X1 U901 ( .A1(n1046), .A2(n1236), .A3(n1068), .ZN(n1238) );
XOR2_X1 U902 ( .A(n1222), .B(n1245), .Z(G3) );
NAND2_X1 U903 ( .A1(KEYINPUT35), .A2(G101), .ZN(n1245) );
NAND3_X1 U904 ( .A1(n1233), .A2(n1220), .A3(n1056), .ZN(n1222) );
NOR2_X1 U905 ( .A1(n1246), .A2(n1068), .ZN(n1233) );
XNOR2_X1 U906 ( .A(G125), .B(n1215), .ZN(G27) );
NAND4_X1 U907 ( .A1(n1047), .A2(n1234), .A3(n1123), .A4(n1247), .ZN(n1215) );
NOR3_X1 U908 ( .A1(n1046), .A2(n1236), .A3(n1248), .ZN(n1247) );
INV_X1 U909 ( .A(n1240), .ZN(n1236) );
NAND2_X1 U910 ( .A1(n1071), .A2(n1249), .ZN(n1240) );
NAND4_X1 U911 ( .A1(G953), .A2(G902), .A3(n1250), .A4(n1103), .ZN(n1249) );
INV_X1 U912 ( .A(G900), .ZN(n1103) );
XNOR2_X1 U913 ( .A(G122), .B(n1216), .ZN(G24) );
NAND4_X1 U914 ( .A1(n1046), .A2(n1220), .A3(n1047), .A4(n1251), .ZN(n1216) );
NOR3_X1 U915 ( .A1(n1248), .A2(n1237), .A3(n1088), .ZN(n1251) );
XNOR2_X1 U916 ( .A(G119), .B(n1217), .ZN(G21) );
NAND4_X1 U917 ( .A1(n1056), .A2(n1047), .A3(n1252), .A4(n1220), .ZN(n1217) );
INV_X1 U918 ( .A(n1253), .ZN(n1220) );
AND2_X1 U919 ( .A1(n1077), .A2(n1254), .ZN(n1252) );
XOR2_X1 U920 ( .A(n1255), .B(n1256), .Z(G18) );
NOR3_X1 U921 ( .A1(n1257), .A2(n1253), .A3(n1063), .ZN(n1256) );
XNOR2_X1 U922 ( .A(KEYINPUT9), .B(n1055), .ZN(n1257) );
NAND2_X1 U923 ( .A1(n1237), .A2(n1258), .ZN(n1055) );
NAND2_X1 U924 ( .A1(KEYINPUT54), .A2(n1259), .ZN(n1255) );
INV_X1 U925 ( .A(G116), .ZN(n1259) );
XOR2_X1 U926 ( .A(G113), .B(n1260), .Z(G15) );
NOR2_X1 U927 ( .A1(KEYINPUT20), .A2(n1261), .ZN(n1260) );
INV_X1 U928 ( .A(n1137), .ZN(n1261) );
NOR3_X1 U929 ( .A1(n1054), .A2(n1253), .A3(n1063), .ZN(n1137) );
NAND2_X1 U930 ( .A1(n1219), .A2(n1047), .ZN(n1063) );
NOR2_X1 U931 ( .A1(n1070), .A2(n1262), .ZN(n1047) );
INV_X1 U932 ( .A(n1069), .ZN(n1262) );
INV_X1 U933 ( .A(n1246), .ZN(n1219) );
NAND2_X1 U934 ( .A1(n1046), .A2(n1077), .ZN(n1246) );
INV_X1 U935 ( .A(n1254), .ZN(n1046) );
INV_X1 U936 ( .A(n1123), .ZN(n1054) );
NOR2_X1 U937 ( .A1(n1258), .A2(n1237), .ZN(n1123) );
XNOR2_X1 U938 ( .A(G110), .B(n1223), .ZN(G12) );
NAND3_X1 U939 ( .A1(n1227), .A2(n1254), .A3(n1056), .ZN(n1223) );
AND2_X1 U940 ( .A1(n1088), .A2(n1237), .ZN(n1056) );
XNOR2_X1 U941 ( .A(n1081), .B(n1263), .ZN(n1237) );
XNOR2_X1 U942 ( .A(KEYINPUT2), .B(n1087), .ZN(n1263) );
INV_X1 U943 ( .A(G475), .ZN(n1087) );
AND2_X1 U944 ( .A1(n1168), .A2(n1264), .ZN(n1081) );
XNOR2_X1 U945 ( .A(n1265), .B(n1266), .ZN(n1168) );
XOR2_X1 U946 ( .A(G104), .B(n1267), .Z(n1266) );
NOR2_X1 U947 ( .A1(KEYINPUT46), .A2(n1268), .ZN(n1267) );
XOR2_X1 U948 ( .A(n1269), .B(n1270), .Z(n1268) );
XNOR2_X1 U949 ( .A(n1271), .B(n1272), .ZN(n1270) );
XNOR2_X1 U950 ( .A(n1273), .B(G143), .ZN(n1272) );
XNOR2_X1 U951 ( .A(n1274), .B(n1275), .ZN(n1269) );
NOR4_X1 U952 ( .A1(KEYINPUT24), .A2(G953), .A3(G237), .A4(n1276), .ZN(n1275) );
NOR2_X1 U953 ( .A1(KEYINPUT31), .A2(n1277), .ZN(n1274) );
XOR2_X1 U954 ( .A(n1278), .B(n1108), .Z(n1277) );
XNOR2_X1 U955 ( .A(G113), .B(G122), .ZN(n1265) );
INV_X1 U956 ( .A(n1258), .ZN(n1088) );
XOR2_X1 U957 ( .A(n1279), .B(n1164), .Z(n1258) );
INV_X1 U958 ( .A(G478), .ZN(n1164) );
OR2_X1 U959 ( .A1(n1163), .A2(G902), .ZN(n1279) );
XNOR2_X1 U960 ( .A(n1280), .B(n1281), .ZN(n1163) );
XOR2_X1 U961 ( .A(n1282), .B(n1283), .Z(n1281) );
XNOR2_X1 U962 ( .A(G107), .B(G122), .ZN(n1283) );
NAND2_X1 U963 ( .A1(n1284), .A2(n1285), .ZN(n1282) );
XOR2_X1 U964 ( .A(KEYINPUT28), .B(G217), .Z(n1285) );
XOR2_X1 U965 ( .A(n1286), .B(n1287), .Z(n1280) );
XOR2_X1 U966 ( .A(n1288), .B(n1159), .Z(n1254) );
NAND2_X1 U967 ( .A1(G217), .A2(n1289), .ZN(n1159) );
OR2_X1 U968 ( .A1(n1158), .A2(G902), .ZN(n1288) );
XNOR2_X1 U969 ( .A(n1290), .B(n1291), .ZN(n1158) );
XNOR2_X1 U970 ( .A(G137), .B(n1292), .ZN(n1291) );
NAND2_X1 U971 ( .A1(n1293), .A2(KEYINPUT25), .ZN(n1292) );
XOR2_X1 U972 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U973 ( .A(n1296), .B(G110), .ZN(n1295) );
INV_X1 U974 ( .A(G119), .ZN(n1296) );
XOR2_X1 U975 ( .A(n1297), .B(n1298), .Z(n1294) );
NAND3_X1 U976 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1297) );
NAND2_X1 U977 ( .A1(KEYINPUT17), .A2(n1302), .ZN(n1301) );
NAND3_X1 U978 ( .A1(n1303), .A2(n1304), .A3(n1273), .ZN(n1300) );
INV_X1 U979 ( .A(KEYINPUT17), .ZN(n1304) );
OR2_X1 U980 ( .A1(n1273), .A2(n1303), .ZN(n1299) );
NOR2_X1 U981 ( .A1(KEYINPUT57), .A2(n1302), .ZN(n1303) );
XNOR2_X1 U982 ( .A(n1108), .B(n1305), .ZN(n1302) );
NOR2_X1 U983 ( .A1(KEYINPUT26), .A2(n1278), .ZN(n1305) );
XOR2_X1 U984 ( .A(G140), .B(KEYINPUT38), .Z(n1278) );
NAND2_X1 U985 ( .A1(G221), .A2(n1284), .ZN(n1290) );
AND2_X1 U986 ( .A1(G234), .A2(n1040), .ZN(n1284) );
NOR3_X1 U987 ( .A1(n1253), .A2(n1248), .A3(n1068), .ZN(n1227) );
NAND2_X1 U988 ( .A1(n1070), .A2(n1069), .ZN(n1068) );
NAND2_X1 U989 ( .A1(G221), .A2(n1289), .ZN(n1069) );
NAND2_X1 U990 ( .A1(n1306), .A2(G234), .ZN(n1289) );
INV_X1 U991 ( .A(n1307), .ZN(n1306) );
XOR2_X1 U992 ( .A(n1078), .B(n1308), .Z(n1070) );
XOR2_X1 U993 ( .A(KEYINPUT21), .B(KEYINPUT19), .Z(n1308) );
XOR2_X1 U994 ( .A(n1309), .B(n1193), .Z(n1078) );
INV_X1 U995 ( .A(G469), .ZN(n1193) );
NAND2_X1 U996 ( .A1(n1310), .A2(n1264), .ZN(n1309) );
XOR2_X1 U997 ( .A(n1311), .B(n1312), .Z(n1310) );
XNOR2_X1 U998 ( .A(n1107), .B(n1194), .ZN(n1312) );
XOR2_X1 U999 ( .A(n1313), .B(G101), .Z(n1194) );
NAND2_X1 U1000 ( .A1(KEYINPUT61), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1001 ( .A(KEYINPUT42), .B(n1315), .Z(n1314) );
XNOR2_X1 U1002 ( .A(n1287), .B(n1273), .ZN(n1107) );
XOR2_X1 U1003 ( .A(G143), .B(n1298), .Z(n1287) );
XOR2_X1 U1004 ( .A(n1316), .B(n1196), .Z(n1311) );
XNOR2_X1 U1005 ( .A(n1317), .B(n1318), .ZN(n1196) );
XNOR2_X1 U1006 ( .A(n1109), .B(G110), .ZN(n1318) );
INV_X1 U1007 ( .A(G140), .ZN(n1109) );
NAND2_X1 U1008 ( .A1(G227), .A2(n1040), .ZN(n1317) );
NAND2_X1 U1009 ( .A1(KEYINPUT8), .A2(n1195), .ZN(n1316) );
XNOR2_X1 U1010 ( .A(n1319), .B(n1117), .ZN(n1195) );
INV_X1 U1011 ( .A(n1048), .ZN(n1248) );
XOR2_X1 U1012 ( .A(n1077), .B(KEYINPUT55), .Z(n1048) );
XOR2_X1 U1013 ( .A(n1320), .B(n1177), .Z(n1077) );
INV_X1 U1014 ( .A(G472), .ZN(n1177) );
NAND2_X1 U1015 ( .A1(n1321), .A2(n1264), .ZN(n1320) );
XOR2_X1 U1016 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1017 ( .A(n1185), .B(n1324), .ZN(n1323) );
XOR2_X1 U1018 ( .A(n1286), .B(n1325), .Z(n1324) );
XNOR2_X1 U1019 ( .A(G116), .B(n1117), .ZN(n1286) );
XOR2_X1 U1020 ( .A(G134), .B(KEYINPUT58), .Z(n1117) );
XOR2_X1 U1021 ( .A(n1326), .B(n1327), .Z(n1185) );
INV_X1 U1022 ( .A(n1319), .ZN(n1327) );
XOR2_X1 U1023 ( .A(n1328), .B(n1113), .Z(n1319) );
INV_X1 U1024 ( .A(G137), .ZN(n1113) );
NAND2_X1 U1025 ( .A1(KEYINPUT5), .A2(n1271), .ZN(n1328) );
INV_X1 U1026 ( .A(G131), .ZN(n1271) );
XOR2_X1 U1027 ( .A(n1182), .B(n1329), .Z(n1322) );
XNOR2_X1 U1028 ( .A(G101), .B(KEYINPUT39), .ZN(n1329) );
OR3_X1 U1029 ( .A1(G237), .A2(G953), .A3(n1207), .ZN(n1182) );
NAND2_X1 U1030 ( .A1(n1234), .A2(n1330), .ZN(n1253) );
NAND2_X1 U1031 ( .A1(n1331), .A2(n1071), .ZN(n1330) );
NAND3_X1 U1032 ( .A1(n1250), .A2(n1040), .A3(G952), .ZN(n1071) );
INV_X1 U1033 ( .A(G953), .ZN(n1040) );
NAND4_X1 U1034 ( .A1(G953), .A2(G902), .A3(n1250), .A4(n1148), .ZN(n1331) );
INV_X1 U1035 ( .A(G898), .ZN(n1148) );
NAND2_X1 U1036 ( .A1(G237), .A2(G234), .ZN(n1250) );
NOR2_X1 U1037 ( .A1(n1061), .A2(n1060), .ZN(n1234) );
NOR2_X1 U1038 ( .A1(n1276), .A2(n1206), .ZN(n1060) );
INV_X1 U1039 ( .A(G214), .ZN(n1276) );
XOR2_X1 U1040 ( .A(n1332), .B(n1333), .Z(n1061) );
NOR2_X1 U1041 ( .A1(n1206), .A2(n1207), .ZN(n1333) );
INV_X1 U1042 ( .A(G210), .ZN(n1207) );
NOR2_X1 U1043 ( .A1(n1307), .A2(G237), .ZN(n1206) );
XOR2_X1 U1044 ( .A(G902), .B(KEYINPUT0), .Z(n1307) );
NAND2_X1 U1045 ( .A1(n1334), .A2(n1264), .ZN(n1332) );
INV_X1 U1046 ( .A(G902), .ZN(n1264) );
XOR2_X1 U1047 ( .A(n1335), .B(n1199), .Z(n1334) );
XNOR2_X1 U1048 ( .A(n1145), .B(n1144), .ZN(n1199) );
INV_X1 U1049 ( .A(n1146), .ZN(n1144) );
XNOR2_X1 U1050 ( .A(n1336), .B(G110), .ZN(n1146) );
NAND2_X1 U1051 ( .A1(KEYINPUT30), .A2(n1337), .ZN(n1336) );
INV_X1 U1052 ( .A(G122), .ZN(n1337) );
XNOR2_X1 U1053 ( .A(n1152), .B(n1142), .ZN(n1145) );
INV_X1 U1054 ( .A(n1151), .ZN(n1142) );
XOR2_X1 U1055 ( .A(G116), .B(n1325), .Z(n1151) );
XOR2_X1 U1056 ( .A(G113), .B(G119), .Z(n1325) );
XOR2_X1 U1057 ( .A(n1315), .B(n1338), .Z(n1152) );
NOR2_X1 U1058 ( .A1(G101), .A2(KEYINPUT36), .ZN(n1338) );
XOR2_X1 U1059 ( .A(G104), .B(n1339), .Z(n1315) );
XNOR2_X1 U1060 ( .A(KEYINPUT45), .B(n1340), .ZN(n1339) );
INV_X1 U1061 ( .A(G107), .ZN(n1340) );
XOR2_X1 U1062 ( .A(n1341), .B(KEYINPUT33), .Z(n1335) );
NAND3_X1 U1063 ( .A1(n1342), .A2(n1343), .A3(n1205), .ZN(n1341) );
NAND2_X1 U1064 ( .A1(n1344), .A2(n1345), .ZN(n1205) );
NAND2_X1 U1065 ( .A1(n1204), .A2(n1346), .ZN(n1343) );
INV_X1 U1066 ( .A(KEYINPUT16), .ZN(n1346) );
NOR2_X1 U1067 ( .A1(n1345), .A2(n1344), .ZN(n1204) );
NOR2_X1 U1068 ( .A1(n1154), .A2(G953), .ZN(n1344) );
INV_X1 U1069 ( .A(G224), .ZN(n1154) );
NAND2_X1 U1070 ( .A1(KEYINPUT16), .A2(n1345), .ZN(n1342) );
XNOR2_X1 U1071 ( .A(n1326), .B(n1108), .ZN(n1345) );
XNOR2_X1 U1072 ( .A(G125), .B(KEYINPUT11), .ZN(n1108) );
NAND2_X1 U1073 ( .A1(n1347), .A2(n1348), .ZN(n1326) );
NAND2_X1 U1074 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
XOR2_X1 U1075 ( .A(n1351), .B(KEYINPUT29), .Z(n1347) );
OR2_X1 U1076 ( .A1(n1350), .A2(n1349), .ZN(n1351) );
XNOR2_X1 U1077 ( .A(n1298), .B(KEYINPUT32), .ZN(n1349) );
XOR2_X1 U1078 ( .A(G128), .B(KEYINPUT15), .Z(n1298) );
NAND2_X1 U1079 ( .A1(n1352), .A2(n1353), .ZN(n1350) );
NAND2_X1 U1080 ( .A1(G143), .A2(n1273), .ZN(n1353) );
XOR2_X1 U1081 ( .A(KEYINPUT47), .B(n1354), .Z(n1352) );
NOR2_X1 U1082 ( .A1(G143), .A2(n1273), .ZN(n1354) );
INV_X1 U1083 ( .A(G146), .ZN(n1273) );
endmodule


