//Key = 1110010011100001001100110111111111001100111110101010100111011111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351;

XNOR2_X1 U749 ( .A(G107), .B(n1038), .ZN(G9) );
NAND3_X1 U750 ( .A1(n1039), .A2(n1040), .A3(KEYINPUT32), .ZN(n1038) );
NOR2_X1 U751 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR4_X1 U752 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
NAND3_X1 U753 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1043) );
NAND2_X1 U754 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND4_X1 U755 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1051) );
NAND3_X1 U756 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NAND2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND2_X1 U758 ( .A1(KEYINPUT56), .A2(n1061), .ZN(n1060) );
NAND2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1054) );
INV_X1 U760 ( .A(KEYINPUT56), .ZN(n1063) );
NAND2_X1 U761 ( .A1(n1058), .A2(n1064), .ZN(n1062) );
NAND2_X1 U762 ( .A1(n1065), .A2(n1066), .ZN(n1053) );
NAND2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND3_X1 U764 ( .A1(n1056), .A2(n1069), .A3(n1070), .ZN(n1068) );
INV_X1 U765 ( .A(n1071), .ZN(n1070) );
NAND2_X1 U766 ( .A1(n1072), .A2(n1073), .ZN(n1069) );
NAND2_X1 U767 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U768 ( .A1(n1058), .A2(n1076), .ZN(n1067) );
NAND2_X1 U769 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
OR3_X1 U770 ( .A1(n1079), .A2(KEYINPUT53), .A3(n1080), .ZN(n1078) );
NAND2_X1 U771 ( .A1(KEYINPUT53), .A2(n1081), .ZN(n1052) );
NAND4_X1 U772 ( .A1(n1058), .A2(n1065), .A3(n1082), .A4(n1083), .ZN(n1081) );
NAND4_X1 U773 ( .A1(n1058), .A2(n1056), .A3(n1065), .A4(n1084), .ZN(n1047) );
NAND2_X1 U774 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U775 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U776 ( .A(n1089), .B(KEYINPUT21), .Z(n1085) );
NOR3_X1 U777 ( .A1(n1090), .A2(n1074), .A3(n1071), .ZN(n1058) );
NOR3_X1 U778 ( .A1(n1045), .A2(G952), .A3(n1091), .ZN(n1041) );
INV_X1 U779 ( .A(n1048), .ZN(n1091) );
NAND4_X1 U780 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1048) );
NOR4_X1 U781 ( .A1(n1096), .A2(n1090), .A3(n1097), .A4(n1098), .ZN(n1095) );
XOR2_X1 U782 ( .A(KEYINPUT38), .B(n1080), .Z(n1098) );
XOR2_X1 U783 ( .A(KEYINPUT35), .B(n1099), .Z(n1097) );
NOR2_X1 U784 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR3_X1 U785 ( .A1(n1083), .A2(n1102), .A3(n1103), .ZN(n1094) );
INV_X1 U786 ( .A(n1079), .ZN(n1083) );
NAND2_X1 U787 ( .A1(n1100), .A2(n1101), .ZN(n1093) );
XOR2_X1 U788 ( .A(n1104), .B(n1105), .Z(G72) );
XOR2_X1 U789 ( .A(n1106), .B(n1107), .Z(n1105) );
NAND2_X1 U790 ( .A1(KEYINPUT18), .A2(n1108), .ZN(n1107) );
NAND2_X1 U791 ( .A1(n1044), .A2(n1109), .ZN(n1108) );
NAND2_X1 U792 ( .A1(n1110), .A2(n1111), .ZN(n1106) );
NAND2_X1 U793 ( .A1(G953), .A2(n1112), .ZN(n1111) );
XOR2_X1 U794 ( .A(n1113), .B(n1114), .Z(n1110) );
XOR2_X1 U795 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U796 ( .A1(KEYINPUT15), .A2(n1117), .ZN(n1115) );
XOR2_X1 U797 ( .A(G134), .B(n1118), .Z(n1117) );
XOR2_X1 U798 ( .A(n1119), .B(n1120), .Z(n1113) );
XOR2_X1 U799 ( .A(G140), .B(G131), .Z(n1120) );
NAND2_X1 U800 ( .A1(G953), .A2(n1121), .ZN(n1104) );
NAND2_X1 U801 ( .A1(G900), .A2(G227), .ZN(n1121) );
NAND2_X1 U802 ( .A1(n1122), .A2(n1123), .ZN(G69) );
NAND2_X1 U803 ( .A1(n1124), .A2(n1109), .ZN(n1123) );
XNOR2_X1 U804 ( .A(n1046), .B(n1125), .ZN(n1124) );
NAND2_X1 U805 ( .A1(n1126), .A2(G953), .ZN(n1122) );
NAND2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U807 ( .A1(n1125), .A2(n1129), .ZN(n1128) );
INV_X1 U808 ( .A(G224), .ZN(n1129) );
NAND2_X1 U809 ( .A1(G224), .A2(n1130), .ZN(n1127) );
NAND2_X1 U810 ( .A1(G898), .A2(n1125), .ZN(n1130) );
NAND2_X1 U811 ( .A1(n1131), .A2(n1132), .ZN(n1125) );
NAND2_X1 U812 ( .A1(G953), .A2(n1133), .ZN(n1132) );
XOR2_X1 U813 ( .A(n1134), .B(n1135), .Z(n1131) );
NOR2_X1 U814 ( .A1(n1136), .A2(n1137), .ZN(G66) );
XOR2_X1 U815 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U816 ( .A1(n1101), .A2(n1140), .ZN(n1139) );
NOR2_X1 U817 ( .A1(n1136), .A2(n1141), .ZN(G63) );
XOR2_X1 U818 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U819 ( .A1(n1144), .A2(n1140), .ZN(n1142) );
INV_X1 U820 ( .A(G478), .ZN(n1144) );
NOR2_X1 U821 ( .A1(n1136), .A2(n1145), .ZN(G60) );
XOR2_X1 U822 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U823 ( .A1(n1148), .A2(n1140), .ZN(n1147) );
INV_X1 U824 ( .A(G475), .ZN(n1148) );
XOR2_X1 U825 ( .A(G104), .B(n1149), .Z(G6) );
NOR3_X1 U826 ( .A1(n1150), .A2(KEYINPUT54), .A3(n1151), .ZN(n1149) );
NOR2_X1 U827 ( .A1(n1136), .A2(n1152), .ZN(G57) );
XOR2_X1 U828 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U829 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U830 ( .A1(n1157), .A2(n1140), .ZN(n1155) );
INV_X1 U831 ( .A(G472), .ZN(n1157) );
XOR2_X1 U832 ( .A(n1158), .B(KEYINPUT0), .Z(n1153) );
NAND3_X1 U833 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1158) );
OR2_X1 U834 ( .A1(n1162), .A2(KEYINPUT31), .ZN(n1161) );
OR3_X1 U835 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1160) );
INV_X1 U836 ( .A(KEYINPUT31), .ZN(n1163) );
NAND2_X1 U837 ( .A1(n1164), .A2(n1165), .ZN(n1159) );
NAND2_X1 U838 ( .A1(KEYINPUT55), .A2(n1162), .ZN(n1164) );
XNOR2_X1 U839 ( .A(n1166), .B(n1167), .ZN(n1162) );
NAND2_X1 U840 ( .A1(KEYINPUT23), .A2(n1168), .ZN(n1166) );
NOR2_X1 U841 ( .A1(n1136), .A2(n1169), .ZN(G54) );
XOR2_X1 U842 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U843 ( .A1(n1172), .A2(n1140), .ZN(n1171) );
INV_X1 U844 ( .A(G469), .ZN(n1172) );
NOR2_X1 U845 ( .A1(n1173), .A2(n1174), .ZN(n1170) );
XOR2_X1 U846 ( .A(n1175), .B(KEYINPUT63), .Z(n1174) );
NAND2_X1 U847 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U848 ( .A(KEYINPUT10), .B(n1178), .Z(n1177) );
NOR2_X1 U849 ( .A1(n1176), .A2(n1179), .ZN(n1173) );
XOR2_X1 U850 ( .A(KEYINPUT8), .B(n1178), .Z(n1179) );
XNOR2_X1 U851 ( .A(n1180), .B(n1181), .ZN(n1178) );
XOR2_X1 U852 ( .A(n1182), .B(n1183), .Z(n1176) );
NOR2_X1 U853 ( .A1(KEYINPUT58), .A2(n1168), .ZN(n1183) );
NOR2_X1 U854 ( .A1(n1109), .A2(G952), .ZN(n1136) );
NOR2_X1 U855 ( .A1(n1184), .A2(n1185), .ZN(G51) );
XOR2_X1 U856 ( .A(n1186), .B(n1187), .Z(n1185) );
XNOR2_X1 U857 ( .A(n1188), .B(n1189), .ZN(n1187) );
XOR2_X1 U858 ( .A(n1190), .B(n1191), .Z(n1186) );
NOR2_X1 U859 ( .A1(n1192), .A2(n1140), .ZN(n1191) );
NAND2_X1 U860 ( .A1(n1193), .A2(n1194), .ZN(n1140) );
OR2_X1 U861 ( .A1(n1044), .A2(n1046), .ZN(n1194) );
NAND4_X1 U862 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1046) );
AND4_X1 U863 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1198) );
NAND2_X1 U864 ( .A1(n1203), .A2(n1204), .ZN(n1197) );
XNOR2_X1 U865 ( .A(KEYINPUT7), .B(n1205), .ZN(n1204) );
NAND2_X1 U866 ( .A1(n1040), .A2(n1206), .ZN(n1195) );
NAND2_X1 U867 ( .A1(n1150), .A2(n1059), .ZN(n1206) );
INV_X1 U868 ( .A(n1151), .ZN(n1040) );
NAND2_X1 U869 ( .A1(n1207), .A2(n1208), .ZN(n1151) );
NAND4_X1 U870 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1044) );
AND4_X1 U871 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1212) );
NOR2_X1 U872 ( .A1(n1217), .A2(n1218), .ZN(n1211) );
NOR3_X1 U873 ( .A1(n1219), .A2(n1150), .A3(n1220), .ZN(n1218) );
XOR2_X1 U874 ( .A(KEYINPUT61), .B(n1203), .Z(n1219) );
XOR2_X1 U875 ( .A(n1221), .B(KEYINPUT52), .Z(n1193) );
NAND2_X1 U876 ( .A1(KEYINPUT5), .A2(G125), .ZN(n1190) );
NOR2_X1 U877 ( .A1(G952), .A2(n1222), .ZN(n1184) );
XOR2_X1 U878 ( .A(KEYINPUT44), .B(G953), .Z(n1222) );
XNOR2_X1 U879 ( .A(G146), .B(n1223), .ZN(G48) );
NAND2_X1 U880 ( .A1(n1224), .A2(n1061), .ZN(n1223) );
XNOR2_X1 U881 ( .A(n1217), .B(n1225), .ZN(G45) );
NAND2_X1 U882 ( .A1(KEYINPUT41), .A2(G143), .ZN(n1225) );
AND4_X1 U883 ( .A1(n1207), .A2(n1203), .A3(n1226), .A4(n1227), .ZN(n1217) );
NOR3_X1 U884 ( .A1(n1092), .A2(n1228), .A3(n1229), .ZN(n1227) );
XOR2_X1 U885 ( .A(n1230), .B(n1209), .Z(G42) );
NAND3_X1 U886 ( .A1(n1050), .A2(n1207), .A3(n1231), .ZN(n1209) );
XNOR2_X1 U887 ( .A(G137), .B(n1215), .ZN(G39) );
NAND3_X1 U888 ( .A1(n1232), .A2(n1050), .A3(n1065), .ZN(n1215) );
INV_X1 U889 ( .A(n1096), .ZN(n1050) );
INV_X1 U890 ( .A(n1220), .ZN(n1232) );
XOR2_X1 U891 ( .A(n1233), .B(n1214), .Z(G36) );
NAND3_X1 U892 ( .A1(n1039), .A2(n1234), .A3(n1235), .ZN(n1214) );
XNOR2_X1 U893 ( .A(G131), .B(n1213), .ZN(G33) );
NAND3_X1 U894 ( .A1(n1235), .A2(n1234), .A3(n1061), .ZN(n1213) );
NOR3_X1 U895 ( .A1(n1096), .A2(n1077), .A3(n1072), .ZN(n1235) );
NAND2_X1 U896 ( .A1(n1088), .A2(n1236), .ZN(n1096) );
XOR2_X1 U897 ( .A(n1237), .B(n1210), .Z(G30) );
NAND2_X1 U898 ( .A1(n1224), .A2(n1039), .ZN(n1210) );
NOR2_X1 U899 ( .A1(n1220), .A2(n1089), .ZN(n1224) );
NAND4_X1 U900 ( .A1(n1074), .A2(n1207), .A3(n1090), .A4(n1234), .ZN(n1220) );
XNOR2_X1 U901 ( .A(G101), .B(n1196), .ZN(G3) );
NAND4_X1 U902 ( .A1(n1065), .A2(n1226), .A3(n1207), .A4(n1238), .ZN(n1196) );
XOR2_X1 U903 ( .A(n1119), .B(n1216), .Z(G27) );
NAND3_X1 U904 ( .A1(n1231), .A2(n1203), .A3(n1056), .ZN(n1216) );
NOR4_X1 U905 ( .A1(n1239), .A2(n1150), .A3(n1090), .A4(n1229), .ZN(n1231) );
INV_X1 U906 ( .A(n1234), .ZN(n1229) );
NAND2_X1 U907 ( .A1(n1071), .A2(n1240), .ZN(n1234) );
NAND4_X1 U908 ( .A1(G953), .A2(G902), .A3(n1241), .A4(n1112), .ZN(n1240) );
INV_X1 U909 ( .A(G900), .ZN(n1112) );
XOR2_X1 U910 ( .A(n1242), .B(n1202), .Z(G24) );
NAND4_X1 U911 ( .A1(n1056), .A2(n1208), .A3(n1243), .A4(n1244), .ZN(n1202) );
AND3_X1 U912 ( .A1(n1075), .A2(n1239), .A3(n1238), .ZN(n1208) );
XOR2_X1 U913 ( .A(n1245), .B(n1201), .Z(G21) );
NAND3_X1 U914 ( .A1(n1056), .A2(n1090), .A3(n1246), .ZN(n1201) );
XOR2_X1 U915 ( .A(G116), .B(n1247), .Z(G18) );
NOR2_X1 U916 ( .A1(n1089), .A2(n1205), .ZN(n1247) );
NAND4_X1 U917 ( .A1(n1056), .A2(n1226), .A3(n1039), .A4(n1248), .ZN(n1205) );
INV_X1 U918 ( .A(n1059), .ZN(n1039) );
NAND2_X1 U919 ( .A1(n1228), .A2(n1243), .ZN(n1059) );
INV_X1 U920 ( .A(n1203), .ZN(n1089) );
XNOR2_X1 U921 ( .A(G113), .B(n1200), .ZN(G15) );
NAND3_X1 U922 ( .A1(n1226), .A2(n1238), .A3(n1064), .ZN(n1200) );
AND2_X1 U923 ( .A1(n1056), .A2(n1061), .ZN(n1064) );
INV_X1 U924 ( .A(n1150), .ZN(n1061) );
NAND2_X1 U925 ( .A1(n1092), .A2(n1244), .ZN(n1150) );
INV_X1 U926 ( .A(n1243), .ZN(n1092) );
AND2_X1 U927 ( .A1(n1082), .A2(n1249), .ZN(n1056) );
INV_X1 U928 ( .A(n1072), .ZN(n1226) );
NAND2_X1 U929 ( .A1(n1090), .A2(n1239), .ZN(n1072) );
INV_X1 U930 ( .A(n1074), .ZN(n1239) );
INV_X1 U931 ( .A(n1075), .ZN(n1090) );
XOR2_X1 U932 ( .A(n1250), .B(n1199), .Z(G12) );
NAND3_X1 U933 ( .A1(n1075), .A2(n1207), .A3(n1246), .ZN(n1199) );
AND3_X1 U934 ( .A1(n1074), .A2(n1238), .A3(n1065), .ZN(n1246) );
NOR2_X1 U935 ( .A1(n1244), .A2(n1243), .ZN(n1065) );
XOR2_X1 U936 ( .A(n1251), .B(n1252), .Z(n1243) );
XOR2_X1 U937 ( .A(KEYINPUT37), .B(G478), .Z(n1252) );
OR2_X1 U938 ( .A1(n1143), .A2(G902), .ZN(n1251) );
XNOR2_X1 U939 ( .A(n1253), .B(n1254), .ZN(n1143) );
XOR2_X1 U940 ( .A(G107), .B(n1255), .Z(n1254) );
XOR2_X1 U941 ( .A(KEYINPUT20), .B(G134), .Z(n1255) );
XNOR2_X1 U942 ( .A(n1256), .B(n1257), .ZN(n1253) );
XOR2_X1 U943 ( .A(n1258), .B(n1259), .Z(n1257) );
NAND3_X1 U944 ( .A1(G217), .A2(n1109), .A3(G234), .ZN(n1259) );
NAND2_X1 U945 ( .A1(n1260), .A2(n1261), .ZN(n1258) );
NAND2_X1 U946 ( .A1(G116), .A2(n1242), .ZN(n1261) );
XOR2_X1 U947 ( .A(n1262), .B(KEYINPUT17), .Z(n1260) );
OR2_X1 U948 ( .A1(n1242), .A2(G116), .ZN(n1262) );
INV_X1 U949 ( .A(n1228), .ZN(n1244) );
NOR2_X1 U950 ( .A1(n1263), .A2(n1103), .ZN(n1228) );
NOR3_X1 U951 ( .A1(G475), .A2(G902), .A3(n1146), .ZN(n1103) );
XOR2_X1 U952 ( .A(n1102), .B(KEYINPUT16), .Z(n1263) );
AND2_X1 U953 ( .A1(G475), .A2(n1264), .ZN(n1102) );
NAND2_X1 U954 ( .A1(n1265), .A2(n1221), .ZN(n1264) );
INV_X1 U955 ( .A(n1146), .ZN(n1265) );
XOR2_X1 U956 ( .A(n1266), .B(n1267), .Z(n1146) );
XOR2_X1 U957 ( .A(G104), .B(n1268), .Z(n1267) );
NOR2_X1 U958 ( .A1(KEYINPUT24), .A2(n1269), .ZN(n1268) );
XOR2_X1 U959 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U960 ( .A(n1272), .B(n1273), .Z(n1271) );
AND3_X1 U961 ( .A1(G214), .A2(n1109), .A3(n1274), .ZN(n1273) );
NOR2_X1 U962 ( .A1(KEYINPUT13), .A2(n1275), .ZN(n1272) );
XOR2_X1 U963 ( .A(n1276), .B(n1277), .Z(n1275) );
NOR2_X1 U964 ( .A1(KEYINPUT12), .A2(n1230), .ZN(n1277) );
XOR2_X1 U965 ( .A(G131), .B(n1278), .Z(n1270) );
XOR2_X1 U966 ( .A(KEYINPUT28), .B(G143), .Z(n1278) );
XOR2_X1 U967 ( .A(G113), .B(n1242), .Z(n1266) );
INV_X1 U968 ( .A(G122), .ZN(n1242) );
AND2_X1 U969 ( .A1(n1203), .A2(n1248), .ZN(n1238) );
NAND2_X1 U970 ( .A1(n1071), .A2(n1279), .ZN(n1248) );
NAND4_X1 U971 ( .A1(G953), .A2(G902), .A3(n1241), .A4(n1133), .ZN(n1279) );
INV_X1 U972 ( .A(G898), .ZN(n1133) );
NAND3_X1 U973 ( .A1(n1280), .A2(n1241), .A3(G952), .ZN(n1071) );
NAND2_X1 U974 ( .A1(G234), .A2(G237), .ZN(n1241) );
INV_X1 U975 ( .A(n1045), .ZN(n1280) );
XOR2_X1 U976 ( .A(n1109), .B(KEYINPUT2), .Z(n1045) );
NOR2_X1 U977 ( .A1(n1088), .A2(n1087), .ZN(n1203) );
INV_X1 U978 ( .A(n1236), .ZN(n1087) );
NAND2_X1 U979 ( .A1(G214), .A2(n1281), .ZN(n1236) );
XNOR2_X1 U980 ( .A(n1282), .B(n1192), .ZN(n1088) );
NAND2_X1 U981 ( .A1(G210), .A2(n1281), .ZN(n1192) );
NAND2_X1 U982 ( .A1(n1283), .A2(n1221), .ZN(n1281) );
NAND2_X1 U983 ( .A1(n1284), .A2(n1221), .ZN(n1282) );
XOR2_X1 U984 ( .A(n1285), .B(n1189), .Z(n1284) );
XNOR2_X1 U985 ( .A(n1286), .B(n1135), .ZN(n1189) );
XOR2_X1 U986 ( .A(G110), .B(G122), .Z(n1135) );
NAND2_X1 U987 ( .A1(KEYINPUT33), .A2(n1134), .ZN(n1286) );
XOR2_X1 U988 ( .A(n1287), .B(n1288), .Z(n1134) );
XOR2_X1 U989 ( .A(G116), .B(n1289), .Z(n1288) );
XOR2_X1 U990 ( .A(KEYINPUT29), .B(G119), .Z(n1289) );
XOR2_X1 U991 ( .A(n1290), .B(n1291), .Z(n1287) );
NAND2_X1 U992 ( .A1(KEYINPUT59), .A2(n1292), .ZN(n1290) );
NAND2_X1 U993 ( .A1(KEYINPUT36), .A2(n1293), .ZN(n1285) );
XOR2_X1 U994 ( .A(G125), .B(n1188), .Z(n1293) );
XNOR2_X1 U995 ( .A(n1294), .B(n1167), .ZN(n1188) );
NAND2_X1 U996 ( .A1(G224), .A2(n1109), .ZN(n1294) );
XNOR2_X1 U997 ( .A(n1295), .B(n1101), .ZN(n1074) );
NAND2_X1 U998 ( .A1(G217), .A2(n1296), .ZN(n1101) );
XNOR2_X1 U999 ( .A(n1100), .B(KEYINPUT9), .ZN(n1295) );
NOR2_X1 U1000 ( .A1(n1138), .A2(G902), .ZN(n1100) );
XOR2_X1 U1001 ( .A(n1297), .B(n1298), .Z(n1138) );
XOR2_X1 U1002 ( .A(n1299), .B(n1300), .Z(n1298) );
NAND2_X1 U1003 ( .A1(KEYINPUT19), .A2(n1301), .ZN(n1300) );
XOR2_X1 U1004 ( .A(n1245), .B(n1302), .Z(n1301) );
NAND2_X1 U1005 ( .A1(KEYINPUT30), .A2(n1237), .ZN(n1302) );
INV_X1 U1006 ( .A(G119), .ZN(n1245) );
NAND3_X1 U1007 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(n1299) );
NAND2_X1 U1008 ( .A1(n1118), .A2(n1306), .ZN(n1305) );
OR3_X1 U1009 ( .A1(n1306), .A2(n1118), .A3(KEYINPUT6), .ZN(n1304) );
NAND2_X1 U1010 ( .A1(KEYINPUT22), .A2(n1307), .ZN(n1306) );
INV_X1 U1011 ( .A(n1308), .ZN(n1307) );
NAND2_X1 U1012 ( .A1(KEYINPUT6), .A2(n1308), .ZN(n1303) );
NAND3_X1 U1013 ( .A1(G234), .A2(n1109), .A3(G221), .ZN(n1308) );
XOR2_X1 U1014 ( .A(n1276), .B(n1181), .Z(n1297) );
XOR2_X1 U1015 ( .A(G110), .B(G140), .Z(n1181) );
XOR2_X1 U1016 ( .A(G146), .B(n1119), .Z(n1276) );
INV_X1 U1017 ( .A(G125), .ZN(n1119) );
INV_X1 U1018 ( .A(n1077), .ZN(n1207) );
NAND2_X1 U1019 ( .A1(n1249), .A2(n1080), .ZN(n1077) );
INV_X1 U1020 ( .A(n1082), .ZN(n1080) );
XOR2_X1 U1021 ( .A(n1309), .B(G469), .Z(n1082) );
NAND2_X1 U1022 ( .A1(n1310), .A2(n1221), .ZN(n1309) );
XOR2_X1 U1023 ( .A(n1311), .B(n1312), .Z(n1310) );
NOR2_X1 U1024 ( .A1(KEYINPUT3), .A2(n1180), .ZN(n1312) );
NAND2_X1 U1025 ( .A1(G227), .A2(n1109), .ZN(n1180) );
XOR2_X1 U1026 ( .A(n1313), .B(n1314), .Z(n1311) );
NOR2_X1 U1027 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NOR2_X1 U1028 ( .A1(n1317), .A2(G110), .ZN(n1316) );
NOR2_X1 U1029 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NOR2_X1 U1030 ( .A1(G140), .A2(n1320), .ZN(n1318) );
NOR2_X1 U1031 ( .A1(n1321), .A2(n1230), .ZN(n1315) );
INV_X1 U1032 ( .A(G140), .ZN(n1230) );
NOR2_X1 U1033 ( .A1(n1322), .A2(n1320), .ZN(n1321) );
INV_X1 U1034 ( .A(KEYINPUT60), .ZN(n1320) );
NOR2_X1 U1035 ( .A1(n1250), .A2(n1319), .ZN(n1322) );
INV_X1 U1036 ( .A(KEYINPUT1), .ZN(n1319) );
NAND2_X1 U1037 ( .A1(n1323), .A2(KEYINPUT57), .ZN(n1313) );
XOR2_X1 U1038 ( .A(n1182), .B(n1324), .Z(n1323) );
XOR2_X1 U1039 ( .A(KEYINPUT50), .B(n1325), .Z(n1324) );
XOR2_X1 U1040 ( .A(n1326), .B(n1327), .Z(n1182) );
XOR2_X1 U1041 ( .A(KEYINPUT51), .B(KEYINPUT34), .Z(n1327) );
XNOR2_X1 U1042 ( .A(n1116), .B(n1291), .ZN(n1326) );
XOR2_X1 U1043 ( .A(G101), .B(n1328), .Z(n1291) );
XOR2_X1 U1044 ( .A(G107), .B(G104), .Z(n1328) );
XNOR2_X1 U1045 ( .A(n1329), .B(n1167), .ZN(n1116) );
XNOR2_X1 U1046 ( .A(KEYINPUT47), .B(KEYINPUT25), .ZN(n1329) );
XOR2_X1 U1047 ( .A(n1079), .B(KEYINPUT49), .Z(n1249) );
NAND2_X1 U1048 ( .A1(G221), .A2(n1296), .ZN(n1079) );
NAND2_X1 U1049 ( .A1(G234), .A2(n1221), .ZN(n1296) );
XOR2_X1 U1050 ( .A(n1330), .B(G472), .Z(n1075) );
NAND2_X1 U1051 ( .A1(n1331), .A2(n1221), .ZN(n1330) );
INV_X1 U1052 ( .A(G902), .ZN(n1221) );
XOR2_X1 U1053 ( .A(n1332), .B(n1333), .Z(n1331) );
XNOR2_X1 U1054 ( .A(KEYINPUT11), .B(n1165), .ZN(n1333) );
NAND2_X1 U1055 ( .A1(n1334), .A2(n1335), .ZN(n1165) );
NAND2_X1 U1056 ( .A1(n1292), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1057 ( .A(n1337), .B(KEYINPUT4), .Z(n1334) );
OR2_X1 U1058 ( .A1(n1336), .A2(n1292), .ZN(n1337) );
XNOR2_X1 U1059 ( .A(G113), .B(KEYINPUT39), .ZN(n1292) );
XNOR2_X1 U1060 ( .A(n1338), .B(n1339), .ZN(n1336) );
XOR2_X1 U1061 ( .A(KEYINPUT27), .B(G119), .Z(n1339) );
NAND2_X1 U1062 ( .A1(KEYINPUT48), .A2(G116), .ZN(n1338) );
XOR2_X1 U1063 ( .A(n1340), .B(n1156), .Z(n1332) );
XNOR2_X1 U1064 ( .A(n1341), .B(G101), .ZN(n1156) );
NAND3_X1 U1065 ( .A1(n1342), .A2(n1109), .A3(G210), .ZN(n1341) );
INV_X1 U1066 ( .A(G953), .ZN(n1109) );
XOR2_X1 U1067 ( .A(KEYINPUT14), .B(n1274), .Z(n1342) );
XNOR2_X1 U1068 ( .A(n1283), .B(KEYINPUT26), .ZN(n1274) );
INV_X1 U1069 ( .A(G237), .ZN(n1283) );
NAND4_X1 U1070 ( .A1(KEYINPUT46), .A2(n1343), .A3(n1344), .A4(n1345), .ZN(n1340) );
NAND3_X1 U1071 ( .A1(n1346), .A2(n1347), .A3(KEYINPUT42), .ZN(n1345) );
INV_X1 U1072 ( .A(n1348), .ZN(n1346) );
OR2_X1 U1073 ( .A1(n1325), .A2(KEYINPUT42), .ZN(n1344) );
NAND2_X1 U1074 ( .A1(n1167), .A2(n1348), .ZN(n1343) );
NAND2_X1 U1075 ( .A1(KEYINPUT40), .A2(n1325), .ZN(n1348) );
INV_X1 U1076 ( .A(n1168), .ZN(n1325) );
XOR2_X1 U1077 ( .A(n1349), .B(n1350), .Z(n1168) );
XOR2_X1 U1078 ( .A(KEYINPUT62), .B(G131), .Z(n1350) );
XOR2_X1 U1079 ( .A(n1351), .B(n1118), .Z(n1349) );
XOR2_X1 U1080 ( .A(G137), .B(KEYINPUT45), .Z(n1118) );
NAND2_X1 U1081 ( .A1(KEYINPUT43), .A2(n1233), .ZN(n1351) );
INV_X1 U1082 ( .A(G134), .ZN(n1233) );
INV_X1 U1083 ( .A(n1347), .ZN(n1167) );
XNOR2_X1 U1084 ( .A(G146), .B(n1256), .ZN(n1347) );
XNOR2_X1 U1085 ( .A(n1237), .B(G143), .ZN(n1256) );
INV_X1 U1086 ( .A(G128), .ZN(n1237) );
INV_X1 U1087 ( .A(G110), .ZN(n1250) );
endmodule


