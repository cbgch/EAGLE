//Key = 0010100010001011100111000110101100010100100011101100110101101101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359;

XOR2_X1 U746 ( .A(n1023), .B(G107), .Z(G9) );
NAND2_X1 U747 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND2_X1 U748 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
INV_X1 U749 ( .A(KEYINPUT38), .ZN(n1027) );
NAND3_X1 U750 ( .A1(n1028), .A2(n1029), .A3(KEYINPUT38), .ZN(n1024) );
NOR2_X1 U751 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR3_X1 U752 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NAND3_X1 U753 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1032) );
NAND2_X1 U754 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U755 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND4_X1 U756 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1041) );
NAND2_X1 U757 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U758 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U759 ( .A1(n1050), .A2(n1051), .ZN(n1040) );
NAND2_X1 U760 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND3_X1 U761 ( .A1(n1044), .A2(n1054), .A3(n1042), .ZN(n1053) );
OR2_X1 U762 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U763 ( .A1(n1043), .A2(n1057), .ZN(n1052) );
NAND2_X1 U764 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U765 ( .A1(n1044), .A2(n1060), .ZN(n1059) );
NAND2_X1 U766 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U767 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U768 ( .A1(n1042), .A2(n1065), .ZN(n1058) );
NAND2_X1 U769 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
INV_X1 U770 ( .A(n1068), .ZN(n1038) );
NOR3_X1 U771 ( .A1(n1069), .A2(G953), .A3(G952), .ZN(n1030) );
INV_X1 U772 ( .A(n1035), .ZN(n1069) );
NAND4_X1 U773 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1035) );
NOR4_X1 U774 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1073) );
XOR2_X1 U775 ( .A(n1078), .B(n1079), .Z(n1077) );
XOR2_X1 U776 ( .A(KEYINPUT20), .B(n1080), .Z(n1079) );
NOR2_X1 U777 ( .A1(KEYINPUT43), .A2(n1081), .ZN(n1078) );
XNOR2_X1 U778 ( .A(G478), .B(KEYINPUT63), .ZN(n1081) );
AND2_X1 U779 ( .A1(n1067), .A2(KEYINPUT6), .ZN(n1075) );
INV_X1 U780 ( .A(n1082), .ZN(n1067) );
NOR2_X1 U781 ( .A1(KEYINPUT6), .A2(n1044), .ZN(n1074) );
NOR2_X1 U782 ( .A1(n1063), .A2(n1083), .ZN(n1072) );
NOR2_X1 U783 ( .A1(G469), .A2(n1084), .ZN(n1083) );
XOR2_X1 U784 ( .A(n1085), .B(n1086), .Z(n1071) );
XNOR2_X1 U785 ( .A(n1087), .B(KEYINPUT24), .ZN(n1086) );
NAND2_X1 U786 ( .A1(KEYINPUT53), .A2(n1088), .ZN(n1087) );
XOR2_X1 U787 ( .A(KEYINPUT31), .B(n1089), .Z(n1070) );
AND2_X1 U788 ( .A1(n1084), .A2(G469), .ZN(n1089) );
XNOR2_X1 U789 ( .A(n1090), .B(KEYINPUT4), .ZN(n1084) );
XOR2_X1 U790 ( .A(n1091), .B(n1092), .Z(G72) );
NOR2_X1 U791 ( .A1(n1093), .A2(n1036), .ZN(n1092) );
AND2_X1 U792 ( .A1(G227), .A2(G900), .ZN(n1093) );
NAND2_X1 U793 ( .A1(n1094), .A2(n1095), .ZN(n1091) );
NAND2_X1 U794 ( .A1(n1096), .A2(n1036), .ZN(n1095) );
XOR2_X1 U795 ( .A(n1034), .B(n1097), .Z(n1096) );
NAND3_X1 U796 ( .A1(n1098), .A2(n1097), .A3(G953), .ZN(n1094) );
XOR2_X1 U797 ( .A(n1099), .B(n1100), .Z(n1097) );
XOR2_X1 U798 ( .A(n1101), .B(n1102), .Z(n1100) );
XNOR2_X1 U799 ( .A(KEYINPUT39), .B(n1103), .ZN(n1102) );
NOR2_X1 U800 ( .A1(KEYINPUT10), .A2(n1104), .ZN(n1101) );
XNOR2_X1 U801 ( .A(n1105), .B(n1106), .ZN(n1099) );
XNOR2_X1 U802 ( .A(G900), .B(KEYINPUT30), .ZN(n1098) );
XOR2_X1 U803 ( .A(n1107), .B(n1108), .Z(G69) );
NOR2_X1 U804 ( .A1(n1109), .A2(n1036), .ZN(n1108) );
NOR2_X1 U805 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U806 ( .A1(n1112), .A2(n1113), .ZN(n1107) );
NAND2_X1 U807 ( .A1(n1114), .A2(n1036), .ZN(n1113) );
XOR2_X1 U808 ( .A(n1033), .B(n1115), .Z(n1114) );
NAND3_X1 U809 ( .A1(G898), .A2(n1115), .A3(G953), .ZN(n1112) );
XOR2_X1 U810 ( .A(n1116), .B(n1117), .Z(n1115) );
XNOR2_X1 U811 ( .A(KEYINPUT32), .B(n1118), .ZN(n1117) );
XNOR2_X1 U812 ( .A(n1119), .B(n1120), .ZN(n1116) );
NOR2_X1 U813 ( .A1(n1121), .A2(n1122), .ZN(G66) );
XOR2_X1 U814 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U815 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NOR2_X1 U816 ( .A1(n1121), .A2(n1127), .ZN(G63) );
NOR3_X1 U817 ( .A1(n1080), .A2(n1128), .A3(n1129), .ZN(n1127) );
AND3_X1 U818 ( .A1(n1130), .A2(G478), .A3(n1131), .ZN(n1129) );
NOR2_X1 U819 ( .A1(n1132), .A2(n1130), .ZN(n1128) );
NOR2_X1 U820 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U821 ( .A1(n1033), .A2(n1034), .ZN(n1133) );
NOR2_X1 U822 ( .A1(n1121), .A2(n1135), .ZN(G60) );
NOR3_X1 U823 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
AND2_X1 U824 ( .A1(n1139), .A2(KEYINPUT54), .ZN(n1138) );
NOR3_X1 U825 ( .A1(KEYINPUT54), .A2(n1140), .A3(n1139), .ZN(n1137) );
AND3_X1 U826 ( .A1(KEYINPUT21), .A2(G475), .A3(n1131), .ZN(n1140) );
NOR3_X1 U827 ( .A1(n1126), .A2(n1141), .A3(n1142), .ZN(n1136) );
NOR2_X1 U828 ( .A1(n1143), .A2(KEYINPUT54), .ZN(n1141) );
AND2_X1 U829 ( .A1(n1139), .A2(KEYINPUT21), .ZN(n1143) );
XNOR2_X1 U830 ( .A(n1144), .B(n1145), .ZN(G6) );
NAND2_X1 U831 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
OR2_X1 U832 ( .A1(n1148), .A2(KEYINPUT27), .ZN(n1147) );
NAND3_X1 U833 ( .A1(n1149), .A2(n1150), .A3(KEYINPUT27), .ZN(n1146) );
NOR2_X1 U834 ( .A1(n1121), .A2(n1151), .ZN(G57) );
XOR2_X1 U835 ( .A(n1152), .B(n1153), .Z(n1151) );
XNOR2_X1 U836 ( .A(G101), .B(n1154), .ZN(n1153) );
NAND2_X1 U837 ( .A1(n1155), .A2(n1156), .ZN(n1152) );
NAND2_X1 U838 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XOR2_X1 U839 ( .A(n1159), .B(KEYINPUT42), .Z(n1155) );
OR2_X1 U840 ( .A1(n1158), .A2(n1157), .ZN(n1159) );
NAND2_X1 U841 ( .A1(n1131), .A2(G472), .ZN(n1157) );
NAND2_X1 U842 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
NAND2_X1 U843 ( .A1(n1118), .A2(n1162), .ZN(n1161) );
XOR2_X1 U844 ( .A(n1163), .B(KEYINPUT41), .Z(n1160) );
NAND2_X1 U845 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NOR2_X1 U846 ( .A1(n1121), .A2(n1166), .ZN(G54) );
XOR2_X1 U847 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U848 ( .A(n1169), .B(n1170), .Z(n1168) );
AND2_X1 U849 ( .A1(G469), .A2(n1131), .ZN(n1170) );
INV_X1 U850 ( .A(n1126), .ZN(n1131) );
NAND2_X1 U851 ( .A1(KEYINPUT49), .A2(n1171), .ZN(n1169) );
XOR2_X1 U852 ( .A(n1172), .B(n1173), .Z(n1171) );
NAND2_X1 U853 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XOR2_X1 U854 ( .A(KEYINPUT62), .B(KEYINPUT2), .Z(n1175) );
INV_X1 U855 ( .A(n1176), .ZN(n1174) );
NAND3_X1 U856 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1172) );
NAND2_X1 U857 ( .A1(G110), .A2(n1180), .ZN(n1179) );
OR3_X1 U858 ( .A1(n1180), .A2(G110), .A3(n1181), .ZN(n1178) );
NAND2_X1 U859 ( .A1(n1182), .A2(n1183), .ZN(n1180) );
XOR2_X1 U860 ( .A(KEYINPUT47), .B(KEYINPUT44), .Z(n1182) );
NAND2_X1 U861 ( .A1(G140), .A2(n1181), .ZN(n1177) );
INV_X1 U862 ( .A(KEYINPUT45), .ZN(n1181) );
NOR2_X1 U863 ( .A1(n1121), .A2(n1184), .ZN(G51) );
XOR2_X1 U864 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U865 ( .A(KEYINPUT23), .B(n1187), .Z(n1186) );
NOR2_X1 U866 ( .A1(n1188), .A2(n1126), .ZN(n1187) );
NAND2_X1 U867 ( .A1(G902), .A2(n1189), .ZN(n1126) );
OR2_X1 U868 ( .A1(n1034), .A2(n1033), .ZN(n1189) );
NAND4_X1 U869 ( .A1(n1148), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1033) );
NOR4_X1 U870 ( .A1(n1026), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1192) );
AND2_X1 U871 ( .A1(n1028), .A2(n1196), .ZN(n1026) );
AND4_X1 U872 ( .A1(n1056), .A2(n1044), .A3(n1149), .A4(n1197), .ZN(n1028) );
AND2_X1 U873 ( .A1(n1198), .A2(n1199), .ZN(n1191) );
NAND2_X1 U874 ( .A1(n1200), .A2(n1149), .ZN(n1148) );
INV_X1 U875 ( .A(n1150), .ZN(n1200) );
NAND4_X1 U876 ( .A1(n1055), .A2(n1044), .A3(n1197), .A4(n1196), .ZN(n1150) );
NAND4_X1 U877 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1034) );
NOR4_X1 U878 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
AND2_X1 U879 ( .A1(n1209), .A2(n1210), .ZN(n1203) );
NAND2_X1 U880 ( .A1(n1211), .A2(n1212), .ZN(n1201) );
XOR2_X1 U881 ( .A(n1213), .B(KEYINPUT15), .Z(n1211) );
NOR2_X1 U882 ( .A1(n1036), .A2(G952), .ZN(n1121) );
XNOR2_X1 U883 ( .A(G146), .B(n1202), .ZN(G48) );
NAND3_X1 U884 ( .A1(n1055), .A2(n1214), .A3(n1215), .ZN(n1202) );
NAND2_X1 U885 ( .A1(n1216), .A2(n1217), .ZN(G45) );
NAND2_X1 U886 ( .A1(G143), .A2(n1210), .ZN(n1217) );
XOR2_X1 U887 ( .A(KEYINPUT40), .B(n1218), .Z(n1216) );
NOR2_X1 U888 ( .A1(G143), .A2(n1210), .ZN(n1218) );
NAND4_X1 U889 ( .A1(n1215), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1210) );
NOR3_X1 U890 ( .A1(n1046), .A2(n1222), .A3(n1061), .ZN(n1215) );
NAND2_X1 U891 ( .A1(n1223), .A2(n1224), .ZN(G42) );
NAND2_X1 U892 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
NAND2_X1 U893 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
OR2_X1 U894 ( .A1(KEYINPUT34), .A2(KEYINPUT46), .ZN(n1228) );
NAND3_X1 U895 ( .A1(n1229), .A2(n1230), .A3(KEYINPUT46), .ZN(n1223) );
NAND2_X1 U896 ( .A1(n1227), .A2(n1231), .ZN(n1230) );
OR2_X1 U897 ( .A1(n1225), .A2(KEYINPUT34), .ZN(n1231) );
INV_X1 U898 ( .A(n1209), .ZN(n1225) );
NAND3_X1 U899 ( .A1(n1055), .A2(n1232), .A3(n1082), .ZN(n1209) );
OR2_X1 U900 ( .A1(n1227), .A2(KEYINPUT34), .ZN(n1229) );
XOR2_X1 U901 ( .A(G140), .B(KEYINPUT11), .Z(n1227) );
XNOR2_X1 U902 ( .A(G137), .B(n1233), .ZN(G39) );
NAND2_X1 U903 ( .A1(KEYINPUT28), .A2(n1208), .ZN(n1233) );
AND3_X1 U904 ( .A1(n1232), .A2(n1214), .A3(n1043), .ZN(n1208) );
XOR2_X1 U905 ( .A(G134), .B(n1207), .Z(G36) );
AND3_X1 U906 ( .A1(n1219), .A2(n1056), .A3(n1232), .ZN(n1207) );
XOR2_X1 U907 ( .A(n1206), .B(n1234), .Z(G33) );
NOR2_X1 U908 ( .A1(KEYINPUT56), .A2(n1103), .ZN(n1234) );
AND3_X1 U909 ( .A1(n1232), .A2(n1219), .A3(n1055), .ZN(n1206) );
NOR3_X1 U910 ( .A1(n1061), .A2(n1222), .A3(n1076), .ZN(n1232) );
INV_X1 U911 ( .A(n1050), .ZN(n1076) );
NOR2_X1 U912 ( .A1(n1235), .A2(n1048), .ZN(n1050) );
INV_X1 U913 ( .A(n1236), .ZN(n1222) );
XOR2_X1 U914 ( .A(G128), .B(n1205), .Z(G30) );
AND4_X1 U915 ( .A1(n1214), .A2(n1056), .A3(n1237), .A4(n1212), .ZN(n1205) );
AND2_X1 U916 ( .A1(n1236), .A2(n1197), .ZN(n1237) );
XNOR2_X1 U917 ( .A(n1238), .B(n1239), .ZN(G3) );
NAND2_X1 U918 ( .A1(n1240), .A2(n1241), .ZN(n1238) );
NAND2_X1 U919 ( .A1(n1193), .A2(n1242), .ZN(n1241) );
INV_X1 U920 ( .A(KEYINPUT7), .ZN(n1242) );
AND2_X1 U921 ( .A1(n1243), .A2(n1219), .ZN(n1193) );
NAND3_X1 U922 ( .A1(n1243), .A2(n1066), .A3(KEYINPUT7), .ZN(n1240) );
XOR2_X1 U923 ( .A(G125), .B(n1244), .Z(G27) );
NOR2_X1 U924 ( .A1(n1046), .A2(n1213), .ZN(n1244) );
NAND4_X1 U925 ( .A1(n1042), .A2(n1082), .A3(n1055), .A4(n1236), .ZN(n1213) );
NAND2_X1 U926 ( .A1(n1068), .A2(n1245), .ZN(n1236) );
NAND4_X1 U927 ( .A1(G953), .A2(G902), .A3(n1246), .A4(n1247), .ZN(n1245) );
INV_X1 U928 ( .A(G900), .ZN(n1247) );
INV_X1 U929 ( .A(n1248), .ZN(n1055) );
INV_X1 U930 ( .A(n1249), .ZN(n1042) );
XNOR2_X1 U931 ( .A(G122), .B(n1190), .ZN(G24) );
NAND4_X1 U932 ( .A1(n1250), .A2(n1044), .A3(n1220), .A4(n1221), .ZN(n1190) );
NOR2_X1 U933 ( .A1(n1251), .A2(n1252), .ZN(n1044) );
XOR2_X1 U934 ( .A(n1199), .B(n1253), .Z(G21) );
XNOR2_X1 U935 ( .A(G119), .B(KEYINPUT36), .ZN(n1253) );
NAND3_X1 U936 ( .A1(n1043), .A2(n1214), .A3(n1250), .ZN(n1199) );
AND2_X1 U937 ( .A1(n1254), .A2(n1251), .ZN(n1214) );
XNOR2_X1 U938 ( .A(KEYINPUT33), .B(n1255), .ZN(n1254) );
XNOR2_X1 U939 ( .A(G116), .B(n1198), .ZN(G18) );
NAND3_X1 U940 ( .A1(n1219), .A2(n1056), .A3(n1250), .ZN(n1198) );
NOR3_X1 U941 ( .A1(n1046), .A2(n1029), .A3(n1249), .ZN(n1250) );
INV_X1 U942 ( .A(n1196), .ZN(n1029) );
INV_X1 U943 ( .A(n1212), .ZN(n1046) );
NOR2_X1 U944 ( .A1(n1256), .A2(n1257), .ZN(n1056) );
XOR2_X1 U945 ( .A(G113), .B(n1195), .Z(G15) );
AND4_X1 U946 ( .A1(n1149), .A2(n1196), .A3(n1219), .A4(n1258), .ZN(n1195) );
NOR2_X1 U947 ( .A1(n1248), .A2(n1249), .ZN(n1258) );
NAND2_X1 U948 ( .A1(n1064), .A2(n1259), .ZN(n1249) );
NAND2_X1 U949 ( .A1(n1221), .A2(n1256), .ZN(n1248) );
XNOR2_X1 U950 ( .A(n1257), .B(KEYINPUT25), .ZN(n1221) );
INV_X1 U951 ( .A(n1066), .ZN(n1219) );
NAND2_X1 U952 ( .A1(n1255), .A2(n1251), .ZN(n1066) );
XOR2_X1 U953 ( .A(G110), .B(n1194), .Z(G12) );
AND2_X1 U954 ( .A1(n1243), .A2(n1082), .ZN(n1194) );
NOR2_X1 U955 ( .A1(n1251), .A2(n1255), .ZN(n1082) );
INV_X1 U956 ( .A(n1252), .ZN(n1255) );
XOR2_X1 U957 ( .A(n1260), .B(n1125), .Z(n1252) );
NAND2_X1 U958 ( .A1(G217), .A2(n1261), .ZN(n1125) );
OR2_X1 U959 ( .A1(n1124), .A2(G902), .ZN(n1260) );
XNOR2_X1 U960 ( .A(n1262), .B(n1263), .ZN(n1124) );
XOR2_X1 U961 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U962 ( .A(G119), .B(G110), .Z(n1265) );
XOR2_X1 U963 ( .A(KEYINPUT19), .B(G137), .Z(n1264) );
XNOR2_X1 U964 ( .A(n1266), .B(n1104), .ZN(n1262) );
XNOR2_X1 U965 ( .A(G125), .B(G140), .ZN(n1104) );
XOR2_X1 U966 ( .A(n1267), .B(n1268), .Z(n1266) );
NAND2_X1 U967 ( .A1(G221), .A2(n1269), .ZN(n1267) );
XNOR2_X1 U968 ( .A(n1270), .B(G472), .ZN(n1251) );
NAND2_X1 U969 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XOR2_X1 U970 ( .A(n1273), .B(n1274), .Z(n1271) );
XNOR2_X1 U971 ( .A(n1164), .B(n1165), .ZN(n1274) );
INV_X1 U972 ( .A(n1162), .ZN(n1164) );
XOR2_X1 U973 ( .A(n1275), .B(n1276), .Z(n1273) );
NOR2_X1 U974 ( .A1(KEYINPUT29), .A2(n1154), .ZN(n1276) );
NAND3_X1 U975 ( .A1(n1277), .A2(n1036), .A3(G210), .ZN(n1154) );
XNOR2_X1 U976 ( .A(G101), .B(KEYINPUT1), .ZN(n1275) );
AND4_X1 U977 ( .A1(n1149), .A2(n1043), .A3(n1197), .A4(n1196), .ZN(n1243) );
NAND2_X1 U978 ( .A1(n1278), .A2(n1279), .ZN(n1196) );
NAND4_X1 U979 ( .A1(G953), .A2(G902), .A3(n1246), .A4(n1111), .ZN(n1279) );
INV_X1 U980 ( .A(G898), .ZN(n1111) );
XNOR2_X1 U981 ( .A(KEYINPUT55), .B(n1068), .ZN(n1278) );
NAND3_X1 U982 ( .A1(n1246), .A2(n1036), .A3(G952), .ZN(n1068) );
NAND2_X1 U983 ( .A1(G237), .A2(G234), .ZN(n1246) );
XNOR2_X1 U984 ( .A(n1061), .B(KEYINPUT50), .ZN(n1197) );
OR2_X1 U985 ( .A1(n1064), .A2(n1063), .ZN(n1061) );
INV_X1 U986 ( .A(n1259), .ZN(n1063) );
NAND2_X1 U987 ( .A1(G221), .A2(n1261), .ZN(n1259) );
NAND2_X1 U988 ( .A1(G234), .A2(n1280), .ZN(n1261) );
XNOR2_X1 U989 ( .A(KEYINPUT12), .B(n1272), .ZN(n1280) );
XOR2_X1 U990 ( .A(n1090), .B(G469), .Z(n1064) );
NAND2_X1 U991 ( .A1(n1281), .A2(n1272), .ZN(n1090) );
XOR2_X1 U992 ( .A(n1167), .B(n1282), .Z(n1281) );
NOR3_X1 U993 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1282) );
NOR2_X1 U994 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NOR2_X1 U995 ( .A1(n1176), .A2(n1288), .ZN(n1286) );
NOR4_X1 U996 ( .A1(n1289), .A2(n1288), .A3(KEYINPUT18), .A4(n1176), .ZN(n1284) );
INV_X1 U997 ( .A(KEYINPUT58), .ZN(n1288) );
INV_X1 U998 ( .A(n1287), .ZN(n1289) );
XOR2_X1 U999 ( .A(G110), .B(n1290), .Z(n1287) );
NOR2_X1 U1000 ( .A1(KEYINPUT59), .A2(n1183), .ZN(n1290) );
AND2_X1 U1001 ( .A1(n1176), .A2(KEYINPUT18), .ZN(n1283) );
NAND2_X1 U1002 ( .A1(G227), .A2(n1036), .ZN(n1176) );
XOR2_X1 U1003 ( .A(n1291), .B(n1292), .Z(n1167) );
XNOR2_X1 U1004 ( .A(n1293), .B(n1162), .ZN(n1292) );
XOR2_X1 U1005 ( .A(n1294), .B(n1295), .Z(n1162) );
XOR2_X1 U1006 ( .A(n1296), .B(KEYINPUT14), .Z(n1294) );
NAND3_X1 U1007 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1296) );
NAND2_X1 U1008 ( .A1(n1106), .A2(n1300), .ZN(n1299) );
NAND2_X1 U1009 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
INV_X1 U1010 ( .A(KEYINPUT13), .ZN(n1302) );
XNOR2_X1 U1011 ( .A(KEYINPUT61), .B(n1103), .ZN(n1301) );
INV_X1 U1012 ( .A(G131), .ZN(n1103) );
OR3_X1 U1013 ( .A1(n1106), .A2(G131), .A3(KEYINPUT13), .ZN(n1298) );
XOR2_X1 U1014 ( .A(G134), .B(G137), .Z(n1106) );
NAND2_X1 U1015 ( .A1(KEYINPUT13), .A2(G131), .ZN(n1297) );
XNOR2_X1 U1016 ( .A(n1303), .B(n1239), .ZN(n1291) );
NAND2_X1 U1017 ( .A1(KEYINPUT57), .A2(n1145), .ZN(n1303) );
NOR2_X1 U1018 ( .A1(n1220), .A2(n1257), .ZN(n1043) );
XNOR2_X1 U1019 ( .A(n1088), .B(n1085), .ZN(n1257) );
XNOR2_X1 U1020 ( .A(n1142), .B(KEYINPUT16), .ZN(n1085) );
INV_X1 U1021 ( .A(G475), .ZN(n1142) );
NOR2_X1 U1022 ( .A1(n1139), .A2(G902), .ZN(n1088) );
XOR2_X1 U1023 ( .A(n1304), .B(n1305), .Z(n1139) );
XOR2_X1 U1024 ( .A(n1306), .B(n1307), .Z(n1305) );
XOR2_X1 U1025 ( .A(n1308), .B(n1309), .Z(n1307) );
NOR2_X1 U1026 ( .A1(G122), .A2(KEYINPUT17), .ZN(n1309) );
NOR3_X1 U1027 ( .A1(n1310), .A2(G953), .A3(G237), .ZN(n1308) );
XOR2_X1 U1028 ( .A(KEYINPUT37), .B(G214), .Z(n1310) );
XNOR2_X1 U1029 ( .A(n1145), .B(n1311), .ZN(n1306) );
NOR2_X1 U1030 ( .A1(KEYINPUT51), .A2(n1312), .ZN(n1311) );
XOR2_X1 U1031 ( .A(n1313), .B(n1314), .Z(n1312) );
XNOR2_X1 U1032 ( .A(G146), .B(KEYINPUT19), .ZN(n1314) );
NAND2_X1 U1033 ( .A1(n1315), .A2(n1316), .ZN(n1313) );
OR2_X1 U1034 ( .A1(n1183), .A2(G125), .ZN(n1316) );
XOR2_X1 U1035 ( .A(n1317), .B(KEYINPUT3), .Z(n1315) );
NAND2_X1 U1036 ( .A1(G125), .A2(n1183), .ZN(n1317) );
INV_X1 U1037 ( .A(G140), .ZN(n1183) );
XOR2_X1 U1038 ( .A(n1318), .B(n1319), .Z(n1304) );
XOR2_X1 U1039 ( .A(KEYINPUT9), .B(G143), .Z(n1319) );
XNOR2_X1 U1040 ( .A(G113), .B(G131), .ZN(n1318) );
INV_X1 U1041 ( .A(n1256), .ZN(n1220) );
XNOR2_X1 U1042 ( .A(n1320), .B(n1080), .ZN(n1256) );
NOR2_X1 U1043 ( .A1(n1130), .A2(G902), .ZN(n1080) );
XNOR2_X1 U1044 ( .A(n1321), .B(n1322), .ZN(n1130) );
XOR2_X1 U1045 ( .A(G128), .B(n1323), .Z(n1322) );
XOR2_X1 U1046 ( .A(G143), .B(G134), .Z(n1323) );
XOR2_X1 U1047 ( .A(n1324), .B(n1325), .Z(n1321) );
AND2_X1 U1048 ( .A1(n1269), .A2(G217), .ZN(n1325) );
AND2_X1 U1049 ( .A1(G234), .A2(n1036), .ZN(n1269) );
INV_X1 U1050 ( .A(G953), .ZN(n1036) );
NAND2_X1 U1051 ( .A1(n1326), .A2(n1327), .ZN(n1324) );
NAND2_X1 U1052 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NAND2_X1 U1053 ( .A1(KEYINPUT8), .A2(n1330), .ZN(n1329) );
OR2_X1 U1054 ( .A1(n1293), .A2(KEYINPUT0), .ZN(n1330) );
INV_X1 U1055 ( .A(n1331), .ZN(n1328) );
NAND2_X1 U1056 ( .A1(n1293), .A2(n1332), .ZN(n1326) );
NAND2_X1 U1057 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
NAND2_X1 U1058 ( .A1(KEYINPUT8), .A2(n1331), .ZN(n1334) );
XNOR2_X1 U1059 ( .A(n1335), .B(G116), .ZN(n1331) );
NAND2_X1 U1060 ( .A1(KEYINPUT26), .A2(n1336), .ZN(n1335) );
INV_X1 U1061 ( .A(KEYINPUT0), .ZN(n1333) );
NAND2_X1 U1062 ( .A1(KEYINPUT48), .A2(n1134), .ZN(n1320) );
INV_X1 U1063 ( .A(G478), .ZN(n1134) );
XNOR2_X1 U1064 ( .A(n1212), .B(KEYINPUT52), .ZN(n1149) );
NOR2_X1 U1065 ( .A1(n1049), .A2(n1048), .ZN(n1212) );
AND2_X1 U1066 ( .A1(G214), .A2(n1337), .ZN(n1048) );
NAND2_X1 U1067 ( .A1(n1277), .A2(n1272), .ZN(n1337) );
INV_X1 U1068 ( .A(G902), .ZN(n1272) );
INV_X1 U1069 ( .A(n1235), .ZN(n1049) );
NAND3_X1 U1070 ( .A1(n1338), .A2(n1339), .A3(n1340), .ZN(n1235) );
NAND2_X1 U1071 ( .A1(n1341), .A2(n1185), .ZN(n1340) );
OR3_X1 U1072 ( .A1(n1185), .A2(n1341), .A3(G902), .ZN(n1339) );
NOR2_X1 U1073 ( .A1(n1277), .A2(n1188), .ZN(n1341) );
INV_X1 U1074 ( .A(G210), .ZN(n1188) );
INV_X1 U1075 ( .A(G237), .ZN(n1277) );
XOR2_X1 U1076 ( .A(n1342), .B(n1343), .Z(n1185) );
XNOR2_X1 U1077 ( .A(n1295), .B(n1120), .ZN(n1343) );
XNOR2_X1 U1078 ( .A(n1336), .B(G110), .ZN(n1120) );
INV_X1 U1079 ( .A(G122), .ZN(n1336) );
INV_X1 U1080 ( .A(n1105), .ZN(n1295) );
XOR2_X1 U1081 ( .A(G143), .B(n1268), .Z(n1105) );
XOR2_X1 U1082 ( .A(G128), .B(G146), .Z(n1268) );
XOR2_X1 U1083 ( .A(n1344), .B(n1345), .Z(n1342) );
NOR2_X1 U1084 ( .A1(G953), .A2(n1110), .ZN(n1345) );
INV_X1 U1085 ( .A(G224), .ZN(n1110) );
XOR2_X1 U1086 ( .A(n1346), .B(G125), .Z(n1344) );
NAND3_X1 U1087 ( .A1(n1347), .A2(n1348), .A3(n1349), .ZN(n1346) );
NAND2_X1 U1088 ( .A1(n1350), .A2(n1118), .ZN(n1349) );
NAND2_X1 U1089 ( .A1(KEYINPUT5), .A2(n1351), .ZN(n1348) );
NAND2_X1 U1090 ( .A1(n1352), .A2(n1119), .ZN(n1351) );
XNOR2_X1 U1091 ( .A(KEYINPUT22), .B(n1118), .ZN(n1352) );
NAND2_X1 U1092 ( .A1(n1353), .A2(n1354), .ZN(n1347) );
INV_X1 U1093 ( .A(KEYINPUT5), .ZN(n1354) );
NAND2_X1 U1094 ( .A1(n1355), .A2(n1356), .ZN(n1353) );
OR3_X1 U1095 ( .A1(n1350), .A2(n1118), .A3(KEYINPUT22), .ZN(n1356) );
INV_X1 U1096 ( .A(n1119), .ZN(n1350) );
XOR2_X1 U1097 ( .A(n1357), .B(n1293), .Z(n1119) );
XNOR2_X1 U1098 ( .A(G107), .B(KEYINPUT60), .ZN(n1293) );
XNOR2_X1 U1099 ( .A(n1358), .B(n1239), .ZN(n1357) );
INV_X1 U1100 ( .A(G101), .ZN(n1239) );
NAND2_X1 U1101 ( .A1(KEYINPUT35), .A2(n1145), .ZN(n1358) );
INV_X1 U1102 ( .A(G104), .ZN(n1145) );
NAND2_X1 U1103 ( .A1(KEYINPUT22), .A2(n1118), .ZN(n1355) );
INV_X1 U1104 ( .A(n1165), .ZN(n1118) );
XOR2_X1 U1105 ( .A(G113), .B(n1359), .Z(n1165) );
XOR2_X1 U1106 ( .A(G119), .B(G116), .Z(n1359) );
NAND2_X1 U1107 ( .A1(G902), .A2(G210), .ZN(n1338) );
endmodule


