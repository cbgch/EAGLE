//Key = 0010111001101011101011111111000101010000010101100110101111100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
n1415, n1416, n1417, n1418, n1419;

XOR2_X1 U776 ( .A(n1075), .B(n1076), .Z(G9) );
NOR2_X1 U777 ( .A1(n1077), .A2(n1078), .ZN(G75) );
XOR2_X1 U778 ( .A(n1079), .B(KEYINPUT2), .Z(n1078) );
NAND3_X1 U779 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
XOR2_X1 U780 ( .A(KEYINPUT16), .B(G952), .Z(n1082) );
NOR4_X1 U781 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1077) );
XOR2_X1 U782 ( .A(n1087), .B(KEYINPUT37), .Z(n1085) );
NAND2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U784 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
NAND2_X1 U785 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NAND4_X1 U786 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1094) );
NAND2_X1 U787 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U788 ( .A1(n1101), .A2(n1102), .ZN(n1097) );
NAND2_X1 U789 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NAND2_X1 U790 ( .A1(n1105), .A2(n1106), .ZN(n1093) );
XOR2_X1 U791 ( .A(n1107), .B(KEYINPUT44), .Z(n1088) );
NAND4_X1 U792 ( .A1(n1092), .A2(n1105), .A3(n1096), .A4(n1108), .ZN(n1107) );
NAND3_X1 U793 ( .A1(n1080), .A2(n1081), .A3(n1109), .ZN(n1083) );
NAND2_X1 U794 ( .A1(n1092), .A2(n1110), .ZN(n1109) );
NAND2_X1 U795 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND3_X1 U796 ( .A1(n1113), .A2(n1090), .A3(n1105), .ZN(n1112) );
NAND2_X1 U797 ( .A1(n1096), .A2(n1114), .ZN(n1111) );
NAND2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U799 ( .A1(n1090), .A2(n1117), .ZN(n1116) );
NAND2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U801 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U802 ( .A1(n1105), .A2(n1122), .ZN(n1115) );
NOR3_X1 U803 ( .A1(n1123), .A2(n1099), .A3(n1100), .ZN(n1105) );
INV_X1 U804 ( .A(n1120), .ZN(n1100) );
INV_X1 U805 ( .A(n1124), .ZN(n1092) );
NAND4_X1 U806 ( .A1(n1125), .A2(n1120), .A3(n1126), .A4(n1127), .ZN(n1080) );
NOR3_X1 U807 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1127) );
XNOR2_X1 U808 ( .A(n1131), .B(n1132), .ZN(n1129) );
NAND2_X1 U809 ( .A1(KEYINPUT49), .A2(n1133), .ZN(n1131) );
NAND3_X1 U810 ( .A1(n1134), .A2(n1135), .A3(n1102), .ZN(n1128) );
NOR4_X1 U811 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1126) );
NOR3_X1 U812 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
AND2_X1 U813 ( .A1(n1140), .A2(n1142), .ZN(n1138) );
INV_X1 U814 ( .A(KEYINPUT9), .ZN(n1140) );
NOR3_X1 U815 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1137) );
INV_X1 U816 ( .A(KEYINPUT45), .ZN(n1143) );
NOR2_X1 U817 ( .A1(KEYINPUT45), .A2(G475), .ZN(n1136) );
NAND3_X1 U818 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(G72) );
NAND2_X1 U819 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
INV_X1 U820 ( .A(KEYINPUT43), .ZN(n1150) );
OR2_X1 U821 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
NAND3_X1 U822 ( .A1(KEYINPUT43), .A2(n1153), .A3(n1154), .ZN(n1147) );
INV_X1 U823 ( .A(n1152), .ZN(n1154) );
NAND2_X1 U824 ( .A1(n1151), .A2(n1155), .ZN(n1153) );
NAND2_X1 U825 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U826 ( .A1(n1152), .A2(n1151), .ZN(n1146) );
NAND2_X1 U827 ( .A1(G953), .A2(n1158), .ZN(n1151) );
NAND2_X1 U828 ( .A1(G900), .A2(G227), .ZN(n1158) );
NOR3_X1 U829 ( .A1(n1156), .A2(n1159), .A3(n1157), .ZN(n1152) );
NAND2_X1 U830 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NOR2_X1 U831 ( .A1(n1081), .A2(G900), .ZN(n1159) );
XNOR2_X1 U832 ( .A(n1162), .B(n1163), .ZN(n1156) );
XOR2_X1 U833 ( .A(KEYINPUT6), .B(n1164), .Z(n1163) );
XOR2_X1 U834 ( .A(n1165), .B(n1166), .Z(G69) );
XOR2_X1 U835 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U836 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
XOR2_X1 U837 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U838 ( .A(n1173), .B(n1174), .Z(n1172) );
NAND2_X1 U839 ( .A1(n1175), .A2(n1176), .ZN(n1173) );
XNOR2_X1 U840 ( .A(KEYINPUT24), .B(KEYINPUT21), .ZN(n1175) );
NOR2_X1 U841 ( .A1(G898), .A2(n1081), .ZN(n1169) );
NOR2_X1 U842 ( .A1(G953), .A2(n1177), .ZN(n1167) );
NOR2_X1 U843 ( .A1(n1178), .A2(n1081), .ZN(n1165) );
NOR2_X1 U844 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NOR2_X1 U845 ( .A1(n1181), .A2(n1182), .ZN(G66) );
XNOR2_X1 U846 ( .A(n1183), .B(n1184), .ZN(n1182) );
NOR2_X1 U847 ( .A1(n1142), .A2(n1185), .ZN(n1184) );
NOR2_X1 U848 ( .A1(n1181), .A2(n1186), .ZN(G63) );
XOR2_X1 U849 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND3_X1 U850 ( .A1(n1189), .A2(n1190), .A3(G478), .ZN(n1187) );
NAND2_X1 U851 ( .A1(KEYINPUT52), .A2(n1185), .ZN(n1190) );
NAND2_X1 U852 ( .A1(n1191), .A2(n1192), .ZN(n1189) );
INV_X1 U853 ( .A(KEYINPUT52), .ZN(n1192) );
OR2_X1 U854 ( .A1(n1084), .A2(n1193), .ZN(n1191) );
NOR2_X1 U855 ( .A1(n1181), .A2(n1194), .ZN(G60) );
XOR2_X1 U856 ( .A(n1195), .B(n1196), .Z(n1194) );
NOR2_X1 U857 ( .A1(n1145), .A2(n1185), .ZN(n1195) );
XNOR2_X1 U858 ( .A(G104), .B(n1197), .ZN(G6) );
NAND2_X1 U859 ( .A1(n1113), .A2(n1198), .ZN(n1197) );
NOR4_X1 U860 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(G57) );
AND3_X1 U861 ( .A1(KEYINPUT8), .A2(n1081), .A3(n1086), .ZN(n1202) );
NOR2_X1 U862 ( .A1(KEYINPUT8), .A2(n1203), .ZN(n1201) );
AND3_X1 U863 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1200) );
OR2_X1 U864 ( .A1(n1207), .A2(n1208), .ZN(n1205) );
XOR2_X1 U865 ( .A(n1209), .B(n1210), .Z(n1208) );
NOR2_X1 U866 ( .A1(n1211), .A2(n1204), .ZN(n1199) );
NAND2_X1 U867 ( .A1(KEYINPUT25), .A2(n1212), .ZN(n1204) );
NOR2_X1 U868 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
NOR2_X1 U869 ( .A1(n1209), .A2(n1206), .ZN(n1214) );
NAND2_X1 U870 ( .A1(n1207), .A2(n1210), .ZN(n1206) );
INV_X1 U871 ( .A(n1215), .ZN(n1207) );
NOR2_X1 U872 ( .A1(n1216), .A2(n1210), .ZN(n1213) );
NAND2_X1 U873 ( .A1(n1217), .A2(n1218), .ZN(n1210) );
XOR2_X1 U874 ( .A(n1219), .B(KEYINPUT34), .Z(n1217) );
NAND3_X1 U875 ( .A1(G210), .A2(n1220), .A3(n1221), .ZN(n1219) );
XOR2_X1 U876 ( .A(KEYINPUT48), .B(G101), .Z(n1220) );
NOR2_X1 U877 ( .A1(n1215), .A2(n1209), .ZN(n1216) );
INV_X1 U878 ( .A(KEYINPUT15), .ZN(n1209) );
NOR2_X1 U879 ( .A1(n1185), .A2(n1133), .ZN(n1215) );
INV_X1 U880 ( .A(G472), .ZN(n1133) );
NOR3_X1 U881 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(G54) );
AND2_X1 U882 ( .A1(n1181), .A2(KEYINPUT56), .ZN(n1224) );
NOR3_X1 U883 ( .A1(KEYINPUT56), .A2(G953), .A3(G952), .ZN(n1223) );
XOR2_X1 U884 ( .A(n1225), .B(n1226), .Z(n1222) );
NOR2_X1 U885 ( .A1(n1227), .A2(n1185), .ZN(n1226) );
INV_X1 U886 ( .A(G469), .ZN(n1227) );
NOR2_X1 U887 ( .A1(n1228), .A2(n1229), .ZN(n1225) );
XOR2_X1 U888 ( .A(KEYINPUT61), .B(n1230), .Z(n1229) );
NOR2_X1 U889 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
AND2_X1 U890 ( .A1(n1231), .A2(n1232), .ZN(n1228) );
XNOR2_X1 U891 ( .A(n1233), .B(n1234), .ZN(n1232) );
NOR2_X1 U892 ( .A1(n1181), .A2(n1235), .ZN(G51) );
XOR2_X1 U893 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U894 ( .A(n1238), .B(n1239), .Z(n1237) );
NOR2_X1 U895 ( .A1(n1240), .A2(n1185), .ZN(n1239) );
NAND2_X1 U896 ( .A1(G902), .A2(n1084), .ZN(n1185) );
NAND3_X1 U897 ( .A1(n1160), .A2(n1241), .A3(n1177), .ZN(n1084) );
AND2_X1 U898 ( .A1(n1242), .A2(n1243), .ZN(n1177) );
AND4_X1 U899 ( .A1(n1244), .A2(n1076), .A3(n1245), .A4(n1246), .ZN(n1243) );
NAND2_X1 U900 ( .A1(n1198), .A2(n1106), .ZN(n1076) );
AND2_X1 U901 ( .A1(n1247), .A2(n1090), .ZN(n1198) );
NOR4_X1 U902 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1242) );
NOR3_X1 U903 ( .A1(n1252), .A2(n1253), .A3(n1118), .ZN(n1251) );
NOR4_X1 U904 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1250) );
XOR2_X1 U905 ( .A(n1258), .B(KEYINPUT20), .Z(n1257) );
XOR2_X1 U906 ( .A(n1259), .B(KEYINPUT29), .Z(n1256) );
NAND2_X1 U907 ( .A1(n1113), .A2(n1090), .ZN(n1254) );
INV_X1 U908 ( .A(n1260), .ZN(n1249) );
XNOR2_X1 U909 ( .A(KEYINPUT54), .B(n1161), .ZN(n1241) );
AND4_X1 U910 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1160) );
AND4_X1 U911 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1264) );
NAND3_X1 U912 ( .A1(n1269), .A2(n1096), .A3(n1270), .ZN(n1263) );
NAND4_X1 U913 ( .A1(n1120), .A2(n1271), .A3(n1272), .A4(n1273), .ZN(n1261) );
XOR2_X1 U914 ( .A(KEYINPUT62), .B(n1121), .Z(n1272) );
INV_X1 U915 ( .A(n1252), .ZN(n1271) );
NAND3_X1 U916 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1238) );
XNOR2_X1 U917 ( .A(KEYINPUT60), .B(KEYINPUT30), .ZN(n1276) );
NAND2_X1 U918 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
XOR2_X1 U919 ( .A(KEYINPUT12), .B(n1279), .Z(n1277) );
NAND2_X1 U920 ( .A1(n1279), .A2(n1280), .ZN(n1274) );
XOR2_X1 U921 ( .A(G125), .B(n1281), .Z(n1279) );
INV_X1 U922 ( .A(n1203), .ZN(n1181) );
NAND2_X1 U923 ( .A1(G953), .A2(n1086), .ZN(n1203) );
INV_X1 U924 ( .A(G952), .ZN(n1086) );
NAND2_X1 U925 ( .A1(n1282), .A2(n1283), .ZN(G48) );
NAND2_X1 U926 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NAND2_X1 U927 ( .A1(n1262), .A2(n1286), .ZN(n1284) );
OR2_X1 U928 ( .A1(KEYINPUT13), .A2(KEYINPUT50), .ZN(n1286) );
NAND3_X1 U929 ( .A1(n1287), .A2(n1288), .A3(KEYINPUT50), .ZN(n1282) );
OR2_X1 U930 ( .A1(n1262), .A2(KEYINPUT13), .ZN(n1288) );
NAND2_X1 U931 ( .A1(n1289), .A2(n1262), .ZN(n1287) );
NAND3_X1 U932 ( .A1(n1269), .A2(n1113), .A3(n1290), .ZN(n1262) );
OR2_X1 U933 ( .A1(n1285), .A2(KEYINPUT13), .ZN(n1289) );
XNOR2_X1 U934 ( .A(G143), .B(n1268), .ZN(G45) );
NAND4_X1 U935 ( .A1(n1290), .A2(n1122), .A3(n1291), .A4(n1292), .ZN(n1268) );
NAND2_X1 U936 ( .A1(n1293), .A2(n1294), .ZN(G42) );
NAND3_X1 U937 ( .A1(n1295), .A2(KEYINPUT23), .A3(n1296), .ZN(n1294) );
INV_X1 U938 ( .A(G140), .ZN(n1296) );
NAND2_X1 U939 ( .A1(G140), .A2(n1297), .ZN(n1293) );
NAND2_X1 U940 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NAND2_X1 U941 ( .A1(n1295), .A2(n1300), .ZN(n1299) );
NAND2_X1 U942 ( .A1(KEYINPUT23), .A2(n1301), .ZN(n1300) );
INV_X1 U943 ( .A(n1267), .ZN(n1295) );
NAND2_X1 U944 ( .A1(n1301), .A2(n1267), .ZN(n1298) );
NAND3_X1 U945 ( .A1(n1113), .A2(n1108), .A3(n1270), .ZN(n1267) );
XOR2_X1 U946 ( .A(KEYINPUT42), .B(KEYINPUT27), .Z(n1301) );
XOR2_X1 U947 ( .A(n1302), .B(n1303), .Z(G39) );
NAND2_X1 U948 ( .A1(KEYINPUT41), .A2(G137), .ZN(n1303) );
NAND3_X1 U949 ( .A1(n1270), .A2(n1269), .A3(n1304), .ZN(n1302) );
XNOR2_X1 U950 ( .A(n1096), .B(KEYINPUT4), .ZN(n1304) );
XOR2_X1 U951 ( .A(G134), .B(n1305), .Z(G36) );
NOR2_X1 U952 ( .A1(n1252), .A2(n1306), .ZN(n1305) );
XOR2_X1 U953 ( .A(n1266), .B(n1307), .Z(G33) );
NOR2_X1 U954 ( .A1(G131), .A2(KEYINPUT3), .ZN(n1307) );
NAND3_X1 U955 ( .A1(n1113), .A2(n1122), .A3(n1270), .ZN(n1266) );
INV_X1 U956 ( .A(n1306), .ZN(n1270) );
NAND3_X1 U957 ( .A1(n1121), .A2(n1273), .A3(n1120), .ZN(n1306) );
NOR2_X1 U958 ( .A1(n1308), .A2(n1103), .ZN(n1120) );
XOR2_X1 U959 ( .A(n1309), .B(n1161), .Z(G30) );
NAND3_X1 U960 ( .A1(n1269), .A2(n1106), .A3(n1290), .ZN(n1161) );
AND3_X1 U961 ( .A1(n1310), .A2(n1273), .A3(n1121), .ZN(n1290) );
INV_X1 U962 ( .A(n1255), .ZN(n1121) );
XOR2_X1 U963 ( .A(n1311), .B(n1260), .Z(G3) );
NAND3_X1 U964 ( .A1(n1247), .A2(n1122), .A3(n1096), .ZN(n1260) );
XNOR2_X1 U965 ( .A(n1265), .B(n1312), .ZN(G27) );
NOR2_X1 U966 ( .A1(KEYINPUT39), .A2(n1313), .ZN(n1312) );
NAND4_X1 U967 ( .A1(n1314), .A2(n1113), .A3(n1108), .A4(n1273), .ZN(n1265) );
NAND2_X1 U968 ( .A1(n1124), .A2(n1315), .ZN(n1273) );
NAND4_X1 U969 ( .A1(G953), .A2(G902), .A3(n1316), .A4(n1317), .ZN(n1315) );
INV_X1 U970 ( .A(G900), .ZN(n1317) );
XOR2_X1 U971 ( .A(n1318), .B(n1248), .Z(G24) );
AND3_X1 U972 ( .A1(n1314), .A2(n1090), .A3(n1319), .ZN(n1248) );
NOR3_X1 U973 ( .A1(n1125), .A2(n1253), .A3(n1320), .ZN(n1319) );
NAND2_X1 U974 ( .A1(KEYINPUT26), .A2(n1321), .ZN(n1318) );
NAND2_X1 U975 ( .A1(n1322), .A2(n1323), .ZN(G21) );
OR2_X1 U976 ( .A1(n1246), .A2(G119), .ZN(n1323) );
XOR2_X1 U977 ( .A(n1324), .B(KEYINPUT40), .Z(n1322) );
NAND2_X1 U978 ( .A1(G119), .A2(n1246), .ZN(n1324) );
NAND4_X1 U979 ( .A1(n1269), .A2(n1314), .A3(n1096), .A4(n1258), .ZN(n1246) );
INV_X1 U980 ( .A(n1118), .ZN(n1314) );
AND2_X1 U981 ( .A1(n1325), .A2(n1326), .ZN(n1269) );
XOR2_X1 U982 ( .A(KEYINPUT17), .B(n1327), .Z(n1325) );
XOR2_X1 U983 ( .A(G116), .B(n1328), .Z(G18) );
NOR3_X1 U984 ( .A1(n1252), .A2(n1329), .A3(n1118), .ZN(n1328) );
NAND3_X1 U985 ( .A1(n1310), .A2(n1102), .A3(n1095), .ZN(n1118) );
XOR2_X1 U986 ( .A(n1258), .B(KEYINPUT57), .Z(n1329) );
NAND2_X1 U987 ( .A1(n1106), .A2(n1122), .ZN(n1252) );
NOR2_X1 U988 ( .A1(n1292), .A2(n1125), .ZN(n1106) );
XNOR2_X1 U989 ( .A(G113), .B(n1245), .ZN(G15) );
NAND4_X1 U990 ( .A1(n1095), .A2(n1122), .A3(n1113), .A4(n1330), .ZN(n1245) );
NOR3_X1 U991 ( .A1(n1259), .A2(n1253), .A3(n1099), .ZN(n1330) );
INV_X1 U992 ( .A(n1102), .ZN(n1099) );
NOR2_X1 U993 ( .A1(n1291), .A2(n1320), .ZN(n1113) );
INV_X1 U994 ( .A(n1292), .ZN(n1320) );
NAND2_X1 U995 ( .A1(n1331), .A2(n1332), .ZN(n1122) );
OR3_X1 U996 ( .A1(n1326), .A2(n1333), .A3(KEYINPUT17), .ZN(n1332) );
NAND2_X1 U997 ( .A1(KEYINPUT17), .A2(n1090), .ZN(n1331) );
NOR2_X1 U998 ( .A1(n1326), .A2(n1327), .ZN(n1090) );
INV_X1 U999 ( .A(n1333), .ZN(n1327) );
XNOR2_X1 U1000 ( .A(G110), .B(n1244), .ZN(G12) );
NAND3_X1 U1001 ( .A1(n1108), .A2(n1247), .A3(n1096), .ZN(n1244) );
NOR2_X1 U1002 ( .A1(n1291), .A2(n1292), .ZN(n1096) );
NAND2_X1 U1003 ( .A1(n1134), .A2(n1334), .ZN(n1292) );
OR2_X1 U1004 ( .A1(n1145), .A2(n1144), .ZN(n1334) );
NAND2_X1 U1005 ( .A1(n1144), .A2(n1145), .ZN(n1134) );
INV_X1 U1006 ( .A(G475), .ZN(n1145) );
NOR2_X1 U1007 ( .A1(n1196), .A2(G902), .ZN(n1144) );
XNOR2_X1 U1008 ( .A(n1335), .B(n1336), .ZN(n1196) );
XNOR2_X1 U1009 ( .A(G104), .B(n1337), .ZN(n1336) );
NAND2_X1 U1010 ( .A1(KEYINPUT58), .A2(n1338), .ZN(n1337) );
XOR2_X1 U1011 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1012 ( .A(n1341), .B(n1342), .Z(n1340) );
NAND2_X1 U1013 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
XNOR2_X1 U1014 ( .A(KEYINPUT33), .B(KEYINPUT18), .ZN(n1343) );
NAND2_X1 U1015 ( .A1(n1345), .A2(n1346), .ZN(n1341) );
NAND2_X1 U1016 ( .A1(G146), .A2(n1164), .ZN(n1346) );
XOR2_X1 U1017 ( .A(KEYINPUT10), .B(n1347), .Z(n1345) );
NOR2_X1 U1018 ( .A1(G146), .A2(n1164), .ZN(n1347) );
XOR2_X1 U1019 ( .A(G140), .B(G125), .Z(n1164) );
XNOR2_X1 U1020 ( .A(G143), .B(n1348), .ZN(n1339) );
NAND2_X1 U1021 ( .A1(n1221), .A2(G214), .ZN(n1348) );
XOR2_X1 U1022 ( .A(G113), .B(n1321), .Z(n1335) );
INV_X1 U1023 ( .A(n1125), .ZN(n1291) );
XOR2_X1 U1024 ( .A(n1349), .B(G478), .Z(n1125) );
NAND2_X1 U1025 ( .A1(n1188), .A2(n1193), .ZN(n1349) );
XNOR2_X1 U1026 ( .A(n1350), .B(n1351), .ZN(n1188) );
XOR2_X1 U1027 ( .A(n1352), .B(n1353), .Z(n1351) );
XOR2_X1 U1028 ( .A(n1354), .B(n1355), .Z(n1350) );
XOR2_X1 U1029 ( .A(G122), .B(G107), .Z(n1355) );
NAND2_X1 U1030 ( .A1(n1356), .A2(G217), .ZN(n1354) );
NOR3_X1 U1031 ( .A1(n1259), .A2(n1253), .A3(n1255), .ZN(n1247) );
NAND2_X1 U1032 ( .A1(n1123), .A2(n1102), .ZN(n1255) );
NAND2_X1 U1033 ( .A1(G221), .A2(n1357), .ZN(n1102) );
INV_X1 U1034 ( .A(n1095), .ZN(n1123) );
XNOR2_X1 U1035 ( .A(n1130), .B(KEYINPUT53), .ZN(n1095) );
XNOR2_X1 U1036 ( .A(n1358), .B(G469), .ZN(n1130) );
NAND2_X1 U1037 ( .A1(n1359), .A2(n1193), .ZN(n1358) );
XNOR2_X1 U1038 ( .A(n1231), .B(n1360), .ZN(n1359) );
XOR2_X1 U1039 ( .A(n1233), .B(n1361), .Z(n1360) );
NAND2_X1 U1040 ( .A1(KEYINPUT63), .A2(n1234), .ZN(n1361) );
NAND2_X1 U1041 ( .A1(G227), .A2(n1081), .ZN(n1233) );
XNOR2_X1 U1042 ( .A(n1162), .B(n1362), .ZN(n1231) );
NOR2_X1 U1043 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
XOR2_X1 U1044 ( .A(KEYINPUT47), .B(n1365), .Z(n1364) );
NOR2_X1 U1045 ( .A1(G101), .A2(n1366), .ZN(n1365) );
AND2_X1 U1046 ( .A1(n1366), .A2(G101), .ZN(n1363) );
XOR2_X1 U1047 ( .A(G104), .B(G107), .Z(n1366) );
XOR2_X1 U1048 ( .A(n1367), .B(n1368), .Z(n1162) );
INV_X1 U1049 ( .A(n1369), .ZN(n1368) );
NAND2_X1 U1050 ( .A1(KEYINPUT14), .A2(n1309), .ZN(n1367) );
INV_X1 U1051 ( .A(n1258), .ZN(n1253) );
NAND2_X1 U1052 ( .A1(n1370), .A2(n1124), .ZN(n1258) );
NAND3_X1 U1053 ( .A1(n1316), .A2(n1081), .A3(G952), .ZN(n1124) );
NAND4_X1 U1054 ( .A1(G953), .A2(G902), .A3(n1316), .A4(n1180), .ZN(n1370) );
INV_X1 U1055 ( .A(G898), .ZN(n1180) );
NAND2_X1 U1056 ( .A1(G237), .A2(G234), .ZN(n1316) );
XNOR2_X1 U1057 ( .A(n1310), .B(KEYINPUT28), .ZN(n1259) );
NOR2_X1 U1058 ( .A1(n1104), .A2(n1103), .ZN(n1310) );
AND2_X1 U1059 ( .A1(G214), .A2(n1371), .ZN(n1103) );
NAND2_X1 U1060 ( .A1(n1193), .A2(n1372), .ZN(n1371) );
INV_X1 U1061 ( .A(n1308), .ZN(n1104) );
NAND3_X1 U1062 ( .A1(n1373), .A2(n1374), .A3(n1375), .ZN(n1308) );
NAND2_X1 U1063 ( .A1(n1376), .A2(n1377), .ZN(n1375) );
OR3_X1 U1064 ( .A1(n1377), .A2(n1376), .A3(G902), .ZN(n1374) );
NOR2_X1 U1065 ( .A1(n1240), .A2(n1372), .ZN(n1376) );
INV_X1 U1066 ( .A(G237), .ZN(n1372) );
INV_X1 U1067 ( .A(G210), .ZN(n1240) );
XOR2_X1 U1068 ( .A(n1236), .B(n1378), .Z(n1377) );
XNOR2_X1 U1069 ( .A(n1281), .B(n1379), .ZN(n1378) );
NAND2_X1 U1070 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
NAND2_X1 U1071 ( .A1(n1280), .A2(n1313), .ZN(n1381) );
INV_X1 U1072 ( .A(n1278), .ZN(n1280) );
XOR2_X1 U1073 ( .A(n1382), .B(KEYINPUT11), .Z(n1380) );
NAND2_X1 U1074 ( .A1(G125), .A2(n1278), .ZN(n1382) );
XOR2_X1 U1075 ( .A(n1383), .B(n1384), .Z(n1278) );
XOR2_X1 U1076 ( .A(n1309), .B(G143), .Z(n1383) );
INV_X1 U1077 ( .A(G128), .ZN(n1309) );
NOR2_X1 U1078 ( .A1(n1179), .A2(G953), .ZN(n1281) );
INV_X1 U1079 ( .A(G224), .ZN(n1179) );
XOR2_X1 U1080 ( .A(n1174), .B(n1385), .Z(n1236) );
NOR2_X1 U1081 ( .A1(KEYINPUT38), .A2(n1386), .ZN(n1385) );
XOR2_X1 U1082 ( .A(n1171), .B(n1176), .Z(n1386) );
XOR2_X1 U1083 ( .A(n1387), .B(G101), .Z(n1176) );
NAND3_X1 U1084 ( .A1(KEYINPUT46), .A2(n1388), .A3(n1389), .ZN(n1387) );
XOR2_X1 U1085 ( .A(n1390), .B(KEYINPUT19), .Z(n1389) );
NAND2_X1 U1086 ( .A1(G104), .A2(n1075), .ZN(n1390) );
OR2_X1 U1087 ( .A1(n1075), .A2(G104), .ZN(n1388) );
INV_X1 U1088 ( .A(G107), .ZN(n1075) );
XNOR2_X1 U1089 ( .A(n1391), .B(n1392), .ZN(n1171) );
NAND2_X1 U1090 ( .A1(KEYINPUT55), .A2(n1393), .ZN(n1391) );
INV_X1 U1091 ( .A(G116), .ZN(n1393) );
XOR2_X1 U1092 ( .A(G110), .B(n1321), .Z(n1174) );
INV_X1 U1093 ( .A(G122), .ZN(n1321) );
NAND2_X1 U1094 ( .A1(G210), .A2(G902), .ZN(n1373) );
AND2_X1 U1095 ( .A1(n1394), .A2(n1326), .ZN(n1108) );
NAND2_X1 U1096 ( .A1(n1135), .A2(n1395), .ZN(n1326) );
OR2_X1 U1097 ( .A1(n1142), .A2(n1141), .ZN(n1395) );
NAND2_X1 U1098 ( .A1(n1141), .A2(n1142), .ZN(n1135) );
NAND2_X1 U1099 ( .A1(G217), .A2(n1357), .ZN(n1142) );
NAND2_X1 U1100 ( .A1(G234), .A2(n1193), .ZN(n1357) );
AND2_X1 U1101 ( .A1(n1193), .A2(n1183), .ZN(n1141) );
NAND2_X1 U1102 ( .A1(n1396), .A2(n1397), .ZN(n1183) );
NAND2_X1 U1103 ( .A1(n1398), .A2(n1399), .ZN(n1397) );
XOR2_X1 U1104 ( .A(KEYINPUT5), .B(n1400), .Z(n1396) );
NOR2_X1 U1105 ( .A1(n1398), .A2(n1399), .ZN(n1400) );
XNOR2_X1 U1106 ( .A(n1401), .B(n1402), .ZN(n1399) );
XNOR2_X1 U1107 ( .A(n1403), .B(n1234), .ZN(n1402) );
XOR2_X1 U1108 ( .A(G110), .B(G140), .Z(n1234) );
NAND2_X1 U1109 ( .A1(KEYINPUT35), .A2(n1313), .ZN(n1403) );
INV_X1 U1110 ( .A(G125), .ZN(n1313) );
XOR2_X1 U1111 ( .A(n1285), .B(n1404), .Z(n1401) );
NOR2_X1 U1112 ( .A1(KEYINPUT51), .A2(n1405), .ZN(n1404) );
XOR2_X1 U1113 ( .A(G119), .B(n1406), .Z(n1405) );
NOR2_X1 U1114 ( .A1(G128), .A2(KEYINPUT36), .ZN(n1406) );
INV_X1 U1115 ( .A(G146), .ZN(n1285) );
XNOR2_X1 U1116 ( .A(n1407), .B(G137), .ZN(n1398) );
NAND2_X1 U1117 ( .A1(n1356), .A2(G221), .ZN(n1407) );
AND2_X1 U1118 ( .A1(G234), .A2(n1081), .ZN(n1356) );
INV_X1 U1119 ( .A(G953), .ZN(n1081) );
XOR2_X1 U1120 ( .A(n1333), .B(KEYINPUT32), .Z(n1394) );
XOR2_X1 U1121 ( .A(n1132), .B(n1408), .Z(n1333) );
XOR2_X1 U1122 ( .A(KEYINPUT0), .B(G472), .Z(n1408) );
NAND2_X1 U1123 ( .A1(n1409), .A2(n1193), .ZN(n1132) );
INV_X1 U1124 ( .A(G902), .ZN(n1193) );
XOR2_X1 U1125 ( .A(n1212), .B(n1410), .Z(n1409) );
XOR2_X1 U1126 ( .A(n1411), .B(KEYINPUT7), .Z(n1410) );
NAND2_X1 U1127 ( .A1(n1412), .A2(n1413), .ZN(n1411) );
NAND3_X1 U1128 ( .A1(G210), .A2(G101), .A3(n1221), .ZN(n1413) );
XOR2_X1 U1129 ( .A(n1218), .B(KEYINPUT1), .Z(n1412) );
NAND2_X1 U1130 ( .A1(n1311), .A2(n1414), .ZN(n1218) );
NAND2_X1 U1131 ( .A1(n1221), .A2(G210), .ZN(n1414) );
NOR2_X1 U1132 ( .A1(G953), .A2(G237), .ZN(n1221) );
INV_X1 U1133 ( .A(G101), .ZN(n1311) );
XOR2_X1 U1134 ( .A(n1415), .B(n1416), .Z(n1212) );
XOR2_X1 U1135 ( .A(KEYINPUT31), .B(n1353), .Z(n1416) );
XOR2_X1 U1136 ( .A(G116), .B(G128), .Z(n1353) );
XOR2_X1 U1137 ( .A(n1369), .B(n1392), .Z(n1415) );
XOR2_X1 U1138 ( .A(G113), .B(n1417), .Z(n1392) );
XOR2_X1 U1139 ( .A(KEYINPUT22), .B(G119), .Z(n1417) );
XOR2_X1 U1140 ( .A(n1418), .B(n1419), .Z(n1369) );
XOR2_X1 U1141 ( .A(n1352), .B(n1384), .Z(n1419) );
XOR2_X1 U1142 ( .A(G146), .B(KEYINPUT59), .Z(n1384) );
XOR2_X1 U1143 ( .A(G134), .B(G143), .Z(n1352) );
XOR2_X1 U1144 ( .A(n1344), .B(G137), .Z(n1418) );
INV_X1 U1145 ( .A(G131), .ZN(n1344) );
endmodule


