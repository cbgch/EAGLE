//Key = 0000110001110100110111101110111011010101011011100010111001001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340;

XOR2_X1 U730 ( .A(G107), .B(n1015), .Z(G9) );
NOR2_X1 U731 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U732 ( .A1(G953), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1017) );
NOR2_X1 U733 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR2_X1 U734 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR3_X1 U735 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1024) );
NOR2_X1 U736 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR2_X1 U737 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR2_X1 U738 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR2_X1 U739 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR2_X1 U740 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U741 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U742 ( .A1(n1040), .A2(n1041), .ZN(n1032) );
NOR2_X1 U743 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U744 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR3_X1 U745 ( .A1(n1041), .A2(n1046), .A3(n1035), .ZN(n1028) );
NOR2_X1 U746 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR4_X1 U747 ( .A1(n1049), .A2(n1035), .A3(n1031), .A4(n1041), .ZN(n1023) );
NOR2_X1 U748 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U749 ( .A1(n1025), .A2(n1052), .ZN(n1050) );
NOR3_X1 U750 ( .A1(n1018), .A2(G953), .A3(G952), .ZN(n1016) );
AND4_X1 U751 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1018) );
NOR4_X1 U752 ( .A1(n1057), .A2(n1026), .A3(n1058), .A4(n1059), .ZN(n1056) );
INV_X1 U753 ( .A(n1060), .ZN(n1059) );
NOR2_X1 U754 ( .A1(n1031), .A2(n1061), .ZN(n1055) );
NAND2_X1 U755 ( .A1(n1062), .A2(n1063), .ZN(n1054) );
NAND2_X1 U756 ( .A1(n1064), .A2(G469), .ZN(n1063) );
INV_X1 U757 ( .A(n1065), .ZN(n1062) );
XOR2_X1 U758 ( .A(G472), .B(n1066), .Z(n1053) );
NOR2_X1 U759 ( .A1(KEYINPUT6), .A2(n1067), .ZN(n1066) );
XNOR2_X1 U760 ( .A(KEYINPUT38), .B(n1068), .ZN(n1067) );
XOR2_X1 U761 ( .A(n1069), .B(n1070), .Z(G72) );
NOR2_X1 U762 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U763 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NAND3_X1 U764 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1069) );
NAND3_X1 U765 ( .A1(n1078), .A2(n1072), .A3(n1079), .ZN(n1077) );
NAND2_X1 U766 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U767 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U768 ( .A1(KEYINPUT3), .A2(n1082), .ZN(n1076) );
NAND3_X1 U769 ( .A1(n1084), .A2(n1080), .A3(n1085), .ZN(n1075) );
INV_X1 U770 ( .A(n1082), .ZN(n1085) );
NAND2_X1 U771 ( .A1(n1086), .A2(n1087), .ZN(n1082) );
NAND2_X1 U772 ( .A1(G953), .A2(n1074), .ZN(n1087) );
XOR2_X1 U773 ( .A(n1088), .B(n1089), .Z(n1086) );
XOR2_X1 U774 ( .A(KEYINPUT18), .B(n1090), .Z(n1089) );
NOR2_X1 U775 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U776 ( .A(n1093), .B(KEYINPUT26), .Z(n1092) );
NAND2_X1 U777 ( .A1(G140), .A2(n1094), .ZN(n1093) );
NOR2_X1 U778 ( .A1(G140), .A2(n1094), .ZN(n1091) );
XOR2_X1 U779 ( .A(KEYINPUT60), .B(G125), .Z(n1094) );
INV_X1 U780 ( .A(KEYINPUT3), .ZN(n1080) );
NAND2_X1 U781 ( .A1(n1083), .A2(n1078), .ZN(n1084) );
NAND2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(n1078) );
INV_X1 U783 ( .A(KEYINPUT58), .ZN(n1083) );
XOR2_X1 U784 ( .A(n1097), .B(n1098), .Z(G69) );
XOR2_X1 U785 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U786 ( .A1(n1101), .A2(n1072), .ZN(n1100) );
NOR2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND3_X1 U788 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1099) );
XOR2_X1 U789 ( .A(KEYINPUT5), .B(n1107), .Z(n1106) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U791 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
NAND2_X1 U792 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U793 ( .A1(G953), .A2(n1103), .ZN(n1104) );
NAND2_X1 U794 ( .A1(n1072), .A2(n1112), .ZN(n1097) );
NAND2_X1 U795 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XNOR2_X1 U796 ( .A(KEYINPUT45), .B(n1115), .ZN(n1114) );
NOR2_X1 U797 ( .A1(n1116), .A2(n1117), .ZN(G66) );
XNOR2_X1 U798 ( .A(n1118), .B(n1119), .ZN(n1117) );
XOR2_X1 U799 ( .A(KEYINPUT51), .B(n1120), .Z(n1119) );
NOR3_X1 U800 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1120) );
XOR2_X1 U801 ( .A(KEYINPUT44), .B(G217), .Z(n1121) );
NOR2_X1 U802 ( .A1(n1116), .A2(n1124), .ZN(G63) );
XOR2_X1 U803 ( .A(n1125), .B(n1126), .Z(n1124) );
AND2_X1 U804 ( .A1(G478), .A2(n1127), .ZN(n1125) );
NOR2_X1 U805 ( .A1(n1116), .A2(n1128), .ZN(G60) );
XOR2_X1 U806 ( .A(n1129), .B(n1130), .Z(n1128) );
AND2_X1 U807 ( .A1(G475), .A2(n1127), .ZN(n1129) );
XNOR2_X1 U808 ( .A(G104), .B(n1115), .ZN(G6) );
NOR2_X1 U809 ( .A1(n1116), .A2(n1131), .ZN(G57) );
XOR2_X1 U810 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U812 ( .A(n1136), .B(n1137), .Z(n1132) );
NOR2_X1 U813 ( .A1(KEYINPUT62), .A2(n1138), .ZN(n1137) );
XOR2_X1 U814 ( .A(n1139), .B(n1140), .Z(n1136) );
AND2_X1 U815 ( .A1(G472), .A2(n1127), .ZN(n1140) );
NOR2_X1 U816 ( .A1(n1116), .A2(n1141), .ZN(G54) );
XOR2_X1 U817 ( .A(n1142), .B(n1143), .Z(n1141) );
XNOR2_X1 U818 ( .A(n1144), .B(n1145), .ZN(n1143) );
NOR2_X1 U819 ( .A1(KEYINPUT36), .A2(n1146), .ZN(n1145) );
XOR2_X1 U820 ( .A(KEYINPUT16), .B(n1147), .Z(n1146) );
NAND3_X1 U821 ( .A1(n1127), .A2(G469), .A3(KEYINPUT63), .ZN(n1144) );
NOR2_X1 U822 ( .A1(n1116), .A2(n1148), .ZN(G51) );
NOR3_X1 U823 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1148) );
NOR2_X1 U824 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NOR2_X1 U825 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
INV_X1 U826 ( .A(KEYINPUT21), .ZN(n1155) );
XOR2_X1 U827 ( .A(n1156), .B(KEYINPUT13), .Z(n1154) );
AND3_X1 U828 ( .A1(n1153), .A2(n1156), .A3(KEYINPUT21), .ZN(n1150) );
XOR2_X1 U829 ( .A(n1157), .B(n1158), .Z(n1153) );
XNOR2_X1 U830 ( .A(n1159), .B(n1160), .ZN(n1158) );
NAND2_X1 U831 ( .A1(KEYINPUT25), .A2(n1161), .ZN(n1159) );
XOR2_X1 U832 ( .A(G125), .B(n1162), .Z(n1161) );
NOR2_X1 U833 ( .A1(n1163), .A2(KEYINPUT7), .ZN(n1162) );
INV_X1 U834 ( .A(n1139), .ZN(n1163) );
XNOR2_X1 U835 ( .A(n1164), .B(KEYINPUT37), .ZN(n1157) );
NOR2_X1 U836 ( .A1(KEYINPUT21), .A2(n1156), .ZN(n1149) );
NAND2_X1 U837 ( .A1(n1127), .A2(G210), .ZN(n1156) );
INV_X1 U838 ( .A(n1123), .ZN(n1127) );
NAND2_X1 U839 ( .A1(G902), .A2(n1020), .ZN(n1123) );
NAND4_X1 U840 ( .A1(n1165), .A2(n1113), .A3(n1095), .A4(n1115), .ZN(n1020) );
NAND2_X1 U841 ( .A1(n1048), .A2(n1166), .ZN(n1115) );
AND4_X1 U842 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1095) );
NOR3_X1 U843 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1170) );
NAND2_X1 U844 ( .A1(n1174), .A2(n1175), .ZN(n1169) );
NAND2_X1 U845 ( .A1(n1037), .A2(n1176), .ZN(n1168) );
NAND3_X1 U846 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1176) );
OR2_X1 U847 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
OR4_X1 U848 ( .A1(n1182), .A2(n1183), .A3(n1051), .A4(KEYINPUT46), .ZN(n1178) );
OR2_X1 U849 ( .A1(n1184), .A2(n1185), .ZN(n1177) );
NAND2_X1 U850 ( .A1(KEYINPUT46), .A2(n1186), .ZN(n1167) );
AND4_X1 U851 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1113) );
NOR4_X1 U852 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1015), .ZN(n1190) );
AND2_X1 U853 ( .A1(n1047), .A2(n1166), .ZN(n1015) );
NOR4_X1 U854 ( .A1(n1194), .A2(n1195), .A3(n1035), .A4(n1196), .ZN(n1166) );
NAND3_X1 U855 ( .A1(n1197), .A2(n1047), .A3(n1043), .ZN(n1189) );
INV_X1 U856 ( .A(n1181), .ZN(n1047) );
NAND4_X1 U857 ( .A1(n1198), .A2(n1037), .A3(n1183), .A4(n1061), .ZN(n1187) );
XOR2_X1 U858 ( .A(n1096), .B(KEYINPUT59), .Z(n1165) );
NAND2_X1 U859 ( .A1(n1199), .A2(n1200), .ZN(n1096) );
XOR2_X1 U860 ( .A(KEYINPUT31), .B(n1037), .Z(n1200) );
NOR2_X1 U861 ( .A1(n1072), .A2(G952), .ZN(n1116) );
XOR2_X1 U862 ( .A(G146), .B(n1186), .Z(G48) );
NOR3_X1 U863 ( .A1(n1201), .A2(n1195), .A3(n1180), .ZN(n1186) );
XOR2_X1 U864 ( .A(G143), .B(n1202), .Z(G45) );
NOR3_X1 U865 ( .A1(n1203), .A2(n1195), .A3(n1184), .ZN(n1202) );
XNOR2_X1 U866 ( .A(KEYINPUT35), .B(n1185), .ZN(n1203) );
XOR2_X1 U867 ( .A(n1204), .B(n1205), .Z(G42) );
NAND2_X1 U868 ( .A1(KEYINPUT9), .A2(G140), .ZN(n1205) );
NAND2_X1 U869 ( .A1(n1175), .A2(n1206), .ZN(n1204) );
XOR2_X1 U870 ( .A(KEYINPUT1), .B(n1174), .Z(n1206) );
NOR3_X1 U871 ( .A1(n1045), .A2(n1194), .A3(n1182), .ZN(n1174) );
XOR2_X1 U872 ( .A(G137), .B(n1171), .Z(G39) );
NOR3_X1 U873 ( .A1(n1041), .A2(n1031), .A3(n1180), .ZN(n1171) );
XOR2_X1 U874 ( .A(G134), .B(n1173), .Z(G36) );
NOR3_X1 U875 ( .A1(n1184), .A2(n1181), .A3(n1041), .ZN(n1173) );
XOR2_X1 U876 ( .A(G131), .B(n1172), .Z(G33) );
NOR3_X1 U877 ( .A1(n1184), .A2(n1201), .A3(n1041), .ZN(n1172) );
INV_X1 U878 ( .A(n1175), .ZN(n1041) );
NOR2_X1 U879 ( .A1(n1038), .A2(n1058), .ZN(n1175) );
INV_X1 U880 ( .A(n1039), .ZN(n1058) );
NAND3_X1 U881 ( .A1(n1051), .A2(n1207), .A3(n1043), .ZN(n1184) );
XOR2_X1 U882 ( .A(G128), .B(n1208), .Z(G30) );
NOR2_X1 U883 ( .A1(n1195), .A2(n1209), .ZN(n1208) );
XOR2_X1 U884 ( .A(KEYINPUT50), .B(n1210), .Z(n1209) );
NOR2_X1 U885 ( .A1(n1181), .A2(n1180), .ZN(n1210) );
NAND4_X1 U886 ( .A1(n1051), .A2(n1045), .A3(n1061), .A4(n1207), .ZN(n1180) );
INV_X1 U887 ( .A(n1194), .ZN(n1051) );
XOR2_X1 U888 ( .A(n1211), .B(n1188), .Z(G3) );
NAND3_X1 U889 ( .A1(n1043), .A2(n1037), .A3(n1198), .ZN(n1188) );
XOR2_X1 U890 ( .A(n1212), .B(n1213), .Z(G27) );
NOR2_X1 U891 ( .A1(n1195), .A2(n1214), .ZN(n1213) );
XOR2_X1 U892 ( .A(KEYINPUT41), .B(n1199), .Z(n1214) );
NOR4_X1 U893 ( .A1(n1182), .A2(n1025), .A3(n1045), .A4(n1026), .ZN(n1199) );
NAND3_X1 U894 ( .A1(n1061), .A2(n1207), .A3(n1048), .ZN(n1182) );
NAND2_X1 U895 ( .A1(n1022), .A2(n1215), .ZN(n1207) );
NAND4_X1 U896 ( .A1(G953), .A2(G902), .A3(n1216), .A4(n1074), .ZN(n1215) );
INV_X1 U897 ( .A(G900), .ZN(n1074) );
NAND2_X1 U898 ( .A1(KEYINPUT33), .A2(n1217), .ZN(n1212) );
INV_X1 U899 ( .A(G125), .ZN(n1217) );
XOR2_X1 U900 ( .A(G122), .B(n1193), .Z(G24) );
NOR3_X1 U901 ( .A1(n1218), .A2(n1035), .A3(n1185), .ZN(n1193) );
NAND2_X1 U902 ( .A1(n1219), .A2(n1220), .ZN(n1185) );
NAND2_X1 U903 ( .A1(n1044), .A2(n1183), .ZN(n1035) );
XOR2_X1 U904 ( .A(G119), .B(n1192), .Z(G21) );
NOR4_X1 U905 ( .A1(n1218), .A2(n1031), .A3(n1183), .A4(n1044), .ZN(n1192) );
XOR2_X1 U906 ( .A(G116), .B(n1221), .Z(G18) );
NOR3_X1 U907 ( .A1(n1222), .A2(n1181), .A3(n1218), .ZN(n1221) );
INV_X1 U908 ( .A(n1197), .ZN(n1218) );
NAND2_X1 U909 ( .A1(n1219), .A2(n1223), .ZN(n1181) );
XOR2_X1 U910 ( .A(n1224), .B(KEYINPUT28), .Z(n1219) );
XOR2_X1 U911 ( .A(KEYINPUT54), .B(n1043), .Z(n1222) );
XOR2_X1 U912 ( .A(G113), .B(n1191), .Z(G15) );
AND3_X1 U913 ( .A1(n1197), .A2(n1048), .A3(n1043), .ZN(n1191) );
NOR2_X1 U914 ( .A1(n1061), .A2(n1183), .ZN(n1043) );
INV_X1 U915 ( .A(n1201), .ZN(n1048) );
NAND2_X1 U916 ( .A1(n1224), .A2(n1220), .ZN(n1201) );
INV_X1 U917 ( .A(n1223), .ZN(n1220) );
NOR4_X1 U918 ( .A1(n1025), .A2(n1195), .A3(n1196), .A4(n1026), .ZN(n1197) );
INV_X1 U919 ( .A(n1052), .ZN(n1026) );
XOR2_X1 U920 ( .A(n1225), .B(n1226), .Z(G12) );
NAND4_X1 U921 ( .A1(n1183), .A2(n1198), .A3(n1227), .A4(n1061), .ZN(n1226) );
INV_X1 U922 ( .A(n1044), .ZN(n1061) );
XOR2_X1 U923 ( .A(n1228), .B(n1229), .Z(n1044) );
NOR2_X1 U924 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U925 ( .A(KEYINPUT2), .B(n1122), .Z(n1231) );
INV_X1 U926 ( .A(n1232), .ZN(n1122) );
NAND2_X1 U927 ( .A1(n1118), .A2(n1233), .ZN(n1228) );
XNOR2_X1 U928 ( .A(n1234), .B(n1235), .ZN(n1118) );
XOR2_X1 U929 ( .A(G119), .B(n1236), .Z(n1235) );
XOR2_X1 U930 ( .A(G137), .B(G128), .Z(n1236) );
XOR2_X1 U931 ( .A(n1237), .B(n1238), .Z(n1234) );
XOR2_X1 U932 ( .A(n1239), .B(n1240), .Z(n1238) );
AND3_X1 U933 ( .A1(G221), .A2(n1072), .A3(G234), .ZN(n1239) );
XOR2_X1 U934 ( .A(KEYINPUT49), .B(n1037), .Z(n1227) );
INV_X1 U935 ( .A(n1195), .ZN(n1037) );
NAND2_X1 U936 ( .A1(n1039), .A2(n1038), .ZN(n1195) );
NAND2_X1 U937 ( .A1(n1241), .A2(n1060), .ZN(n1038) );
NAND3_X1 U938 ( .A1(n1242), .A2(n1243), .A3(G210), .ZN(n1060) );
XNOR2_X1 U939 ( .A(n1057), .B(KEYINPUT12), .ZN(n1241) );
NOR2_X1 U940 ( .A1(n1243), .A2(n1244), .ZN(n1057) );
AND2_X1 U941 ( .A1(G237), .A2(G210), .ZN(n1244) );
NAND3_X1 U942 ( .A1(n1245), .A2(n1233), .A3(n1246), .ZN(n1243) );
XOR2_X1 U943 ( .A(n1247), .B(KEYINPUT15), .Z(n1246) );
NAND2_X1 U944 ( .A1(n1248), .A2(n1160), .ZN(n1247) );
OR2_X1 U945 ( .A1(n1160), .A2(n1248), .ZN(n1245) );
XNOR2_X1 U946 ( .A(n1249), .B(n1250), .ZN(n1248) );
XOR2_X1 U947 ( .A(KEYINPUT24), .B(G125), .Z(n1250) );
XOR2_X1 U948 ( .A(n1139), .B(n1164), .Z(n1249) );
NOR2_X1 U949 ( .A1(n1102), .A2(G953), .ZN(n1164) );
INV_X1 U950 ( .A(G224), .ZN(n1102) );
XNOR2_X1 U951 ( .A(n1251), .B(n1252), .ZN(n1160) );
NOR2_X1 U952 ( .A1(KEYINPUT48), .A2(n1108), .ZN(n1252) );
XOR2_X1 U953 ( .A(n1253), .B(KEYINPUT30), .Z(n1108) );
NAND3_X1 U954 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1253) );
OR2_X1 U955 ( .A1(n1225), .A2(KEYINPUT4), .ZN(n1256) );
NAND3_X1 U956 ( .A1(KEYINPUT4), .A2(n1257), .A3(n1258), .ZN(n1255) );
OR2_X1 U957 ( .A1(n1258), .A2(n1257), .ZN(n1254) );
NOR2_X1 U958 ( .A1(G110), .A2(KEYINPUT23), .ZN(n1257) );
XNOR2_X1 U959 ( .A(n1259), .B(KEYINPUT42), .ZN(n1258) );
INV_X1 U960 ( .A(G122), .ZN(n1259) );
NAND2_X1 U961 ( .A1(n1260), .A2(n1111), .ZN(n1251) );
NAND2_X1 U962 ( .A1(n1261), .A2(n1262), .ZN(n1111) );
XOR2_X1 U963 ( .A(n1263), .B(n1264), .Z(n1261) );
XOR2_X1 U964 ( .A(n1110), .B(KEYINPUT56), .Z(n1260) );
NAND2_X1 U965 ( .A1(n1265), .A2(n1266), .ZN(n1110) );
XNOR2_X1 U966 ( .A(n1264), .B(n1263), .ZN(n1265) );
NOR2_X1 U967 ( .A1(KEYINPUT27), .A2(G113), .ZN(n1263) );
NAND2_X1 U968 ( .A1(G214), .A2(n1242), .ZN(n1039) );
NAND2_X1 U969 ( .A1(n1267), .A2(n1233), .ZN(n1242) );
NOR3_X1 U970 ( .A1(n1194), .A2(n1196), .A3(n1031), .ZN(n1198) );
NAND2_X1 U971 ( .A1(n1223), .A2(n1224), .ZN(n1031) );
XOR2_X1 U972 ( .A(n1268), .B(G478), .Z(n1224) );
OR2_X1 U973 ( .A1(n1126), .A2(G902), .ZN(n1268) );
XNOR2_X1 U974 ( .A(n1269), .B(n1270), .ZN(n1126) );
XOR2_X1 U975 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U976 ( .A(G122), .B(G107), .Z(n1272) );
XOR2_X1 U977 ( .A(G134), .B(G128), .Z(n1271) );
XNOR2_X1 U978 ( .A(n1273), .B(n1274), .ZN(n1269) );
XOR2_X1 U979 ( .A(n1275), .B(n1276), .Z(n1274) );
NAND2_X1 U980 ( .A1(KEYINPUT11), .A2(G143), .ZN(n1276) );
NAND3_X1 U981 ( .A1(G234), .A2(n1072), .A3(n1277), .ZN(n1275) );
XOR2_X1 U982 ( .A(n1230), .B(KEYINPUT39), .Z(n1277) );
INV_X1 U983 ( .A(G217), .ZN(n1230) );
XOR2_X1 U984 ( .A(n1278), .B(G475), .Z(n1223) );
OR2_X1 U985 ( .A1(n1130), .A2(G902), .ZN(n1278) );
XNOR2_X1 U986 ( .A(n1279), .B(n1280), .ZN(n1130) );
NOR2_X1 U987 ( .A1(KEYINPUT34), .A2(n1281), .ZN(n1280) );
XNOR2_X1 U988 ( .A(G104), .B(n1282), .ZN(n1281) );
XOR2_X1 U989 ( .A(G122), .B(G113), .Z(n1282) );
NAND3_X1 U990 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1279) );
NAND2_X1 U991 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND2_X1 U992 ( .A1(KEYINPUT17), .A2(n1288), .ZN(n1287) );
XOR2_X1 U993 ( .A(G140), .B(n1289), .Z(n1286) );
OR2_X1 U994 ( .A1(n1288), .A2(KEYINPUT32), .ZN(n1284) );
NAND4_X1 U995 ( .A1(n1290), .A2(n1288), .A3(KEYINPUT17), .A4(KEYINPUT32), .ZN(n1283) );
XNOR2_X1 U996 ( .A(n1291), .B(G131), .ZN(n1288) );
NAND2_X1 U997 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND4_X1 U998 ( .A1(G214), .A2(G143), .A3(n1267), .A4(n1072), .ZN(n1293) );
XOR2_X1 U999 ( .A(n1294), .B(KEYINPUT14), .Z(n1292) );
NAND2_X1 U1000 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
NAND3_X1 U1001 ( .A1(n1267), .A2(n1072), .A3(G214), .ZN(n1296) );
XOR2_X1 U1002 ( .A(G140), .B(n1237), .Z(n1290) );
INV_X1 U1003 ( .A(n1289), .ZN(n1237) );
XOR2_X1 U1004 ( .A(G146), .B(G125), .Z(n1289) );
AND2_X1 U1005 ( .A1(n1022), .A2(n1297), .ZN(n1196) );
NAND4_X1 U1006 ( .A1(n1298), .A2(G953), .A3(G902), .A4(n1103), .ZN(n1297) );
INV_X1 U1007 ( .A(G898), .ZN(n1103) );
XOR2_X1 U1008 ( .A(n1216), .B(KEYINPUT43), .Z(n1298) );
NAND3_X1 U1009 ( .A1(n1216), .A2(n1072), .A3(G952), .ZN(n1022) );
NAND2_X1 U1010 ( .A1(G237), .A2(G234), .ZN(n1216) );
NAND2_X1 U1011 ( .A1(n1052), .A2(n1025), .ZN(n1194) );
NAND3_X1 U1012 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1025) );
XOR2_X1 U1013 ( .A(n1302), .B(KEYINPUT19), .Z(n1301) );
NAND2_X1 U1014 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND3_X1 U1015 ( .A1(G469), .A2(n1305), .A3(n1306), .ZN(n1304) );
INV_X1 U1016 ( .A(KEYINPUT0), .ZN(n1306) );
NAND2_X1 U1017 ( .A1(n1065), .A2(KEYINPUT0), .ZN(n1303) );
OR3_X1 U1018 ( .A1(n1305), .A2(G469), .A3(KEYINPUT47), .ZN(n1300) );
NAND2_X1 U1019 ( .A1(KEYINPUT47), .A2(n1065), .ZN(n1299) );
NOR2_X1 U1020 ( .A1(n1064), .A2(G469), .ZN(n1065) );
INV_X1 U1021 ( .A(n1305), .ZN(n1064) );
NAND2_X1 U1022 ( .A1(n1307), .A2(n1233), .ZN(n1305) );
XOR2_X1 U1023 ( .A(n1147), .B(n1308), .Z(n1307) );
INV_X1 U1024 ( .A(n1142), .ZN(n1308) );
XOR2_X1 U1025 ( .A(n1088), .B(n1262), .Z(n1142) );
INV_X1 U1026 ( .A(n1266), .ZN(n1262) );
XOR2_X1 U1027 ( .A(n1211), .B(n1309), .Z(n1266) );
XOR2_X1 U1028 ( .A(G107), .B(G104), .Z(n1309) );
INV_X1 U1029 ( .A(G101), .ZN(n1211) );
XNOR2_X1 U1030 ( .A(n1134), .B(n1310), .ZN(n1088) );
NOR2_X1 U1031 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U1032 ( .A(n1313), .B(KEYINPUT22), .Z(n1312) );
NAND2_X1 U1033 ( .A1(G128), .A2(n1314), .ZN(n1313) );
NOR2_X1 U1034 ( .A1(G128), .A2(n1314), .ZN(n1311) );
NAND2_X1 U1035 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND2_X1 U1036 ( .A1(G146), .A2(n1295), .ZN(n1316) );
XOR2_X1 U1037 ( .A(n1317), .B(KEYINPUT40), .Z(n1315) );
OR2_X1 U1038 ( .A1(n1295), .A2(G146), .ZN(n1317) );
AND2_X1 U1039 ( .A1(n1318), .A2(n1319), .ZN(n1147) );
NAND2_X1 U1040 ( .A1(n1240), .A2(n1320), .ZN(n1319) );
NAND2_X1 U1041 ( .A1(G227), .A2(n1072), .ZN(n1320) );
OR3_X1 U1042 ( .A1(n1073), .A2(G953), .A3(n1240), .ZN(n1318) );
XNOR2_X1 U1043 ( .A(n1225), .B(G140), .ZN(n1240) );
INV_X1 U1044 ( .A(G227), .ZN(n1073) );
NAND2_X1 U1045 ( .A1(G221), .A2(n1232), .ZN(n1052) );
NAND2_X1 U1046 ( .A1(G234), .A2(n1321), .ZN(n1232) );
XOR2_X1 U1047 ( .A(KEYINPUT10), .B(G902), .Z(n1321) );
INV_X1 U1048 ( .A(n1045), .ZN(n1183) );
XNOR2_X1 U1049 ( .A(n1068), .B(G472), .ZN(n1045) );
NAND2_X1 U1050 ( .A1(n1322), .A2(n1233), .ZN(n1068) );
INV_X1 U1051 ( .A(G902), .ZN(n1233) );
XOR2_X1 U1052 ( .A(n1323), .B(n1324), .Z(n1322) );
XNOR2_X1 U1053 ( .A(n1138), .B(n1135), .ZN(n1324) );
XOR2_X1 U1054 ( .A(G101), .B(n1325), .Z(n1135) );
AND3_X1 U1055 ( .A1(G210), .A2(n1072), .A3(n1267), .ZN(n1325) );
INV_X1 U1056 ( .A(G237), .ZN(n1267) );
INV_X1 U1057 ( .A(G953), .ZN(n1072) );
XNOR2_X1 U1058 ( .A(n1326), .B(n1264), .ZN(n1138) );
XOR2_X1 U1059 ( .A(G119), .B(n1273), .Z(n1264) );
XOR2_X1 U1060 ( .A(G116), .B(KEYINPUT20), .Z(n1273) );
NAND2_X1 U1061 ( .A1(KEYINPUT29), .A2(n1327), .ZN(n1326) );
INV_X1 U1062 ( .A(G113), .ZN(n1327) );
XOR2_X1 U1063 ( .A(n1328), .B(KEYINPUT8), .Z(n1323) );
NAND2_X1 U1064 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
NAND2_X1 U1065 ( .A1(n1331), .A2(n1139), .ZN(n1330) );
XOR2_X1 U1066 ( .A(KEYINPUT61), .B(n1332), .Z(n1329) );
NOR2_X1 U1067 ( .A1(n1139), .A2(n1331), .ZN(n1332) );
XOR2_X1 U1068 ( .A(KEYINPUT55), .B(n1134), .Z(n1331) );
XNOR2_X1 U1069 ( .A(n1333), .B(n1334), .ZN(n1134) );
XOR2_X1 U1070 ( .A(KEYINPUT53), .B(G137), .Z(n1334) );
XOR2_X1 U1071 ( .A(G131), .B(n1335), .Z(n1333) );
INV_X1 U1072 ( .A(G134), .ZN(n1335) );
NAND2_X1 U1073 ( .A1(n1336), .A2(n1337), .ZN(n1139) );
NAND2_X1 U1074 ( .A1(n1338), .A2(G128), .ZN(n1337) );
XOR2_X1 U1075 ( .A(KEYINPUT57), .B(n1339), .Z(n1336) );
NOR2_X1 U1076 ( .A1(G128), .A2(n1338), .ZN(n1339) );
XOR2_X1 U1077 ( .A(n1340), .B(G146), .Z(n1338) );
NAND2_X1 U1078 ( .A1(KEYINPUT52), .A2(n1295), .ZN(n1340) );
INV_X1 U1079 ( .A(G143), .ZN(n1295) );
INV_X1 U1080 ( .A(G110), .ZN(n1225) );
endmodule


