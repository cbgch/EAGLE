//Key = 1001100001011101000100010011010110000111101001001001110110000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355;

XNOR2_X1 U757 ( .A(n1041), .B(n1042), .ZN(G9) );
NOR3_X1 U758 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
XNOR2_X1 U759 ( .A(KEYINPUT0), .B(n1046), .ZN(n1043) );
NOR2_X1 U760 ( .A1(n1047), .A2(n1048), .ZN(G75) );
NOR4_X1 U761 ( .A1(n1049), .A2(n1050), .A3(G953), .A4(n1051), .ZN(n1048) );
NOR3_X1 U762 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1050) );
NOR2_X1 U763 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR3_X1 U764 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1055) );
NAND3_X1 U765 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1049) );
NAND2_X1 U766 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NAND3_X1 U767 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
XOR2_X1 U768 ( .A(n1068), .B(KEYINPUT30), .Z(n1067) );
NAND4_X1 U769 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1068) );
NAND4_X1 U770 ( .A1(n1073), .A2(n1074), .A3(n1069), .A4(n1075), .ZN(n1066) );
NOR2_X1 U771 ( .A1(n1054), .A2(n1076), .ZN(n1075) );
NAND2_X1 U772 ( .A1(n1077), .A2(n1078), .ZN(n1074) );
OR2_X1 U773 ( .A1(n1078), .A2(n1072), .ZN(n1073) );
NAND2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1065) );
NAND2_X1 U775 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
OR2_X1 U776 ( .A1(n1046), .A2(KEYINPUT16), .ZN(n1082) );
XOR2_X1 U777 ( .A(n1083), .B(KEYINPUT58), .Z(n1081) );
NAND2_X1 U778 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U779 ( .A1(KEYINPUT16), .A2(n1086), .ZN(n1060) );
NAND3_X1 U780 ( .A1(n1063), .A2(n1087), .A3(n1079), .ZN(n1086) );
INV_X1 U781 ( .A(n1052), .ZN(n1079) );
NAND4_X1 U782 ( .A1(n1069), .A2(n1072), .A3(n1088), .A4(n1078), .ZN(n1052) );
INV_X1 U783 ( .A(n1089), .ZN(n1069) );
NOR3_X1 U784 ( .A1(n1051), .A2(G953), .A3(G952), .ZN(n1047) );
AND4_X1 U785 ( .A1(n1090), .A2(n1057), .A3(n1072), .A4(n1091), .ZN(n1051) );
NOR4_X1 U786 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1091) );
XNOR2_X1 U787 ( .A(KEYINPUT34), .B(n1088), .ZN(n1095) );
XOR2_X1 U788 ( .A(n1096), .B(n1097), .Z(n1094) );
XNOR2_X1 U789 ( .A(n1098), .B(KEYINPUT56), .ZN(n1097) );
NAND2_X1 U790 ( .A1(KEYINPUT53), .A2(n1099), .ZN(n1096) );
AND2_X1 U791 ( .A1(n1054), .A2(KEYINPUT19), .ZN(n1093) );
NOR2_X1 U792 ( .A1(KEYINPUT19), .A2(n1087), .ZN(n1092) );
XOR2_X1 U793 ( .A(KEYINPUT43), .B(n1100), .Z(n1090) );
NOR2_X1 U794 ( .A1(n1058), .A2(n1101), .ZN(n1100) );
XNOR2_X1 U795 ( .A(n1059), .B(KEYINPUT13), .ZN(n1101) );
INV_X1 U796 ( .A(n1102), .ZN(n1058) );
XOR2_X1 U797 ( .A(n1103), .B(n1104), .Z(G72) );
XOR2_X1 U798 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U799 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U800 ( .A(n1109), .B(n1110), .ZN(n1108) );
XOR2_X1 U801 ( .A(n1111), .B(n1112), .Z(n1110) );
NAND2_X1 U802 ( .A1(n1113), .A2(KEYINPUT23), .ZN(n1112) );
XNOR2_X1 U803 ( .A(n1114), .B(KEYINPUT33), .ZN(n1113) );
NOR2_X1 U804 ( .A1(G900), .A2(n1115), .ZN(n1107) );
NAND2_X1 U805 ( .A1(n1115), .A2(n1116), .ZN(n1105) );
NAND2_X1 U806 ( .A1(G953), .A2(n1117), .ZN(n1103) );
NAND2_X1 U807 ( .A1(G900), .A2(G227), .ZN(n1117) );
XOR2_X1 U808 ( .A(n1118), .B(n1119), .Z(G69) );
XOR2_X1 U809 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U810 ( .A1(G953), .A2(n1122), .ZN(n1121) );
NAND2_X1 U811 ( .A1(G898), .A2(G224), .ZN(n1122) );
NAND2_X1 U812 ( .A1(n1123), .A2(n1124), .ZN(n1120) );
XNOR2_X1 U813 ( .A(G953), .B(KEYINPUT47), .ZN(n1123) );
NOR2_X1 U814 ( .A1(n1125), .A2(n1126), .ZN(n1118) );
NOR2_X1 U815 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XNOR2_X1 U816 ( .A(n1129), .B(n1130), .ZN(n1128) );
XOR2_X1 U817 ( .A(n1131), .B(KEYINPUT39), .Z(n1130) );
NAND2_X1 U818 ( .A1(n1132), .A2(n1098), .ZN(n1131) );
NOR2_X1 U819 ( .A1(n1127), .A2(n1133), .ZN(G63) );
XOR2_X1 U820 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U821 ( .A1(n1136), .A2(KEYINPUT62), .ZN(n1134) );
AND2_X1 U822 ( .A1(G478), .A2(n1132), .ZN(n1136) );
NOR2_X1 U823 ( .A1(n1127), .A2(n1137), .ZN(G60) );
XOR2_X1 U824 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U825 ( .A1(n1132), .A2(G475), .ZN(n1138) );
XOR2_X1 U826 ( .A(G104), .B(n1140), .Z(G6) );
NOR3_X1 U827 ( .A1(n1141), .A2(n1044), .A3(n1142), .ZN(n1140) );
XNOR2_X1 U828 ( .A(KEYINPUT11), .B(n1046), .ZN(n1141) );
NOR3_X1 U829 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(G57) );
AND3_X1 U830 ( .A1(KEYINPUT57), .A2(G953), .A3(G952), .ZN(n1145) );
NOR2_X1 U831 ( .A1(KEYINPUT57), .A2(n1146), .ZN(n1144) );
INV_X1 U832 ( .A(n1127), .ZN(n1146) );
XOR2_X1 U833 ( .A(n1147), .B(n1148), .Z(n1143) );
XOR2_X1 U834 ( .A(n1149), .B(n1150), .Z(n1148) );
NAND2_X1 U835 ( .A1(n1132), .A2(G472), .ZN(n1150) );
NAND2_X1 U836 ( .A1(KEYINPUT52), .A2(n1151), .ZN(n1149) );
XOR2_X1 U837 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U838 ( .A1(G101), .A2(KEYINPUT22), .ZN(n1153) );
NOR2_X1 U839 ( .A1(n1127), .A2(n1154), .ZN(G54) );
XOR2_X1 U840 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U841 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NOR2_X1 U842 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U843 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U844 ( .A(KEYINPUT35), .B(KEYINPUT2), .ZN(n1162) );
NOR2_X1 U845 ( .A1(n1163), .A2(n1161), .ZN(n1157) );
XOR2_X1 U846 ( .A(n1164), .B(G140), .Z(n1161) );
NAND2_X1 U847 ( .A1(KEYINPUT26), .A2(n1165), .ZN(n1164) );
INV_X1 U848 ( .A(n1159), .ZN(n1163) );
XNOR2_X1 U849 ( .A(n1166), .B(KEYINPUT9), .ZN(n1159) );
XOR2_X1 U850 ( .A(n1167), .B(n1168), .Z(n1155) );
NAND2_X1 U851 ( .A1(n1132), .A2(G469), .ZN(n1167) );
NOR2_X1 U852 ( .A1(n1127), .A2(n1169), .ZN(G51) );
NOR2_X1 U853 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U854 ( .A(KEYINPUT14), .B(n1172), .Z(n1171) );
NOR2_X1 U855 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
AND2_X1 U856 ( .A1(n1174), .A2(n1173), .ZN(n1170) );
XOR2_X1 U857 ( .A(n1175), .B(n1176), .Z(n1173) );
XOR2_X1 U858 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U859 ( .A(n1179), .B(KEYINPUT45), .Z(n1178) );
XNOR2_X1 U860 ( .A(n1180), .B(n1126), .ZN(n1175) );
INV_X1 U861 ( .A(n1181), .ZN(n1126) );
NAND2_X1 U862 ( .A1(KEYINPUT12), .A2(n1182), .ZN(n1180) );
INV_X1 U863 ( .A(G125), .ZN(n1182) );
NAND2_X1 U864 ( .A1(n1132), .A2(G210), .ZN(n1174) );
NOR2_X1 U865 ( .A1(n1183), .A2(n1062), .ZN(n1132) );
NOR2_X1 U866 ( .A1(n1124), .A2(n1116), .ZN(n1062) );
NAND4_X1 U867 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1116) );
NOR3_X1 U868 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
NOR2_X1 U869 ( .A1(n1077), .A2(n1191), .ZN(n1190) );
NOR2_X1 U870 ( .A1(n1192), .A2(n1193), .ZN(n1189) );
NOR3_X1 U871 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1192) );
NOR3_X1 U872 ( .A1(n1197), .A2(KEYINPUT15), .A3(n1087), .ZN(n1196) );
NOR2_X1 U873 ( .A1(n1045), .A2(n1198), .ZN(n1194) );
AND2_X1 U874 ( .A1(n1199), .A2(KEYINPUT15), .ZN(n1188) );
NAND2_X1 U875 ( .A1(n1056), .A2(n1200), .ZN(n1186) );
XOR2_X1 U876 ( .A(KEYINPUT20), .B(n1201), .Z(n1200) );
NAND4_X1 U877 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1124) );
NOR3_X1 U878 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1205) );
NOR3_X1 U879 ( .A1(n1209), .A2(n1044), .A3(n1054), .ZN(n1208) );
INV_X1 U880 ( .A(n1210), .ZN(n1207) );
NOR2_X1 U881 ( .A1(n1211), .A2(n1046), .ZN(n1206) );
NOR2_X1 U882 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NOR2_X1 U883 ( .A1(n1077), .A2(n1044), .ZN(n1213) );
NOR2_X1 U884 ( .A1(n1214), .A2(n1215), .ZN(n1077) );
NOR3_X1 U885 ( .A1(n1216), .A2(n1076), .A3(n1078), .ZN(n1212) );
NOR2_X1 U886 ( .A1(n1115), .A2(G952), .ZN(n1127) );
NAND2_X1 U887 ( .A1(n1217), .A2(n1218), .ZN(G48) );
NAND2_X1 U888 ( .A1(KEYINPUT61), .A2(n1219), .ZN(n1218) );
XOR2_X1 U889 ( .A(n1220), .B(n1221), .Z(n1217) );
NOR2_X1 U890 ( .A1(KEYINPUT61), .A2(n1219), .ZN(n1221) );
XNOR2_X1 U891 ( .A(KEYINPUT55), .B(n1222), .ZN(n1219) );
OR2_X1 U892 ( .A1(n1191), .A2(n1142), .ZN(n1220) );
XNOR2_X1 U893 ( .A(n1223), .B(n1184), .ZN(G45) );
OR3_X1 U894 ( .A1(n1209), .A2(n1224), .A3(n1198), .ZN(n1184) );
NAND2_X1 U895 ( .A1(KEYINPUT42), .A2(n1225), .ZN(n1223) );
XOR2_X1 U896 ( .A(G140), .B(n1199), .Z(G42) );
NOR3_X1 U897 ( .A1(n1193), .A2(n1046), .A3(n1197), .ZN(n1199) );
INV_X1 U898 ( .A(n1087), .ZN(n1046) );
XNOR2_X1 U899 ( .A(G137), .B(n1226), .ZN(G39) );
NAND2_X1 U900 ( .A1(n1063), .A2(n1227), .ZN(n1226) );
XOR2_X1 U901 ( .A(KEYINPUT46), .B(n1195), .Z(n1227) );
AND2_X1 U902 ( .A1(n1228), .A2(n1072), .ZN(n1195) );
XOR2_X1 U903 ( .A(G134), .B(n1229), .Z(G36) );
NOR3_X1 U904 ( .A1(n1198), .A2(n1230), .A3(n1045), .ZN(n1229) );
INV_X1 U905 ( .A(n1215), .ZN(n1045) );
XNOR2_X1 U906 ( .A(n1063), .B(KEYINPUT18), .ZN(n1230) );
INV_X1 U907 ( .A(n1193), .ZN(n1063) );
XNOR2_X1 U908 ( .A(G131), .B(n1185), .ZN(G33) );
OR3_X1 U909 ( .A1(n1198), .A2(n1142), .A3(n1193), .ZN(n1185) );
NAND3_X1 U910 ( .A1(n1102), .A2(n1057), .A3(n1231), .ZN(n1193) );
NAND3_X1 U911 ( .A1(n1087), .A2(n1232), .A3(n1070), .ZN(n1198) );
XNOR2_X1 U912 ( .A(n1233), .B(n1234), .ZN(G30) );
NOR3_X1 U913 ( .A1(n1191), .A2(KEYINPUT28), .A3(n1235), .ZN(n1234) );
XNOR2_X1 U914 ( .A(n1215), .B(KEYINPUT50), .ZN(n1235) );
NAND2_X1 U915 ( .A1(n1228), .A2(n1056), .ZN(n1191) );
AND4_X1 U916 ( .A1(n1236), .A2(n1087), .A3(n1076), .A4(n1232), .ZN(n1228) );
NAND2_X1 U917 ( .A1(n1237), .A2(n1238), .ZN(G3) );
NAND2_X1 U918 ( .A1(G101), .A2(n1210), .ZN(n1238) );
XOR2_X1 U919 ( .A(n1239), .B(KEYINPUT10), .Z(n1237) );
OR2_X1 U920 ( .A1(n1210), .A2(G101), .ZN(n1239) );
NAND3_X1 U921 ( .A1(n1240), .A2(n1087), .A3(n1070), .ZN(n1210) );
NOR2_X1 U922 ( .A1(n1088), .A2(n1236), .ZN(n1070) );
XNOR2_X1 U923 ( .A(G125), .B(n1241), .ZN(G27) );
NAND2_X1 U924 ( .A1(n1201), .A2(n1056), .ZN(n1241) );
NOR2_X1 U925 ( .A1(n1197), .A2(n1054), .ZN(n1201) );
NAND4_X1 U926 ( .A1(n1236), .A2(n1214), .A3(n1088), .A4(n1232), .ZN(n1197) );
NAND2_X1 U927 ( .A1(n1089), .A2(n1242), .ZN(n1232) );
NAND4_X1 U928 ( .A1(G902), .A2(G953), .A3(n1243), .A4(n1244), .ZN(n1242) );
INV_X1 U929 ( .A(G900), .ZN(n1244) );
XOR2_X1 U930 ( .A(n1245), .B(n1246), .Z(G24) );
NOR2_X1 U931 ( .A1(KEYINPUT8), .A2(n1247), .ZN(n1246) );
NOR4_X1 U932 ( .A1(n1248), .A2(n1249), .A3(n1054), .A4(n1209), .ZN(n1245) );
NAND2_X1 U933 ( .A1(n1250), .A2(n1251), .ZN(n1209) );
NOR2_X1 U934 ( .A1(KEYINPUT4), .A2(n1252), .ZN(n1249) );
AND4_X1 U935 ( .A1(n1224), .A2(n1253), .A3(n1078), .A4(n1088), .ZN(n1252) );
AND2_X1 U936 ( .A1(n1044), .A2(KEYINPUT4), .ZN(n1248) );
NAND2_X1 U937 ( .A1(n1254), .A2(n1088), .ZN(n1044) );
NAND2_X1 U938 ( .A1(n1255), .A2(n1256), .ZN(G21) );
NAND2_X1 U939 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XOR2_X1 U940 ( .A(KEYINPUT38), .B(n1259), .Z(n1255) );
NOR2_X1 U941 ( .A1(n1257), .A2(n1258), .ZN(n1259) );
INV_X1 U942 ( .A(n1204), .ZN(n1257) );
NAND4_X1 U943 ( .A1(n1236), .A2(n1240), .A3(n1071), .A4(n1076), .ZN(n1204) );
XNOR2_X1 U944 ( .A(n1202), .B(n1260), .ZN(G18) );
NOR2_X1 U945 ( .A1(KEYINPUT7), .A2(n1261), .ZN(n1260) );
NAND2_X1 U946 ( .A1(n1262), .A2(n1215), .ZN(n1202) );
NOR2_X1 U947 ( .A1(n1250), .A2(n1263), .ZN(n1215) );
XNOR2_X1 U948 ( .A(G113), .B(n1203), .ZN(G15) );
NAND2_X1 U949 ( .A1(n1214), .A2(n1262), .ZN(n1203) );
AND3_X1 U950 ( .A1(n1254), .A2(n1076), .A3(n1071), .ZN(n1262) );
INV_X1 U951 ( .A(n1054), .ZN(n1071) );
NAND2_X1 U952 ( .A1(n1085), .A2(n1264), .ZN(n1054) );
AND3_X1 U953 ( .A1(n1078), .A2(n1253), .A3(n1056), .ZN(n1254) );
INV_X1 U954 ( .A(n1142), .ZN(n1214) );
NAND2_X1 U955 ( .A1(n1263), .A2(n1250), .ZN(n1142) );
INV_X1 U956 ( .A(n1251), .ZN(n1263) );
XNOR2_X1 U957 ( .A(G110), .B(n1265), .ZN(G12) );
NAND4_X1 U958 ( .A1(n1266), .A2(n1240), .A3(n1236), .A4(n1088), .ZN(n1265) );
INV_X1 U959 ( .A(n1076), .ZN(n1088) );
XNOR2_X1 U960 ( .A(n1267), .B(G472), .ZN(n1076) );
NAND2_X1 U961 ( .A1(n1268), .A2(n1183), .ZN(n1267) );
XOR2_X1 U962 ( .A(n1147), .B(n1269), .Z(n1268) );
XNOR2_X1 U963 ( .A(G101), .B(n1270), .ZN(n1269) );
NAND2_X1 U964 ( .A1(KEYINPUT37), .A2(n1152), .ZN(n1270) );
AND3_X1 U965 ( .A1(n1271), .A2(n1115), .A3(G210), .ZN(n1152) );
XNOR2_X1 U966 ( .A(n1272), .B(n1273), .ZN(n1147) );
XNOR2_X1 U967 ( .A(n1274), .B(n1275), .ZN(n1273) );
INV_X1 U968 ( .A(n1114), .ZN(n1274) );
XNOR2_X1 U969 ( .A(n1179), .B(n1261), .ZN(n1272) );
INV_X1 U970 ( .A(G116), .ZN(n1261) );
INV_X1 U971 ( .A(n1078), .ZN(n1236) );
XNOR2_X1 U972 ( .A(n1276), .B(n1277), .ZN(n1078) );
NOR2_X1 U973 ( .A1(n1098), .A2(KEYINPUT17), .ZN(n1277) );
AND2_X1 U974 ( .A1(G217), .A2(n1278), .ZN(n1098) );
XOR2_X1 U975 ( .A(n1099), .B(KEYINPUT49), .Z(n1276) );
NAND2_X1 U976 ( .A1(n1129), .A2(n1183), .ZN(n1099) );
XNOR2_X1 U977 ( .A(n1279), .B(n1280), .ZN(n1129) );
XOR2_X1 U978 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR2_X1 U979 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
INV_X1 U980 ( .A(G221), .ZN(n1284) );
NOR2_X1 U981 ( .A1(KEYINPUT25), .A2(n1285), .ZN(n1281) );
XOR2_X1 U982 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U983 ( .A(n1288), .B(n1289), .Z(n1287) );
NOR2_X1 U984 ( .A1(G110), .A2(KEYINPUT36), .ZN(n1289) );
NOR2_X1 U985 ( .A1(n1290), .A2(n1291), .ZN(n1288) );
XOR2_X1 U986 ( .A(KEYINPUT54), .B(n1292), .Z(n1291) );
NOR2_X1 U987 ( .A1(G119), .A2(n1233), .ZN(n1292) );
NOR2_X1 U988 ( .A1(G128), .A2(n1258), .ZN(n1290) );
INV_X1 U989 ( .A(G119), .ZN(n1258) );
NOR2_X1 U990 ( .A1(KEYINPUT1), .A2(n1293), .ZN(n1286) );
XNOR2_X1 U991 ( .A(n1222), .B(n1109), .ZN(n1293) );
NAND2_X1 U992 ( .A1(KEYINPUT27), .A2(G137), .ZN(n1279) );
INV_X1 U993 ( .A(n1216), .ZN(n1240) );
NAND3_X1 U994 ( .A1(n1056), .A2(n1253), .A3(n1072), .ZN(n1216) );
NOR2_X1 U995 ( .A1(n1251), .A2(n1250), .ZN(n1072) );
XNOR2_X1 U996 ( .A(n1294), .B(G475), .ZN(n1250) );
NAND2_X1 U997 ( .A1(n1139), .A2(n1183), .ZN(n1294) );
XOR2_X1 U998 ( .A(n1295), .B(n1296), .Z(n1139) );
XOR2_X1 U999 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U1000 ( .A(n1299), .B(n1300), .Z(n1298) );
NOR2_X1 U1001 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
XOR2_X1 U1002 ( .A(KEYINPUT63), .B(n1303), .Z(n1302) );
NOR2_X1 U1003 ( .A1(G146), .A2(n1109), .ZN(n1303) );
NOR2_X1 U1004 ( .A1(n1304), .A2(n1222), .ZN(n1301) );
INV_X1 U1005 ( .A(n1109), .ZN(n1304) );
XOR2_X1 U1006 ( .A(G125), .B(G140), .Z(n1109) );
NOR2_X1 U1007 ( .A1(KEYINPUT6), .A2(n1305), .ZN(n1299) );
XOR2_X1 U1008 ( .A(G104), .B(n1306), .Z(n1305) );
XNOR2_X1 U1009 ( .A(n1247), .B(G113), .ZN(n1306) );
NOR4_X1 U1010 ( .A1(KEYINPUT24), .A2(G953), .A3(G237), .A4(n1307), .ZN(n1297) );
INV_X1 U1011 ( .A(G214), .ZN(n1307) );
XNOR2_X1 U1012 ( .A(G131), .B(n1308), .ZN(n1295) );
XNOR2_X1 U1013 ( .A(KEYINPUT41), .B(n1225), .ZN(n1308) );
XNOR2_X1 U1014 ( .A(n1309), .B(G478), .ZN(n1251) );
NAND2_X1 U1015 ( .A1(n1135), .A2(n1183), .ZN(n1309) );
XNOR2_X1 U1016 ( .A(n1310), .B(n1311), .ZN(n1135) );
NOR2_X1 U1017 ( .A1(n1283), .A2(n1312), .ZN(n1311) );
INV_X1 U1018 ( .A(G217), .ZN(n1312) );
NAND2_X1 U1019 ( .A1(n1313), .A2(n1115), .ZN(n1283) );
XOR2_X1 U1020 ( .A(KEYINPUT5), .B(G234), .Z(n1313) );
NAND3_X1 U1021 ( .A1(n1314), .A2(n1315), .A3(KEYINPUT51), .ZN(n1310) );
NAND2_X1 U1022 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
NAND2_X1 U1023 ( .A1(KEYINPUT31), .A2(n1041), .ZN(n1317) );
XOR2_X1 U1024 ( .A(n1318), .B(n1319), .Z(n1316) );
AND2_X1 U1025 ( .A1(n1320), .A2(KEYINPUT32), .ZN(n1318) );
NAND3_X1 U1026 ( .A1(n1321), .A2(n1041), .A3(KEYINPUT31), .ZN(n1314) );
INV_X1 U1027 ( .A(G107), .ZN(n1041) );
XOR2_X1 U1028 ( .A(n1322), .B(n1319), .Z(n1321) );
XOR2_X1 U1029 ( .A(G134), .B(n1323), .Z(n1319) );
NOR2_X1 U1030 ( .A1(n1324), .A2(n1320), .ZN(n1322) );
INV_X1 U1031 ( .A(KEYINPUT32), .ZN(n1324) );
NAND2_X1 U1032 ( .A1(n1089), .A2(n1325), .ZN(n1253) );
NAND3_X1 U1033 ( .A1(n1125), .A2(n1243), .A3(G902), .ZN(n1325) );
NOR2_X1 U1034 ( .A1(n1115), .A2(G898), .ZN(n1125) );
NAND3_X1 U1035 ( .A1(n1243), .A2(n1115), .A3(G952), .ZN(n1089) );
NAND2_X1 U1036 ( .A1(G237), .A2(G234), .ZN(n1243) );
INV_X1 U1037 ( .A(n1224), .ZN(n1056) );
NAND2_X1 U1038 ( .A1(n1057), .A2(n1326), .ZN(n1224) );
NAND2_X1 U1039 ( .A1(n1231), .A2(n1102), .ZN(n1326) );
NAND3_X1 U1040 ( .A1(n1327), .A2(n1328), .A3(G210), .ZN(n1102) );
INV_X1 U1041 ( .A(n1059), .ZN(n1231) );
NOR2_X1 U1042 ( .A1(n1328), .A2(n1329), .ZN(n1059) );
AND2_X1 U1043 ( .A1(G237), .A2(G210), .ZN(n1329) );
NAND2_X1 U1044 ( .A1(n1330), .A2(n1183), .ZN(n1328) );
XOR2_X1 U1045 ( .A(n1331), .B(n1332), .Z(n1330) );
XNOR2_X1 U1046 ( .A(n1177), .B(n1333), .ZN(n1332) );
NOR2_X1 U1047 ( .A1(KEYINPUT21), .A2(n1181), .ZN(n1333) );
XNOR2_X1 U1048 ( .A(n1334), .B(n1335), .ZN(n1181) );
XOR2_X1 U1049 ( .A(n1336), .B(n1337), .Z(n1335) );
XNOR2_X1 U1050 ( .A(KEYINPUT59), .B(n1165), .ZN(n1337) );
NOR2_X1 U1051 ( .A1(G101), .A2(KEYINPUT44), .ZN(n1336) );
XNOR2_X1 U1052 ( .A(n1320), .B(n1338), .ZN(n1334) );
XOR2_X1 U1053 ( .A(n1339), .B(n1275), .Z(n1338) );
XOR2_X1 U1054 ( .A(G113), .B(G119), .Z(n1275) );
XNOR2_X1 U1055 ( .A(G116), .B(n1247), .ZN(n1320) );
INV_X1 U1056 ( .A(G122), .ZN(n1247) );
NAND2_X1 U1057 ( .A1(n1340), .A2(n1115), .ZN(n1177) );
XNOR2_X1 U1058 ( .A(G224), .B(KEYINPUT40), .ZN(n1340) );
XNOR2_X1 U1059 ( .A(G125), .B(n1179), .ZN(n1331) );
NAND2_X1 U1060 ( .A1(n1341), .A2(n1342), .ZN(n1179) );
NAND2_X1 U1061 ( .A1(n1343), .A2(n1222), .ZN(n1342) );
XNOR2_X1 U1062 ( .A(KEYINPUT60), .B(n1323), .ZN(n1343) );
XNOR2_X1 U1063 ( .A(n1233), .B(G143), .ZN(n1323) );
NAND2_X1 U1064 ( .A1(G214), .A2(n1327), .ZN(n1057) );
NAND2_X1 U1065 ( .A1(n1271), .A2(n1183), .ZN(n1327) );
INV_X1 U1066 ( .A(G237), .ZN(n1271) );
XNOR2_X1 U1067 ( .A(n1087), .B(KEYINPUT48), .ZN(n1266) );
NOR2_X1 U1068 ( .A1(n1085), .A2(n1084), .ZN(n1087) );
INV_X1 U1069 ( .A(n1264), .ZN(n1084) );
NAND2_X1 U1070 ( .A1(G221), .A2(n1278), .ZN(n1264) );
NAND2_X1 U1071 ( .A1(G234), .A2(n1183), .ZN(n1278) );
XOR2_X1 U1072 ( .A(n1344), .B(G469), .Z(n1085) );
NAND2_X1 U1073 ( .A1(n1345), .A2(n1183), .ZN(n1344) );
INV_X1 U1074 ( .A(G902), .ZN(n1183) );
XOR2_X1 U1075 ( .A(n1346), .B(n1347), .Z(n1345) );
XNOR2_X1 U1076 ( .A(n1166), .B(n1168), .ZN(n1347) );
XNOR2_X1 U1077 ( .A(n1348), .B(n1349), .ZN(n1168) );
XOR2_X1 U1078 ( .A(n1111), .B(n1350), .Z(n1349) );
NAND2_X1 U1079 ( .A1(KEYINPUT29), .A2(G101), .ZN(n1350) );
NAND2_X1 U1080 ( .A1(n1341), .A2(n1351), .ZN(n1111) );
NAND2_X1 U1081 ( .A1(n1352), .A2(n1222), .ZN(n1351) );
INV_X1 U1082 ( .A(G146), .ZN(n1222) );
XOR2_X1 U1083 ( .A(KEYINPUT3), .B(n1353), .Z(n1352) );
NAND2_X1 U1084 ( .A1(G146), .A2(n1353), .ZN(n1341) );
XNOR2_X1 U1085 ( .A(n1233), .B(n1354), .ZN(n1353) );
XNOR2_X1 U1086 ( .A(KEYINPUT60), .B(n1225), .ZN(n1354) );
INV_X1 U1087 ( .A(G143), .ZN(n1225) );
INV_X1 U1088 ( .A(G128), .ZN(n1233) );
XNOR2_X1 U1089 ( .A(n1114), .B(n1339), .ZN(n1348) );
XOR2_X1 U1090 ( .A(G104), .B(G107), .Z(n1339) );
XOR2_X1 U1091 ( .A(G131), .B(n1355), .Z(n1114) );
XOR2_X1 U1092 ( .A(G137), .B(G134), .Z(n1355) );
NAND2_X1 U1093 ( .A1(G227), .A2(n1115), .ZN(n1166) );
INV_X1 U1094 ( .A(G953), .ZN(n1115) );
XNOR2_X1 U1095 ( .A(G140), .B(n1165), .ZN(n1346) );
INV_X1 U1096 ( .A(G110), .ZN(n1165) );
endmodule


