//Key = 1000000110101001000100101111111101100100111011010111001010000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325;

XOR2_X1 U731 ( .A(n1004), .B(n1005), .Z(G9) );
XOR2_X1 U732 ( .A(KEYINPUT26), .B(G107), .Z(n1005) );
NOR2_X1 U733 ( .A1(n1006), .A2(n1007), .ZN(G75) );
NOR3_X1 U734 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1007) );
NAND3_X1 U735 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1008) );
NAND2_X1 U736 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND2_X1 U737 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NAND4_X1 U738 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
NAND2_X1 U739 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND3_X1 U740 ( .A1(n1024), .A2(n1025), .A3(KEYINPUT38), .ZN(n1023) );
NAND3_X1 U741 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1020) );
NAND2_X1 U742 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NAND2_X1 U743 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U744 ( .A1(n1024), .A2(n1033), .ZN(n1026) );
NAND2_X1 U745 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U746 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U747 ( .A1(n1024), .A2(n1038), .A3(n1029), .ZN(n1016) );
NAND3_X1 U748 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NAND2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U750 ( .A1(n1019), .A2(n1044), .ZN(n1039) );
NAND2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
OR3_X1 U752 ( .A1(n1047), .A2(KEYINPUT38), .A3(n1028), .ZN(n1046) );
NOR3_X1 U753 ( .A1(n1048), .A2(G953), .A3(G952), .ZN(n1006) );
INV_X1 U754 ( .A(n1011), .ZN(n1048) );
NAND4_X1 U755 ( .A1(n1049), .A2(n1024), .A3(n1050), .A4(n1051), .ZN(n1011) );
NOR4_X1 U756 ( .A1(n1036), .A2(n1022), .A3(n1052), .A4(n1053), .ZN(n1051) );
XOR2_X1 U757 ( .A(n1054), .B(n1055), .Z(n1052) );
NOR2_X1 U758 ( .A1(G475), .A2(KEYINPUT57), .ZN(n1055) );
NAND2_X1 U759 ( .A1(n1056), .A2(n1057), .ZN(G72) );
NAND2_X1 U760 ( .A1(n1058), .A2(n1012), .ZN(n1057) );
XOR2_X1 U761 ( .A(n1059), .B(n1060), .Z(n1058) );
NAND2_X1 U762 ( .A1(KEYINPUT37), .A2(n1010), .ZN(n1060) );
NAND2_X1 U763 ( .A1(n1061), .A2(G953), .ZN(n1056) );
XOR2_X1 U764 ( .A(n1059), .B(n1062), .Z(n1061) );
NOR2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1059) );
NAND2_X1 U767 ( .A1(G953), .A2(n1064), .ZN(n1066) );
XOR2_X1 U768 ( .A(n1067), .B(n1068), .Z(n1065) );
XOR2_X1 U769 ( .A(n1069), .B(n1070), .Z(n1068) );
XNOR2_X1 U770 ( .A(KEYINPUT25), .B(KEYINPUT11), .ZN(n1070) );
XOR2_X1 U771 ( .A(n1071), .B(n1072), .Z(n1067) );
XOR2_X1 U772 ( .A(n1073), .B(n1074), .Z(n1071) );
XOR2_X1 U773 ( .A(n1075), .B(n1076), .Z(G69) );
XOR2_X1 U774 ( .A(n1077), .B(n1078), .Z(n1076) );
AND2_X1 U775 ( .A1(n1009), .A2(n1012), .ZN(n1078) );
NOR2_X1 U776 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
XOR2_X1 U777 ( .A(KEYINPUT24), .B(G953), .Z(n1080) );
AND2_X1 U778 ( .A1(G224), .A2(G898), .ZN(n1079) );
NOR2_X1 U779 ( .A1(n1081), .A2(n1082), .ZN(n1075) );
NOR2_X1 U780 ( .A1(n1083), .A2(n1084), .ZN(G66) );
XOR2_X1 U781 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U782 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U783 ( .A1(KEYINPUT30), .A2(n1089), .ZN(n1085) );
NOR2_X1 U784 ( .A1(n1083), .A2(n1090), .ZN(G63) );
XOR2_X1 U785 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U786 ( .A1(n1093), .A2(G478), .ZN(n1091) );
NOR2_X1 U787 ( .A1(n1083), .A2(n1094), .ZN(G60) );
XOR2_X1 U788 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND2_X1 U789 ( .A1(n1093), .A2(G475), .ZN(n1095) );
XOR2_X1 U790 ( .A(n1097), .B(n1098), .Z(G6) );
NOR2_X1 U791 ( .A1(KEYINPUT62), .A2(n1099), .ZN(n1098) );
NOR2_X1 U792 ( .A1(n1083), .A2(n1100), .ZN(G57) );
XOR2_X1 U793 ( .A(n1101), .B(n1102), .Z(n1100) );
XOR2_X1 U794 ( .A(n1103), .B(n1104), .Z(n1102) );
XOR2_X1 U795 ( .A(n1105), .B(n1106), .Z(n1103) );
NOR2_X1 U796 ( .A1(G101), .A2(KEYINPUT48), .ZN(n1106) );
NAND2_X1 U797 ( .A1(n1093), .A2(G472), .ZN(n1105) );
XOR2_X1 U798 ( .A(n1107), .B(n1108), .Z(n1101) );
NOR2_X1 U799 ( .A1(KEYINPUT18), .A2(n1109), .ZN(n1108) );
XOR2_X1 U800 ( .A(n1110), .B(KEYINPUT1), .Z(n1107) );
NOR2_X1 U801 ( .A1(n1083), .A2(n1111), .ZN(G54) );
XOR2_X1 U802 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U803 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U804 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U805 ( .A(n1118), .B(n1119), .Z(n1117) );
INV_X1 U806 ( .A(KEYINPUT36), .ZN(n1116) );
NOR2_X1 U807 ( .A1(KEYINPUT36), .A2(n1120), .ZN(n1114) );
XOR2_X1 U808 ( .A(n1118), .B(n1121), .Z(n1120) );
XNOR2_X1 U809 ( .A(n1122), .B(n1123), .ZN(n1118) );
NAND2_X1 U810 ( .A1(KEYINPUT56), .A2(n1124), .ZN(n1123) );
INV_X1 U811 ( .A(G140), .ZN(n1124) );
NAND2_X1 U812 ( .A1(KEYINPUT40), .A2(n1125), .ZN(n1122) );
XOR2_X1 U813 ( .A(n1126), .B(n1127), .Z(n1112) );
NAND2_X1 U814 ( .A1(n1128), .A2(n1093), .ZN(n1126) );
XNOR2_X1 U815 ( .A(G469), .B(KEYINPUT19), .ZN(n1128) );
NOR2_X1 U816 ( .A1(n1083), .A2(n1129), .ZN(G51) );
XOR2_X1 U817 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U818 ( .A(n1132), .B(n1082), .Z(n1131) );
XOR2_X1 U819 ( .A(n1133), .B(n1134), .Z(n1130) );
NOR3_X1 U820 ( .A1(n1135), .A2(G953), .A3(n1136), .ZN(n1134) );
INV_X1 U821 ( .A(G224), .ZN(n1136) );
XOR2_X1 U822 ( .A(KEYINPUT5), .B(KEYINPUT17), .Z(n1135) );
NAND2_X1 U823 ( .A1(n1093), .A2(n1137), .ZN(n1133) );
INV_X1 U824 ( .A(n1088), .ZN(n1093) );
NAND2_X1 U825 ( .A1(G902), .A2(n1138), .ZN(n1088) );
OR2_X1 U826 ( .A1(n1010), .A2(n1009), .ZN(n1138) );
NAND4_X1 U827 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1009) );
NOR4_X1 U828 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1097), .ZN(n1142) );
AND3_X1 U829 ( .A1(n1024), .A2(n1146), .A3(n1147), .ZN(n1097) );
OR2_X1 U830 ( .A1(n1004), .A2(KEYINPUT52), .ZN(n1141) );
NAND3_X1 U831 ( .A1(n1024), .A2(n1146), .A3(n1043), .ZN(n1004) );
NAND2_X1 U832 ( .A1(n1148), .A2(n1149), .ZN(n1140) );
NAND2_X1 U833 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
NAND4_X1 U834 ( .A1(KEYINPUT52), .A2(n1043), .A3(n1152), .A4(n1024), .ZN(n1151) );
NOR2_X1 U835 ( .A1(n1153), .A2(n1045), .ZN(n1152) );
NAND3_X1 U836 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1150) );
XOR2_X1 U837 ( .A(KEYINPUT35), .B(n1153), .Z(n1155) );
NAND2_X1 U838 ( .A1(n1019), .A2(n1157), .ZN(n1139) );
NAND2_X1 U839 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U840 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U841 ( .A1(n1162), .A2(n1146), .ZN(n1158) );
NAND4_X1 U842 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1010) );
AND3_X1 U843 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1166) );
NAND2_X1 U844 ( .A1(n1153), .A2(n1170), .ZN(n1165) );
NAND2_X1 U845 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XOR2_X1 U846 ( .A(KEYINPUT45), .B(n1173), .Z(n1171) );
NAND3_X1 U847 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1163) );
NAND2_X1 U848 ( .A1(n1177), .A2(n1031), .ZN(n1175) );
XOR2_X1 U849 ( .A(KEYINPUT44), .B(n1154), .Z(n1177) );
NOR2_X1 U850 ( .A1(n1012), .A2(G952), .ZN(n1083) );
XNOR2_X1 U851 ( .A(G146), .B(n1164), .ZN(G48) );
NAND3_X1 U852 ( .A1(n1178), .A2(n1153), .A3(n1147), .ZN(n1164) );
XNOR2_X1 U853 ( .A(G143), .B(n1167), .ZN(G45) );
NAND4_X1 U854 ( .A1(n1153), .A2(n1174), .A3(n1154), .A4(n1179), .ZN(n1167) );
NOR3_X1 U855 ( .A1(n1050), .A2(n1180), .A3(n1181), .ZN(n1179) );
XOR2_X1 U856 ( .A(G140), .B(n1182), .Z(G42) );
NOR3_X1 U857 ( .A1(n1031), .A2(n1183), .A3(n1184), .ZN(n1182) );
XOR2_X1 U858 ( .A(n1045), .B(KEYINPUT4), .Z(n1183) );
INV_X1 U859 ( .A(n1162), .ZN(n1031) );
NAND2_X1 U860 ( .A1(n1185), .A2(n1186), .ZN(G39) );
NAND2_X1 U861 ( .A1(G137), .A2(n1169), .ZN(n1186) );
XOR2_X1 U862 ( .A(KEYINPUT7), .B(n1187), .Z(n1185) );
NOR2_X1 U863 ( .A1(G137), .A2(n1169), .ZN(n1187) );
NAND3_X1 U864 ( .A1(n1178), .A2(n1029), .A3(n1019), .ZN(n1169) );
XOR2_X1 U865 ( .A(n1188), .B(n1168), .Z(G36) );
NAND4_X1 U866 ( .A1(n1154), .A2(n1029), .A3(n1189), .A4(n1043), .ZN(n1168) );
NOR2_X1 U867 ( .A1(n1180), .A2(n1045), .ZN(n1189) );
INV_X1 U868 ( .A(n1190), .ZN(n1180) );
XOR2_X1 U869 ( .A(n1069), .B(n1191), .Z(G33) );
NAND3_X1 U870 ( .A1(n1154), .A2(n1174), .A3(n1176), .ZN(n1191) );
INV_X1 U871 ( .A(n1184), .ZN(n1176) );
NAND3_X1 U872 ( .A1(n1029), .A2(n1190), .A3(n1147), .ZN(n1184) );
INV_X1 U873 ( .A(n1025), .ZN(n1029) );
NAND2_X1 U874 ( .A1(n1037), .A2(n1192), .ZN(n1025) );
XOR2_X1 U875 ( .A(n1193), .B(n1194), .Z(G30) );
NAND2_X1 U876 ( .A1(n1173), .A2(n1153), .ZN(n1194) );
AND2_X1 U877 ( .A1(n1178), .A2(n1043), .ZN(n1173) );
AND3_X1 U878 ( .A1(n1174), .A2(n1190), .A3(n1161), .ZN(n1178) );
INV_X1 U879 ( .A(n1045), .ZN(n1174) );
XOR2_X1 U880 ( .A(G101), .B(n1145), .Z(G3) );
AND3_X1 U881 ( .A1(n1154), .A2(n1146), .A3(n1019), .ZN(n1145) );
NOR3_X1 U882 ( .A1(n1045), .A2(n1195), .A3(n1034), .ZN(n1146) );
XOR2_X1 U883 ( .A(n1196), .B(n1197), .Z(G27) );
XOR2_X1 U884 ( .A(KEYINPUT43), .B(G125), .Z(n1197) );
NOR2_X1 U885 ( .A1(n1198), .A2(n1034), .ZN(n1196) );
XOR2_X1 U886 ( .A(n1172), .B(KEYINPUT39), .Z(n1198) );
NAND3_X1 U887 ( .A1(n1156), .A2(n1190), .A3(n1162), .ZN(n1172) );
NAND2_X1 U888 ( .A1(n1199), .A2(n1200), .ZN(n1190) );
NAND4_X1 U889 ( .A1(n1201), .A2(G953), .A3(G902), .A4(n1015), .ZN(n1200) );
XOR2_X1 U890 ( .A(n1064), .B(KEYINPUT14), .Z(n1201) );
INV_X1 U891 ( .A(G900), .ZN(n1064) );
XOR2_X1 U892 ( .A(G122), .B(n1144), .Z(G24) );
AND4_X1 U893 ( .A1(n1160), .A2(n1024), .A3(n1202), .A4(n1203), .ZN(n1144) );
NOR2_X1 U894 ( .A1(n1204), .A2(n1205), .ZN(n1024) );
XNOR2_X1 U895 ( .A(G119), .B(n1206), .ZN(G21) );
NAND3_X1 U896 ( .A1(n1019), .A2(n1207), .A3(n1160), .ZN(n1206) );
XOR2_X1 U897 ( .A(KEYINPUT21), .B(n1161), .Z(n1207) );
AND2_X1 U898 ( .A1(n1205), .A2(n1204), .ZN(n1161) );
XOR2_X1 U899 ( .A(n1143), .B(n1208), .Z(G18) );
NOR2_X1 U900 ( .A1(KEYINPUT23), .A2(n1209), .ZN(n1208) );
AND3_X1 U901 ( .A1(n1154), .A2(n1043), .A3(n1160), .ZN(n1143) );
AND3_X1 U902 ( .A1(n1153), .A2(n1149), .A3(n1042), .ZN(n1160) );
NOR2_X1 U903 ( .A1(n1203), .A2(n1050), .ZN(n1043) );
XOR2_X1 U904 ( .A(n1210), .B(n1211), .Z(G15) );
NAND4_X1 U905 ( .A1(n1212), .A2(n1156), .A3(n1154), .A4(n1153), .ZN(n1211) );
INV_X1 U906 ( .A(n1032), .ZN(n1154) );
NAND2_X1 U907 ( .A1(n1213), .A2(n1204), .ZN(n1032) );
XOR2_X1 U908 ( .A(KEYINPUT31), .B(n1205), .Z(n1213) );
INV_X1 U909 ( .A(n1214), .ZN(n1205) );
INV_X1 U910 ( .A(n1040), .ZN(n1156) );
NAND2_X1 U911 ( .A1(n1042), .A2(n1147), .ZN(n1040) );
NOR2_X1 U912 ( .A1(n1202), .A2(n1181), .ZN(n1147) );
NOR2_X1 U913 ( .A1(n1047), .A2(n1022), .ZN(n1042) );
INV_X1 U914 ( .A(n1028), .ZN(n1022) );
XOR2_X1 U915 ( .A(n1149), .B(KEYINPUT6), .Z(n1212) );
XNOR2_X1 U916 ( .A(G110), .B(n1215), .ZN(G12) );
NAND3_X1 U917 ( .A1(n1162), .A2(n1019), .A3(n1216), .ZN(n1215) );
NOR3_X1 U918 ( .A1(n1045), .A2(n1195), .A3(n1217), .ZN(n1216) );
XOR2_X1 U919 ( .A(n1034), .B(KEYINPUT13), .Z(n1217) );
INV_X1 U920 ( .A(n1153), .ZN(n1034) );
NOR2_X1 U921 ( .A1(n1037), .A2(n1036), .ZN(n1153) );
INV_X1 U922 ( .A(n1192), .ZN(n1036) );
NAND2_X1 U923 ( .A1(G214), .A2(n1218), .ZN(n1192) );
XOR2_X1 U924 ( .A(n1053), .B(KEYINPUT27), .Z(n1037) );
XNOR2_X1 U925 ( .A(n1219), .B(n1137), .ZN(n1053) );
AND2_X1 U926 ( .A1(G210), .A2(n1218), .ZN(n1137) );
NAND2_X1 U927 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
XOR2_X1 U928 ( .A(KEYINPUT15), .B(G237), .Z(n1220) );
NAND2_X1 U929 ( .A1(n1222), .A2(n1223), .ZN(n1219) );
XNOR2_X1 U930 ( .A(n1224), .B(n1082), .ZN(n1222) );
XNOR2_X1 U931 ( .A(n1225), .B(n1226), .ZN(n1082) );
XOR2_X1 U932 ( .A(n1227), .B(n1228), .Z(n1226) );
NAND2_X1 U933 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
OR2_X1 U934 ( .A1(n1231), .A2(KEYINPUT58), .ZN(n1230) );
NAND3_X1 U935 ( .A1(G104), .A2(n1232), .A3(KEYINPUT58), .ZN(n1229) );
NAND3_X1 U936 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(n1227) );
OR2_X1 U937 ( .A1(n1210), .A2(n1236), .ZN(n1235) );
NAND2_X1 U938 ( .A1(n1237), .A2(n1238), .ZN(n1234) );
INV_X1 U939 ( .A(KEYINPUT29), .ZN(n1238) );
NAND2_X1 U940 ( .A1(n1236), .A2(n1239), .ZN(n1237) );
XOR2_X1 U941 ( .A(KEYINPUT33), .B(G113), .Z(n1239) );
NAND2_X1 U942 ( .A1(KEYINPUT29), .A2(n1240), .ZN(n1233) );
NAND2_X1 U943 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
OR2_X1 U944 ( .A1(n1210), .A2(KEYINPUT33), .ZN(n1242) );
NAND3_X1 U945 ( .A1(n1236), .A2(n1210), .A3(KEYINPUT33), .ZN(n1241) );
INV_X1 U946 ( .A(G113), .ZN(n1210) );
XNOR2_X1 U947 ( .A(G101), .B(n1243), .ZN(n1225) );
XOR2_X1 U948 ( .A(G122), .B(G110), .Z(n1243) );
NAND3_X1 U949 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1224) );
NAND2_X1 U950 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
OR3_X1 U951 ( .A1(n1248), .A2(n1247), .A3(KEYINPUT32), .ZN(n1245) );
XNOR2_X1 U952 ( .A(n1132), .B(KEYINPUT47), .ZN(n1247) );
XOR2_X1 U953 ( .A(G125), .B(n1109), .Z(n1132) );
NAND2_X1 U954 ( .A1(KEYINPUT41), .A2(n1249), .ZN(n1248) );
NAND2_X1 U955 ( .A1(G224), .A2(n1012), .ZN(n1249) );
NAND3_X1 U956 ( .A1(G224), .A2(n1012), .A3(KEYINPUT32), .ZN(n1244) );
INV_X1 U957 ( .A(n1149), .ZN(n1195) );
NAND2_X1 U958 ( .A1(n1199), .A2(n1250), .ZN(n1149) );
NAND3_X1 U959 ( .A1(G902), .A2(n1015), .A3(n1081), .ZN(n1250) );
NOR2_X1 U960 ( .A1(n1012), .A2(G898), .ZN(n1081) );
NAND3_X1 U961 ( .A1(n1015), .A2(n1012), .A3(G952), .ZN(n1199) );
NAND2_X1 U962 ( .A1(G237), .A2(n1251), .ZN(n1015) );
NAND2_X1 U963 ( .A1(n1047), .A2(n1028), .ZN(n1045) );
NAND2_X1 U964 ( .A1(G221), .A2(n1252), .ZN(n1028) );
INV_X1 U965 ( .A(n1018), .ZN(n1047) );
XOR2_X1 U966 ( .A(n1049), .B(KEYINPUT20), .Z(n1018) );
XOR2_X1 U967 ( .A(n1253), .B(n1254), .Z(n1049) );
XOR2_X1 U968 ( .A(KEYINPUT63), .B(G469), .Z(n1254) );
NAND2_X1 U969 ( .A1(n1255), .A2(n1223), .ZN(n1253) );
XOR2_X1 U970 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U971 ( .A(G140), .B(n1127), .Z(n1257) );
XOR2_X1 U972 ( .A(G110), .B(n1258), .Z(n1127) );
NOR2_X1 U973 ( .A1(G953), .A2(n1063), .ZN(n1258) );
INV_X1 U974 ( .A(G227), .ZN(n1063) );
NOR2_X1 U975 ( .A1(n1259), .A2(n1260), .ZN(n1256) );
NOR2_X1 U976 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
INV_X1 U977 ( .A(n1121), .ZN(n1261) );
NOR2_X1 U978 ( .A1(n1121), .A2(n1263), .ZN(n1259) );
XOR2_X1 U979 ( .A(n1262), .B(KEYINPUT8), .Z(n1263) );
XOR2_X1 U980 ( .A(n1125), .B(KEYINPUT0), .Z(n1262) );
NOR2_X1 U981 ( .A1(n1119), .A2(n1264), .ZN(n1121) );
AND2_X1 U982 ( .A1(n1265), .A2(n1074), .ZN(n1264) );
NOR2_X1 U983 ( .A1(n1074), .A2(n1265), .ZN(n1119) );
XNOR2_X1 U984 ( .A(G101), .B(n1231), .ZN(n1265) );
XNOR2_X1 U985 ( .A(n1099), .B(G107), .ZN(n1231) );
INV_X1 U986 ( .A(G104), .ZN(n1099) );
XNOR2_X1 U987 ( .A(n1266), .B(n1267), .ZN(n1074) );
NAND2_X1 U988 ( .A1(KEYINPUT50), .A2(n1268), .ZN(n1266) );
XOR2_X1 U989 ( .A(KEYINPUT3), .B(n1269), .Z(n1268) );
NOR2_X1 U990 ( .A1(n1202), .A2(n1203), .ZN(n1019) );
INV_X1 U991 ( .A(n1181), .ZN(n1203) );
XOR2_X1 U992 ( .A(n1054), .B(G475), .Z(n1181) );
NAND2_X1 U993 ( .A1(n1096), .A2(n1223), .ZN(n1054) );
XNOR2_X1 U994 ( .A(n1270), .B(n1271), .ZN(n1096) );
XOR2_X1 U995 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U996 ( .A(G113), .B(G104), .Z(n1273) );
XOR2_X1 U997 ( .A(G131), .B(G122), .Z(n1272) );
XOR2_X1 U998 ( .A(n1274), .B(n1275), .Z(n1270) );
XOR2_X1 U999 ( .A(n1276), .B(n1269), .Z(n1274) );
NAND2_X1 U1000 ( .A1(G214), .A2(n1277), .ZN(n1276) );
INV_X1 U1001 ( .A(n1050), .ZN(n1202) );
XOR2_X1 U1002 ( .A(n1278), .B(G478), .Z(n1050) );
NAND2_X1 U1003 ( .A1(n1092), .A2(n1223), .ZN(n1278) );
NAND2_X1 U1004 ( .A1(n1279), .A2(n1280), .ZN(n1092) );
NAND2_X1 U1005 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XOR2_X1 U1006 ( .A(n1283), .B(KEYINPUT46), .Z(n1281) );
NAND2_X1 U1007 ( .A1(n1284), .A2(n1285), .ZN(n1279) );
INV_X1 U1008 ( .A(n1282), .ZN(n1285) );
XOR2_X1 U1009 ( .A(n1232), .B(n1286), .Z(n1282) );
XOR2_X1 U1010 ( .A(G122), .B(G116), .Z(n1286) );
INV_X1 U1011 ( .A(G107), .ZN(n1232) );
XOR2_X1 U1012 ( .A(KEYINPUT55), .B(n1287), .Z(n1284) );
INV_X1 U1013 ( .A(n1283), .ZN(n1287) );
XOR2_X1 U1014 ( .A(n1288), .B(n1289), .Z(n1283) );
XOR2_X1 U1015 ( .A(n1290), .B(n1291), .Z(n1289) );
NAND2_X1 U1016 ( .A1(G217), .A2(n1292), .ZN(n1291) );
NAND2_X1 U1017 ( .A1(KEYINPUT12), .A2(n1193), .ZN(n1290) );
INV_X1 U1018 ( .A(G128), .ZN(n1193) );
XOR2_X1 U1019 ( .A(G143), .B(n1188), .Z(n1288) );
NOR2_X1 U1020 ( .A1(n1204), .A2(n1214), .ZN(n1162) );
XNOR2_X1 U1021 ( .A(n1293), .B(n1087), .ZN(n1214) );
NAND2_X1 U1022 ( .A1(G217), .A2(n1252), .ZN(n1087) );
NAND2_X1 U1023 ( .A1(n1294), .A2(n1251), .ZN(n1252) );
XOR2_X1 U1024 ( .A(G234), .B(KEYINPUT2), .Z(n1251) );
XOR2_X1 U1025 ( .A(n1221), .B(KEYINPUT53), .Z(n1294) );
INV_X1 U1026 ( .A(G902), .ZN(n1221) );
NAND2_X1 U1027 ( .A1(n1089), .A2(n1223), .ZN(n1293) );
XNOR2_X1 U1028 ( .A(n1295), .B(n1296), .ZN(n1089) );
XOR2_X1 U1029 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U1030 ( .A(G137), .B(G128), .Z(n1298) );
XOR2_X1 U1031 ( .A(KEYINPUT9), .B(G146), .Z(n1297) );
XOR2_X1 U1032 ( .A(n1299), .B(n1300), .Z(n1295) );
XOR2_X1 U1033 ( .A(G119), .B(G110), .Z(n1300) );
XOR2_X1 U1034 ( .A(n1301), .B(n1275), .Z(n1299) );
XOR2_X1 U1035 ( .A(n1072), .B(KEYINPUT16), .Z(n1275) );
XOR2_X1 U1036 ( .A(G125), .B(G140), .Z(n1072) );
NAND2_X1 U1037 ( .A1(G221), .A2(n1292), .ZN(n1301) );
AND2_X1 U1038 ( .A1(G234), .A2(n1012), .ZN(n1292) );
INV_X1 U1039 ( .A(G953), .ZN(n1012) );
XNOR2_X1 U1040 ( .A(n1302), .B(G472), .ZN(n1204) );
NAND2_X1 U1041 ( .A1(n1303), .A2(n1223), .ZN(n1302) );
XOR2_X1 U1042 ( .A(G902), .B(KEYINPUT22), .Z(n1223) );
XNOR2_X1 U1043 ( .A(n1110), .B(n1304), .ZN(n1303) );
XNOR2_X1 U1044 ( .A(G101), .B(n1305), .ZN(n1304) );
NAND2_X1 U1045 ( .A1(KEYINPUT54), .A2(n1306), .ZN(n1305) );
XOR2_X1 U1046 ( .A(n1307), .B(n1104), .Z(n1306) );
XNOR2_X1 U1047 ( .A(n1308), .B(n1309), .ZN(n1104) );
NOR2_X1 U1048 ( .A1(KEYINPUT61), .A2(n1236), .ZN(n1309) );
XOR2_X1 U1049 ( .A(n1209), .B(G119), .Z(n1236) );
INV_X1 U1050 ( .A(G116), .ZN(n1209) );
XOR2_X1 U1051 ( .A(n1125), .B(G113), .Z(n1308) );
NAND3_X1 U1052 ( .A1(n1310), .A2(n1311), .A3(n1312), .ZN(n1125) );
NAND2_X1 U1053 ( .A1(G131), .A2(n1313), .ZN(n1312) );
NAND2_X1 U1054 ( .A1(KEYINPUT42), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1055 ( .A(n1315), .B(n1316), .Z(n1314) );
NAND3_X1 U1056 ( .A1(KEYINPUT51), .A2(n1317), .A3(n1316), .ZN(n1311) );
INV_X1 U1057 ( .A(n1318), .ZN(n1316) );
NAND2_X1 U1058 ( .A1(KEYINPUT34), .A2(n1319), .ZN(n1317) );
NAND3_X1 U1059 ( .A1(n1320), .A2(n1321), .A3(n1318), .ZN(n1310) );
NAND2_X1 U1060 ( .A1(n1322), .A2(n1323), .ZN(n1318) );
NAND2_X1 U1061 ( .A1(KEYINPUT10), .A2(n1073), .ZN(n1323) );
XOR2_X1 U1062 ( .A(n1188), .B(G137), .Z(n1073) );
OR3_X1 U1063 ( .A1(n1188), .A2(G137), .A3(KEYINPUT10), .ZN(n1322) );
INV_X1 U1064 ( .A(G134), .ZN(n1188) );
INV_X1 U1065 ( .A(KEYINPUT51), .ZN(n1321) );
NAND2_X1 U1066 ( .A1(n1315), .A2(n1319), .ZN(n1320) );
NAND2_X1 U1067 ( .A1(KEYINPUT42), .A2(n1069), .ZN(n1319) );
INV_X1 U1068 ( .A(G131), .ZN(n1069) );
INV_X1 U1069 ( .A(KEYINPUT34), .ZN(n1315) );
NOR2_X1 U1070 ( .A1(KEYINPUT59), .A2(n1324), .ZN(n1307) );
XOR2_X1 U1071 ( .A(n1109), .B(KEYINPUT60), .Z(n1324) );
XOR2_X1 U1072 ( .A(n1325), .B(n1267), .Z(n1109) );
XOR2_X1 U1073 ( .A(G128), .B(KEYINPUT49), .Z(n1267) );
NAND2_X1 U1074 ( .A1(KEYINPUT28), .A2(n1269), .ZN(n1325) );
XOR2_X1 U1075 ( .A(G143), .B(G146), .Z(n1269) );
NAND2_X1 U1076 ( .A1(G210), .A2(n1277), .ZN(n1110) );
NOR2_X1 U1077 ( .A1(G953), .A2(G237), .ZN(n1277) );
endmodule


