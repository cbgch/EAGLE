//Key = 1000000111100011000000001111101100000100010011100110010101100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383;

XOR2_X1 U761 ( .A(n1054), .B(n1055), .Z(G9) );
NOR2_X1 U762 ( .A1(KEYINPUT34), .A2(G107), .ZN(n1055) );
NAND4_X1 U763 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1054) );
NOR2_X1 U764 ( .A1(n1060), .A2(n1061), .ZN(G75) );
NOR4_X1 U765 ( .A1(G953), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1061) );
NOR2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NOR2_X1 U767 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR3_X1 U768 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1068) );
NOR2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U772 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U773 ( .A1(n1080), .A2(n1056), .ZN(n1078) );
NOR2_X1 U774 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR3_X1 U775 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1076) );
INV_X1 U776 ( .A(n1086), .ZN(n1084) );
XNOR2_X1 U777 ( .A(KEYINPUT62), .B(n1087), .ZN(n1083) );
NOR2_X1 U778 ( .A1(n1088), .A2(n1087), .ZN(n1072) );
NOR2_X1 U779 ( .A1(n1089), .A2(n1058), .ZN(n1088) );
NOR2_X1 U780 ( .A1(n1090), .A2(n1079), .ZN(n1089) );
NOR2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR4_X1 U782 ( .A1(n1093), .A2(n1075), .A3(n1087), .A4(n1079), .ZN(n1067) );
NOR3_X1 U783 ( .A1(n1062), .A2(G953), .A3(G952), .ZN(n1060) );
AND4_X1 U784 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1062) );
NOR4_X1 U785 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
XOR2_X1 U786 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U787 ( .A(n1104), .B(n1105), .Z(n1100) );
XOR2_X1 U788 ( .A(KEYINPUT56), .B(n1106), .Z(n1099) );
NOR3_X1 U789 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1096) );
INV_X1 U790 ( .A(n1082), .ZN(n1109) );
NAND2_X1 U791 ( .A1(G469), .A2(n1110), .ZN(n1095) );
XOR2_X1 U792 ( .A(n1111), .B(n1112), .Z(n1094) );
XOR2_X1 U793 ( .A(KEYINPUT30), .B(G478), .Z(n1112) );
NOR2_X1 U794 ( .A1(KEYINPUT16), .A2(n1113), .ZN(n1111) );
XOR2_X1 U795 ( .A(n1114), .B(n1115), .Z(G72) );
NOR2_X1 U796 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
AND2_X1 U797 ( .A1(G227), .A2(G900), .ZN(n1116) );
NAND2_X1 U798 ( .A1(n1118), .A2(n1119), .ZN(n1114) );
NAND2_X1 U799 ( .A1(n1120), .A2(n1117), .ZN(n1119) );
XOR2_X1 U800 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U801 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
OR3_X1 U802 ( .A1(n1125), .A2(n1122), .A3(n1117), .ZN(n1118) );
XNOR2_X1 U803 ( .A(n1126), .B(n1127), .ZN(n1122) );
XOR2_X1 U804 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U805 ( .A(n1130), .B(n1131), .Z(n1126) );
NOR2_X1 U806 ( .A1(G131), .A2(KEYINPUT12), .ZN(n1131) );
XOR2_X1 U807 ( .A(n1132), .B(KEYINPUT37), .Z(n1130) );
NAND2_X1 U808 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U809 ( .A1(G125), .A2(n1135), .ZN(n1134) );
XOR2_X1 U810 ( .A(n1136), .B(KEYINPUT13), .Z(n1133) );
NAND2_X1 U811 ( .A1(G140), .A2(n1137), .ZN(n1136) );
NAND3_X1 U812 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(G69) );
XOR2_X1 U813 ( .A(n1141), .B(KEYINPUT1), .Z(n1140) );
NAND3_X1 U814 ( .A1(n1142), .A2(n1143), .A3(G953), .ZN(n1141) );
NAND2_X1 U815 ( .A1(G898), .A2(G224), .ZN(n1142) );
NAND2_X1 U816 ( .A1(n1144), .A2(n1117), .ZN(n1139) );
XOR2_X1 U817 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND3_X1 U818 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1145) );
XOR2_X1 U819 ( .A(KEYINPUT63), .B(n1150), .Z(n1147) );
NAND3_X1 U820 ( .A1(n1146), .A2(G224), .A3(G953), .ZN(n1138) );
INV_X1 U821 ( .A(n1143), .ZN(n1146) );
NAND2_X1 U822 ( .A1(n1151), .A2(n1152), .ZN(n1143) );
NAND2_X1 U823 ( .A1(G953), .A2(n1153), .ZN(n1152) );
XOR2_X1 U824 ( .A(n1154), .B(n1155), .Z(n1151) );
NOR2_X1 U825 ( .A1(KEYINPUT43), .A2(n1156), .ZN(n1155) );
XNOR2_X1 U826 ( .A(n1157), .B(n1158), .ZN(n1156) );
NOR3_X1 U827 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(G66) );
AND3_X1 U828 ( .A1(KEYINPUT23), .A2(G953), .A3(G952), .ZN(n1161) );
NOR2_X1 U829 ( .A1(KEYINPUT23), .A2(n1162), .ZN(n1160) );
INV_X1 U830 ( .A(n1163), .ZN(n1162) );
XOR2_X1 U831 ( .A(n1164), .B(n1165), .Z(n1159) );
NOR2_X1 U832 ( .A1(KEYINPUT47), .A2(n1166), .ZN(n1165) );
NAND2_X1 U833 ( .A1(n1167), .A2(n1168), .ZN(n1164) );
NOR2_X1 U834 ( .A1(n1163), .A2(n1169), .ZN(G63) );
XOR2_X1 U835 ( .A(n1170), .B(n1171), .Z(n1169) );
AND2_X1 U836 ( .A1(G478), .A2(n1167), .ZN(n1170) );
NOR2_X1 U837 ( .A1(n1163), .A2(n1172), .ZN(G60) );
XOR2_X1 U838 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U839 ( .A1(KEYINPUT17), .A2(n1175), .ZN(n1174) );
NOR2_X1 U840 ( .A1(n1104), .A2(n1176), .ZN(n1173) );
XNOR2_X1 U841 ( .A(G104), .B(n1177), .ZN(G6) );
NAND4_X1 U842 ( .A1(n1178), .A2(n1179), .A3(n1056), .A4(n1058), .ZN(n1177) );
XOR2_X1 U843 ( .A(n1059), .B(KEYINPUT3), .Z(n1178) );
NOR2_X1 U844 ( .A1(n1163), .A2(n1180), .ZN(G57) );
XOR2_X1 U845 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U846 ( .A(n1183), .B(n1184), .Z(n1182) );
XNOR2_X1 U847 ( .A(n1185), .B(n1186), .ZN(n1184) );
NOR3_X1 U848 ( .A1(n1176), .A2(KEYINPUT35), .A3(n1187), .ZN(n1186) );
INV_X1 U849 ( .A(G472), .ZN(n1187) );
XOR2_X1 U850 ( .A(n1188), .B(n1189), .Z(n1181) );
NOR2_X1 U851 ( .A1(n1163), .A2(n1190), .ZN(G54) );
NOR2_X1 U852 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U853 ( .A(KEYINPUT36), .B(n1193), .Z(n1192) );
NOR2_X1 U854 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
XNOR2_X1 U855 ( .A(n1196), .B(KEYINPUT39), .ZN(n1195) );
INV_X1 U856 ( .A(n1197), .ZN(n1194) );
NOR2_X1 U857 ( .A1(n1196), .A2(n1197), .ZN(n1191) );
NAND2_X1 U858 ( .A1(n1167), .A2(G469), .ZN(n1197) );
INV_X1 U859 ( .A(n1176), .ZN(n1167) );
XNOR2_X1 U860 ( .A(n1198), .B(n1199), .ZN(n1196) );
XNOR2_X1 U861 ( .A(n1185), .B(n1200), .ZN(n1199) );
XOR2_X1 U862 ( .A(n1201), .B(n1202), .Z(n1198) );
NOR2_X1 U863 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NOR2_X1 U864 ( .A1(G110), .A2(n1135), .ZN(n1203) );
INV_X1 U865 ( .A(G140), .ZN(n1135) );
NAND2_X1 U866 ( .A1(KEYINPUT27), .A2(n1205), .ZN(n1201) );
NOR2_X1 U867 ( .A1(n1163), .A2(n1206), .ZN(G51) );
XNOR2_X1 U868 ( .A(n1207), .B(n1208), .ZN(n1206) );
XOR2_X1 U869 ( .A(n1209), .B(n1210), .Z(n1208) );
NOR2_X1 U870 ( .A1(n1103), .A2(n1176), .ZN(n1210) );
NAND2_X1 U871 ( .A1(G902), .A2(n1064), .ZN(n1176) );
NAND4_X1 U872 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1149), .ZN(n1064) );
AND4_X1 U873 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1149) );
NOR2_X1 U874 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NOR3_X1 U875 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1219) );
NOR3_X1 U876 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1222) );
AND2_X1 U877 ( .A1(n1058), .A2(n1179), .ZN(n1225) );
NOR3_X1 U878 ( .A1(n1226), .A2(KEYINPUT15), .A3(n1227), .ZN(n1224) );
NOR2_X1 U879 ( .A1(n1228), .A2(n1059), .ZN(n1221) );
NOR3_X1 U880 ( .A1(n1079), .A2(KEYINPUT61), .A3(n1229), .ZN(n1228) );
NOR2_X1 U881 ( .A1(n1230), .A2(n1231), .ZN(n1218) );
NOR2_X1 U882 ( .A1(n1232), .A2(n1233), .ZN(n1230) );
NOR2_X1 U883 ( .A1(n1229), .A2(n1234), .ZN(n1233) );
INV_X1 U884 ( .A(KEYINPUT61), .ZN(n1234) );
AND2_X1 U885 ( .A1(n1235), .A2(KEYINPUT15), .ZN(n1232) );
NOR2_X1 U886 ( .A1(n1150), .A2(n1236), .ZN(n1213) );
XOR2_X1 U887 ( .A(n1148), .B(KEYINPUT9), .Z(n1236) );
NAND3_X1 U888 ( .A1(n1237), .A2(n1179), .A3(n1238), .ZN(n1148) );
XOR2_X1 U889 ( .A(n1239), .B(KEYINPUT57), .Z(n1238) );
AND4_X1 U890 ( .A1(n1057), .A2(n1058), .A3(n1240), .A4(n1059), .ZN(n1150) );
XOR2_X1 U891 ( .A(KEYINPUT54), .B(n1056), .Z(n1240) );
NOR3_X1 U892 ( .A1(n1107), .A2(n1086), .A3(n1075), .ZN(n1058) );
INV_X1 U893 ( .A(n1124), .ZN(n1212) );
NAND4_X1 U894 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1124) );
NOR3_X1 U895 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1244) );
NAND2_X1 U896 ( .A1(n1056), .A2(n1248), .ZN(n1243) );
XNOR2_X1 U897 ( .A(KEYINPUT29), .B(n1249), .ZN(n1248) );
OR3_X1 U898 ( .A1(n1250), .A2(n1093), .A3(n1239), .ZN(n1241) );
NOR2_X1 U899 ( .A1(n1179), .A2(n1057), .ZN(n1093) );
XNOR2_X1 U900 ( .A(n1123), .B(KEYINPUT18), .ZN(n1211) );
NAND2_X1 U901 ( .A1(n1251), .A2(n1252), .ZN(n1209) );
INV_X1 U902 ( .A(n1253), .ZN(n1252) );
NAND2_X1 U903 ( .A1(n1254), .A2(n1255), .ZN(n1251) );
NOR2_X1 U904 ( .A1(n1117), .A2(G952), .ZN(n1163) );
XOR2_X1 U905 ( .A(G146), .B(n1246), .Z(G48) );
AND2_X1 U906 ( .A1(n1179), .A2(n1256), .ZN(n1246) );
XOR2_X1 U907 ( .A(n1257), .B(n1242), .Z(G45) );
NAND3_X1 U908 ( .A1(n1092), .A2(n1258), .A3(n1259), .ZN(n1242) );
NOR3_X1 U909 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1259) );
XOR2_X1 U910 ( .A(G140), .B(n1123), .Z(G42) );
AND3_X1 U911 ( .A1(n1263), .A2(n1179), .A3(n1091), .ZN(n1123) );
NAND2_X1 U912 ( .A1(n1264), .A2(n1265), .ZN(G39) );
NAND2_X1 U913 ( .A1(n1247), .A2(n1266), .ZN(n1265) );
XOR2_X1 U914 ( .A(n1267), .B(KEYINPUT22), .Z(n1264) );
OR2_X1 U915 ( .A1(n1266), .A2(n1247), .ZN(n1267) );
NOR2_X1 U916 ( .A1(n1250), .A2(n1229), .ZN(n1247) );
INV_X1 U917 ( .A(G137), .ZN(n1266) );
XNOR2_X1 U918 ( .A(G134), .B(n1268), .ZN(G36) );
NOR2_X1 U919 ( .A1(n1269), .A2(KEYINPUT48), .ZN(n1268) );
NOR2_X1 U920 ( .A1(n1250), .A2(n1226), .ZN(n1269) );
XOR2_X1 U921 ( .A(G131), .B(n1270), .Z(G33) );
NOR3_X1 U922 ( .A1(n1271), .A2(KEYINPUT21), .A3(n1250), .ZN(n1270) );
INV_X1 U923 ( .A(n1263), .ZN(n1250) );
NOR4_X1 U924 ( .A1(n1087), .A2(n1261), .A3(n1107), .A4(n1086), .ZN(n1263) );
INV_X1 U925 ( .A(n1272), .ZN(n1261) );
NAND2_X1 U926 ( .A1(n1273), .A2(n1082), .ZN(n1087) );
XOR2_X1 U927 ( .A(G128), .B(n1245), .Z(G30) );
AND2_X1 U928 ( .A1(n1256), .A2(n1057), .ZN(n1245) );
AND4_X1 U929 ( .A1(n1274), .A2(n1258), .A3(n1106), .A4(n1272), .ZN(n1256) );
XOR2_X1 U930 ( .A(n1275), .B(n1216), .Z(G3) );
NAND3_X1 U931 ( .A1(n1092), .A2(n1258), .A3(n1276), .ZN(n1216) );
XOR2_X1 U932 ( .A(G125), .B(n1277), .Z(G27) );
NOR2_X1 U933 ( .A1(n1220), .A2(n1249), .ZN(n1277) );
NAND4_X1 U934 ( .A1(n1227), .A2(n1091), .A3(n1179), .A4(n1272), .ZN(n1249) );
NAND2_X1 U935 ( .A1(n1066), .A2(n1278), .ZN(n1272) );
NAND4_X1 U936 ( .A1(G953), .A2(G902), .A3(n1279), .A4(n1125), .ZN(n1278) );
INV_X1 U937 ( .A(G900), .ZN(n1125) );
XNOR2_X1 U938 ( .A(G122), .B(n1214), .ZN(G24) );
OR4_X1 U939 ( .A1(n1231), .A2(n1075), .A3(n1260), .A4(n1262), .ZN(n1214) );
NAND2_X1 U940 ( .A1(n1280), .A2(n1281), .ZN(n1075) );
XOR2_X1 U941 ( .A(G119), .B(n1282), .Z(G21) );
NOR2_X1 U942 ( .A1(n1229), .A2(n1231), .ZN(n1282) );
NAND4_X1 U943 ( .A1(n1274), .A2(n1262), .A3(n1283), .A4(n1106), .ZN(n1229) );
INV_X1 U944 ( .A(n1281), .ZN(n1106) );
XOR2_X1 U945 ( .A(n1280), .B(KEYINPUT55), .Z(n1274) );
XOR2_X1 U946 ( .A(n1284), .B(n1285), .Z(G18) );
NAND3_X1 U947 ( .A1(n1235), .A2(n1237), .A3(KEYINPUT7), .ZN(n1285) );
INV_X1 U948 ( .A(n1231), .ZN(n1237) );
INV_X1 U949 ( .A(n1226), .ZN(n1235) );
NAND2_X1 U950 ( .A1(n1092), .A2(n1057), .ZN(n1226) );
NOR2_X1 U951 ( .A1(n1069), .A2(n1260), .ZN(n1057) );
XOR2_X1 U952 ( .A(n1283), .B(KEYINPUT5), .Z(n1260) );
XOR2_X1 U953 ( .A(G113), .B(n1286), .Z(G15) );
NOR3_X1 U954 ( .A1(n1271), .A2(KEYINPUT4), .A3(n1231), .ZN(n1286) );
NAND3_X1 U955 ( .A1(n1056), .A2(n1059), .A3(n1227), .ZN(n1231) );
INV_X1 U956 ( .A(n1079), .ZN(n1227) );
NAND2_X1 U957 ( .A1(n1086), .A2(n1085), .ZN(n1079) );
INV_X1 U958 ( .A(n1220), .ZN(n1056) );
NAND2_X1 U959 ( .A1(n1092), .A2(n1179), .ZN(n1271) );
NOR2_X1 U960 ( .A1(n1071), .A2(n1262), .ZN(n1179) );
INV_X1 U961 ( .A(n1239), .ZN(n1092) );
NAND2_X1 U962 ( .A1(n1281), .A2(n1098), .ZN(n1239) );
XOR2_X1 U963 ( .A(n1287), .B(n1215), .Z(G12) );
NAND3_X1 U964 ( .A1(n1091), .A2(n1258), .A3(n1276), .ZN(n1215) );
NOR3_X1 U965 ( .A1(n1071), .A2(n1223), .A3(n1069), .ZN(n1276) );
INV_X1 U966 ( .A(n1262), .ZN(n1069) );
XOR2_X1 U967 ( .A(n1105), .B(n1288), .Z(n1262) );
NOR2_X1 U968 ( .A1(KEYINPUT38), .A2(n1104), .ZN(n1288) );
INV_X1 U969 ( .A(G475), .ZN(n1104) );
NAND2_X1 U970 ( .A1(n1289), .A2(n1290), .ZN(n1105) );
XOR2_X1 U971 ( .A(KEYINPUT52), .B(n1175), .Z(n1289) );
XNOR2_X1 U972 ( .A(n1291), .B(n1292), .ZN(n1175) );
XOR2_X1 U973 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U974 ( .A(G122), .B(G113), .Z(n1294) );
XOR2_X1 U975 ( .A(KEYINPUT49), .B(G143), .Z(n1293) );
XOR2_X1 U976 ( .A(n1295), .B(n1296), .Z(n1291) );
XNOR2_X1 U977 ( .A(G104), .B(n1297), .ZN(n1296) );
NAND2_X1 U978 ( .A1(n1298), .A2(G214), .ZN(n1297) );
XNOR2_X1 U979 ( .A(n1299), .B(n1300), .ZN(n1295) );
NOR2_X1 U980 ( .A1(G131), .A2(KEYINPUT6), .ZN(n1300) );
INV_X1 U981 ( .A(n1059), .ZN(n1223) );
NAND2_X1 U982 ( .A1(n1066), .A2(n1301), .ZN(n1059) );
NAND4_X1 U983 ( .A1(G953), .A2(G902), .A3(n1279), .A4(n1153), .ZN(n1301) );
INV_X1 U984 ( .A(G898), .ZN(n1153) );
NAND3_X1 U985 ( .A1(n1279), .A2(n1117), .A3(G952), .ZN(n1066) );
NAND2_X1 U986 ( .A1(G237), .A2(G234), .ZN(n1279) );
INV_X1 U987 ( .A(n1283), .ZN(n1071) );
XOR2_X1 U988 ( .A(n1113), .B(G478), .Z(n1283) );
OR2_X1 U989 ( .A1(n1171), .A2(G902), .ZN(n1113) );
XNOR2_X1 U990 ( .A(n1302), .B(n1303), .ZN(n1171) );
XNOR2_X1 U991 ( .A(n1304), .B(n1305), .ZN(n1303) );
XOR2_X1 U992 ( .A(n1306), .B(n1307), .Z(n1305) );
AND3_X1 U993 ( .A1(G234), .A2(n1117), .A3(G217), .ZN(n1307) );
NAND2_X1 U994 ( .A1(KEYINPUT45), .A2(G128), .ZN(n1306) );
XOR2_X1 U995 ( .A(n1308), .B(n1309), .Z(n1302) );
XOR2_X1 U996 ( .A(G143), .B(G122), .Z(n1309) );
XOR2_X1 U997 ( .A(G107), .B(n1284), .Z(n1308) );
NOR3_X1 U998 ( .A1(n1107), .A2(n1086), .A3(n1220), .ZN(n1258) );
NAND2_X1 U999 ( .A1(n1081), .A2(n1082), .ZN(n1220) );
NAND2_X1 U1000 ( .A1(G214), .A2(n1310), .ZN(n1082) );
INV_X1 U1001 ( .A(n1273), .ZN(n1081) );
XOR2_X1 U1002 ( .A(n1102), .B(n1311), .Z(n1273) );
NOR2_X1 U1003 ( .A1(KEYINPUT33), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U1004 ( .A(KEYINPUT24), .B(n1103), .ZN(n1312) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1310), .ZN(n1103) );
NAND2_X1 U1006 ( .A1(n1313), .A2(n1314), .ZN(n1310) );
INV_X1 U1007 ( .A(G237), .ZN(n1314) );
NAND2_X1 U1008 ( .A1(n1315), .A2(n1290), .ZN(n1102) );
XOR2_X1 U1009 ( .A(n1316), .B(n1317), .Z(n1315) );
NOR2_X1 U1010 ( .A1(KEYINPUT19), .A2(n1207), .ZN(n1317) );
XNOR2_X1 U1011 ( .A(n1154), .B(n1318), .ZN(n1207) );
XNOR2_X1 U1012 ( .A(n1319), .B(n1157), .ZN(n1318) );
XOR2_X1 U1013 ( .A(n1275), .B(n1320), .Z(n1157) );
INV_X1 U1014 ( .A(G101), .ZN(n1275) );
NAND2_X1 U1015 ( .A1(KEYINPUT26), .A2(n1158), .ZN(n1319) );
XNOR2_X1 U1016 ( .A(G113), .B(n1321), .ZN(n1158) );
XOR2_X1 U1017 ( .A(G119), .B(G116), .Z(n1321) );
XOR2_X1 U1018 ( .A(n1287), .B(n1322), .Z(n1154) );
NOR2_X1 U1019 ( .A1(G122), .A2(KEYINPUT2), .ZN(n1322) );
NOR2_X1 U1020 ( .A1(n1253), .A2(n1323), .ZN(n1316) );
NOR2_X1 U1021 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
XOR2_X1 U1022 ( .A(n1255), .B(KEYINPUT14), .Z(n1324) );
NOR2_X1 U1023 ( .A1(n1255), .A2(n1254), .ZN(n1253) );
INV_X1 U1024 ( .A(n1325), .ZN(n1254) );
XNOR2_X1 U1025 ( .A(n1188), .B(G125), .ZN(n1325) );
NAND2_X1 U1026 ( .A1(G224), .A2(n1117), .ZN(n1255) );
NOR2_X1 U1027 ( .A1(n1326), .A2(n1108), .ZN(n1086) );
NOR2_X1 U1028 ( .A1(n1110), .A2(G469), .ZN(n1108) );
AND2_X1 U1029 ( .A1(n1327), .A2(n1110), .ZN(n1326) );
NAND2_X1 U1030 ( .A1(n1328), .A2(n1290), .ZN(n1110) );
XOR2_X1 U1031 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1032 ( .A(n1331), .B(n1200), .Z(n1330) );
XOR2_X1 U1033 ( .A(n1332), .B(n1129), .Z(n1200) );
XOR2_X1 U1034 ( .A(G128), .B(n1333), .Z(n1129) );
NOR2_X1 U1035 ( .A1(KEYINPUT20), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1036 ( .A(n1257), .B(n1335), .Z(n1334) );
NAND2_X1 U1037 ( .A1(KEYINPUT31), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1038 ( .A(n1337), .B(G101), .Z(n1332) );
NAND2_X1 U1039 ( .A1(KEYINPUT58), .A2(n1320), .ZN(n1337) );
XNOR2_X1 U1040 ( .A(G104), .B(G107), .ZN(n1320) );
NAND2_X1 U1041 ( .A1(KEYINPUT10), .A2(n1338), .ZN(n1331) );
XNOR2_X1 U1042 ( .A(n1339), .B(n1205), .ZN(n1338) );
NAND2_X1 U1043 ( .A1(G227), .A2(n1117), .ZN(n1205) );
NOR2_X1 U1044 ( .A1(n1204), .A2(n1340), .ZN(n1339) );
XOR2_X1 U1045 ( .A(n1341), .B(KEYINPUT44), .Z(n1340) );
NAND2_X1 U1046 ( .A1(n1342), .A2(n1287), .ZN(n1341) );
XOR2_X1 U1047 ( .A(KEYINPUT51), .B(G140), .Z(n1342) );
NOR2_X1 U1048 ( .A1(n1287), .A2(G140), .ZN(n1204) );
NAND2_X1 U1049 ( .A1(n1343), .A2(n1344), .ZN(n1329) );
NAND2_X1 U1050 ( .A1(KEYINPUT11), .A2(n1185), .ZN(n1344) );
OR2_X1 U1051 ( .A1(KEYINPUT32), .A2(n1185), .ZN(n1343) );
XNOR2_X1 U1052 ( .A(G469), .B(KEYINPUT8), .ZN(n1327) );
INV_X1 U1053 ( .A(n1085), .ZN(n1107) );
NAND2_X1 U1054 ( .A1(G221), .A2(n1345), .ZN(n1085) );
NOR2_X1 U1055 ( .A1(n1098), .A2(n1281), .ZN(n1091) );
XOR2_X1 U1056 ( .A(n1346), .B(n1168), .Z(n1281) );
AND2_X1 U1057 ( .A1(G217), .A2(n1345), .ZN(n1168) );
NAND2_X1 U1058 ( .A1(n1313), .A2(n1347), .ZN(n1345) );
XOR2_X1 U1059 ( .A(KEYINPUT60), .B(G234), .Z(n1347) );
XOR2_X1 U1060 ( .A(n1290), .B(KEYINPUT42), .Z(n1313) );
OR2_X1 U1061 ( .A1(n1166), .A2(G902), .ZN(n1346) );
XOR2_X1 U1062 ( .A(n1348), .B(n1349), .Z(n1166) );
XOR2_X1 U1063 ( .A(n1350), .B(n1351), .Z(n1349) );
XOR2_X1 U1064 ( .A(G119), .B(G110), .Z(n1351) );
XOR2_X1 U1065 ( .A(KEYINPUT41), .B(G137), .Z(n1350) );
XOR2_X1 U1066 ( .A(n1352), .B(n1299), .Z(n1348) );
XNOR2_X1 U1067 ( .A(n1137), .B(n1353), .ZN(n1299) );
XOR2_X1 U1068 ( .A(G146), .B(G140), .Z(n1353) );
INV_X1 U1069 ( .A(G125), .ZN(n1137) );
XOR2_X1 U1070 ( .A(n1354), .B(n1355), .Z(n1352) );
AND3_X1 U1071 ( .A1(G221), .A2(n1117), .A3(G234), .ZN(n1355) );
INV_X1 U1072 ( .A(G953), .ZN(n1117) );
NAND2_X1 U1073 ( .A1(KEYINPUT50), .A2(n1356), .ZN(n1354) );
XOR2_X1 U1074 ( .A(KEYINPUT25), .B(G128), .Z(n1356) );
INV_X1 U1075 ( .A(n1280), .ZN(n1098) );
XOR2_X1 U1076 ( .A(n1357), .B(G472), .Z(n1280) );
NAND2_X1 U1077 ( .A1(n1358), .A2(n1290), .ZN(n1357) );
INV_X1 U1078 ( .A(G902), .ZN(n1290) );
XOR2_X1 U1079 ( .A(n1359), .B(n1183), .Z(n1358) );
XOR2_X1 U1080 ( .A(n1360), .B(G101), .Z(n1183) );
NAND2_X1 U1081 ( .A1(n1298), .A2(G210), .ZN(n1360) );
NOR2_X1 U1082 ( .A1(G953), .A2(G237), .ZN(n1298) );
NAND2_X1 U1083 ( .A1(n1361), .A2(n1362), .ZN(n1359) );
NAND2_X1 U1084 ( .A1(n1189), .A2(n1363), .ZN(n1362) );
XOR2_X1 U1085 ( .A(n1364), .B(KEYINPUT40), .Z(n1361) );
OR2_X1 U1086 ( .A1(n1363), .A2(n1189), .ZN(n1364) );
AND2_X1 U1087 ( .A1(n1365), .A2(n1366), .ZN(n1189) );
NAND2_X1 U1088 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
INV_X1 U1089 ( .A(G113), .ZN(n1368) );
XOR2_X1 U1090 ( .A(n1284), .B(n1369), .Z(n1367) );
INV_X1 U1091 ( .A(G116), .ZN(n1284) );
NAND2_X1 U1092 ( .A1(G113), .A2(n1370), .ZN(n1365) );
XOR2_X1 U1093 ( .A(n1369), .B(G116), .Z(n1370) );
NAND2_X1 U1094 ( .A1(KEYINPUT46), .A2(n1371), .ZN(n1369) );
INV_X1 U1095 ( .A(G119), .ZN(n1371) );
XNOR2_X1 U1096 ( .A(n1372), .B(n1373), .ZN(n1363) );
INV_X1 U1097 ( .A(n1188), .ZN(n1373) );
XOR2_X1 U1098 ( .A(n1374), .B(G128), .Z(n1188) );
NAND3_X1 U1099 ( .A1(n1375), .A2(n1376), .A3(n1377), .ZN(n1374) );
NAND2_X1 U1100 ( .A1(G146), .A2(n1257), .ZN(n1377) );
NAND2_X1 U1101 ( .A1(n1378), .A2(n1379), .ZN(n1376) );
INV_X1 U1102 ( .A(KEYINPUT28), .ZN(n1379) );
NAND2_X1 U1103 ( .A1(n1380), .A2(G143), .ZN(n1378) );
XOR2_X1 U1104 ( .A(KEYINPUT59), .B(n1336), .Z(n1380) );
INV_X1 U1105 ( .A(G146), .ZN(n1336) );
NAND2_X1 U1106 ( .A1(KEYINPUT28), .A2(n1381), .ZN(n1375) );
NAND2_X1 U1107 ( .A1(n1382), .A2(n1383), .ZN(n1381) );
OR3_X1 U1108 ( .A1(n1257), .A2(G146), .A3(KEYINPUT59), .ZN(n1383) );
INV_X1 U1109 ( .A(G143), .ZN(n1257) );
NAND2_X1 U1110 ( .A1(KEYINPUT59), .A2(G146), .ZN(n1382) );
NAND2_X1 U1111 ( .A1(KEYINPUT53), .A2(n1185), .ZN(n1372) );
XOR2_X1 U1112 ( .A(G131), .B(n1128), .Z(n1185) );
XOR2_X1 U1113 ( .A(G137), .B(n1304), .Z(n1128) );
XOR2_X1 U1114 ( .A(G134), .B(KEYINPUT0), .Z(n1304) );
INV_X1 U1115 ( .A(G110), .ZN(n1287) );
endmodule


