//Key = 1100010110011110110011101011110101000111100110010000001010101110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417, n1418, n1419;

XNOR2_X1 U777 ( .A(G107), .B(n1077), .ZN(G9) );
NOR2_X1 U778 ( .A1(n1078), .A2(n1079), .ZN(G75) );
AND3_X1 U779 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NOR3_X1 U780 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1078) );
XOR2_X1 U781 ( .A(n1086), .B(KEYINPUT33), .Z(n1084) );
NAND4_X1 U782 ( .A1(n1087), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1086) );
NOR2_X1 U783 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
XNOR2_X1 U784 ( .A(n1093), .B(KEYINPUT46), .ZN(n1091) );
NAND3_X1 U785 ( .A1(n1094), .A2(n1081), .A3(n1080), .ZN(n1083) );
NAND4_X1 U786 ( .A1(n1095), .A2(n1087), .A3(n1096), .A4(n1097), .ZN(n1080) );
NOR4_X1 U787 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
XNOR2_X1 U788 ( .A(G478), .B(n1102), .ZN(n1100) );
NOR2_X1 U789 ( .A1(n1103), .A2(KEYINPUT25), .ZN(n1102) );
NOR2_X1 U790 ( .A1(n1104), .A2(n1105), .ZN(n1099) );
XNOR2_X1 U791 ( .A(G472), .B(KEYINPUT52), .ZN(n1105) );
INV_X1 U792 ( .A(n1106), .ZN(n1104) );
XOR2_X1 U793 ( .A(n1107), .B(n1108), .Z(n1096) );
NOR2_X1 U794 ( .A1(KEYINPUT53), .A2(n1109), .ZN(n1108) );
XNOR2_X1 U795 ( .A(n1110), .B(n1111), .ZN(n1095) );
NAND2_X1 U796 ( .A1(n1093), .A2(n1112), .ZN(n1094) );
NAND2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND3_X1 U798 ( .A1(n1090), .A2(n1115), .A3(n1116), .ZN(n1114) );
NAND2_X1 U799 ( .A1(n1117), .A2(n1118), .ZN(n1115) );
NAND2_X1 U800 ( .A1(n1087), .A2(n1119), .ZN(n1118) );
OR2_X1 U801 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U802 ( .A1(n1088), .A2(n1122), .ZN(n1117) );
NAND2_X1 U803 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
OR3_X1 U804 ( .A1(n1125), .A2(KEYINPUT18), .A3(n1126), .ZN(n1124) );
NAND3_X1 U805 ( .A1(n1088), .A2(n1127), .A3(n1087), .ZN(n1113) );
NAND2_X1 U806 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND3_X1 U807 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1129) );
XNOR2_X1 U808 ( .A(n1090), .B(KEYINPUT60), .ZN(n1132) );
NAND2_X1 U809 ( .A1(n1116), .A2(n1133), .ZN(n1128) );
NAND3_X1 U810 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1133) );
NAND2_X1 U811 ( .A1(KEYINPUT18), .A2(n1090), .ZN(n1136) );
INV_X1 U812 ( .A(n1137), .ZN(n1093) );
XOR2_X1 U813 ( .A(n1138), .B(n1139), .Z(G72) );
NOR2_X1 U814 ( .A1(n1140), .A2(n1081), .ZN(n1139) );
NOR2_X1 U815 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XOR2_X1 U816 ( .A(KEYINPUT14), .B(G227), .Z(n1142) );
NAND2_X1 U817 ( .A1(n1143), .A2(n1144), .ZN(n1138) );
NAND3_X1 U818 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(n1144) );
NAND2_X1 U819 ( .A1(G953), .A2(n1141), .ZN(n1146) );
OR2_X1 U820 ( .A1(n1145), .A2(n1147), .ZN(n1143) );
NAND2_X1 U821 ( .A1(n1081), .A2(n1148), .ZN(n1147) );
NAND3_X1 U822 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1148) );
XOR2_X1 U823 ( .A(KEYINPUT32), .B(n1152), .Z(n1150) );
XNOR2_X1 U824 ( .A(KEYINPUT61), .B(n1153), .ZN(n1149) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1145) );
NOR3_X1 U826 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1155) );
NOR2_X1 U827 ( .A1(KEYINPUT24), .A2(n1159), .ZN(n1158) );
INV_X1 U828 ( .A(n1160), .ZN(n1159) );
AND3_X1 U829 ( .A1(KEYINPUT24), .A2(n1161), .A3(n1162), .ZN(n1157) );
NOR2_X1 U830 ( .A1(n1162), .A2(n1161), .ZN(n1156) );
NOR2_X1 U831 ( .A1(KEYINPUT48), .A2(n1160), .ZN(n1162) );
XOR2_X1 U832 ( .A(G125), .B(KEYINPUT55), .Z(n1160) );
NAND2_X1 U833 ( .A1(n1163), .A2(n1164), .ZN(n1154) );
OR2_X1 U834 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XOR2_X1 U835 ( .A(n1167), .B(KEYINPUT51), .Z(n1163) );
NAND2_X1 U836 ( .A1(n1168), .A2(n1165), .ZN(n1167) );
XOR2_X1 U837 ( .A(n1169), .B(n1170), .Z(n1165) );
XNOR2_X1 U838 ( .A(n1166), .B(KEYINPUT37), .ZN(n1168) );
XOR2_X1 U839 ( .A(n1171), .B(n1172), .Z(G69) );
NOR2_X1 U840 ( .A1(n1173), .A2(n1081), .ZN(n1172) );
AND2_X1 U841 ( .A1(G224), .A2(G898), .ZN(n1173) );
NAND2_X1 U842 ( .A1(n1174), .A2(n1175), .ZN(n1171) );
NAND2_X1 U843 ( .A1(n1176), .A2(n1081), .ZN(n1175) );
XOR2_X1 U844 ( .A(n1177), .B(n1178), .Z(n1176) );
OR3_X1 U845 ( .A1(n1179), .A2(n1178), .A3(n1081), .ZN(n1174) );
XOR2_X1 U846 ( .A(n1180), .B(n1181), .Z(n1178) );
NOR2_X1 U847 ( .A1(n1182), .A2(n1183), .ZN(G66) );
XOR2_X1 U848 ( .A(n1184), .B(n1185), .Z(n1183) );
AND2_X1 U849 ( .A1(G217), .A2(n1186), .ZN(n1184) );
NOR2_X1 U850 ( .A1(n1182), .A2(n1187), .ZN(G63) );
XOR2_X1 U851 ( .A(n1188), .B(n1189), .Z(n1187) );
NOR2_X1 U852 ( .A1(n1190), .A2(n1191), .ZN(n1188) );
NOR2_X1 U853 ( .A1(n1182), .A2(n1192), .ZN(G60) );
XOR2_X1 U854 ( .A(n1193), .B(n1194), .Z(n1192) );
NAND3_X1 U855 ( .A1(n1186), .A2(G475), .A3(KEYINPUT47), .ZN(n1193) );
XOR2_X1 U856 ( .A(G104), .B(n1195), .Z(G6) );
NOR2_X1 U857 ( .A1(n1182), .A2(n1196), .ZN(G57) );
XOR2_X1 U858 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U859 ( .A(n1199), .B(n1200), .Z(n1198) );
XOR2_X1 U860 ( .A(n1201), .B(n1202), .Z(n1197) );
AND2_X1 U861 ( .A1(G472), .A2(n1186), .ZN(n1202) );
NAND3_X1 U862 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1201) );
NAND2_X1 U863 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U864 ( .A1(KEYINPUT57), .A2(n1208), .ZN(n1204) );
NAND2_X1 U865 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XNOR2_X1 U866 ( .A(KEYINPUT49), .B(n1206), .ZN(n1209) );
NAND2_X1 U867 ( .A1(n1211), .A2(n1212), .ZN(n1203) );
INV_X1 U868 ( .A(KEYINPUT57), .ZN(n1212) );
NAND2_X1 U869 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
OR3_X1 U870 ( .A1(n1206), .A2(n1207), .A3(KEYINPUT49), .ZN(n1214) );
NAND2_X1 U871 ( .A1(KEYINPUT49), .A2(n1206), .ZN(n1213) );
NOR3_X1 U872 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(G54) );
AND2_X1 U873 ( .A1(KEYINPUT12), .A2(n1182), .ZN(n1217) );
NOR3_X1 U874 ( .A1(KEYINPUT12), .A2(n1081), .A3(n1082), .ZN(n1216) );
INV_X1 U875 ( .A(G952), .ZN(n1082) );
XOR2_X1 U876 ( .A(n1218), .B(n1219), .Z(n1215) );
XOR2_X1 U877 ( .A(n1220), .B(n1221), .Z(n1219) );
NAND2_X1 U878 ( .A1(KEYINPUT1), .A2(n1222), .ZN(n1221) );
NAND3_X1 U879 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1220) );
NAND2_X1 U880 ( .A1(n1226), .A2(n1207), .ZN(n1225) );
NAND2_X1 U881 ( .A1(n1227), .A2(n1228), .ZN(n1224) );
INV_X1 U882 ( .A(KEYINPUT21), .ZN(n1228) );
NAND2_X1 U883 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
XNOR2_X1 U884 ( .A(KEYINPUT35), .B(n1207), .ZN(n1229) );
NAND2_X1 U885 ( .A1(KEYINPUT21), .A2(n1231), .ZN(n1223) );
NAND2_X1 U886 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
OR3_X1 U887 ( .A1(n1226), .A2(n1207), .A3(KEYINPUT35), .ZN(n1233) );
INV_X1 U888 ( .A(n1230), .ZN(n1226) );
XOR2_X1 U889 ( .A(n1166), .B(n1234), .Z(n1230) );
NAND2_X1 U890 ( .A1(KEYINPUT35), .A2(n1207), .ZN(n1232) );
XOR2_X1 U891 ( .A(n1235), .B(n1236), .Z(n1218) );
AND2_X1 U892 ( .A1(G469), .A2(n1186), .ZN(n1236) );
INV_X1 U893 ( .A(n1191), .ZN(n1186) );
NOR2_X1 U894 ( .A1(n1182), .A2(n1237), .ZN(G51) );
XOR2_X1 U895 ( .A(n1238), .B(n1239), .Z(n1237) );
NOR2_X1 U896 ( .A1(n1240), .A2(n1191), .ZN(n1239) );
NAND2_X1 U897 ( .A1(G902), .A2(n1085), .ZN(n1191) );
NAND4_X1 U898 ( .A1(n1152), .A2(n1177), .A3(n1151), .A4(n1153), .ZN(n1085) );
AND3_X1 U899 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1151) );
NAND2_X1 U900 ( .A1(n1116), .A2(n1244), .ZN(n1243) );
XNOR2_X1 U901 ( .A(KEYINPUT9), .B(n1245), .ZN(n1244) );
AND4_X1 U902 ( .A1(n1246), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1177) );
NOR4_X1 U903 ( .A1(n1195), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1249) );
NOR2_X1 U904 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NOR2_X1 U905 ( .A1(n1255), .A2(n1256), .ZN(n1251) );
NOR2_X1 U906 ( .A1(n1257), .A2(n1258), .ZN(n1255) );
NOR3_X1 U907 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1258) );
NOR3_X1 U908 ( .A1(n1262), .A2(n1123), .A3(n1135), .ZN(n1257) );
INV_X1 U909 ( .A(n1263), .ZN(n1135) );
NAND3_X1 U910 ( .A1(n1092), .A2(n1254), .A3(n1264), .ZN(n1262) );
INV_X1 U911 ( .A(KEYINPUT43), .ZN(n1254) );
AND3_X1 U912 ( .A1(n1090), .A2(n1265), .A3(n1120), .ZN(n1195) );
AND2_X1 U913 ( .A1(n1077), .A2(n1266), .ZN(n1248) );
NAND3_X1 U914 ( .A1(n1090), .A2(n1265), .A3(n1121), .ZN(n1077) );
AND3_X1 U915 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(n1152) );
NAND2_X1 U916 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U917 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NAND4_X1 U918 ( .A1(n1274), .A2(n1275), .A3(n1276), .A4(n1277), .ZN(n1273) );
XOR2_X1 U919 ( .A(n1278), .B(n1279), .Z(n1238) );
NOR2_X1 U920 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
XOR2_X1 U921 ( .A(KEYINPUT6), .B(n1282), .Z(n1281) );
NOR2_X1 U922 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
AND2_X1 U923 ( .A1(n1283), .A2(n1284), .ZN(n1280) );
NAND2_X1 U924 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND2_X1 U925 ( .A1(G125), .A2(n1287), .ZN(n1286) );
XOR2_X1 U926 ( .A(n1288), .B(KEYINPUT59), .Z(n1285) );
NAND2_X1 U927 ( .A1(n1206), .A2(n1289), .ZN(n1288) );
INV_X1 U928 ( .A(n1287), .ZN(n1206) );
NOR2_X1 U929 ( .A1(n1081), .A2(G952), .ZN(n1182) );
XNOR2_X1 U930 ( .A(G146), .B(n1267), .ZN(G48) );
NAND3_X1 U931 ( .A1(n1290), .A2(n1275), .A3(n1120), .ZN(n1267) );
XOR2_X1 U932 ( .A(n1291), .B(n1292), .Z(G45) );
XNOR2_X1 U933 ( .A(KEYINPUT38), .B(n1293), .ZN(n1292) );
NAND3_X1 U934 ( .A1(KEYINPUT31), .A2(n1294), .A3(n1295), .ZN(n1291) );
NOR3_X1 U935 ( .A1(n1092), .A2(n1296), .A3(n1297), .ZN(n1295) );
XNOR2_X1 U936 ( .A(n1161), .B(n1298), .ZN(G42) );
NOR3_X1 U937 ( .A1(n1272), .A2(KEYINPUT3), .A3(n1299), .ZN(n1298) );
NAND3_X1 U938 ( .A1(n1120), .A2(n1116), .A3(n1263), .ZN(n1272) );
XNOR2_X1 U939 ( .A(G137), .B(n1268), .ZN(G39) );
NAND3_X1 U940 ( .A1(n1290), .A2(n1116), .A3(n1088), .ZN(n1268) );
XNOR2_X1 U941 ( .A(G134), .B(n1153), .ZN(G36) );
NAND3_X1 U942 ( .A1(n1116), .A2(n1121), .A3(n1294), .ZN(n1153) );
INV_X1 U943 ( .A(n1101), .ZN(n1116) );
XOR2_X1 U944 ( .A(G131), .B(n1300), .Z(G33) );
NOR2_X1 U945 ( .A1(n1101), .A2(n1245), .ZN(n1300) );
NAND2_X1 U946 ( .A1(n1294), .A2(n1120), .ZN(n1245) );
NOR2_X1 U947 ( .A1(n1134), .A2(n1299), .ZN(n1294) );
INV_X1 U948 ( .A(n1274), .ZN(n1134) );
NAND2_X1 U949 ( .A1(n1130), .A2(n1301), .ZN(n1101) );
XNOR2_X1 U950 ( .A(G128), .B(n1241), .ZN(G30) );
NAND3_X1 U951 ( .A1(n1121), .A2(n1275), .A3(n1290), .ZN(n1241) );
NOR3_X1 U952 ( .A1(n1261), .A2(n1260), .A3(n1299), .ZN(n1290) );
INV_X1 U953 ( .A(n1270), .ZN(n1299) );
NOR2_X1 U954 ( .A1(n1123), .A2(n1302), .ZN(n1270) );
XOR2_X1 U955 ( .A(n1303), .B(G101), .Z(G3) );
NAND2_X1 U956 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND2_X1 U957 ( .A1(n1250), .A2(n1306), .ZN(n1305) );
INV_X1 U958 ( .A(KEYINPUT4), .ZN(n1306) );
NOR2_X1 U959 ( .A1(n1307), .A2(n1092), .ZN(n1250) );
NAND3_X1 U960 ( .A1(n1275), .A2(n1307), .A3(KEYINPUT4), .ZN(n1304) );
NAND4_X1 U961 ( .A1(n1274), .A2(n1088), .A3(n1308), .A4(n1264), .ZN(n1307) );
XNOR2_X1 U962 ( .A(G125), .B(n1242), .ZN(G27) );
NAND4_X1 U963 ( .A1(n1087), .A2(n1263), .A3(n1309), .A4(n1120), .ZN(n1242) );
NOR2_X1 U964 ( .A1(n1302), .A2(n1092), .ZN(n1309) );
INV_X1 U965 ( .A(n1275), .ZN(n1092) );
AND2_X1 U966 ( .A1(n1137), .A2(n1310), .ZN(n1302) );
NAND4_X1 U967 ( .A1(G953), .A2(G902), .A3(n1311), .A4(n1141), .ZN(n1310) );
INV_X1 U968 ( .A(G900), .ZN(n1141) );
NAND2_X1 U969 ( .A1(n1312), .A2(n1313), .ZN(G24) );
OR2_X1 U970 ( .A1(n1314), .A2(G122), .ZN(n1313) );
NAND2_X1 U971 ( .A1(G122), .A2(n1315), .ZN(n1312) );
NAND2_X1 U972 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
OR2_X1 U973 ( .A1(n1246), .A2(KEYINPUT54), .ZN(n1317) );
NAND2_X1 U974 ( .A1(KEYINPUT54), .A2(n1314), .ZN(n1316) );
NAND2_X1 U975 ( .A1(KEYINPUT26), .A2(n1318), .ZN(n1314) );
INV_X1 U976 ( .A(n1246), .ZN(n1318) );
NAND4_X1 U977 ( .A1(n1319), .A2(n1090), .A3(n1276), .A4(n1277), .ZN(n1246) );
NOR2_X1 U978 ( .A1(n1320), .A2(n1321), .ZN(n1090) );
XNOR2_X1 U979 ( .A(G119), .B(n1322), .ZN(G21) );
NAND3_X1 U980 ( .A1(KEYINPUT11), .A2(n1319), .A3(n1323), .ZN(n1322) );
NOR3_X1 U981 ( .A1(n1256), .A2(n1260), .A3(n1261), .ZN(n1323) );
INV_X1 U982 ( .A(n1088), .ZN(n1256) );
XNOR2_X1 U983 ( .A(G116), .B(n1247), .ZN(G18) );
NAND3_X1 U984 ( .A1(n1274), .A2(n1121), .A3(n1319), .ZN(n1247) );
NOR2_X1 U985 ( .A1(n1276), .A2(n1296), .ZN(n1121) );
INV_X1 U986 ( .A(n1277), .ZN(n1296) );
XNOR2_X1 U987 ( .A(G113), .B(n1266), .ZN(G15) );
NAND3_X1 U988 ( .A1(n1274), .A2(n1120), .A3(n1319), .ZN(n1266) );
INV_X1 U989 ( .A(n1259), .ZN(n1319) );
NAND3_X1 U990 ( .A1(n1275), .A2(n1264), .A3(n1087), .ZN(n1259) );
NOR2_X1 U991 ( .A1(n1125), .A2(n1324), .ZN(n1087) );
INV_X1 U992 ( .A(n1126), .ZN(n1324) );
NOR2_X1 U993 ( .A1(n1277), .A2(n1297), .ZN(n1120) );
INV_X1 U994 ( .A(n1276), .ZN(n1297) );
NOR2_X1 U995 ( .A1(n1321), .A2(n1260), .ZN(n1274) );
INV_X1 U996 ( .A(n1261), .ZN(n1321) );
XNOR2_X1 U997 ( .A(G110), .B(n1253), .ZN(G12) );
NAND3_X1 U998 ( .A1(n1088), .A2(n1265), .A3(n1263), .ZN(n1253) );
NOR2_X1 U999 ( .A1(n1261), .A2(n1320), .ZN(n1263) );
INV_X1 U1000 ( .A(n1260), .ZN(n1320) );
NOR2_X1 U1001 ( .A1(n1325), .A2(n1098), .ZN(n1260) );
NOR2_X1 U1002 ( .A1(n1106), .A2(G472), .ZN(n1098) );
AND2_X1 U1003 ( .A1(G472), .A2(n1106), .ZN(n1325) );
NAND2_X1 U1004 ( .A1(n1326), .A2(n1327), .ZN(n1106) );
XOR2_X1 U1005 ( .A(n1328), .B(n1329), .Z(n1326) );
XNOR2_X1 U1006 ( .A(n1330), .B(n1200), .ZN(n1329) );
XNOR2_X1 U1007 ( .A(n1331), .B(n1332), .ZN(n1200) );
NAND3_X1 U1008 ( .A1(n1333), .A2(n1081), .A3(G210), .ZN(n1331) );
XNOR2_X1 U1009 ( .A(n1334), .B(n1207), .ZN(n1328) );
INV_X1 U1010 ( .A(n1210), .ZN(n1207) );
XNOR2_X1 U1011 ( .A(n1335), .B(n1336), .ZN(n1334) );
XOR2_X1 U1012 ( .A(n1337), .B(n1107), .Z(n1261) );
NAND2_X1 U1013 ( .A1(n1338), .A2(G217), .ZN(n1107) );
XOR2_X1 U1014 ( .A(n1339), .B(KEYINPUT50), .Z(n1338) );
NAND2_X1 U1015 ( .A1(KEYINPUT0), .A2(n1109), .ZN(n1337) );
OR2_X1 U1016 ( .A1(n1185), .A2(G902), .ZN(n1109) );
XNOR2_X1 U1017 ( .A(n1340), .B(n1341), .ZN(n1185) );
XOR2_X1 U1018 ( .A(n1342), .B(n1343), .Z(n1341) );
XNOR2_X1 U1019 ( .A(n1336), .B(G110), .ZN(n1343) );
XNOR2_X1 U1020 ( .A(G137), .B(n1289), .ZN(n1342) );
XNOR2_X1 U1021 ( .A(n1344), .B(n1345), .ZN(n1340) );
XNOR2_X1 U1022 ( .A(n1346), .B(n1347), .ZN(n1345) );
NOR2_X1 U1023 ( .A1(KEYINPUT19), .A2(G140), .ZN(n1347) );
NAND4_X1 U1024 ( .A1(KEYINPUT27), .A2(G221), .A3(G234), .A4(n1081), .ZN(n1346) );
AND3_X1 U1025 ( .A1(n1275), .A2(n1264), .A3(n1308), .ZN(n1265) );
INV_X1 U1026 ( .A(n1123), .ZN(n1308) );
NAND2_X1 U1027 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NAND2_X1 U1028 ( .A1(G221), .A2(n1339), .ZN(n1126) );
NAND2_X1 U1029 ( .A1(n1348), .A2(n1327), .ZN(n1339) );
XNOR2_X1 U1030 ( .A(KEYINPUT16), .B(n1349), .ZN(n1348) );
XNOR2_X1 U1031 ( .A(n1350), .B(G469), .ZN(n1125) );
NAND2_X1 U1032 ( .A1(n1351), .A2(n1327), .ZN(n1350) );
XOR2_X1 U1033 ( .A(n1352), .B(n1353), .Z(n1351) );
XNOR2_X1 U1034 ( .A(n1354), .B(n1222), .ZN(n1353) );
XNOR2_X1 U1035 ( .A(G110), .B(n1161), .ZN(n1222) );
INV_X1 U1036 ( .A(G140), .ZN(n1161) );
NAND2_X1 U1037 ( .A1(KEYINPUT7), .A2(n1210), .ZN(n1354) );
XNOR2_X1 U1038 ( .A(n1355), .B(n1170), .ZN(n1210) );
XOR2_X1 U1039 ( .A(G131), .B(KEYINPUT44), .Z(n1170) );
NAND2_X1 U1040 ( .A1(n1356), .A2(KEYINPUT58), .ZN(n1355) );
XNOR2_X1 U1041 ( .A(n1357), .B(n1358), .ZN(n1356) );
INV_X1 U1042 ( .A(n1169), .ZN(n1358) );
XOR2_X1 U1043 ( .A(G134), .B(G137), .Z(n1169) );
XNOR2_X1 U1044 ( .A(KEYINPUT29), .B(KEYINPUT23), .ZN(n1357) );
XNOR2_X1 U1045 ( .A(n1359), .B(n1235), .ZN(n1352) );
NAND2_X1 U1046 ( .A1(G227), .A2(n1081), .ZN(n1235) );
NAND2_X1 U1047 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
OR2_X1 U1048 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
XOR2_X1 U1049 ( .A(n1364), .B(KEYINPUT45), .Z(n1360) );
NAND2_X1 U1050 ( .A1(n1363), .A2(n1362), .ZN(n1364) );
XOR2_X1 U1051 ( .A(n1234), .B(KEYINPUT34), .Z(n1362) );
XOR2_X1 U1052 ( .A(G101), .B(n1365), .Z(n1234) );
XNOR2_X1 U1053 ( .A(n1366), .B(G104), .ZN(n1365) );
INV_X1 U1054 ( .A(n1166), .ZN(n1363) );
XNOR2_X1 U1055 ( .A(n1367), .B(n1368), .ZN(n1166) );
XOR2_X1 U1056 ( .A(n1369), .B(n1344), .Z(n1368) );
XNOR2_X1 U1057 ( .A(G128), .B(n1370), .ZN(n1344) );
NOR2_X1 U1058 ( .A1(KEYINPUT30), .A2(n1293), .ZN(n1369) );
XNOR2_X1 U1059 ( .A(KEYINPUT36), .B(KEYINPUT13), .ZN(n1367) );
NAND2_X1 U1060 ( .A1(n1137), .A2(n1371), .ZN(n1264) );
NAND4_X1 U1061 ( .A1(G953), .A2(G902), .A3(n1311), .A4(n1179), .ZN(n1371) );
INV_X1 U1062 ( .A(G898), .ZN(n1179) );
NAND3_X1 U1063 ( .A1(n1311), .A2(n1081), .A3(n1372), .ZN(n1137) );
XNOR2_X1 U1064 ( .A(G952), .B(KEYINPUT39), .ZN(n1372) );
NAND2_X1 U1065 ( .A1(G237), .A2(n1349), .ZN(n1311) );
XNOR2_X1 U1066 ( .A(G234), .B(KEYINPUT40), .ZN(n1349) );
NOR2_X1 U1067 ( .A1(n1130), .A2(n1131), .ZN(n1275) );
INV_X1 U1068 ( .A(n1301), .ZN(n1131) );
NAND2_X1 U1069 ( .A1(G214), .A2(n1373), .ZN(n1301) );
XNOR2_X1 U1070 ( .A(n1374), .B(n1240), .ZN(n1130) );
NAND2_X1 U1071 ( .A1(G210), .A2(n1373), .ZN(n1240) );
NAND2_X1 U1072 ( .A1(n1333), .A2(n1327), .ZN(n1373) );
NAND2_X1 U1073 ( .A1(n1375), .A2(n1327), .ZN(n1374) );
XOR2_X1 U1074 ( .A(n1376), .B(n1377), .Z(n1375) );
XNOR2_X1 U1075 ( .A(n1283), .B(n1287), .ZN(n1377) );
XNOR2_X1 U1076 ( .A(n1335), .B(G128), .ZN(n1287) );
NAND2_X1 U1077 ( .A1(n1378), .A2(n1379), .ZN(n1335) );
NAND2_X1 U1078 ( .A1(G143), .A2(n1370), .ZN(n1379) );
XOR2_X1 U1079 ( .A(KEYINPUT8), .B(n1380), .Z(n1378) );
NOR2_X1 U1080 ( .A1(G143), .A2(n1370), .ZN(n1380) );
NAND2_X1 U1081 ( .A1(G224), .A2(n1081), .ZN(n1283) );
XNOR2_X1 U1082 ( .A(G125), .B(n1278), .ZN(n1376) );
NAND2_X1 U1083 ( .A1(n1381), .A2(n1382), .ZN(n1278) );
NAND2_X1 U1084 ( .A1(n1181), .A2(n1383), .ZN(n1382) );
XOR2_X1 U1085 ( .A(KEYINPUT20), .B(n1384), .Z(n1381) );
NOR2_X1 U1086 ( .A1(n1181), .A2(n1383), .ZN(n1384) );
XOR2_X1 U1087 ( .A(n1180), .B(KEYINPUT22), .Z(n1383) );
XOR2_X1 U1088 ( .A(n1385), .B(n1386), .Z(n1180) );
XNOR2_X1 U1089 ( .A(n1387), .B(n1332), .ZN(n1386) );
XOR2_X1 U1090 ( .A(G101), .B(G113), .Z(n1332) );
NAND2_X1 U1091 ( .A1(n1388), .A2(KEYINPUT28), .ZN(n1387) );
XNOR2_X1 U1092 ( .A(G107), .B(n1389), .ZN(n1388) );
NOR2_X1 U1093 ( .A1(G104), .A2(KEYINPUT10), .ZN(n1389) );
NAND2_X1 U1094 ( .A1(n1390), .A2(n1391), .ZN(n1385) );
OR2_X1 U1095 ( .A1(n1392), .A2(n1199), .ZN(n1391) );
XOR2_X1 U1096 ( .A(G119), .B(n1393), .Z(n1199) );
NAND3_X1 U1097 ( .A1(n1393), .A2(n1336), .A3(n1392), .ZN(n1390) );
INV_X1 U1098 ( .A(KEYINPUT62), .ZN(n1392) );
INV_X1 U1099 ( .A(G119), .ZN(n1336) );
XNOR2_X1 U1100 ( .A(G110), .B(G122), .ZN(n1181) );
NOR2_X1 U1101 ( .A1(n1277), .A2(n1276), .ZN(n1088) );
XNOR2_X1 U1102 ( .A(n1110), .B(n1394), .ZN(n1276) );
NOR2_X1 U1103 ( .A1(KEYINPUT41), .A2(n1111), .ZN(n1394) );
INV_X1 U1104 ( .A(G475), .ZN(n1111) );
NAND2_X1 U1105 ( .A1(n1194), .A2(n1327), .ZN(n1110) );
INV_X1 U1106 ( .A(G902), .ZN(n1327) );
XNOR2_X1 U1107 ( .A(n1395), .B(n1396), .ZN(n1194) );
XOR2_X1 U1108 ( .A(n1397), .B(n1398), .Z(n1396) );
XOR2_X1 U1109 ( .A(G104), .B(n1399), .Z(n1398) );
NOR2_X1 U1110 ( .A1(KEYINPUT15), .A2(n1400), .ZN(n1399) );
XNOR2_X1 U1111 ( .A(n1289), .B(n1401), .ZN(n1400) );
XNOR2_X1 U1112 ( .A(n1370), .B(G140), .ZN(n1401) );
INV_X1 U1113 ( .A(G146), .ZN(n1370) );
INV_X1 U1114 ( .A(G125), .ZN(n1289) );
NOR2_X1 U1115 ( .A1(n1402), .A2(n1403), .ZN(n1397) );
XOR2_X1 U1116 ( .A(KEYINPUT42), .B(n1404), .Z(n1403) );
NOR2_X1 U1117 ( .A1(G131), .A2(n1405), .ZN(n1404) );
AND2_X1 U1118 ( .A1(n1405), .A2(G131), .ZN(n1402) );
NAND2_X1 U1119 ( .A1(n1406), .A2(n1407), .ZN(n1405) );
NAND2_X1 U1120 ( .A1(n1408), .A2(n1293), .ZN(n1407) );
XOR2_X1 U1121 ( .A(KEYINPUT5), .B(n1409), .Z(n1406) );
NOR2_X1 U1122 ( .A1(n1293), .A2(n1408), .ZN(n1409) );
NAND3_X1 U1123 ( .A1(n1333), .A2(n1081), .A3(G214), .ZN(n1408) );
INV_X1 U1124 ( .A(G237), .ZN(n1333) );
XNOR2_X1 U1125 ( .A(G113), .B(n1410), .ZN(n1395) );
XOR2_X1 U1126 ( .A(KEYINPUT63), .B(G122), .Z(n1410) );
NAND2_X1 U1127 ( .A1(n1411), .A2(n1412), .ZN(n1277) );
NAND2_X1 U1128 ( .A1(n1103), .A2(n1190), .ZN(n1412) );
XOR2_X1 U1129 ( .A(KEYINPUT56), .B(n1413), .Z(n1411) );
NOR2_X1 U1130 ( .A1(n1103), .A2(n1190), .ZN(n1413) );
INV_X1 U1131 ( .A(G478), .ZN(n1190) );
NOR2_X1 U1132 ( .A1(n1189), .A2(G902), .ZN(n1103) );
XNOR2_X1 U1133 ( .A(n1414), .B(n1415), .ZN(n1189) );
XOR2_X1 U1134 ( .A(G122), .B(n1416), .Z(n1415) );
XNOR2_X1 U1135 ( .A(n1293), .B(G134), .ZN(n1416) );
INV_X1 U1136 ( .A(G143), .ZN(n1293) );
XOR2_X1 U1137 ( .A(n1417), .B(n1330), .Z(n1414) );
XOR2_X1 U1138 ( .A(G128), .B(n1393), .Z(n1330) );
XOR2_X1 U1139 ( .A(G116), .B(KEYINPUT2), .Z(n1393) );
XOR2_X1 U1140 ( .A(n1418), .B(n1419), .Z(n1417) );
AND3_X1 U1141 ( .A1(G234), .A2(n1081), .A3(G217), .ZN(n1419) );
INV_X1 U1142 ( .A(G953), .ZN(n1081) );
NAND2_X1 U1143 ( .A1(KEYINPUT17), .A2(n1366), .ZN(n1418) );
INV_X1 U1144 ( .A(G107), .ZN(n1366) );
endmodule


