//Key = 1000000001100001101111010101110110010101110111010000111001110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371;

XNOR2_X1 U750 ( .A(G107), .B(n1032), .ZN(G9) );
NOR2_X1 U751 ( .A1(n1033), .A2(n1034), .ZN(G75) );
NOR2_X1 U752 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND4_X1 U753 ( .A1(KEYINPUT10), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1036) );
NAND4_X1 U754 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1035) );
NAND3_X1 U755 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1042) );
INV_X1 U756 ( .A(KEYINPUT54), .ZN(n1045) );
NAND4_X1 U757 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1044) );
NAND2_X1 U758 ( .A1(n1047), .A2(n1051), .ZN(n1041) );
NAND2_X1 U759 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND3_X1 U760 ( .A1(n1054), .A2(n1055), .A3(n1046), .ZN(n1053) );
NAND2_X1 U761 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
INV_X1 U762 ( .A(n1049), .ZN(n1057) );
NAND3_X1 U763 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1056) );
INV_X1 U764 ( .A(KEYINPUT37), .ZN(n1059) );
NAND3_X1 U765 ( .A1(n1061), .A2(n1062), .A3(n1049), .ZN(n1054) );
NAND2_X1 U766 ( .A1(n1050), .A2(n1063), .ZN(n1062) );
NAND2_X1 U767 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U768 ( .A1(KEYINPUT54), .A2(n1048), .ZN(n1065) );
NAND2_X1 U769 ( .A1(n1058), .A2(n1066), .ZN(n1061) );
NAND2_X1 U770 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U771 ( .A1(KEYINPUT37), .A2(n1060), .ZN(n1068) );
NAND3_X1 U772 ( .A1(n1050), .A2(n1069), .A3(n1058), .ZN(n1052) );
NAND3_X1 U773 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
NAND2_X1 U774 ( .A1(n1046), .A2(n1073), .ZN(n1072) );
NAND2_X1 U775 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U776 ( .A1(KEYINPUT9), .A2(n1076), .ZN(n1075) );
NAND2_X1 U777 ( .A1(n1077), .A2(n1078), .ZN(n1074) );
NAND3_X1 U778 ( .A1(n1079), .A2(n1080), .A3(n1049), .ZN(n1070) );
NAND2_X1 U779 ( .A1(n1081), .A2(n1082), .ZN(n1040) );
INV_X1 U780 ( .A(KEYINPUT9), .ZN(n1082) );
NAND4_X1 U781 ( .A1(n1047), .A2(n1046), .A3(n1083), .A4(n1058), .ZN(n1081) );
AND2_X1 U782 ( .A1(n1076), .A2(n1050), .ZN(n1083) );
INV_X1 U783 ( .A(n1084), .ZN(n1047) );
AND3_X1 U784 ( .A1(n1038), .A2(n1085), .A3(n1043), .ZN(n1033) );
NAND4_X1 U785 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1043) );
NOR4_X1 U786 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1089) );
XNOR2_X1 U787 ( .A(G475), .B(n1094), .ZN(n1093) );
XNOR2_X1 U788 ( .A(n1095), .B(n1096), .ZN(n1090) );
NOR3_X1 U789 ( .A1(n1077), .A2(n1080), .A3(n1097), .ZN(n1088) );
NAND2_X1 U790 ( .A1(n1098), .A2(G469), .ZN(n1087) );
XNOR2_X1 U791 ( .A(n1099), .B(KEYINPUT6), .ZN(n1098) );
XNOR2_X1 U792 ( .A(n1100), .B(n1101), .ZN(n1086) );
NAND2_X1 U793 ( .A1(KEYINPUT52), .A2(n1102), .ZN(n1101) );
XOR2_X1 U794 ( .A(n1103), .B(n1104), .Z(G72) );
NOR2_X1 U795 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NOR2_X1 U796 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
NAND2_X1 U797 ( .A1(n1109), .A2(n1110), .ZN(n1103) );
NAND2_X1 U798 ( .A1(n1111), .A2(n1106), .ZN(n1110) );
XNOR2_X1 U799 ( .A(n1039), .B(n1112), .ZN(n1111) );
NAND3_X1 U800 ( .A1(G900), .A2(n1112), .A3(G953), .ZN(n1109) );
XOR2_X1 U801 ( .A(n1113), .B(n1114), .Z(n1112) );
XNOR2_X1 U802 ( .A(n1115), .B(n1116), .ZN(n1114) );
XOR2_X1 U803 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U804 ( .A1(n1119), .A2(KEYINPUT0), .ZN(n1117) );
XOR2_X1 U805 ( .A(n1120), .B(G134), .Z(n1119) );
NAND2_X1 U806 ( .A1(KEYINPUT58), .A2(n1121), .ZN(n1120) );
XNOR2_X1 U807 ( .A(n1122), .B(n1123), .ZN(n1113) );
XNOR2_X1 U808 ( .A(KEYINPUT5), .B(KEYINPUT29), .ZN(n1122) );
XOR2_X1 U809 ( .A(n1124), .B(n1125), .Z(G69) );
NOR2_X1 U810 ( .A1(KEYINPUT33), .A2(n1126), .ZN(n1125) );
XOR2_X1 U811 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U812 ( .A1(n1037), .A2(G953), .ZN(n1128) );
NAND3_X1 U813 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1127) );
NAND2_X1 U814 ( .A1(G953), .A2(n1132), .ZN(n1131) );
NAND2_X1 U815 ( .A1(n1133), .A2(n1134), .ZN(n1130) );
NAND2_X1 U816 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U817 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XNOR2_X1 U818 ( .A(n1139), .B(KEYINPUT1), .ZN(n1135) );
NAND2_X1 U819 ( .A1(n1140), .A2(n1141), .ZN(n1129) );
NAND2_X1 U820 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
OR2_X1 U821 ( .A1(n1144), .A2(KEYINPUT1), .ZN(n1143) );
NAND2_X1 U822 ( .A1(n1139), .A2(KEYINPUT1), .ZN(n1142) );
NOR2_X1 U823 ( .A1(n1106), .A2(n1145), .ZN(n1124) );
XOR2_X1 U824 ( .A(KEYINPUT12), .B(n1146), .Z(n1145) );
NOR2_X1 U825 ( .A1(n1147), .A2(n1132), .ZN(n1146) );
NOR2_X1 U826 ( .A1(n1148), .A2(n1149), .ZN(G66) );
XOR2_X1 U827 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U828 ( .A1(n1102), .A2(n1152), .ZN(n1151) );
NOR2_X1 U829 ( .A1(n1153), .A2(n1154), .ZN(G63) );
XNOR2_X1 U830 ( .A(n1155), .B(n1156), .ZN(n1154) );
NOR2_X1 U831 ( .A1(n1157), .A2(n1152), .ZN(n1156) );
NOR2_X1 U832 ( .A1(n1106), .A2(n1158), .ZN(n1153) );
XNOR2_X1 U833 ( .A(KEYINPUT30), .B(n1085), .ZN(n1158) );
INV_X1 U834 ( .A(G952), .ZN(n1085) );
NOR2_X1 U835 ( .A1(n1148), .A2(n1159), .ZN(G60) );
XNOR2_X1 U836 ( .A(n1160), .B(n1161), .ZN(n1159) );
NOR3_X1 U837 ( .A1(n1152), .A2(KEYINPUT8), .A3(n1162), .ZN(n1161) );
XOR2_X1 U838 ( .A(G104), .B(n1163), .Z(G6) );
NOR2_X1 U839 ( .A1(n1148), .A2(n1164), .ZN(G57) );
NOR2_X1 U840 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XOR2_X1 U841 ( .A(KEYINPUT56), .B(n1167), .Z(n1166) );
AND2_X1 U842 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U843 ( .A1(n1169), .A2(n1168), .ZN(n1165) );
XOR2_X1 U844 ( .A(n1170), .B(n1171), .Z(n1168) );
NOR2_X1 U845 ( .A1(n1172), .A2(n1152), .ZN(n1171) );
NOR2_X1 U846 ( .A1(n1148), .A2(n1173), .ZN(G54) );
XOR2_X1 U847 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U848 ( .A1(n1176), .A2(n1152), .ZN(n1175) );
NOR2_X1 U849 ( .A1(n1177), .A2(n1178), .ZN(n1174) );
XOR2_X1 U850 ( .A(n1179), .B(KEYINPUT45), .Z(n1178) );
NAND2_X1 U851 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NOR2_X1 U852 ( .A1(n1181), .A2(n1180), .ZN(n1177) );
XNOR2_X1 U853 ( .A(n1182), .B(n1183), .ZN(n1180) );
XOR2_X1 U854 ( .A(n1184), .B(n1185), .Z(n1181) );
XOR2_X1 U855 ( .A(G140), .B(n1186), .Z(n1185) );
NAND2_X1 U856 ( .A1(KEYINPUT31), .A2(n1187), .ZN(n1184) );
NOR2_X1 U857 ( .A1(n1148), .A2(n1188), .ZN(G51) );
XOR2_X1 U858 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR3_X1 U859 ( .A1(n1152), .A2(KEYINPUT50), .A3(n1191), .ZN(n1190) );
NAND2_X1 U860 ( .A1(n1192), .A2(n1193), .ZN(n1152) );
NAND2_X1 U861 ( .A1(n1037), .A2(n1039), .ZN(n1193) );
AND4_X1 U862 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1039) );
NOR3_X1 U863 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1197) );
NOR2_X1 U864 ( .A1(KEYINPUT46), .A2(n1201), .ZN(n1200) );
NOR2_X1 U865 ( .A1(KEYINPUT38), .A2(n1202), .ZN(n1199) );
NAND4_X1 U866 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1198) );
NAND3_X1 U867 ( .A1(n1207), .A2(n1067), .A3(n1208), .ZN(n1206) );
INV_X1 U868 ( .A(KEYINPUT20), .ZN(n1208) );
NAND2_X1 U869 ( .A1(n1209), .A2(KEYINPUT20), .ZN(n1205) );
NAND2_X1 U870 ( .A1(n1210), .A2(n1211), .ZN(n1204) );
INV_X1 U871 ( .A(KEYINPUT22), .ZN(n1211) );
NAND3_X1 U872 ( .A1(n1046), .A2(n1212), .A3(KEYINPUT22), .ZN(n1203) );
AND3_X1 U873 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1196) );
NAND3_X1 U874 ( .A1(n1048), .A2(n1216), .A3(n1060), .ZN(n1194) );
NAND2_X1 U875 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NAND3_X1 U876 ( .A1(n1219), .A2(n1220), .A3(KEYINPUT38), .ZN(n1218) );
NAND3_X1 U877 ( .A1(n1221), .A2(n1222), .A3(KEYINPUT46), .ZN(n1217) );
AND4_X1 U878 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1037) );
NOR4_X1 U879 ( .A1(n1227), .A2(n1228), .A3(n1163), .A4(n1229), .ZN(n1226) );
NOR4_X1 U880 ( .A1(n1230), .A2(n1231), .A3(n1067), .A4(n1232), .ZN(n1229) );
XOR2_X1 U881 ( .A(KEYINPUT32), .B(n1233), .Z(n1232) );
INV_X1 U882 ( .A(n1234), .ZN(n1067) );
XNOR2_X1 U883 ( .A(n1076), .B(KEYINPUT51), .ZN(n1230) );
AND3_X1 U884 ( .A1(n1050), .A2(n1235), .A3(n1048), .ZN(n1163) );
AND2_X1 U885 ( .A1(n1032), .A2(n1236), .ZN(n1225) );
NAND3_X1 U886 ( .A1(n1237), .A2(n1235), .A3(n1050), .ZN(n1032) );
XNOR2_X1 U887 ( .A(G902), .B(KEYINPUT21), .ZN(n1192) );
NOR2_X1 U888 ( .A1(n1106), .A2(G952), .ZN(n1148) );
XNOR2_X1 U889 ( .A(G146), .B(n1195), .ZN(G48) );
NAND3_X1 U890 ( .A1(n1238), .A2(n1233), .A3(n1239), .ZN(n1195) );
XOR2_X1 U891 ( .A(n1209), .B(n1240), .Z(G45) );
NOR2_X1 U892 ( .A1(KEYINPUT26), .A2(n1241), .ZN(n1240) );
AND2_X1 U893 ( .A1(n1207), .A2(n1234), .ZN(n1209) );
AND4_X1 U894 ( .A1(n1242), .A2(n1219), .A3(n1243), .A4(n1233), .ZN(n1207) );
XNOR2_X1 U895 ( .A(G140), .B(n1202), .ZN(G42) );
NAND3_X1 U896 ( .A1(n1046), .A2(n1060), .A3(n1239), .ZN(n1202) );
XNOR2_X1 U897 ( .A(G137), .B(n1213), .ZN(G39) );
NAND4_X1 U898 ( .A1(n1046), .A2(n1219), .A3(n1238), .A4(n1058), .ZN(n1213) );
XNOR2_X1 U899 ( .A(G134), .B(n1215), .ZN(G36) );
NAND4_X1 U900 ( .A1(n1046), .A2(n1219), .A3(n1234), .A4(n1237), .ZN(n1215) );
INV_X1 U901 ( .A(n1220), .ZN(n1046) );
XOR2_X1 U902 ( .A(n1210), .B(n1244), .Z(G33) );
NOR2_X1 U903 ( .A1(KEYINPUT49), .A2(n1123), .ZN(n1244) );
NOR2_X1 U904 ( .A1(n1212), .A2(n1220), .ZN(n1210) );
NAND2_X1 U905 ( .A1(n1079), .A2(n1245), .ZN(n1220) );
INV_X1 U906 ( .A(n1092), .ZN(n1079) );
NAND2_X1 U907 ( .A1(n1239), .A2(n1234), .ZN(n1212) );
AND2_X1 U908 ( .A1(n1219), .A2(n1048), .ZN(n1239) );
XNOR2_X1 U909 ( .A(G128), .B(n1214), .ZN(G30) );
NAND4_X1 U910 ( .A1(n1219), .A2(n1238), .A3(n1237), .A4(n1233), .ZN(n1214) );
NOR2_X1 U911 ( .A1(n1246), .A2(n1221), .ZN(n1219) );
INV_X1 U912 ( .A(n1247), .ZN(n1221) );
INV_X1 U913 ( .A(n1076), .ZN(n1246) );
XNOR2_X1 U914 ( .A(G101), .B(n1248), .ZN(G3) );
NAND4_X1 U915 ( .A1(n1249), .A2(n1234), .A3(n1250), .A4(n1233), .ZN(n1248) );
XNOR2_X1 U916 ( .A(n1076), .B(KEYINPUT47), .ZN(n1249) );
XNOR2_X1 U917 ( .A(n1251), .B(n1201), .ZN(G27) );
NAND4_X1 U918 ( .A1(n1060), .A2(n1048), .A3(n1222), .A4(n1247), .ZN(n1201) );
NAND2_X1 U919 ( .A1(n1084), .A2(n1252), .ZN(n1247) );
NAND4_X1 U920 ( .A1(G902), .A2(G953), .A3(n1253), .A4(n1108), .ZN(n1252) );
INV_X1 U921 ( .A(G900), .ZN(n1108) );
XNOR2_X1 U922 ( .A(G125), .B(KEYINPUT25), .ZN(n1251) );
XOR2_X1 U923 ( .A(G122), .B(n1228), .Z(G24) );
AND4_X1 U924 ( .A1(n1243), .A2(n1254), .A3(n1050), .A4(n1255), .ZN(n1228) );
NOR2_X1 U925 ( .A1(n1071), .A2(n1256), .ZN(n1255) );
NOR2_X1 U926 ( .A1(n1091), .A2(n1257), .ZN(n1050) );
XNOR2_X1 U927 ( .A(n1258), .B(n1227), .ZN(G21) );
AND3_X1 U928 ( .A1(n1250), .A2(n1222), .A3(n1238), .ZN(n1227) );
AND2_X1 U929 ( .A1(n1257), .A2(n1091), .ZN(n1238) );
INV_X1 U930 ( .A(n1231), .ZN(n1250) );
NAND2_X1 U931 ( .A1(n1058), .A2(n1254), .ZN(n1231) );
XNOR2_X1 U932 ( .A(G116), .B(n1223), .ZN(G18) );
NAND2_X1 U933 ( .A1(n1259), .A2(n1237), .ZN(n1223) );
INV_X1 U934 ( .A(n1064), .ZN(n1237) );
NAND2_X1 U935 ( .A1(n1243), .A2(n1256), .ZN(n1064) );
XNOR2_X1 U936 ( .A(G113), .B(n1224), .ZN(G15) );
NAND2_X1 U937 ( .A1(n1259), .A2(n1048), .ZN(n1224) );
NOR2_X1 U938 ( .A1(n1256), .A2(n1243), .ZN(n1048) );
AND3_X1 U939 ( .A1(n1222), .A2(n1254), .A3(n1234), .ZN(n1259) );
NOR2_X1 U940 ( .A1(n1257), .A2(n1260), .ZN(n1234) );
INV_X1 U941 ( .A(n1071), .ZN(n1222) );
NAND2_X1 U942 ( .A1(n1049), .A2(n1233), .ZN(n1071) );
NOR2_X1 U943 ( .A1(n1261), .A2(n1077), .ZN(n1049) );
XNOR2_X1 U944 ( .A(G110), .B(n1236), .ZN(G12) );
NAND3_X1 U945 ( .A1(n1058), .A2(n1235), .A3(n1060), .ZN(n1236) );
AND2_X1 U946 ( .A1(n1260), .A2(n1257), .ZN(n1060) );
XNOR2_X1 U947 ( .A(n1102), .B(n1100), .ZN(n1257) );
NOR2_X1 U948 ( .A1(n1150), .A2(G902), .ZN(n1100) );
NAND2_X1 U949 ( .A1(n1262), .A2(n1263), .ZN(n1150) );
NAND2_X1 U950 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NAND2_X1 U951 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
INV_X1 U952 ( .A(KEYINPUT42), .ZN(n1267) );
OR2_X1 U953 ( .A1(n1268), .A2(KEYINPUT24), .ZN(n1266) );
NAND2_X1 U954 ( .A1(n1268), .A2(n1269), .ZN(n1262) );
NAND2_X1 U955 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
INV_X1 U956 ( .A(KEYINPUT24), .ZN(n1271) );
OR2_X1 U957 ( .A1(n1264), .A2(KEYINPUT42), .ZN(n1270) );
XNOR2_X1 U958 ( .A(n1272), .B(n1273), .ZN(n1264) );
NAND2_X1 U959 ( .A1(G221), .A2(n1274), .ZN(n1272) );
XNOR2_X1 U960 ( .A(n1275), .B(n1276), .ZN(n1268) );
XNOR2_X1 U961 ( .A(n1187), .B(n1277), .ZN(n1276) );
NOR2_X1 U962 ( .A1(KEYINPUT4), .A2(n1278), .ZN(n1277) );
XOR2_X1 U963 ( .A(n1279), .B(n1280), .Z(n1278) );
XNOR2_X1 U964 ( .A(n1281), .B(n1115), .ZN(n1280) );
NAND2_X1 U965 ( .A1(KEYINPUT16), .A2(n1282), .ZN(n1281) );
XOR2_X1 U966 ( .A(KEYINPUT62), .B(KEYINPUT48), .Z(n1279) );
INV_X1 U967 ( .A(G110), .ZN(n1187) );
XNOR2_X1 U968 ( .A(G119), .B(G128), .ZN(n1275) );
NAND2_X1 U969 ( .A1(G217), .A2(n1283), .ZN(n1102) );
INV_X1 U970 ( .A(n1091), .ZN(n1260) );
XOR2_X1 U971 ( .A(n1284), .B(n1172), .Z(n1091) );
INV_X1 U972 ( .A(G472), .ZN(n1172) );
NAND2_X1 U973 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
XNOR2_X1 U974 ( .A(n1287), .B(n1288), .ZN(n1285) );
INV_X1 U975 ( .A(n1170), .ZN(n1288) );
XNOR2_X1 U976 ( .A(n1289), .B(n1290), .ZN(n1170) );
XNOR2_X1 U977 ( .A(n1291), .B(n1292), .ZN(n1290) );
XOR2_X1 U978 ( .A(KEYINPUT23), .B(n1293), .Z(n1292) );
XOR2_X1 U979 ( .A(n1294), .B(n1295), .Z(n1289) );
NAND2_X1 U980 ( .A1(KEYINPUT35), .A2(n1169), .ZN(n1287) );
XOR2_X1 U981 ( .A(n1296), .B(G101), .Z(n1169) );
NAND3_X1 U982 ( .A1(n1297), .A2(n1106), .A3(G210), .ZN(n1296) );
XNOR2_X1 U983 ( .A(KEYINPUT15), .B(n1298), .ZN(n1297) );
AND3_X1 U984 ( .A1(n1233), .A2(n1254), .A3(n1076), .ZN(n1235) );
NOR2_X1 U985 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
INV_X1 U986 ( .A(n1261), .ZN(n1078) );
NAND3_X1 U987 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1261) );
INV_X1 U988 ( .A(n1097), .ZN(n1301) );
NOR2_X1 U989 ( .A1(n1302), .A2(G469), .ZN(n1097) );
NAND2_X1 U990 ( .A1(n1303), .A2(n1304), .ZN(n1300) );
INV_X1 U991 ( .A(KEYINPUT59), .ZN(n1304) );
NAND2_X1 U992 ( .A1(n1305), .A2(n1302), .ZN(n1303) );
XNOR2_X1 U993 ( .A(KEYINPUT17), .B(n1176), .ZN(n1305) );
NAND2_X1 U994 ( .A1(KEYINPUT59), .A2(n1306), .ZN(n1299) );
NAND2_X1 U995 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
OR3_X1 U996 ( .A1(n1176), .A2(n1099), .A3(KEYINPUT17), .ZN(n1308) );
INV_X1 U997 ( .A(n1302), .ZN(n1099) );
NAND2_X1 U998 ( .A1(n1309), .A2(n1286), .ZN(n1302) );
XOR2_X1 U999 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1000 ( .A(n1312), .B(n1183), .Z(n1311) );
XNOR2_X1 U1001 ( .A(n1313), .B(n1314), .ZN(n1183) );
XOR2_X1 U1002 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1003 ( .A(KEYINPUT14), .B(G104), .Z(n1316) );
NOR2_X1 U1004 ( .A1(KEYINPUT3), .A2(n1317), .ZN(n1315) );
INV_X1 U1005 ( .A(G101), .ZN(n1317) );
XOR2_X1 U1006 ( .A(n1318), .B(n1118), .Z(n1313) );
AND2_X1 U1007 ( .A1(n1319), .A2(n1320), .ZN(n1118) );
NAND3_X1 U1008 ( .A1(n1321), .A2(n1322), .A3(G128), .ZN(n1320) );
XOR2_X1 U1009 ( .A(KEYINPUT27), .B(n1323), .Z(n1319) );
NOR2_X1 U1010 ( .A1(G128), .A2(n1324), .ZN(n1323) );
AND2_X1 U1011 ( .A1(n1321), .A2(n1322), .ZN(n1324) );
NAND2_X1 U1012 ( .A1(n1325), .A2(n1326), .ZN(n1322) );
INV_X1 U1013 ( .A(KEYINPUT2), .ZN(n1326) );
XNOR2_X1 U1014 ( .A(G143), .B(G146), .ZN(n1325) );
NAND3_X1 U1015 ( .A1(G143), .A2(n1282), .A3(KEYINPUT2), .ZN(n1321) );
NAND2_X1 U1016 ( .A1(KEYINPUT43), .A2(n1327), .ZN(n1318) );
XOR2_X1 U1017 ( .A(KEYINPUT63), .B(G107), .Z(n1327) );
NOR2_X1 U1018 ( .A1(KEYINPUT13), .A2(n1291), .ZN(n1312) );
INV_X1 U1019 ( .A(n1182), .ZN(n1291) );
XOR2_X1 U1020 ( .A(n1328), .B(n1123), .Z(n1182) );
NAND2_X1 U1021 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
NAND2_X1 U1022 ( .A1(G134), .A2(n1273), .ZN(n1330) );
XOR2_X1 U1023 ( .A(KEYINPUT44), .B(n1331), .Z(n1329) );
NOR2_X1 U1024 ( .A1(G134), .A2(n1273), .ZN(n1331) );
INV_X1 U1025 ( .A(n1121), .ZN(n1273) );
XOR2_X1 U1026 ( .A(G137), .B(KEYINPUT7), .Z(n1121) );
NOR2_X1 U1027 ( .A1(n1332), .A2(n1333), .ZN(n1310) );
NOR2_X1 U1028 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
INV_X1 U1029 ( .A(n1336), .ZN(n1335) );
XOR2_X1 U1030 ( .A(KEYINPUT40), .B(n1186), .Z(n1334) );
NOR2_X1 U1031 ( .A1(n1336), .A2(n1337), .ZN(n1332) );
XOR2_X1 U1032 ( .A(KEYINPUT55), .B(n1186), .Z(n1337) );
NOR2_X1 U1033 ( .A1(n1107), .A2(G953), .ZN(n1186) );
INV_X1 U1034 ( .A(G227), .ZN(n1107) );
XOR2_X1 U1035 ( .A(G110), .B(G140), .Z(n1336) );
NAND2_X1 U1036 ( .A1(KEYINPUT17), .A2(n1176), .ZN(n1307) );
INV_X1 U1037 ( .A(G469), .ZN(n1176) );
AND2_X1 U1038 ( .A1(G221), .A2(n1283), .ZN(n1077) );
NAND2_X1 U1039 ( .A1(G234), .A2(n1286), .ZN(n1283) );
NAND2_X1 U1040 ( .A1(n1338), .A2(n1084), .ZN(n1254) );
NAND3_X1 U1041 ( .A1(n1038), .A2(n1253), .A3(G952), .ZN(n1084) );
XOR2_X1 U1042 ( .A(n1106), .B(KEYINPUT11), .Z(n1038) );
XOR2_X1 U1043 ( .A(KEYINPUT41), .B(n1339), .Z(n1338) );
AND4_X1 U1044 ( .A1(n1132), .A2(n1253), .A3(G953), .A4(G902), .ZN(n1339) );
NAND2_X1 U1045 ( .A1(G234), .A2(G237), .ZN(n1253) );
INV_X1 U1046 ( .A(G898), .ZN(n1132) );
AND2_X1 U1047 ( .A1(n1245), .A2(n1092), .ZN(n1233) );
XOR2_X1 U1048 ( .A(n1340), .B(n1191), .Z(n1092) );
NAND2_X1 U1049 ( .A1(G210), .A2(n1341), .ZN(n1191) );
NAND2_X1 U1050 ( .A1(n1342), .A2(n1286), .ZN(n1340) );
XOR2_X1 U1051 ( .A(n1189), .B(KEYINPUT19), .Z(n1342) );
XOR2_X1 U1052 ( .A(n1343), .B(n1344), .Z(n1189) );
XOR2_X1 U1053 ( .A(n1144), .B(n1345), .Z(n1344) );
XNOR2_X1 U1054 ( .A(G146), .B(n1346), .ZN(n1345) );
NOR2_X1 U1055 ( .A1(G953), .A2(n1147), .ZN(n1346) );
INV_X1 U1056 ( .A(G224), .ZN(n1147) );
OR2_X1 U1057 ( .A1(n1139), .A2(n1347), .ZN(n1144) );
AND2_X1 U1058 ( .A1(n1137), .A2(n1138), .ZN(n1347) );
NOR2_X1 U1059 ( .A1(n1138), .A2(n1137), .ZN(n1139) );
XOR2_X1 U1060 ( .A(G101), .B(n1348), .Z(n1137) );
XOR2_X1 U1061 ( .A(G107), .B(G104), .Z(n1348) );
XNOR2_X1 U1062 ( .A(n1349), .B(n1293), .ZN(n1138) );
XNOR2_X1 U1063 ( .A(n1258), .B(KEYINPUT60), .ZN(n1293) );
INV_X1 U1064 ( .A(G119), .ZN(n1258) );
XNOR2_X1 U1065 ( .A(G113), .B(G116), .ZN(n1349) );
XNOR2_X1 U1066 ( .A(n1350), .B(n1351), .ZN(n1343) );
XNOR2_X1 U1067 ( .A(n1141), .B(n1352), .ZN(n1351) );
INV_X1 U1068 ( .A(n1133), .ZN(n1141) );
XOR2_X1 U1069 ( .A(G110), .B(G122), .Z(n1133) );
XOR2_X1 U1070 ( .A(KEYINPUT28), .B(n1080), .Z(n1245) );
AND2_X1 U1071 ( .A1(G214), .A2(n1341), .ZN(n1080) );
NAND2_X1 U1072 ( .A1(n1298), .A2(n1286), .ZN(n1341) );
NOR2_X1 U1073 ( .A1(n1243), .A2(n1242), .ZN(n1058) );
INV_X1 U1074 ( .A(n1256), .ZN(n1242) );
XOR2_X1 U1075 ( .A(n1353), .B(n1094), .Z(n1256) );
NAND2_X1 U1076 ( .A1(n1160), .A2(n1286), .ZN(n1094) );
XNOR2_X1 U1077 ( .A(n1354), .B(n1355), .ZN(n1160) );
XOR2_X1 U1078 ( .A(G104), .B(n1356), .Z(n1355) );
XNOR2_X1 U1079 ( .A(n1123), .B(G122), .ZN(n1356) );
INV_X1 U1080 ( .A(G131), .ZN(n1123) );
XOR2_X1 U1081 ( .A(n1357), .B(n1358), .Z(n1354) );
NOR2_X1 U1082 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
NOR2_X1 U1083 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
XNOR2_X1 U1084 ( .A(KEYINPUT39), .B(n1241), .ZN(n1361) );
NOR2_X1 U1085 ( .A1(n1363), .A2(n1364), .ZN(n1359) );
XNOR2_X1 U1086 ( .A(KEYINPUT34), .B(n1241), .ZN(n1364) );
INV_X1 U1087 ( .A(n1362), .ZN(n1363) );
NAND3_X1 U1088 ( .A1(n1298), .A2(n1106), .A3(G214), .ZN(n1362) );
INV_X1 U1089 ( .A(G237), .ZN(n1298) );
XOR2_X1 U1090 ( .A(n1365), .B(n1295), .Z(n1357) );
XNOR2_X1 U1091 ( .A(G113), .B(n1282), .ZN(n1295) );
INV_X1 U1092 ( .A(G146), .ZN(n1282) );
NAND2_X1 U1093 ( .A1(KEYINPUT57), .A2(n1115), .ZN(n1365) );
XNOR2_X1 U1094 ( .A(G140), .B(n1366), .ZN(n1115) );
INV_X1 U1095 ( .A(n1350), .ZN(n1366) );
XOR2_X1 U1096 ( .A(G125), .B(KEYINPUT36), .Z(n1350) );
NAND2_X1 U1097 ( .A1(KEYINPUT53), .A2(n1162), .ZN(n1353) );
INV_X1 U1098 ( .A(G475), .ZN(n1162) );
XOR2_X1 U1099 ( .A(n1095), .B(n1367), .Z(n1243) );
NOR2_X1 U1100 ( .A1(KEYINPUT61), .A2(n1096), .ZN(n1367) );
XOR2_X1 U1101 ( .A(n1157), .B(KEYINPUT18), .Z(n1096) );
INV_X1 U1102 ( .A(G478), .ZN(n1157) );
NAND2_X1 U1103 ( .A1(n1155), .A2(n1286), .ZN(n1095) );
INV_X1 U1104 ( .A(G902), .ZN(n1286) );
XNOR2_X1 U1105 ( .A(n1368), .B(n1369), .ZN(n1155) );
XOR2_X1 U1106 ( .A(G107), .B(n1370), .Z(n1369) );
XOR2_X1 U1107 ( .A(G134), .B(G122), .Z(n1370) );
XOR2_X1 U1108 ( .A(n1294), .B(n1371), .Z(n1368) );
AND2_X1 U1109 ( .A1(G217), .A2(n1274), .ZN(n1371) );
AND2_X1 U1110 ( .A1(G234), .A2(n1106), .ZN(n1274) );
INV_X1 U1111 ( .A(G953), .ZN(n1106) );
XNOR2_X1 U1112 ( .A(G116), .B(n1352), .ZN(n1294) );
XNOR2_X1 U1113 ( .A(G128), .B(n1241), .ZN(n1352) );
INV_X1 U1114 ( .A(G143), .ZN(n1241) );
endmodule


