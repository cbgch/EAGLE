//Key = 1010100010011101110000010011010100110010001100101000101100011101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;

XNOR2_X1 U733 ( .A(G107), .B(n1010), .ZN(G9) );
NOR2_X1 U734 ( .A1(n1011), .A2(n1012), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
INV_X1 U736 ( .A(G952), .ZN(n1016) );
NOR2_X1 U737 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NOR3_X1 U738 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1017) );
NOR2_X1 U739 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NOR2_X1 U740 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR3_X1 U741 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NOR3_X1 U742 ( .A1(n1029), .A2(KEYINPUT7), .A3(n1030), .ZN(n1024) );
NOR3_X1 U743 ( .A1(n1029), .A2(n1031), .A3(n1028), .ZN(n1020) );
NOR2_X1 U744 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U745 ( .A1(n1034), .A2(n1035), .ZN(n1019) );
INV_X1 U746 ( .A(KEYINPUT7), .ZN(n1035) );
NOR3_X1 U747 ( .A1(n1029), .A2(n1030), .A3(n1023), .ZN(n1034) );
INV_X1 U748 ( .A(n1036), .ZN(n1030) );
INV_X1 U749 ( .A(n1037), .ZN(n1029) );
NAND3_X1 U750 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1013) );
NAND3_X1 U751 ( .A1(n1041), .A2(n1042), .A3(n1037), .ZN(n1040) );
NOR3_X1 U752 ( .A1(n1043), .A2(n1044), .A3(n1026), .ZN(n1037) );
NAND2_X1 U753 ( .A1(n1045), .A2(n1046), .ZN(n1042) );
NAND3_X1 U754 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
XOR2_X1 U755 ( .A(n1018), .B(KEYINPUT13), .Z(n1049) );
NAND2_X1 U756 ( .A1(n1050), .A2(n1051), .ZN(n1045) );
NAND2_X1 U757 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U758 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR3_X1 U759 ( .A1(n1056), .A2(G953), .A3(n1057), .ZN(n1011) );
INV_X1 U760 ( .A(n1038), .ZN(n1057) );
NAND4_X1 U761 ( .A1(n1047), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1038) );
XOR2_X1 U762 ( .A(KEYINPUT51), .B(n1061), .Z(n1059) );
NOR4_X1 U763 ( .A1(n1043), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1061) );
XOR2_X1 U764 ( .A(G478), .B(n1065), .Z(n1064) );
XNOR2_X1 U765 ( .A(n1066), .B(n1067), .ZN(n1063) );
XOR2_X1 U766 ( .A(KEYINPUT22), .B(G952), .Z(n1056) );
XOR2_X1 U767 ( .A(n1068), .B(n1069), .Z(G72) );
XOR2_X1 U768 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U770 ( .A(n1074), .B(n1075), .Z(n1073) );
XOR2_X1 U771 ( .A(n1076), .B(n1077), .Z(n1075) );
XOR2_X1 U772 ( .A(n1078), .B(n1079), .Z(n1074) );
XNOR2_X1 U773 ( .A(KEYINPUT59), .B(KEYINPUT38), .ZN(n1079) );
NAND2_X1 U774 ( .A1(KEYINPUT35), .A2(n1080), .ZN(n1078) );
XNOR2_X1 U775 ( .A(n1081), .B(n1082), .ZN(n1080) );
XNOR2_X1 U776 ( .A(KEYINPUT8), .B(KEYINPUT21), .ZN(n1082) );
XOR2_X1 U777 ( .A(n1083), .B(KEYINPUT41), .Z(n1072) );
NAND2_X1 U778 ( .A1(n1084), .A2(G953), .ZN(n1083) );
XOR2_X1 U779 ( .A(n1085), .B(KEYINPUT3), .Z(n1084) );
NAND2_X1 U780 ( .A1(KEYINPUT42), .A2(n1086), .ZN(n1070) );
NAND2_X1 U781 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U782 ( .A(n1039), .B(KEYINPUT30), .Z(n1087) );
NAND2_X1 U783 ( .A1(G953), .A2(n1089), .ZN(n1068) );
NAND2_X1 U784 ( .A1(G900), .A2(G227), .ZN(n1089) );
XOR2_X1 U785 ( .A(n1090), .B(n1091), .Z(G69) );
NOR2_X1 U786 ( .A1(n1092), .A2(n1039), .ZN(n1091) );
NOR2_X1 U787 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U788 ( .A(n1095), .B(KEYINPUT56), .Z(n1093) );
NAND2_X1 U789 ( .A1(n1096), .A2(n1097), .ZN(n1090) );
NAND2_X1 U790 ( .A1(n1098), .A2(n1039), .ZN(n1097) );
XNOR2_X1 U791 ( .A(n1099), .B(n1100), .ZN(n1098) );
OR3_X1 U792 ( .A1(n1095), .A2(n1100), .A3(n1039), .ZN(n1096) );
XOR2_X1 U793 ( .A(n1101), .B(n1102), .Z(n1100) );
XOR2_X1 U794 ( .A(n1103), .B(n1104), .Z(n1101) );
NOR2_X1 U795 ( .A1(n1105), .A2(n1106), .ZN(G66) );
XOR2_X1 U796 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND2_X1 U797 ( .A1(n1109), .A2(n1067), .ZN(n1107) );
NOR2_X1 U798 ( .A1(n1105), .A2(n1110), .ZN(G63) );
NOR3_X1 U799 ( .A1(n1111), .A2(n1065), .A3(n1112), .ZN(n1110) );
NOR2_X1 U800 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U801 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
XOR2_X1 U802 ( .A(n1117), .B(KEYINPUT31), .Z(n1111) );
NAND3_X1 U803 ( .A1(G478), .A2(n1114), .A3(n1109), .ZN(n1117) );
NOR2_X1 U804 ( .A1(n1105), .A2(n1118), .ZN(G60) );
XNOR2_X1 U805 ( .A(n1119), .B(n1120), .ZN(n1118) );
AND2_X1 U806 ( .A1(G475), .A2(n1109), .ZN(n1120) );
XNOR2_X1 U807 ( .A(G104), .B(n1121), .ZN(G6) );
NOR2_X1 U808 ( .A1(n1105), .A2(n1122), .ZN(G57) );
NOR3_X1 U809 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1122) );
NOR2_X1 U810 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NOR2_X1 U811 ( .A1(KEYINPUT62), .A2(n1128), .ZN(n1127) );
XOR2_X1 U812 ( .A(KEYINPUT33), .B(n1129), .Z(n1128) );
INV_X1 U813 ( .A(n1130), .ZN(n1126) );
NOR3_X1 U814 ( .A1(n1130), .A2(KEYINPUT62), .A3(n1129), .ZN(n1124) );
NAND2_X1 U815 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U816 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U817 ( .A1(n1109), .A2(G472), .ZN(n1134) );
XOR2_X1 U818 ( .A(KEYINPUT43), .B(n1135), .Z(n1131) );
NOR3_X1 U819 ( .A1(n1136), .A2(n1133), .A3(n1137), .ZN(n1135) );
INV_X1 U820 ( .A(G472), .ZN(n1137) );
AND2_X1 U821 ( .A1(n1138), .A2(n1139), .ZN(n1133) );
NAND2_X1 U822 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U823 ( .A1(n1142), .A2(n1143), .ZN(n1138) );
XOR2_X1 U824 ( .A(n1141), .B(KEYINPUT2), .Z(n1142) );
XNOR2_X1 U825 ( .A(n1081), .B(n1144), .ZN(n1141) );
AND2_X1 U826 ( .A1(n1129), .A2(KEYINPUT62), .ZN(n1123) );
NOR2_X1 U827 ( .A1(n1105), .A2(n1145), .ZN(G54) );
NOR2_X1 U828 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U829 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U830 ( .A1(KEYINPUT46), .A2(n1150), .ZN(n1149) );
NAND2_X1 U831 ( .A1(n1109), .A2(G469), .ZN(n1148) );
INV_X1 U832 ( .A(n1136), .ZN(n1109) );
NOR2_X1 U833 ( .A1(KEYINPUT46), .A2(n1150), .ZN(n1146) );
XOR2_X1 U834 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U835 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U836 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U837 ( .A1(n1157), .A2(n1158), .ZN(n1153) );
XOR2_X1 U838 ( .A(n1155), .B(KEYINPUT63), .Z(n1158) );
INV_X1 U839 ( .A(n1156), .ZN(n1157) );
XNOR2_X1 U840 ( .A(n1159), .B(KEYINPUT24), .ZN(n1156) );
XOR2_X1 U841 ( .A(n1160), .B(KEYINPUT55), .Z(n1151) );
NOR2_X1 U842 ( .A1(n1105), .A2(n1161), .ZN(G51) );
XNOR2_X1 U843 ( .A(n1162), .B(n1163), .ZN(n1161) );
XOR2_X1 U844 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U845 ( .A1(KEYINPUT45), .A2(n1166), .ZN(n1165) );
NOR2_X1 U846 ( .A1(n1167), .A2(n1136), .ZN(n1164) );
NAND2_X1 U847 ( .A1(G902), .A2(n1014), .ZN(n1136) );
INV_X1 U848 ( .A(n1115), .ZN(n1014) );
NOR2_X1 U849 ( .A1(n1099), .A2(n1088), .ZN(n1115) );
NAND4_X1 U850 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1088) );
NOR4_X1 U851 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1171) );
NOR2_X1 U852 ( .A1(n1176), .A2(n1177), .ZN(n1170) );
NOR2_X1 U853 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
INV_X1 U854 ( .A(KEYINPUT4), .ZN(n1179) );
NAND2_X1 U855 ( .A1(n1180), .A2(n1181), .ZN(n1169) );
NAND3_X1 U856 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1181) );
OR2_X1 U857 ( .A1(n1185), .A2(KEYINPUT20), .ZN(n1184) );
NAND4_X1 U858 ( .A1(n1186), .A2(n1033), .A3(n1187), .A4(n1188), .ZN(n1182) );
NOR2_X1 U859 ( .A1(KEYINPUT4), .A2(n1050), .ZN(n1187) );
NAND3_X1 U860 ( .A1(KEYINPUT20), .A2(n1189), .A3(n1052), .ZN(n1168) );
INV_X1 U861 ( .A(n1185), .ZN(n1189) );
NAND4_X1 U862 ( .A1(n1190), .A2(n1121), .A3(n1191), .A4(n1192), .ZN(n1099) );
AND4_X1 U863 ( .A1(n1010), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1192) );
NAND3_X1 U864 ( .A1(n1032), .A2(n1196), .A3(n1036), .ZN(n1010) );
NAND2_X1 U865 ( .A1(n1197), .A2(n1180), .ZN(n1191) );
NAND3_X1 U866 ( .A1(n1036), .A2(n1196), .A3(n1033), .ZN(n1121) );
OR2_X1 U867 ( .A1(n1198), .A2(n1027), .ZN(n1190) );
NOR2_X1 U868 ( .A1(n1186), .A2(n1199), .ZN(n1027) );
NOR2_X1 U869 ( .A1(n1039), .A2(G952), .ZN(n1105) );
XNOR2_X1 U870 ( .A(n1175), .B(n1200), .ZN(G48) );
NAND2_X1 U871 ( .A1(G146), .A2(n1201), .ZN(n1200) );
XOR2_X1 U872 ( .A(KEYINPUT58), .B(KEYINPUT0), .Z(n1201) );
AND3_X1 U873 ( .A1(n1202), .A2(n1036), .A3(n1203), .ZN(n1175) );
NAND2_X1 U874 ( .A1(n1204), .A2(n1205), .ZN(G45) );
OR2_X1 U875 ( .A1(G143), .A2(KEYINPUT27), .ZN(n1205) );
XOR2_X1 U876 ( .A(n1206), .B(n1207), .Z(n1204) );
NOR2_X1 U877 ( .A1(n1052), .A2(n1185), .ZN(n1207) );
NAND4_X1 U878 ( .A1(n1208), .A2(n1199), .A3(n1209), .A4(n1036), .ZN(n1185) );
AND2_X1 U879 ( .A1(n1188), .A2(n1210), .ZN(n1209) );
NAND2_X1 U880 ( .A1(KEYINPUT27), .A2(G143), .ZN(n1206) );
NAND2_X1 U881 ( .A1(n1211), .A2(n1212), .ZN(G42) );
NAND2_X1 U882 ( .A1(G140), .A2(n1213), .ZN(n1212) );
XOR2_X1 U883 ( .A(n1214), .B(KEYINPUT28), .Z(n1211) );
NAND2_X1 U884 ( .A1(n1176), .A2(n1215), .ZN(n1214) );
INV_X1 U885 ( .A(n1213), .ZN(n1176) );
NAND3_X1 U886 ( .A1(n1216), .A2(n1033), .A3(n1186), .ZN(n1213) );
XOR2_X1 U887 ( .A(G137), .B(n1174), .Z(G39) );
AND3_X1 U888 ( .A1(n1202), .A2(n1041), .A3(n1216), .ZN(n1174) );
XOR2_X1 U889 ( .A(G134), .B(n1173), .Z(G36) );
AND3_X1 U890 ( .A1(n1199), .A2(n1032), .A3(n1216), .ZN(n1173) );
XOR2_X1 U891 ( .A(G131), .B(n1172), .Z(G33) );
AND3_X1 U892 ( .A1(n1033), .A2(n1199), .A3(n1216), .ZN(n1172) );
AND3_X1 U893 ( .A1(n1036), .A2(n1188), .A3(n1058), .ZN(n1216) );
INV_X1 U894 ( .A(n1018), .ZN(n1058) );
NAND2_X1 U895 ( .A1(n1055), .A2(n1217), .ZN(n1018) );
INV_X1 U896 ( .A(n1218), .ZN(n1199) );
XNOR2_X1 U897 ( .A(G128), .B(n1219), .ZN(G30) );
NAND2_X1 U898 ( .A1(n1220), .A2(n1180), .ZN(n1219) );
XOR2_X1 U899 ( .A(n1183), .B(KEYINPUT61), .Z(n1220) );
NAND4_X1 U900 ( .A1(n1202), .A2(n1036), .A3(n1032), .A4(n1188), .ZN(n1183) );
XOR2_X1 U901 ( .A(n1221), .B(n1222), .Z(G3) );
NOR2_X1 U902 ( .A1(KEYINPUT19), .A2(n1223), .ZN(n1222) );
NOR2_X1 U903 ( .A1(n1218), .A2(n1198), .ZN(n1221) );
XNOR2_X1 U904 ( .A(G125), .B(n1178), .ZN(G27) );
NAND3_X1 U905 ( .A1(n1203), .A2(n1050), .A3(n1186), .ZN(n1178) );
AND3_X1 U906 ( .A1(n1180), .A2(n1188), .A3(n1033), .ZN(n1203) );
NAND2_X1 U907 ( .A1(n1026), .A2(n1224), .ZN(n1188) );
NAND4_X1 U908 ( .A1(G953), .A2(G902), .A3(n1225), .A4(n1085), .ZN(n1224) );
INV_X1 U909 ( .A(G900), .ZN(n1085) );
NAND2_X1 U910 ( .A1(n1226), .A2(n1227), .ZN(G24) );
OR2_X1 U911 ( .A1(n1195), .A2(G122), .ZN(n1227) );
XOR2_X1 U912 ( .A(n1228), .B(KEYINPUT9), .Z(n1226) );
NAND2_X1 U913 ( .A1(G122), .A2(n1195), .ZN(n1228) );
NAND4_X1 U914 ( .A1(n1208), .A2(n1050), .A3(n1210), .A4(n1196), .ZN(n1195) );
NOR4_X1 U915 ( .A1(n1052), .A2(n1044), .A3(n1043), .A4(n1229), .ZN(n1196) );
XNOR2_X1 U916 ( .A(G119), .B(n1194), .ZN(G21) );
NAND3_X1 U917 ( .A1(n1202), .A2(n1050), .A3(n1230), .ZN(n1194) );
INV_X1 U918 ( .A(n1028), .ZN(n1050) );
NOR2_X1 U919 ( .A1(n1231), .A2(n1232), .ZN(n1202) );
INV_X1 U920 ( .A(n1043), .ZN(n1232) );
XNOR2_X1 U921 ( .A(G116), .B(n1233), .ZN(G18) );
NAND2_X1 U922 ( .A1(n1180), .A2(n1234), .ZN(n1233) );
XOR2_X1 U923 ( .A(KEYINPUT40), .B(n1197), .Z(n1234) );
AND2_X1 U924 ( .A1(n1235), .A2(n1032), .ZN(n1197) );
AND2_X1 U925 ( .A1(n1210), .A2(n1236), .ZN(n1032) );
XNOR2_X1 U926 ( .A(G113), .B(n1193), .ZN(G15) );
NAND3_X1 U927 ( .A1(n1235), .A2(n1180), .A3(n1033), .ZN(n1193) );
NOR2_X1 U928 ( .A1(n1236), .A2(n1210), .ZN(n1033) );
INV_X1 U929 ( .A(n1208), .ZN(n1236) );
NOR3_X1 U930 ( .A1(n1218), .A2(n1229), .A3(n1028), .ZN(n1235) );
NAND2_X1 U931 ( .A1(n1237), .A2(n1047), .ZN(n1028) );
XOR2_X1 U932 ( .A(KEYINPUT5), .B(n1060), .Z(n1237) );
NAND2_X1 U933 ( .A1(n1238), .A2(n1043), .ZN(n1218) );
XNOR2_X1 U934 ( .A(KEYINPUT57), .B(n1044), .ZN(n1238) );
XOR2_X1 U935 ( .A(G110), .B(n1239), .Z(G12) );
NOR2_X1 U936 ( .A1(n1198), .A2(n1240), .ZN(n1239) );
XOR2_X1 U937 ( .A(KEYINPUT12), .B(n1186), .Z(n1240) );
NOR2_X1 U938 ( .A1(n1043), .A2(n1231), .ZN(n1186) );
XOR2_X1 U939 ( .A(n1044), .B(KEYINPUT26), .Z(n1231) );
NAND3_X1 U940 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1044) );
OR2_X1 U941 ( .A1(n1066), .A2(n1067), .ZN(n1243) );
NAND2_X1 U942 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
INV_X1 U943 ( .A(KEYINPUT17), .ZN(n1245) );
NAND2_X1 U944 ( .A1(n1246), .A2(n1066), .ZN(n1244) );
XNOR2_X1 U945 ( .A(n1067), .B(KEYINPUT15), .ZN(n1246) );
NAND2_X1 U946 ( .A1(KEYINPUT17), .A2(n1247), .ZN(n1241) );
NAND2_X1 U947 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
OR2_X1 U948 ( .A1(n1067), .A2(KEYINPUT15), .ZN(n1249) );
NAND3_X1 U949 ( .A1(n1067), .A2(n1066), .A3(KEYINPUT15), .ZN(n1248) );
NAND2_X1 U950 ( .A1(n1108), .A2(n1250), .ZN(n1066) );
XOR2_X1 U951 ( .A(n1251), .B(n1252), .Z(n1108) );
XOR2_X1 U952 ( .A(n1253), .B(n1254), .Z(n1252) );
NOR2_X1 U953 ( .A1(n1255), .A2(n1256), .ZN(n1253) );
INV_X1 U954 ( .A(G221), .ZN(n1255) );
XOR2_X1 U955 ( .A(n1257), .B(n1258), .Z(n1251) );
NOR2_X1 U956 ( .A1(KEYINPUT14), .A2(n1259), .ZN(n1258) );
XOR2_X1 U957 ( .A(n1260), .B(n1261), .Z(n1259) );
NOR2_X1 U958 ( .A1(KEYINPUT49), .A2(G110), .ZN(n1261) );
XNOR2_X1 U959 ( .A(G119), .B(G128), .ZN(n1260) );
XNOR2_X1 U960 ( .A(G137), .B(KEYINPUT37), .ZN(n1257) );
AND2_X1 U961 ( .A1(G217), .A2(n1262), .ZN(n1067) );
XNOR2_X1 U962 ( .A(n1263), .B(n1264), .ZN(n1043) );
XOR2_X1 U963 ( .A(KEYINPUT32), .B(G472), .Z(n1264) );
NAND2_X1 U964 ( .A1(n1265), .A2(n1250), .ZN(n1263) );
XOR2_X1 U965 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U966 ( .A(n1140), .B(n1144), .Z(n1267) );
INV_X1 U967 ( .A(n1143), .ZN(n1140) );
XOR2_X1 U968 ( .A(n1268), .B(G113), .Z(n1143) );
NAND2_X1 U969 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
OR2_X1 U970 ( .A1(n1271), .A2(G119), .ZN(n1270) );
XOR2_X1 U971 ( .A(n1272), .B(KEYINPUT50), .Z(n1269) );
NAND2_X1 U972 ( .A1(G119), .A2(n1271), .ZN(n1272) );
XOR2_X1 U973 ( .A(G116), .B(KEYINPUT60), .Z(n1271) );
XNOR2_X1 U974 ( .A(n1129), .B(n1273), .ZN(n1266) );
XNOR2_X1 U975 ( .A(n1274), .B(KEYINPUT11), .ZN(n1273) );
NAND2_X1 U976 ( .A1(KEYINPUT52), .A2(n1081), .ZN(n1274) );
XNOR2_X1 U977 ( .A(n1275), .B(G101), .ZN(n1129) );
NAND2_X1 U978 ( .A1(G210), .A2(n1276), .ZN(n1275) );
NAND2_X1 U979 ( .A1(n1230), .A2(n1036), .ZN(n1198) );
NOR2_X1 U980 ( .A1(n1277), .A2(n1047), .ZN(n1036) );
XOR2_X1 U981 ( .A(n1278), .B(G469), .Z(n1047) );
NAND2_X1 U982 ( .A1(n1279), .A2(n1250), .ZN(n1278) );
XOR2_X1 U983 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U984 ( .A(n1282), .B(n1159), .Z(n1281) );
XOR2_X1 U985 ( .A(n1283), .B(n1215), .Z(n1159) );
INV_X1 U986 ( .A(G140), .ZN(n1215) );
INV_X1 U987 ( .A(G110), .ZN(n1283) );
INV_X1 U988 ( .A(n1160), .ZN(n1282) );
XOR2_X1 U989 ( .A(n1284), .B(n1285), .Z(n1160) );
XNOR2_X1 U990 ( .A(n1286), .B(n1077), .ZN(n1285) );
XNOR2_X1 U991 ( .A(n1287), .B(n1288), .ZN(n1077) );
XOR2_X1 U992 ( .A(n1289), .B(KEYINPUT44), .Z(n1287) );
XNOR2_X1 U993 ( .A(n1081), .B(n1290), .ZN(n1284) );
XOR2_X1 U994 ( .A(KEYINPUT39), .B(G101), .Z(n1290) );
XNOR2_X1 U995 ( .A(n1291), .B(n1292), .ZN(n1081) );
XOR2_X1 U996 ( .A(KEYINPUT47), .B(G137), .Z(n1292) );
XNOR2_X1 U997 ( .A(G131), .B(n1293), .ZN(n1291) );
XOR2_X1 U998 ( .A(KEYINPUT18), .B(n1294), .Z(n1280) );
NOR2_X1 U999 ( .A1(KEYINPUT36), .A2(n1155), .ZN(n1294) );
NAND2_X1 U1000 ( .A1(G227), .A2(n1039), .ZN(n1155) );
XOR2_X1 U1001 ( .A(KEYINPUT5), .B(n1048), .Z(n1277) );
INV_X1 U1002 ( .A(n1060), .ZN(n1048) );
NAND2_X1 U1003 ( .A1(G221), .A2(n1262), .ZN(n1060) );
NAND2_X1 U1004 ( .A1(G234), .A2(n1250), .ZN(n1262) );
NOR3_X1 U1005 ( .A1(n1052), .A2(n1229), .A3(n1023), .ZN(n1230) );
INV_X1 U1006 ( .A(n1041), .ZN(n1023) );
NOR2_X1 U1007 ( .A1(n1208), .A2(n1210), .ZN(n1041) );
XOR2_X1 U1008 ( .A(n1295), .B(n1065), .Z(n1210) );
NOR2_X1 U1009 ( .A1(n1114), .A2(G902), .ZN(n1065) );
XNOR2_X1 U1010 ( .A(n1296), .B(n1297), .ZN(n1114) );
XOR2_X1 U1011 ( .A(n1298), .B(n1299), .Z(n1297) );
NOR2_X1 U1012 ( .A1(n1256), .A2(n1300), .ZN(n1299) );
INV_X1 U1013 ( .A(G217), .ZN(n1300) );
NAND2_X1 U1014 ( .A1(G234), .A2(n1039), .ZN(n1256) );
NOR2_X1 U1015 ( .A1(G116), .A2(KEYINPUT25), .ZN(n1298) );
XOR2_X1 U1016 ( .A(n1301), .B(n1302), .Z(n1296) );
NOR2_X1 U1017 ( .A1(KEYINPUT10), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1018 ( .A(n1304), .B(n1293), .Z(n1303) );
XOR2_X1 U1019 ( .A(G134), .B(KEYINPUT53), .Z(n1293) );
XOR2_X1 U1020 ( .A(G128), .B(n1289), .Z(n1304) );
XNOR2_X1 U1021 ( .A(G107), .B(G122), .ZN(n1301) );
NAND2_X1 U1022 ( .A1(KEYINPUT16), .A2(n1116), .ZN(n1295) );
INV_X1 U1023 ( .A(G478), .ZN(n1116) );
XNOR2_X1 U1024 ( .A(n1062), .B(KEYINPUT34), .ZN(n1208) );
XNOR2_X1 U1025 ( .A(n1305), .B(G475), .ZN(n1062) );
NAND2_X1 U1026 ( .A1(n1119), .A2(n1250), .ZN(n1305) );
XNOR2_X1 U1027 ( .A(n1306), .B(n1307), .ZN(n1119) );
XOR2_X1 U1028 ( .A(G104), .B(n1308), .Z(n1307) );
XOR2_X1 U1029 ( .A(G122), .B(G113), .Z(n1308) );
XOR2_X1 U1030 ( .A(n1309), .B(n1254), .Z(n1306) );
XOR2_X1 U1031 ( .A(G146), .B(n1076), .Z(n1254) );
XOR2_X1 U1032 ( .A(G125), .B(G140), .Z(n1076) );
NAND2_X1 U1033 ( .A1(KEYINPUT29), .A2(n1310), .ZN(n1309) );
XOR2_X1 U1034 ( .A(n1311), .B(n1312), .Z(n1310) );
XOR2_X1 U1035 ( .A(G131), .B(n1289), .Z(n1312) );
NAND2_X1 U1036 ( .A1(G214), .A2(n1276), .ZN(n1311) );
NOR2_X1 U1037 ( .A1(G953), .A2(G237), .ZN(n1276) );
AND2_X1 U1038 ( .A1(n1026), .A2(n1313), .ZN(n1229) );
NAND4_X1 U1039 ( .A1(G953), .A2(G902), .A3(n1225), .A4(n1095), .ZN(n1313) );
INV_X1 U1040 ( .A(G898), .ZN(n1095) );
NAND3_X1 U1041 ( .A1(n1225), .A2(n1039), .A3(G952), .ZN(n1026) );
INV_X1 U1042 ( .A(G953), .ZN(n1039) );
NAND2_X1 U1043 ( .A1(G237), .A2(G234), .ZN(n1225) );
INV_X1 U1044 ( .A(n1180), .ZN(n1052) );
NOR2_X1 U1045 ( .A1(n1055), .A2(n1054), .ZN(n1180) );
INV_X1 U1046 ( .A(n1217), .ZN(n1054) );
NAND2_X1 U1047 ( .A1(G214), .A2(n1314), .ZN(n1217) );
XNOR2_X1 U1048 ( .A(n1315), .B(n1167), .ZN(n1055) );
NAND2_X1 U1049 ( .A1(G210), .A2(n1314), .ZN(n1167) );
NAND2_X1 U1050 ( .A1(n1316), .A2(n1250), .ZN(n1314) );
INV_X1 U1051 ( .A(G237), .ZN(n1316) );
NAND2_X1 U1052 ( .A1(n1317), .A2(n1250), .ZN(n1315) );
INV_X1 U1053 ( .A(G902), .ZN(n1250) );
XNOR2_X1 U1054 ( .A(n1166), .B(n1162), .ZN(n1317) );
XNOR2_X1 U1055 ( .A(n1318), .B(n1319), .ZN(n1162) );
XNOR2_X1 U1056 ( .A(n1103), .B(n1320), .ZN(n1319) );
NOR2_X1 U1057 ( .A1(KEYINPUT1), .A2(n1104), .ZN(n1320) );
XOR2_X1 U1058 ( .A(G110), .B(G122), .Z(n1104) );
NAND2_X1 U1059 ( .A1(n1321), .A2(n1322), .ZN(n1103) );
NAND2_X1 U1060 ( .A1(n1286), .A2(n1223), .ZN(n1322) );
XOR2_X1 U1061 ( .A(KEYINPUT54), .B(n1323), .Z(n1321) );
NOR2_X1 U1062 ( .A1(n1286), .A2(n1223), .ZN(n1323) );
INV_X1 U1063 ( .A(G101), .ZN(n1223) );
XNOR2_X1 U1064 ( .A(G104), .B(G107), .ZN(n1286) );
NAND2_X1 U1065 ( .A1(KEYINPUT23), .A2(n1102), .ZN(n1318) );
XNOR2_X1 U1066 ( .A(G113), .B(n1324), .ZN(n1102) );
NOR2_X1 U1067 ( .A1(KEYINPUT6), .A2(n1325), .ZN(n1324) );
XNOR2_X1 U1068 ( .A(G116), .B(G119), .ZN(n1325) );
XOR2_X1 U1069 ( .A(n1144), .B(n1326), .Z(n1166) );
XOR2_X1 U1070 ( .A(G125), .B(n1327), .Z(n1326) );
NOR2_X1 U1071 ( .A1(G953), .A2(n1094), .ZN(n1327) );
INV_X1 U1072 ( .A(G224), .ZN(n1094) );
XNOR2_X1 U1073 ( .A(n1328), .B(n1288), .ZN(n1144) );
XOR2_X1 U1074 ( .A(G146), .B(G128), .Z(n1288) );
NAND2_X1 U1075 ( .A1(KEYINPUT48), .A2(n1289), .ZN(n1328) );
INV_X1 U1076 ( .A(G143), .ZN(n1289) );
endmodule


