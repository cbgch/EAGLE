//Key = 1101011111001101111111111100101010000100110110011111101110100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393;

XOR2_X1 U771 ( .A(G107), .B(n1063), .Z(G9) );
NOR2_X1 U772 ( .A1(n1064), .A2(n1065), .ZN(G75) );
NOR4_X1 U773 ( .A1(G953), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1065) );
NOR2_X1 U774 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR2_X1 U775 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR3_X1 U776 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
NOR2_X1 U777 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U778 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U779 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR2_X1 U780 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U781 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
AND2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1080) );
NOR2_X1 U784 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NOR3_X1 U786 ( .A1(n1089), .A2(n1094), .A3(n1083), .ZN(n1076) );
NOR2_X1 U787 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR4_X1 U788 ( .A1(n1097), .A2(n1079), .A3(n1083), .A4(n1089), .ZN(n1071) );
NOR2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U790 ( .A1(n1100), .A2(n1075), .ZN(n1098) );
NOR3_X1 U791 ( .A1(n1066), .A2(G953), .A3(G952), .ZN(n1064) );
AND4_X1 U792 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1066) );
NOR4_X1 U793 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1104) );
NOR2_X1 U794 ( .A1(G478), .A2(n1109), .ZN(n1108) );
AND3_X1 U795 ( .A1(n1109), .A2(n1110), .A3(G478), .ZN(n1107) );
INV_X1 U796 ( .A(KEYINPUT10), .ZN(n1109) );
XOR2_X1 U797 ( .A(KEYINPUT27), .B(n1073), .Z(n1106) );
NAND3_X1 U798 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1105) );
XOR2_X1 U799 ( .A(n1114), .B(n1115), .Z(n1112) );
NOR2_X1 U800 ( .A1(G475), .A2(KEYINPUT38), .ZN(n1115) );
XOR2_X1 U801 ( .A(n1116), .B(n1117), .Z(n1111) );
XOR2_X1 U802 ( .A(n1118), .B(KEYINPUT57), .Z(n1117) );
NAND2_X1 U803 ( .A1(KEYINPUT5), .A2(n1119), .ZN(n1116) );
NOR3_X1 U804 ( .A1(n1087), .A2(n1120), .A3(n1121), .ZN(n1103) );
INV_X1 U805 ( .A(n1093), .ZN(n1121) );
NAND2_X1 U806 ( .A1(n1122), .A2(n1123), .ZN(n1102) );
XOR2_X1 U807 ( .A(KEYINPUT9), .B(n1124), .Z(n1101) );
NOR2_X1 U808 ( .A1(n1122), .A2(n1125), .ZN(n1124) );
XOR2_X1 U809 ( .A(n1123), .B(KEYINPUT2), .Z(n1125) );
XOR2_X1 U810 ( .A(n1126), .B(n1127), .Z(G72) );
XOR2_X1 U811 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U812 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XNOR2_X1 U813 ( .A(n1132), .B(n1133), .ZN(n1131) );
XNOR2_X1 U814 ( .A(n1134), .B(n1135), .ZN(n1133) );
NOR2_X1 U815 ( .A1(G900), .A2(n1136), .ZN(n1130) );
NAND2_X1 U816 ( .A1(n1137), .A2(n1136), .ZN(n1128) );
XOR2_X1 U817 ( .A(KEYINPUT30), .B(n1138), .Z(n1137) );
NAND2_X1 U818 ( .A1(G953), .A2(n1139), .ZN(n1126) );
NAND2_X1 U819 ( .A1(G900), .A2(G227), .ZN(n1139) );
XOR2_X1 U820 ( .A(n1140), .B(n1141), .Z(G69) );
NOR2_X1 U821 ( .A1(n1136), .A2(n1142), .ZN(n1141) );
XOR2_X1 U822 ( .A(KEYINPUT60), .B(n1143), .Z(n1142) );
NOR2_X1 U823 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND2_X1 U824 ( .A1(n1146), .A2(n1147), .ZN(n1140) );
NAND2_X1 U825 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U826 ( .A(n1150), .B(n1151), .Z(n1146) );
NOR2_X1 U827 ( .A1(n1152), .A2(G953), .ZN(n1151) );
OR2_X1 U828 ( .A1(n1149), .A2(n1148), .ZN(n1150) );
NAND2_X1 U829 ( .A1(n1153), .A2(n1154), .ZN(n1148) );
NAND2_X1 U830 ( .A1(G953), .A2(n1145), .ZN(n1154) );
XOR2_X1 U831 ( .A(n1155), .B(n1156), .Z(n1153) );
INV_X1 U832 ( .A(KEYINPUT3), .ZN(n1149) );
NOR2_X1 U833 ( .A1(n1157), .A2(n1158), .ZN(G66) );
XNOR2_X1 U834 ( .A(n1159), .B(n1160), .ZN(n1158) );
NOR2_X1 U835 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U836 ( .A1(n1157), .A2(n1163), .ZN(G63) );
XOR2_X1 U837 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U838 ( .A(n1166), .B(KEYINPUT45), .Z(n1165) );
NAND3_X1 U839 ( .A1(n1167), .A2(n1168), .A3(G478), .ZN(n1166) );
NAND2_X1 U840 ( .A1(KEYINPUT18), .A2(n1162), .ZN(n1168) );
NAND2_X1 U841 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
INV_X1 U842 ( .A(KEYINPUT18), .ZN(n1170) );
NAND2_X1 U843 ( .A1(n1171), .A2(G902), .ZN(n1169) );
NOR2_X1 U844 ( .A1(n1157), .A2(n1172), .ZN(G60) );
NOR3_X1 U845 ( .A1(n1114), .A2(n1173), .A3(n1174), .ZN(n1172) );
NOR3_X1 U846 ( .A1(n1175), .A2(n1176), .A3(n1162), .ZN(n1174) );
NOR2_X1 U847 ( .A1(n1177), .A2(n1178), .ZN(n1173) );
NOR2_X1 U848 ( .A1(n1171), .A2(n1176), .ZN(n1177) );
INV_X1 U849 ( .A(G475), .ZN(n1176) );
INV_X1 U850 ( .A(n1068), .ZN(n1171) );
XOR2_X1 U851 ( .A(n1179), .B(G104), .Z(G6) );
NAND2_X1 U852 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NAND3_X1 U853 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1181) );
OR2_X1 U854 ( .A1(n1185), .A2(n1184), .ZN(n1180) );
INV_X1 U855 ( .A(KEYINPUT51), .ZN(n1184) );
NOR2_X1 U856 ( .A1(n1157), .A2(n1186), .ZN(G57) );
XOR2_X1 U857 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U858 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U859 ( .A1(n1191), .A2(n1162), .ZN(n1190) );
INV_X1 U860 ( .A(G472), .ZN(n1191) );
NOR2_X1 U861 ( .A1(n1192), .A2(n1193), .ZN(n1189) );
XOR2_X1 U862 ( .A(KEYINPUT26), .B(n1194), .Z(n1193) );
NOR2_X1 U863 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NOR2_X1 U864 ( .A1(n1197), .A2(n1198), .ZN(n1192) );
XOR2_X1 U865 ( .A(n1199), .B(n1200), .Z(n1187) );
NAND2_X1 U866 ( .A1(KEYINPUT20), .A2(n1201), .ZN(n1199) );
NOR2_X1 U867 ( .A1(n1157), .A2(n1202), .ZN(G54) );
XOR2_X1 U868 ( .A(n1203), .B(n1204), .Z(n1202) );
XOR2_X1 U869 ( .A(n1205), .B(n1206), .Z(n1204) );
NOR2_X1 U870 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U871 ( .A(n1209), .B(KEYINPUT55), .Z(n1208) );
NAND2_X1 U872 ( .A1(n1210), .A2(n1196), .ZN(n1209) );
NOR2_X1 U873 ( .A1(n1196), .A2(n1210), .ZN(n1207) );
XOR2_X1 U874 ( .A(n1211), .B(n1134), .Z(n1210) );
NOR3_X1 U875 ( .A1(n1212), .A2(KEYINPUT34), .A3(n1213), .ZN(n1205) );
INV_X1 U876 ( .A(n1214), .ZN(n1213) );
NAND3_X1 U877 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1212) );
NAND3_X1 U878 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1216) );
NAND3_X1 U879 ( .A1(n1221), .A2(n1219), .A3(G140), .ZN(n1215) );
NOR2_X1 U880 ( .A1(n1119), .A2(n1162), .ZN(n1203) );
INV_X1 U881 ( .A(G469), .ZN(n1119) );
NOR2_X1 U882 ( .A1(n1157), .A2(n1222), .ZN(G51) );
XNOR2_X1 U883 ( .A(n1223), .B(n1224), .ZN(n1222) );
XOR2_X1 U884 ( .A(n1225), .B(n1226), .Z(n1223) );
NOR2_X1 U885 ( .A1(n1227), .A2(n1162), .ZN(n1226) );
NAND2_X1 U886 ( .A1(G902), .A2(n1068), .ZN(n1162) );
NAND2_X1 U887 ( .A1(n1152), .A2(n1138), .ZN(n1068) );
AND4_X1 U888 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1138) );
AND4_X1 U889 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1231) );
NOR2_X1 U890 ( .A1(n1236), .A2(n1237), .ZN(n1230) );
NAND3_X1 U891 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1228) );
NAND2_X1 U892 ( .A1(KEYINPUT61), .A2(n1241), .ZN(n1239) );
NAND2_X1 U893 ( .A1(n1242), .A2(n1243), .ZN(n1238) );
INV_X1 U894 ( .A(KEYINPUT61), .ZN(n1243) );
NAND2_X1 U895 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
AND4_X1 U896 ( .A1(n1246), .A2(n1185), .A3(n1247), .A4(n1248), .ZN(n1152) );
AND4_X1 U897 ( .A1(n1249), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1248) );
NOR3_X1 U898 ( .A1(n1063), .A2(n1253), .A3(n1254), .ZN(n1247) );
NOR3_X1 U899 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1254) );
AND2_X1 U900 ( .A1(n1255), .A2(n1258), .ZN(n1253) );
INV_X1 U901 ( .A(KEYINPUT39), .ZN(n1255) );
AND2_X1 U902 ( .A1(n1095), .A2(n1182), .ZN(n1063) );
NAND2_X1 U903 ( .A1(n1096), .A2(n1182), .ZN(n1185) );
AND3_X1 U904 ( .A1(n1100), .A2(n1259), .A3(n1091), .ZN(n1182) );
NAND2_X1 U905 ( .A1(KEYINPUT50), .A2(n1260), .ZN(n1225) );
XOR2_X1 U906 ( .A(n1261), .B(n1262), .Z(n1260) );
XNOR2_X1 U907 ( .A(G125), .B(n1263), .ZN(n1262) );
NAND2_X1 U908 ( .A1(KEYINPUT63), .A2(n1195), .ZN(n1261) );
NOR2_X1 U909 ( .A1(n1136), .A2(G952), .ZN(n1157) );
XOR2_X1 U910 ( .A(G146), .B(n1237), .Z(G48) );
AND3_X1 U911 ( .A1(n1096), .A2(n1085), .A3(n1264), .ZN(n1237) );
XOR2_X1 U912 ( .A(n1265), .B(n1229), .Z(G45) );
NAND4_X1 U913 ( .A1(n1266), .A2(n1085), .A3(n1267), .A4(n1268), .ZN(n1229) );
XNOR2_X1 U914 ( .A(n1236), .B(n1269), .ZN(G42) );
XOR2_X1 U915 ( .A(KEYINPUT15), .B(G140), .Z(n1269) );
AND4_X1 U916 ( .A1(n1240), .A2(n1099), .A3(n1091), .A4(n1270), .ZN(n1236) );
XNOR2_X1 U917 ( .A(G137), .B(n1235), .ZN(G39) );
NAND3_X1 U918 ( .A1(n1264), .A2(n1271), .A3(n1272), .ZN(n1235) );
XOR2_X1 U919 ( .A(n1234), .B(n1273), .Z(G36) );
NAND2_X1 U920 ( .A1(KEYINPUT41), .A2(G134), .ZN(n1273) );
NAND3_X1 U921 ( .A1(n1266), .A2(n1095), .A3(n1272), .ZN(n1234) );
INV_X1 U922 ( .A(n1089), .ZN(n1272) );
XOR2_X1 U923 ( .A(G131), .B(n1274), .Z(G33) );
AND2_X1 U924 ( .A1(n1266), .A2(n1240), .ZN(n1274) );
NOR2_X1 U925 ( .A1(n1089), .A2(n1183), .ZN(n1240) );
NAND2_X1 U926 ( .A1(n1086), .A2(n1275), .ZN(n1089) );
INV_X1 U927 ( .A(n1241), .ZN(n1266) );
NAND2_X1 U928 ( .A1(n1244), .A2(n1091), .ZN(n1241) );
AND3_X1 U929 ( .A1(n1073), .A2(n1270), .A3(n1113), .ZN(n1244) );
XOR2_X1 U930 ( .A(n1276), .B(n1233), .Z(G30) );
NAND3_X1 U931 ( .A1(n1095), .A2(n1085), .A3(n1264), .ZN(n1233) );
AND4_X1 U932 ( .A1(n1091), .A2(n1073), .A3(n1075), .A4(n1270), .ZN(n1264) );
XOR2_X1 U933 ( .A(n1277), .B(n1252), .Z(G3) );
NAND3_X1 U934 ( .A1(n1271), .A2(n1091), .A3(n1278), .ZN(n1252) );
XOR2_X1 U935 ( .A(n1232), .B(n1279), .Z(G27) );
XNOR2_X1 U936 ( .A(G125), .B(KEYINPUT53), .ZN(n1279) );
NAND4_X1 U937 ( .A1(n1085), .A2(n1270), .A3(n1099), .A4(n1280), .ZN(n1232) );
NOR2_X1 U938 ( .A1(n1083), .A2(n1183), .ZN(n1280) );
NAND2_X1 U939 ( .A1(n1281), .A2(n1070), .ZN(n1270) );
XOR2_X1 U940 ( .A(KEYINPUT58), .B(n1282), .Z(n1281) );
NOR4_X1 U941 ( .A1(G900), .A2(n1283), .A3(n1284), .A4(n1136), .ZN(n1282) );
INV_X1 U942 ( .A(n1285), .ZN(n1283) );
XOR2_X1 U943 ( .A(n1286), .B(n1287), .Z(G24) );
NOR2_X1 U944 ( .A1(n1258), .A2(KEYINPUT31), .ZN(n1287) );
NOR2_X1 U945 ( .A1(n1257), .A2(n1083), .ZN(n1258) );
NAND4_X1 U946 ( .A1(n1100), .A2(n1259), .A3(n1267), .A4(n1268), .ZN(n1257) );
XOR2_X1 U947 ( .A(n1251), .B(n1288), .Z(G21) );
NAND2_X1 U948 ( .A1(KEYINPUT23), .A2(G119), .ZN(n1288) );
NAND4_X1 U949 ( .A1(n1073), .A2(n1075), .A3(n1289), .A4(n1290), .ZN(n1251) );
NOR2_X1 U950 ( .A1(n1079), .A2(n1083), .ZN(n1290) );
INV_X1 U951 ( .A(n1271), .ZN(n1079) );
INV_X1 U952 ( .A(n1113), .ZN(n1075) );
XNOR2_X1 U953 ( .A(G116), .B(n1250), .ZN(G18) );
NAND3_X1 U954 ( .A1(n1256), .A2(n1095), .A3(n1278), .ZN(n1250) );
NOR2_X1 U955 ( .A1(n1267), .A2(n1291), .ZN(n1095) );
XOR2_X1 U956 ( .A(n1292), .B(G113), .Z(G15) );
NAND3_X1 U957 ( .A1(n1293), .A2(n1294), .A3(KEYINPUT0), .ZN(n1292) );
NAND4_X1 U958 ( .A1(n1278), .A2(n1083), .A3(n1096), .A4(n1295), .ZN(n1294) );
OR2_X1 U959 ( .A1(n1246), .A2(n1295), .ZN(n1293) );
INV_X1 U960 ( .A(KEYINPUT43), .ZN(n1295) );
NAND3_X1 U961 ( .A1(n1278), .A2(n1256), .A3(n1096), .ZN(n1246) );
INV_X1 U962 ( .A(n1183), .ZN(n1096) );
NAND2_X1 U963 ( .A1(n1291), .A2(n1267), .ZN(n1183) );
INV_X1 U964 ( .A(n1083), .ZN(n1256) );
NAND2_X1 U965 ( .A1(n1296), .A2(n1093), .ZN(n1083) );
AND2_X1 U966 ( .A1(n1259), .A2(n1073), .ZN(n1278) );
AND2_X1 U967 ( .A1(n1289), .A2(n1113), .ZN(n1259) );
NAND2_X1 U968 ( .A1(n1297), .A2(n1298), .ZN(G12) );
NAND2_X1 U969 ( .A1(n1299), .A2(n1219), .ZN(n1298) );
XOR2_X1 U970 ( .A(KEYINPUT12), .B(n1300), .Z(n1297) );
NOR2_X1 U971 ( .A1(n1299), .A2(n1219), .ZN(n1300) );
INV_X1 U972 ( .A(n1249), .ZN(n1299) );
NAND4_X1 U973 ( .A1(n1271), .A2(n1099), .A3(n1091), .A4(n1289), .ZN(n1249) );
AND2_X1 U974 ( .A1(n1085), .A2(n1301), .ZN(n1289) );
NAND2_X1 U975 ( .A1(n1070), .A2(n1302), .ZN(n1301) );
NAND4_X1 U976 ( .A1(G953), .A2(G902), .A3(n1285), .A4(n1145), .ZN(n1302) );
INV_X1 U977 ( .A(G898), .ZN(n1145) );
NAND3_X1 U978 ( .A1(n1285), .A2(n1136), .A3(G952), .ZN(n1070) );
NAND2_X1 U979 ( .A1(G237), .A2(G234), .ZN(n1285) );
NOR2_X1 U980 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
INV_X1 U981 ( .A(n1275), .ZN(n1087) );
NAND2_X1 U982 ( .A1(G214), .A2(n1303), .ZN(n1275) );
XOR2_X1 U983 ( .A(n1123), .B(n1122), .Z(n1086) );
INV_X1 U984 ( .A(n1227), .ZN(n1122) );
NAND2_X1 U985 ( .A1(G210), .A2(n1303), .ZN(n1227) );
NAND2_X1 U986 ( .A1(n1304), .A2(n1284), .ZN(n1303) );
NAND2_X1 U987 ( .A1(n1305), .A2(n1284), .ZN(n1123) );
XOR2_X1 U988 ( .A(n1306), .B(n1307), .Z(n1305) );
XOR2_X1 U989 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U990 ( .A(KEYINPUT8), .B(n1263), .Z(n1309) );
NOR2_X1 U991 ( .A1(n1144), .A2(G953), .ZN(n1263) );
INV_X1 U992 ( .A(G224), .ZN(n1144) );
NOR2_X1 U993 ( .A1(G125), .A2(KEYINPUT14), .ZN(n1308) );
XOR2_X1 U994 ( .A(n1224), .B(n1198), .Z(n1306) );
INV_X1 U995 ( .A(n1195), .ZN(n1198) );
NAND2_X1 U996 ( .A1(n1310), .A2(n1311), .ZN(n1224) );
NAND2_X1 U997 ( .A1(n1156), .A2(n1155), .ZN(n1311) );
NAND2_X1 U998 ( .A1(n1312), .A2(n1313), .ZN(n1310) );
XOR2_X1 U999 ( .A(n1156), .B(KEYINPUT24), .Z(n1313) );
XOR2_X1 U1000 ( .A(n1314), .B(n1315), .Z(n1156) );
XOR2_X1 U1001 ( .A(G110), .B(n1316), .Z(n1315) );
XOR2_X1 U1002 ( .A(G122), .B(G113), .Z(n1316) );
XOR2_X1 U1003 ( .A(n1317), .B(n1318), .Z(n1314) );
NAND2_X1 U1004 ( .A1(KEYINPUT47), .A2(G119), .ZN(n1317) );
INV_X1 U1005 ( .A(n1155), .ZN(n1312) );
XOR2_X1 U1006 ( .A(n1319), .B(n1320), .Z(n1155) );
NAND2_X1 U1007 ( .A1(KEYINPUT49), .A2(n1277), .ZN(n1319) );
INV_X1 U1008 ( .A(n1245), .ZN(n1091) );
NAND2_X1 U1009 ( .A1(n1092), .A2(n1093), .ZN(n1245) );
NAND2_X1 U1010 ( .A1(G221), .A2(n1321), .ZN(n1093) );
INV_X1 U1011 ( .A(n1296), .ZN(n1092) );
XOR2_X1 U1012 ( .A(n1118), .B(G469), .Z(n1296) );
NAND3_X1 U1013 ( .A1(n1322), .A2(n1284), .A3(n1323), .ZN(n1118) );
NAND2_X1 U1014 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
XOR2_X1 U1015 ( .A(KEYINPUT35), .B(n1326), .Z(n1325) );
XOR2_X1 U1016 ( .A(n1327), .B(n1211), .Z(n1324) );
NAND2_X1 U1017 ( .A1(n1328), .A2(n1329), .ZN(n1322) );
XNOR2_X1 U1018 ( .A(n1211), .B(n1327), .ZN(n1329) );
XNOR2_X1 U1019 ( .A(n1330), .B(n1331), .ZN(n1327) );
NAND2_X1 U1020 ( .A1(KEYINPUT21), .A2(n1134), .ZN(n1331) );
XNOR2_X1 U1021 ( .A(n1276), .B(n1332), .ZN(n1134) );
NAND2_X1 U1022 ( .A1(KEYINPUT19), .A2(n1196), .ZN(n1330) );
XNOR2_X1 U1023 ( .A(n1277), .B(n1320), .ZN(n1211) );
XOR2_X1 U1024 ( .A(G104), .B(n1333), .Z(n1320) );
INV_X1 U1025 ( .A(G101), .ZN(n1277) );
XOR2_X1 U1026 ( .A(KEYINPUT6), .B(n1326), .Z(n1328) );
AND4_X1 U1027 ( .A1(n1217), .A2(n1214), .A3(n1334), .A4(n1335), .ZN(n1326) );
NAND3_X1 U1028 ( .A1(n1336), .A2(n1219), .A3(n1221), .ZN(n1335) );
XOR2_X1 U1029 ( .A(KEYINPUT13), .B(n1220), .Z(n1336) );
NAND3_X1 U1030 ( .A1(n1337), .A2(n1219), .A3(n1218), .ZN(n1334) );
INV_X1 U1031 ( .A(G110), .ZN(n1219) );
XOR2_X1 U1032 ( .A(KEYINPUT13), .B(G140), .Z(n1337) );
NAND3_X1 U1033 ( .A1(n1221), .A2(n1220), .A3(G110), .ZN(n1214) );
INV_X1 U1034 ( .A(G140), .ZN(n1220) );
NAND3_X1 U1035 ( .A1(G110), .A2(G140), .A3(n1218), .ZN(n1217) );
INV_X1 U1036 ( .A(n1221), .ZN(n1218) );
NAND2_X1 U1037 ( .A1(G227), .A2(n1136), .ZN(n1221) );
NOR2_X1 U1038 ( .A1(n1073), .A2(n1113), .ZN(n1099) );
XNOR2_X1 U1039 ( .A(n1338), .B(n1161), .ZN(n1113) );
NAND2_X1 U1040 ( .A1(G217), .A2(n1321), .ZN(n1161) );
NAND2_X1 U1041 ( .A1(G234), .A2(n1284), .ZN(n1321) );
NAND2_X1 U1042 ( .A1(n1159), .A2(n1284), .ZN(n1338) );
XNOR2_X1 U1043 ( .A(n1339), .B(n1340), .ZN(n1159) );
XOR2_X1 U1044 ( .A(n1341), .B(n1342), .Z(n1340) );
NOR2_X1 U1045 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
XOR2_X1 U1046 ( .A(n1345), .B(KEYINPUT40), .Z(n1344) );
NAND2_X1 U1047 ( .A1(G110), .A2(n1346), .ZN(n1345) );
XOR2_X1 U1048 ( .A(KEYINPUT42), .B(n1347), .Z(n1346) );
NOR2_X1 U1049 ( .A1(G110), .A2(n1347), .ZN(n1343) );
XOR2_X1 U1050 ( .A(G119), .B(G128), .Z(n1347) );
NOR2_X1 U1051 ( .A1(KEYINPUT59), .A2(n1348), .ZN(n1341) );
XOR2_X1 U1052 ( .A(n1349), .B(n1350), .Z(n1348) );
XOR2_X1 U1053 ( .A(KEYINPUT22), .B(n1351), .Z(n1350) );
AND3_X1 U1054 ( .A1(G221), .A2(n1136), .A3(G234), .ZN(n1351) );
NOR2_X1 U1055 ( .A1(G137), .A2(KEYINPUT46), .ZN(n1349) );
NAND3_X1 U1056 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1339) );
NAND2_X1 U1057 ( .A1(G146), .A2(n1355), .ZN(n1354) );
OR3_X1 U1058 ( .A1(n1355), .A2(G146), .A3(KEYINPUT11), .ZN(n1353) );
NAND2_X1 U1059 ( .A1(KEYINPUT28), .A2(n1356), .ZN(n1355) );
NAND2_X1 U1060 ( .A1(KEYINPUT11), .A2(n1357), .ZN(n1352) );
INV_X1 U1061 ( .A(n1356), .ZN(n1357) );
INV_X1 U1062 ( .A(n1100), .ZN(n1073) );
XOR2_X1 U1063 ( .A(n1358), .B(G472), .Z(n1100) );
NAND2_X1 U1064 ( .A1(n1359), .A2(n1284), .ZN(n1358) );
XOR2_X1 U1065 ( .A(n1360), .B(n1361), .Z(n1359) );
XOR2_X1 U1066 ( .A(n1362), .B(n1196), .Z(n1361) );
INV_X1 U1067 ( .A(n1197), .ZN(n1196) );
XOR2_X1 U1068 ( .A(n1363), .B(n1364), .Z(n1197) );
XOR2_X1 U1069 ( .A(KEYINPUT16), .B(G131), .Z(n1364) );
NAND2_X1 U1070 ( .A1(KEYINPUT37), .A2(n1135), .ZN(n1363) );
XOR2_X1 U1071 ( .A(G134), .B(G137), .Z(n1135) );
XOR2_X1 U1072 ( .A(n1200), .B(n1195), .Z(n1362) );
XNOR2_X1 U1073 ( .A(n1332), .B(n1365), .ZN(n1195) );
NOR2_X1 U1074 ( .A1(KEYINPUT36), .A2(n1276), .ZN(n1365) );
INV_X1 U1075 ( .A(G128), .ZN(n1276) );
XOR2_X1 U1076 ( .A(n1265), .B(n1366), .Z(n1332) );
INV_X1 U1077 ( .A(G146), .ZN(n1366) );
XNOR2_X1 U1078 ( .A(n1367), .B(n1368), .ZN(n1200) );
XOR2_X1 U1079 ( .A(KEYINPUT4), .B(G113), .Z(n1368) );
XOR2_X1 U1080 ( .A(n1369), .B(G101), .Z(n1367) );
NAND2_X1 U1081 ( .A1(KEYINPUT62), .A2(n1370), .ZN(n1369) );
XNOR2_X1 U1082 ( .A(n1371), .B(n1318), .ZN(n1370) );
NAND2_X1 U1083 ( .A1(KEYINPUT48), .A2(n1372), .ZN(n1371) );
INV_X1 U1084 ( .A(G119), .ZN(n1372) );
XOR2_X1 U1085 ( .A(n1373), .B(n1374), .Z(n1360) );
XOR2_X1 U1086 ( .A(KEYINPUT1), .B(n1201), .Z(n1374) );
AND3_X1 U1087 ( .A1(n1304), .A2(n1136), .A3(G210), .ZN(n1201) );
XNOR2_X1 U1088 ( .A(KEYINPUT33), .B(KEYINPUT29), .ZN(n1373) );
NOR2_X1 U1089 ( .A1(n1268), .A2(n1267), .ZN(n1271) );
XOR2_X1 U1090 ( .A(n1114), .B(G475), .Z(n1267) );
NOR2_X1 U1091 ( .A1(n1178), .A2(G902), .ZN(n1114) );
INV_X1 U1092 ( .A(n1175), .ZN(n1178) );
XOR2_X1 U1093 ( .A(n1375), .B(n1376), .Z(n1175) );
XNOR2_X1 U1094 ( .A(G104), .B(n1377), .ZN(n1376) );
NAND2_X1 U1095 ( .A1(n1378), .A2(KEYINPUT25), .ZN(n1377) );
XOR2_X1 U1096 ( .A(n1379), .B(n1380), .Z(n1378) );
XOR2_X1 U1097 ( .A(KEYINPUT52), .B(G146), .Z(n1380) );
XOR2_X1 U1098 ( .A(n1381), .B(n1132), .Z(n1379) );
XOR2_X1 U1099 ( .A(G131), .B(n1356), .Z(n1132) );
XOR2_X1 U1100 ( .A(G125), .B(G140), .Z(n1356) );
NAND2_X1 U1101 ( .A1(n1382), .A2(KEYINPUT44), .ZN(n1381) );
XOR2_X1 U1102 ( .A(n1265), .B(n1383), .Z(n1382) );
AND3_X1 U1103 ( .A1(G214), .A2(n1136), .A3(n1304), .ZN(n1383) );
INV_X1 U1104 ( .A(G237), .ZN(n1304) );
INV_X1 U1105 ( .A(G143), .ZN(n1265) );
XOR2_X1 U1106 ( .A(G113), .B(n1286), .Z(n1375) );
INV_X1 U1107 ( .A(n1291), .ZN(n1268) );
NOR2_X1 U1108 ( .A1(n1384), .A2(n1120), .ZN(n1291) );
NOR2_X1 U1109 ( .A1(n1110), .A2(G478), .ZN(n1120) );
AND2_X1 U1110 ( .A1(G478), .A2(n1110), .ZN(n1384) );
NAND2_X1 U1111 ( .A1(n1164), .A2(n1284), .ZN(n1110) );
INV_X1 U1112 ( .A(G902), .ZN(n1284) );
XOR2_X1 U1113 ( .A(n1385), .B(n1386), .Z(n1164) );
XOR2_X1 U1114 ( .A(G128), .B(n1387), .Z(n1386) );
AND3_X1 U1115 ( .A1(G234), .A2(n1136), .A3(G217), .ZN(n1387) );
INV_X1 U1116 ( .A(G953), .ZN(n1136) );
XOR2_X1 U1117 ( .A(n1388), .B(n1389), .Z(n1385) );
XOR2_X1 U1118 ( .A(n1390), .B(n1391), .Z(n1389) );
XOR2_X1 U1119 ( .A(n1392), .B(n1333), .Z(n1391) );
XOR2_X1 U1120 ( .A(G107), .B(KEYINPUT32), .Z(n1333) );
XNOR2_X1 U1121 ( .A(G134), .B(n1318), .ZN(n1392) );
XOR2_X1 U1122 ( .A(G116), .B(KEYINPUT17), .Z(n1318) );
XOR2_X1 U1123 ( .A(n1393), .B(G143), .Z(n1390) );
XNOR2_X1 U1124 ( .A(KEYINPUT56), .B(KEYINPUT54), .ZN(n1393) );
NAND2_X1 U1125 ( .A1(KEYINPUT7), .A2(n1286), .ZN(n1388) );
INV_X1 U1126 ( .A(G122), .ZN(n1286) );
endmodule


