//Key = 1011100011110101110000101110110001000100101000011101000011000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362;

XNOR2_X1 U756 ( .A(G107), .B(n1046), .ZN(G9) );
NAND2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U758 ( .A1(n1049), .A2(n1050), .ZN(G75) );
NOR4_X1 U759 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1050) );
NOR4_X1 U760 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1053) );
NOR4_X1 U761 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1056) );
AND2_X1 U762 ( .A1(n1047), .A2(n1063), .ZN(n1062) );
NOR2_X1 U763 ( .A1(n1064), .A2(n1065), .ZN(n1061) );
NOR2_X1 U764 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
AND2_X1 U765 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U766 ( .A1(KEYINPUT58), .A2(n1070), .ZN(n1060) );
NOR2_X1 U767 ( .A1(n1071), .A2(n1072), .ZN(n1055) );
AND2_X1 U768 ( .A1(n1073), .A2(KEYINPUT58), .ZN(n1072) );
NAND3_X1 U769 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1051) );
NAND4_X1 U770 ( .A1(n1071), .A2(n1063), .A3(n1077), .A4(n1078), .ZN(n1076) );
NAND2_X1 U771 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND3_X1 U772 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1080) );
NAND2_X1 U773 ( .A1(n1057), .A2(n1084), .ZN(n1082) );
INV_X1 U774 ( .A(n1085), .ZN(n1057) );
NAND3_X1 U775 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1081) );
NAND2_X1 U776 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NAND2_X1 U777 ( .A1(n1091), .A2(n1085), .ZN(n1079) );
INV_X1 U778 ( .A(n1059), .ZN(n1071) );
NOR3_X1 U779 ( .A1(n1092), .A2(G953), .A3(n1093), .ZN(n1049) );
XNOR2_X1 U780 ( .A(KEYINPUT20), .B(n1054), .ZN(n1093) );
INV_X1 U781 ( .A(G952), .ZN(n1054) );
XNOR2_X1 U782 ( .A(KEYINPUT19), .B(n1074), .ZN(n1092) );
NAND4_X1 U783 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1074) );
NOR4_X1 U784 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
XNOR2_X1 U785 ( .A(n1102), .B(n1103), .ZN(n1101) );
XNOR2_X1 U786 ( .A(n1104), .B(KEYINPUT40), .ZN(n1098) );
NOR2_X1 U787 ( .A1(n1069), .A2(n1089), .ZN(n1096) );
XNOR2_X1 U788 ( .A(n1105), .B(n1106), .ZN(n1095) );
NOR2_X1 U789 ( .A1(G469), .A2(KEYINPUT50), .ZN(n1106) );
XNOR2_X1 U790 ( .A(n1107), .B(n1108), .ZN(n1094) );
NOR2_X1 U791 ( .A1(n1109), .A2(KEYINPUT39), .ZN(n1108) );
XOR2_X1 U792 ( .A(n1110), .B(n1111), .Z(G72) );
XOR2_X1 U793 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND2_X1 U794 ( .A1(G953), .A2(n1114), .ZN(n1113) );
NAND2_X1 U795 ( .A1(G900), .A2(G227), .ZN(n1114) );
NAND2_X1 U796 ( .A1(n1115), .A2(n1116), .ZN(n1112) );
NAND2_X1 U797 ( .A1(G953), .A2(n1117), .ZN(n1116) );
XOR2_X1 U798 ( .A(n1118), .B(n1119), .Z(n1115) );
NAND2_X1 U799 ( .A1(KEYINPUT33), .A2(n1120), .ZN(n1118) );
XOR2_X1 U800 ( .A(n1121), .B(n1122), .Z(n1120) );
XNOR2_X1 U801 ( .A(n1123), .B(n1124), .ZN(n1122) );
NAND2_X1 U802 ( .A1(KEYINPUT4), .A2(n1125), .ZN(n1123) );
NOR2_X1 U803 ( .A1(n1126), .A2(G953), .ZN(n1110) );
XOR2_X1 U804 ( .A(n1127), .B(n1128), .Z(G69) );
XOR2_X1 U805 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U806 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XNOR2_X1 U807 ( .A(n1133), .B(KEYINPUT22), .ZN(n1132) );
NOR2_X1 U808 ( .A1(G898), .A2(n1075), .ZN(n1131) );
NOR2_X1 U809 ( .A1(G953), .A2(n1134), .ZN(n1129) );
NOR3_X1 U810 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1134) );
XOR2_X1 U811 ( .A(n1138), .B(KEYINPUT17), .Z(n1137) );
NOR2_X1 U812 ( .A1(n1139), .A2(n1075), .ZN(n1127) );
AND2_X1 U813 ( .A1(G224), .A2(G898), .ZN(n1139) );
NOR2_X1 U814 ( .A1(n1140), .A2(n1141), .ZN(G66) );
NOR3_X1 U815 ( .A1(n1102), .A2(n1142), .A3(n1143), .ZN(n1141) );
NOR3_X1 U816 ( .A1(n1144), .A2(n1103), .A3(n1145), .ZN(n1143) );
NOR2_X1 U817 ( .A1(n1146), .A2(n1147), .ZN(n1142) );
NOR2_X1 U818 ( .A1(n1148), .A2(n1103), .ZN(n1146) );
INV_X1 U819 ( .A(n1052), .ZN(n1148) );
NOR2_X1 U820 ( .A1(n1140), .A2(n1149), .ZN(G63) );
XOR2_X1 U821 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U822 ( .A1(n1107), .A2(n1145), .ZN(n1151) );
NAND2_X1 U823 ( .A1(KEYINPUT9), .A2(n1152), .ZN(n1150) );
NOR2_X1 U824 ( .A1(n1140), .A2(n1153), .ZN(G60) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U826 ( .A1(n1156), .A2(n1145), .ZN(n1154) );
XNOR2_X1 U827 ( .A(n1157), .B(n1158), .ZN(G6) );
NAND2_X1 U828 ( .A1(n1159), .A2(KEYINPUT62), .ZN(n1158) );
XNOR2_X1 U829 ( .A(G104), .B(KEYINPUT51), .ZN(n1159) );
NOR2_X1 U830 ( .A1(n1140), .A2(n1160), .ZN(G57) );
XOR2_X1 U831 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U832 ( .A(n1125), .B(n1163), .ZN(n1162) );
XOR2_X1 U833 ( .A(n1164), .B(n1165), .Z(n1161) );
XOR2_X1 U834 ( .A(n1166), .B(n1167), .Z(n1164) );
NOR2_X1 U835 ( .A1(n1168), .A2(n1145), .ZN(n1167) );
XNOR2_X1 U836 ( .A(G472), .B(KEYINPUT12), .ZN(n1168) );
NOR3_X1 U837 ( .A1(n1169), .A2(n1170), .A3(n1171), .ZN(G54) );
NOR3_X1 U838 ( .A1(n1172), .A2(G953), .A3(G952), .ZN(n1171) );
AND2_X1 U839 ( .A1(n1172), .A2(n1140), .ZN(n1170) );
INV_X1 U840 ( .A(KEYINPUT43), .ZN(n1172) );
XOR2_X1 U841 ( .A(n1173), .B(n1174), .Z(n1169) );
XNOR2_X1 U842 ( .A(n1175), .B(n1176), .ZN(n1174) );
NAND3_X1 U843 ( .A1(G469), .A2(n1052), .A3(n1177), .ZN(n1175) );
XNOR2_X1 U844 ( .A(G902), .B(KEYINPUT3), .ZN(n1177) );
XOR2_X1 U845 ( .A(n1178), .B(n1179), .Z(n1173) );
NOR2_X1 U846 ( .A1(KEYINPUT32), .A2(n1125), .ZN(n1179) );
XNOR2_X1 U847 ( .A(n1180), .B(n1181), .ZN(n1178) );
NAND2_X1 U848 ( .A1(KEYINPUT29), .A2(n1182), .ZN(n1180) );
XOR2_X1 U849 ( .A(G140), .B(G110), .Z(n1182) );
NOR2_X1 U850 ( .A1(n1140), .A2(n1183), .ZN(G51) );
XOR2_X1 U851 ( .A(n1184), .B(n1185), .Z(n1183) );
XOR2_X1 U852 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U853 ( .A(n1188), .B(n1166), .Z(n1187) );
NOR2_X1 U854 ( .A1(n1189), .A2(n1145), .ZN(n1186) );
NAND2_X1 U855 ( .A1(G902), .A2(n1052), .ZN(n1145) );
NAND4_X1 U856 ( .A1(n1126), .A2(n1190), .A3(n1191), .A4(n1138), .ZN(n1052) );
NAND4_X1 U857 ( .A1(n1047), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1138) );
NAND2_X1 U858 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
INV_X1 U859 ( .A(KEYINPUT31), .ZN(n1196) );
NAND2_X1 U860 ( .A1(KEYINPUT31), .A2(n1197), .ZN(n1193) );
NAND2_X1 U861 ( .A1(n1198), .A2(n1087), .ZN(n1197) );
XOR2_X1 U862 ( .A(KEYINPUT28), .B(n1136), .Z(n1191) );
INV_X1 U863 ( .A(n1135), .ZN(n1190) );
NAND4_X1 U864 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1135) );
NOR3_X1 U865 ( .A1(n1203), .A2(n1204), .A3(n1157), .ZN(n1202) );
AND2_X1 U866 ( .A1(n1205), .A2(n1048), .ZN(n1157) );
NOR2_X1 U867 ( .A1(n1195), .A2(n1058), .ZN(n1048) );
INV_X1 U868 ( .A(n1192), .ZN(n1058) );
NOR4_X1 U869 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1070), .ZN(n1203) );
XNOR2_X1 U870 ( .A(n1209), .B(KEYINPUT7), .ZN(n1207) );
AND4_X1 U871 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1126) );
AND4_X1 U872 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1213) );
AND2_X1 U873 ( .A1(n1218), .A2(n1219), .ZN(n1212) );
XOR2_X1 U874 ( .A(n1220), .B(n1221), .Z(n1184) );
NOR2_X1 U875 ( .A1(G125), .A2(KEYINPUT52), .ZN(n1221) );
NAND2_X1 U876 ( .A1(KEYINPUT0), .A2(n1133), .ZN(n1220) );
NOR2_X1 U877 ( .A1(n1075), .A2(G952), .ZN(n1140) );
XNOR2_X1 U878 ( .A(G146), .B(n1218), .ZN(G48) );
NAND3_X1 U879 ( .A1(n1222), .A2(n1209), .A3(n1205), .ZN(n1218) );
XOR2_X1 U880 ( .A(n1210), .B(n1223), .Z(G45) );
NAND2_X1 U881 ( .A1(KEYINPUT48), .A2(G143), .ZN(n1223) );
NAND4_X1 U882 ( .A1(n1224), .A2(n1209), .A3(n1104), .A4(n1225), .ZN(n1210) );
XNOR2_X1 U883 ( .A(n1211), .B(n1226), .ZN(G42) );
NOR2_X1 U884 ( .A1(KEYINPUT23), .A2(n1227), .ZN(n1226) );
XOR2_X1 U885 ( .A(KEYINPUT13), .B(G140), .Z(n1227) );
NAND4_X1 U886 ( .A1(n1205), .A2(n1228), .A3(n1083), .A4(n1085), .ZN(n1211) );
XNOR2_X1 U887 ( .A(G137), .B(n1217), .ZN(G39) );
NAND3_X1 U888 ( .A1(n1222), .A2(n1085), .A3(n1077), .ZN(n1217) );
XOR2_X1 U889 ( .A(n1216), .B(n1229), .Z(G36) );
NOR2_X1 U890 ( .A1(G134), .A2(KEYINPUT18), .ZN(n1229) );
NAND3_X1 U891 ( .A1(n1047), .A2(n1085), .A3(n1224), .ZN(n1216) );
XNOR2_X1 U892 ( .A(G131), .B(n1215), .ZN(G33) );
NAND3_X1 U893 ( .A1(n1224), .A2(n1085), .A3(n1205), .ZN(n1215) );
NAND2_X1 U894 ( .A1(n1230), .A2(n1231), .ZN(n1085) );
OR2_X1 U895 ( .A1(n1087), .A2(KEYINPUT42), .ZN(n1231) );
NAND3_X1 U896 ( .A1(n1090), .A2(n1232), .A3(KEYINPUT42), .ZN(n1230) );
AND3_X1 U897 ( .A1(n1067), .A2(n1233), .A3(n1091), .ZN(n1224) );
XNOR2_X1 U898 ( .A(G128), .B(n1214), .ZN(G30) );
NAND3_X1 U899 ( .A1(n1047), .A2(n1209), .A3(n1222), .ZN(n1214) );
AND2_X1 U900 ( .A1(n1228), .A2(n1099), .ZN(n1222) );
AND3_X1 U901 ( .A1(n1084), .A2(n1233), .A3(n1067), .ZN(n1228) );
NAND3_X1 U902 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(G3) );
OR2_X1 U903 ( .A1(n1237), .A2(n1204), .ZN(n1236) );
NAND2_X1 U904 ( .A1(KEYINPUT53), .A2(n1238), .ZN(n1235) );
NAND2_X1 U905 ( .A1(n1239), .A2(n1237), .ZN(n1238) );
XNOR2_X1 U906 ( .A(n1204), .B(KEYINPUT49), .ZN(n1239) );
NAND2_X1 U907 ( .A1(n1240), .A2(n1241), .ZN(n1234) );
INV_X1 U908 ( .A(KEYINPUT53), .ZN(n1241) );
NAND2_X1 U909 ( .A1(n1242), .A2(n1243), .ZN(n1240) );
OR2_X1 U910 ( .A1(n1204), .A2(KEYINPUT49), .ZN(n1243) );
NAND3_X1 U911 ( .A1(n1204), .A2(n1237), .A3(KEYINPUT49), .ZN(n1242) );
NOR3_X1 U912 ( .A1(n1208), .A2(n1195), .A3(n1065), .ZN(n1204) );
INV_X1 U913 ( .A(n1091), .ZN(n1208) );
XNOR2_X1 U914 ( .A(G125), .B(n1219), .ZN(G27) );
NAND3_X1 U915 ( .A1(n1083), .A2(n1073), .A3(n1244), .ZN(n1219) );
AND3_X1 U916 ( .A1(n1209), .A2(n1233), .A3(n1084), .ZN(n1244) );
NAND2_X1 U917 ( .A1(n1059), .A2(n1245), .ZN(n1233) );
NAND4_X1 U918 ( .A1(G953), .A2(G902), .A3(n1246), .A4(n1117), .ZN(n1245) );
INV_X1 U919 ( .A(G900), .ZN(n1117) );
XNOR2_X1 U920 ( .A(G122), .B(n1201), .ZN(G24) );
NAND4_X1 U921 ( .A1(n1247), .A2(n1192), .A3(n1104), .A4(n1225), .ZN(n1201) );
NOR2_X1 U922 ( .A1(n1084), .A2(n1099), .ZN(n1192) );
NAND3_X1 U923 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(G21) );
OR2_X1 U924 ( .A1(n1199), .A2(G119), .ZN(n1250) );
NAND2_X1 U925 ( .A1(KEYINPUT54), .A2(n1251), .ZN(n1249) );
NAND2_X1 U926 ( .A1(G119), .A2(n1252), .ZN(n1251) );
XNOR2_X1 U927 ( .A(KEYINPUT37), .B(n1199), .ZN(n1252) );
NAND2_X1 U928 ( .A1(n1253), .A2(n1254), .ZN(n1248) );
INV_X1 U929 ( .A(KEYINPUT54), .ZN(n1254) );
NAND2_X1 U930 ( .A1(n1255), .A2(n1256), .ZN(n1253) );
NAND3_X1 U931 ( .A1(KEYINPUT37), .A2(G119), .A3(n1199), .ZN(n1256) );
OR2_X1 U932 ( .A1(n1199), .A2(KEYINPUT37), .ZN(n1255) );
NAND4_X1 U933 ( .A1(n1247), .A2(n1077), .A3(n1099), .A4(n1084), .ZN(n1199) );
XOR2_X1 U934 ( .A(n1200), .B(n1257), .Z(G18) );
NOR2_X1 U935 ( .A1(G116), .A2(KEYINPUT34), .ZN(n1257) );
NAND3_X1 U936 ( .A1(n1091), .A2(n1047), .A3(n1247), .ZN(n1200) );
NOR3_X1 U937 ( .A1(n1087), .A2(n1206), .A3(n1258), .ZN(n1247) );
INV_X1 U938 ( .A(n1259), .ZN(n1206) );
INV_X1 U939 ( .A(n1209), .ZN(n1087) );
NOR2_X1 U940 ( .A1(n1104), .A2(n1260), .ZN(n1047) );
XNOR2_X1 U941 ( .A(G113), .B(n1261), .ZN(G15) );
NAND4_X1 U942 ( .A1(n1073), .A2(n1091), .A3(n1209), .A4(n1259), .ZN(n1261) );
NOR2_X1 U943 ( .A1(n1084), .A2(n1083), .ZN(n1091) );
INV_X1 U944 ( .A(n1099), .ZN(n1083) );
INV_X1 U945 ( .A(n1070), .ZN(n1073) );
NAND2_X1 U946 ( .A1(n1063), .A2(n1205), .ZN(n1070) );
AND2_X1 U947 ( .A1(n1260), .A2(n1104), .ZN(n1205) );
INV_X1 U948 ( .A(n1225), .ZN(n1260) );
INV_X1 U949 ( .A(n1258), .ZN(n1063) );
NAND2_X1 U950 ( .A1(n1068), .A2(n1262), .ZN(n1258) );
XOR2_X1 U951 ( .A(G110), .B(n1136), .Z(G12) );
NOR4_X1 U952 ( .A1(n1065), .A2(n1195), .A3(n1099), .A4(n1088), .ZN(n1136) );
INV_X1 U953 ( .A(n1084), .ZN(n1088) );
XOR2_X1 U954 ( .A(n1102), .B(n1263), .Z(n1084) );
NOR2_X1 U955 ( .A1(KEYINPUT63), .A2(n1103), .ZN(n1263) );
NAND2_X1 U956 ( .A1(G217), .A2(n1264), .ZN(n1103) );
NOR2_X1 U957 ( .A1(n1147), .A2(G902), .ZN(n1102) );
INV_X1 U958 ( .A(n1144), .ZN(n1147) );
XNOR2_X1 U959 ( .A(n1265), .B(n1266), .ZN(n1144) );
XOR2_X1 U960 ( .A(n1267), .B(n1268), .Z(n1266) );
NAND2_X1 U961 ( .A1(KEYINPUT16), .A2(G137), .ZN(n1268) );
NAND2_X1 U962 ( .A1(n1269), .A2(n1270), .ZN(n1267) );
NAND2_X1 U963 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XOR2_X1 U964 ( .A(n1273), .B(KEYINPUT38), .Z(n1269) );
OR2_X1 U965 ( .A1(n1272), .A2(n1271), .ZN(n1273) );
XOR2_X1 U966 ( .A(n1274), .B(n1275), .Z(n1271) );
XOR2_X1 U967 ( .A(KEYINPUT57), .B(G119), .Z(n1275) );
XOR2_X1 U968 ( .A(n1276), .B(G110), .Z(n1274) );
NAND2_X1 U969 ( .A1(KEYINPUT26), .A2(n1124), .ZN(n1276) );
XNOR2_X1 U970 ( .A(n1277), .B(n1278), .ZN(n1272) );
XOR2_X1 U971 ( .A(KEYINPUT35), .B(KEYINPUT27), .Z(n1278) );
XOR2_X1 U972 ( .A(G146), .B(n1119), .Z(n1277) );
XOR2_X1 U973 ( .A(n1279), .B(KEYINPUT56), .Z(n1265) );
NAND2_X1 U974 ( .A1(G221), .A2(n1280), .ZN(n1279) );
XNOR2_X1 U975 ( .A(n1281), .B(G472), .ZN(n1099) );
NAND2_X1 U976 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
XNOR2_X1 U977 ( .A(n1165), .B(n1284), .ZN(n1282) );
NOR2_X1 U978 ( .A1(KEYINPUT1), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U979 ( .A(n1286), .B(n1125), .ZN(n1285) );
INV_X1 U980 ( .A(n1287), .ZN(n1125) );
XNOR2_X1 U981 ( .A(n1288), .B(n1289), .ZN(n1286) );
NOR2_X1 U982 ( .A1(KEYINPUT60), .A2(n1163), .ZN(n1289) );
XOR2_X1 U983 ( .A(n1290), .B(n1291), .Z(n1163) );
NOR2_X1 U984 ( .A1(KEYINPUT59), .A2(n1292), .ZN(n1291) );
XNOR2_X1 U985 ( .A(G116), .B(G119), .ZN(n1290) );
NOR2_X1 U986 ( .A1(KEYINPUT36), .A2(n1166), .ZN(n1288) );
XOR2_X1 U987 ( .A(G101), .B(n1293), .Z(n1165) );
AND3_X1 U988 ( .A1(G210), .A2(n1075), .A3(n1294), .ZN(n1293) );
NAND2_X1 U989 ( .A1(n1209), .A2(n1198), .ZN(n1195) );
AND2_X1 U990 ( .A1(n1067), .A2(n1259), .ZN(n1198) );
NAND2_X1 U991 ( .A1(n1059), .A2(n1295), .ZN(n1259) );
NAND4_X1 U992 ( .A1(G953), .A2(G902), .A3(n1246), .A4(n1296), .ZN(n1295) );
INV_X1 U993 ( .A(G898), .ZN(n1296) );
NAND3_X1 U994 ( .A1(n1246), .A2(n1075), .A3(G952), .ZN(n1059) );
NAND2_X1 U995 ( .A1(G237), .A2(G234), .ZN(n1246) );
NOR2_X1 U996 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
INV_X1 U997 ( .A(n1262), .ZN(n1069) );
NAND2_X1 U998 ( .A1(G221), .A2(n1264), .ZN(n1262) );
NAND2_X1 U999 ( .A1(n1297), .A2(G234), .ZN(n1264) );
XNOR2_X1 U1000 ( .A(G902), .B(KEYINPUT5), .ZN(n1297) );
XOR2_X1 U1001 ( .A(n1105), .B(G469), .Z(n1068) );
NAND2_X1 U1002 ( .A1(n1298), .A2(n1283), .ZN(n1105) );
XOR2_X1 U1003 ( .A(n1299), .B(n1300), .Z(n1298) );
XOR2_X1 U1004 ( .A(G140), .B(n1301), .Z(n1300) );
NOR2_X1 U1005 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
XOR2_X1 U1006 ( .A(n1304), .B(KEYINPUT10), .Z(n1303) );
NAND2_X1 U1007 ( .A1(n1176), .A2(n1287), .ZN(n1304) );
NOR2_X1 U1008 ( .A1(n1176), .A2(n1287), .ZN(n1302) );
XOR2_X1 U1009 ( .A(G131), .B(n1305), .Z(n1287) );
XOR2_X1 U1010 ( .A(G137), .B(G134), .Z(n1305) );
XOR2_X1 U1011 ( .A(n1306), .B(n1307), .Z(n1176) );
XNOR2_X1 U1012 ( .A(n1124), .B(G101), .ZN(n1307) );
XOR2_X1 U1013 ( .A(n1308), .B(n1309), .Z(n1306) );
NAND2_X1 U1014 ( .A1(KEYINPUT2), .A2(n1310), .ZN(n1308) );
XNOR2_X1 U1015 ( .A(n1311), .B(n1312), .ZN(n1299) );
NOR2_X1 U1016 ( .A1(G110), .A2(KEYINPUT55), .ZN(n1312) );
NOR2_X1 U1017 ( .A1(KEYINPUT14), .A2(n1181), .ZN(n1311) );
NAND2_X1 U1018 ( .A1(G227), .A2(n1075), .ZN(n1181) );
NOR2_X1 U1019 ( .A1(n1090), .A2(n1089), .ZN(n1209) );
INV_X1 U1020 ( .A(n1232), .ZN(n1089) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1313), .ZN(n1232) );
XOR2_X1 U1022 ( .A(KEYINPUT24), .B(n1314), .Z(n1313) );
NOR2_X1 U1023 ( .A1(G237), .A2(G902), .ZN(n1314) );
INV_X1 U1024 ( .A(n1100), .ZN(n1090) );
XOR2_X1 U1025 ( .A(n1315), .B(n1189), .Z(n1100) );
NAND2_X1 U1026 ( .A1(G210), .A2(n1316), .ZN(n1189) );
NAND2_X1 U1027 ( .A1(n1294), .A2(n1283), .ZN(n1316) );
NAND2_X1 U1028 ( .A1(n1317), .A2(n1283), .ZN(n1315) );
XOR2_X1 U1029 ( .A(n1318), .B(n1319), .Z(n1317) );
XNOR2_X1 U1030 ( .A(n1166), .B(n1133), .ZN(n1319) );
XNOR2_X1 U1031 ( .A(n1320), .B(n1321), .ZN(n1133) );
XOR2_X1 U1032 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1033 ( .A(G110), .B(n1310), .ZN(n1323) );
INV_X1 U1034 ( .A(G107), .ZN(n1310) );
XNOR2_X1 U1035 ( .A(G119), .B(n1292), .ZN(n1322) );
XOR2_X1 U1036 ( .A(n1324), .B(n1325), .Z(n1320) );
XNOR2_X1 U1037 ( .A(n1326), .B(n1327), .ZN(n1325) );
NOR2_X1 U1038 ( .A1(KEYINPUT46), .A2(n1328), .ZN(n1327) );
INV_X1 U1039 ( .A(G116), .ZN(n1328) );
NAND2_X1 U1040 ( .A1(KEYINPUT47), .A2(n1329), .ZN(n1326) );
INV_X1 U1041 ( .A(G104), .ZN(n1329) );
XNOR2_X1 U1042 ( .A(n1330), .B(n1237), .ZN(n1324) );
INV_X1 U1043 ( .A(G101), .ZN(n1237) );
NAND2_X1 U1044 ( .A1(KEYINPUT11), .A2(n1331), .ZN(n1330) );
NAND3_X1 U1045 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1166) );
NAND2_X1 U1046 ( .A1(G128), .A2(n1335), .ZN(n1334) );
OR3_X1 U1047 ( .A1(n1335), .A2(G128), .A3(KEYINPUT21), .ZN(n1333) );
OR2_X1 U1048 ( .A1(KEYINPUT45), .A2(n1121), .ZN(n1335) );
NAND2_X1 U1049 ( .A1(KEYINPUT21), .A2(n1121), .ZN(n1332) );
XNOR2_X1 U1050 ( .A(n1188), .B(n1336), .ZN(n1318) );
XNOR2_X1 U1051 ( .A(KEYINPUT8), .B(n1337), .ZN(n1336) );
INV_X1 U1052 ( .A(G125), .ZN(n1337) );
NAND2_X1 U1053 ( .A1(G224), .A2(n1075), .ZN(n1188) );
INV_X1 U1054 ( .A(n1077), .ZN(n1065) );
NOR2_X1 U1055 ( .A1(n1225), .A2(n1104), .ZN(n1077) );
XOR2_X1 U1056 ( .A(n1338), .B(n1156), .Z(n1104) );
INV_X1 U1057 ( .A(G475), .ZN(n1156) );
OR2_X1 U1058 ( .A1(n1155), .A2(G902), .ZN(n1338) );
XNOR2_X1 U1059 ( .A(n1339), .B(n1340), .ZN(n1155) );
XNOR2_X1 U1060 ( .A(n1309), .B(n1341), .ZN(n1340) );
XOR2_X1 U1061 ( .A(n1342), .B(n1343), .Z(n1341) );
NOR2_X1 U1062 ( .A1(G131), .A2(KEYINPUT44), .ZN(n1343) );
NAND2_X1 U1063 ( .A1(n1344), .A2(n1345), .ZN(n1342) );
NAND2_X1 U1064 ( .A1(G113), .A2(n1331), .ZN(n1345) );
INV_X1 U1065 ( .A(G122), .ZN(n1331) );
XOR2_X1 U1066 ( .A(n1346), .B(KEYINPUT6), .Z(n1344) );
NAND2_X1 U1067 ( .A1(G122), .A2(n1292), .ZN(n1346) );
INV_X1 U1068 ( .A(G113), .ZN(n1292) );
XNOR2_X1 U1069 ( .A(G104), .B(n1121), .ZN(n1309) );
XNOR2_X1 U1070 ( .A(G143), .B(G146), .ZN(n1121) );
XOR2_X1 U1071 ( .A(n1347), .B(n1348), .Z(n1339) );
XOR2_X1 U1072 ( .A(KEYINPUT35), .B(KEYINPUT30), .Z(n1348) );
XOR2_X1 U1073 ( .A(n1349), .B(n1350), .Z(n1347) );
AND3_X1 U1074 ( .A1(G214), .A2(n1075), .A3(n1294), .ZN(n1350) );
INV_X1 U1075 ( .A(G237), .ZN(n1294) );
NAND2_X1 U1076 ( .A1(KEYINPUT25), .A2(n1119), .ZN(n1349) );
XNOR2_X1 U1077 ( .A(G125), .B(G140), .ZN(n1119) );
NAND2_X1 U1078 ( .A1(n1351), .A2(n1352), .ZN(n1225) );
NAND2_X1 U1079 ( .A1(n1109), .A2(n1107), .ZN(n1352) );
INV_X1 U1080 ( .A(G478), .ZN(n1107) );
INV_X1 U1081 ( .A(n1353), .ZN(n1109) );
XOR2_X1 U1082 ( .A(n1354), .B(KEYINPUT41), .Z(n1351) );
NAND2_X1 U1083 ( .A1(G478), .A2(n1353), .ZN(n1354) );
NAND2_X1 U1084 ( .A1(n1152), .A2(n1283), .ZN(n1353) );
INV_X1 U1085 ( .A(G902), .ZN(n1283) );
XOR2_X1 U1086 ( .A(n1355), .B(n1356), .Z(n1152) );
XOR2_X1 U1087 ( .A(n1357), .B(n1358), .Z(n1356) );
XNOR2_X1 U1088 ( .A(G134), .B(n1124), .ZN(n1358) );
INV_X1 U1089 ( .A(G128), .ZN(n1124) );
XOR2_X1 U1090 ( .A(KEYINPUT15), .B(G143), .Z(n1357) );
XOR2_X1 U1091 ( .A(n1359), .B(n1360), .Z(n1355) );
XOR2_X1 U1092 ( .A(n1361), .B(n1362), .Z(n1360) );
NAND2_X1 U1093 ( .A1(G217), .A2(n1280), .ZN(n1362) );
AND2_X1 U1094 ( .A1(G234), .A2(n1075), .ZN(n1280) );
INV_X1 U1095 ( .A(G953), .ZN(n1075) );
NAND2_X1 U1096 ( .A1(KEYINPUT61), .A2(G116), .ZN(n1361) );
XNOR2_X1 U1097 ( .A(G107), .B(G122), .ZN(n1359) );
endmodule


