//Key = 1101001110101011000000010101100101000110010001111100100011010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384;

XNOR2_X1 U759 ( .A(n1048), .B(n1049), .ZN(G9) );
NAND2_X1 U760 ( .A1(KEYINPUT6), .A2(G107), .ZN(n1049) );
NAND3_X1 U761 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(G75) );
NAND2_X1 U762 ( .A1(G952), .A2(n1053), .ZN(n1052) );
NAND4_X1 U763 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1053) );
NAND2_X1 U764 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U765 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND3_X1 U766 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
XNOR2_X1 U767 ( .A(n1065), .B(KEYINPUT49), .ZN(n1064) );
NAND2_X1 U768 ( .A1(n1065), .A2(n1066), .ZN(n1060) );
NAND2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1056) );
NAND3_X1 U770 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1068) );
XOR2_X1 U771 ( .A(KEYINPUT14), .B(n1072), .Z(n1071) );
AND2_X1 U772 ( .A1(n1073), .A2(n1058), .ZN(n1072) );
NAND4_X1 U773 ( .A1(n1065), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1070) );
NAND2_X1 U774 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U775 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND4_X1 U776 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1075) );
NAND2_X1 U777 ( .A1(n1085), .A2(n1079), .ZN(n1083) );
NAND3_X1 U778 ( .A1(n1080), .A2(n1086), .A3(n1087), .ZN(n1081) );
NAND2_X1 U779 ( .A1(n1058), .A2(n1088), .ZN(n1069) );
AND4_X1 U780 ( .A1(n1080), .A2(n1079), .A3(n1084), .A4(n1074), .ZN(n1058) );
XNOR2_X1 U781 ( .A(n1089), .B(KEYINPUT25), .ZN(n1074) );
NAND4_X1 U782 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1050) );
NOR4_X1 U783 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1093) );
NOR2_X1 U784 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
NOR2_X1 U785 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
XOR2_X1 U786 ( .A(KEYINPUT21), .B(G475), .Z(n1101) );
XNOR2_X1 U787 ( .A(n1102), .B(n1103), .ZN(n1095) );
NAND4_X1 U788 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1094) );
NAND3_X1 U789 ( .A1(KEYINPUT45), .A2(n1099), .A3(n1108), .ZN(n1107) );
XOR2_X1 U790 ( .A(n1109), .B(KEYINPUT41), .Z(n1099) );
NAND2_X1 U791 ( .A1(G475), .A2(n1100), .ZN(n1106) );
INV_X1 U792 ( .A(KEYINPUT45), .ZN(n1100) );
OR3_X1 U793 ( .A1(n1110), .A2(n1111), .A3(KEYINPUT26), .ZN(n1105) );
NAND2_X1 U794 ( .A1(KEYINPUT26), .A2(n1110), .ZN(n1104) );
NOR3_X1 U795 ( .A1(n1112), .A2(n1063), .A3(n1113), .ZN(n1092) );
XOR2_X1 U796 ( .A(n1114), .B(n1115), .Z(n1091) );
NOR2_X1 U797 ( .A1(n1116), .A2(KEYINPUT4), .ZN(n1115) );
NOR2_X1 U798 ( .A1(n1087), .A2(n1117), .ZN(n1090) );
NOR2_X1 U799 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U800 ( .A1(G902), .A2(n1120), .ZN(n1118) );
XOR2_X1 U801 ( .A(n1121), .B(n1122), .Z(G72) );
XOR2_X1 U802 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U803 ( .A1(G953), .A2(n1125), .ZN(n1124) );
NAND2_X1 U804 ( .A1(G900), .A2(n1126), .ZN(n1125) );
XOR2_X1 U805 ( .A(KEYINPUT16), .B(G227), .Z(n1126) );
NAND2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(n1123) );
NAND2_X1 U807 ( .A1(G953), .A2(n1129), .ZN(n1128) );
XOR2_X1 U808 ( .A(n1130), .B(n1131), .Z(n1127) );
XOR2_X1 U809 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U810 ( .A(n1134), .B(n1135), .Z(n1130) );
XOR2_X1 U811 ( .A(G131), .B(G128), .Z(n1135) );
NAND3_X1 U812 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1134) );
OR2_X1 U813 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NAND3_X1 U814 ( .A1(n1140), .A2(n1139), .A3(KEYINPUT57), .ZN(n1137) );
NOR2_X1 U815 ( .A1(KEYINPUT34), .A2(n1141), .ZN(n1140) );
OR2_X1 U816 ( .A1(n1142), .A2(KEYINPUT57), .ZN(n1136) );
NOR2_X1 U817 ( .A1(n1055), .A2(G953), .ZN(n1121) );
XOR2_X1 U818 ( .A(n1143), .B(n1144), .Z(G69) );
XOR2_X1 U819 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR2_X1 U820 ( .A1(n1147), .A2(n1051), .ZN(n1146) );
AND2_X1 U821 ( .A1(G224), .A2(G898), .ZN(n1147) );
NAND2_X1 U822 ( .A1(n1148), .A2(n1149), .ZN(n1145) );
NAND2_X1 U823 ( .A1(G953), .A2(n1150), .ZN(n1149) );
XOR2_X1 U824 ( .A(n1151), .B(n1152), .Z(n1148) );
NAND2_X1 U825 ( .A1(n1051), .A2(n1153), .ZN(n1143) );
NOR2_X1 U826 ( .A1(n1154), .A2(n1155), .ZN(G66) );
XNOR2_X1 U827 ( .A(n1156), .B(n1157), .ZN(n1155) );
NOR2_X1 U828 ( .A1(n1102), .A2(n1158), .ZN(n1157) );
NOR2_X1 U829 ( .A1(n1154), .A2(n1159), .ZN(G63) );
XOR2_X1 U830 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U831 ( .A1(n1110), .A2(n1158), .ZN(n1160) );
NOR2_X1 U832 ( .A1(n1154), .A2(n1162), .ZN(G60) );
XNOR2_X1 U833 ( .A(n1163), .B(n1164), .ZN(n1162) );
NOR2_X1 U834 ( .A1(n1108), .A2(n1158), .ZN(n1164) );
XOR2_X1 U835 ( .A(G104), .B(n1165), .Z(G6) );
NOR2_X1 U836 ( .A1(n1154), .A2(n1166), .ZN(G57) );
XOR2_X1 U837 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U838 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U839 ( .A1(KEYINPUT24), .A2(n1171), .ZN(n1170) );
NOR2_X1 U840 ( .A1(n1172), .A2(n1158), .ZN(n1169) );
INV_X1 U841 ( .A(G472), .ZN(n1172) );
XOR2_X1 U842 ( .A(n1173), .B(n1174), .Z(n1167) );
NOR2_X1 U843 ( .A1(n1154), .A2(n1175), .ZN(G54) );
XOR2_X1 U844 ( .A(n1176), .B(n1177), .Z(n1175) );
OR2_X1 U845 ( .A1(n1158), .A2(n1119), .ZN(n1177) );
INV_X1 U846 ( .A(G469), .ZN(n1119) );
NAND2_X1 U847 ( .A1(KEYINPUT31), .A2(n1178), .ZN(n1176) );
XOR2_X1 U848 ( .A(n1179), .B(n1180), .Z(n1178) );
XNOR2_X1 U849 ( .A(n1181), .B(n1182), .ZN(n1180) );
NAND3_X1 U850 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1181) );
NAND2_X1 U851 ( .A1(G140), .A2(n1186), .ZN(n1185) );
NAND2_X1 U852 ( .A1(KEYINPUT44), .A2(n1187), .ZN(n1184) );
NAND2_X1 U853 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U854 ( .A(KEYINPUT51), .B(G110), .Z(n1188) );
NAND2_X1 U855 ( .A1(n1190), .A2(n1191), .ZN(n1183) );
INV_X1 U856 ( .A(KEYINPUT44), .ZN(n1191) );
NAND2_X1 U857 ( .A1(n1192), .A2(n1193), .ZN(n1190) );
OR3_X1 U858 ( .A1(n1186), .A2(G140), .A3(KEYINPUT51), .ZN(n1193) );
NAND2_X1 U859 ( .A1(KEYINPUT51), .A2(n1186), .ZN(n1192) );
NOR3_X1 U860 ( .A1(n1154), .A2(n1194), .A3(n1195), .ZN(G51) );
NOR2_X1 U861 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
XOR2_X1 U862 ( .A(n1198), .B(n1199), .Z(n1197) );
AND2_X1 U863 ( .A1(n1200), .A2(KEYINPUT52), .ZN(n1199) );
INV_X1 U864 ( .A(KEYINPUT40), .ZN(n1196) );
NOR2_X1 U865 ( .A1(KEYINPUT40), .A2(n1201), .ZN(n1194) );
XOR2_X1 U866 ( .A(n1198), .B(n1202), .Z(n1201) );
NOR2_X1 U867 ( .A1(n1200), .A2(n1203), .ZN(n1202) );
INV_X1 U868 ( .A(KEYINPUT52), .ZN(n1203) );
XOR2_X1 U869 ( .A(n1204), .B(n1205), .Z(n1198) );
XOR2_X1 U870 ( .A(n1206), .B(n1207), .Z(n1205) );
NOR2_X1 U871 ( .A1(n1208), .A2(n1158), .ZN(n1206) );
NAND2_X1 U872 ( .A1(n1209), .A2(n1210), .ZN(n1158) );
NAND2_X1 U873 ( .A1(n1054), .A2(n1055), .ZN(n1210) );
AND4_X1 U874 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1055) );
NOR4_X1 U875 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
NOR2_X1 U876 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
XOR2_X1 U877 ( .A(KEYINPUT22), .B(n1221), .Z(n1220) );
INV_X1 U878 ( .A(n1222), .ZN(n1215) );
NOR2_X1 U879 ( .A1(n1223), .A2(n1224), .ZN(n1213) );
INV_X1 U880 ( .A(n1153), .ZN(n1054) );
NAND4_X1 U881 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1153) );
NOR4_X1 U882 ( .A1(n1229), .A2(n1230), .A3(n1165), .A4(n1048), .ZN(n1228) );
AND2_X1 U883 ( .A1(n1231), .A2(n1073), .ZN(n1048) );
AND2_X1 U884 ( .A1(n1088), .A2(n1231), .ZN(n1165) );
NOR2_X1 U885 ( .A1(n1232), .A2(n1082), .ZN(n1231) );
NOR2_X1 U886 ( .A1(n1233), .A2(n1234), .ZN(n1227) );
NOR2_X1 U887 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XOR2_X1 U888 ( .A(KEYINPUT12), .B(n1237), .Z(n1236) );
NOR2_X1 U889 ( .A1(n1082), .A2(n1238), .ZN(n1237) );
NAND2_X1 U890 ( .A1(n1239), .A2(n1080), .ZN(n1082) );
INV_X1 U891 ( .A(n1240), .ZN(n1233) );
XOR2_X1 U892 ( .A(KEYINPUT13), .B(G902), .Z(n1209) );
XOR2_X1 U893 ( .A(n1241), .B(n1242), .Z(n1204) );
NAND2_X1 U894 ( .A1(KEYINPUT37), .A2(n1243), .ZN(n1241) );
NOR2_X1 U895 ( .A1(n1051), .A2(G952), .ZN(n1154) );
XOR2_X1 U896 ( .A(G146), .B(n1217), .Z(G48) );
AND3_X1 U897 ( .A1(n1088), .A2(n1066), .A3(n1244), .ZN(n1217) );
XOR2_X1 U898 ( .A(G143), .B(n1216), .Z(G45) );
AND4_X1 U899 ( .A1(n1245), .A2(n1246), .A3(n1247), .A4(n1248), .ZN(n1216) );
NOR2_X1 U900 ( .A1(n1235), .A2(n1249), .ZN(n1248) );
XOR2_X1 U901 ( .A(n1189), .B(n1222), .Z(G42) );
NAND3_X1 U902 ( .A1(n1250), .A2(n1239), .A3(n1067), .ZN(n1222) );
INV_X1 U903 ( .A(G140), .ZN(n1189) );
XOR2_X1 U904 ( .A(n1139), .B(n1211), .Z(G39) );
NAND3_X1 U905 ( .A1(n1244), .A2(n1065), .A3(n1067), .ZN(n1211) );
XOR2_X1 U906 ( .A(n1251), .B(n1252), .Z(G36) );
NOR2_X1 U907 ( .A1(n1221), .A2(n1219), .ZN(n1252) );
NAND3_X1 U908 ( .A1(n1253), .A2(n1073), .A3(n1067), .ZN(n1219) );
INV_X1 U909 ( .A(n1247), .ZN(n1221) );
NOR2_X1 U910 ( .A1(KEYINPUT61), .A2(n1254), .ZN(n1251) );
NAND2_X1 U911 ( .A1(n1255), .A2(n1256), .ZN(G33) );
NAND2_X1 U912 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND2_X1 U913 ( .A1(G131), .A2(n1259), .ZN(n1255) );
NAND2_X1 U914 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
OR2_X1 U915 ( .A1(n1212), .A2(KEYINPUT3), .ZN(n1261) );
NAND2_X1 U916 ( .A1(KEYINPUT3), .A2(n1262), .ZN(n1260) );
INV_X1 U917 ( .A(n1257), .ZN(n1262) );
NOR2_X1 U918 ( .A1(KEYINPUT54), .A2(n1212), .ZN(n1257) );
NAND4_X1 U919 ( .A1(n1067), .A2(n1253), .A3(n1088), .A4(n1247), .ZN(n1212) );
AND2_X1 U920 ( .A1(n1062), .A2(n1263), .ZN(n1067) );
XOR2_X1 U921 ( .A(G128), .B(n1224), .Z(G30) );
AND3_X1 U922 ( .A1(n1073), .A2(n1066), .A3(n1244), .ZN(n1224) );
AND4_X1 U923 ( .A1(n1085), .A2(n1239), .A3(n1077), .A4(n1247), .ZN(n1244) );
XOR2_X1 U924 ( .A(n1264), .B(n1240), .Z(G3) );
NAND4_X1 U925 ( .A1(n1253), .A2(n1065), .A3(n1066), .A4(n1265), .ZN(n1240) );
INV_X1 U926 ( .A(n1249), .ZN(n1253) );
NAND3_X1 U927 ( .A1(n1084), .A2(n1239), .A3(n1085), .ZN(n1249) );
XOR2_X1 U928 ( .A(G125), .B(n1223), .Z(G27) );
AND3_X1 U929 ( .A1(n1079), .A2(n1066), .A3(n1250), .ZN(n1223) );
AND4_X1 U930 ( .A1(n1080), .A2(n1088), .A3(n1077), .A4(n1247), .ZN(n1250) );
NAND2_X1 U931 ( .A1(n1266), .A2(n1267), .ZN(n1247) );
NAND2_X1 U932 ( .A1(n1268), .A2(n1129), .ZN(n1267) );
INV_X1 U933 ( .A(G900), .ZN(n1129) );
INV_X1 U934 ( .A(n1269), .ZN(n1079) );
XNOR2_X1 U935 ( .A(G122), .B(n1225), .ZN(G24) );
NAND4_X1 U936 ( .A1(n1080), .A2(n1270), .A3(n1245), .A4(n1246), .ZN(n1225) );
XOR2_X1 U937 ( .A(n1230), .B(n1271), .Z(G21) );
NOR2_X1 U938 ( .A1(KEYINPUT43), .A2(n1272), .ZN(n1271) );
NOR4_X1 U939 ( .A1(n1273), .A2(n1238), .A3(n1269), .A4(n1235), .ZN(n1230) );
INV_X1 U940 ( .A(n1085), .ZN(n1273) );
XNOR2_X1 U941 ( .A(n1229), .B(n1274), .ZN(G18) );
XOR2_X1 U942 ( .A(KEYINPUT33), .B(G116), .Z(n1274) );
AND3_X1 U943 ( .A1(n1085), .A2(n1073), .A3(n1270), .ZN(n1229) );
NOR2_X1 U944 ( .A1(n1245), .A2(n1275), .ZN(n1073) );
NAND2_X1 U945 ( .A1(n1276), .A2(n1277), .ZN(G15) );
OR2_X1 U946 ( .A1(n1226), .A2(G113), .ZN(n1277) );
XOR2_X1 U947 ( .A(n1278), .B(KEYINPUT32), .Z(n1276) );
NAND2_X1 U948 ( .A1(G113), .A2(n1226), .ZN(n1278) );
NAND3_X1 U949 ( .A1(n1085), .A2(n1270), .A3(n1088), .ZN(n1226) );
AND2_X1 U950 ( .A1(n1275), .A2(n1245), .ZN(n1088) );
NOR2_X1 U951 ( .A1(n1269), .A2(n1232), .ZN(n1270) );
NAND3_X1 U952 ( .A1(n1084), .A2(n1265), .A3(n1066), .ZN(n1232) );
NAND2_X1 U953 ( .A1(n1086), .A2(n1279), .ZN(n1269) );
XOR2_X1 U954 ( .A(n1080), .B(KEYINPUT56), .Z(n1085) );
XOR2_X1 U955 ( .A(G110), .B(n1280), .Z(G12) );
NOR4_X1 U956 ( .A1(n1281), .A2(n1282), .A3(n1238), .A4(n1097), .ZN(n1280) );
INV_X1 U957 ( .A(n1080), .ZN(n1097) );
XOR2_X1 U958 ( .A(n1283), .B(G472), .Z(n1080) );
NAND2_X1 U959 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XNOR2_X1 U960 ( .A(n1171), .B(n1286), .ZN(n1284) );
XOR2_X1 U961 ( .A(n1287), .B(n1173), .Z(n1286) );
XOR2_X1 U962 ( .A(n1288), .B(n1289), .Z(n1173) );
XOR2_X1 U963 ( .A(G119), .B(G116), .Z(n1289) );
XNOR2_X1 U964 ( .A(n1207), .B(G113), .ZN(n1288) );
NAND2_X1 U965 ( .A1(n1290), .A2(KEYINPUT0), .ZN(n1287) );
XNOR2_X1 U966 ( .A(n1174), .B(KEYINPUT63), .ZN(n1290) );
XNOR2_X1 U967 ( .A(n1291), .B(G101), .ZN(n1174) );
NAND3_X1 U968 ( .A1(G210), .A2(n1051), .A3(n1292), .ZN(n1291) );
NAND3_X1 U969 ( .A1(n1077), .A2(n1265), .A3(n1065), .ZN(n1238) );
NOR2_X1 U970 ( .A1(n1246), .A2(n1245), .ZN(n1065) );
NAND3_X1 U971 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(n1245) );
NAND2_X1 U972 ( .A1(KEYINPUT36), .A2(n1296), .ZN(n1295) );
NAND2_X1 U973 ( .A1(n1109), .A2(n1297), .ZN(n1296) );
NAND2_X1 U974 ( .A1(G475), .A2(n1298), .ZN(n1297) );
NAND4_X1 U975 ( .A1(n1109), .A2(n1299), .A3(KEYINPUT62), .A4(G475), .ZN(n1294) );
NAND2_X1 U976 ( .A1(n1300), .A2(n1108), .ZN(n1293) );
INV_X1 U977 ( .A(G475), .ZN(n1108) );
NAND3_X1 U978 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1300) );
NAND2_X1 U979 ( .A1(KEYINPUT62), .A2(KEYINPUT36), .ZN(n1303) );
NAND2_X1 U980 ( .A1(KEYINPUT35), .A2(n1109), .ZN(n1302) );
NAND2_X1 U981 ( .A1(n1304), .A2(n1305), .ZN(n1301) );
INV_X1 U982 ( .A(KEYINPUT35), .ZN(n1305) );
NAND2_X1 U983 ( .A1(n1109), .A2(n1306), .ZN(n1304) );
NAND2_X1 U984 ( .A1(n1299), .A2(n1298), .ZN(n1306) );
INV_X1 U985 ( .A(KEYINPUT62), .ZN(n1298) );
INV_X1 U986 ( .A(KEYINPUT36), .ZN(n1299) );
NAND2_X1 U987 ( .A1(n1163), .A2(n1285), .ZN(n1109) );
XNOR2_X1 U988 ( .A(n1307), .B(n1308), .ZN(n1163) );
XOR2_X1 U989 ( .A(G104), .B(n1309), .Z(n1308) );
XOR2_X1 U990 ( .A(G131), .B(G113), .Z(n1309) );
XOR2_X1 U991 ( .A(n1310), .B(n1311), .Z(n1307) );
XOR2_X1 U992 ( .A(n1312), .B(n1313), .Z(n1310) );
NAND2_X1 U993 ( .A1(n1314), .A2(n1315), .ZN(n1312) );
NAND4_X1 U994 ( .A1(n1292), .A2(G214), .A3(G143), .A4(n1051), .ZN(n1315) );
XOR2_X1 U995 ( .A(n1316), .B(KEYINPUT50), .Z(n1314) );
NAND2_X1 U996 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND3_X1 U997 ( .A1(G214), .A2(n1051), .A3(n1292), .ZN(n1318) );
XOR2_X1 U998 ( .A(n1319), .B(KEYINPUT18), .Z(n1292) );
INV_X1 U999 ( .A(n1275), .ZN(n1246) );
NOR2_X1 U1000 ( .A1(n1112), .A2(n1320), .ZN(n1275) );
NOR2_X1 U1001 ( .A1(n1110), .A2(n1111), .ZN(n1320) );
AND2_X1 U1002 ( .A1(n1111), .A2(n1110), .ZN(n1112) );
INV_X1 U1003 ( .A(G478), .ZN(n1110) );
NOR2_X1 U1004 ( .A1(n1161), .A2(G902), .ZN(n1111) );
XNOR2_X1 U1005 ( .A(n1321), .B(n1322), .ZN(n1161) );
XOR2_X1 U1006 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1007 ( .A(G116), .B(n1317), .Z(n1324) );
NAND3_X1 U1008 ( .A1(G234), .A2(n1051), .A3(G217), .ZN(n1323) );
XNOR2_X1 U1009 ( .A(n1325), .B(n1326), .ZN(n1321) );
XOR2_X1 U1010 ( .A(n1142), .B(n1313), .Z(n1326) );
NAND2_X1 U1011 ( .A1(n1266), .A2(n1327), .ZN(n1265) );
NAND2_X1 U1012 ( .A1(n1268), .A2(n1150), .ZN(n1327) );
INV_X1 U1013 ( .A(G898), .ZN(n1150) );
AND3_X1 U1014 ( .A1(G902), .A2(n1089), .A3(G953), .ZN(n1268) );
NAND3_X1 U1015 ( .A1(n1089), .A2(n1051), .A3(G952), .ZN(n1266) );
NAND2_X1 U1016 ( .A1(G237), .A2(G234), .ZN(n1089) );
INV_X1 U1017 ( .A(n1084), .ZN(n1077) );
XNOR2_X1 U1018 ( .A(n1328), .B(n1102), .ZN(n1084) );
NAND2_X1 U1019 ( .A1(G217), .A2(n1329), .ZN(n1102) );
NAND2_X1 U1020 ( .A1(KEYINPUT10), .A2(n1103), .ZN(n1328) );
AND2_X1 U1021 ( .A1(n1285), .A2(n1156), .ZN(n1103) );
NAND2_X1 U1022 ( .A1(n1330), .A2(n1331), .ZN(n1156) );
NAND2_X1 U1023 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
XOR2_X1 U1024 ( .A(KEYINPUT28), .B(n1334), .Z(n1330) );
NOR2_X1 U1025 ( .A1(n1333), .A2(n1332), .ZN(n1334) );
XOR2_X1 U1026 ( .A(n1335), .B(n1336), .Z(n1332) );
OR2_X1 U1027 ( .A1(KEYINPUT29), .A2(n1139), .ZN(n1336) );
INV_X1 U1028 ( .A(G137), .ZN(n1139) );
NAND3_X1 U1029 ( .A1(G234), .A2(n1051), .A3(G221), .ZN(n1335) );
XOR2_X1 U1030 ( .A(n1311), .B(n1337), .Z(n1333) );
XOR2_X1 U1031 ( .A(G110), .B(n1338), .Z(n1337) );
NOR2_X1 U1032 ( .A1(KEYINPUT5), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1033 ( .A(G119), .B(n1340), .Z(n1339) );
XOR2_X1 U1034 ( .A(KEYINPUT9), .B(G128), .Z(n1340) );
XOR2_X1 U1035 ( .A(G146), .B(n1132), .Z(n1311) );
XOR2_X1 U1036 ( .A(G125), .B(G140), .Z(n1132) );
XNOR2_X1 U1037 ( .A(n1239), .B(KEYINPUT11), .ZN(n1282) );
NOR2_X1 U1038 ( .A1(n1087), .A2(n1086), .ZN(n1239) );
NOR2_X1 U1039 ( .A1(n1341), .A2(n1113), .ZN(n1086) );
NOR3_X1 U1040 ( .A1(G469), .A2(G902), .A3(n1120), .ZN(n1113) );
AND2_X1 U1041 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
OR2_X1 U1042 ( .A1(n1120), .A2(G902), .ZN(n1343) );
XOR2_X1 U1043 ( .A(n1344), .B(n1345), .Z(n1120) );
XOR2_X1 U1044 ( .A(G140), .B(G110), .Z(n1345) );
XOR2_X1 U1045 ( .A(n1179), .B(n1346), .Z(n1344) );
NOR2_X1 U1046 ( .A1(KEYINPUT60), .A2(n1182), .ZN(n1346) );
NAND2_X1 U1047 ( .A1(G227), .A2(n1051), .ZN(n1182) );
XOR2_X1 U1048 ( .A(n1347), .B(n1348), .Z(n1179) );
XOR2_X1 U1049 ( .A(G101), .B(n1349), .Z(n1348) );
XOR2_X1 U1050 ( .A(KEYINPUT23), .B(G104), .Z(n1349) );
XOR2_X1 U1051 ( .A(n1171), .B(n1350), .Z(n1347) );
XOR2_X1 U1052 ( .A(n1325), .B(n1133), .Z(n1350) );
XOR2_X1 U1053 ( .A(G107), .B(G128), .Z(n1325) );
XOR2_X1 U1054 ( .A(n1351), .B(n1352), .Z(n1171) );
XOR2_X1 U1055 ( .A(KEYINPUT58), .B(G137), .Z(n1352) );
XOR2_X1 U1056 ( .A(n1258), .B(n1142), .Z(n1351) );
INV_X1 U1057 ( .A(n1141), .ZN(n1142) );
XOR2_X1 U1058 ( .A(n1254), .B(KEYINPUT15), .Z(n1141) );
INV_X1 U1059 ( .A(G134), .ZN(n1254) );
INV_X1 U1060 ( .A(G131), .ZN(n1258) );
XOR2_X1 U1061 ( .A(KEYINPUT17), .B(G469), .Z(n1342) );
INV_X1 U1062 ( .A(n1279), .ZN(n1087) );
NAND2_X1 U1063 ( .A1(G221), .A2(n1329), .ZN(n1279) );
NAND2_X1 U1064 ( .A1(G234), .A2(n1285), .ZN(n1329) );
XOR2_X1 U1065 ( .A(n1235), .B(KEYINPUT30), .Z(n1281) );
INV_X1 U1066 ( .A(n1066), .ZN(n1235) );
NOR2_X1 U1067 ( .A1(n1353), .A2(n1062), .ZN(n1066) );
XOR2_X1 U1068 ( .A(n1354), .B(n1355), .Z(n1062) );
XOR2_X1 U1069 ( .A(KEYINPUT55), .B(n1116), .Z(n1355) );
AND2_X1 U1070 ( .A1(n1356), .A2(n1285), .ZN(n1116) );
XOR2_X1 U1071 ( .A(n1357), .B(n1358), .Z(n1356) );
XOR2_X1 U1072 ( .A(KEYINPUT53), .B(KEYINPUT27), .Z(n1358) );
XNOR2_X1 U1073 ( .A(n1200), .B(n1359), .ZN(n1357) );
NOR2_X1 U1074 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NOR2_X1 U1075 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
XOR2_X1 U1076 ( .A(n1364), .B(n1243), .Z(n1363) );
XOR2_X1 U1077 ( .A(n1365), .B(KEYINPUT2), .Z(n1362) );
NOR2_X1 U1078 ( .A1(n1366), .A2(n1367), .ZN(n1360) );
XOR2_X1 U1079 ( .A(KEYINPUT39), .B(n1242), .Z(n1367) );
INV_X1 U1080 ( .A(n1365), .ZN(n1242) );
NAND2_X1 U1081 ( .A1(G224), .A2(n1051), .ZN(n1365) );
INV_X1 U1082 ( .A(G953), .ZN(n1051) );
XOR2_X1 U1083 ( .A(n1364), .B(n1368), .Z(n1366) );
INV_X1 U1084 ( .A(n1243), .ZN(n1368) );
XOR2_X1 U1085 ( .A(n1369), .B(KEYINPUT42), .Z(n1243) );
INV_X1 U1086 ( .A(G125), .ZN(n1369) );
NAND2_X1 U1087 ( .A1(KEYINPUT47), .A2(n1207), .ZN(n1364) );
XNOR2_X1 U1088 ( .A(n1370), .B(n1133), .ZN(n1207) );
XNOR2_X1 U1089 ( .A(G146), .B(n1317), .ZN(n1133) );
INV_X1 U1090 ( .A(G143), .ZN(n1317) );
NAND2_X1 U1091 ( .A1(KEYINPUT7), .A2(n1371), .ZN(n1370) );
INV_X1 U1092 ( .A(G128), .ZN(n1371) );
XNOR2_X1 U1093 ( .A(n1372), .B(n1373), .ZN(n1200) );
INV_X1 U1094 ( .A(n1151), .ZN(n1373) );
XOR2_X1 U1095 ( .A(n1374), .B(n1375), .Z(n1151) );
XOR2_X1 U1096 ( .A(n1376), .B(n1377), .Z(n1375) );
NAND2_X1 U1097 ( .A1(KEYINPUT1), .A2(n1272), .ZN(n1377) );
INV_X1 U1098 ( .A(G119), .ZN(n1272) );
NAND2_X1 U1099 ( .A1(n1378), .A2(n1379), .ZN(n1376) );
NAND2_X1 U1100 ( .A1(n1380), .A2(n1264), .ZN(n1379) );
XOR2_X1 U1101 ( .A(n1381), .B(KEYINPUT19), .Z(n1378) );
OR2_X1 U1102 ( .A1(n1264), .A2(n1380), .ZN(n1381) );
XNOR2_X1 U1103 ( .A(n1382), .B(G107), .ZN(n1380) );
NAND2_X1 U1104 ( .A1(KEYINPUT59), .A2(n1383), .ZN(n1382) );
INV_X1 U1105 ( .A(G104), .ZN(n1383) );
INV_X1 U1106 ( .A(G101), .ZN(n1264) );
XNOR2_X1 U1107 ( .A(G113), .B(G116), .ZN(n1374) );
NAND2_X1 U1108 ( .A1(KEYINPUT38), .A2(n1152), .ZN(n1372) );
XOR2_X1 U1109 ( .A(n1186), .B(n1313), .Z(n1152) );
XOR2_X1 U1110 ( .A(G122), .B(KEYINPUT20), .Z(n1313) );
INV_X1 U1111 ( .A(G110), .ZN(n1186) );
NAND2_X1 U1112 ( .A1(KEYINPUT46), .A2(n1114), .ZN(n1354) );
INV_X1 U1113 ( .A(n1208), .ZN(n1114) );
NAND2_X1 U1114 ( .A1(G210), .A2(n1384), .ZN(n1208) );
XOR2_X1 U1115 ( .A(n1263), .B(KEYINPUT48), .Z(n1353) );
XOR2_X1 U1116 ( .A(n1063), .B(KEYINPUT8), .Z(n1263) );
AND2_X1 U1117 ( .A1(G214), .A2(n1384), .ZN(n1063) );
NAND2_X1 U1118 ( .A1(n1319), .A2(n1285), .ZN(n1384) );
INV_X1 U1119 ( .A(G902), .ZN(n1285) );
INV_X1 U1120 ( .A(G237), .ZN(n1319) );
endmodule


