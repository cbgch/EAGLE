//Key = 0111001001011000100010101110011000001011001110100101111100111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307;

NAND2_X1 U710 ( .A1(n992), .A2(n993), .ZN(G9) );
NAND2_X1 U711 ( .A1(G107), .A2(n994), .ZN(n993) );
NAND2_X1 U712 ( .A1(n995), .A2(n996), .ZN(n992) );
XOR2_X1 U713 ( .A(KEYINPUT3), .B(G107), .Z(n996) );
XOR2_X1 U714 ( .A(n994), .B(KEYINPUT16), .Z(n995) );
NAND2_X1 U715 ( .A1(n997), .A2(n998), .ZN(n994) );
XNOR2_X1 U716 ( .A(KEYINPUT35), .B(n999), .ZN(n998) );
NAND4_X1 U717 ( .A1(n1000), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(G75) );
NAND2_X1 U718 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NAND2_X1 U719 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NAND2_X1 U720 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND2_X1 U721 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND4_X1 U722 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1011) );
NAND2_X1 U723 ( .A1(n1016), .A2(n1017), .ZN(n1010) );
NAND2_X1 U724 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND2_X1 U725 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U726 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U727 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND2_X1 U728 ( .A1(n1013), .A2(n1026), .ZN(n1018) );
NAND2_X1 U729 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U730 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
INV_X1 U731 ( .A(n1031), .ZN(n1008) );
NAND4_X1 U732 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1006) );
NOR4_X1 U733 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
XOR2_X1 U734 ( .A(n1040), .B(n1041), .Z(n1039) );
NOR2_X1 U735 ( .A1(KEYINPUT5), .A2(n1013), .ZN(n1037) );
AND2_X1 U736 ( .A1(n1022), .A2(KEYINPUT5), .ZN(n1036) );
INV_X1 U737 ( .A(n1042), .ZN(n1022) );
NAND2_X1 U738 ( .A1(G475), .A2(n1043), .ZN(n1034) );
NOR2_X1 U739 ( .A1(G953), .A2(n1044), .ZN(n1002) );
NOR4_X1 U740 ( .A1(n1045), .A2(n1046), .A3(n1014), .A4(n1031), .ZN(n1044) );
INV_X1 U741 ( .A(n1013), .ZN(n1046) );
NOR2_X1 U742 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR3_X1 U743 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
NOR3_X1 U744 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1051) );
NOR2_X1 U745 ( .A1(n1055), .A2(n1015), .ZN(n1054) );
INV_X1 U746 ( .A(KEYINPUT52), .ZN(n1015) );
NOR2_X1 U747 ( .A1(n1056), .A2(n1057), .ZN(n1050) );
AND2_X1 U748 ( .A1(n1016), .A2(KEYINPUT1), .ZN(n1056) );
NOR2_X1 U749 ( .A1(n1058), .A2(n1059), .ZN(n1047) );
INV_X1 U750 ( .A(n1016), .ZN(n1059) );
NOR2_X1 U751 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U752 ( .A1(KEYINPUT1), .A2(n1062), .ZN(n1060) );
XOR2_X1 U753 ( .A(n1063), .B(n1064), .Z(G72) );
XOR2_X1 U754 ( .A(n1065), .B(n1066), .Z(n1064) );
NOR2_X1 U755 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
AND2_X1 U756 ( .A1(G227), .A2(G900), .ZN(n1067) );
NAND2_X1 U757 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
NAND2_X1 U758 ( .A1(G953), .A2(n1071), .ZN(n1070) );
XOR2_X1 U759 ( .A(n1072), .B(n1073), .Z(n1069) );
XNOR2_X1 U760 ( .A(n1074), .B(n1075), .ZN(n1073) );
NAND2_X1 U761 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NAND2_X1 U762 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XOR2_X1 U763 ( .A(n1080), .B(n1081), .Z(n1079) );
XOR2_X1 U764 ( .A(KEYINPUT44), .B(n1082), .Z(n1078) );
XOR2_X1 U765 ( .A(n1083), .B(KEYINPUT47), .Z(n1076) );
NAND2_X1 U766 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XOR2_X1 U767 ( .A(G137), .B(n1081), .Z(n1085) );
XOR2_X1 U768 ( .A(KEYINPUT44), .B(G131), .Z(n1084) );
NAND2_X1 U769 ( .A1(n1068), .A2(n1086), .ZN(n1063) );
XOR2_X1 U770 ( .A(n1087), .B(n1088), .Z(G69) );
NOR2_X1 U771 ( .A1(n1089), .A2(n1068), .ZN(n1088) );
NOR2_X1 U772 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U773 ( .A1(n1092), .A2(n1093), .ZN(n1087) );
NAND2_X1 U774 ( .A1(n1094), .A2(n1068), .ZN(n1093) );
XOR2_X1 U775 ( .A(n1095), .B(n1000), .Z(n1094) );
NAND3_X1 U776 ( .A1(G898), .A2(n1096), .A3(G953), .ZN(n1092) );
INV_X1 U777 ( .A(n1095), .ZN(n1096) );
NOR2_X1 U778 ( .A1(n1097), .A2(n1098), .ZN(G66) );
XOR2_X1 U779 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U780 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR2_X1 U781 ( .A1(n1097), .A2(n1103), .ZN(G63) );
XOR2_X1 U782 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR3_X1 U783 ( .A1(n1102), .A2(KEYINPUT7), .A3(n1106), .ZN(n1105) );
NOR2_X1 U784 ( .A1(n1097), .A2(n1107), .ZN(G60) );
XOR2_X1 U785 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U786 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
AND2_X1 U787 ( .A1(KEYINPUT17), .A2(n1112), .ZN(n1111) );
NOR2_X1 U788 ( .A1(KEYINPUT41), .A2(n1112), .ZN(n1110) );
NAND2_X1 U789 ( .A1(n1113), .A2(G475), .ZN(n1112) );
XOR2_X1 U790 ( .A(n1114), .B(n1115), .Z(G6) );
NOR2_X1 U791 ( .A1(n1097), .A2(n1116), .ZN(G57) );
XOR2_X1 U792 ( .A(n1117), .B(n1118), .Z(n1116) );
XNOR2_X1 U793 ( .A(n1119), .B(n1120), .ZN(n1118) );
NOR2_X1 U794 ( .A1(KEYINPUT34), .A2(n1121), .ZN(n1119) );
NOR2_X1 U795 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XOR2_X1 U796 ( .A(n1124), .B(KEYINPUT30), .Z(n1123) );
NAND2_X1 U797 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR2_X1 U798 ( .A1(n1125), .A2(n1126), .ZN(n1122) );
XNOR2_X1 U799 ( .A(n1127), .B(n1128), .ZN(n1126) );
XOR2_X1 U800 ( .A(n1129), .B(n1130), .Z(n1128) );
AND2_X1 U801 ( .A1(n1113), .A2(G472), .ZN(n1125) );
XOR2_X1 U802 ( .A(n1131), .B(KEYINPUT26), .Z(n1117) );
NOR2_X1 U803 ( .A1(n1097), .A2(n1132), .ZN(G54) );
XOR2_X1 U804 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U805 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U806 ( .A(n1137), .B(n1138), .Z(n1135) );
NOR2_X1 U807 ( .A1(KEYINPUT28), .A2(n1139), .ZN(n1138) );
XOR2_X1 U808 ( .A(n1140), .B(n1141), .Z(n1133) );
XOR2_X1 U809 ( .A(KEYINPUT10), .B(n1142), .Z(n1141) );
AND2_X1 U810 ( .A1(G469), .A2(n1113), .ZN(n1142) );
INV_X1 U811 ( .A(n1102), .ZN(n1113) );
NAND2_X1 U812 ( .A1(KEYINPUT54), .A2(n1143), .ZN(n1140) );
NOR2_X1 U813 ( .A1(n1097), .A2(n1144), .ZN(G51) );
XOR2_X1 U814 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U815 ( .A(n1095), .B(n1147), .Z(n1146) );
XOR2_X1 U816 ( .A(n1148), .B(n1149), .Z(n1145) );
XOR2_X1 U817 ( .A(KEYINPUT38), .B(n1150), .Z(n1149) );
NOR2_X1 U818 ( .A1(n1041), .A2(n1102), .ZN(n1148) );
NAND2_X1 U819 ( .A1(n1151), .A2(n1152), .ZN(n1102) );
NAND2_X1 U820 ( .A1(n1000), .A2(n1001), .ZN(n1152) );
INV_X1 U821 ( .A(n1086), .ZN(n1001) );
NAND4_X1 U822 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1086) );
NOR4_X1 U823 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1156) );
AND2_X1 U824 ( .A1(n1161), .A2(n1162), .ZN(n1155) );
AND2_X1 U825 ( .A1(n1163), .A2(n1164), .ZN(n1000) );
AND4_X1 U826 ( .A1(n1165), .A2(n1115), .A3(n1166), .A4(n1167), .ZN(n1164) );
NAND4_X1 U827 ( .A1(n1013), .A2(n1168), .A3(n1061), .A4(n1169), .ZN(n1115) );
NOR2_X1 U828 ( .A1(n1027), .A2(n1055), .ZN(n1169) );
AND4_X1 U829 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1163) );
OR2_X1 U830 ( .A1(n999), .A2(n1027), .ZN(n1173) );
INV_X1 U831 ( .A(n997), .ZN(n1027) );
NAND4_X1 U832 ( .A1(n1061), .A2(n1053), .A3(n1013), .A4(n1168), .ZN(n999) );
XOR2_X1 U833 ( .A(KEYINPUT31), .B(G902), .Z(n1151) );
NOR2_X1 U834 ( .A1(n1068), .A2(G952), .ZN(n1097) );
NAND2_X1 U835 ( .A1(n1174), .A2(n1175), .ZN(G48) );
NAND2_X1 U836 ( .A1(G146), .A2(n1153), .ZN(n1175) );
XOR2_X1 U837 ( .A(n1176), .B(KEYINPUT45), .Z(n1174) );
OR2_X1 U838 ( .A1(n1153), .A2(G146), .ZN(n1176) );
NAND3_X1 U839 ( .A1(n1012), .A2(n997), .A3(n1177), .ZN(n1153) );
XOR2_X1 U840 ( .A(n1178), .B(n1154), .Z(G45) );
NAND4_X1 U841 ( .A1(n1179), .A2(n997), .A3(n1038), .A4(n1180), .ZN(n1154) );
XNOR2_X1 U842 ( .A(n1160), .B(n1181), .ZN(G42) );
NAND2_X1 U843 ( .A1(KEYINPUT49), .A2(G140), .ZN(n1181) );
AND3_X1 U844 ( .A1(n1182), .A2(n1061), .A3(n1020), .ZN(n1160) );
XOR2_X1 U845 ( .A(G137), .B(n1159), .Z(G39) );
AND3_X1 U846 ( .A1(n1177), .A2(n1016), .A3(n1020), .ZN(n1159) );
NAND2_X1 U847 ( .A1(n1183), .A2(n1184), .ZN(G36) );
NAND2_X1 U848 ( .A1(G134), .A2(n1162), .ZN(n1184) );
XOR2_X1 U849 ( .A(n1185), .B(KEYINPUT23), .Z(n1183) );
OR2_X1 U850 ( .A1(n1162), .A2(G134), .ZN(n1185) );
NAND3_X1 U851 ( .A1(n1020), .A2(n1053), .A3(n1179), .ZN(n1162) );
XOR2_X1 U852 ( .A(n1082), .B(n1161), .Z(G33) );
NAND3_X1 U853 ( .A1(n1020), .A2(n1012), .A3(n1179), .ZN(n1161) );
AND3_X1 U854 ( .A1(n1061), .A2(n1186), .A3(n1042), .ZN(n1179) );
INV_X1 U855 ( .A(n1014), .ZN(n1020) );
NAND2_X1 U856 ( .A1(n1030), .A2(n1032), .ZN(n1014) );
XOR2_X1 U857 ( .A(G128), .B(n1158), .Z(G30) );
AND3_X1 U858 ( .A1(n997), .A2(n1053), .A3(n1177), .ZN(n1158) );
AND4_X1 U859 ( .A1(n1061), .A2(n1025), .A3(n1187), .A4(n1186), .ZN(n1177) );
XOR2_X1 U860 ( .A(n1131), .B(n1172), .Z(G3) );
NAND2_X1 U861 ( .A1(n1042), .A2(n1188), .ZN(n1172) );
XOR2_X1 U862 ( .A(G125), .B(n1157), .Z(G27) );
AND3_X1 U863 ( .A1(n1004), .A2(n997), .A3(n1182), .ZN(n1157) );
AND4_X1 U864 ( .A1(n1024), .A2(n1012), .A3(n1025), .A4(n1186), .ZN(n1182) );
NAND2_X1 U865 ( .A1(n1031), .A2(n1189), .ZN(n1186) );
NAND4_X1 U866 ( .A1(G953), .A2(G902), .A3(n1190), .A4(n1071), .ZN(n1189) );
INV_X1 U867 ( .A(G900), .ZN(n1071) );
XNOR2_X1 U868 ( .A(n1165), .B(n1191), .ZN(G24) );
NOR2_X1 U869 ( .A1(KEYINPUT56), .A2(n1192), .ZN(n1191) );
INV_X1 U870 ( .A(G122), .ZN(n1192) );
NAND4_X1 U871 ( .A1(n1193), .A2(n1013), .A3(n1038), .A4(n1180), .ZN(n1165) );
NOR2_X1 U872 ( .A1(n1187), .A2(n1025), .ZN(n1013) );
XOR2_X1 U873 ( .A(n1194), .B(n1171), .Z(G21) );
NAND4_X1 U874 ( .A1(n1016), .A2(n1193), .A3(n1025), .A4(n1187), .ZN(n1171) );
INV_X1 U875 ( .A(n1024), .ZN(n1187) );
XNOR2_X1 U876 ( .A(G116), .B(n1170), .ZN(G18) );
NAND3_X1 U877 ( .A1(n1193), .A2(n1053), .A3(n1042), .ZN(n1170) );
NOR2_X1 U878 ( .A1(n1180), .A2(n1195), .ZN(n1053) );
XNOR2_X1 U879 ( .A(G113), .B(n1167), .ZN(G15) );
NAND3_X1 U880 ( .A1(n1012), .A2(n1193), .A3(n1042), .ZN(n1167) );
NOR2_X1 U881 ( .A1(n1025), .A2(n1024), .ZN(n1042) );
AND3_X1 U882 ( .A1(n997), .A2(n1168), .A3(n1004), .ZN(n1193) );
NOR2_X1 U883 ( .A1(n1049), .A2(n1052), .ZN(n1004) );
INV_X1 U884 ( .A(n1062), .ZN(n1049) );
INV_X1 U885 ( .A(n1055), .ZN(n1012) );
NAND2_X1 U886 ( .A1(n1196), .A2(n1180), .ZN(n1055) );
XOR2_X1 U887 ( .A(n1195), .B(KEYINPUT32), .Z(n1196) );
XOR2_X1 U888 ( .A(n1166), .B(n1197), .Z(G12) );
NOR2_X1 U889 ( .A1(G110), .A2(KEYINPUT48), .ZN(n1197) );
NAND3_X1 U890 ( .A1(n1024), .A2(n1025), .A3(n1188), .ZN(n1166) );
AND4_X1 U891 ( .A1(n1016), .A2(n997), .A3(n1061), .A4(n1168), .ZN(n1188) );
NAND2_X1 U892 ( .A1(n1031), .A2(n1198), .ZN(n1168) );
NAND4_X1 U893 ( .A1(G953), .A2(G902), .A3(n1190), .A4(n1091), .ZN(n1198) );
INV_X1 U894 ( .A(G898), .ZN(n1091) );
NAND3_X1 U895 ( .A1(n1190), .A2(n1068), .A3(G952), .ZN(n1031) );
NAND2_X1 U896 ( .A1(G237), .A2(G234), .ZN(n1190) );
NOR2_X1 U897 ( .A1(n1062), .A2(n1052), .ZN(n1061) );
INV_X1 U898 ( .A(n1057), .ZN(n1052) );
NAND2_X1 U899 ( .A1(G221), .A2(n1199), .ZN(n1057) );
XOR2_X1 U900 ( .A(n1200), .B(G469), .Z(n1062) );
NAND2_X1 U901 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
XOR2_X1 U902 ( .A(n1203), .B(n1204), .Z(n1201) );
XOR2_X1 U903 ( .A(n1137), .B(n1205), .Z(n1203) );
NOR2_X1 U904 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
XOR2_X1 U905 ( .A(KEYINPUT57), .B(n1208), .Z(n1207) );
NOR2_X1 U906 ( .A1(n1209), .A2(n1139), .ZN(n1208) );
AND2_X1 U907 ( .A1(n1139), .A2(n1209), .ZN(n1206) );
XOR2_X1 U908 ( .A(n1210), .B(n1143), .Z(n1209) );
INV_X1 U909 ( .A(G140), .ZN(n1143) );
INV_X1 U910 ( .A(G110), .ZN(n1210) );
NAND2_X1 U911 ( .A1(G227), .A2(n1068), .ZN(n1139) );
XOR2_X1 U912 ( .A(n1211), .B(n1072), .Z(n1137) );
XNOR2_X1 U913 ( .A(n1212), .B(n1213), .ZN(n1072) );
XOR2_X1 U914 ( .A(n1214), .B(G143), .Z(n1212) );
NAND2_X1 U915 ( .A1(KEYINPUT63), .A2(n1215), .ZN(n1214) );
XOR2_X1 U916 ( .A(n1216), .B(n1130), .Z(n1211) );
INV_X1 U917 ( .A(n1217), .ZN(n1130) );
NAND2_X1 U918 ( .A1(KEYINPUT55), .A2(n1218), .ZN(n1216) );
NOR2_X1 U919 ( .A1(n1030), .A2(n1029), .ZN(n997) );
INV_X1 U920 ( .A(n1032), .ZN(n1029) );
NAND2_X1 U921 ( .A1(G214), .A2(n1219), .ZN(n1032) );
XNOR2_X1 U922 ( .A(n1040), .B(n1220), .ZN(n1030) );
NOR2_X1 U923 ( .A1(n1221), .A2(KEYINPUT13), .ZN(n1220) );
INV_X1 U924 ( .A(n1041), .ZN(n1221) );
NAND2_X1 U925 ( .A1(G210), .A2(n1219), .ZN(n1041) );
NAND2_X1 U926 ( .A1(n1222), .A2(n1223), .ZN(n1219) );
INV_X1 U927 ( .A(G237), .ZN(n1222) );
NAND3_X1 U928 ( .A1(n1224), .A2(n1225), .A3(n1202), .ZN(n1040) );
NAND2_X1 U929 ( .A1(n1226), .A2(n1095), .ZN(n1225) );
NAND2_X1 U930 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NAND2_X1 U931 ( .A1(KEYINPUT39), .A2(n1229), .ZN(n1228) );
NAND2_X1 U932 ( .A1(n1230), .A2(n1231), .ZN(n1227) );
INV_X1 U933 ( .A(KEYINPUT39), .ZN(n1231) );
OR2_X1 U934 ( .A1(n1229), .A2(n1095), .ZN(n1224) );
XOR2_X1 U935 ( .A(n1232), .B(n1233), .Z(n1095) );
XOR2_X1 U936 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U937 ( .A(G122), .B(G119), .Z(n1235) );
XNOR2_X1 U938 ( .A(n1136), .B(n1218), .ZN(n1232) );
XOR2_X1 U939 ( .A(G101), .B(KEYINPUT43), .Z(n1218) );
XOR2_X1 U940 ( .A(n1204), .B(G110), .Z(n1136) );
XNOR2_X1 U941 ( .A(n1114), .B(n1236), .ZN(n1204) );
XOR2_X1 U942 ( .A(KEYINPUT4), .B(G107), .Z(n1236) );
INV_X1 U943 ( .A(G104), .ZN(n1114) );
NAND2_X1 U944 ( .A1(KEYINPUT42), .A2(n1230), .ZN(n1229) );
XNOR2_X1 U945 ( .A(n1237), .B(n1238), .ZN(n1230) );
XOR2_X1 U946 ( .A(KEYINPUT9), .B(n1150), .Z(n1238) );
NOR2_X1 U947 ( .A1(n1090), .A2(G953), .ZN(n1150) );
INV_X1 U948 ( .A(G224), .ZN(n1090) );
NAND2_X1 U949 ( .A1(KEYINPUT6), .A2(n1147), .ZN(n1237) );
XNOR2_X1 U950 ( .A(n1129), .B(G125), .ZN(n1147) );
NOR2_X1 U951 ( .A1(n1038), .A2(n1180), .ZN(n1016) );
NAND3_X1 U952 ( .A1(n1239), .A2(n1240), .A3(n1033), .ZN(n1180) );
OR2_X1 U953 ( .A1(n1043), .A2(G475), .ZN(n1033) );
OR2_X1 U954 ( .A1(G475), .A2(KEYINPUT36), .ZN(n1240) );
NAND3_X1 U955 ( .A1(G475), .A2(n1043), .A3(KEYINPUT36), .ZN(n1239) );
NAND2_X1 U956 ( .A1(n1109), .A2(n1202), .ZN(n1043) );
XNOR2_X1 U957 ( .A(n1241), .B(n1242), .ZN(n1109) );
XNOR2_X1 U958 ( .A(n1243), .B(n1244), .ZN(n1242) );
XOR2_X1 U959 ( .A(n1245), .B(n1075), .Z(n1244) );
NAND2_X1 U960 ( .A1(KEYINPUT51), .A2(n1246), .ZN(n1245) );
XOR2_X1 U961 ( .A(G113), .B(n1247), .Z(n1246) );
XOR2_X1 U962 ( .A(KEYINPUT21), .B(G122), .Z(n1247) );
XOR2_X1 U963 ( .A(n1248), .B(n1249), .Z(n1241) );
XOR2_X1 U964 ( .A(KEYINPUT60), .B(G131), .Z(n1249) );
XOR2_X1 U965 ( .A(n1250), .B(G104), .Z(n1248) );
NAND2_X1 U966 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
OR2_X1 U967 ( .A1(n1253), .A2(KEYINPUT12), .ZN(n1252) );
XOR2_X1 U968 ( .A(n1254), .B(n1255), .Z(n1251) );
AND2_X1 U969 ( .A1(G214), .A2(n1256), .ZN(n1255) );
NAND2_X1 U970 ( .A1(KEYINPUT12), .A2(n1253), .ZN(n1254) );
XNOR2_X1 U971 ( .A(n1178), .B(KEYINPUT24), .ZN(n1253) );
INV_X1 U972 ( .A(n1195), .ZN(n1038) );
XOR2_X1 U973 ( .A(n1106), .B(n1257), .Z(n1195) );
NOR2_X1 U974 ( .A1(n1258), .A2(n1104), .ZN(n1257) );
XOR2_X1 U975 ( .A(n1259), .B(n1260), .Z(n1104) );
NOR2_X1 U976 ( .A1(KEYINPUT14), .A2(n1261), .ZN(n1260) );
XOR2_X1 U977 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U978 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U979 ( .A(G122), .B(G116), .Z(n1265) );
XOR2_X1 U980 ( .A(KEYINPUT33), .B(G128), .Z(n1264) );
XOR2_X1 U981 ( .A(n1266), .B(n1081), .Z(n1262) );
XOR2_X1 U982 ( .A(n1267), .B(G107), .Z(n1266) );
NAND2_X1 U983 ( .A1(KEYINPUT59), .A2(n1178), .ZN(n1267) );
INV_X1 U984 ( .A(G143), .ZN(n1178) );
NAND2_X1 U985 ( .A1(G217), .A2(n1268), .ZN(n1259) );
INV_X1 U986 ( .A(G478), .ZN(n1106) );
XOR2_X1 U987 ( .A(n1269), .B(n1101), .Z(n1025) );
NAND2_X1 U988 ( .A1(G217), .A2(n1199), .ZN(n1101) );
NAND2_X1 U989 ( .A1(G234), .A2(n1223), .ZN(n1199) );
OR2_X1 U990 ( .A1(n1100), .A2(n1258), .ZN(n1269) );
XNOR2_X1 U991 ( .A(n1270), .B(n1271), .ZN(n1100) );
AND2_X1 U992 ( .A1(G221), .A2(n1268), .ZN(n1271) );
AND2_X1 U993 ( .A1(G234), .A2(n1068), .ZN(n1268) );
INV_X1 U994 ( .A(G953), .ZN(n1068) );
XNOR2_X1 U995 ( .A(n1272), .B(n1273), .ZN(n1270) );
NOR2_X1 U996 ( .A1(G137), .A2(KEYINPUT37), .ZN(n1273) );
NOR2_X1 U997 ( .A1(KEYINPUT40), .A2(n1274), .ZN(n1272) );
NOR2_X1 U998 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
XOR2_X1 U999 ( .A(KEYINPUT19), .B(n1277), .Z(n1276) );
AND2_X1 U1000 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NOR2_X1 U1001 ( .A1(n1279), .A2(n1278), .ZN(n1275) );
XOR2_X1 U1002 ( .A(n1075), .B(n1280), .Z(n1278) );
NOR2_X1 U1003 ( .A1(KEYINPUT15), .A2(n1243), .ZN(n1280) );
XOR2_X1 U1004 ( .A(n1213), .B(KEYINPUT11), .Z(n1243) );
XOR2_X1 U1005 ( .A(G125), .B(G140), .Z(n1075) );
XNOR2_X1 U1006 ( .A(n1281), .B(n1282), .ZN(n1279) );
XOR2_X1 U1007 ( .A(KEYINPUT2), .B(G110), .Z(n1282) );
NAND3_X1 U1008 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1281) );
OR2_X1 U1009 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND3_X1 U1010 ( .A1(n1287), .A2(n1286), .A3(KEYINPUT25), .ZN(n1284) );
XNOR2_X1 U1011 ( .A(G128), .B(KEYINPUT27), .ZN(n1286) );
NOR2_X1 U1012 ( .A1(G119), .A2(KEYINPUT8), .ZN(n1287) );
OR2_X1 U1013 ( .A1(n1194), .A2(KEYINPUT25), .ZN(n1283) );
XOR2_X1 U1014 ( .A(n1288), .B(G472), .Z(n1024) );
NAND2_X1 U1015 ( .A1(n1289), .A2(n1202), .ZN(n1288) );
INV_X1 U1016 ( .A(n1258), .ZN(n1202) );
XOR2_X1 U1017 ( .A(n1223), .B(KEYINPUT61), .Z(n1258) );
INV_X1 U1018 ( .A(G902), .ZN(n1223) );
XOR2_X1 U1019 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U1020 ( .A(n1292), .B(n1217), .Z(n1291) );
XNOR2_X1 U1021 ( .A(n1081), .B(n1293), .ZN(n1217) );
XNOR2_X1 U1022 ( .A(n1294), .B(n1295), .ZN(n1293) );
NOR2_X1 U1023 ( .A1(KEYINPUT62), .A2(n1082), .ZN(n1295) );
INV_X1 U1024 ( .A(G131), .ZN(n1082) );
NAND2_X1 U1025 ( .A1(KEYINPUT29), .A2(n1080), .ZN(n1294) );
INV_X1 U1026 ( .A(G137), .ZN(n1080) );
XOR2_X1 U1027 ( .A(G134), .B(KEYINPUT22), .Z(n1081) );
NAND2_X1 U1028 ( .A1(KEYINPUT58), .A2(n1127), .ZN(n1292) );
AND2_X1 U1029 ( .A1(n1296), .A2(n1297), .ZN(n1127) );
NAND2_X1 U1030 ( .A1(n1298), .A2(n1194), .ZN(n1297) );
INV_X1 U1031 ( .A(G119), .ZN(n1194) );
XOR2_X1 U1032 ( .A(KEYINPUT20), .B(n1234), .Z(n1298) );
NAND2_X1 U1033 ( .A1(n1234), .A2(G119), .ZN(n1296) );
XOR2_X1 U1034 ( .A(G113), .B(G116), .Z(n1234) );
XOR2_X1 U1035 ( .A(n1299), .B(n1300), .Z(n1290) );
NOR2_X1 U1036 ( .A1(KEYINPUT50), .A2(n1129), .ZN(n1300) );
XNOR2_X1 U1037 ( .A(n1301), .B(n1302), .ZN(n1129) );
NOR2_X1 U1038 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NOR2_X1 U1039 ( .A1(KEYINPUT53), .A2(n1213), .ZN(n1304) );
AND2_X1 U1040 ( .A1(KEYINPUT46), .A2(n1213), .ZN(n1303) );
XOR2_X1 U1041 ( .A(G146), .B(KEYINPUT18), .Z(n1213) );
XOR2_X1 U1042 ( .A(n1215), .B(G143), .Z(n1301) );
INV_X1 U1043 ( .A(G128), .ZN(n1215) );
NOR2_X1 U1044 ( .A1(n1305), .A2(n1306), .ZN(n1299) );
XOR2_X1 U1045 ( .A(KEYINPUT0), .B(n1307), .Z(n1306) );
NOR2_X1 U1046 ( .A1(n1131), .A2(n1120), .ZN(n1307) );
AND2_X1 U1047 ( .A1(n1131), .A2(n1120), .ZN(n1305) );
NAND2_X1 U1048 ( .A1(n1256), .A2(G210), .ZN(n1120) );
NOR2_X1 U1049 ( .A1(G953), .A2(G237), .ZN(n1256) );
INV_X1 U1050 ( .A(G101), .ZN(n1131) );
endmodule


