//Key = 1010001010010111010111001011100100000011101100101100110011101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385;

XOR2_X1 U772 ( .A(G107), .B(n1062), .Z(G9) );
NOR2_X1 U773 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U774 ( .A1(n1065), .A2(n1066), .ZN(G75) );
NOR4_X1 U775 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
NOR2_X1 U776 ( .A1(n1064), .A2(n1071), .ZN(n1069) );
NAND4_X1 U777 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1067) );
NAND3_X1 U778 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1073) );
XNOR2_X1 U779 ( .A(KEYINPUT44), .B(n1071), .ZN(n1077) );
NAND4_X1 U780 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1082), .ZN(n1071) );
NAND3_X1 U781 ( .A1(n1083), .A2(n1084), .A3(n1079), .ZN(n1072) );
INV_X1 U782 ( .A(n1085), .ZN(n1079) );
NAND3_X1 U783 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1084) );
NAND2_X1 U784 ( .A1(n1081), .A2(n1089), .ZN(n1088) );
NAND2_X1 U785 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U786 ( .A1(n1082), .A2(n1092), .ZN(n1091) );
OR2_X1 U787 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U788 ( .A1(n1095), .A2(n1080), .ZN(n1090) );
XNOR2_X1 U789 ( .A(n1096), .B(KEYINPUT13), .ZN(n1095) );
NAND2_X1 U790 ( .A1(n1080), .A2(n1097), .ZN(n1087) );
NAND2_X1 U791 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U792 ( .A1(n1082), .A2(n1100), .ZN(n1099) );
NAND2_X1 U793 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U794 ( .A1(KEYINPUT31), .A2(n1103), .ZN(n1102) );
OR2_X1 U795 ( .A1(n1104), .A2(n1105), .ZN(n1101) );
NAND2_X1 U796 ( .A1(n1081), .A2(n1106), .ZN(n1098) );
NAND4_X1 U797 ( .A1(n1103), .A2(n1107), .A3(n1082), .A4(n1108), .ZN(n1086) );
INV_X1 U798 ( .A(KEYINPUT31), .ZN(n1107) );
NOR3_X1 U799 ( .A1(n1109), .A2(G953), .A3(G952), .ZN(n1065) );
INV_X1 U800 ( .A(n1074), .ZN(n1109) );
NAND4_X1 U801 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1074) );
NOR3_X1 U802 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1113) );
XOR2_X1 U803 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U804 ( .A1(KEYINPUT11), .A2(n1119), .ZN(n1117) );
XOR2_X1 U805 ( .A(n1120), .B(n1121), .Z(n1115) );
XOR2_X1 U806 ( .A(KEYINPUT60), .B(n1122), .Z(n1121) );
NAND2_X1 U807 ( .A1(KEYINPUT6), .A2(n1123), .ZN(n1120) );
NAND3_X1 U808 ( .A1(n1104), .A2(n1124), .A3(n1125), .ZN(n1114) );
NAND2_X1 U809 ( .A1(G469), .A2(n1126), .ZN(n1125) );
NOR3_X1 U810 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1112) );
NOR2_X1 U811 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
INV_X1 U812 ( .A(KEYINPUT42), .ZN(n1131) );
NOR2_X1 U813 ( .A1(n1132), .A2(n1133), .ZN(n1130) );
NOR3_X1 U814 ( .A1(n1126), .A2(KEYINPUT59), .A3(G469), .ZN(n1133) );
AND2_X1 U815 ( .A1(n1126), .A2(KEYINPUT59), .ZN(n1132) );
NOR2_X1 U816 ( .A1(KEYINPUT42), .A2(n1134), .ZN(n1128) );
NOR2_X1 U817 ( .A1(G469), .A2(n1135), .ZN(n1134) );
XOR2_X1 U818 ( .A(n1126), .B(KEYINPUT59), .Z(n1135) );
XNOR2_X1 U819 ( .A(G472), .B(n1136), .ZN(n1127) );
XOR2_X1 U820 ( .A(KEYINPUT5), .B(n1137), .Z(n1111) );
XOR2_X1 U821 ( .A(n1138), .B(n1139), .Z(G72) );
XOR2_X1 U822 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U823 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
INV_X1 U824 ( .A(n1144), .ZN(n1143) );
XOR2_X1 U825 ( .A(n1145), .B(n1146), .Z(n1142) );
XOR2_X1 U826 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U827 ( .A(n1149), .B(n1150), .Z(n1145) );
NOR2_X1 U828 ( .A1(KEYINPUT33), .A2(n1151), .ZN(n1150) );
XNOR2_X1 U829 ( .A(KEYINPUT8), .B(KEYINPUT39), .ZN(n1149) );
NAND2_X1 U830 ( .A1(G953), .A2(n1152), .ZN(n1140) );
NAND2_X1 U831 ( .A1(G227), .A2(n1153), .ZN(n1152) );
XOR2_X1 U832 ( .A(KEYINPUT47), .B(G900), .Z(n1153) );
NOR2_X1 U833 ( .A1(n1154), .A2(G953), .ZN(n1138) );
XOR2_X1 U834 ( .A(n1155), .B(n1156), .Z(G69) );
NOR2_X1 U835 ( .A1(n1157), .A2(n1075), .ZN(n1156) );
NOR2_X1 U836 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NOR2_X1 U837 ( .A1(KEYINPUT50), .A2(n1160), .ZN(n1155) );
XOR2_X1 U838 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U839 ( .A1(n1163), .A2(G953), .ZN(n1162) );
NAND2_X1 U840 ( .A1(n1164), .A2(n1165), .ZN(n1161) );
NAND2_X1 U841 ( .A1(G953), .A2(n1159), .ZN(n1165) );
XOR2_X1 U842 ( .A(n1166), .B(n1167), .Z(n1164) );
XOR2_X1 U843 ( .A(n1168), .B(KEYINPUT61), .Z(n1167) );
NAND2_X1 U844 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
OR2_X1 U845 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U846 ( .A1(n1173), .A2(n1174), .ZN(G66) );
NOR3_X1 U847 ( .A1(n1118), .A2(n1175), .A3(n1176), .ZN(n1174) );
NOR3_X1 U848 ( .A1(n1177), .A2(n1119), .A3(n1178), .ZN(n1176) );
INV_X1 U849 ( .A(n1179), .ZN(n1177) );
NOR2_X1 U850 ( .A1(n1180), .A2(n1179), .ZN(n1175) );
NOR2_X1 U851 ( .A1(n1181), .A2(n1119), .ZN(n1180) );
NOR2_X1 U852 ( .A1(n1070), .A2(n1068), .ZN(n1181) );
NOR2_X1 U853 ( .A1(n1173), .A2(n1182), .ZN(G63) );
XOR2_X1 U854 ( .A(n1183), .B(n1184), .Z(n1182) );
AND2_X1 U855 ( .A1(G478), .A2(n1185), .ZN(n1184) );
NOR2_X1 U856 ( .A1(KEYINPUT30), .A2(n1186), .ZN(n1183) );
XOR2_X1 U857 ( .A(KEYINPUT15), .B(n1187), .Z(n1186) );
NOR2_X1 U858 ( .A1(n1173), .A2(n1188), .ZN(G60) );
XNOR2_X1 U859 ( .A(n1189), .B(n1190), .ZN(n1188) );
AND2_X1 U860 ( .A1(G475), .A2(n1185), .ZN(n1190) );
XOR2_X1 U861 ( .A(G104), .B(n1191), .Z(G6) );
NOR2_X1 U862 ( .A1(KEYINPUT9), .A2(n1192), .ZN(n1191) );
NOR3_X1 U863 ( .A1(n1193), .A2(n1173), .A3(n1194), .ZN(G57) );
NOR3_X1 U864 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1194) );
XNOR2_X1 U865 ( .A(n1198), .B(n1199), .ZN(n1196) );
NOR2_X1 U866 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
INV_X1 U867 ( .A(KEYINPUT63), .ZN(n1201) );
NOR2_X1 U868 ( .A1(n1202), .A2(n1203), .ZN(n1193) );
XOR2_X1 U869 ( .A(n1204), .B(n1198), .Z(n1203) );
XOR2_X1 U870 ( .A(n1205), .B(G101), .Z(n1198) );
NAND2_X1 U871 ( .A1(n1200), .A2(KEYINPUT63), .ZN(n1204) );
AND2_X1 U872 ( .A1(n1185), .A2(G472), .ZN(n1200) );
NOR2_X1 U873 ( .A1(n1197), .A2(n1195), .ZN(n1202) );
INV_X1 U874 ( .A(KEYINPUT0), .ZN(n1195) );
XNOR2_X1 U875 ( .A(n1206), .B(n1207), .ZN(n1197) );
NAND2_X1 U876 ( .A1(n1208), .A2(n1209), .ZN(n1206) );
OR2_X1 U877 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U878 ( .A(n1212), .B(KEYINPUT16), .Z(n1208) );
NAND2_X1 U879 ( .A1(n1210), .A2(n1211), .ZN(n1212) );
NOR2_X1 U880 ( .A1(n1173), .A2(n1213), .ZN(G54) );
XOR2_X1 U881 ( .A(n1214), .B(n1215), .Z(n1213) );
XNOR2_X1 U882 ( .A(n1210), .B(n1216), .ZN(n1215) );
XOR2_X1 U883 ( .A(n1217), .B(n1218), .Z(n1214) );
XOR2_X1 U884 ( .A(n1219), .B(n1220), .Z(n1218) );
NAND2_X1 U885 ( .A1(n1221), .A2(KEYINPUT17), .ZN(n1220) );
XOR2_X1 U886 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR2_X1 U887 ( .A1(G110), .A2(KEYINPUT34), .ZN(n1223) );
INV_X1 U888 ( .A(G140), .ZN(n1222) );
AND2_X1 U889 ( .A1(G469), .A2(n1185), .ZN(n1217) );
NOR3_X1 U890 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(G51) );
NOR3_X1 U891 ( .A1(n1227), .A2(G953), .A3(G952), .ZN(n1226) );
AND2_X1 U892 ( .A1(n1227), .A2(n1173), .ZN(n1225) );
NOR2_X1 U893 ( .A1(n1075), .A2(G952), .ZN(n1173) );
INV_X1 U894 ( .A(KEYINPUT35), .ZN(n1227) );
XOR2_X1 U895 ( .A(n1228), .B(n1229), .Z(n1224) );
XOR2_X1 U896 ( .A(n1230), .B(n1231), .Z(n1229) );
NOR2_X1 U897 ( .A1(KEYINPUT18), .A2(n1232), .ZN(n1231) );
XNOR2_X1 U898 ( .A(KEYINPUT58), .B(n1233), .ZN(n1232) );
NAND2_X1 U899 ( .A1(n1185), .A2(n1122), .ZN(n1230) );
INV_X1 U900 ( .A(n1178), .ZN(n1185) );
NAND2_X1 U901 ( .A1(G902), .A2(n1234), .ZN(n1178) );
NAND2_X1 U902 ( .A1(n1154), .A2(n1163), .ZN(n1234) );
INV_X1 U903 ( .A(n1070), .ZN(n1163) );
NAND4_X1 U904 ( .A1(n1192), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1070) );
AND4_X1 U905 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1237) );
NOR3_X1 U906 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1236) );
NOR2_X1 U907 ( .A1(n1064), .A2(n1245), .ZN(n1244) );
XNOR2_X1 U908 ( .A(KEYINPUT57), .B(n1063), .ZN(n1245) );
NAND4_X1 U909 ( .A1(n1094), .A2(n1082), .A3(n1103), .A4(n1246), .ZN(n1063) );
NOR4_X1 U910 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1108), .ZN(n1243) );
INV_X1 U911 ( .A(n1106), .ZN(n1249) );
NAND3_X1 U912 ( .A1(n1246), .A2(n1250), .A3(n1103), .ZN(n1248) );
NOR2_X1 U913 ( .A1(n1251), .A2(n1250), .ZN(n1242) );
INV_X1 U914 ( .A(KEYINPUT43), .ZN(n1250) );
NAND3_X1 U915 ( .A1(n1093), .A2(n1082), .A3(n1252), .ZN(n1192) );
INV_X1 U916 ( .A(n1068), .ZN(n1154) );
NAND4_X1 U917 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1068) );
NOR4_X1 U918 ( .A1(n1257), .A2(n1258), .A3(n1259), .A4(n1260), .ZN(n1256) );
INV_X1 U919 ( .A(n1261), .ZN(n1258) );
NOR2_X1 U920 ( .A1(n1262), .A2(n1263), .ZN(n1255) );
NAND3_X1 U921 ( .A1(n1264), .A2(n1103), .A3(n1265), .ZN(n1253) );
XOR2_X1 U922 ( .A(n1266), .B(KEYINPUT1), .Z(n1265) );
INV_X1 U923 ( .A(n1267), .ZN(n1264) );
XOR2_X1 U924 ( .A(G146), .B(n1257), .Z(G48) );
AND3_X1 U925 ( .A1(n1268), .A2(n1247), .A3(n1093), .ZN(n1257) );
XOR2_X1 U926 ( .A(n1269), .B(n1254), .Z(G45) );
NAND4_X1 U927 ( .A1(n1270), .A2(n1247), .A3(n1096), .A4(n1271), .ZN(n1254) );
NOR3_X1 U928 ( .A1(n1272), .A2(n1273), .A3(n1110), .ZN(n1271) );
XOR2_X1 U929 ( .A(G140), .B(n1263), .Z(G42) );
AND2_X1 U930 ( .A1(n1274), .A2(n1106), .ZN(n1263) );
XOR2_X1 U931 ( .A(G137), .B(n1262), .Z(G39) );
AND3_X1 U932 ( .A1(n1083), .A2(n1268), .A3(n1080), .ZN(n1262) );
XOR2_X1 U933 ( .A(n1275), .B(n1276), .Z(G36) );
NOR2_X1 U934 ( .A1(KEYINPUT23), .A2(n1277), .ZN(n1276) );
INV_X1 U935 ( .A(G134), .ZN(n1277) );
NOR3_X1 U936 ( .A1(n1267), .A2(n1273), .A3(n1278), .ZN(n1275) );
XOR2_X1 U937 ( .A(n1272), .B(KEYINPUT7), .Z(n1278) );
INV_X1 U938 ( .A(n1266), .ZN(n1273) );
NAND3_X1 U939 ( .A1(n1083), .A2(n1094), .A3(n1096), .ZN(n1267) );
XOR2_X1 U940 ( .A(G131), .B(n1260), .Z(G33) );
AND2_X1 U941 ( .A1(n1096), .A2(n1274), .ZN(n1260) );
AND4_X1 U942 ( .A1(n1083), .A2(n1093), .A3(n1103), .A4(n1266), .ZN(n1274) );
NOR2_X1 U943 ( .A1(n1279), .A2(n1078), .ZN(n1083) );
INV_X1 U944 ( .A(n1124), .ZN(n1078) );
XOR2_X1 U945 ( .A(G128), .B(n1259), .Z(G30) );
AND3_X1 U946 ( .A1(n1247), .A2(n1094), .A3(n1268), .ZN(n1259) );
AND4_X1 U947 ( .A1(n1103), .A2(n1280), .A3(n1281), .A4(n1266), .ZN(n1268) );
XOR2_X1 U948 ( .A(n1282), .B(n1235), .Z(G3) );
NAND3_X1 U949 ( .A1(n1080), .A2(n1096), .A3(n1252), .ZN(n1235) );
XOR2_X1 U950 ( .A(n1283), .B(n1261), .Z(G27) );
NAND3_X1 U951 ( .A1(n1081), .A2(n1106), .A3(n1284), .ZN(n1261) );
AND3_X1 U952 ( .A1(n1093), .A2(n1266), .A3(n1247), .ZN(n1284) );
NAND2_X1 U953 ( .A1(n1285), .A2(n1085), .ZN(n1266) );
NAND3_X1 U954 ( .A1(G902), .A2(n1286), .A3(n1144), .ZN(n1285) );
NOR2_X1 U955 ( .A1(n1075), .A2(G900), .ZN(n1144) );
XOR2_X1 U956 ( .A(n1287), .B(n1241), .Z(G24) );
NAND4_X1 U957 ( .A1(n1270), .A2(n1288), .A3(n1082), .A4(n1289), .ZN(n1241) );
NOR2_X1 U958 ( .A1(n1281), .A2(n1280), .ZN(n1082) );
XOR2_X1 U959 ( .A(n1290), .B(n1240), .Z(G21) );
NAND4_X1 U960 ( .A1(n1288), .A2(n1080), .A3(n1280), .A4(n1281), .ZN(n1240) );
INV_X1 U961 ( .A(n1291), .ZN(n1280) );
XOR2_X1 U962 ( .A(n1239), .B(n1292), .Z(G18) );
XNOR2_X1 U963 ( .A(G116), .B(KEYINPUT10), .ZN(n1292) );
NAND3_X1 U964 ( .A1(n1096), .A2(n1094), .A3(n1288), .ZN(n1239) );
NOR2_X1 U965 ( .A1(n1270), .A2(n1110), .ZN(n1094) );
XOR2_X1 U966 ( .A(n1238), .B(n1293), .Z(G15) );
XOR2_X1 U967 ( .A(KEYINPUT38), .B(G113), .Z(n1293) );
NAND3_X1 U968 ( .A1(n1096), .A2(n1093), .A3(n1288), .ZN(n1238) );
AND3_X1 U969 ( .A1(n1247), .A2(n1246), .A3(n1081), .ZN(n1288) );
NOR2_X1 U970 ( .A1(n1105), .A2(n1294), .ZN(n1081) );
INV_X1 U971 ( .A(n1104), .ZN(n1294) );
NOR2_X1 U972 ( .A1(n1289), .A2(n1137), .ZN(n1093) );
INV_X1 U973 ( .A(n1110), .ZN(n1289) );
AND2_X1 U974 ( .A1(n1291), .A2(n1281), .ZN(n1096) );
XOR2_X1 U975 ( .A(n1251), .B(n1295), .Z(G12) );
NAND2_X1 U976 ( .A1(KEYINPUT2), .A2(G110), .ZN(n1295) );
NAND3_X1 U977 ( .A1(n1080), .A2(n1106), .A3(n1252), .ZN(n1251) );
AND3_X1 U978 ( .A1(n1103), .A2(n1246), .A3(n1247), .ZN(n1252) );
INV_X1 U979 ( .A(n1064), .ZN(n1247) );
NAND2_X1 U980 ( .A1(n1279), .A2(n1124), .ZN(n1064) );
NAND2_X1 U981 ( .A1(G214), .A2(n1296), .ZN(n1124) );
INV_X1 U982 ( .A(n1076), .ZN(n1279) );
XNOR2_X1 U983 ( .A(n1123), .B(n1122), .ZN(n1076) );
AND2_X1 U984 ( .A1(G210), .A2(n1296), .ZN(n1122) );
NAND2_X1 U985 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XOR2_X1 U986 ( .A(n1299), .B(KEYINPUT12), .Z(n1297) );
AND2_X1 U987 ( .A1(n1300), .A2(n1298), .ZN(n1123) );
XOR2_X1 U988 ( .A(n1301), .B(n1302), .Z(n1300) );
XNOR2_X1 U989 ( .A(n1303), .B(KEYINPUT29), .ZN(n1302) );
NAND2_X1 U990 ( .A1(KEYINPUT27), .A2(n1233), .ZN(n1303) );
XNOR2_X1 U991 ( .A(n1304), .B(n1211), .ZN(n1233) );
XOR2_X1 U992 ( .A(n1283), .B(n1305), .Z(n1304) );
NOR2_X1 U993 ( .A1(G953), .A2(n1158), .ZN(n1305) );
INV_X1 U994 ( .A(G224), .ZN(n1158) );
INV_X1 U995 ( .A(n1228), .ZN(n1301) );
XOR2_X1 U996 ( .A(n1306), .B(n1307), .Z(n1228) );
INV_X1 U997 ( .A(n1166), .ZN(n1307) );
XNOR2_X1 U998 ( .A(G110), .B(n1308), .ZN(n1166) );
XOR2_X1 U999 ( .A(KEYINPUT53), .B(G122), .Z(n1308) );
NAND3_X1 U1000 ( .A1(n1309), .A2(n1310), .A3(n1169), .ZN(n1306) );
NAND2_X1 U1001 ( .A1(n1172), .A2(n1171), .ZN(n1169) );
OR3_X1 U1002 ( .A1(n1171), .A2(n1172), .A3(KEYINPUT51), .ZN(n1310) );
AND2_X1 U1003 ( .A1(n1311), .A2(n1312), .ZN(n1172) );
NAND2_X1 U1004 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U1005 ( .A(KEYINPUT40), .B(G113), .Z(n1314) );
XOR2_X1 U1006 ( .A(G119), .B(G116), .Z(n1313) );
NAND2_X1 U1007 ( .A1(n1315), .A2(n1316), .ZN(n1311) );
XNOR2_X1 U1008 ( .A(G113), .B(KEYINPUT49), .ZN(n1316) );
XOR2_X1 U1009 ( .A(G116), .B(n1290), .Z(n1315) );
NAND2_X1 U1010 ( .A1(KEYINPUT51), .A2(n1171), .ZN(n1309) );
NAND2_X1 U1011 ( .A1(n1085), .A2(n1317), .ZN(n1246) );
NAND4_X1 U1012 ( .A1(G953), .A2(G902), .A3(n1286), .A4(n1159), .ZN(n1317) );
INV_X1 U1013 ( .A(G898), .ZN(n1159) );
NAND3_X1 U1014 ( .A1(n1286), .A2(n1075), .A3(G952), .ZN(n1085) );
NAND2_X1 U1015 ( .A1(G234), .A2(G237), .ZN(n1286) );
INV_X1 U1016 ( .A(n1272), .ZN(n1103) );
NAND2_X1 U1017 ( .A1(n1105), .A2(n1104), .ZN(n1272) );
NAND2_X1 U1018 ( .A1(G221), .A2(n1318), .ZN(n1104) );
XNOR2_X1 U1019 ( .A(n1126), .B(G469), .ZN(n1105) );
NAND2_X1 U1020 ( .A1(n1319), .A2(n1298), .ZN(n1126) );
XOR2_X1 U1021 ( .A(n1210), .B(n1320), .Z(n1319) );
XNOR2_X1 U1022 ( .A(n1321), .B(n1322), .ZN(n1320) );
NAND2_X1 U1023 ( .A1(KEYINPUT46), .A2(n1216), .ZN(n1322) );
XNOR2_X1 U1024 ( .A(n1171), .B(n1151), .ZN(n1216) );
XNOR2_X1 U1025 ( .A(n1323), .B(n1324), .ZN(n1151) );
XOR2_X1 U1026 ( .A(G146), .B(n1325), .Z(n1324) );
NOR2_X1 U1027 ( .A1(KEYINPUT32), .A2(n1269), .ZN(n1325) );
INV_X1 U1028 ( .A(G143), .ZN(n1269) );
XNOR2_X1 U1029 ( .A(n1326), .B(n1327), .ZN(n1171) );
XOR2_X1 U1030 ( .A(KEYINPUT52), .B(G104), .Z(n1327) );
XOR2_X1 U1031 ( .A(n1282), .B(n1328), .Z(n1326) );
INV_X1 U1032 ( .A(G101), .ZN(n1282) );
NAND2_X1 U1033 ( .A1(n1329), .A2(KEYINPUT20), .ZN(n1321) );
XOR2_X1 U1034 ( .A(n1219), .B(n1330), .Z(n1329) );
XOR2_X1 U1035 ( .A(G140), .B(G110), .Z(n1330) );
NAND2_X1 U1036 ( .A1(G227), .A2(n1075), .ZN(n1219) );
NOR2_X1 U1037 ( .A1(n1281), .A2(n1291), .ZN(n1106) );
XOR2_X1 U1038 ( .A(n1119), .B(n1118), .Z(n1291) );
NOR2_X1 U1039 ( .A1(n1179), .A2(G902), .ZN(n1118) );
NAND3_X1 U1040 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(n1179) );
OR2_X1 U1041 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NAND3_X1 U1042 ( .A1(n1336), .A2(n1334), .A3(n1337), .ZN(n1332) );
INV_X1 U1043 ( .A(KEYINPUT3), .ZN(n1334) );
OR2_X1 U1044 ( .A1(n1337), .A2(n1336), .ZN(n1331) );
AND2_X1 U1045 ( .A1(KEYINPUT28), .A2(n1335), .ZN(n1336) );
XNOR2_X1 U1046 ( .A(n1338), .B(n1339), .ZN(n1335) );
NOR2_X1 U1047 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
INV_X1 U1048 ( .A(G221), .ZN(n1341) );
INV_X1 U1049 ( .A(G137), .ZN(n1338) );
XNOR2_X1 U1050 ( .A(n1342), .B(n1343), .ZN(n1337) );
XOR2_X1 U1051 ( .A(G110), .B(n1344), .Z(n1343) );
NOR2_X1 U1052 ( .A1(KEYINPUT36), .A2(n1345), .ZN(n1344) );
XOR2_X1 U1053 ( .A(n1346), .B(n1347), .Z(n1345) );
XOR2_X1 U1054 ( .A(n1348), .B(G140), .Z(n1347) );
NAND2_X1 U1055 ( .A1(KEYINPUT21), .A2(G146), .ZN(n1348) );
NAND2_X1 U1056 ( .A1(KEYINPUT26), .A2(n1283), .ZN(n1346) );
INV_X1 U1057 ( .A(G125), .ZN(n1283) );
XOR2_X1 U1058 ( .A(n1290), .B(G128), .Z(n1342) );
NAND2_X1 U1059 ( .A1(G217), .A2(n1318), .ZN(n1119) );
NAND2_X1 U1060 ( .A1(G234), .A2(n1298), .ZN(n1318) );
NAND2_X1 U1061 ( .A1(n1349), .A2(n1350), .ZN(n1281) );
NAND2_X1 U1062 ( .A1(G472), .A2(n1136), .ZN(n1350) );
XOR2_X1 U1063 ( .A(n1351), .B(KEYINPUT45), .Z(n1349) );
OR2_X1 U1064 ( .A1(n1136), .A2(G472), .ZN(n1351) );
NAND2_X1 U1065 ( .A1(n1352), .A2(n1298), .ZN(n1136) );
XOR2_X1 U1066 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1067 ( .A(n1355), .B(G101), .Z(n1354) );
NAND2_X1 U1068 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
NAND2_X1 U1069 ( .A1(n1358), .A2(n1207), .ZN(n1357) );
XOR2_X1 U1070 ( .A(n1359), .B(KEYINPUT62), .Z(n1356) );
OR2_X1 U1071 ( .A1(n1207), .A2(n1358), .ZN(n1359) );
XOR2_X1 U1072 ( .A(n1210), .B(n1211), .Z(n1358) );
XOR2_X1 U1073 ( .A(n1360), .B(n1323), .Z(n1211) );
XOR2_X1 U1074 ( .A(G128), .B(KEYINPUT22), .Z(n1323) );
XNOR2_X1 U1075 ( .A(n1147), .B(KEYINPUT4), .ZN(n1210) );
XOR2_X1 U1076 ( .A(G131), .B(n1361), .Z(n1147) );
XOR2_X1 U1077 ( .A(G137), .B(G134), .Z(n1361) );
XOR2_X1 U1078 ( .A(G113), .B(n1362), .Z(n1207) );
NOR2_X1 U1079 ( .A1(KEYINPUT55), .A2(n1363), .ZN(n1362) );
XNOR2_X1 U1080 ( .A(G116), .B(n1364), .ZN(n1363) );
NAND2_X1 U1081 ( .A1(KEYINPUT14), .A2(n1290), .ZN(n1364) );
INV_X1 U1082 ( .A(G119), .ZN(n1290) );
NAND2_X1 U1083 ( .A1(KEYINPUT19), .A2(n1205), .ZN(n1353) );
AND3_X1 U1084 ( .A1(n1299), .A2(n1075), .A3(G210), .ZN(n1205) );
INV_X1 U1085 ( .A(n1108), .ZN(n1080) );
NAND2_X1 U1086 ( .A1(n1110), .A2(n1137), .ZN(n1108) );
INV_X1 U1087 ( .A(n1270), .ZN(n1137) );
XOR2_X1 U1088 ( .A(n1365), .B(n1366), .Z(n1270) );
XOR2_X1 U1089 ( .A(KEYINPUT56), .B(G475), .Z(n1366) );
NAND2_X1 U1090 ( .A1(n1189), .A2(n1298), .ZN(n1365) );
INV_X1 U1091 ( .A(G902), .ZN(n1298) );
XNOR2_X1 U1092 ( .A(n1367), .B(n1368), .ZN(n1189) );
XOR2_X1 U1093 ( .A(n1369), .B(n1370), .Z(n1368) );
XNOR2_X1 U1094 ( .A(G104), .B(G131), .ZN(n1370) );
NAND2_X1 U1095 ( .A1(n1371), .A2(KEYINPUT48), .ZN(n1369) );
XNOR2_X1 U1096 ( .A(G113), .B(n1372), .ZN(n1371) );
NOR2_X1 U1097 ( .A1(G122), .A2(KEYINPUT37), .ZN(n1372) );
XOR2_X1 U1098 ( .A(n1373), .B(n1148), .Z(n1367) );
XOR2_X1 U1099 ( .A(G125), .B(G140), .Z(n1148) );
XNOR2_X1 U1100 ( .A(n1374), .B(n1360), .ZN(n1373) );
XNOR2_X1 U1101 ( .A(G143), .B(G146), .ZN(n1360) );
NAND3_X1 U1102 ( .A1(n1299), .A2(n1075), .A3(G214), .ZN(n1374) );
INV_X1 U1103 ( .A(G237), .ZN(n1299) );
XOR2_X1 U1104 ( .A(n1375), .B(G478), .Z(n1110) );
OR2_X1 U1105 ( .A1(n1187), .A2(G902), .ZN(n1375) );
XNOR2_X1 U1106 ( .A(n1376), .B(n1377), .ZN(n1187) );
XNOR2_X1 U1107 ( .A(n1378), .B(n1328), .ZN(n1377) );
XOR2_X1 U1108 ( .A(G107), .B(KEYINPUT54), .Z(n1328) );
NAND2_X1 U1109 ( .A1(KEYINPUT24), .A2(n1379), .ZN(n1378) );
XOR2_X1 U1110 ( .A(n1380), .B(n1381), .Z(n1379) );
XOR2_X1 U1111 ( .A(G143), .B(G134), .Z(n1381) );
NOR2_X1 U1112 ( .A1(G128), .A2(KEYINPUT25), .ZN(n1380) );
XOR2_X1 U1113 ( .A(n1382), .B(n1383), .Z(n1376) );
NOR2_X1 U1114 ( .A1(n1340), .A2(n1384), .ZN(n1383) );
INV_X1 U1115 ( .A(G217), .ZN(n1384) );
NAND2_X1 U1116 ( .A1(n1385), .A2(n1075), .ZN(n1340) );
INV_X1 U1117 ( .A(G953), .ZN(n1075) );
XOR2_X1 U1118 ( .A(KEYINPUT41), .B(G234), .Z(n1385) );
XOR2_X1 U1119 ( .A(G116), .B(n1287), .Z(n1382) );
INV_X1 U1120 ( .A(G122), .ZN(n1287) );
endmodule


