//Key = 0011101010111110111011100100110000100000000100101001010001011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;

XNOR2_X1 U723 ( .A(G107), .B(n995), .ZN(G9) );
NOR2_X1 U724 ( .A1(n996), .A2(n997), .ZN(G75) );
NOR4_X1 U725 ( .A1(G953), .A2(n998), .A3(n999), .A4(n1000), .ZN(n997) );
NOR2_X1 U726 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NOR2_X1 U727 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
NOR4_X1 U728 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1004) );
NOR4_X1 U729 ( .A1(n1009), .A2(n1010), .A3(n1011), .A4(n1012), .ZN(n1006) );
NOR2_X1 U730 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NOR3_X1 U731 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1011) );
NOR2_X1 U732 ( .A1(n1018), .A2(n1019), .ZN(n1005) );
NOR2_X1 U733 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
NOR4_X1 U734 ( .A1(n1009), .A2(n1020), .A3(n1014), .A4(n1015), .ZN(n1003) );
NOR2_X1 U735 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U736 ( .A1(n1023), .A2(n1008), .ZN(n1022) );
INV_X1 U737 ( .A(n1024), .ZN(n1008) );
NOR2_X1 U738 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
AND2_X1 U739 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR2_X1 U740 ( .A1(n1029), .A2(n1007), .ZN(n1021) );
NOR2_X1 U741 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR3_X1 U742 ( .A1(n998), .A2(G953), .A3(G952), .ZN(n996) );
AND4_X1 U743 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n998) );
NOR4_X1 U744 ( .A1(n1009), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1035) );
XOR2_X1 U745 ( .A(n1039), .B(G475), .Z(n1038) );
NAND2_X1 U746 ( .A1(KEYINPUT10), .A2(n1040), .ZN(n1039) );
XNOR2_X1 U747 ( .A(n1041), .B(n1042), .ZN(n1037) );
NOR2_X1 U748 ( .A1(G478), .A2(KEYINPUT44), .ZN(n1042) );
INV_X1 U749 ( .A(n1019), .ZN(n1009) );
NOR2_X1 U750 ( .A1(n1043), .A2(n1044), .ZN(n1034) );
NOR3_X1 U751 ( .A1(n1045), .A2(G469), .A3(n1046), .ZN(n1044) );
NOR2_X1 U752 ( .A1(n1047), .A2(n1048), .ZN(n1043) );
NOR2_X1 U753 ( .A1(G469), .A2(n1046), .ZN(n1048) );
INV_X1 U754 ( .A(KEYINPUT22), .ZN(n1046) );
XOR2_X1 U755 ( .A(KEYINPUT11), .B(n1049), .Z(n1033) );
NAND2_X1 U756 ( .A1(n1050), .A2(n1051), .ZN(G72) );
NAND2_X1 U757 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U758 ( .A1(G953), .A2(n1054), .ZN(n1053) );
NAND3_X1 U759 ( .A1(G953), .A2(n1055), .A3(n1056), .ZN(n1050) );
INV_X1 U760 ( .A(n1052), .ZN(n1056) );
XNOR2_X1 U761 ( .A(n1057), .B(n1058), .ZN(n1052) );
NOR2_X1 U762 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XOR2_X1 U763 ( .A(n1061), .B(n1062), .Z(n1060) );
XNOR2_X1 U764 ( .A(n1063), .B(n1064), .ZN(n1062) );
XOR2_X1 U765 ( .A(n1065), .B(n1066), .Z(n1061) );
NOR2_X1 U766 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XOR2_X1 U767 ( .A(n1069), .B(KEYINPUT17), .Z(n1068) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR2_X1 U769 ( .A1(n1070), .A2(n1071), .ZN(n1067) );
XNOR2_X1 U770 ( .A(G134), .B(n1072), .ZN(n1070) );
XNOR2_X1 U771 ( .A(KEYINPUT33), .B(n1073), .ZN(n1072) );
XNOR2_X1 U772 ( .A(G140), .B(KEYINPUT32), .ZN(n1065) );
NOR2_X1 U773 ( .A1(G900), .A2(n1074), .ZN(n1059) );
NAND3_X1 U774 ( .A1(n1075), .A2(n1074), .A3(KEYINPUT48), .ZN(n1057) );
NAND2_X1 U775 ( .A1(G900), .A2(G227), .ZN(n1055) );
XOR2_X1 U776 ( .A(n1076), .B(n1077), .Z(G69) );
XOR2_X1 U777 ( .A(n1078), .B(n1079), .Z(n1077) );
NAND2_X1 U778 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XNOR2_X1 U779 ( .A(n1082), .B(n1083), .ZN(n1081) );
XNOR2_X1 U780 ( .A(n1084), .B(KEYINPUT24), .ZN(n1080) );
NAND2_X1 U781 ( .A1(n1085), .A2(n1086), .ZN(n1078) );
NAND2_X1 U782 ( .A1(G898), .A2(G224), .ZN(n1086) );
XNOR2_X1 U783 ( .A(G953), .B(KEYINPUT16), .ZN(n1085) );
NOR2_X1 U784 ( .A1(G953), .A2(n1087), .ZN(n1076) );
NOR3_X1 U785 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1087) );
NAND3_X1 U786 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1088) );
NOR2_X1 U787 ( .A1(n1094), .A2(n1095), .ZN(G66) );
XNOR2_X1 U788 ( .A(n1096), .B(n1097), .ZN(n1095) );
NAND2_X1 U789 ( .A1(n1098), .A2(G217), .ZN(n1096) );
NOR2_X1 U790 ( .A1(n1094), .A2(n1099), .ZN(G63) );
NOR3_X1 U791 ( .A1(n1041), .A2(n1100), .A3(n1101), .ZN(n1099) );
AND3_X1 U792 ( .A1(n1102), .A2(G478), .A3(n1098), .ZN(n1101) );
NOR2_X1 U793 ( .A1(n1103), .A2(n1102), .ZN(n1100) );
AND2_X1 U794 ( .A1(n1000), .A2(G478), .ZN(n1103) );
NOR2_X1 U795 ( .A1(n1094), .A2(n1104), .ZN(G60) );
XOR2_X1 U796 ( .A(n1105), .B(n1106), .Z(n1104) );
XOR2_X1 U797 ( .A(n1107), .B(KEYINPUT35), .Z(n1105) );
NAND2_X1 U798 ( .A1(n1098), .A2(G475), .ZN(n1107) );
XNOR2_X1 U799 ( .A(n1108), .B(n1109), .ZN(G6) );
XNOR2_X1 U800 ( .A(KEYINPUT9), .B(n1110), .ZN(n1109) );
NOR2_X1 U801 ( .A1(n1094), .A2(n1111), .ZN(G57) );
XOR2_X1 U802 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U803 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U804 ( .A1(n1098), .A2(G472), .ZN(n1115) );
NAND3_X1 U805 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1114) );
OR2_X1 U806 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND3_X1 U807 ( .A1(n1120), .A2(n1119), .A3(KEYINPUT2), .ZN(n1117) );
AND2_X1 U808 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U809 ( .A(KEYINPUT7), .B(KEYINPUT29), .Z(n1121) );
OR2_X1 U810 ( .A1(n1122), .A2(KEYINPUT2), .ZN(n1116) );
XOR2_X1 U811 ( .A(n1123), .B(n1124), .Z(n1112) );
XNOR2_X1 U812 ( .A(KEYINPUT13), .B(n1125), .ZN(n1124) );
NOR2_X1 U813 ( .A1(n1094), .A2(n1126), .ZN(G54) );
XOR2_X1 U814 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U815 ( .A(n1129), .B(n1130), .Z(n1128) );
XNOR2_X1 U816 ( .A(n1131), .B(n1132), .ZN(n1130) );
NOR2_X1 U817 ( .A1(KEYINPUT61), .A2(n1133), .ZN(n1132) );
NOR2_X1 U818 ( .A1(KEYINPUT54), .A2(n1134), .ZN(n1131) );
XNOR2_X1 U819 ( .A(n1135), .B(n1136), .ZN(n1134) );
XNOR2_X1 U820 ( .A(n1137), .B(G110), .ZN(n1136) );
NAND2_X1 U821 ( .A1(n1098), .A2(G469), .ZN(n1129) );
INV_X1 U822 ( .A(n1138), .ZN(n1098) );
XOR2_X1 U823 ( .A(n1139), .B(n1064), .Z(n1127) );
NOR2_X1 U824 ( .A1(n1094), .A2(n1140), .ZN(G51) );
XOR2_X1 U825 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U826 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U827 ( .A(n1145), .B(n1146), .ZN(n1144) );
NOR2_X1 U828 ( .A1(KEYINPUT58), .A2(n1063), .ZN(n1146) );
NAND2_X1 U829 ( .A1(KEYINPUT25), .A2(n1147), .ZN(n1145) );
XOR2_X1 U830 ( .A(n1148), .B(n1149), .Z(n1141) );
NOR3_X1 U831 ( .A1(n1138), .A2(KEYINPUT56), .A3(n1150), .ZN(n1149) );
NAND2_X1 U832 ( .A1(G902), .A2(n1000), .ZN(n1138) );
OR3_X1 U833 ( .A1(n1090), .A2(n1151), .A3(n1075), .ZN(n1000) );
NAND4_X1 U834 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1075) );
NOR4_X1 U835 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
NOR2_X1 U836 ( .A1(n1160), .A2(n1161), .ZN(n1154) );
NAND3_X1 U837 ( .A1(n1031), .A2(n1162), .A3(n1163), .ZN(n1152) );
XOR2_X1 U838 ( .A(KEYINPUT1), .B(n1164), .Z(n1162) );
XNOR2_X1 U839 ( .A(KEYINPUT38), .B(n1165), .ZN(n1151) );
AND4_X1 U840 ( .A1(n1092), .A2(n1091), .A3(n1093), .A4(n1166), .ZN(n1165) );
XNOR2_X1 U841 ( .A(KEYINPUT39), .B(n1089), .ZN(n1166) );
NAND3_X1 U842 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1092) );
XNOR2_X1 U843 ( .A(KEYINPUT45), .B(n1014), .ZN(n1168) );
INV_X1 U844 ( .A(n1170), .ZN(n1014) );
NAND4_X1 U845 ( .A1(n1108), .A2(n1171), .A3(n1172), .A4(n995), .ZN(n1090) );
NAND3_X1 U846 ( .A1(n1030), .A2(n1032), .A3(n1173), .ZN(n995) );
NAND3_X1 U847 ( .A1(n1173), .A2(n1032), .A3(n1031), .ZN(n1108) );
XOR2_X1 U848 ( .A(n1174), .B(KEYINPUT34), .Z(n1148) );
NOR2_X1 U849 ( .A1(n1074), .A2(G952), .ZN(n1094) );
XNOR2_X1 U850 ( .A(G146), .B(n1175), .ZN(G48) );
NAND4_X1 U851 ( .A1(KEYINPUT53), .A2(n1164), .A3(n1163), .A4(n1031), .ZN(n1175) );
NAND2_X1 U852 ( .A1(n1176), .A2(n1177), .ZN(G45) );
NAND2_X1 U853 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XOR2_X1 U854 ( .A(n1180), .B(KEYINPUT42), .Z(n1176) );
OR2_X1 U855 ( .A1(n1179), .A2(n1178), .ZN(n1180) );
INV_X1 U856 ( .A(n1153), .ZN(n1178) );
NAND4_X1 U857 ( .A1(n1163), .A2(n1026), .A3(n1181), .A4(n1182), .ZN(n1153) );
XOR2_X1 U858 ( .A(G143), .B(KEYINPUT20), .Z(n1179) );
XNOR2_X1 U859 ( .A(n1137), .B(n1161), .ZN(G42) );
AND2_X1 U860 ( .A1(n1183), .A2(n1184), .ZN(n1161) );
NAND3_X1 U861 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(G39) );
NAND2_X1 U862 ( .A1(n1160), .A2(n1073), .ZN(n1187) );
INV_X1 U863 ( .A(n1188), .ZN(n1160) );
NAND2_X1 U864 ( .A1(KEYINPUT40), .A2(n1189), .ZN(n1186) );
NAND2_X1 U865 ( .A1(G137), .A2(n1190), .ZN(n1189) );
XNOR2_X1 U866 ( .A(KEYINPUT3), .B(n1188), .ZN(n1190) );
NAND2_X1 U867 ( .A1(n1191), .A2(n1192), .ZN(n1185) );
INV_X1 U868 ( .A(KEYINPUT40), .ZN(n1192) );
NAND2_X1 U869 ( .A1(n1193), .A2(n1194), .ZN(n1191) );
NAND3_X1 U870 ( .A1(KEYINPUT3), .A2(G137), .A3(n1188), .ZN(n1194) );
OR2_X1 U871 ( .A1(n1188), .A2(KEYINPUT3), .ZN(n1193) );
NAND2_X1 U872 ( .A1(n1169), .A2(n1184), .ZN(n1188) );
INV_X1 U873 ( .A(n1195), .ZN(n1169) );
XNOR2_X1 U874 ( .A(n1196), .B(n1157), .ZN(G36) );
AND3_X1 U875 ( .A1(n1184), .A2(n1030), .A3(n1026), .ZN(n1157) );
XNOR2_X1 U876 ( .A(n1071), .B(n1156), .ZN(G33) );
AND3_X1 U877 ( .A1(n1184), .A2(n1031), .A3(n1026), .ZN(n1156) );
AND3_X1 U878 ( .A1(n1197), .A2(n1019), .A3(n1010), .ZN(n1184) );
AND3_X1 U879 ( .A1(n1016), .A2(n1017), .A3(n1013), .ZN(n1010) );
INV_X1 U880 ( .A(n1015), .ZN(n1013) );
XOR2_X1 U881 ( .A(G128), .B(n1159), .Z(G30) );
AND3_X1 U882 ( .A1(n1163), .A2(n1030), .A3(n1164), .ZN(n1159) );
AND3_X1 U883 ( .A1(n1016), .A2(n1017), .A3(n1198), .ZN(n1163) );
XNOR2_X1 U884 ( .A(G101), .B(n1171), .ZN(G3) );
NAND3_X1 U885 ( .A1(n1026), .A2(n1173), .A3(n1024), .ZN(n1171) );
XOR2_X1 U886 ( .A(G125), .B(n1158), .Z(G27) );
AND3_X1 U887 ( .A1(n1183), .A2(n1198), .A3(n1170), .ZN(n1158) );
AND3_X1 U888 ( .A1(n1197), .A2(n1019), .A3(n1015), .ZN(n1198) );
NAND2_X1 U889 ( .A1(n1002), .A2(n1199), .ZN(n1197) );
NAND4_X1 U890 ( .A1(G902), .A2(G953), .A3(n1200), .A4(n1201), .ZN(n1199) );
INV_X1 U891 ( .A(G900), .ZN(n1201) );
AND3_X1 U892 ( .A1(n1028), .A2(n1027), .A3(n1031), .ZN(n1183) );
XNOR2_X1 U893 ( .A(G122), .B(n1093), .ZN(G24) );
NAND4_X1 U894 ( .A1(n1202), .A2(n1032), .A3(n1181), .A4(n1182), .ZN(n1093) );
INV_X1 U895 ( .A(n1007), .ZN(n1032) );
NAND2_X1 U896 ( .A1(n1203), .A2(n1028), .ZN(n1007) );
XOR2_X1 U897 ( .A(G119), .B(n1204), .Z(G21) );
NOR2_X1 U898 ( .A1(n1195), .A2(n1205), .ZN(n1204) );
NAND2_X1 U899 ( .A1(n1024), .A2(n1164), .ZN(n1195) );
NOR2_X1 U900 ( .A1(n1028), .A2(n1203), .ZN(n1164) );
INV_X1 U901 ( .A(n1027), .ZN(n1203) );
XOR2_X1 U902 ( .A(n1206), .B(n1207), .Z(G18) );
XOR2_X1 U903 ( .A(KEYINPUT47), .B(G116), .Z(n1207) );
NOR2_X1 U904 ( .A1(KEYINPUT27), .A2(n1091), .ZN(n1206) );
NAND3_X1 U905 ( .A1(n1026), .A2(n1030), .A3(n1202), .ZN(n1091) );
AND2_X1 U906 ( .A1(n1208), .A2(n1182), .ZN(n1030) );
XNOR2_X1 U907 ( .A(n1089), .B(n1209), .ZN(G15) );
XOR2_X1 U908 ( .A(KEYINPUT4), .B(G113), .Z(n1209) );
AND3_X1 U909 ( .A1(n1026), .A2(n1031), .A3(n1202), .ZN(n1089) );
INV_X1 U910 ( .A(n1205), .ZN(n1202) );
NAND2_X1 U911 ( .A1(n1170), .A2(n1167), .ZN(n1205) );
NOR2_X1 U912 ( .A1(n1016), .A2(n1036), .ZN(n1170) );
INV_X1 U913 ( .A(n1017), .ZN(n1036) );
NOR2_X1 U914 ( .A1(n1182), .A2(n1208), .ZN(n1031) );
INV_X1 U915 ( .A(n1181), .ZN(n1208) );
NOR2_X1 U916 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
XNOR2_X1 U917 ( .A(G110), .B(n1172), .ZN(G12) );
NAND4_X1 U918 ( .A1(n1024), .A2(n1173), .A3(n1028), .A4(n1027), .ZN(n1172) );
NAND3_X1 U919 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1027) );
NAND2_X1 U920 ( .A1(n1213), .A2(n1097), .ZN(n1212) );
OR3_X1 U921 ( .A1(n1097), .A2(n1213), .A3(G902), .ZN(n1211) );
NOR2_X1 U922 ( .A1(n1214), .A2(G234), .ZN(n1213) );
INV_X1 U923 ( .A(G217), .ZN(n1214) );
XOR2_X1 U924 ( .A(n1215), .B(n1216), .Z(n1097) );
XOR2_X1 U925 ( .A(n1217), .B(n1218), .Z(n1216) );
XOR2_X1 U926 ( .A(G110), .B(n1219), .Z(n1218) );
AND3_X1 U927 ( .A1(G221), .A2(n1074), .A3(G234), .ZN(n1219) );
XOR2_X1 U928 ( .A(KEYINPUT55), .B(G119), .Z(n1217) );
XNOR2_X1 U929 ( .A(n1220), .B(n1221), .ZN(n1215) );
XOR2_X1 U930 ( .A(n1222), .B(n1223), .Z(n1220) );
NOR2_X1 U931 ( .A1(KEYINPUT23), .A2(n1137), .ZN(n1223) );
NAND2_X1 U932 ( .A1(G217), .A2(G902), .ZN(n1210) );
XOR2_X1 U933 ( .A(n1224), .B(G472), .Z(n1028) );
NAND2_X1 U934 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U935 ( .A(n1227), .B(n1228), .Z(n1225) );
XOR2_X1 U936 ( .A(KEYINPUT12), .B(n1229), .Z(n1228) );
NOR2_X1 U937 ( .A1(KEYINPUT30), .A2(n1230), .ZN(n1229) );
XNOR2_X1 U938 ( .A(n1123), .B(n1231), .ZN(n1230) );
NOR2_X1 U939 ( .A1(KEYINPUT63), .A2(n1125), .ZN(n1231) );
INV_X1 U940 ( .A(G101), .ZN(n1125) );
NAND2_X1 U941 ( .A1(n1232), .A2(G210), .ZN(n1123) );
XNOR2_X1 U942 ( .A(n1122), .B(n1119), .ZN(n1227) );
XOR2_X1 U943 ( .A(n1233), .B(n1234), .Z(n1119) );
INV_X1 U944 ( .A(n1235), .ZN(n1234) );
NAND2_X1 U945 ( .A1(KEYINPUT18), .A2(G113), .ZN(n1233) );
XOR2_X1 U946 ( .A(n1236), .B(n1237), .Z(n1122) );
XOR2_X1 U947 ( .A(n1222), .B(n1238), .Z(n1236) );
XNOR2_X1 U948 ( .A(G137), .B(n1239), .ZN(n1222) );
AND3_X1 U949 ( .A1(n1016), .A2(n1017), .A3(n1167), .ZN(n1173) );
AND3_X1 U950 ( .A1(n1240), .A2(n1019), .A3(n1015), .ZN(n1167) );
XOR2_X1 U951 ( .A(n1049), .B(KEYINPUT31), .Z(n1015) );
XOR2_X1 U952 ( .A(n1241), .B(n1150), .Z(n1049) );
NAND2_X1 U953 ( .A1(G210), .A2(n1242), .ZN(n1150) );
NAND2_X1 U954 ( .A1(n1243), .A2(n1226), .ZN(n1241) );
XOR2_X1 U955 ( .A(n1244), .B(n1245), .Z(n1243) );
XNOR2_X1 U956 ( .A(n1147), .B(n1246), .ZN(n1245) );
NOR2_X1 U957 ( .A1(KEYINPUT52), .A2(n1247), .ZN(n1246) );
XNOR2_X1 U958 ( .A(n1063), .B(n1143), .ZN(n1247) );
XNOR2_X1 U959 ( .A(n1237), .B(n1239), .ZN(n1143) );
XOR2_X1 U960 ( .A(G128), .B(G146), .Z(n1239) );
XNOR2_X1 U961 ( .A(G143), .B(KEYINPUT37), .ZN(n1237) );
AND2_X1 U962 ( .A1(n1248), .A2(n1249), .ZN(n1147) );
NAND2_X1 U963 ( .A1(n1250), .A2(n1083), .ZN(n1249) );
INV_X1 U964 ( .A(n1251), .ZN(n1083) );
XNOR2_X1 U965 ( .A(KEYINPUT49), .B(n1252), .ZN(n1250) );
NAND2_X1 U966 ( .A1(n1253), .A2(n1251), .ZN(n1248) );
XOR2_X1 U967 ( .A(n1235), .B(n1254), .Z(n1251) );
NOR2_X1 U968 ( .A1(G113), .A2(KEYINPUT50), .ZN(n1254) );
XOR2_X1 U969 ( .A(G116), .B(G119), .Z(n1235) );
XNOR2_X1 U970 ( .A(KEYINPUT51), .B(n1252), .ZN(n1253) );
INV_X1 U971 ( .A(n1082), .ZN(n1252) );
XNOR2_X1 U972 ( .A(n1255), .B(G122), .ZN(n1082) );
XNOR2_X1 U973 ( .A(n1256), .B(n1174), .ZN(n1244) );
NAND2_X1 U974 ( .A1(G224), .A2(n1074), .ZN(n1174) );
XNOR2_X1 U975 ( .A(KEYINPUT59), .B(KEYINPUT46), .ZN(n1256) );
NAND2_X1 U976 ( .A1(G214), .A2(n1242), .ZN(n1019) );
NAND2_X1 U977 ( .A1(n1257), .A2(n1226), .ZN(n1242) );
INV_X1 U978 ( .A(G237), .ZN(n1257) );
NAND2_X1 U979 ( .A1(n1258), .A2(n1002), .ZN(n1240) );
NAND3_X1 U980 ( .A1(n1200), .A2(n1074), .A3(G952), .ZN(n1002) );
XOR2_X1 U981 ( .A(n1259), .B(KEYINPUT41), .Z(n1258) );
NAND3_X1 U982 ( .A1(n1084), .A2(n1200), .A3(G902), .ZN(n1259) );
NAND2_X1 U983 ( .A1(G237), .A2(G234), .ZN(n1200) );
NOR2_X1 U984 ( .A1(n1074), .A2(G898), .ZN(n1084) );
NAND2_X1 U985 ( .A1(G221), .A2(n1260), .ZN(n1017) );
NAND2_X1 U986 ( .A1(G234), .A2(n1226), .ZN(n1260) );
XOR2_X1 U987 ( .A(n1047), .B(G469), .Z(n1016) );
INV_X1 U988 ( .A(n1045), .ZN(n1047) );
NAND2_X1 U989 ( .A1(n1261), .A2(n1226), .ZN(n1045) );
XOR2_X1 U990 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U991 ( .A(n1264), .B(n1265), .Z(n1263) );
XNOR2_X1 U992 ( .A(n1266), .B(n1137), .ZN(n1265) );
NAND2_X1 U993 ( .A1(KEYINPUT8), .A2(n1064), .ZN(n1266) );
XNOR2_X1 U994 ( .A(n1267), .B(G128), .ZN(n1064) );
NAND2_X1 U995 ( .A1(KEYINPUT62), .A2(n1268), .ZN(n1267) );
XNOR2_X1 U996 ( .A(n1269), .B(G143), .ZN(n1268) );
NAND2_X1 U997 ( .A1(KEYINPUT14), .A2(n1135), .ZN(n1264) );
NOR2_X1 U998 ( .A1(n1054), .A2(G953), .ZN(n1135) );
INV_X1 U999 ( .A(G227), .ZN(n1054) );
XOR2_X1 U1000 ( .A(n1255), .B(n1133), .Z(n1262) );
XNOR2_X1 U1001 ( .A(n1073), .B(n1238), .ZN(n1133) );
XNOR2_X1 U1002 ( .A(n1270), .B(n1271), .ZN(n1238) );
NOR2_X1 U1003 ( .A1(KEYINPUT36), .A2(n1071), .ZN(n1271) );
NAND2_X1 U1004 ( .A1(KEYINPUT43), .A2(n1196), .ZN(n1270) );
INV_X1 U1005 ( .A(G134), .ZN(n1196) );
INV_X1 U1006 ( .A(G137), .ZN(n1073) );
XOR2_X1 U1007 ( .A(n1139), .B(G110), .Z(n1255) );
XNOR2_X1 U1008 ( .A(G101), .B(n1272), .ZN(n1139) );
XNOR2_X1 U1009 ( .A(G107), .B(n1110), .ZN(n1272) );
NOR2_X1 U1010 ( .A1(n1182), .A2(n1181), .ZN(n1024) );
XNOR2_X1 U1011 ( .A(n1040), .B(n1273), .ZN(n1181) );
XOR2_X1 U1012 ( .A(KEYINPUT5), .B(G475), .Z(n1273) );
NAND2_X1 U1013 ( .A1(n1106), .A2(n1226), .ZN(n1040) );
INV_X1 U1014 ( .A(G902), .ZN(n1226) );
XNOR2_X1 U1015 ( .A(n1274), .B(KEYINPUT57), .ZN(n1106) );
XOR2_X1 U1016 ( .A(n1275), .B(n1276), .Z(n1274) );
XOR2_X1 U1017 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U1018 ( .A(G122), .B(G113), .Z(n1278) );
XNOR2_X1 U1019 ( .A(G143), .B(n1071), .ZN(n1277) );
INV_X1 U1020 ( .A(G131), .ZN(n1071) );
XOR2_X1 U1021 ( .A(n1279), .B(n1280), .Z(n1275) );
XOR2_X1 U1022 ( .A(n1281), .B(n1282), .Z(n1280) );
NAND2_X1 U1023 ( .A1(KEYINPUT60), .A2(n1269), .ZN(n1282) );
INV_X1 U1024 ( .A(G146), .ZN(n1269) );
NAND3_X1 U1025 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1281) );
NAND2_X1 U1026 ( .A1(G140), .A2(n1221), .ZN(n1285) );
INV_X1 U1027 ( .A(n1063), .ZN(n1221) );
NAND2_X1 U1028 ( .A1(KEYINPUT19), .A2(n1286), .ZN(n1284) );
NAND2_X1 U1029 ( .A1(n1287), .A2(n1137), .ZN(n1286) );
XNOR2_X1 U1030 ( .A(KEYINPUT21), .B(n1063), .ZN(n1287) );
NAND2_X1 U1031 ( .A1(n1288), .A2(n1289), .ZN(n1283) );
INV_X1 U1032 ( .A(KEYINPUT19), .ZN(n1289) );
NAND2_X1 U1033 ( .A1(n1290), .A2(n1291), .ZN(n1288) );
OR2_X1 U1034 ( .A1(n1063), .A2(KEYINPUT21), .ZN(n1291) );
NAND3_X1 U1035 ( .A1(n1063), .A2(n1137), .A3(KEYINPUT21), .ZN(n1290) );
INV_X1 U1036 ( .A(G140), .ZN(n1137) );
XOR2_X1 U1037 ( .A(G125), .B(KEYINPUT0), .Z(n1063) );
XOR2_X1 U1038 ( .A(n1292), .B(n1293), .Z(n1279) );
AND2_X1 U1039 ( .A1(G214), .A2(n1232), .ZN(n1293) );
NOR2_X1 U1040 ( .A1(G953), .A2(G237), .ZN(n1232) );
NAND2_X1 U1041 ( .A1(KEYINPUT28), .A2(n1110), .ZN(n1292) );
INV_X1 U1042 ( .A(G104), .ZN(n1110) );
XOR2_X1 U1043 ( .A(n1041), .B(G478), .Z(n1182) );
NOR2_X1 U1044 ( .A1(n1102), .A2(G902), .ZN(n1041) );
XOR2_X1 U1045 ( .A(n1294), .B(n1295), .Z(n1102) );
XOR2_X1 U1046 ( .A(n1296), .B(n1297), .Z(n1295) );
XNOR2_X1 U1047 ( .A(n1298), .B(n1299), .ZN(n1297) );
NOR2_X1 U1048 ( .A1(G134), .A2(KEYINPUT26), .ZN(n1299) );
NAND2_X1 U1049 ( .A1(KEYINPUT6), .A2(n1300), .ZN(n1298) );
XOR2_X1 U1050 ( .A(G122), .B(G116), .Z(n1300) );
NOR2_X1 U1051 ( .A1(G128), .A2(KEYINPUT15), .ZN(n1296) );
XOR2_X1 U1052 ( .A(n1301), .B(n1302), .Z(n1294) );
XOR2_X1 U1053 ( .A(G143), .B(G107), .Z(n1302) );
NAND3_X1 U1054 ( .A1(G234), .A2(n1074), .A3(G217), .ZN(n1301) );
INV_X1 U1055 ( .A(G953), .ZN(n1074) );
endmodule


