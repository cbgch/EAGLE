//Key = 0000100100110000001110101011111001100101111101001000000101110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413;

XOR2_X1 U783 ( .A(n1087), .B(n1088), .Z(G9) );
NAND2_X1 U784 ( .A1(KEYINPUT18), .A2(G107), .ZN(n1088) );
OR2_X1 U785 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR2_X1 U786 ( .A1(n1091), .A2(n1092), .ZN(G75) );
NOR4_X1 U787 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1092) );
XNOR2_X1 U788 ( .A(n1097), .B(KEYINPUT44), .ZN(n1096) );
NOR2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
NOR2_X1 U790 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
XOR2_X1 U791 ( .A(KEYINPUT53), .B(n1102), .Z(n1101) );
AND4_X1 U792 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1102) );
NOR2_X1 U793 ( .A1(n1107), .A2(n1108), .ZN(n1100) );
NOR2_X1 U794 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
NOR2_X1 U795 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
INV_X1 U796 ( .A(n1105), .ZN(n1112) );
NOR2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U799 ( .A1(n1117), .A2(n1118), .ZN(n1115) );
NOR2_X1 U800 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NOR2_X1 U801 ( .A1(n1121), .A2(n1122), .ZN(n1113) );
XNOR2_X1 U802 ( .A(n1123), .B(KEYINPUT43), .ZN(n1122) );
NOR3_X1 U803 ( .A1(n1121), .A2(n1124), .A3(n1116), .ZN(n1109) );
NOR2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND3_X1 U805 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1093) );
NAND4_X1 U806 ( .A1(n1106), .A2(n1105), .A3(n1130), .A4(n1131), .ZN(n1129) );
NAND3_X1 U807 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
NAND2_X1 U808 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
INV_X1 U809 ( .A(KEYINPUT62), .ZN(n1136) );
NAND3_X1 U810 ( .A1(KEYINPUT62), .A2(n1137), .A3(n1121), .ZN(n1133) );
NAND3_X1 U811 ( .A1(n1138), .A2(n1139), .A3(n1103), .ZN(n1132) );
INV_X1 U812 ( .A(n1108), .ZN(n1106) );
AND3_X1 U813 ( .A1(n1127), .A2(n1128), .A3(n1140), .ZN(n1091) );
NAND4_X1 U814 ( .A1(n1141), .A2(n1103), .A3(n1142), .A4(n1143), .ZN(n1127) );
NOR4_X1 U815 ( .A1(n1138), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1143) );
XOR2_X1 U816 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U817 ( .A1(G472), .A2(KEYINPUT25), .ZN(n1148) );
XOR2_X1 U818 ( .A(n1139), .B(KEYINPUT58), .Z(n1145) );
XNOR2_X1 U819 ( .A(n1149), .B(n1150), .ZN(n1144) );
NOR2_X1 U820 ( .A1(G475), .A2(KEYINPUT3), .ZN(n1150) );
XNOR2_X1 U821 ( .A(n1151), .B(G478), .ZN(n1142) );
XOR2_X1 U822 ( .A(n1152), .B(n1153), .Z(G72) );
XOR2_X1 U823 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U824 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XNOR2_X1 U825 ( .A(KEYINPUT21), .B(n1128), .ZN(n1157) );
NAND2_X1 U826 ( .A1(n1158), .A2(n1159), .ZN(n1154) );
INV_X1 U827 ( .A(n1160), .ZN(n1159) );
XOR2_X1 U828 ( .A(n1161), .B(n1162), .Z(n1158) );
XOR2_X1 U829 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U830 ( .A1(KEYINPUT38), .A2(n1165), .ZN(n1164) );
XNOR2_X1 U831 ( .A(G131), .B(n1166), .ZN(n1161) );
NOR2_X1 U832 ( .A1(KEYINPUT35), .A2(n1167), .ZN(n1166) );
XNOR2_X1 U833 ( .A(G134), .B(G137), .ZN(n1167) );
NAND2_X1 U834 ( .A1(G953), .A2(n1168), .ZN(n1152) );
NAND2_X1 U835 ( .A1(G900), .A2(G227), .ZN(n1168) );
XOR2_X1 U836 ( .A(n1169), .B(n1170), .Z(G69) );
NAND2_X1 U837 ( .A1(G953), .A2(n1171), .ZN(n1170) );
NAND2_X1 U838 ( .A1(G898), .A2(G224), .ZN(n1171) );
NAND2_X1 U839 ( .A1(KEYINPUT10), .A2(n1172), .ZN(n1169) );
XOR2_X1 U840 ( .A(n1173), .B(n1174), .Z(n1172) );
NAND2_X1 U841 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND2_X1 U842 ( .A1(G953), .A2(n1177), .ZN(n1176) );
XOR2_X1 U843 ( .A(n1178), .B(n1179), .Z(n1175) );
NAND2_X1 U844 ( .A1(KEYINPUT28), .A2(n1180), .ZN(n1178) );
NAND3_X1 U845 ( .A1(n1181), .A2(n1182), .A3(n1128), .ZN(n1173) );
OR3_X1 U846 ( .A1(n1183), .A2(n1184), .A3(KEYINPUT27), .ZN(n1182) );
NAND2_X1 U847 ( .A1(KEYINPUT27), .A2(n1097), .ZN(n1181) );
NOR3_X1 U848 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(G66) );
AND2_X1 U849 ( .A1(KEYINPUT37), .A2(n1188), .ZN(n1187) );
NOR3_X1 U850 ( .A1(KEYINPUT37), .A2(G953), .A3(G952), .ZN(n1186) );
XOR2_X1 U851 ( .A(n1189), .B(n1190), .Z(n1185) );
NAND2_X1 U852 ( .A1(n1191), .A2(n1192), .ZN(n1189) );
NOR3_X1 U853 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(G63) );
NOR3_X1 U854 ( .A1(n1196), .A2(n1128), .A3(n1140), .ZN(n1195) );
INV_X1 U855 ( .A(G952), .ZN(n1140) );
AND2_X1 U856 ( .A1(n1196), .A2(n1188), .ZN(n1194) );
INV_X1 U857 ( .A(KEYINPUT32), .ZN(n1196) );
NOR3_X1 U858 ( .A1(n1151), .A2(n1197), .A3(n1198), .ZN(n1193) );
AND3_X1 U859 ( .A1(n1199), .A2(G478), .A3(n1191), .ZN(n1198) );
NOR2_X1 U860 ( .A1(n1200), .A2(n1199), .ZN(n1197) );
NOR2_X1 U861 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
INV_X1 U862 ( .A(G478), .ZN(n1202) );
NOR2_X1 U863 ( .A1(n1188), .A2(n1203), .ZN(G60) );
NOR3_X1 U864 ( .A1(n1149), .A2(n1204), .A3(n1205), .ZN(n1203) );
AND3_X1 U865 ( .A1(n1206), .A2(n1191), .A3(G475), .ZN(n1205) );
NOR2_X1 U866 ( .A1(n1207), .A2(n1206), .ZN(n1204) );
NOR2_X1 U867 ( .A1(n1201), .A2(n1208), .ZN(n1207) );
INV_X1 U868 ( .A(G475), .ZN(n1208) );
NOR2_X1 U869 ( .A1(n1209), .A2(n1094), .ZN(n1201) );
INV_X1 U870 ( .A(n1097), .ZN(n1209) );
XOR2_X1 U871 ( .A(G104), .B(n1210), .Z(G6) );
NOR2_X1 U872 ( .A1(n1188), .A2(n1211), .ZN(G57) );
XOR2_X1 U873 ( .A(n1212), .B(n1213), .Z(n1211) );
XNOR2_X1 U874 ( .A(n1214), .B(n1215), .ZN(n1213) );
NAND2_X1 U875 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U876 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
INV_X1 U877 ( .A(KEYINPUT15), .ZN(n1219) );
NAND2_X1 U878 ( .A1(n1220), .A2(KEYINPUT15), .ZN(n1216) );
XOR2_X1 U879 ( .A(n1221), .B(n1222), .Z(n1212) );
NAND2_X1 U880 ( .A1(n1191), .A2(G472), .ZN(n1221) );
NOR2_X1 U881 ( .A1(n1188), .A2(n1223), .ZN(G54) );
XOR2_X1 U882 ( .A(n1224), .B(n1225), .Z(n1223) );
XOR2_X1 U883 ( .A(n1226), .B(n1227), .Z(n1225) );
NAND2_X1 U884 ( .A1(n1191), .A2(G469), .ZN(n1226) );
XOR2_X1 U885 ( .A(n1228), .B(n1229), .Z(n1224) );
XNOR2_X1 U886 ( .A(n1230), .B(n1163), .ZN(n1229) );
NAND2_X1 U887 ( .A1(KEYINPUT45), .A2(n1231), .ZN(n1230) );
NAND2_X1 U888 ( .A1(n1232), .A2(KEYINPUT34), .ZN(n1228) );
XNOR2_X1 U889 ( .A(n1233), .B(n1234), .ZN(n1232) );
XOR2_X1 U890 ( .A(KEYINPUT4), .B(KEYINPUT0), .Z(n1234) );
NOR2_X1 U891 ( .A1(n1188), .A2(n1235), .ZN(G51) );
XOR2_X1 U892 ( .A(n1236), .B(n1237), .Z(n1235) );
NAND2_X1 U893 ( .A1(n1191), .A2(G210), .ZN(n1237) );
AND2_X1 U894 ( .A1(G902), .A2(n1238), .ZN(n1191) );
NAND2_X1 U895 ( .A1(n1156), .A2(n1097), .ZN(n1238) );
NOR2_X1 U896 ( .A1(n1184), .A2(n1239), .ZN(n1097) );
NAND4_X1 U897 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1184) );
AND3_X1 U898 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1243) );
NAND2_X1 U899 ( .A1(KEYINPUT7), .A2(n1210), .ZN(n1242) );
AND4_X1 U900 ( .A1(n1126), .A2(n1137), .A3(n1130), .A4(n1247), .ZN(n1210) );
NAND3_X1 U901 ( .A1(n1125), .A2(n1248), .A3(n1249), .ZN(n1241) );
NAND2_X1 U902 ( .A1(n1137), .A2(n1250), .ZN(n1240) );
NAND2_X1 U903 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U904 ( .A1(n1247), .A2(n1253), .ZN(n1252) );
NAND2_X1 U905 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
OR3_X1 U906 ( .A1(n1126), .A2(KEYINPUT7), .A3(n1116), .ZN(n1255) );
INV_X1 U907 ( .A(n1130), .ZN(n1116) );
NAND2_X1 U908 ( .A1(n1105), .A2(n1104), .ZN(n1254) );
XOR2_X1 U909 ( .A(n1090), .B(KEYINPUT8), .Z(n1251) );
NAND3_X1 U910 ( .A1(n1125), .A2(n1247), .A3(n1130), .ZN(n1090) );
INV_X1 U911 ( .A(n1094), .ZN(n1156) );
NAND4_X1 U912 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1094) );
NOR4_X1 U913 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(n1259) );
NOR3_X1 U914 ( .A1(n1264), .A2(n1089), .A3(n1265), .ZN(n1263) );
NOR2_X1 U915 ( .A1(n1266), .A2(n1267), .ZN(n1258) );
INV_X1 U916 ( .A(n1268), .ZN(n1266) );
NAND2_X1 U917 ( .A1(n1269), .A2(n1270), .ZN(n1236) );
NAND2_X1 U918 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XOR2_X1 U919 ( .A(n1273), .B(KEYINPUT56), .Z(n1269) );
OR2_X1 U920 ( .A1(n1272), .A2(n1271), .ZN(n1273) );
XNOR2_X1 U921 ( .A(n1274), .B(n1275), .ZN(n1272) );
XOR2_X1 U922 ( .A(n1276), .B(n1277), .Z(n1274) );
NOR2_X1 U923 ( .A1(n1128), .A2(G952), .ZN(n1188) );
XOR2_X1 U924 ( .A(n1278), .B(n1261), .Z(G48) );
AND3_X1 U925 ( .A1(n1126), .A2(n1137), .A3(n1279), .ZN(n1261) );
XNOR2_X1 U926 ( .A(G146), .B(KEYINPUT59), .ZN(n1278) );
XNOR2_X1 U927 ( .A(G143), .B(n1280), .ZN(G45) );
NAND3_X1 U928 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1280) );
XNOR2_X1 U929 ( .A(n1137), .B(KEYINPUT41), .ZN(n1283) );
XOR2_X1 U930 ( .A(G140), .B(n1260), .Z(G42) );
AND3_X1 U931 ( .A1(n1284), .A2(n1118), .A3(n1285), .ZN(n1260) );
XNOR2_X1 U932 ( .A(G137), .B(n1256), .ZN(G39) );
NAND3_X1 U933 ( .A1(n1285), .A2(n1279), .A3(n1105), .ZN(n1256) );
NAND2_X1 U934 ( .A1(n1286), .A2(n1287), .ZN(G36) );
NAND2_X1 U935 ( .A1(G134), .A2(n1257), .ZN(n1287) );
XOR2_X1 U936 ( .A(KEYINPUT26), .B(n1288), .Z(n1286) );
NOR2_X1 U937 ( .A1(G134), .A2(n1257), .ZN(n1288) );
NAND3_X1 U938 ( .A1(n1282), .A2(n1265), .A3(n1285), .ZN(n1257) );
INV_X1 U939 ( .A(n1264), .ZN(n1282) );
NAND2_X1 U940 ( .A1(n1289), .A2(n1290), .ZN(n1264) );
XOR2_X1 U941 ( .A(G131), .B(n1262), .Z(G33) );
AND3_X1 U942 ( .A1(n1289), .A2(n1126), .A3(n1285), .ZN(n1262) );
INV_X1 U943 ( .A(n1099), .ZN(n1285) );
NAND2_X1 U944 ( .A1(n1139), .A2(n1291), .ZN(n1099) );
AND3_X1 U945 ( .A1(n1248), .A2(n1292), .A3(n1118), .ZN(n1289) );
XOR2_X1 U946 ( .A(G128), .B(n1267), .Z(G30) );
AND3_X1 U947 ( .A1(n1137), .A2(n1125), .A3(n1279), .ZN(n1267) );
AND4_X1 U948 ( .A1(n1118), .A2(n1293), .A3(n1294), .A4(n1292), .ZN(n1279) );
NAND2_X1 U949 ( .A1(n1295), .A2(n1296), .ZN(G3) );
NAND2_X1 U950 ( .A1(G101), .A2(n1244), .ZN(n1296) );
XOR2_X1 U951 ( .A(KEYINPUT61), .B(n1297), .Z(n1295) );
NOR2_X1 U952 ( .A1(G101), .A2(n1244), .ZN(n1297) );
NAND4_X1 U953 ( .A1(n1105), .A2(n1137), .A3(n1247), .A4(n1248), .ZN(n1244) );
XNOR2_X1 U954 ( .A(G125), .B(n1268), .ZN(G27) );
NAND2_X1 U955 ( .A1(n1135), .A2(n1284), .ZN(n1268) );
AND3_X1 U956 ( .A1(n1104), .A2(n1292), .A3(n1126), .ZN(n1284) );
NAND2_X1 U957 ( .A1(n1108), .A2(n1298), .ZN(n1292) );
NAND3_X1 U958 ( .A1(G902), .A2(n1299), .A3(n1160), .ZN(n1298) );
NOR2_X1 U959 ( .A1(n1128), .A2(G900), .ZN(n1160) );
XOR2_X1 U960 ( .A(n1246), .B(n1300), .Z(G24) );
NOR2_X1 U961 ( .A1(G122), .A2(KEYINPUT16), .ZN(n1300) );
NAND4_X1 U962 ( .A1(n1281), .A2(n1249), .A3(n1290), .A4(n1130), .ZN(n1246) );
XOR2_X1 U963 ( .A(G119), .B(n1239), .Z(G21) );
INV_X1 U964 ( .A(n1183), .ZN(n1239) );
NAND4_X1 U965 ( .A1(n1249), .A2(n1105), .A3(n1293), .A4(n1294), .ZN(n1183) );
NAND3_X1 U966 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(G18) );
NAND2_X1 U967 ( .A1(G116), .A2(n1304), .ZN(n1303) );
NAND2_X1 U968 ( .A1(KEYINPUT14), .A2(n1305), .ZN(n1302) );
NAND2_X1 U969 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XNOR2_X1 U970 ( .A(KEYINPUT13), .B(n1304), .ZN(n1306) );
NAND2_X1 U971 ( .A1(n1308), .A2(n1309), .ZN(n1301) );
INV_X1 U972 ( .A(KEYINPUT14), .ZN(n1309) );
NAND2_X1 U973 ( .A1(n1310), .A2(n1311), .ZN(n1308) );
NAND2_X1 U974 ( .A1(KEYINPUT13), .A2(n1304), .ZN(n1311) );
OR3_X1 U975 ( .A1(G116), .A2(KEYINPUT13), .A3(n1304), .ZN(n1310) );
NAND3_X1 U976 ( .A1(n1103), .A2(n1125), .A3(n1312), .ZN(n1304) );
NOR3_X1 U977 ( .A1(n1313), .A2(n1123), .A3(n1314), .ZN(n1312) );
XOR2_X1 U978 ( .A(n1315), .B(KEYINPUT22), .Z(n1314) );
INV_X1 U979 ( .A(n1248), .ZN(n1123) );
XNOR2_X1 U980 ( .A(n1137), .B(KEYINPUT31), .ZN(n1313) );
AND2_X1 U981 ( .A1(n1290), .A2(n1265), .ZN(n1125) );
INV_X1 U982 ( .A(n1121), .ZN(n1103) );
XNOR2_X1 U983 ( .A(n1245), .B(n1316), .ZN(G15) );
NOR2_X1 U984 ( .A1(KEYINPUT60), .A2(n1317), .ZN(n1316) );
NAND3_X1 U985 ( .A1(n1126), .A2(n1248), .A3(n1249), .ZN(n1245) );
AND2_X1 U986 ( .A1(n1135), .A2(n1315), .ZN(n1249) );
NOR2_X1 U987 ( .A1(n1121), .A2(n1089), .ZN(n1135) );
NAND2_X1 U988 ( .A1(n1318), .A2(n1120), .ZN(n1121) );
INV_X1 U989 ( .A(n1119), .ZN(n1318) );
NAND2_X1 U990 ( .A1(n1319), .A2(n1320), .ZN(n1248) );
NAND3_X1 U991 ( .A1(n1294), .A2(n1141), .A3(n1321), .ZN(n1320) );
INV_X1 U992 ( .A(KEYINPUT46), .ZN(n1321) );
NAND2_X1 U993 ( .A1(KEYINPUT46), .A2(n1130), .ZN(n1319) );
NOR2_X1 U994 ( .A1(n1294), .A2(n1293), .ZN(n1130) );
NOR2_X1 U995 ( .A1(n1265), .A2(n1290), .ZN(n1126) );
XOR2_X1 U996 ( .A(n1322), .B(n1323), .Z(G12) );
NAND2_X1 U997 ( .A1(KEYINPUT30), .A2(G110), .ZN(n1323) );
NAND4_X1 U998 ( .A1(n1105), .A2(n1104), .A3(n1247), .A4(n1324), .ZN(n1322) );
XNOR2_X1 U999 ( .A(KEYINPUT12), .B(n1089), .ZN(n1324) );
INV_X1 U1000 ( .A(n1137), .ZN(n1089) );
NOR2_X1 U1001 ( .A1(n1139), .A2(n1138), .ZN(n1137) );
INV_X1 U1002 ( .A(n1291), .ZN(n1138) );
NAND2_X1 U1003 ( .A1(G214), .A2(n1325), .ZN(n1291) );
XOR2_X1 U1004 ( .A(n1326), .B(n1327), .Z(n1139) );
AND2_X1 U1005 ( .A1(n1325), .A2(G210), .ZN(n1327) );
NAND2_X1 U1006 ( .A1(n1328), .A2(n1329), .ZN(n1325) );
XNOR2_X1 U1007 ( .A(G237), .B(KEYINPUT52), .ZN(n1328) );
NAND2_X1 U1008 ( .A1(n1330), .A2(n1329), .ZN(n1326) );
XNOR2_X1 U1009 ( .A(n1331), .B(n1271), .ZN(n1330) );
XOR2_X1 U1010 ( .A(n1179), .B(n1332), .Z(n1271) );
NOR2_X1 U1011 ( .A1(KEYINPUT54), .A2(n1180), .ZN(n1332) );
XNOR2_X1 U1012 ( .A(n1333), .B(G122), .ZN(n1180) );
XOR2_X1 U1013 ( .A(n1334), .B(n1335), .Z(n1179) );
XNOR2_X1 U1014 ( .A(KEYINPUT33), .B(n1336), .ZN(n1335) );
XNOR2_X1 U1015 ( .A(n1222), .B(n1337), .ZN(n1334) );
NAND2_X1 U1016 ( .A1(n1338), .A2(n1339), .ZN(n1331) );
NAND2_X1 U1017 ( .A1(n1340), .A2(n1276), .ZN(n1339) );
XOR2_X1 U1018 ( .A(n1341), .B(KEYINPUT6), .Z(n1338) );
OR2_X1 U1019 ( .A1(n1276), .A2(n1340), .ZN(n1341) );
XNOR2_X1 U1020 ( .A(n1275), .B(n1342), .ZN(n1340) );
XNOR2_X1 U1021 ( .A(n1343), .B(KEYINPUT48), .ZN(n1342) );
NAND2_X1 U1022 ( .A1(KEYINPUT57), .A2(n1277), .ZN(n1343) );
XOR2_X1 U1023 ( .A(G125), .B(KEYINPUT40), .Z(n1275) );
NAND2_X1 U1024 ( .A1(G224), .A2(n1128), .ZN(n1276) );
AND2_X1 U1025 ( .A1(n1118), .A2(n1315), .ZN(n1247) );
NAND2_X1 U1026 ( .A1(n1108), .A2(n1344), .ZN(n1315) );
NAND4_X1 U1027 ( .A1(G953), .A2(G902), .A3(n1299), .A4(n1177), .ZN(n1344) );
INV_X1 U1028 ( .A(G898), .ZN(n1177) );
NAND3_X1 U1029 ( .A1(n1299), .A2(n1128), .A3(G952), .ZN(n1108) );
NAND2_X1 U1030 ( .A1(G234), .A2(G237), .ZN(n1299) );
AND2_X1 U1031 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U1032 ( .A1(G221), .A2(n1345), .ZN(n1120) );
XNOR2_X1 U1033 ( .A(n1346), .B(G469), .ZN(n1119) );
NAND2_X1 U1034 ( .A1(n1347), .A2(n1329), .ZN(n1346) );
XOR2_X1 U1035 ( .A(n1348), .B(n1349), .Z(n1347) );
XOR2_X1 U1036 ( .A(n1163), .B(n1233), .Z(n1349) );
XNOR2_X1 U1037 ( .A(n1350), .B(n1351), .ZN(n1233) );
XNOR2_X1 U1038 ( .A(G140), .B(n1333), .ZN(n1351) );
NAND2_X1 U1039 ( .A1(G227), .A2(n1128), .ZN(n1350) );
NAND2_X1 U1040 ( .A1(n1352), .A2(n1353), .ZN(n1163) );
NAND2_X1 U1041 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
XOR2_X1 U1042 ( .A(KEYINPUT42), .B(n1356), .Z(n1352) );
NOR2_X1 U1043 ( .A1(n1355), .A2(n1354), .ZN(n1356) );
XOR2_X1 U1044 ( .A(KEYINPUT17), .B(G128), .Z(n1354) );
XNOR2_X1 U1045 ( .A(n1357), .B(G146), .ZN(n1355) );
XNOR2_X1 U1046 ( .A(n1358), .B(n1359), .ZN(n1348) );
NOR2_X1 U1047 ( .A1(KEYINPUT51), .A2(n1227), .ZN(n1359) );
NAND2_X1 U1048 ( .A1(n1360), .A2(n1361), .ZN(n1227) );
NAND2_X1 U1049 ( .A1(n1337), .A2(G107), .ZN(n1361) );
NAND2_X1 U1050 ( .A1(n1362), .A2(n1336), .ZN(n1360) );
XNOR2_X1 U1051 ( .A(n1337), .B(KEYINPUT36), .ZN(n1362) );
XOR2_X1 U1052 ( .A(G104), .B(G101), .Z(n1337) );
NOR2_X1 U1053 ( .A1(KEYINPUT47), .A2(n1231), .ZN(n1358) );
NOR2_X1 U1054 ( .A1(n1294), .A2(n1141), .ZN(n1104) );
INV_X1 U1055 ( .A(n1293), .ZN(n1141) );
XNOR2_X1 U1056 ( .A(n1363), .B(n1192), .ZN(n1293) );
AND2_X1 U1057 ( .A1(G217), .A2(n1345), .ZN(n1192) );
NAND2_X1 U1058 ( .A1(G234), .A2(n1329), .ZN(n1345) );
NAND2_X1 U1059 ( .A1(n1190), .A2(n1329), .ZN(n1363) );
XNOR2_X1 U1060 ( .A(n1364), .B(n1365), .ZN(n1190) );
XOR2_X1 U1061 ( .A(n1366), .B(n1367), .Z(n1365) );
AND2_X1 U1062 ( .A1(n1368), .A2(G221), .ZN(n1366) );
XOR2_X1 U1063 ( .A(n1369), .B(n1370), .Z(n1364) );
XOR2_X1 U1064 ( .A(KEYINPUT19), .B(G137), .Z(n1370) );
NAND2_X1 U1065 ( .A1(n1371), .A2(n1372), .ZN(n1369) );
NAND2_X1 U1066 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
NAND2_X1 U1067 ( .A1(n1375), .A2(n1376), .ZN(n1374) );
NAND2_X1 U1068 ( .A1(G110), .A2(n1377), .ZN(n1376) );
INV_X1 U1069 ( .A(KEYINPUT1), .ZN(n1375) );
NAND2_X1 U1070 ( .A1(n1378), .A2(n1333), .ZN(n1371) );
INV_X1 U1071 ( .A(G110), .ZN(n1333) );
NAND2_X1 U1072 ( .A1(n1377), .A2(n1379), .ZN(n1378) );
OR2_X1 U1073 ( .A1(n1373), .A2(KEYINPUT1), .ZN(n1379) );
XOR2_X1 U1074 ( .A(G119), .B(n1380), .Z(n1373) );
XOR2_X1 U1075 ( .A(KEYINPUT29), .B(G128), .Z(n1380) );
INV_X1 U1076 ( .A(KEYINPUT23), .ZN(n1377) );
XNOR2_X1 U1077 ( .A(n1147), .B(G472), .ZN(n1294) );
NAND2_X1 U1078 ( .A1(n1381), .A2(n1329), .ZN(n1147) );
INV_X1 U1079 ( .A(G902), .ZN(n1329) );
XOR2_X1 U1080 ( .A(n1382), .B(n1222), .Z(n1381) );
XOR2_X1 U1081 ( .A(G113), .B(n1383), .Z(n1222) );
XNOR2_X1 U1082 ( .A(G119), .B(n1307), .ZN(n1383) );
XOR2_X1 U1083 ( .A(n1384), .B(n1218), .Z(n1382) );
NOR2_X1 U1084 ( .A1(n1220), .A2(n1385), .ZN(n1218) );
AND2_X1 U1085 ( .A1(n1386), .A2(G101), .ZN(n1385) );
NOR2_X1 U1086 ( .A1(n1386), .A2(G101), .ZN(n1220) );
AND3_X1 U1087 ( .A1(n1387), .A2(n1128), .A3(G210), .ZN(n1386) );
NAND2_X1 U1088 ( .A1(KEYINPUT39), .A2(n1214), .ZN(n1384) );
XNOR2_X1 U1089 ( .A(n1231), .B(n1277), .ZN(n1214) );
XNOR2_X1 U1090 ( .A(n1388), .B(n1389), .ZN(n1277) );
NOR2_X1 U1091 ( .A1(G146), .A2(KEYINPUT2), .ZN(n1389) );
XNOR2_X1 U1092 ( .A(G143), .B(G128), .ZN(n1388) );
XOR2_X1 U1093 ( .A(n1390), .B(n1391), .Z(n1231) );
XOR2_X1 U1094 ( .A(G137), .B(G131), .Z(n1391) );
NAND2_X1 U1095 ( .A1(KEYINPUT20), .A2(G134), .ZN(n1390) );
NOR2_X1 U1096 ( .A1(n1290), .A2(n1281), .ZN(n1105) );
INV_X1 U1097 ( .A(n1265), .ZN(n1281) );
XOR2_X1 U1098 ( .A(n1149), .B(n1392), .Z(n1265) );
NOR2_X1 U1099 ( .A1(G475), .A2(KEYINPUT9), .ZN(n1392) );
NOR2_X1 U1100 ( .A1(n1206), .A2(G902), .ZN(n1149) );
XNOR2_X1 U1101 ( .A(n1393), .B(n1394), .ZN(n1206) );
XOR2_X1 U1102 ( .A(n1395), .B(n1396), .Z(n1394) );
XOR2_X1 U1103 ( .A(G122), .B(G104), .Z(n1396) );
XNOR2_X1 U1104 ( .A(n1357), .B(G131), .ZN(n1395) );
XOR2_X1 U1105 ( .A(n1397), .B(n1398), .Z(n1393) );
XNOR2_X1 U1106 ( .A(n1399), .B(n1400), .ZN(n1398) );
NOR2_X1 U1107 ( .A1(KEYINPUT63), .A2(n1401), .ZN(n1400) );
NOR3_X1 U1108 ( .A1(n1402), .A2(G953), .A3(n1403), .ZN(n1401) );
INV_X1 U1109 ( .A(G214), .ZN(n1403) );
XNOR2_X1 U1110 ( .A(KEYINPUT5), .B(n1387), .ZN(n1402) );
INV_X1 U1111 ( .A(G237), .ZN(n1387) );
NAND2_X1 U1112 ( .A1(n1404), .A2(KEYINPUT24), .ZN(n1399) );
XNOR2_X1 U1113 ( .A(n1367), .B(KEYINPUT50), .ZN(n1404) );
XOR2_X1 U1114 ( .A(G146), .B(n1165), .Z(n1367) );
XNOR2_X1 U1115 ( .A(n1405), .B(G140), .ZN(n1165) );
INV_X1 U1116 ( .A(G125), .ZN(n1405) );
NAND2_X1 U1117 ( .A1(KEYINPUT11), .A2(n1317), .ZN(n1397) );
INV_X1 U1118 ( .A(G113), .ZN(n1317) );
XNOR2_X1 U1119 ( .A(n1151), .B(n1406), .ZN(n1290) );
NOR2_X1 U1120 ( .A1(G478), .A2(KEYINPUT49), .ZN(n1406) );
NOR2_X1 U1121 ( .A1(n1199), .A2(G902), .ZN(n1151) );
XNOR2_X1 U1122 ( .A(n1407), .B(n1408), .ZN(n1199) );
XOR2_X1 U1123 ( .A(n1409), .B(n1410), .Z(n1408) );
XNOR2_X1 U1124 ( .A(n1411), .B(n1307), .ZN(n1410) );
INV_X1 U1125 ( .A(G116), .ZN(n1307) );
NAND2_X1 U1126 ( .A1(KEYINPUT55), .A2(n1336), .ZN(n1411) );
INV_X1 U1127 ( .A(G107), .ZN(n1336) );
NAND2_X1 U1128 ( .A1(n1368), .A2(G217), .ZN(n1409) );
AND2_X1 U1129 ( .A1(G234), .A2(n1128), .ZN(n1368) );
INV_X1 U1130 ( .A(G953), .ZN(n1128) );
XOR2_X1 U1131 ( .A(n1412), .B(n1413), .Z(n1407) );
XNOR2_X1 U1132 ( .A(n1357), .B(G134), .ZN(n1413) );
INV_X1 U1133 ( .A(G143), .ZN(n1357) );
XNOR2_X1 U1134 ( .A(G122), .B(G128), .ZN(n1412) );
endmodule


