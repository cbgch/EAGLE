//Key = 0111111101111000000101011001010110011010011101100101100101111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319;

XOR2_X1 U721 ( .A(G107), .B(n997), .Z(G9) );
NOR2_X1 U722 ( .A1(n998), .A2(n999), .ZN(n997) );
XOR2_X1 U723 ( .A(n1000), .B(KEYINPUT60), .Z(n999) );
NOR2_X1 U724 ( .A1(n1001), .A2(n1002), .ZN(G75) );
NOR4_X1 U725 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1002) );
NOR3_X1 U726 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1005) );
NOR2_X1 U727 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NOR2_X1 U728 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR2_X1 U729 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR2_X1 U730 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR3_X1 U731 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1016) );
NOR2_X1 U732 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U733 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
AND2_X1 U734 ( .A1(n1025), .A2(KEYINPUT24), .ZN(n1024) );
NOR2_X1 U735 ( .A1(n1026), .A2(n1027), .ZN(n1023) );
XOR2_X1 U736 ( .A(n1028), .B(KEYINPUT6), .Z(n1026) );
NOR3_X1 U737 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1019) );
XOR2_X1 U738 ( .A(n1032), .B(KEYINPUT35), .Z(n1029) );
NOR2_X1 U739 ( .A1(KEYINPUT56), .A2(n1033), .ZN(n1018) );
NOR2_X1 U740 ( .A1(n1034), .A2(n1022), .ZN(n1014) );
NOR2_X1 U741 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U742 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U743 ( .A1(n1039), .A2(n1000), .ZN(n1037) );
NOR3_X1 U744 ( .A1(n1040), .A2(KEYINPUT24), .A3(n1041), .ZN(n1035) );
NOR3_X1 U745 ( .A1(n1022), .A2(n1038), .A3(n1042), .ZN(n1010) );
NAND4_X1 U746 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1003) );
NAND3_X1 U747 ( .A1(n1047), .A2(n1048), .A3(KEYINPUT56), .ZN(n1044) );
NAND3_X1 U748 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
INV_X1 U749 ( .A(n1013), .ZN(n1050) );
NAND3_X1 U750 ( .A1(n1052), .A2(n1053), .A3(n1051), .ZN(n1043) );
NOR3_X1 U751 ( .A1(n1009), .A2(n1038), .A3(n1017), .ZN(n1051) );
INV_X1 U752 ( .A(n1032), .ZN(n1038) );
NOR3_X1 U753 ( .A1(n1054), .A2(G953), .A3(G952), .ZN(n1001) );
INV_X1 U754 ( .A(n1045), .ZN(n1054) );
NAND4_X1 U755 ( .A1(n1055), .A2(n1028), .A3(n1056), .A4(n1057), .ZN(n1045) );
NOR3_X1 U756 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
XNOR2_X1 U757 ( .A(n1061), .B(KEYINPUT51), .ZN(n1059) );
NAND3_X1 U758 ( .A1(n1030), .A2(n1027), .A3(n1062), .ZN(n1058) );
NAND2_X1 U759 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR3_X1 U760 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1056) );
NOR2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
INV_X1 U762 ( .A(KEYINPUT27), .ZN(n1069) );
NOR2_X1 U763 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR3_X1 U764 ( .A1(n1072), .A2(n1063), .A3(n1064), .ZN(n1071) );
INV_X1 U765 ( .A(KEYINPUT4), .ZN(n1072) );
NOR2_X1 U766 ( .A1(KEYINPUT4), .A2(n1073), .ZN(n1070) );
NOR2_X1 U767 ( .A1(KEYINPUT27), .A2(n1074), .ZN(n1066) );
NOR2_X1 U768 ( .A1(n1063), .A2(n1075), .ZN(n1074) );
XOR2_X1 U769 ( .A(KEYINPUT4), .B(n1073), .Z(n1075) );
XOR2_X1 U770 ( .A(KEYINPUT34), .B(n1007), .Z(n1065) );
XOR2_X1 U771 ( .A(n1076), .B(n1077), .Z(n1055) );
NOR2_X1 U772 ( .A1(KEYINPUT50), .A2(n1078), .ZN(n1077) );
XOR2_X1 U773 ( .A(n1079), .B(n1080), .Z(G72) );
XOR2_X1 U774 ( .A(n1081), .B(n1082), .Z(n1080) );
NOR3_X1 U775 ( .A1(n1083), .A2(KEYINPUT22), .A3(n1084), .ZN(n1082) );
NOR2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
INV_X1 U777 ( .A(n1087), .ZN(n1083) );
NAND2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(n1081) );
NAND2_X1 U779 ( .A1(G953), .A2(n1086), .ZN(n1089) );
XOR2_X1 U780 ( .A(n1090), .B(n1091), .Z(n1088) );
XOR2_X1 U781 ( .A(n1092), .B(n1093), .Z(n1091) );
XOR2_X1 U782 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U783 ( .A1(n1096), .A2(KEYINPUT12), .ZN(n1095) );
XOR2_X1 U784 ( .A(n1097), .B(KEYINPUT43), .Z(n1096) );
INV_X1 U785 ( .A(G125), .ZN(n1097) );
XOR2_X1 U786 ( .A(n1098), .B(n1099), .Z(n1090) );
NOR2_X1 U787 ( .A1(KEYINPUT40), .A2(G131), .ZN(n1099) );
XOR2_X1 U788 ( .A(n1100), .B(KEYINPUT44), .Z(n1098) );
INV_X1 U789 ( .A(G140), .ZN(n1100) );
NAND2_X1 U790 ( .A1(n1046), .A2(n1006), .ZN(n1079) );
XOR2_X1 U791 ( .A(n1101), .B(n1102), .Z(G69) );
XOR2_X1 U792 ( .A(n1103), .B(n1104), .Z(n1102) );
NAND2_X1 U793 ( .A1(n1087), .A2(n1105), .ZN(n1104) );
NAND2_X1 U794 ( .A1(G898), .A2(G224), .ZN(n1105) );
XOR2_X1 U795 ( .A(n1046), .B(KEYINPUT49), .Z(n1087) );
NAND2_X1 U796 ( .A1(n1106), .A2(n1107), .ZN(n1103) );
NAND2_X1 U797 ( .A1(G953), .A2(n1108), .ZN(n1107) );
XOR2_X1 U798 ( .A(n1109), .B(n1110), .Z(n1106) );
XNOR2_X1 U799 ( .A(n1111), .B(KEYINPUT17), .ZN(n1110) );
NAND2_X1 U800 ( .A1(KEYINPUT52), .A2(n1112), .ZN(n1111) );
XOR2_X1 U801 ( .A(n1113), .B(n1114), .Z(n1109) );
AND2_X1 U802 ( .A1(n1004), .A2(n1046), .ZN(n1101) );
NOR2_X1 U803 ( .A1(n1115), .A2(n1116), .ZN(G66) );
XOR2_X1 U804 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND3_X1 U805 ( .A1(n1119), .A2(n1120), .A3(KEYINPUT42), .ZN(n1118) );
NOR2_X1 U806 ( .A1(n1115), .A2(n1121), .ZN(G63) );
XOR2_X1 U807 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U808 ( .A1(n1076), .A2(n1124), .ZN(n1122) );
INV_X1 U809 ( .A(G478), .ZN(n1076) );
NOR2_X1 U810 ( .A1(n1115), .A2(n1125), .ZN(G60) );
XNOR2_X1 U811 ( .A(n1126), .B(n1127), .ZN(n1125) );
AND2_X1 U812 ( .A1(G475), .A2(n1119), .ZN(n1127) );
XOR2_X1 U813 ( .A(G104), .B(n1128), .Z(G6) );
NOR2_X1 U814 ( .A1(n1115), .A2(n1129), .ZN(G57) );
XOR2_X1 U815 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U816 ( .A1(n1132), .A2(KEYINPUT57), .ZN(n1130) );
XOR2_X1 U817 ( .A(n1133), .B(n1134), .Z(n1132) );
AND2_X1 U818 ( .A1(G472), .A2(n1119), .ZN(n1134) );
NOR2_X1 U819 ( .A1(n1115), .A2(n1135), .ZN(G54) );
XOR2_X1 U820 ( .A(n1136), .B(n1137), .Z(n1135) );
NOR2_X1 U821 ( .A1(KEYINPUT53), .A2(n1138), .ZN(n1137) );
XOR2_X1 U822 ( .A(n1139), .B(n1140), .Z(n1138) );
XNOR2_X1 U823 ( .A(n1141), .B(n1142), .ZN(n1140) );
XOR2_X1 U824 ( .A(n1143), .B(n1144), .Z(n1139) );
XOR2_X1 U825 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND2_X1 U826 ( .A1(n1147), .A2(n1148), .ZN(n1145) );
NAND2_X1 U827 ( .A1(G140), .A2(n1149), .ZN(n1148) );
XOR2_X1 U828 ( .A(KEYINPUT10), .B(n1150), .Z(n1147) );
NOR2_X1 U829 ( .A1(G140), .A2(n1149), .ZN(n1150) );
NAND2_X1 U830 ( .A1(KEYINPUT41), .A2(n1151), .ZN(n1143) );
NAND2_X1 U831 ( .A1(n1119), .A2(G469), .ZN(n1136) );
INV_X1 U832 ( .A(n1124), .ZN(n1119) );
NOR2_X1 U833 ( .A1(n1115), .A2(n1152), .ZN(G51) );
XOR2_X1 U834 ( .A(n1153), .B(n1154), .Z(n1152) );
XNOR2_X1 U835 ( .A(KEYINPUT47), .B(n1155), .ZN(n1154) );
NOR3_X1 U836 ( .A1(n1124), .A2(KEYINPUT14), .A3(n1064), .ZN(n1155) );
NAND2_X1 U837 ( .A1(G902), .A2(n1156), .ZN(n1124) );
OR2_X1 U838 ( .A1(n1004), .A2(n1006), .ZN(n1156) );
NAND4_X1 U839 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1006) );
NOR4_X1 U840 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1160) );
INV_X1 U841 ( .A(n1165), .ZN(n1164) );
NAND2_X1 U842 ( .A1(n1052), .A2(n1166), .ZN(n1159) );
NAND2_X1 U843 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND2_X1 U844 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
XOR2_X1 U845 ( .A(KEYINPUT63), .B(n1025), .Z(n1170) );
INV_X1 U846 ( .A(n1171), .ZN(n1169) );
NAND2_X1 U847 ( .A1(n1172), .A2(n1000), .ZN(n1167) );
OR3_X1 U848 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1157) );
NAND4_X1 U849 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1004) );
NOR4_X1 U850 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1179) );
NOR2_X1 U851 ( .A1(n1184), .A2(n1128), .ZN(n1178) );
NOR2_X1 U852 ( .A1(n1173), .A2(n998), .ZN(n1128) );
NOR2_X1 U853 ( .A1(n1185), .A2(n998), .ZN(n1184) );
OR3_X1 U854 ( .A1(n1007), .A2(n1013), .A3(n1186), .ZN(n998) );
NAND2_X1 U855 ( .A1(n1187), .A2(n1047), .ZN(n1176) );
XOR2_X1 U856 ( .A(n1188), .B(KEYINPUT2), .Z(n1187) );
NOR2_X1 U857 ( .A1(n1046), .A2(G952), .ZN(n1115) );
XOR2_X1 U858 ( .A(G146), .B(n1189), .Z(G48) );
NOR4_X1 U859 ( .A1(KEYINPUT62), .A2(n1174), .A3(n1173), .A4(n1175), .ZN(n1189) );
NAND2_X1 U860 ( .A1(n1190), .A2(n1191), .ZN(G45) );
NAND2_X1 U861 ( .A1(n1192), .A2(n1158), .ZN(n1191) );
XOR2_X1 U862 ( .A(KEYINPUT11), .B(n1193), .Z(n1190) );
NOR2_X1 U863 ( .A1(n1192), .A2(n1158), .ZN(n1193) );
NAND2_X1 U864 ( .A1(n1172), .A2(n1194), .ZN(n1158) );
XNOR2_X1 U865 ( .A(KEYINPUT58), .B(G143), .ZN(n1192) );
XOR2_X1 U866 ( .A(G140), .B(n1195), .Z(G42) );
NOR3_X1 U867 ( .A1(n1022), .A2(n1040), .A3(n1171), .ZN(n1195) );
XOR2_X1 U868 ( .A(G137), .B(n1162), .Z(G39) );
NOR3_X1 U869 ( .A1(n1022), .A2(n1017), .A3(n1175), .ZN(n1162) );
XOR2_X1 U870 ( .A(G134), .B(n1196), .Z(G36) );
NOR3_X1 U871 ( .A1(n1197), .A2(n1185), .A3(n1198), .ZN(n1196) );
XOR2_X1 U872 ( .A(n1022), .B(KEYINPUT18), .Z(n1198) );
INV_X1 U873 ( .A(n1052), .ZN(n1022) );
XOR2_X1 U874 ( .A(n1199), .B(G131), .Z(G33) );
NAND2_X1 U875 ( .A1(KEYINPUT59), .A2(n1165), .ZN(n1199) );
NAND3_X1 U876 ( .A1(n1052), .A2(n1039), .A3(n1172), .ZN(n1165) );
INV_X1 U877 ( .A(n1197), .ZN(n1172) );
NAND3_X1 U878 ( .A1(n1025), .A2(n1200), .A3(n1053), .ZN(n1197) );
NOR2_X1 U879 ( .A1(n1031), .A2(n1201), .ZN(n1052) );
INV_X1 U880 ( .A(n1030), .ZN(n1201) );
XOR2_X1 U881 ( .A(G128), .B(n1163), .Z(G30) );
NOR3_X1 U882 ( .A1(n1174), .A2(n1185), .A3(n1175), .ZN(n1163) );
NAND4_X1 U883 ( .A1(n1025), .A2(n1061), .A3(n1007), .A4(n1200), .ZN(n1175) );
XOR2_X1 U884 ( .A(G101), .B(n1183), .Z(G3) );
NOR3_X1 U885 ( .A1(n1017), .A2(n1186), .A3(n1202), .ZN(n1183) );
XOR2_X1 U886 ( .A(G125), .B(n1161), .Z(G27) );
NOR2_X1 U887 ( .A1(n1171), .A2(n1033), .ZN(n1161) );
NAND4_X1 U888 ( .A1(n1049), .A2(n1039), .A3(n1061), .A4(n1200), .ZN(n1171) );
NAND2_X1 U889 ( .A1(n1009), .A2(n1203), .ZN(n1200) );
NAND4_X1 U890 ( .A1(G953), .A2(G902), .A3(n1204), .A4(n1086), .ZN(n1203) );
INV_X1 U891 ( .A(G900), .ZN(n1086) );
NAND2_X1 U892 ( .A1(n1205), .A2(n1206), .ZN(G24) );
OR2_X1 U893 ( .A1(n1177), .A2(G122), .ZN(n1206) );
XOR2_X1 U894 ( .A(n1207), .B(KEYINPUT28), .Z(n1205) );
NAND2_X1 U895 ( .A1(G122), .A2(n1177), .ZN(n1207) );
NAND4_X1 U896 ( .A1(n1049), .A2(n1194), .A3(n1208), .A4(n1032), .ZN(n1177) );
NOR2_X1 U897 ( .A1(n1209), .A2(n1013), .ZN(n1208) );
XNOR2_X1 U898 ( .A(n1210), .B(KEYINPUT25), .ZN(n1013) );
NOR3_X1 U899 ( .A1(n1174), .A2(n1211), .A3(n1212), .ZN(n1194) );
XNOR2_X1 U900 ( .A(G119), .B(n1213), .ZN(G21) );
NOR2_X1 U901 ( .A1(n1182), .A2(KEYINPUT39), .ZN(n1213) );
NOR4_X1 U902 ( .A1(n1033), .A2(n1042), .A3(n1049), .A4(n1209), .ZN(n1182) );
XNOR2_X1 U903 ( .A(G116), .B(n1214), .ZN(G18) );
NAND2_X1 U904 ( .A1(KEYINPUT31), .A2(n1181), .ZN(n1214) );
NOR4_X1 U905 ( .A1(n1202), .A2(n1033), .A3(n1185), .A4(n1209), .ZN(n1181) );
INV_X1 U906 ( .A(n1215), .ZN(n1209) );
INV_X1 U907 ( .A(n1000), .ZN(n1185) );
NAND2_X1 U908 ( .A1(n1216), .A2(n1217), .ZN(n1000) );
OR3_X1 U909 ( .A1(n1211), .A2(n1218), .A3(KEYINPUT54), .ZN(n1217) );
NAND2_X1 U910 ( .A1(KEYINPUT54), .A2(n1041), .ZN(n1216) );
NAND2_X1 U911 ( .A1(n1047), .A2(n1032), .ZN(n1033) );
XNOR2_X1 U912 ( .A(G113), .B(n1219), .ZN(G15) );
NAND2_X1 U913 ( .A1(n1220), .A2(n1047), .ZN(n1219) );
XOR2_X1 U914 ( .A(n1188), .B(KEYINPUT1), .Z(n1220) );
NAND4_X1 U915 ( .A1(n1039), .A2(n1053), .A3(n1032), .A4(n1215), .ZN(n1188) );
NAND2_X1 U916 ( .A1(n1221), .A2(n1222), .ZN(n1032) );
OR2_X1 U917 ( .A1(n1040), .A2(KEYINPUT6), .ZN(n1222) );
NAND3_X1 U918 ( .A1(n1028), .A2(n1027), .A3(KEYINPUT6), .ZN(n1221) );
INV_X1 U919 ( .A(n1202), .ZN(n1053) );
NAND2_X1 U920 ( .A1(n1210), .A2(n1007), .ZN(n1202) );
XOR2_X1 U921 ( .A(n1061), .B(KEYINPUT61), .Z(n1210) );
INV_X1 U922 ( .A(n1173), .ZN(n1039) );
NAND2_X1 U923 ( .A1(n1218), .A2(n1211), .ZN(n1173) );
XOR2_X1 U924 ( .A(n1149), .B(n1223), .Z(G12) );
NOR2_X1 U925 ( .A1(n1180), .A2(KEYINPUT37), .ZN(n1223) );
NOR3_X1 U926 ( .A1(n1007), .A2(n1186), .A3(n1042), .ZN(n1180) );
NAND2_X1 U927 ( .A1(n1041), .A2(n1061), .ZN(n1042) );
XNOR2_X1 U928 ( .A(n1224), .B(n1120), .ZN(n1061) );
AND2_X1 U929 ( .A1(G217), .A2(n1225), .ZN(n1120) );
NAND2_X1 U930 ( .A1(n1226), .A2(n1117), .ZN(n1224) );
NAND3_X1 U931 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1117) );
NAND2_X1 U932 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND2_X1 U933 ( .A1(KEYINPUT33), .A2(n1232), .ZN(n1228) );
NAND2_X1 U934 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
XNOR2_X1 U935 ( .A(KEYINPUT8), .B(n1230), .ZN(n1233) );
NAND2_X1 U936 ( .A1(n1235), .A2(n1236), .ZN(n1227) );
INV_X1 U937 ( .A(KEYINPUT33), .ZN(n1236) );
NAND2_X1 U938 ( .A1(n1237), .A2(n1238), .ZN(n1235) );
OR3_X1 U939 ( .A1(n1231), .A2(n1230), .A3(KEYINPUT8), .ZN(n1238) );
INV_X1 U940 ( .A(n1234), .ZN(n1231) );
XOR2_X1 U941 ( .A(n1239), .B(n1240), .Z(n1234) );
XOR2_X1 U942 ( .A(n1241), .B(n1242), .Z(n1240) );
NOR2_X1 U943 ( .A1(G119), .A2(KEYINPUT20), .ZN(n1241) );
XOR2_X1 U944 ( .A(n1243), .B(n1244), .Z(n1239) );
NOR2_X1 U945 ( .A1(KEYINPUT0), .A2(n1245), .ZN(n1244) );
XOR2_X1 U946 ( .A(n1246), .B(G110), .Z(n1243) );
NAND2_X1 U947 ( .A1(KEYINPUT8), .A2(n1230), .ZN(n1237) );
AND2_X1 U948 ( .A1(n1247), .A2(n1248), .ZN(n1230) );
NAND2_X1 U949 ( .A1(n1249), .A2(G137), .ZN(n1248) );
XOR2_X1 U950 ( .A(KEYINPUT45), .B(n1250), .Z(n1247) );
NOR2_X1 U951 ( .A1(n1249), .A2(G137), .ZN(n1250) );
AND3_X1 U952 ( .A1(n1251), .A2(n1046), .A3(G234), .ZN(n1249) );
XOR2_X1 U953 ( .A(KEYINPUT26), .B(G221), .Z(n1251) );
INV_X1 U954 ( .A(n1017), .ZN(n1041) );
NAND2_X1 U955 ( .A1(n1211), .A2(n1212), .ZN(n1017) );
INV_X1 U956 ( .A(n1218), .ZN(n1212) );
XNOR2_X1 U957 ( .A(n1060), .B(KEYINPUT9), .ZN(n1218) );
XNOR2_X1 U958 ( .A(n1252), .B(G475), .ZN(n1060) );
NAND2_X1 U959 ( .A1(n1126), .A2(n1226), .ZN(n1252) );
XNOR2_X1 U960 ( .A(n1253), .B(n1254), .ZN(n1126) );
XOR2_X1 U961 ( .A(G131), .B(n1255), .Z(n1254) );
XOR2_X1 U962 ( .A(G146), .B(G143), .Z(n1255) );
XOR2_X1 U963 ( .A(n1256), .B(n1242), .Z(n1253) );
XOR2_X1 U964 ( .A(G125), .B(G140), .Z(n1242) );
XOR2_X1 U965 ( .A(n1257), .B(n1258), .Z(n1256) );
AND2_X1 U966 ( .A1(G214), .A2(n1259), .ZN(n1258) );
NAND2_X1 U967 ( .A1(n1260), .A2(n1261), .ZN(n1257) );
NAND2_X1 U968 ( .A1(G104), .A2(n1262), .ZN(n1261) );
XOR2_X1 U969 ( .A(KEYINPUT46), .B(n1263), .Z(n1260) );
NOR2_X1 U970 ( .A1(G104), .A2(n1262), .ZN(n1263) );
XOR2_X1 U971 ( .A(G122), .B(G113), .Z(n1262) );
XOR2_X1 U972 ( .A(n1078), .B(G478), .Z(n1211) );
OR2_X1 U973 ( .A1(n1123), .A2(G902), .ZN(n1078) );
XNOR2_X1 U974 ( .A(n1264), .B(n1265), .ZN(n1123) );
XOR2_X1 U975 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U976 ( .A(n1268), .B(G107), .Z(n1267) );
NAND2_X1 U977 ( .A1(KEYINPUT5), .A2(n1269), .ZN(n1268) );
NAND2_X1 U978 ( .A1(n1270), .A2(KEYINPUT19), .ZN(n1266) );
XOR2_X1 U979 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U980 ( .A(n1273), .B(n1274), .Z(n1264) );
NAND3_X1 U981 ( .A1(G234), .A2(n1046), .A3(G217), .ZN(n1273) );
NAND3_X1 U982 ( .A1(n1025), .A2(n1215), .A3(n1047), .ZN(n1186) );
INV_X1 U983 ( .A(n1174), .ZN(n1047) );
NAND2_X1 U984 ( .A1(n1031), .A2(n1030), .ZN(n1174) );
NAND2_X1 U985 ( .A1(G214), .A2(n1275), .ZN(n1030) );
XOR2_X1 U986 ( .A(n1063), .B(n1073), .Z(n1031) );
INV_X1 U987 ( .A(n1064), .ZN(n1073) );
NAND2_X1 U988 ( .A1(G210), .A2(n1275), .ZN(n1064) );
NAND2_X1 U989 ( .A1(n1276), .A2(n1226), .ZN(n1275) );
INV_X1 U990 ( .A(G237), .ZN(n1276) );
AND2_X1 U991 ( .A1(n1153), .A2(n1226), .ZN(n1063) );
XOR2_X1 U992 ( .A(n1277), .B(n1278), .Z(n1153) );
XOR2_X1 U993 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U994 ( .A(KEYINPUT7), .B(G125), .Z(n1280) );
AND2_X1 U995 ( .A1(n1046), .A2(G224), .ZN(n1279) );
XOR2_X1 U996 ( .A(n1281), .B(n1282), .Z(n1277) );
INV_X1 U997 ( .A(n1113), .ZN(n1282) );
XOR2_X1 U998 ( .A(n1283), .B(n1284), .Z(n1113) );
NOR2_X1 U999 ( .A1(KEYINPUT30), .A2(n1285), .ZN(n1284) );
NAND2_X1 U1000 ( .A1(n1286), .A2(n1287), .ZN(n1283) );
NAND2_X1 U1001 ( .A1(G110), .A2(n1271), .ZN(n1287) );
XOR2_X1 U1002 ( .A(KEYINPUT55), .B(n1288), .Z(n1286) );
NOR2_X1 U1003 ( .A1(G110), .A2(n1271), .ZN(n1288) );
INV_X1 U1004 ( .A(G122), .ZN(n1271) );
XOR2_X1 U1005 ( .A(n1289), .B(n1112), .Z(n1281) );
XNOR2_X1 U1006 ( .A(n1290), .B(n1291), .ZN(n1112) );
NAND2_X1 U1007 ( .A1(KEYINPUT23), .A2(n1292), .ZN(n1290) );
NAND2_X1 U1008 ( .A1(n1293), .A2(n1294), .ZN(n1215) );
NAND4_X1 U1009 ( .A1(G953), .A2(G902), .A3(n1204), .A4(n1108), .ZN(n1294) );
INV_X1 U1010 ( .A(G898), .ZN(n1108) );
XOR2_X1 U1011 ( .A(n1009), .B(KEYINPUT16), .Z(n1293) );
NAND3_X1 U1012 ( .A1(n1204), .A2(n1046), .A3(G952), .ZN(n1009) );
INV_X1 U1013 ( .A(G953), .ZN(n1046) );
NAND2_X1 U1014 ( .A1(G237), .A2(G234), .ZN(n1204) );
INV_X1 U1015 ( .A(n1040), .ZN(n1025) );
NAND2_X1 U1016 ( .A1(n1295), .A2(n1027), .ZN(n1040) );
NAND2_X1 U1017 ( .A1(G221), .A2(n1225), .ZN(n1027) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1226), .ZN(n1225) );
INV_X1 U1019 ( .A(n1028), .ZN(n1295) );
XOR2_X1 U1020 ( .A(n1296), .B(G469), .Z(n1028) );
NAND2_X1 U1021 ( .A1(n1297), .A2(n1226), .ZN(n1296) );
XOR2_X1 U1022 ( .A(n1298), .B(n1299), .Z(n1297) );
XOR2_X1 U1023 ( .A(n1151), .B(n1142), .Z(n1299) );
XOR2_X1 U1024 ( .A(n1291), .B(n1292), .Z(n1142) );
XOR2_X1 U1025 ( .A(G107), .B(G104), .Z(n1292) );
XOR2_X1 U1026 ( .A(G101), .B(KEYINPUT48), .Z(n1291) );
XNOR2_X1 U1027 ( .A(n1300), .B(n1301), .ZN(n1298) );
NAND2_X1 U1028 ( .A1(KEYINPUT21), .A2(n1141), .ZN(n1301) );
XOR2_X1 U1029 ( .A(n1094), .B(KEYINPUT29), .Z(n1141) );
NAND2_X1 U1030 ( .A1(n1302), .A2(n1303), .ZN(n1094) );
NAND2_X1 U1031 ( .A1(n1304), .A2(n1245), .ZN(n1303) );
XOR2_X1 U1032 ( .A(KEYINPUT13), .B(n1305), .Z(n1304) );
NAND2_X1 U1033 ( .A1(KEYINPUT3), .A2(n1306), .ZN(n1300) );
XOR2_X1 U1034 ( .A(n1146), .B(n1307), .Z(n1306) );
XOR2_X1 U1035 ( .A(G140), .B(G110), .Z(n1307) );
NOR2_X1 U1036 ( .A1(n1085), .A2(G953), .ZN(n1146) );
INV_X1 U1037 ( .A(G227), .ZN(n1085) );
INV_X1 U1038 ( .A(n1049), .ZN(n1007) );
XOR2_X1 U1039 ( .A(n1308), .B(G472), .Z(n1049) );
NAND2_X1 U1040 ( .A1(n1309), .A2(n1226), .ZN(n1308) );
INV_X1 U1041 ( .A(G902), .ZN(n1226) );
XOR2_X1 U1042 ( .A(n1133), .B(n1310), .Z(n1309) );
XOR2_X1 U1043 ( .A(KEYINPUT38), .B(n1311), .Z(n1310) );
INV_X1 U1044 ( .A(n1131), .ZN(n1311) );
XOR2_X1 U1045 ( .A(n1312), .B(G101), .Z(n1131) );
NAND2_X1 U1046 ( .A1(n1259), .A2(G210), .ZN(n1312) );
NOR2_X1 U1047 ( .A1(G953), .A2(G237), .ZN(n1259) );
XNOR2_X1 U1048 ( .A(n1313), .B(n1151), .ZN(n1133) );
XNOR2_X1 U1049 ( .A(G131), .B(n1314), .ZN(n1151) );
INV_X1 U1050 ( .A(n1092), .ZN(n1314) );
XOR2_X1 U1051 ( .A(n1269), .B(G137), .Z(n1092) );
INV_X1 U1052 ( .A(G134), .ZN(n1269) );
XOR2_X1 U1053 ( .A(n1289), .B(n1315), .Z(n1313) );
NOR2_X1 U1054 ( .A1(KEYINPUT15), .A2(n1272), .ZN(n1315) );
INV_X1 U1055 ( .A(n1285), .ZN(n1272) );
XNOR2_X1 U1056 ( .A(G116), .B(KEYINPUT36), .ZN(n1285) );
XOR2_X1 U1057 ( .A(n1316), .B(n1114), .Z(n1289) );
XOR2_X1 U1058 ( .A(G119), .B(G113), .Z(n1114) );
NAND2_X1 U1059 ( .A1(n1302), .A2(n1317), .ZN(n1316) );
NAND2_X1 U1060 ( .A1(n1318), .A2(n1245), .ZN(n1317) );
XOR2_X1 U1061 ( .A(KEYINPUT32), .B(n1274), .Z(n1318) );
XOR2_X1 U1062 ( .A(G128), .B(G143), .Z(n1274) );
OR2_X1 U1063 ( .A1(n1245), .A2(n1305), .ZN(n1302) );
XNOR2_X1 U1064 ( .A(n1246), .B(n1319), .ZN(n1305) );
XOR2_X1 U1065 ( .A(KEYINPUT32), .B(G143), .Z(n1319) );
INV_X1 U1066 ( .A(G128), .ZN(n1246) );
INV_X1 U1067 ( .A(G146), .ZN(n1245) );
INV_X1 U1068 ( .A(G110), .ZN(n1149) );
endmodule


