//Key = 1011111110111011111110101011111100101010010010001010101010011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388;

NAND3_X1 U768 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(G9) );
NAND2_X1 U769 ( .A1(KEYINPUT58), .A2(n1062), .ZN(n1061) );
NAND3_X1 U770 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1060) );
NAND2_X1 U771 ( .A1(G107), .A2(n1066), .ZN(n1059) );
NAND2_X1 U772 ( .A1(n1067), .A2(n1064), .ZN(n1066) );
INV_X1 U773 ( .A(KEYINPUT58), .ZN(n1064) );
XNOR2_X1 U774 ( .A(KEYINPUT37), .B(n1062), .ZN(n1067) );
NOR2_X1 U775 ( .A1(n1068), .A2(n1069), .ZN(G75) );
NOR4_X1 U776 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
XOR2_X1 U777 ( .A(n1074), .B(KEYINPUT10), .Z(n1073) );
NAND4_X1 U778 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
XNOR2_X1 U779 ( .A(n1079), .B(KEYINPUT4), .ZN(n1075) );
NOR2_X1 U780 ( .A1(n1080), .A2(n1081), .ZN(n1072) );
NOR3_X1 U781 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1080) );
NOR2_X1 U782 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U783 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR2_X1 U784 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR2_X1 U785 ( .A1(n1091), .A2(n1092), .ZN(n1087) );
XOR2_X1 U786 ( .A(KEYINPUT5), .B(n1093), .Z(n1092) );
NOR3_X1 U787 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1083) );
XNOR2_X1 U788 ( .A(n1079), .B(KEYINPUT42), .ZN(n1094) );
NOR2_X1 U789 ( .A1(n1097), .A2(n1098), .ZN(n1082) );
NAND4_X1 U790 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1070) );
NAND4_X1 U791 ( .A1(n1103), .A2(n1104), .A3(n1079), .A4(n1105), .ZN(n1100) );
NOR3_X1 U792 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
NOR3_X1 U793 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1108) );
NOR2_X1 U794 ( .A1(n1077), .A2(n1112), .ZN(n1107) );
INV_X1 U795 ( .A(n1097), .ZN(n1079) );
NAND3_X1 U796 ( .A1(n1113), .A2(n1090), .A3(n1114), .ZN(n1099) );
INV_X1 U797 ( .A(KEYINPUT12), .ZN(n1090) );
OR2_X1 U798 ( .A1(n1081), .A2(n1086), .ZN(n1113) );
INV_X1 U799 ( .A(n1104), .ZN(n1086) );
NAND4_X1 U800 ( .A1(n1076), .A2(n1077), .A3(n1103), .A4(n1112), .ZN(n1081) );
INV_X1 U801 ( .A(n1106), .ZN(n1076) );
NOR3_X1 U802 ( .A1(n1115), .A2(G953), .A3(G952), .ZN(n1068) );
INV_X1 U803 ( .A(n1101), .ZN(n1115) );
NAND4_X1 U804 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1101) );
NOR4_X1 U805 ( .A1(n1109), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1119) );
XNOR2_X1 U806 ( .A(n1123), .B(KEYINPUT3), .ZN(n1122) );
XNOR2_X1 U807 ( .A(n1124), .B(n1125), .ZN(n1121) );
NOR2_X1 U808 ( .A1(KEYINPUT61), .A2(n1126), .ZN(n1125) );
XNOR2_X1 U809 ( .A(G478), .B(KEYINPUT59), .ZN(n1126) );
NOR2_X1 U810 ( .A1(n1127), .A2(n1128), .ZN(n1118) );
XNOR2_X1 U811 ( .A(n1129), .B(n1130), .ZN(n1116) );
XOR2_X1 U812 ( .A(KEYINPUT53), .B(G472), .Z(n1130) );
XOR2_X1 U813 ( .A(n1131), .B(n1132), .Z(G72) );
XOR2_X1 U814 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U815 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U816 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U817 ( .A(KEYINPUT25), .B(n1139), .Z(n1138) );
NOR3_X1 U818 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
NOR2_X1 U819 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NOR2_X1 U820 ( .A1(n1145), .A2(n1146), .ZN(n1143) );
INV_X1 U821 ( .A(KEYINPUT7), .ZN(n1146) );
XOR2_X1 U822 ( .A(n1147), .B(KEYINPUT38), .Z(n1145) );
AND3_X1 U823 ( .A1(n1144), .A2(n1147), .A3(KEYINPUT7), .ZN(n1141) );
XOR2_X1 U824 ( .A(n1148), .B(n1149), .Z(n1144) );
NOR2_X1 U825 ( .A1(KEYINPUT13), .A2(n1150), .ZN(n1149) );
NOR2_X1 U826 ( .A1(KEYINPUT7), .A2(n1147), .ZN(n1140) );
NOR2_X1 U827 ( .A1(n1151), .A2(n1152), .ZN(n1133) );
XNOR2_X1 U828 ( .A(KEYINPUT52), .B(n1102), .ZN(n1152) );
AND2_X1 U829 ( .A1(G227), .A2(G900), .ZN(n1151) );
NOR3_X1 U830 ( .A1(n1153), .A2(KEYINPUT62), .A3(G953), .ZN(n1131) );
NAND3_X1 U831 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(G69) );
OR2_X1 U832 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND3_X1 U833 ( .A1(n1158), .A2(n1157), .A3(G953), .ZN(n1155) );
NAND2_X1 U834 ( .A1(n1159), .A2(G224), .ZN(n1158) );
XNOR2_X1 U835 ( .A(G898), .B(KEYINPUT28), .ZN(n1159) );
NAND2_X1 U836 ( .A1(n1160), .A2(n1102), .ZN(n1154) );
NAND2_X1 U837 ( .A1(n1157), .A2(n1161), .ZN(n1160) );
OR2_X1 U838 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND3_X1 U839 ( .A1(n1164), .A2(n1165), .A3(n1162), .ZN(n1157) );
XOR2_X1 U840 ( .A(n1166), .B(n1167), .Z(n1162) );
NAND2_X1 U841 ( .A1(KEYINPUT11), .A2(n1168), .ZN(n1166) );
NAND2_X1 U842 ( .A1(G953), .A2(n1169), .ZN(n1165) );
XOR2_X1 U843 ( .A(KEYINPUT22), .B(n1170), .Z(n1164) );
NOR2_X1 U844 ( .A1(n1163), .A2(G953), .ZN(n1170) );
NOR2_X1 U845 ( .A1(n1171), .A2(n1172), .ZN(G66) );
XOR2_X1 U846 ( .A(n1173), .B(n1174), .Z(n1172) );
NAND3_X1 U847 ( .A1(n1175), .A2(n1176), .A3(G902), .ZN(n1173) );
XNOR2_X1 U848 ( .A(KEYINPUT6), .B(n1071), .ZN(n1176) );
NOR2_X1 U849 ( .A1(n1171), .A2(n1177), .ZN(G63) );
NOR3_X1 U850 ( .A1(n1124), .A2(n1178), .A3(n1179), .ZN(n1177) );
NOR3_X1 U851 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1179) );
NOR2_X1 U852 ( .A1(n1183), .A2(n1184), .ZN(n1178) );
AND2_X1 U853 ( .A1(n1071), .A2(G478), .ZN(n1183) );
NOR2_X1 U854 ( .A1(n1171), .A2(n1185), .ZN(G60) );
XOR2_X1 U855 ( .A(n1186), .B(n1187), .Z(n1185) );
NAND2_X1 U856 ( .A1(n1188), .A2(G475), .ZN(n1186) );
XNOR2_X1 U857 ( .A(n1189), .B(n1190), .ZN(G6) );
NOR2_X1 U858 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XNOR2_X1 U859 ( .A(n1114), .B(KEYINPUT57), .ZN(n1191) );
NOR2_X1 U860 ( .A1(n1171), .A2(n1193), .ZN(G57) );
NOR2_X1 U861 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
XOR2_X1 U862 ( .A(n1196), .B(KEYINPUT50), .Z(n1195) );
NAND2_X1 U863 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NOR2_X1 U864 ( .A1(n1197), .A2(n1198), .ZN(n1194) );
AND2_X1 U865 ( .A1(n1199), .A2(n1200), .ZN(n1197) );
NAND4_X1 U866 ( .A1(n1188), .A2(G472), .A3(n1201), .A4(n1202), .ZN(n1200) );
NAND2_X1 U867 ( .A1(n1203), .A2(n1204), .ZN(n1199) );
NAND2_X1 U868 ( .A1(n1201), .A2(n1202), .ZN(n1204) );
NAND2_X1 U869 ( .A1(n1205), .A2(n1206), .ZN(n1202) );
XNOR2_X1 U870 ( .A(n1207), .B(n1208), .ZN(n1205) );
INV_X1 U871 ( .A(n1209), .ZN(n1207) );
XNOR2_X1 U872 ( .A(n1210), .B(KEYINPUT17), .ZN(n1201) );
NAND2_X1 U873 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
INV_X1 U874 ( .A(n1206), .ZN(n1212) );
XNOR2_X1 U875 ( .A(n1209), .B(n1208), .ZN(n1211) );
NAND2_X1 U876 ( .A1(n1188), .A2(G472), .ZN(n1203) );
NOR2_X1 U877 ( .A1(n1171), .A2(n1213), .ZN(G54) );
XOR2_X1 U878 ( .A(n1214), .B(n1215), .Z(n1213) );
XOR2_X1 U879 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U880 ( .A(n1147), .B(n1218), .Z(n1217) );
XNOR2_X1 U881 ( .A(KEYINPUT31), .B(KEYINPUT23), .ZN(n1216) );
XOR2_X1 U882 ( .A(n1219), .B(n1220), .Z(n1214) );
XNOR2_X1 U883 ( .A(n1221), .B(n1208), .ZN(n1220) );
NAND2_X1 U884 ( .A1(n1188), .A2(G469), .ZN(n1221) );
XOR2_X1 U885 ( .A(n1222), .B(n1223), .Z(n1219) );
NOR2_X1 U886 ( .A1(n1171), .A2(n1224), .ZN(G51) );
XOR2_X1 U887 ( .A(n1225), .B(n1226), .Z(n1224) );
XOR2_X1 U888 ( .A(n1227), .B(n1228), .Z(n1226) );
XNOR2_X1 U889 ( .A(G125), .B(n1229), .ZN(n1228) );
NAND2_X1 U890 ( .A1(n1188), .A2(n1230), .ZN(n1227) );
INV_X1 U891 ( .A(n1182), .ZN(n1188) );
NAND2_X1 U892 ( .A1(G902), .A2(n1071), .ZN(n1182) );
NAND2_X1 U893 ( .A1(n1153), .A2(n1163), .ZN(n1071) );
AND4_X1 U894 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1163) );
NOR4_X1 U895 ( .A1(n1235), .A2(n1236), .A3(n1237), .A4(n1063), .ZN(n1234) );
INV_X1 U896 ( .A(n1062), .ZN(n1063) );
NAND4_X1 U897 ( .A1(n1114), .A2(n1110), .A3(n1078), .A4(n1238), .ZN(n1062) );
NAND2_X1 U898 ( .A1(n1114), .A2(n1239), .ZN(n1233) );
NAND2_X1 U899 ( .A1(n1240), .A2(n1192), .ZN(n1239) );
NAND3_X1 U900 ( .A1(n1078), .A2(n1238), .A3(n1111), .ZN(n1192) );
AND2_X1 U901 ( .A1(n1241), .A2(n1104), .ZN(n1078) );
XOR2_X1 U902 ( .A(n1242), .B(KEYINPUT43), .Z(n1240) );
AND4_X1 U903 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1153) );
NOR4_X1 U904 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1246) );
NOR2_X1 U905 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
INV_X1 U906 ( .A(KEYINPUT36), .ZN(n1252) );
NOR3_X1 U907 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1249) );
INV_X1 U908 ( .A(n1110), .ZN(n1255) );
NOR2_X1 U909 ( .A1(n1256), .A2(n1257), .ZN(n1254) );
NOR3_X1 U910 ( .A1(n1097), .A2(KEYINPUT36), .A3(n1258), .ZN(n1257) );
NOR2_X1 U911 ( .A1(n1259), .A2(n1260), .ZN(n1256) );
XNOR2_X1 U912 ( .A(KEYINPUT63), .B(n1089), .ZN(n1260) );
XOR2_X1 U913 ( .A(KEYINPUT24), .B(n1261), .Z(n1259) );
INV_X1 U914 ( .A(n1262), .ZN(n1247) );
AND2_X1 U915 ( .A1(n1263), .A2(n1264), .ZN(n1245) );
XNOR2_X1 U916 ( .A(n1209), .B(n1265), .ZN(n1225) );
NOR2_X1 U917 ( .A1(KEYINPUT21), .A2(n1266), .ZN(n1265) );
NOR2_X1 U918 ( .A1(n1102), .A2(G952), .ZN(n1171) );
XNOR2_X1 U919 ( .A(n1248), .B(n1267), .ZN(G48) );
XNOR2_X1 U920 ( .A(G146), .B(KEYINPUT9), .ZN(n1267) );
AND4_X1 U921 ( .A1(n1261), .A2(n1268), .A3(n1111), .A4(n1114), .ZN(n1248) );
XNOR2_X1 U922 ( .A(G143), .B(n1262), .ZN(G45) );
NAND4_X1 U923 ( .A1(n1127), .A2(n1269), .A3(n1114), .A4(n1270), .ZN(n1262) );
NOR2_X1 U924 ( .A1(n1253), .A2(n1098), .ZN(n1270) );
INV_X1 U925 ( .A(n1258), .ZN(n1098) );
XNOR2_X1 U926 ( .A(G140), .B(n1271), .ZN(G42) );
NAND2_X1 U927 ( .A1(KEYINPUT30), .A2(n1272), .ZN(n1271) );
INV_X1 U928 ( .A(n1243), .ZN(n1272) );
NAND4_X1 U929 ( .A1(n1273), .A2(n1111), .A3(n1123), .A4(n1274), .ZN(n1243) );
XNOR2_X1 U930 ( .A(G137), .B(n1244), .ZN(G39) );
NAND3_X1 U931 ( .A1(n1261), .A2(n1273), .A3(n1077), .ZN(n1244) );
XOR2_X1 U932 ( .A(n1251), .B(n1275), .Z(G36) );
NAND2_X1 U933 ( .A1(KEYINPUT18), .A2(G134), .ZN(n1275) );
NAND3_X1 U934 ( .A1(n1273), .A2(n1110), .A3(n1258), .ZN(n1251) );
XOR2_X1 U935 ( .A(n1264), .B(n1276), .Z(G33) );
NAND2_X1 U936 ( .A1(KEYINPUT14), .A2(G131), .ZN(n1276) );
NAND3_X1 U937 ( .A1(n1273), .A2(n1111), .A3(n1258), .ZN(n1264) );
NOR2_X1 U938 ( .A1(n1253), .A2(n1097), .ZN(n1273) );
NAND2_X1 U939 ( .A1(n1093), .A2(n1091), .ZN(n1097) );
XNOR2_X1 U940 ( .A(n1277), .B(n1278), .ZN(G30) );
NAND2_X1 U941 ( .A1(KEYINPUT34), .A2(n1279), .ZN(n1277) );
NAND4_X1 U942 ( .A1(n1261), .A2(n1268), .A3(n1114), .A4(n1110), .ZN(n1279) );
INV_X1 U943 ( .A(n1253), .ZN(n1268) );
NAND2_X1 U944 ( .A1(n1241), .A2(n1280), .ZN(n1253) );
XOR2_X1 U945 ( .A(G101), .B(n1281), .Z(G3) );
NOR2_X1 U946 ( .A1(n1089), .A2(n1242), .ZN(n1281) );
NAND4_X1 U947 ( .A1(n1077), .A2(n1258), .A3(n1241), .A4(n1238), .ZN(n1242) );
NOR2_X1 U948 ( .A1(n1103), .A2(n1109), .ZN(n1241) );
XNOR2_X1 U949 ( .A(G125), .B(n1263), .ZN(G27) );
NAND4_X1 U950 ( .A1(n1111), .A2(n1282), .A3(n1103), .A4(n1280), .ZN(n1263) );
NAND2_X1 U951 ( .A1(n1283), .A2(n1106), .ZN(n1280) );
NAND2_X1 U952 ( .A1(n1135), .A2(n1284), .ZN(n1283) );
NOR2_X1 U953 ( .A1(n1102), .A2(G900), .ZN(n1135) );
XNOR2_X1 U954 ( .A(G122), .B(n1231), .ZN(G24) );
NAND4_X1 U955 ( .A1(n1285), .A2(n1104), .A3(n1127), .A4(n1269), .ZN(n1231) );
NOR2_X1 U956 ( .A1(n1123), .A2(n1095), .ZN(n1104) );
XOR2_X1 U957 ( .A(G119), .B(n1237), .Z(G21) );
AND3_X1 U958 ( .A1(n1077), .A2(n1261), .A3(n1285), .ZN(n1237) );
NOR2_X1 U959 ( .A1(n1274), .A2(n1096), .ZN(n1261) );
XNOR2_X1 U960 ( .A(n1286), .B(n1236), .ZN(G18) );
AND3_X1 U961 ( .A1(n1258), .A2(n1110), .A3(n1285), .ZN(n1236) );
NOR2_X1 U962 ( .A1(n1127), .A2(n1287), .ZN(n1110) );
NAND2_X1 U963 ( .A1(n1288), .A2(n1289), .ZN(G15) );
NAND2_X1 U964 ( .A1(n1235), .A2(n1290), .ZN(n1289) );
XOR2_X1 U965 ( .A(KEYINPUT29), .B(n1291), .Z(n1288) );
NOR2_X1 U966 ( .A1(n1235), .A2(n1290), .ZN(n1291) );
INV_X1 U967 ( .A(G113), .ZN(n1290) );
AND3_X1 U968 ( .A1(n1258), .A2(n1111), .A3(n1285), .ZN(n1235) );
AND4_X1 U969 ( .A1(n1103), .A2(n1114), .A3(n1238), .A4(n1112), .ZN(n1285) );
INV_X1 U970 ( .A(n1292), .ZN(n1103) );
AND2_X1 U971 ( .A1(n1287), .A2(n1127), .ZN(n1111) );
INV_X1 U972 ( .A(n1269), .ZN(n1287) );
NOR2_X1 U973 ( .A1(n1274), .A2(n1123), .ZN(n1258) );
XNOR2_X1 U974 ( .A(G110), .B(n1232), .ZN(G12) );
NAND4_X1 U975 ( .A1(n1077), .A2(n1282), .A3(n1292), .A4(n1238), .ZN(n1232) );
NAND2_X1 U976 ( .A1(n1293), .A2(n1106), .ZN(n1238) );
NAND3_X1 U977 ( .A1(n1294), .A2(n1102), .A3(G952), .ZN(n1106) );
XOR2_X1 U978 ( .A(n1295), .B(KEYINPUT55), .Z(n1293) );
NAND3_X1 U979 ( .A1(n1284), .A2(n1169), .A3(G953), .ZN(n1295) );
INV_X1 U980 ( .A(G898), .ZN(n1169) );
AND2_X1 U981 ( .A1(G902), .A2(n1294), .ZN(n1284) );
NAND2_X1 U982 ( .A1(G237), .A2(G234), .ZN(n1294) );
XNOR2_X1 U983 ( .A(n1117), .B(KEYINPUT40), .ZN(n1292) );
XOR2_X1 U984 ( .A(n1296), .B(G469), .Z(n1117) );
NAND2_X1 U985 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XOR2_X1 U986 ( .A(n1299), .B(n1300), .Z(n1297) );
XNOR2_X1 U987 ( .A(n1301), .B(n1302), .ZN(n1300) );
NAND2_X1 U988 ( .A1(KEYINPUT2), .A2(n1303), .ZN(n1302) );
NAND2_X1 U989 ( .A1(n1304), .A2(KEYINPUT56), .ZN(n1301) );
XNOR2_X1 U990 ( .A(n1223), .B(KEYINPUT15), .ZN(n1304) );
XOR2_X1 U991 ( .A(n1305), .B(n1218), .Z(n1299) );
AND2_X1 U992 ( .A1(G227), .A2(n1102), .ZN(n1218) );
NAND2_X1 U993 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U994 ( .A1(n1222), .A2(n1147), .ZN(n1307) );
XOR2_X1 U995 ( .A(KEYINPUT48), .B(n1308), .Z(n1306) );
NOR2_X1 U996 ( .A1(n1222), .A2(n1147), .ZN(n1308) );
NAND3_X1 U997 ( .A1(n1309), .A2(n1310), .A3(n1311), .ZN(n1147) );
OR2_X1 U998 ( .A1(n1312), .A2(KEYINPUT16), .ZN(n1311) );
NAND3_X1 U999 ( .A1(KEYINPUT16), .A2(n1312), .A3(G128), .ZN(n1310) );
NAND2_X1 U1000 ( .A1(n1313), .A2(n1278), .ZN(n1309) );
NAND2_X1 U1001 ( .A1(n1314), .A2(KEYINPUT16), .ZN(n1313) );
XNOR2_X1 U1002 ( .A(n1312), .B(KEYINPUT26), .ZN(n1314) );
XOR2_X1 U1003 ( .A(n1315), .B(n1316), .Z(n1222) );
XNOR2_X1 U1004 ( .A(n1189), .B(G101), .ZN(n1316) );
XNOR2_X1 U1005 ( .A(n1317), .B(n1065), .ZN(n1315) );
XNOR2_X1 U1006 ( .A(KEYINPUT51), .B(KEYINPUT32), .ZN(n1317) );
NOR4_X1 U1007 ( .A1(n1089), .A2(n1096), .A3(n1095), .A4(n1109), .ZN(n1282) );
INV_X1 U1008 ( .A(n1112), .ZN(n1109) );
NAND2_X1 U1009 ( .A1(G221), .A2(n1318), .ZN(n1112) );
INV_X1 U1010 ( .A(n1274), .ZN(n1095) );
XOR2_X1 U1011 ( .A(G472), .B(n1319), .Z(n1274) );
NOR2_X1 U1012 ( .A1(n1129), .A2(KEYINPUT46), .ZN(n1319) );
AND2_X1 U1013 ( .A1(n1320), .A2(n1298), .ZN(n1129) );
XOR2_X1 U1014 ( .A(n1321), .B(n1322), .Z(n1320) );
XNOR2_X1 U1015 ( .A(n1208), .B(n1198), .ZN(n1322) );
XOR2_X1 U1016 ( .A(n1323), .B(G101), .Z(n1198) );
NAND2_X1 U1017 ( .A1(n1324), .A2(G210), .ZN(n1323) );
INV_X1 U1018 ( .A(n1303), .ZN(n1208) );
XOR2_X1 U1019 ( .A(n1148), .B(n1150), .Z(n1303) );
XNOR2_X1 U1020 ( .A(G134), .B(G137), .ZN(n1150) );
XOR2_X1 U1021 ( .A(n1325), .B(n1326), .Z(n1321) );
NOR2_X1 U1022 ( .A1(KEYINPUT47), .A2(n1327), .ZN(n1326) );
XNOR2_X1 U1023 ( .A(n1206), .B(KEYINPUT41), .ZN(n1327) );
XNOR2_X1 U1024 ( .A(n1328), .B(n1329), .ZN(n1206) );
NOR2_X1 U1025 ( .A1(G119), .A2(KEYINPUT49), .ZN(n1329) );
XNOR2_X1 U1026 ( .A(G116), .B(G113), .ZN(n1328) );
NOR2_X1 U1027 ( .A1(n1209), .A2(n1330), .ZN(n1325) );
XOR2_X1 U1028 ( .A(KEYINPUT8), .B(KEYINPUT27), .Z(n1330) );
INV_X1 U1029 ( .A(n1123), .ZN(n1096) );
XNOR2_X1 U1030 ( .A(n1331), .B(n1175), .ZN(n1123) );
AND2_X1 U1031 ( .A1(G217), .A2(n1318), .ZN(n1175) );
NAND2_X1 U1032 ( .A1(G234), .A2(n1298), .ZN(n1318) );
NAND2_X1 U1033 ( .A1(n1174), .A2(n1298), .ZN(n1331) );
XNOR2_X1 U1034 ( .A(n1332), .B(n1333), .ZN(n1174) );
XOR2_X1 U1035 ( .A(n1334), .B(n1335), .Z(n1333) );
XNOR2_X1 U1036 ( .A(n1278), .B(G125), .ZN(n1335) );
XOR2_X1 U1037 ( .A(G146), .B(G137), .Z(n1334) );
XOR2_X1 U1038 ( .A(n1336), .B(n1223), .Z(n1332) );
XNOR2_X1 U1039 ( .A(G140), .B(n1337), .ZN(n1223) );
XOR2_X1 U1040 ( .A(n1338), .B(G119), .Z(n1336) );
NAND2_X1 U1041 ( .A1(G221), .A2(n1339), .ZN(n1338) );
INV_X1 U1042 ( .A(n1114), .ZN(n1089) );
NOR2_X1 U1043 ( .A1(n1093), .A2(n1120), .ZN(n1114) );
INV_X1 U1044 ( .A(n1091), .ZN(n1120) );
NAND2_X1 U1045 ( .A1(G214), .A2(n1340), .ZN(n1091) );
XOR2_X1 U1046 ( .A(n1128), .B(KEYINPUT44), .Z(n1093) );
XNOR2_X1 U1047 ( .A(n1341), .B(n1230), .ZN(n1128) );
AND2_X1 U1048 ( .A1(G210), .A2(n1340), .ZN(n1230) );
NAND2_X1 U1049 ( .A1(n1342), .A2(n1298), .ZN(n1340) );
INV_X1 U1050 ( .A(G237), .ZN(n1342) );
NAND2_X1 U1051 ( .A1(n1343), .A2(n1298), .ZN(n1341) );
XNOR2_X1 U1052 ( .A(n1344), .B(n1266), .ZN(n1343) );
XNOR2_X1 U1053 ( .A(n1167), .B(n1168), .ZN(n1266) );
AND2_X1 U1054 ( .A1(n1345), .A2(n1346), .ZN(n1168) );
NAND2_X1 U1055 ( .A1(G122), .A2(n1337), .ZN(n1346) );
XOR2_X1 U1056 ( .A(KEYINPUT20), .B(n1347), .Z(n1345) );
NOR2_X1 U1057 ( .A1(G122), .A2(n1337), .ZN(n1347) );
INV_X1 U1058 ( .A(G110), .ZN(n1337) );
XNOR2_X1 U1059 ( .A(n1348), .B(n1349), .ZN(n1167) );
NOR2_X1 U1060 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
XOR2_X1 U1061 ( .A(KEYINPUT39), .B(n1352), .Z(n1351) );
NOR2_X1 U1062 ( .A1(G113), .A2(n1353), .ZN(n1352) );
AND2_X1 U1063 ( .A1(n1353), .A2(G113), .ZN(n1350) );
XOR2_X1 U1064 ( .A(G116), .B(G119), .Z(n1353) );
XOR2_X1 U1065 ( .A(n1354), .B(G101), .Z(n1348) );
NAND2_X1 U1066 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
NAND2_X1 U1067 ( .A1(G104), .A2(n1065), .ZN(n1356) );
INV_X1 U1068 ( .A(G107), .ZN(n1065) );
XOR2_X1 U1069 ( .A(n1357), .B(KEYINPUT1), .Z(n1355) );
NAND2_X1 U1070 ( .A1(G107), .A2(n1189), .ZN(n1357) );
INV_X1 U1071 ( .A(G104), .ZN(n1189) );
NAND2_X1 U1072 ( .A1(n1358), .A2(n1359), .ZN(n1344) );
NAND2_X1 U1073 ( .A1(n1229), .A2(n1360), .ZN(n1359) );
XOR2_X1 U1074 ( .A(KEYINPUT19), .B(n1361), .Z(n1358) );
NOR2_X1 U1075 ( .A1(n1360), .A2(n1362), .ZN(n1361) );
XOR2_X1 U1076 ( .A(KEYINPUT45), .B(n1229), .Z(n1362) );
AND2_X1 U1077 ( .A1(G224), .A2(n1102), .ZN(n1229) );
XOR2_X1 U1078 ( .A(G125), .B(n1363), .Z(n1360) );
NOR2_X1 U1079 ( .A1(KEYINPUT33), .A2(n1209), .ZN(n1363) );
XOR2_X1 U1080 ( .A(G128), .B(n1312), .Z(n1209) );
XOR2_X1 U1081 ( .A(G143), .B(G146), .Z(n1312) );
NOR2_X1 U1082 ( .A1(n1269), .A2(n1127), .ZN(n1077) );
XNOR2_X1 U1083 ( .A(n1364), .B(G475), .ZN(n1127) );
NAND2_X1 U1084 ( .A1(n1187), .A2(n1298), .ZN(n1364) );
INV_X1 U1085 ( .A(G902), .ZN(n1298) );
XNOR2_X1 U1086 ( .A(n1365), .B(n1366), .ZN(n1187) );
XOR2_X1 U1087 ( .A(n1367), .B(n1368), .Z(n1366) );
XNOR2_X1 U1088 ( .A(G104), .B(G143), .ZN(n1368) );
NAND2_X1 U1089 ( .A1(KEYINPUT0), .A2(n1369), .ZN(n1367) );
XOR2_X1 U1090 ( .A(G146), .B(n1137), .Z(n1369) );
XOR2_X1 U1091 ( .A(G140), .B(G125), .Z(n1137) );
XNOR2_X1 U1092 ( .A(n1370), .B(n1371), .ZN(n1365) );
INV_X1 U1093 ( .A(n1148), .ZN(n1371) );
XOR2_X1 U1094 ( .A(G131), .B(KEYINPUT54), .Z(n1148) );
XOR2_X1 U1095 ( .A(n1372), .B(n1373), .Z(n1370) );
AND2_X1 U1096 ( .A1(G214), .A2(n1324), .ZN(n1373) );
NOR2_X1 U1097 ( .A1(G953), .A2(G237), .ZN(n1324) );
NAND2_X1 U1098 ( .A1(n1374), .A2(n1375), .ZN(n1372) );
NAND2_X1 U1099 ( .A1(G113), .A2(n1376), .ZN(n1375) );
XOR2_X1 U1100 ( .A(KEYINPUT60), .B(n1377), .Z(n1374) );
NOR2_X1 U1101 ( .A1(G113), .A2(n1376), .ZN(n1377) );
INV_X1 U1102 ( .A(G122), .ZN(n1376) );
NAND2_X1 U1103 ( .A1(n1378), .A2(n1379), .ZN(n1269) );
NAND2_X1 U1104 ( .A1(G478), .A2(n1380), .ZN(n1379) );
INV_X1 U1105 ( .A(n1124), .ZN(n1380) );
XOR2_X1 U1106 ( .A(n1381), .B(KEYINPUT35), .Z(n1378) );
NAND2_X1 U1107 ( .A1(n1124), .A2(n1181), .ZN(n1381) );
INV_X1 U1108 ( .A(G478), .ZN(n1181) );
NOR2_X1 U1109 ( .A1(n1184), .A2(G902), .ZN(n1124) );
INV_X1 U1110 ( .A(n1180), .ZN(n1184) );
XNOR2_X1 U1111 ( .A(n1382), .B(n1383), .ZN(n1180) );
XOR2_X1 U1112 ( .A(n1384), .B(n1385), .Z(n1383) );
XNOR2_X1 U1113 ( .A(n1278), .B(G122), .ZN(n1385) );
INV_X1 U1114 ( .A(G128), .ZN(n1278) );
XNOR2_X1 U1115 ( .A(n1386), .B(G134), .ZN(n1384) );
INV_X1 U1116 ( .A(G143), .ZN(n1386) );
XOR2_X1 U1117 ( .A(n1387), .B(n1388), .Z(n1382) );
XNOR2_X1 U1118 ( .A(n1286), .B(G107), .ZN(n1388) );
INV_X1 U1119 ( .A(G116), .ZN(n1286) );
NAND2_X1 U1120 ( .A1(G217), .A2(n1339), .ZN(n1387) );
AND2_X1 U1121 ( .A1(G234), .A2(n1102), .ZN(n1339) );
INV_X1 U1122 ( .A(G953), .ZN(n1102) );
endmodule


