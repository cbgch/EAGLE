//Key = 1001000011111110000110001111101100001001100001101000101010011111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
n1456, n1457, n1458, n1459, n1460, n1461, n1462;

XOR2_X1 U807 ( .A(n1116), .B(n1117), .Z(G9) );
XNOR2_X1 U808 ( .A(G107), .B(KEYINPUT33), .ZN(n1117) );
NAND2_X1 U809 ( .A1(KEYINPUT40), .A2(n1118), .ZN(n1116) );
NOR2_X1 U810 ( .A1(n1119), .A2(n1120), .ZN(G75) );
NOR3_X1 U811 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1120) );
NOR2_X1 U812 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
NOR3_X1 U813 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1124) );
NOR2_X1 U814 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
INV_X1 U815 ( .A(n1131), .ZN(n1130) );
NOR2_X1 U816 ( .A1(n1132), .A2(n1133), .ZN(n1129) );
NOR2_X1 U817 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NOR2_X1 U818 ( .A1(n1136), .A2(n1137), .ZN(n1134) );
NOR2_X1 U819 ( .A1(n1138), .A2(n1139), .ZN(n1136) );
NOR2_X1 U820 ( .A1(n1140), .A2(n1141), .ZN(n1132) );
XNOR2_X1 U821 ( .A(KEYINPUT52), .B(n1142), .ZN(n1141) );
NOR4_X1 U822 ( .A1(n1143), .A2(n1142), .A3(n1135), .A4(n1144), .ZN(n1127) );
INV_X1 U823 ( .A(n1145), .ZN(n1142) );
NOR2_X1 U824 ( .A1(n1146), .A2(n1147), .ZN(n1143) );
XOR2_X1 U825 ( .A(n1148), .B(KEYINPUT59), .Z(n1126) );
NAND4_X1 U826 ( .A1(n1149), .A2(n1131), .A3(n1150), .A4(n1145), .ZN(n1148) );
NAND3_X1 U827 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1121) );
NAND4_X1 U828 ( .A1(n1131), .A2(n1154), .A3(n1145), .A4(n1155), .ZN(n1153) );
NAND2_X1 U829 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U830 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NOR2_X1 U831 ( .A1(n1144), .A2(n1160), .ZN(n1131) );
NOR3_X1 U832 ( .A1(n1161), .A2(G953), .A3(G952), .ZN(n1119) );
INV_X1 U833 ( .A(n1151), .ZN(n1161) );
NAND4_X1 U834 ( .A1(n1162), .A2(n1154), .A3(n1163), .A4(n1164), .ZN(n1151) );
NOR4_X1 U835 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
XOR2_X1 U836 ( .A(n1169), .B(G472), .Z(n1167) );
NAND2_X1 U837 ( .A1(KEYINPUT26), .A2(n1170), .ZN(n1169) );
AND2_X1 U838 ( .A1(n1171), .A2(n1172), .ZN(n1166) );
XOR2_X1 U839 ( .A(n1173), .B(n1174), .Z(G72) );
XOR2_X1 U840 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U841 ( .A1(G953), .A2(n1177), .ZN(n1176) );
NAND2_X1 U842 ( .A1(G900), .A2(G227), .ZN(n1177) );
NAND3_X1 U843 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1175) );
XOR2_X1 U844 ( .A(n1181), .B(KEYINPUT58), .Z(n1180) );
NAND3_X1 U845 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1181) );
XNOR2_X1 U846 ( .A(n1185), .B(n1186), .ZN(n1184) );
NAND3_X1 U847 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1179) );
NAND2_X1 U848 ( .A1(n1186), .A2(n1185), .ZN(n1189) );
NAND2_X1 U849 ( .A1(n1182), .A2(n1183), .ZN(n1187) );
NAND2_X1 U850 ( .A1(n1190), .A2(n1191), .ZN(n1183) );
XNOR2_X1 U851 ( .A(n1192), .B(KEYINPUT42), .ZN(n1190) );
OR2_X1 U852 ( .A1(n1191), .A2(n1193), .ZN(n1182) );
XOR2_X1 U853 ( .A(n1194), .B(n1195), .Z(n1191) );
NOR2_X1 U854 ( .A1(KEYINPUT6), .A2(G131), .ZN(n1195) );
NAND2_X1 U855 ( .A1(G953), .A2(n1196), .ZN(n1178) );
XNOR2_X1 U856 ( .A(KEYINPUT9), .B(n1197), .ZN(n1196) );
NOR2_X1 U857 ( .A1(n1198), .A2(G953), .ZN(n1173) );
NOR2_X1 U858 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U859 ( .A(n1201), .B(n1202), .Z(G69) );
NOR2_X1 U860 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NOR2_X1 U861 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XNOR2_X1 U862 ( .A(KEYINPUT15), .B(n1207), .ZN(n1206) );
NOR2_X1 U863 ( .A1(n1207), .A2(n1208), .ZN(n1203) );
XNOR2_X1 U864 ( .A(KEYINPUT7), .B(n1205), .ZN(n1208) );
NAND2_X1 U865 ( .A1(n1152), .A2(n1209), .ZN(n1205) );
NAND3_X1 U866 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1207) );
XOR2_X1 U867 ( .A(n1213), .B(KEYINPUT18), .Z(n1212) );
OR2_X1 U868 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND2_X1 U869 ( .A1(n1214), .A2(n1215), .ZN(n1211) );
XNOR2_X1 U870 ( .A(n1216), .B(n1217), .ZN(n1214) );
NAND2_X1 U871 ( .A1(KEYINPUT31), .A2(n1218), .ZN(n1216) );
NAND2_X1 U872 ( .A1(G953), .A2(n1219), .ZN(n1210) );
NAND2_X1 U873 ( .A1(G953), .A2(n1220), .ZN(n1201) );
NAND2_X1 U874 ( .A1(G898), .A2(G224), .ZN(n1220) );
NOR3_X1 U875 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(G66) );
AND3_X1 U876 ( .A1(KEYINPUT29), .A2(G953), .A3(G952), .ZN(n1223) );
NOR2_X1 U877 ( .A1(KEYINPUT29), .A2(n1224), .ZN(n1222) );
INV_X1 U878 ( .A(n1225), .ZN(n1224) );
XOR2_X1 U879 ( .A(n1226), .B(n1227), .Z(n1221) );
NOR2_X1 U880 ( .A1(n1171), .A2(n1228), .ZN(n1227) );
NOR2_X1 U881 ( .A1(n1225), .A2(n1229), .ZN(G63) );
XNOR2_X1 U882 ( .A(n1230), .B(n1231), .ZN(n1229) );
AND2_X1 U883 ( .A1(G478), .A2(n1232), .ZN(n1231) );
NOR2_X1 U884 ( .A1(n1225), .A2(n1233), .ZN(G60) );
XOR2_X1 U885 ( .A(n1234), .B(n1235), .Z(n1233) );
AND2_X1 U886 ( .A1(G475), .A2(n1232), .ZN(n1234) );
XOR2_X1 U887 ( .A(G104), .B(n1236), .Z(G6) );
NOR2_X1 U888 ( .A1(KEYINPUT21), .A2(n1237), .ZN(n1236) );
NOR2_X1 U889 ( .A1(n1238), .A2(n1239), .ZN(G57) );
XOR2_X1 U890 ( .A(n1240), .B(n1241), .Z(n1239) );
XNOR2_X1 U891 ( .A(n1242), .B(n1243), .ZN(n1241) );
XOR2_X1 U892 ( .A(n1244), .B(n1245), .Z(n1240) );
AND2_X1 U893 ( .A1(G472), .A2(n1232), .ZN(n1245) );
XNOR2_X1 U894 ( .A(n1225), .B(KEYINPUT28), .ZN(n1238) );
NOR2_X1 U895 ( .A1(n1225), .A2(n1246), .ZN(G54) );
NOR2_X1 U896 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
XOR2_X1 U897 ( .A(n1249), .B(n1250), .Z(n1248) );
NOR2_X1 U898 ( .A1(KEYINPUT34), .A2(n1251), .ZN(n1250) );
AND2_X1 U899 ( .A1(G469), .A2(n1232), .ZN(n1249) );
AND2_X1 U900 ( .A1(n1251), .A2(KEYINPUT34), .ZN(n1247) );
XNOR2_X1 U901 ( .A(n1252), .B(n1253), .ZN(n1251) );
XOR2_X1 U902 ( .A(n1254), .B(n1255), .Z(n1252) );
NAND3_X1 U903 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1254) );
NAND2_X1 U904 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
INV_X1 U905 ( .A(KEYINPUT63), .ZN(n1260) );
XNOR2_X1 U906 ( .A(n1261), .B(n1262), .ZN(n1259) );
NOR2_X1 U907 ( .A1(n1193), .A2(n1263), .ZN(n1262) );
NAND2_X1 U908 ( .A1(KEYINPUT63), .A2(n1264), .ZN(n1256) );
NOR2_X1 U909 ( .A1(n1225), .A2(n1265), .ZN(G51) );
XOR2_X1 U910 ( .A(n1266), .B(n1267), .Z(n1265) );
NAND2_X1 U911 ( .A1(n1232), .A2(G210), .ZN(n1267) );
INV_X1 U912 ( .A(n1228), .ZN(n1232) );
NAND2_X1 U913 ( .A1(G902), .A2(n1123), .ZN(n1228) );
OR3_X1 U914 ( .A1(n1268), .A2(n1209), .A3(n1200), .ZN(n1123) );
NAND4_X1 U915 ( .A1(n1269), .A2(n1270), .A3(n1271), .A4(n1272), .ZN(n1200) );
AND4_X1 U916 ( .A1(n1273), .A2(n1274), .A3(n1275), .A4(n1276), .ZN(n1272) );
OR2_X1 U917 ( .A1(n1277), .A2(n1125), .ZN(n1271) );
NAND4_X1 U918 ( .A1(n1278), .A2(n1279), .A3(n1280), .A4(n1281), .ZN(n1209) );
AND4_X1 U919 ( .A1(n1282), .A2(n1283), .A3(n1284), .A4(n1237), .ZN(n1281) );
NAND3_X1 U920 ( .A1(n1285), .A2(n1145), .A3(n1147), .ZN(n1237) );
INV_X1 U921 ( .A(n1286), .ZN(n1282) );
NOR2_X1 U922 ( .A1(n1287), .A2(n1118), .ZN(n1280) );
AND3_X1 U923 ( .A1(n1146), .A2(n1145), .A3(n1285), .ZN(n1118) );
NOR4_X1 U924 ( .A1(n1288), .A2(n1289), .A3(n1160), .A4(n1290), .ZN(n1287) );
INV_X1 U925 ( .A(n1291), .ZN(n1160) );
NOR2_X1 U926 ( .A1(KEYINPUT46), .A2(n1292), .ZN(n1289) );
NOR3_X1 U927 ( .A1(n1293), .A2(n1294), .A3(n1156), .ZN(n1292) );
INV_X1 U928 ( .A(n1295), .ZN(n1156) );
INV_X1 U929 ( .A(n1296), .ZN(n1294) );
NOR2_X1 U930 ( .A1(n1285), .A2(n1297), .ZN(n1288) );
INV_X1 U931 ( .A(KEYINPUT46), .ZN(n1297) );
XNOR2_X1 U932 ( .A(n1199), .B(KEYINPUT25), .ZN(n1268) );
NAND2_X1 U933 ( .A1(n1298), .A2(n1299), .ZN(n1199) );
NAND4_X1 U934 ( .A1(n1300), .A2(n1147), .A3(n1301), .A4(n1302), .ZN(n1299) );
NOR2_X1 U935 ( .A1(n1290), .A2(n1303), .ZN(n1301) );
OR2_X1 U936 ( .A1(n1304), .A2(n1302), .ZN(n1298) );
INV_X1 U937 ( .A(KEYINPUT24), .ZN(n1302) );
NAND2_X1 U938 ( .A1(n1305), .A2(KEYINPUT20), .ZN(n1266) );
XNOR2_X1 U939 ( .A(n1306), .B(n1307), .ZN(n1305) );
NOR3_X1 U940 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1307) );
NOR2_X1 U941 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
INV_X1 U942 ( .A(KEYINPUT10), .ZN(n1312) );
NOR2_X1 U943 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
NOR2_X1 U944 ( .A1(KEYINPUT13), .A2(n1315), .ZN(n1314) );
NOR3_X1 U945 ( .A1(n1186), .A2(n1244), .A3(n1316), .ZN(n1313) );
INV_X1 U946 ( .A(KEYINPUT13), .ZN(n1316) );
NOR2_X1 U947 ( .A1(KEYINPUT10), .A2(n1317), .ZN(n1309) );
NOR2_X1 U948 ( .A1(n1318), .A2(n1244), .ZN(n1317) );
XNOR2_X1 U949 ( .A(KEYINPUT13), .B(n1186), .ZN(n1318) );
NOR2_X1 U950 ( .A1(n1152), .A2(G952), .ZN(n1225) );
XNOR2_X1 U951 ( .A(G146), .B(n1269), .ZN(G48) );
NAND4_X1 U952 ( .A1(n1319), .A2(n1295), .A3(n1320), .A4(n1321), .ZN(n1269) );
XNOR2_X1 U953 ( .A(G143), .B(n1270), .ZN(G45) );
NAND4_X1 U954 ( .A1(n1322), .A2(n1323), .A3(n1295), .A4(n1324), .ZN(n1270) );
XNOR2_X1 U955 ( .A(G140), .B(n1276), .ZN(G42) );
NAND3_X1 U956 ( .A1(n1325), .A2(n1319), .A3(n1300), .ZN(n1276) );
NAND2_X1 U957 ( .A1(n1326), .A2(n1327), .ZN(G39) );
NAND2_X1 U958 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
XOR2_X1 U959 ( .A(KEYINPUT56), .B(n1330), .Z(n1326) );
NOR2_X1 U960 ( .A1(n1328), .A2(n1329), .ZN(n1330) );
INV_X1 U961 ( .A(n1275), .ZN(n1328) );
NAND3_X1 U962 ( .A1(n1300), .A2(n1303), .A3(n1331), .ZN(n1275) );
NOR2_X1 U963 ( .A1(n1125), .A2(n1140), .ZN(n1300) );
INV_X1 U964 ( .A(n1320), .ZN(n1140) );
INV_X1 U965 ( .A(n1163), .ZN(n1125) );
XNOR2_X1 U966 ( .A(G134), .B(n1332), .ZN(G36) );
NAND2_X1 U967 ( .A1(n1333), .A2(n1163), .ZN(n1332) );
XOR2_X1 U968 ( .A(n1277), .B(KEYINPUT3), .Z(n1333) );
NAND2_X1 U969 ( .A1(n1323), .A2(n1146), .ZN(n1277) );
XNOR2_X1 U970 ( .A(G131), .B(n1304), .ZN(G33) );
NAND3_X1 U971 ( .A1(n1147), .A2(n1163), .A3(n1323), .ZN(n1304) );
AND3_X1 U972 ( .A1(n1320), .A2(n1303), .A3(n1137), .ZN(n1323) );
XOR2_X1 U973 ( .A(n1296), .B(KEYINPUT49), .Z(n1320) );
NOR2_X1 U974 ( .A1(n1334), .A2(n1158), .ZN(n1163) );
NAND2_X1 U975 ( .A1(n1335), .A2(n1336), .ZN(G30) );
NAND2_X1 U976 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
NAND2_X1 U977 ( .A1(n1339), .A2(G128), .ZN(n1335) );
NAND2_X1 U978 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
NAND2_X1 U979 ( .A1(KEYINPUT44), .A2(n1342), .ZN(n1341) );
INV_X1 U980 ( .A(n1274), .ZN(n1342) );
OR2_X1 U981 ( .A1(n1337), .A2(KEYINPUT44), .ZN(n1340) );
NOR2_X1 U982 ( .A1(KEYINPUT57), .A2(n1274), .ZN(n1337) );
NAND4_X1 U983 ( .A1(n1303), .A2(n1343), .A3(n1321), .A4(n1344), .ZN(n1274) );
AND3_X1 U984 ( .A1(n1146), .A2(n1296), .A3(n1295), .ZN(n1344) );
XNOR2_X1 U985 ( .A(n1345), .B(n1346), .ZN(G3) );
NOR2_X1 U986 ( .A1(n1290), .A2(n1347), .ZN(n1346) );
XNOR2_X1 U987 ( .A(G125), .B(n1273), .ZN(G27) );
NAND4_X1 U988 ( .A1(n1319), .A2(n1154), .A3(n1325), .A4(n1295), .ZN(n1273) );
INV_X1 U989 ( .A(n1139), .ZN(n1325) );
AND3_X1 U990 ( .A1(n1303), .A2(n1343), .A3(n1147), .ZN(n1319) );
NAND2_X1 U991 ( .A1(n1144), .A2(n1348), .ZN(n1303) );
NAND4_X1 U992 ( .A1(G953), .A2(G902), .A3(n1349), .A4(n1197), .ZN(n1348) );
INV_X1 U993 ( .A(G900), .ZN(n1197) );
XNOR2_X1 U994 ( .A(G122), .B(n1278), .ZN(G24) );
NAND4_X1 U995 ( .A1(n1350), .A2(n1145), .A3(n1322), .A4(n1324), .ZN(n1278) );
NOR2_X1 U996 ( .A1(n1343), .A2(n1139), .ZN(n1145) );
XNOR2_X1 U997 ( .A(G119), .B(n1279), .ZN(G21) );
NAND2_X1 U998 ( .A1(n1350), .A2(n1331), .ZN(n1279) );
AND3_X1 U999 ( .A1(n1321), .A2(n1343), .A3(n1291), .ZN(n1331) );
INV_X1 U1000 ( .A(n1138), .ZN(n1343) );
XNOR2_X1 U1001 ( .A(G116), .B(n1284), .ZN(G18) );
NAND3_X1 U1002 ( .A1(n1137), .A2(n1146), .A3(n1350), .ZN(n1284) );
AND2_X1 U1003 ( .A1(n1162), .A2(n1322), .ZN(n1146) );
XNOR2_X1 U1004 ( .A(G113), .B(n1283), .ZN(G15) );
NAND3_X1 U1005 ( .A1(n1137), .A2(n1147), .A3(n1350), .ZN(n1283) );
AND3_X1 U1006 ( .A1(n1295), .A2(n1293), .A3(n1154), .ZN(n1350) );
INV_X1 U1007 ( .A(n1135), .ZN(n1154) );
NAND2_X1 U1008 ( .A1(n1150), .A2(n1351), .ZN(n1135) );
NOR2_X1 U1009 ( .A1(n1322), .A2(n1162), .ZN(n1147) );
INV_X1 U1010 ( .A(n1324), .ZN(n1162) );
INV_X1 U1011 ( .A(n1290), .ZN(n1137) );
NAND2_X1 U1012 ( .A1(n1138), .A2(n1321), .ZN(n1290) );
NAND3_X1 U1013 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(G12) );
NAND2_X1 U1014 ( .A1(n1286), .A2(n1355), .ZN(n1354) );
NAND2_X1 U1015 ( .A1(KEYINPUT35), .A2(n1356), .ZN(n1353) );
NAND2_X1 U1016 ( .A1(n1357), .A2(G110), .ZN(n1356) );
XNOR2_X1 U1017 ( .A(n1286), .B(KEYINPUT23), .ZN(n1357) );
NAND2_X1 U1018 ( .A1(n1358), .A2(n1359), .ZN(n1352) );
INV_X1 U1019 ( .A(KEYINPUT35), .ZN(n1359) );
NAND2_X1 U1020 ( .A1(n1360), .A2(n1361), .ZN(n1358) );
OR3_X1 U1021 ( .A1(n1355), .A2(n1286), .A3(KEYINPUT23), .ZN(n1361) );
INV_X1 U1022 ( .A(G110), .ZN(n1355) );
NAND2_X1 U1023 ( .A1(KEYINPUT23), .A2(n1286), .ZN(n1360) );
NOR3_X1 U1024 ( .A1(n1139), .A2(n1138), .A3(n1347), .ZN(n1286) );
NAND2_X1 U1025 ( .A1(n1291), .A2(n1285), .ZN(n1347) );
AND3_X1 U1026 ( .A1(n1296), .A2(n1293), .A3(n1295), .ZN(n1285) );
NOR2_X1 U1027 ( .A1(n1159), .A2(n1158), .ZN(n1295) );
AND2_X1 U1028 ( .A1(G214), .A2(n1362), .ZN(n1158) );
NAND2_X1 U1029 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
INV_X1 U1030 ( .A(n1334), .ZN(n1159) );
NAND3_X1 U1031 ( .A1(n1365), .A2(n1366), .A3(n1367), .ZN(n1334) );
NAND2_X1 U1032 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
OR3_X1 U1033 ( .A1(n1369), .A2(n1368), .A3(G902), .ZN(n1366) );
AND2_X1 U1034 ( .A1(G237), .A2(G210), .ZN(n1368) );
XOR2_X1 U1035 ( .A(n1370), .B(n1371), .Z(n1369) );
INV_X1 U1036 ( .A(n1306), .ZN(n1371) );
XNOR2_X1 U1037 ( .A(n1372), .B(n1373), .ZN(n1306) );
XOR2_X1 U1038 ( .A(n1374), .B(n1217), .Z(n1373) );
AND2_X1 U1039 ( .A1(n1375), .A2(G224), .ZN(n1374) );
XNOR2_X1 U1040 ( .A(n1215), .B(n1218), .ZN(n1372) );
XNOR2_X1 U1041 ( .A(n1376), .B(KEYINPUT39), .ZN(n1218) );
XOR2_X1 U1042 ( .A(G122), .B(n1377), .Z(n1215) );
NOR2_X1 U1043 ( .A1(KEYINPUT2), .A2(n1378), .ZN(n1377) );
XNOR2_X1 U1044 ( .A(KEYINPUT41), .B(n1379), .ZN(n1370) );
NOR2_X1 U1045 ( .A1(KEYINPUT5), .A2(n1380), .ZN(n1379) );
NOR2_X1 U1046 ( .A1(n1381), .A2(n1308), .ZN(n1380) );
AND2_X1 U1047 ( .A1(n1186), .A2(n1244), .ZN(n1308) );
NOR2_X1 U1048 ( .A1(n1186), .A2(n1244), .ZN(n1381) );
NAND2_X1 U1049 ( .A1(G902), .A2(G210), .ZN(n1365) );
NAND2_X1 U1050 ( .A1(n1144), .A2(n1382), .ZN(n1293) );
NAND4_X1 U1051 ( .A1(G953), .A2(G902), .A3(n1349), .A4(n1219), .ZN(n1382) );
INV_X1 U1052 ( .A(G898), .ZN(n1219) );
NAND3_X1 U1053 ( .A1(n1349), .A2(n1152), .A3(G952), .ZN(n1144) );
INV_X1 U1054 ( .A(G953), .ZN(n1152) );
NAND2_X1 U1055 ( .A1(G234), .A2(n1383), .ZN(n1349) );
XNOR2_X1 U1056 ( .A(KEYINPUT47), .B(n1363), .ZN(n1383) );
NOR2_X1 U1057 ( .A1(n1150), .A2(n1149), .ZN(n1296) );
INV_X1 U1058 ( .A(n1351), .ZN(n1149) );
NAND2_X1 U1059 ( .A1(G221), .A2(n1384), .ZN(n1351) );
XOR2_X1 U1060 ( .A(n1385), .B(G469), .Z(n1150) );
NAND2_X1 U1061 ( .A1(n1386), .A2(n1364), .ZN(n1385) );
XOR2_X1 U1062 ( .A(n1387), .B(n1388), .Z(n1386) );
XOR2_X1 U1063 ( .A(n1389), .B(n1255), .Z(n1388) );
AND2_X1 U1064 ( .A1(G227), .A2(n1375), .ZN(n1255) );
NAND2_X1 U1065 ( .A1(n1390), .A2(n1258), .ZN(n1389) );
NAND3_X1 U1066 ( .A1(n1193), .A2(n1263), .A3(n1391), .ZN(n1258) );
INV_X1 U1067 ( .A(n1192), .ZN(n1193) );
INV_X1 U1068 ( .A(n1264), .ZN(n1390) );
NAND2_X1 U1069 ( .A1(n1392), .A2(n1393), .ZN(n1264) );
NAND2_X1 U1070 ( .A1(n1261), .A2(n1394), .ZN(n1393) );
XNOR2_X1 U1071 ( .A(n1263), .B(n1192), .ZN(n1394) );
NAND3_X1 U1072 ( .A1(n1192), .A2(n1376), .A3(n1391), .ZN(n1392) );
INV_X1 U1073 ( .A(n1263), .ZN(n1376) );
XNOR2_X1 U1074 ( .A(n1395), .B(n1396), .ZN(n1263) );
XOR2_X1 U1075 ( .A(KEYINPUT62), .B(G107), .Z(n1396) );
XNOR2_X1 U1076 ( .A(G101), .B(G104), .ZN(n1395) );
XNOR2_X1 U1077 ( .A(n1397), .B(n1398), .ZN(n1192) );
XNOR2_X1 U1078 ( .A(G146), .B(KEYINPUT43), .ZN(n1397) );
NAND2_X1 U1079 ( .A1(n1399), .A2(n1400), .ZN(n1387) );
NAND2_X1 U1080 ( .A1(n1253), .A2(n1401), .ZN(n1400) );
INV_X1 U1081 ( .A(KEYINPUT4), .ZN(n1401) );
XNOR2_X1 U1082 ( .A(n1185), .B(n1402), .ZN(n1253) );
INV_X1 U1083 ( .A(G140), .ZN(n1185) );
NAND3_X1 U1084 ( .A1(G140), .A2(n1402), .A3(KEYINPUT4), .ZN(n1399) );
NOR2_X1 U1085 ( .A1(n1324), .A2(n1322), .ZN(n1291) );
XNOR2_X1 U1086 ( .A(n1168), .B(KEYINPUT54), .ZN(n1322) );
XNOR2_X1 U1087 ( .A(n1403), .B(G478), .ZN(n1168) );
NAND2_X1 U1088 ( .A1(n1230), .A2(n1364), .ZN(n1403) );
XNOR2_X1 U1089 ( .A(n1404), .B(n1405), .ZN(n1230) );
XOR2_X1 U1090 ( .A(n1406), .B(n1407), .Z(n1405) );
XOR2_X1 U1091 ( .A(G134), .B(G122), .Z(n1407) );
XOR2_X1 U1092 ( .A(KEYINPUT50), .B(KEYINPUT1), .Z(n1406) );
XOR2_X1 U1093 ( .A(n1408), .B(n1409), .Z(n1404) );
XOR2_X1 U1094 ( .A(G116), .B(G107), .Z(n1409) );
XOR2_X1 U1095 ( .A(n1410), .B(n1398), .Z(n1408) );
XNOR2_X1 U1096 ( .A(G143), .B(n1338), .ZN(n1398) );
NAND3_X1 U1097 ( .A1(G217), .A2(n1411), .A3(KEYINPUT19), .ZN(n1410) );
XNOR2_X1 U1098 ( .A(n1412), .B(G475), .ZN(n1324) );
OR2_X1 U1099 ( .A1(n1235), .A2(G902), .ZN(n1412) );
XNOR2_X1 U1100 ( .A(n1413), .B(n1414), .ZN(n1235) );
XOR2_X1 U1101 ( .A(n1415), .B(n1416), .Z(n1414) );
XOR2_X1 U1102 ( .A(n1417), .B(n1418), .Z(n1416) );
NOR2_X1 U1103 ( .A1(n1419), .A2(n1420), .ZN(n1418) );
XOR2_X1 U1104 ( .A(n1421), .B(KEYINPUT48), .Z(n1420) );
NAND2_X1 U1105 ( .A1(G104), .A2(n1422), .ZN(n1421) );
NOR2_X1 U1106 ( .A1(G104), .A2(n1422), .ZN(n1419) );
XOR2_X1 U1107 ( .A(G122), .B(G113), .Z(n1422) );
NAND4_X1 U1108 ( .A1(n1423), .A2(n1188), .A3(n1424), .A4(n1425), .ZN(n1417) );
OR4_X1 U1109 ( .A1(G140), .A2(KEYINPUT53), .A3(n1315), .A4(KEYINPUT37), .ZN(n1425) );
NAND2_X1 U1110 ( .A1(KEYINPUT37), .A2(G140), .ZN(n1424) );
NAND2_X1 U1111 ( .A1(KEYINPUT53), .A2(n1315), .ZN(n1423) );
NAND2_X1 U1112 ( .A1(n1426), .A2(G214), .ZN(n1415) );
XOR2_X1 U1113 ( .A(n1427), .B(n1428), .Z(n1413) );
XOR2_X1 U1114 ( .A(KEYINPUT27), .B(G146), .Z(n1428) );
XNOR2_X1 U1115 ( .A(G131), .B(G143), .ZN(n1427) );
NOR2_X1 U1116 ( .A1(n1429), .A2(n1165), .ZN(n1138) );
NOR2_X1 U1117 ( .A1(n1171), .A2(n1172), .ZN(n1165) );
AND2_X1 U1118 ( .A1(n1172), .A2(n1430), .ZN(n1429) );
XNOR2_X1 U1119 ( .A(KEYINPUT60), .B(n1171), .ZN(n1430) );
NAND2_X1 U1120 ( .A1(G217), .A2(n1384), .ZN(n1171) );
NAND2_X1 U1121 ( .A1(G234), .A2(n1364), .ZN(n1384) );
NOR2_X1 U1122 ( .A1(n1226), .A2(G902), .ZN(n1172) );
XOR2_X1 U1123 ( .A(n1431), .B(n1432), .Z(n1226) );
XNOR2_X1 U1124 ( .A(n1329), .B(n1433), .ZN(n1432) );
NOR4_X1 U1125 ( .A1(n1434), .A2(n1435), .A3(KEYINPUT51), .A4(n1436), .ZN(n1433) );
NOR2_X1 U1126 ( .A1(G140), .A2(n1437), .ZN(n1436) );
XNOR2_X1 U1127 ( .A(n1186), .B(n1438), .ZN(n1437) );
XNOR2_X1 U1128 ( .A(KEYINPUT45), .B(n1439), .ZN(n1438) );
NOR2_X1 U1129 ( .A1(n1439), .A2(n1188), .ZN(n1435) );
NAND2_X1 U1130 ( .A1(G140), .A2(n1315), .ZN(n1188) );
INV_X1 U1131 ( .A(n1186), .ZN(n1315) );
AND3_X1 U1132 ( .A1(n1439), .A2(n1186), .A3(G140), .ZN(n1434) );
XOR2_X1 U1133 ( .A(G125), .B(KEYINPUT36), .Z(n1186) );
XNOR2_X1 U1134 ( .A(G146), .B(KEYINPUT0), .ZN(n1439) );
XOR2_X1 U1135 ( .A(n1440), .B(n1441), .Z(n1431) );
AND2_X1 U1136 ( .A1(G221), .A2(n1411), .ZN(n1441) );
AND2_X1 U1137 ( .A1(G234), .A2(n1375), .ZN(n1411) );
NAND2_X1 U1138 ( .A1(n1442), .A2(n1443), .ZN(n1440) );
NAND2_X1 U1139 ( .A1(n1378), .A2(n1444), .ZN(n1443) );
XOR2_X1 U1140 ( .A(n1445), .B(KEYINPUT38), .Z(n1442) );
OR2_X1 U1141 ( .A1(n1444), .A2(n1378), .ZN(n1445) );
INV_X1 U1142 ( .A(n1402), .ZN(n1378) );
XOR2_X1 U1143 ( .A(G110), .B(KEYINPUT11), .Z(n1402) );
XOR2_X1 U1144 ( .A(G128), .B(n1446), .Z(n1444) );
XOR2_X1 U1145 ( .A(n1321), .B(KEYINPUT16), .Z(n1139) );
XNOR2_X1 U1146 ( .A(n1170), .B(n1447), .ZN(n1321) );
XOR2_X1 U1147 ( .A(KEYINPUT22), .B(G472), .Z(n1447) );
NAND2_X1 U1148 ( .A1(n1448), .A2(n1364), .ZN(n1170) );
INV_X1 U1149 ( .A(G902), .ZN(n1364) );
XNOR2_X1 U1150 ( .A(n1243), .B(n1449), .ZN(n1448) );
XOR2_X1 U1151 ( .A(n1450), .B(n1242), .Z(n1449) );
XNOR2_X1 U1152 ( .A(n1217), .B(n1391), .ZN(n1242) );
INV_X1 U1153 ( .A(n1261), .ZN(n1391) );
XNOR2_X1 U1154 ( .A(n1194), .B(n1451), .ZN(n1261) );
XNOR2_X1 U1155 ( .A(KEYINPUT61), .B(n1452), .ZN(n1451) );
INV_X1 U1156 ( .A(G131), .ZN(n1452) );
XNOR2_X1 U1157 ( .A(G134), .B(n1453), .ZN(n1194) );
XNOR2_X1 U1158 ( .A(KEYINPUT12), .B(n1329), .ZN(n1453) );
INV_X1 U1159 ( .A(G137), .ZN(n1329) );
XNOR2_X1 U1160 ( .A(n1454), .B(n1446), .ZN(n1217) );
XOR2_X1 U1161 ( .A(G119), .B(KEYINPUT17), .Z(n1446) );
XNOR2_X1 U1162 ( .A(G116), .B(G113), .ZN(n1454) );
NAND2_X1 U1163 ( .A1(KEYINPUT8), .A2(n1244), .ZN(n1450) );
NAND3_X1 U1164 ( .A1(n1455), .A2(n1456), .A3(n1457), .ZN(n1244) );
OR2_X1 U1165 ( .A1(n1338), .A2(n1458), .ZN(n1457) );
NAND3_X1 U1166 ( .A1(n1458), .A2(n1338), .A3(KEYINPUT30), .ZN(n1456) );
INV_X1 U1167 ( .A(G128), .ZN(n1338) );
NOR2_X1 U1168 ( .A1(KEYINPUT32), .A2(n1459), .ZN(n1458) );
NAND2_X1 U1169 ( .A1(n1459), .A2(n1460), .ZN(n1455) );
INV_X1 U1170 ( .A(KEYINPUT30), .ZN(n1460) );
XOR2_X1 U1171 ( .A(n1461), .B(G143), .Z(n1459) );
NAND2_X1 U1172 ( .A1(KEYINPUT14), .A2(G146), .ZN(n1461) );
XOR2_X1 U1173 ( .A(n1462), .B(n1345), .Z(n1243) );
INV_X1 U1174 ( .A(G101), .ZN(n1345) );
NAND2_X1 U1175 ( .A1(n1426), .A2(G210), .ZN(n1462) );
AND2_X1 U1176 ( .A1(n1375), .A2(n1363), .ZN(n1426) );
INV_X1 U1177 ( .A(G237), .ZN(n1363) );
XNOR2_X1 U1178 ( .A(G953), .B(KEYINPUT55), .ZN(n1375) );
endmodule


