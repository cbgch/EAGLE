//Key = 1001000101101010000001111011011000001111000000011100000101101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414, n1415;

NAND2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(G9) );
NAND2_X1 U779 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U780 ( .A(KEYINPUT29), .B(n1085), .Z(n1081) );
NOR2_X1 U781 ( .A1(n1083), .A2(n1084), .ZN(n1085) );
INV_X1 U782 ( .A(G107), .ZN(n1084) );
NOR2_X1 U783 ( .A1(n1086), .A2(n1087), .ZN(G75) );
NOR3_X1 U784 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1087) );
NOR2_X1 U785 ( .A1(KEYINPUT62), .A2(n1091), .ZN(n1089) );
AND4_X1 U786 ( .A1(n1092), .A2(KEYINPUT26), .A3(n1093), .A4(n1094), .ZN(n1091) );
AND3_X1 U787 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1092) );
NAND3_X1 U788 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1088) );
NAND3_X1 U789 ( .A1(n1101), .A2(n1096), .A3(KEYINPUT26), .ZN(n1100) );
NAND2_X1 U790 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND3_X1 U791 ( .A1(n1097), .A2(n1104), .A3(n1093), .ZN(n1103) );
NAND2_X1 U792 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U793 ( .A1(n1094), .A2(n1107), .ZN(n1106) );
NAND2_X1 U794 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U795 ( .A1(KEYINPUT62), .A2(n1095), .ZN(n1109) );
NAND2_X1 U796 ( .A1(n1110), .A2(n1111), .ZN(n1105) );
NAND2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U798 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND3_X1 U799 ( .A1(n1110), .A2(n1116), .A3(n1094), .ZN(n1102) );
NAND2_X1 U800 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U801 ( .A1(n1093), .A2(n1119), .ZN(n1118) );
NAND2_X1 U802 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U803 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U804 ( .A1(n1097), .A2(n1124), .ZN(n1117) );
NAND2_X1 U805 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
AND3_X1 U807 ( .A1(n1098), .A2(n1099), .A3(n1129), .ZN(n1086) );
NAND4_X1 U808 ( .A1(n1130), .A2(n1093), .A3(n1131), .A4(n1132), .ZN(n1098) );
NOR4_X1 U809 ( .A1(n1133), .A2(n1114), .A3(n1134), .A4(n1123), .ZN(n1132) );
XOR2_X1 U810 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U811 ( .A1(n1137), .A2(KEYINPUT13), .ZN(n1136) );
NOR3_X1 U812 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1131) );
AND3_X1 U813 ( .A1(KEYINPUT36), .A2(n1141), .A3(G478), .ZN(n1140) );
NOR2_X1 U814 ( .A1(KEYINPUT36), .A2(G478), .ZN(n1139) );
XOR2_X1 U815 ( .A(n1142), .B(n1143), .Z(n1138) );
NAND3_X1 U816 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(G72) );
NAND2_X1 U817 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U818 ( .A1(n1149), .A2(n1150), .ZN(n1147) );
XOR2_X1 U819 ( .A(n1151), .B(n1152), .Z(n1149) );
NAND2_X1 U820 ( .A1(KEYINPUT58), .A2(n1153), .ZN(n1152) );
OR4_X1 U821 ( .A1(n1151), .A2(KEYINPUT25), .A3(n1148), .A4(n1153), .ZN(n1145) );
NAND4_X1 U822 ( .A1(n1154), .A2(n1150), .A3(n1155), .A4(n1153), .ZN(n1144) );
NAND2_X1 U823 ( .A1(n1156), .A2(n1157), .ZN(n1153) );
NAND2_X1 U824 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XNOR2_X1 U825 ( .A(KEYINPUT44), .B(n1160), .ZN(n1159) );
INV_X1 U826 ( .A(n1161), .ZN(n1158) );
XOR2_X1 U827 ( .A(n1099), .B(KEYINPUT15), .Z(n1156) );
INV_X1 U828 ( .A(n1148), .ZN(n1155) );
NAND2_X1 U829 ( .A1(G953), .A2(n1162), .ZN(n1148) );
NAND2_X1 U830 ( .A1(G900), .A2(G227), .ZN(n1162) );
INV_X1 U831 ( .A(KEYINPUT25), .ZN(n1150) );
XNOR2_X1 U832 ( .A(KEYINPUT58), .B(n1151), .ZN(n1154) );
NAND2_X1 U833 ( .A1(n1163), .A2(n1164), .ZN(n1151) );
NAND2_X1 U834 ( .A1(G953), .A2(n1165), .ZN(n1164) );
XOR2_X1 U835 ( .A(n1166), .B(n1167), .Z(n1163) );
XOR2_X1 U836 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U837 ( .A(n1170), .B(n1171), .Z(n1166) );
XOR2_X1 U838 ( .A(KEYINPUT8), .B(G134), .Z(n1171) );
XOR2_X1 U839 ( .A(n1172), .B(n1173), .Z(G69) );
XOR2_X1 U840 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR3_X1 U841 ( .A1(n1176), .A2(KEYINPUT63), .A3(G953), .ZN(n1175) );
NOR3_X1 U842 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1176) );
INV_X1 U843 ( .A(n1180), .ZN(n1178) );
XOR2_X1 U844 ( .A(KEYINPUT11), .B(n1181), .Z(n1177) );
NAND2_X1 U845 ( .A1(n1182), .A2(n1183), .ZN(n1174) );
NAND2_X1 U846 ( .A1(G953), .A2(n1184), .ZN(n1183) );
XNOR2_X1 U847 ( .A(n1185), .B(n1186), .ZN(n1182) );
XNOR2_X1 U848 ( .A(KEYINPUT4), .B(n1187), .ZN(n1186) );
NOR2_X1 U849 ( .A1(n1188), .A2(KEYINPUT28), .ZN(n1187) );
NOR2_X1 U850 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U851 ( .A(KEYINPUT59), .B(n1191), .Z(n1190) );
NOR2_X1 U852 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
AND2_X1 U853 ( .A1(n1192), .A2(n1193), .ZN(n1189) );
NAND2_X1 U854 ( .A1(G953), .A2(n1194), .ZN(n1172) );
NAND2_X1 U855 ( .A1(G898), .A2(G224), .ZN(n1194) );
NOR2_X1 U856 ( .A1(n1195), .A2(n1196), .ZN(G66) );
XOR2_X1 U857 ( .A(n1197), .B(n1198), .Z(n1196) );
NOR2_X1 U858 ( .A1(n1199), .A2(n1200), .ZN(n1197) );
NOR2_X1 U859 ( .A1(n1195), .A2(n1201), .ZN(G63) );
XOR2_X1 U860 ( .A(n1202), .B(n1203), .Z(n1201) );
AND2_X1 U861 ( .A1(G478), .A2(n1204), .ZN(n1202) );
NOR2_X1 U862 ( .A1(n1195), .A2(n1205), .ZN(G60) );
NOR3_X1 U863 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1205) );
NOR3_X1 U864 ( .A1(n1209), .A2(n1142), .A3(n1200), .ZN(n1208) );
NOR2_X1 U865 ( .A1(n1210), .A2(n1211), .ZN(n1207) );
AND2_X1 U866 ( .A1(n1090), .A2(G475), .ZN(n1210) );
XOR2_X1 U867 ( .A(G104), .B(n1212), .Z(G6) );
NOR2_X1 U868 ( .A1(n1195), .A2(n1213), .ZN(G57) );
XOR2_X1 U869 ( .A(n1214), .B(n1215), .Z(n1213) );
XOR2_X1 U870 ( .A(G101), .B(n1216), .Z(n1215) );
NAND2_X1 U871 ( .A1(n1217), .A2(n1218), .ZN(n1214) );
OR2_X1 U872 ( .A1(n1219), .A2(KEYINPUT24), .ZN(n1218) );
XOR2_X1 U873 ( .A(n1220), .B(n1221), .Z(n1217) );
NOR2_X1 U874 ( .A1(n1135), .A2(n1200), .ZN(n1221) );
INV_X1 U875 ( .A(G472), .ZN(n1135) );
NAND2_X1 U876 ( .A1(KEYINPUT24), .A2(n1219), .ZN(n1220) );
XOR2_X1 U877 ( .A(n1222), .B(n1223), .Z(n1219) );
NOR3_X1 U878 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(G54) );
AND2_X1 U879 ( .A1(KEYINPUT23), .A2(n1195), .ZN(n1226) );
NOR3_X1 U880 ( .A1(KEYINPUT23), .A2(n1099), .A3(n1129), .ZN(n1225) );
INV_X1 U881 ( .A(G952), .ZN(n1129) );
XOR2_X1 U882 ( .A(n1227), .B(n1228), .Z(n1224) );
XOR2_X1 U883 ( .A(n1229), .B(n1230), .Z(n1228) );
NAND2_X1 U884 ( .A1(KEYINPUT47), .A2(n1223), .ZN(n1230) );
NAND2_X1 U885 ( .A1(n1231), .A2(n1232), .ZN(n1229) );
NAND2_X1 U886 ( .A1(n1233), .A2(n1234), .ZN(n1231) );
NAND2_X1 U887 ( .A1(G227), .A2(n1099), .ZN(n1234) );
XOR2_X1 U888 ( .A(n1235), .B(n1236), .Z(n1227) );
AND2_X1 U889 ( .A1(G469), .A2(n1204), .ZN(n1236) );
NOR2_X1 U890 ( .A1(n1195), .A2(n1237), .ZN(G51) );
XOR2_X1 U891 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U892 ( .A(n1240), .B(n1241), .Z(n1238) );
NOR2_X1 U893 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U894 ( .A(KEYINPUT56), .B(n1244), .Z(n1243) );
NAND3_X1 U895 ( .A1(n1204), .A2(n1245), .A3(KEYINPUT0), .ZN(n1240) );
INV_X1 U896 ( .A(n1200), .ZN(n1204) );
NAND2_X1 U897 ( .A1(G902), .A2(n1090), .ZN(n1200) );
NAND3_X1 U898 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1090) );
NOR3_X1 U899 ( .A1(n1161), .A2(n1181), .A3(n1160), .ZN(n1248) );
NAND4_X1 U900 ( .A1(n1249), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1160) );
AND2_X1 U901 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NAND3_X1 U902 ( .A1(n1093), .A2(n1255), .A3(n1256), .ZN(n1251) );
XOR2_X1 U903 ( .A(KEYINPUT20), .B(n1257), .Z(n1255) );
NAND2_X1 U904 ( .A1(n1258), .A2(n1259), .ZN(n1250) );
INV_X1 U905 ( .A(KEYINPUT45), .ZN(n1259) );
NAND4_X1 U906 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(KEYINPUT45), .ZN(n1249) );
NAND4_X1 U907 ( .A1(n1263), .A2(n1264), .A3(n1265), .A4(n1266), .ZN(n1161) );
INV_X1 U908 ( .A(n1179), .ZN(n1247) );
NAND4_X1 U909 ( .A1(n1267), .A2(n1268), .A3(n1269), .A4(n1270), .ZN(n1179) );
NOR3_X1 U910 ( .A1(n1083), .A2(n1271), .A3(n1212), .ZN(n1270) );
NOR3_X1 U911 ( .A1(n1272), .A2(n1273), .A3(n1108), .ZN(n1212) );
AND3_X1 U912 ( .A1(n1095), .A2(n1274), .A3(n1097), .ZN(n1083) );
NAND3_X1 U913 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1269) );
INV_X1 U914 ( .A(KEYINPUT42), .ZN(n1276) );
NAND4_X1 U915 ( .A1(n1278), .A2(n1279), .A3(n1097), .A4(n1280), .ZN(n1268) );
NAND3_X1 U916 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1267) );
NAND2_X1 U917 ( .A1(n1284), .A2(n1285), .ZN(n1282) );
NAND4_X1 U918 ( .A1(KEYINPUT42), .A2(n1275), .A3(n1286), .A4(n1287), .ZN(n1285) );
NAND2_X1 U919 ( .A1(n1122), .A2(n1273), .ZN(n1281) );
XOR2_X1 U920 ( .A(n1180), .B(KEYINPUT51), .Z(n1246) );
NOR2_X1 U921 ( .A1(n1099), .A2(G952), .ZN(n1195) );
XOR2_X1 U922 ( .A(n1258), .B(n1288), .Z(G48) );
NOR2_X1 U923 ( .A1(KEYINPUT17), .A2(n1289), .ZN(n1288) );
INV_X1 U924 ( .A(G146), .ZN(n1289) );
AND3_X1 U925 ( .A1(n1261), .A2(n1290), .A3(n1260), .ZN(n1258) );
XNOR2_X1 U926 ( .A(G143), .B(n1254), .ZN(G45) );
NAND3_X1 U927 ( .A1(n1278), .A2(n1291), .A3(n1292), .ZN(n1254) );
NOR3_X1 U928 ( .A1(n1120), .A2(n1293), .A3(n1262), .ZN(n1292) );
INV_X1 U929 ( .A(n1290), .ZN(n1262) );
INV_X1 U930 ( .A(n1294), .ZN(n1120) );
XNOR2_X1 U931 ( .A(G140), .B(n1295), .ZN(G42) );
NAND2_X1 U932 ( .A1(n1093), .A2(n1296), .ZN(n1295) );
XOR2_X1 U933 ( .A(KEYINPUT19), .B(n1297), .Z(n1296) );
NOR2_X1 U934 ( .A1(n1112), .A2(n1298), .ZN(n1297) );
XNOR2_X1 U935 ( .A(G137), .B(n1253), .ZN(G39) );
NAND3_X1 U936 ( .A1(n1283), .A2(n1284), .A3(n1299), .ZN(n1253) );
INV_X1 U937 ( .A(n1300), .ZN(n1283) );
XOR2_X1 U938 ( .A(n1301), .B(G134), .Z(G36) );
NAND2_X1 U939 ( .A1(KEYINPUT9), .A2(n1266), .ZN(n1301) );
NAND3_X1 U940 ( .A1(n1095), .A2(n1294), .A3(n1299), .ZN(n1266) );
XNOR2_X1 U941 ( .A(G131), .B(n1263), .ZN(G33) );
NAND3_X1 U942 ( .A1(n1261), .A2(n1294), .A3(n1299), .ZN(n1263) );
AND3_X1 U943 ( .A1(n1257), .A2(n1290), .A3(n1093), .ZN(n1299) );
NOR2_X1 U944 ( .A1(n1302), .A2(n1127), .ZN(n1093) );
INV_X1 U945 ( .A(n1128), .ZN(n1302) );
XNOR2_X1 U946 ( .A(G128), .B(n1264), .ZN(G30) );
NAND3_X1 U947 ( .A1(n1095), .A2(n1290), .A3(n1260), .ZN(n1264) );
AND3_X1 U948 ( .A1(n1284), .A2(n1123), .A3(n1291), .ZN(n1260) );
XOR2_X1 U949 ( .A(n1181), .B(n1303), .Z(G3) );
NOR2_X1 U950 ( .A1(KEYINPUT5), .A2(n1304), .ZN(n1303) );
AND3_X1 U951 ( .A1(n1274), .A2(n1294), .A3(n1110), .ZN(n1181) );
INV_X1 U952 ( .A(n1273), .ZN(n1274) );
XNOR2_X1 U953 ( .A(G125), .B(n1265), .ZN(G27) );
NAND3_X1 U954 ( .A1(n1094), .A2(n1275), .A3(n1256), .ZN(n1265) );
INV_X1 U955 ( .A(n1298), .ZN(n1256) );
NAND4_X1 U956 ( .A1(n1122), .A2(n1261), .A3(n1123), .A4(n1290), .ZN(n1298) );
NAND2_X1 U957 ( .A1(n1305), .A2(n1306), .ZN(n1290) );
NAND2_X1 U958 ( .A1(n1307), .A2(n1165), .ZN(n1306) );
INV_X1 U959 ( .A(G900), .ZN(n1165) );
XNOR2_X1 U960 ( .A(G122), .B(n1308), .ZN(G24) );
NAND4_X1 U961 ( .A1(n1278), .A2(n1094), .A3(n1309), .A4(n1310), .ZN(n1308) );
NOR3_X1 U962 ( .A1(n1272), .A2(n1311), .A3(n1293), .ZN(n1310) );
INV_X1 U963 ( .A(n1097), .ZN(n1272) );
XOR2_X1 U964 ( .A(n1125), .B(KEYINPUT14), .Z(n1309) );
INV_X1 U965 ( .A(n1286), .ZN(n1094) );
NAND2_X1 U966 ( .A1(n1312), .A2(n1313), .ZN(G21) );
OR2_X1 U967 ( .A1(n1314), .A2(G119), .ZN(n1313) );
XOR2_X1 U968 ( .A(n1315), .B(KEYINPUT33), .Z(n1312) );
NAND2_X1 U969 ( .A1(G119), .A2(n1314), .ZN(n1315) );
NAND2_X1 U970 ( .A1(n1275), .A2(n1316), .ZN(n1314) );
XOR2_X1 U971 ( .A(KEYINPUT54), .B(n1277), .Z(n1316) );
NOR4_X1 U972 ( .A1(n1300), .A2(n1286), .A3(n1122), .A4(n1311), .ZN(n1277) );
XOR2_X1 U973 ( .A(n1317), .B(n1180), .Z(G18) );
NAND3_X1 U974 ( .A1(n1095), .A2(n1294), .A3(n1279), .ZN(n1180) );
NOR2_X1 U975 ( .A1(n1278), .A2(n1293), .ZN(n1095) );
XOR2_X1 U976 ( .A(G113), .B(n1271), .Z(G15) );
AND3_X1 U977 ( .A1(n1279), .A2(n1294), .A3(n1261), .ZN(n1271) );
INV_X1 U978 ( .A(n1108), .ZN(n1261) );
NAND2_X1 U979 ( .A1(n1278), .A2(n1293), .ZN(n1108) );
NAND2_X1 U980 ( .A1(n1318), .A2(n1319), .ZN(n1294) );
OR3_X1 U981 ( .A1(n1122), .A2(n1123), .A3(KEYINPUT2), .ZN(n1319) );
INV_X1 U982 ( .A(n1284), .ZN(n1122) );
NAND2_X1 U983 ( .A1(KEYINPUT2), .A2(n1097), .ZN(n1318) );
NOR2_X1 U984 ( .A1(n1123), .A2(n1284), .ZN(n1097) );
NOR3_X1 U985 ( .A1(n1125), .A2(n1311), .A3(n1286), .ZN(n1279) );
NAND2_X1 U986 ( .A1(n1115), .A2(n1320), .ZN(n1286) );
INV_X1 U987 ( .A(n1287), .ZN(n1311) );
XNOR2_X1 U988 ( .A(G110), .B(n1321), .ZN(G12) );
NOR2_X1 U989 ( .A1(KEYINPUT31), .A2(n1322), .ZN(n1321) );
NOR3_X1 U990 ( .A1(n1300), .A2(n1273), .A3(n1284), .ZN(n1322) );
XOR2_X1 U991 ( .A(n1137), .B(G472), .Z(n1284) );
AND2_X1 U992 ( .A1(n1323), .A2(n1324), .ZN(n1137) );
XOR2_X1 U993 ( .A(n1325), .B(n1326), .Z(n1323) );
XOR2_X1 U994 ( .A(n1327), .B(n1222), .Z(n1326) );
XOR2_X1 U995 ( .A(n1328), .B(n1329), .Z(n1222) );
XOR2_X1 U996 ( .A(G113), .B(n1330), .Z(n1329) );
XOR2_X1 U997 ( .A(KEYINPUT53), .B(G116), .Z(n1330) );
XOR2_X1 U998 ( .A(n1331), .B(n1332), .Z(n1328) );
NAND2_X1 U999 ( .A1(KEYINPUT27), .A2(G119), .ZN(n1331) );
NAND2_X1 U1000 ( .A1(KEYINPUT12), .A2(n1223), .ZN(n1327) );
XOR2_X1 U1001 ( .A(KEYINPUT43), .B(n1333), .Z(n1325) );
NOR2_X1 U1002 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
XOR2_X1 U1003 ( .A(KEYINPUT40), .B(n1336), .Z(n1335) );
NOR2_X1 U1004 ( .A1(n1337), .A2(n1304), .ZN(n1336) );
NOR2_X1 U1005 ( .A1(G101), .A2(n1216), .ZN(n1334) );
INV_X1 U1006 ( .A(n1337), .ZN(n1216) );
NAND2_X1 U1007 ( .A1(G210), .A2(n1338), .ZN(n1337) );
NAND2_X1 U1008 ( .A1(n1291), .A2(n1287), .ZN(n1273) );
NAND2_X1 U1009 ( .A1(n1305), .A2(n1339), .ZN(n1287) );
NAND2_X1 U1010 ( .A1(n1307), .A2(n1184), .ZN(n1339) );
INV_X1 U1011 ( .A(G898), .ZN(n1184) );
AND3_X1 U1012 ( .A1(G902), .A2(n1096), .A3(G953), .ZN(n1307) );
NAND3_X1 U1013 ( .A1(n1096), .A2(n1099), .A3(G952), .ZN(n1305) );
NAND2_X1 U1014 ( .A1(G237), .A2(G234), .ZN(n1096) );
NOR2_X1 U1015 ( .A1(n1125), .A2(n1112), .ZN(n1291) );
INV_X1 U1016 ( .A(n1257), .ZN(n1112) );
NOR2_X1 U1017 ( .A1(n1115), .A2(n1114), .ZN(n1257) );
INV_X1 U1018 ( .A(n1320), .ZN(n1114) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1340), .ZN(n1320) );
XNOR2_X1 U1020 ( .A(n1130), .B(KEYINPUT48), .ZN(n1115) );
XOR2_X1 U1021 ( .A(n1341), .B(G469), .Z(n1130) );
NAND2_X1 U1022 ( .A1(n1342), .A2(n1324), .ZN(n1341) );
XNOR2_X1 U1023 ( .A(n1343), .B(n1223), .ZN(n1342) );
XOR2_X1 U1024 ( .A(n1344), .B(G131), .Z(n1223) );
NAND3_X1 U1025 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1344) );
NAND2_X1 U1026 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
NAND2_X1 U1027 ( .A1(n1350), .A2(KEYINPUT10), .ZN(n1349) );
XOR2_X1 U1028 ( .A(n1351), .B(KEYINPUT50), .Z(n1350) );
NAND3_X1 U1029 ( .A1(KEYINPUT10), .A2(n1352), .A3(n1351), .ZN(n1346) );
OR2_X1 U1030 ( .A1(n1351), .A2(KEYINPUT10), .ZN(n1345) );
INV_X1 U1031 ( .A(G134), .ZN(n1351) );
XOR2_X1 U1032 ( .A(n1235), .B(n1353), .Z(n1343) );
NOR2_X1 U1033 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NOR2_X1 U1034 ( .A1(KEYINPUT61), .A2(n1232), .ZN(n1355) );
NAND3_X1 U1035 ( .A1(G227), .A2(n1099), .A3(n1356), .ZN(n1232) );
NOR2_X1 U1036 ( .A1(n1357), .A2(n1356), .ZN(n1354) );
INV_X1 U1037 ( .A(n1233), .ZN(n1356) );
XOR2_X1 U1038 ( .A(G110), .B(G140), .Z(n1233) );
NOR3_X1 U1039 ( .A1(n1358), .A2(KEYINPUT61), .A3(G953), .ZN(n1357) );
INV_X1 U1040 ( .A(G227), .ZN(n1358) );
XOR2_X1 U1041 ( .A(n1359), .B(n1360), .Z(n1235) );
XOR2_X1 U1042 ( .A(n1170), .B(n1361), .Z(n1359) );
NOR2_X1 U1043 ( .A1(KEYINPUT1), .A2(n1362), .ZN(n1361) );
XNOR2_X1 U1044 ( .A(n1332), .B(KEYINPUT39), .ZN(n1170) );
INV_X1 U1045 ( .A(n1275), .ZN(n1125) );
NOR2_X1 U1046 ( .A1(n1128), .A2(n1127), .ZN(n1275) );
AND2_X1 U1047 ( .A1(G214), .A2(n1363), .ZN(n1127) );
XOR2_X1 U1048 ( .A(n1364), .B(n1245), .Z(n1128) );
AND2_X1 U1049 ( .A1(G210), .A2(n1363), .ZN(n1245) );
OR2_X1 U1050 ( .A1(G902), .A2(G237), .ZN(n1363) );
NAND2_X1 U1051 ( .A1(n1365), .A2(n1324), .ZN(n1364) );
XOR2_X1 U1052 ( .A(n1366), .B(n1239), .Z(n1365) );
XNOR2_X1 U1053 ( .A(n1367), .B(n1185), .ZN(n1239) );
XNOR2_X1 U1054 ( .A(n1368), .B(n1369), .ZN(n1185) );
XOR2_X1 U1055 ( .A(G122), .B(G110), .Z(n1369) );
XNOR2_X1 U1056 ( .A(KEYINPUT46), .B(KEYINPUT41), .ZN(n1368) );
XOR2_X1 U1057 ( .A(n1193), .B(n1192), .Z(n1367) );
NAND2_X1 U1058 ( .A1(n1370), .A2(n1371), .ZN(n1192) );
NAND2_X1 U1059 ( .A1(G113), .A2(n1372), .ZN(n1371) );
XOR2_X1 U1060 ( .A(KEYINPUT3), .B(n1373), .Z(n1370) );
NOR2_X1 U1061 ( .A1(G113), .A2(n1372), .ZN(n1373) );
XOR2_X1 U1062 ( .A(G116), .B(n1374), .Z(n1372) );
XOR2_X1 U1063 ( .A(KEYINPUT16), .B(G119), .Z(n1374) );
XOR2_X1 U1064 ( .A(n1360), .B(n1362), .Z(n1193) );
XNOR2_X1 U1065 ( .A(n1375), .B(KEYINPUT18), .ZN(n1362) );
XNOR2_X1 U1066 ( .A(n1304), .B(n1376), .ZN(n1360) );
INV_X1 U1067 ( .A(G101), .ZN(n1304) );
NOR2_X1 U1068 ( .A1(n1244), .A2(n1242), .ZN(n1366) );
AND3_X1 U1069 ( .A1(G224), .A2(n1099), .A3(n1377), .ZN(n1242) );
XNOR2_X1 U1070 ( .A(n1332), .B(G125), .ZN(n1377) );
AND2_X1 U1071 ( .A1(n1378), .A2(n1379), .ZN(n1244) );
NAND2_X1 U1072 ( .A1(G224), .A2(n1099), .ZN(n1379) );
XOR2_X1 U1073 ( .A(G125), .B(n1332), .Z(n1378) );
XOR2_X1 U1074 ( .A(G143), .B(n1380), .Z(n1332) );
NAND2_X1 U1075 ( .A1(n1110), .A2(n1123), .ZN(n1300) );
XOR2_X1 U1076 ( .A(n1381), .B(n1199), .Z(n1123) );
NAND2_X1 U1077 ( .A1(G217), .A2(n1340), .ZN(n1199) );
NAND2_X1 U1078 ( .A1(G234), .A2(n1324), .ZN(n1340) );
OR2_X1 U1079 ( .A1(n1198), .A2(G902), .ZN(n1381) );
XNOR2_X1 U1080 ( .A(n1382), .B(n1383), .ZN(n1198) );
XOR2_X1 U1081 ( .A(n1384), .B(n1385), .Z(n1383) );
XNOR2_X1 U1082 ( .A(G110), .B(G119), .ZN(n1385) );
NAND2_X1 U1083 ( .A1(G221), .A2(n1386), .ZN(n1384) );
XNOR2_X1 U1084 ( .A(n1169), .B(n1387), .ZN(n1382) );
XNOR2_X1 U1085 ( .A(n1388), .B(n1380), .ZN(n1387) );
XOR2_X1 U1086 ( .A(G128), .B(G146), .Z(n1380) );
NAND2_X1 U1087 ( .A1(KEYINPUT60), .A2(G140), .ZN(n1388) );
XOR2_X1 U1088 ( .A(G125), .B(n1348), .Z(n1169) );
INV_X1 U1089 ( .A(n1352), .ZN(n1348) );
XNOR2_X1 U1090 ( .A(G137), .B(KEYINPUT49), .ZN(n1352) );
NOR2_X1 U1091 ( .A1(n1280), .A2(n1278), .ZN(n1110) );
AND2_X1 U1092 ( .A1(n1389), .A2(n1390), .ZN(n1278) );
NAND2_X1 U1093 ( .A1(n1391), .A2(n1142), .ZN(n1390) );
INV_X1 U1094 ( .A(G475), .ZN(n1142) );
XOR2_X1 U1095 ( .A(KEYINPUT37), .B(n1206), .Z(n1391) );
NAND2_X1 U1096 ( .A1(n1392), .A2(G475), .ZN(n1389) );
XOR2_X1 U1097 ( .A(KEYINPUT35), .B(n1206), .Z(n1392) );
INV_X1 U1098 ( .A(n1143), .ZN(n1206) );
NAND2_X1 U1099 ( .A1(n1209), .A2(n1324), .ZN(n1143) );
INV_X1 U1100 ( .A(G902), .ZN(n1324) );
INV_X1 U1101 ( .A(n1211), .ZN(n1209) );
XOR2_X1 U1102 ( .A(n1393), .B(n1394), .Z(n1211) );
XOR2_X1 U1103 ( .A(n1395), .B(n1396), .Z(n1394) );
XOR2_X1 U1104 ( .A(n1397), .B(G146), .Z(n1396) );
NAND2_X1 U1105 ( .A1(KEYINPUT21), .A2(n1398), .ZN(n1397) );
XNOR2_X1 U1106 ( .A(n1375), .B(n1399), .ZN(n1398) );
XOR2_X1 U1107 ( .A(G122), .B(G113), .Z(n1399) );
XNOR2_X1 U1108 ( .A(G104), .B(KEYINPUT6), .ZN(n1375) );
NAND2_X1 U1109 ( .A1(KEYINPUT38), .A2(n1400), .ZN(n1395) );
XOR2_X1 U1110 ( .A(n1401), .B(n1402), .Z(n1400) );
NOR2_X1 U1111 ( .A1(G143), .A2(n1403), .ZN(n1402) );
XOR2_X1 U1112 ( .A(KEYINPUT57), .B(KEYINPUT55), .Z(n1403) );
AND2_X1 U1113 ( .A1(n1338), .A2(G214), .ZN(n1401) );
AND2_X1 U1114 ( .A1(n1404), .A2(n1099), .ZN(n1338) );
XOR2_X1 U1115 ( .A(KEYINPUT30), .B(G237), .Z(n1404) );
XNOR2_X1 U1116 ( .A(n1168), .B(n1405), .ZN(n1393) );
NOR2_X1 U1117 ( .A1(G125), .A2(KEYINPUT34), .ZN(n1405) );
XOR2_X1 U1118 ( .A(G131), .B(G140), .Z(n1168) );
INV_X1 U1119 ( .A(n1293), .ZN(n1280) );
NOR2_X1 U1120 ( .A1(n1133), .A2(n1406), .ZN(n1293) );
AND2_X1 U1121 ( .A1(G478), .A2(n1141), .ZN(n1406) );
NOR2_X1 U1122 ( .A1(n1141), .A2(G478), .ZN(n1133) );
OR2_X1 U1123 ( .A1(n1203), .A2(G902), .ZN(n1141) );
XNOR2_X1 U1124 ( .A(n1407), .B(n1408), .ZN(n1203) );
AND2_X1 U1125 ( .A1(G217), .A2(n1386), .ZN(n1408) );
AND2_X1 U1126 ( .A1(G234), .A2(n1099), .ZN(n1386) );
INV_X1 U1127 ( .A(G953), .ZN(n1099) );
NAND2_X1 U1128 ( .A1(n1409), .A2(KEYINPUT22), .ZN(n1407) );
XOR2_X1 U1129 ( .A(n1410), .B(n1376), .Z(n1409) );
XOR2_X1 U1130 ( .A(G107), .B(KEYINPUT7), .Z(n1376) );
XNOR2_X1 U1131 ( .A(n1411), .B(n1412), .ZN(n1410) );
NOR2_X1 U1132 ( .A1(KEYINPUT32), .A2(n1413), .ZN(n1412) );
XOR2_X1 U1133 ( .A(G128), .B(n1414), .Z(n1413) );
XOR2_X1 U1134 ( .A(G143), .B(G134), .Z(n1414) );
NOR2_X1 U1135 ( .A1(KEYINPUT52), .A2(n1415), .ZN(n1411) );
XOR2_X1 U1136 ( .A(n1317), .B(G122), .Z(n1415) );
INV_X1 U1137 ( .A(G116), .ZN(n1317) );
endmodule


