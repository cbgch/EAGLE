//Key = 1010001111110111100000010000111111001100010001110011000010110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361;

XNOR2_X1 U742 ( .A(G107), .B(n1026), .ZN(G9) );
NAND4_X1 U743 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
NOR2_X1 U744 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
XNOR2_X1 U745 ( .A(n1033), .B(KEYINPUT54), .ZN(n1032) );
NOR2_X1 U746 ( .A1(n1034), .A2(n1035), .ZN(G75) );
NOR4_X1 U747 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
XOR2_X1 U748 ( .A(n1040), .B(KEYINPUT49), .Z(n1039) );
NAND2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND4_X1 U750 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
OR2_X1 U751 ( .A1(n1047), .A2(n1028), .ZN(n1046) );
NAND2_X1 U752 ( .A1(n1048), .A2(n1047), .ZN(n1045) );
NAND2_X1 U753 ( .A1(n1049), .A2(n1050), .ZN(n1041) );
NAND2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND3_X1 U755 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NAND2_X1 U756 ( .A1(n1056), .A2(n1030), .ZN(n1051) );
INV_X1 U757 ( .A(n1057), .ZN(n1049) );
NOR2_X1 U758 ( .A1(n1058), .A2(n1057), .ZN(n1038) );
NAND4_X1 U759 ( .A1(n1043), .A2(n1059), .A3(n1028), .A4(n1047), .ZN(n1057) );
INV_X1 U760 ( .A(n1060), .ZN(n1059) );
NOR2_X1 U761 ( .A1(n1061), .A2(n1062), .ZN(n1058) );
NOR2_X1 U762 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U763 ( .A1(n1065), .A2(n1066), .ZN(n1061) );
INV_X1 U764 ( .A(n1067), .ZN(n1037) );
NAND3_X1 U765 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1036) );
NAND2_X1 U766 ( .A1(n1044), .A2(n1071), .ZN(n1070) );
NAND2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND3_X1 U768 ( .A1(n1074), .A2(n1047), .A3(n1043), .ZN(n1073) );
NAND2_X1 U769 ( .A1(n1028), .A2(n1033), .ZN(n1072) );
NOR3_X1 U770 ( .A1(n1065), .A2(n1063), .A3(n1060), .ZN(n1044) );
INV_X1 U771 ( .A(n1053), .ZN(n1063) );
NOR3_X1 U772 ( .A1(n1075), .A2(G953), .A3(G952), .ZN(n1034) );
INV_X1 U773 ( .A(n1068), .ZN(n1075) );
NAND4_X1 U774 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1068) );
NOR4_X1 U775 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1055), .ZN(n1079) );
NAND2_X1 U776 ( .A1(n1083), .A2(n1047), .ZN(n1080) );
NOR3_X1 U777 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1078) );
XNOR2_X1 U778 ( .A(n1087), .B(n1088), .ZN(n1085) );
NOR2_X1 U779 ( .A1(n1089), .A2(KEYINPUT57), .ZN(n1088) );
XOR2_X1 U780 ( .A(n1090), .B(n1091), .Z(n1077) );
XOR2_X1 U781 ( .A(KEYINPUT53), .B(G469), .Z(n1091) );
XNOR2_X1 U782 ( .A(n1092), .B(KEYINPUT34), .ZN(n1076) );
XOR2_X1 U783 ( .A(n1093), .B(n1094), .Z(G72) );
XOR2_X1 U784 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U785 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U786 ( .A(n1099), .B(n1100), .Z(n1098) );
XNOR2_X1 U787 ( .A(KEYINPUT30), .B(n1101), .ZN(n1100) );
NOR2_X1 U788 ( .A1(G900), .A2(n1102), .ZN(n1097) );
XNOR2_X1 U789 ( .A(G953), .B(KEYINPUT21), .ZN(n1102) );
NAND3_X1 U790 ( .A1(n1103), .A2(n1069), .A3(KEYINPUT59), .ZN(n1095) );
NAND2_X1 U791 ( .A1(G953), .A2(n1104), .ZN(n1093) );
NAND2_X1 U792 ( .A1(G900), .A2(G227), .ZN(n1104) );
XOR2_X1 U793 ( .A(n1105), .B(n1106), .Z(G69) );
NOR2_X1 U794 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XOR2_X1 U795 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U796 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U797 ( .A1(G953), .A2(n1113), .ZN(n1109) );
NOR3_X1 U798 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1113) );
NAND3_X1 U799 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1114) );
AND2_X1 U800 ( .A1(n1112), .A2(n1111), .ZN(n1107) );
NAND2_X1 U801 ( .A1(n1120), .A2(n1121), .ZN(n1111) );
NAND2_X1 U802 ( .A1(G953), .A2(n1122), .ZN(n1121) );
XOR2_X1 U803 ( .A(n1123), .B(n1124), .Z(n1120) );
NAND2_X1 U804 ( .A1(KEYINPUT33), .A2(n1125), .ZN(n1123) );
INV_X1 U805 ( .A(KEYINPUT7), .ZN(n1112) );
NAND3_X1 U806 ( .A1(G953), .A2(n1126), .A3(KEYINPUT46), .ZN(n1105) );
NAND2_X1 U807 ( .A1(G224), .A2(G898), .ZN(n1126) );
NOR2_X1 U808 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XNOR2_X1 U809 ( .A(n1129), .B(n1130), .ZN(n1128) );
NOR2_X1 U810 ( .A1(KEYINPUT25), .A2(n1131), .ZN(n1130) );
NOR2_X1 U811 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XNOR2_X1 U812 ( .A(G217), .B(KEYINPUT44), .ZN(n1132) );
NOR2_X1 U813 ( .A1(n1127), .A2(n1134), .ZN(G63) );
XOR2_X1 U814 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U815 ( .A1(KEYINPUT55), .A2(n1137), .ZN(n1136) );
AND2_X1 U816 ( .A1(G478), .A2(n1138), .ZN(n1135) );
NOR2_X1 U817 ( .A1(n1127), .A2(n1139), .ZN(G60) );
XOR2_X1 U818 ( .A(n1140), .B(n1141), .Z(n1139) );
AND2_X1 U819 ( .A1(G475), .A2(n1138), .ZN(n1140) );
XNOR2_X1 U820 ( .A(G104), .B(n1142), .ZN(G6) );
NOR2_X1 U821 ( .A1(n1127), .A2(n1143), .ZN(G57) );
XOR2_X1 U822 ( .A(n1144), .B(n1145), .Z(n1143) );
XNOR2_X1 U823 ( .A(n1146), .B(n1147), .ZN(n1145) );
XOR2_X1 U824 ( .A(n1148), .B(n1149), .Z(n1144) );
NAND2_X1 U825 ( .A1(KEYINPUT23), .A2(n1150), .ZN(n1149) );
NAND3_X1 U826 ( .A1(n1151), .A2(n1152), .A3(G472), .ZN(n1148) );
NAND2_X1 U827 ( .A1(KEYINPUT36), .A2(n1133), .ZN(n1152) );
NAND2_X1 U828 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
INV_X1 U829 ( .A(KEYINPUT36), .ZN(n1154) );
NOR2_X1 U830 ( .A1(n1127), .A2(n1155), .ZN(G54) );
XOR2_X1 U831 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U832 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U833 ( .A(n1160), .B(n1161), .Z(n1159) );
NAND2_X1 U834 ( .A1(n1138), .A2(G469), .ZN(n1161) );
XOR2_X1 U835 ( .A(n1162), .B(n1163), .Z(n1158) );
NOR2_X1 U836 ( .A1(G110), .A2(KEYINPUT24), .ZN(n1163) );
XOR2_X1 U837 ( .A(n1164), .B(n1165), .Z(n1156) );
XOR2_X1 U838 ( .A(KEYINPUT15), .B(G140), .Z(n1165) );
XNOR2_X1 U839 ( .A(n1166), .B(n1167), .ZN(n1164) );
NAND2_X1 U840 ( .A1(n1168), .A2(n1169), .ZN(n1166) );
NAND2_X1 U841 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NAND2_X1 U842 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NAND2_X1 U843 ( .A1(KEYINPUT14), .A2(n1174), .ZN(n1173) );
INV_X1 U844 ( .A(n1175), .ZN(n1174) );
NAND2_X1 U845 ( .A1(n1175), .A2(n1176), .ZN(n1168) );
NAND2_X1 U846 ( .A1(KEYINPUT14), .A2(n1177), .ZN(n1176) );
NAND2_X1 U847 ( .A1(n1178), .A2(n1172), .ZN(n1177) );
INV_X1 U848 ( .A(KEYINPUT39), .ZN(n1172) );
XNOR2_X1 U849 ( .A(n1179), .B(n1180), .ZN(n1175) );
NOR2_X1 U850 ( .A1(n1127), .A2(n1181), .ZN(G51) );
XOR2_X1 U851 ( .A(n1182), .B(n1183), .Z(n1181) );
NAND3_X1 U852 ( .A1(n1184), .A2(n1185), .A3(n1087), .ZN(n1183) );
INV_X1 U853 ( .A(n1186), .ZN(n1087) );
NAND2_X1 U854 ( .A1(KEYINPUT32), .A2(n1133), .ZN(n1185) );
INV_X1 U855 ( .A(n1138), .ZN(n1133) );
NOR2_X1 U856 ( .A1(n1187), .A2(n1067), .ZN(n1138) );
NAND2_X1 U857 ( .A1(n1153), .A2(n1188), .ZN(n1184) );
INV_X1 U858 ( .A(KEYINPUT32), .ZN(n1188) );
NAND2_X1 U859 ( .A1(n1067), .A2(G902), .ZN(n1153) );
NOR3_X1 U860 ( .A1(n1116), .A2(n1189), .A3(n1103), .ZN(n1067) );
NAND4_X1 U861 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1103) );
NOR4_X1 U862 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
NOR3_X1 U863 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1192) );
NOR2_X1 U864 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
INV_X1 U865 ( .A(KEYINPUT63), .ZN(n1201) );
NOR2_X1 U866 ( .A1(KEYINPUT63), .A2(n1203), .ZN(n1199) );
NAND4_X1 U867 ( .A1(n1204), .A2(n1030), .A3(n1205), .A4(n1064), .ZN(n1203) );
XNOR2_X1 U868 ( .A(KEYINPUT38), .B(n1206), .ZN(n1189) );
AND4_X1 U869 ( .A1(n1118), .A2(n1117), .A3(n1119), .A4(n1207), .ZN(n1206) );
XOR2_X1 U870 ( .A(n1115), .B(KEYINPUT0), .Z(n1207) );
NAND4_X1 U871 ( .A1(n1208), .A2(n1209), .A3(n1142), .A4(n1210), .ZN(n1116) );
NAND3_X1 U872 ( .A1(n1211), .A2(n1028), .A3(n1212), .ZN(n1142) );
NAND4_X1 U873 ( .A1(n1027), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1209) );
NAND2_X1 U874 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND3_X1 U875 ( .A1(n1053), .A2(n1218), .A3(n1074), .ZN(n1216) );
INV_X1 U876 ( .A(KEYINPUT13), .ZN(n1218) );
NAND2_X1 U877 ( .A1(n1033), .A2(n1219), .ZN(n1214) );
NAND2_X1 U878 ( .A1(n1028), .A2(n1030), .ZN(n1219) );
NAND2_X1 U879 ( .A1(KEYINPUT13), .A2(n1220), .ZN(n1208) );
NAND3_X1 U880 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1182) );
OR2_X1 U881 ( .A1(n1224), .A2(KEYINPUT6), .ZN(n1223) );
NAND3_X1 U882 ( .A1(KEYINPUT6), .A2(n1224), .A3(n1225), .ZN(n1222) );
NAND2_X1 U883 ( .A1(n1226), .A2(n1227), .ZN(n1221) );
NAND2_X1 U884 ( .A1(KEYINPUT6), .A2(n1228), .ZN(n1227) );
XOR2_X1 U885 ( .A(KEYINPUT48), .B(n1224), .Z(n1228) );
XNOR2_X1 U886 ( .A(n1229), .B(n1230), .ZN(n1224) );
NOR2_X1 U887 ( .A1(KEYINPUT52), .A2(n1231), .ZN(n1230) );
NOR2_X1 U888 ( .A1(n1069), .A2(G952), .ZN(n1127) );
NAND2_X1 U889 ( .A1(n1232), .A2(n1233), .ZN(G48) );
NAND2_X1 U890 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U891 ( .A(KEYINPUT56), .B(G146), .Z(n1235) );
XOR2_X1 U892 ( .A(KEYINPUT51), .B(n1236), .Z(n1232) );
NOR2_X1 U893 ( .A1(n1234), .A2(n1237), .ZN(n1236) );
XOR2_X1 U894 ( .A(KEYINPUT47), .B(G146), .Z(n1237) );
INV_X1 U895 ( .A(n1190), .ZN(n1234) );
NAND3_X1 U896 ( .A1(n1211), .A2(n1205), .A3(n1238), .ZN(n1190) );
XNOR2_X1 U897 ( .A(G143), .B(n1239), .ZN(G45) );
NAND2_X1 U898 ( .A1(KEYINPUT37), .A2(n1240), .ZN(n1239) );
INV_X1 U899 ( .A(n1191), .ZN(n1240) );
NAND4_X1 U900 ( .A1(n1238), .A2(n1074), .A3(n1084), .A4(n1241), .ZN(n1191) );
XOR2_X1 U901 ( .A(G140), .B(n1197), .Z(G42) );
AND3_X1 U902 ( .A1(n1211), .A2(n1242), .A3(n1243), .ZN(n1197) );
XNOR2_X1 U903 ( .A(G137), .B(n1244), .ZN(G39) );
NOR2_X1 U904 ( .A1(n1196), .A2(KEYINPUT26), .ZN(n1244) );
AND3_X1 U905 ( .A1(n1205), .A2(n1053), .A3(n1243), .ZN(n1196) );
NAND3_X1 U906 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(G36) );
OR2_X1 U907 ( .A1(n1167), .A2(KEYINPUT31), .ZN(n1247) );
NAND3_X1 U908 ( .A1(KEYINPUT31), .A2(n1167), .A3(n1198), .ZN(n1246) );
INV_X1 U909 ( .A(n1248), .ZN(n1198) );
NAND2_X1 U910 ( .A1(n1249), .A2(n1248), .ZN(n1245) );
NAND3_X1 U911 ( .A1(n1030), .A2(n1074), .A3(n1243), .ZN(n1248) );
NAND2_X1 U912 ( .A1(KEYINPUT31), .A2(n1250), .ZN(n1249) );
XNOR2_X1 U913 ( .A(KEYINPUT9), .B(n1167), .ZN(n1250) );
XOR2_X1 U914 ( .A(G131), .B(n1195), .Z(G33) );
AND3_X1 U915 ( .A1(n1211), .A2(n1074), .A3(n1243), .ZN(n1195) );
AND4_X1 U916 ( .A1(n1043), .A2(n1027), .A3(n1251), .A4(n1047), .ZN(n1243) );
XNOR2_X1 U917 ( .A(G128), .B(n1202), .ZN(G30) );
NAND3_X1 U918 ( .A1(n1030), .A2(n1205), .A3(n1238), .ZN(n1202) );
AND2_X1 U919 ( .A1(n1204), .A2(n1027), .ZN(n1238) );
XOR2_X1 U920 ( .A(G101), .B(n1220), .Z(G3) );
AND3_X1 U921 ( .A1(n1074), .A2(n1053), .A3(n1212), .ZN(n1220) );
XOR2_X1 U922 ( .A(G125), .B(n1194), .Z(G27) );
AND4_X1 U923 ( .A1(n1211), .A2(n1204), .A3(n1242), .A4(n1056), .ZN(n1194) );
INV_X1 U924 ( .A(n1065), .ZN(n1056) );
AND2_X1 U925 ( .A1(n1033), .A2(n1251), .ZN(n1204) );
NAND2_X1 U926 ( .A1(n1060), .A2(n1252), .ZN(n1251) );
NAND4_X1 U927 ( .A1(G953), .A2(G902), .A3(n1253), .A4(n1254), .ZN(n1252) );
INV_X1 U928 ( .A(G900), .ZN(n1254) );
XNOR2_X1 U929 ( .A(G122), .B(n1119), .ZN(G24) );
NAND4_X1 U930 ( .A1(n1255), .A2(n1028), .A3(n1084), .A4(n1241), .ZN(n1119) );
INV_X1 U931 ( .A(n1256), .ZN(n1241) );
XNOR2_X1 U932 ( .A(G119), .B(n1117), .ZN(G21) );
NAND3_X1 U933 ( .A1(n1205), .A2(n1053), .A3(n1255), .ZN(n1117) );
NAND2_X1 U934 ( .A1(n1257), .A2(n1258), .ZN(n1205) );
NAND2_X1 U935 ( .A1(n1242), .A2(n1259), .ZN(n1258) );
NAND3_X1 U936 ( .A1(n1086), .A2(n1260), .A3(KEYINPUT8), .ZN(n1257) );
XNOR2_X1 U937 ( .A(G116), .B(n1118), .ZN(G18) );
NAND3_X1 U938 ( .A1(n1030), .A2(n1074), .A3(n1255), .ZN(n1118) );
AND2_X1 U939 ( .A1(n1261), .A2(n1262), .ZN(n1030) );
XNOR2_X1 U940 ( .A(n1256), .B(KEYINPUT62), .ZN(n1262) );
XNOR2_X1 U941 ( .A(n1084), .B(KEYINPUT29), .ZN(n1261) );
XOR2_X1 U942 ( .A(G113), .B(n1115), .Z(G15) );
AND3_X1 U943 ( .A1(n1211), .A2(n1074), .A3(n1255), .ZN(n1115) );
NOR3_X1 U944 ( .A1(n1217), .A2(n1031), .A3(n1065), .ZN(n1255) );
NAND2_X1 U945 ( .A1(n1054), .A2(n1263), .ZN(n1065) );
NAND2_X1 U946 ( .A1(n1264), .A2(n1265), .ZN(n1074) );
NAND2_X1 U947 ( .A1(n1028), .A2(n1259), .ZN(n1265) );
NOR2_X1 U948 ( .A1(n1260), .A2(n1086), .ZN(n1028) );
OR3_X1 U949 ( .A1(n1260), .A2(n1266), .A3(n1259), .ZN(n1264) );
INV_X1 U950 ( .A(KEYINPUT8), .ZN(n1259) );
NAND2_X1 U951 ( .A1(n1267), .A2(n1268), .ZN(G12) );
NAND3_X1 U952 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1268) );
NAND2_X1 U953 ( .A1(G110), .A2(n1272), .ZN(n1267) );
NAND2_X1 U954 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
OR2_X1 U955 ( .A1(n1275), .A2(n1210), .ZN(n1274) );
NAND2_X1 U956 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
NAND2_X1 U957 ( .A1(n1269), .A2(n1270), .ZN(n1276) );
INV_X1 U958 ( .A(KEYINPUT3), .ZN(n1270) );
INV_X1 U959 ( .A(n1210), .ZN(n1269) );
NAND3_X1 U960 ( .A1(n1242), .A2(n1053), .A3(n1212), .ZN(n1210) );
NOR3_X1 U961 ( .A1(n1217), .A2(n1031), .A3(n1064), .ZN(n1212) );
INV_X1 U962 ( .A(n1027), .ZN(n1064) );
NOR2_X1 U963 ( .A1(n1054), .A2(n1055), .ZN(n1027) );
INV_X1 U964 ( .A(n1263), .ZN(n1055) );
NAND2_X1 U965 ( .A1(G221), .A2(n1277), .ZN(n1263) );
NAND2_X1 U966 ( .A1(G234), .A2(n1187), .ZN(n1277) );
NAND3_X1 U967 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1054) );
OR2_X1 U968 ( .A1(n1090), .A2(KEYINPUT16), .ZN(n1280) );
OR3_X1 U969 ( .A1(n1281), .A2(n1282), .A3(G469), .ZN(n1279) );
INV_X1 U970 ( .A(KEYINPUT16), .ZN(n1281) );
NAND2_X1 U971 ( .A1(G469), .A2(n1282), .ZN(n1278) );
NAND2_X1 U972 ( .A1(KEYINPUT28), .A2(n1090), .ZN(n1282) );
NAND2_X1 U973 ( .A1(n1283), .A2(n1187), .ZN(n1090) );
XOR2_X1 U974 ( .A(n1284), .B(n1285), .Z(n1283) );
XOR2_X1 U975 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U976 ( .A(KEYINPUT35), .B(KEYINPUT20), .Z(n1287) );
NOR2_X1 U977 ( .A1(n1288), .A2(n1289), .ZN(n1286) );
XOR2_X1 U978 ( .A(KEYINPUT1), .B(n1290), .Z(n1289) );
NOR2_X1 U979 ( .A1(n1291), .A2(n1160), .ZN(n1290) );
AND2_X1 U980 ( .A1(n1160), .A2(n1291), .ZN(n1288) );
XNOR2_X1 U981 ( .A(G140), .B(n1271), .ZN(n1291) );
INV_X1 U982 ( .A(G110), .ZN(n1271) );
NAND2_X1 U983 ( .A1(G227), .A2(n1069), .ZN(n1160) );
XNOR2_X1 U984 ( .A(n1099), .B(n1178), .ZN(n1284) );
INV_X1 U985 ( .A(n1170), .ZN(n1178) );
XNOR2_X1 U986 ( .A(n1292), .B(n1293), .ZN(n1170) );
XNOR2_X1 U987 ( .A(G101), .B(KEYINPUT22), .ZN(n1292) );
XOR2_X1 U988 ( .A(n1179), .B(n1294), .Z(n1099) );
NAND2_X1 U989 ( .A1(KEYINPUT50), .A2(n1295), .ZN(n1179) );
INV_X1 U990 ( .A(n1213), .ZN(n1031) );
NAND2_X1 U991 ( .A1(n1060), .A2(n1296), .ZN(n1213) );
NAND4_X1 U992 ( .A1(G953), .A2(G902), .A3(n1122), .A4(n1253), .ZN(n1296) );
XOR2_X1 U993 ( .A(KEYINPUT41), .B(G898), .Z(n1122) );
NAND3_X1 U994 ( .A1(n1253), .A2(n1069), .A3(G952), .ZN(n1060) );
NAND2_X1 U995 ( .A1(G237), .A2(G234), .ZN(n1253) );
INV_X1 U996 ( .A(n1033), .ZN(n1217) );
NOR2_X1 U997 ( .A1(n1043), .A2(n1297), .ZN(n1033) );
INV_X1 U998 ( .A(n1047), .ZN(n1297) );
NAND2_X1 U999 ( .A1(G214), .A2(n1298), .ZN(n1047) );
XOR2_X1 U1000 ( .A(n1089), .B(n1186), .Z(n1043) );
NAND2_X1 U1001 ( .A1(G210), .A2(n1298), .ZN(n1186) );
NAND2_X1 U1002 ( .A1(n1299), .A2(n1187), .ZN(n1298) );
INV_X1 U1003 ( .A(G237), .ZN(n1299) );
AND3_X1 U1004 ( .A1(n1300), .A2(n1187), .A3(n1301), .ZN(n1089) );
XOR2_X1 U1005 ( .A(n1302), .B(KEYINPUT5), .Z(n1301) );
NAND2_X1 U1006 ( .A1(n1225), .A2(n1303), .ZN(n1302) );
XNOR2_X1 U1007 ( .A(n1304), .B(n1305), .ZN(n1303) );
INV_X1 U1008 ( .A(n1226), .ZN(n1225) );
NAND2_X1 U1009 ( .A1(n1306), .A2(n1226), .ZN(n1300) );
XOR2_X1 U1010 ( .A(n1124), .B(n1125), .Z(n1226) );
XOR2_X1 U1011 ( .A(n1307), .B(n1308), .Z(n1124) );
XOR2_X1 U1012 ( .A(n1309), .B(n1293), .Z(n1308) );
XOR2_X1 U1013 ( .A(G104), .B(G107), .Z(n1293) );
NOR2_X1 U1014 ( .A1(G122), .A2(KEYINPUT43), .ZN(n1309) );
XNOR2_X1 U1015 ( .A(G110), .B(n1310), .ZN(n1307) );
NOR2_X1 U1016 ( .A1(G101), .A2(KEYINPUT17), .ZN(n1310) );
XNOR2_X1 U1017 ( .A(n1304), .B(n1229), .ZN(n1306) );
INV_X1 U1018 ( .A(n1305), .ZN(n1229) );
XOR2_X1 U1019 ( .A(G125), .B(n1311), .Z(n1305) );
AND2_X1 U1020 ( .A1(n1069), .A2(G224), .ZN(n1311) );
INV_X1 U1021 ( .A(G953), .ZN(n1069) );
NAND2_X1 U1022 ( .A1(KEYINPUT2), .A2(n1231), .ZN(n1304) );
XNOR2_X1 U1023 ( .A(n1180), .B(n1295), .ZN(n1231) );
NAND2_X1 U1024 ( .A1(n1312), .A2(n1313), .ZN(n1053) );
OR2_X1 U1025 ( .A1(n1066), .A2(KEYINPUT62), .ZN(n1313) );
INV_X1 U1026 ( .A(n1211), .ZN(n1066) );
NOR2_X1 U1027 ( .A1(n1084), .A2(n1256), .ZN(n1211) );
NAND3_X1 U1028 ( .A1(n1256), .A2(n1314), .A3(KEYINPUT62), .ZN(n1312) );
INV_X1 U1029 ( .A(n1084), .ZN(n1314) );
XNOR2_X1 U1030 ( .A(n1315), .B(G478), .ZN(n1084) );
NAND2_X1 U1031 ( .A1(n1316), .A2(n1137), .ZN(n1315) );
XNOR2_X1 U1032 ( .A(n1317), .B(n1318), .ZN(n1137) );
XOR2_X1 U1033 ( .A(G116), .B(n1319), .Z(n1318) );
XNOR2_X1 U1034 ( .A(n1320), .B(G122), .ZN(n1319) );
INV_X1 U1035 ( .A(G143), .ZN(n1320) );
XOR2_X1 U1036 ( .A(n1321), .B(n1322), .Z(n1317) );
XNOR2_X1 U1037 ( .A(n1323), .B(n1324), .ZN(n1321) );
INV_X1 U1038 ( .A(G107), .ZN(n1324) );
NAND2_X1 U1039 ( .A1(G217), .A2(n1325), .ZN(n1323) );
XNOR2_X1 U1040 ( .A(KEYINPUT58), .B(n1187), .ZN(n1316) );
NOR2_X1 U1041 ( .A1(n1092), .A2(n1082), .ZN(n1256) );
NOR3_X1 U1042 ( .A1(G475), .A2(G902), .A3(n1141), .ZN(n1082) );
AND2_X1 U1043 ( .A1(G475), .A2(n1326), .ZN(n1092) );
OR2_X1 U1044 ( .A1(n1141), .A2(G902), .ZN(n1326) );
XNOR2_X1 U1045 ( .A(n1327), .B(KEYINPUT42), .ZN(n1141) );
XOR2_X1 U1046 ( .A(n1328), .B(n1329), .Z(n1327) );
XOR2_X1 U1047 ( .A(n1330), .B(n1331), .Z(n1329) );
XOR2_X1 U1048 ( .A(n1332), .B(G113), .Z(n1331) );
NAND2_X1 U1049 ( .A1(G214), .A2(n1333), .ZN(n1332) );
XNOR2_X1 U1050 ( .A(G131), .B(KEYINPUT10), .ZN(n1330) );
XOR2_X1 U1051 ( .A(n1334), .B(n1335), .Z(n1328) );
XNOR2_X1 U1052 ( .A(n1295), .B(n1101), .ZN(n1335) );
XNOR2_X1 U1053 ( .A(n1336), .B(n1337), .ZN(n1334) );
NOR2_X1 U1054 ( .A1(G122), .A2(KEYINPUT61), .ZN(n1337) );
NOR2_X1 U1055 ( .A1(G104), .A2(KEYINPUT60), .ZN(n1336) );
INV_X1 U1056 ( .A(n1048), .ZN(n1242) );
NAND2_X1 U1057 ( .A1(n1266), .A2(n1260), .ZN(n1048) );
NAND2_X1 U1058 ( .A1(n1338), .A2(n1083), .ZN(n1260) );
NAND2_X1 U1059 ( .A1(G217), .A2(n1339), .ZN(n1083) );
NAND2_X1 U1060 ( .A1(n1187), .A2(n1340), .ZN(n1339) );
NAND2_X1 U1061 ( .A1(n1129), .A2(n1341), .ZN(n1340) );
XOR2_X1 U1062 ( .A(KEYINPUT11), .B(n1081), .Z(n1338) );
AND3_X1 U1063 ( .A1(n1342), .A2(n1187), .A3(n1343), .ZN(n1081) );
INV_X1 U1064 ( .A(n1129), .ZN(n1343) );
XNOR2_X1 U1065 ( .A(n1344), .B(n1345), .ZN(n1129) );
XNOR2_X1 U1066 ( .A(n1180), .B(n1346), .ZN(n1345) );
XNOR2_X1 U1067 ( .A(n1347), .B(n1348), .ZN(n1346) );
NOR2_X1 U1068 ( .A1(KEYINPUT12), .A2(n1101), .ZN(n1348) );
XNOR2_X1 U1069 ( .A(G125), .B(G140), .ZN(n1101) );
NOR2_X1 U1070 ( .A1(KEYINPUT19), .A2(n1349), .ZN(n1347) );
XNOR2_X1 U1071 ( .A(n1350), .B(n1351), .ZN(n1349) );
INV_X1 U1072 ( .A(G137), .ZN(n1351) );
NAND2_X1 U1073 ( .A1(n1325), .A2(G221), .ZN(n1350) );
NOR2_X1 U1074 ( .A1(n1341), .A2(G953), .ZN(n1325) );
XOR2_X1 U1075 ( .A(n1352), .B(n1353), .Z(n1344) );
XOR2_X1 U1076 ( .A(KEYINPUT10), .B(G146), .Z(n1353) );
XNOR2_X1 U1077 ( .A(G119), .B(G110), .ZN(n1352) );
NAND2_X1 U1078 ( .A1(G217), .A2(n1341), .ZN(n1342) );
INV_X1 U1079 ( .A(G234), .ZN(n1341) );
INV_X1 U1080 ( .A(n1086), .ZN(n1266) );
XNOR2_X1 U1081 ( .A(n1354), .B(G472), .ZN(n1086) );
NAND2_X1 U1082 ( .A1(n1355), .A2(n1187), .ZN(n1354) );
INV_X1 U1083 ( .A(G902), .ZN(n1187) );
XOR2_X1 U1084 ( .A(n1356), .B(n1357), .Z(n1355) );
XOR2_X1 U1085 ( .A(KEYINPUT27), .B(n1150), .Z(n1357) );
XNOR2_X1 U1086 ( .A(n1125), .B(KEYINPUT45), .ZN(n1150) );
XNOR2_X1 U1087 ( .A(G113), .B(n1358), .ZN(n1125) );
XNOR2_X1 U1088 ( .A(n1359), .B(G116), .ZN(n1358) );
INV_X1 U1089 ( .A(G119), .ZN(n1359) );
XNOR2_X1 U1090 ( .A(n1147), .B(n1360), .ZN(n1356) );
INV_X1 U1091 ( .A(n1146), .ZN(n1360) );
XNOR2_X1 U1092 ( .A(n1361), .B(G101), .ZN(n1146) );
NAND2_X1 U1093 ( .A1(G210), .A2(n1333), .ZN(n1361) );
NOR2_X1 U1094 ( .A1(G953), .A2(G237), .ZN(n1333) );
XNOR2_X1 U1095 ( .A(n1295), .B(n1294), .ZN(n1147) );
XNOR2_X1 U1096 ( .A(n1162), .B(n1322), .ZN(n1294) );
XNOR2_X1 U1097 ( .A(n1167), .B(n1180), .ZN(n1322) );
XOR2_X1 U1098 ( .A(G128), .B(KEYINPUT4), .Z(n1180) );
INV_X1 U1099 ( .A(G134), .ZN(n1167) );
XNOR2_X1 U1100 ( .A(G131), .B(G137), .ZN(n1162) );
XOR2_X1 U1101 ( .A(G143), .B(G146), .Z(n1295) );
XNOR2_X1 U1102 ( .A(KEYINPUT40), .B(KEYINPUT18), .ZN(n1275) );
endmodule


