//Key = 0100010111001001100011000000101110101000010010001010100100111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339;

XOR2_X1 U734 ( .A(n1016), .B(G107), .Z(G9) );
NAND2_X1 U735 ( .A1(KEYINPUT28), .A2(n1017), .ZN(n1016) );
NOR2_X1 U736 ( .A1(n1018), .A2(n1019), .ZN(G75) );
NOR4_X1 U737 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1019) );
INV_X1 U738 ( .A(G952), .ZN(n1022) );
NAND3_X1 U739 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1020) );
NAND2_X1 U740 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U741 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND3_X1 U742 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
NAND2_X1 U743 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NAND2_X1 U744 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U745 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U747 ( .A1(n1042), .A2(n1043), .ZN(n1034) );
NAND2_X1 U748 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U749 ( .A1(n1036), .A2(n1046), .A3(n1042), .ZN(n1029) );
NAND2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U751 ( .A1(n1031), .A2(n1049), .ZN(n1048) );
NAND2_X1 U752 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U753 ( .A1(n1033), .A2(n1052), .ZN(n1047) );
NAND2_X1 U754 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U755 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
INV_X1 U756 ( .A(n1057), .ZN(n1055) );
INV_X1 U757 ( .A(n1058), .ZN(n1027) );
NOR3_X1 U758 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1018) );
NOR2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
INV_X1 U760 ( .A(KEYINPUT21), .ZN(n1063) );
NOR2_X1 U761 ( .A1(G953), .A2(G952), .ZN(n1062) );
NOR2_X1 U762 ( .A1(KEYINPUT21), .A2(n1064), .ZN(n1060) );
INV_X1 U763 ( .A(n1024), .ZN(n1059) );
NAND4_X1 U764 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1024) );
NOR3_X1 U765 ( .A1(n1069), .A2(n1040), .A3(n1070), .ZN(n1068) );
NOR2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U767 ( .A1(n1073), .A2(n1074), .A3(n1057), .ZN(n1069) );
NOR3_X1 U768 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1067) );
XOR2_X1 U769 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U770 ( .A1(G472), .A2(KEYINPUT6), .ZN(n1079) );
NOR2_X1 U771 ( .A1(n1080), .A2(n1081), .ZN(n1076) );
XNOR2_X1 U772 ( .A(n1082), .B(n1083), .ZN(n1075) );
NOR2_X1 U773 ( .A1(n1084), .A2(KEYINPUT18), .ZN(n1083) );
XNOR2_X1 U774 ( .A(n1085), .B(KEYINPUT26), .ZN(n1065) );
XOR2_X1 U775 ( .A(n1086), .B(n1087), .Z(G72) );
XOR2_X1 U776 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
AND2_X1 U778 ( .A1(G227), .A2(G900), .ZN(n1090) );
NAND2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1088) );
NAND2_X1 U780 ( .A1(G953), .A2(n1094), .ZN(n1093) );
XOR2_X1 U781 ( .A(n1095), .B(n1096), .Z(n1092) );
XOR2_X1 U782 ( .A(n1097), .B(n1098), .Z(n1096) );
XNOR2_X1 U783 ( .A(n1099), .B(n1100), .ZN(n1098) );
XNOR2_X1 U784 ( .A(KEYINPUT15), .B(n1101), .ZN(n1095) );
XNOR2_X1 U785 ( .A(KEYINPUT51), .B(KEYINPUT16), .ZN(n1101) );
NAND2_X1 U786 ( .A1(n1025), .A2(n1021), .ZN(n1086) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(G69) );
NOR2_X1 U788 ( .A1(n1104), .A2(n1091), .ZN(n1103) );
XNOR2_X1 U789 ( .A(G953), .B(KEYINPUT22), .ZN(n1091) );
AND2_X1 U790 ( .A1(G224), .A2(G898), .ZN(n1104) );
NAND2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1102) );
NAND2_X1 U792 ( .A1(n1107), .A2(n1025), .ZN(n1106) );
XOR2_X1 U793 ( .A(n1023), .B(n1108), .Z(n1107) );
NAND3_X1 U794 ( .A1(G898), .A2(n1108), .A3(G953), .ZN(n1105) );
NAND2_X1 U795 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
OR2_X1 U796 ( .A1(n1111), .A2(KEYINPUT42), .ZN(n1110) );
NAND2_X1 U797 ( .A1(n1112), .A2(KEYINPUT42), .ZN(n1109) );
NOR2_X1 U798 ( .A1(n1064), .A2(n1113), .ZN(G66) );
XOR2_X1 U799 ( .A(n1114), .B(n1115), .Z(n1113) );
AND3_X1 U800 ( .A1(n1116), .A2(n1117), .A3(G217), .ZN(n1115) );
NAND2_X1 U801 ( .A1(KEYINPUT55), .A2(n1118), .ZN(n1114) );
NOR2_X1 U802 ( .A1(n1064), .A2(n1119), .ZN(G63) );
XNOR2_X1 U803 ( .A(n1120), .B(n1121), .ZN(n1119) );
NOR3_X1 U804 ( .A1(n1122), .A2(KEYINPUT53), .A3(n1123), .ZN(n1121) );
NOR2_X1 U805 ( .A1(n1064), .A2(n1124), .ZN(G60) );
XOR2_X1 U806 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND2_X1 U807 ( .A1(n1116), .A2(G475), .ZN(n1125) );
XNOR2_X1 U808 ( .A(G104), .B(n1127), .ZN(G6) );
NOR2_X1 U809 ( .A1(n1064), .A2(n1128), .ZN(G57) );
XOR2_X1 U810 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U811 ( .A(n1131), .B(n1132), .Z(n1129) );
NOR3_X1 U812 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
NOR3_X1 U813 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(n1134) );
INV_X1 U815 ( .A(n1141), .ZN(n1133) );
NAND2_X1 U816 ( .A1(n1116), .A2(G472), .ZN(n1131) );
NOR2_X1 U817 ( .A1(n1142), .A2(n1143), .ZN(G54) );
XOR2_X1 U818 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U819 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U820 ( .A1(n1148), .A2(KEYINPUT46), .ZN(n1147) );
AND2_X1 U821 ( .A1(G469), .A2(n1116), .ZN(n1148) );
INV_X1 U822 ( .A(n1122), .ZN(n1116) );
NOR2_X1 U823 ( .A1(n1149), .A2(n1150), .ZN(n1146) );
XOR2_X1 U824 ( .A(KEYINPUT61), .B(n1151), .Z(n1150) );
NOR2_X1 U825 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
AND2_X1 U826 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
XNOR2_X1 U827 ( .A(n1154), .B(KEYINPUT9), .ZN(n1153) );
XNOR2_X1 U828 ( .A(n1064), .B(KEYINPUT1), .ZN(n1142) );
NOR2_X1 U829 ( .A1(n1064), .A2(n1155), .ZN(G51) );
XOR2_X1 U830 ( .A(KEYINPUT27), .B(n1156), .Z(n1155) );
NOR2_X1 U831 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NOR2_X1 U832 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U833 ( .A(KEYINPUT10), .B(n1161), .Z(n1159) );
AND2_X1 U834 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NOR2_X1 U835 ( .A1(n1122), .A2(n1162), .ZN(n1161) );
NAND2_X1 U836 ( .A1(G902), .A2(n1163), .ZN(n1122) );
OR2_X1 U837 ( .A1(n1021), .A2(n1023), .ZN(n1163) );
NAND4_X1 U838 ( .A1(n1164), .A2(n1127), .A3(n1165), .A4(n1166), .ZN(n1023) );
AND4_X1 U839 ( .A1(n1017), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1166) );
NAND3_X1 U840 ( .A1(n1170), .A2(n1036), .A3(n1171), .ZN(n1017) );
NAND2_X1 U841 ( .A1(n1172), .A2(n1173), .ZN(n1165) );
XOR2_X1 U842 ( .A(n1174), .B(KEYINPUT58), .Z(n1172) );
NAND3_X1 U843 ( .A1(n1171), .A2(n1036), .A3(n1175), .ZN(n1127) );
NAND3_X1 U844 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1164) );
NAND2_X1 U845 ( .A1(n1179), .A2(n1050), .ZN(n1177) );
XNOR2_X1 U846 ( .A(n1170), .B(KEYINPUT13), .ZN(n1179) );
NAND2_X1 U847 ( .A1(n1180), .A2(n1181), .ZN(n1021) );
AND4_X1 U848 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181) );
NOR4_X1 U849 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1180) );
XOR2_X1 U850 ( .A(n1190), .B(n1191), .Z(n1160) );
XNOR2_X1 U851 ( .A(n1192), .B(n1193), .ZN(n1190) );
NAND2_X1 U852 ( .A1(KEYINPUT59), .A2(n1111), .ZN(n1192) );
INV_X1 U853 ( .A(n1194), .ZN(n1111) );
NOR2_X1 U854 ( .A1(n1025), .A2(G952), .ZN(n1064) );
XOR2_X1 U855 ( .A(G146), .B(n1189), .Z(G48) );
AND3_X1 U856 ( .A1(n1175), .A2(n1173), .A3(n1195), .ZN(n1189) );
XNOR2_X1 U857 ( .A(G143), .B(n1196), .ZN(G45) );
NAND2_X1 U858 ( .A1(KEYINPUT50), .A2(n1188), .ZN(n1196) );
AND3_X1 U859 ( .A1(n1197), .A2(n1173), .A3(n1198), .ZN(n1188) );
NOR3_X1 U860 ( .A1(n1066), .A2(n1199), .A3(n1200), .ZN(n1198) );
XOR2_X1 U861 ( .A(G140), .B(n1187), .Z(G42) );
AND3_X1 U862 ( .A1(n1201), .A2(n1175), .A3(n1202), .ZN(n1187) );
XOR2_X1 U863 ( .A(G137), .B(n1186), .Z(G39) );
AND3_X1 U864 ( .A1(n1031), .A2(n1195), .A3(n1033), .ZN(n1186) );
NAND2_X1 U865 ( .A1(n1203), .A2(n1204), .ZN(G36) );
NAND2_X1 U866 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NAND2_X1 U867 ( .A1(G134), .A2(n1207), .ZN(n1203) );
NAND2_X1 U868 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U869 ( .A1(KEYINPUT40), .A2(n1210), .ZN(n1209) );
INV_X1 U870 ( .A(n1185), .ZN(n1210) );
OR2_X1 U871 ( .A1(n1205), .A2(KEYINPUT40), .ZN(n1208) );
NOR2_X1 U872 ( .A1(KEYINPUT63), .A2(n1185), .ZN(n1205) );
NAND2_X1 U873 ( .A1(n1211), .A2(n1202), .ZN(n1185) );
XNOR2_X1 U874 ( .A(G131), .B(n1184), .ZN(G33) );
NAND3_X1 U875 ( .A1(n1175), .A2(n1176), .A3(n1202), .ZN(n1184) );
AND3_X1 U876 ( .A1(n1212), .A2(n1213), .A3(n1031), .ZN(n1202) );
AND2_X1 U877 ( .A1(n1056), .A2(n1057), .ZN(n1031) );
XNOR2_X1 U878 ( .A(n1214), .B(KEYINPUT44), .ZN(n1056) );
NAND2_X1 U879 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XNOR2_X1 U880 ( .A(G128), .B(n1183), .ZN(G30) );
NAND3_X1 U881 ( .A1(n1170), .A2(n1173), .A3(n1195), .ZN(n1183) );
AND4_X1 U882 ( .A1(n1212), .A2(n1217), .A3(n1218), .A4(n1213), .ZN(n1195) );
XNOR2_X1 U883 ( .A(n1219), .B(n1220), .ZN(G3) );
NOR3_X1 U884 ( .A1(n1053), .A2(KEYINPUT33), .A3(n1221), .ZN(n1220) );
XOR2_X1 U885 ( .A(n1174), .B(KEYINPUT17), .Z(n1221) );
NAND3_X1 U886 ( .A1(n1033), .A2(n1222), .A3(n1197), .ZN(n1174) );
NOR2_X1 U887 ( .A1(n1045), .A2(n1038), .ZN(n1197) );
XNOR2_X1 U888 ( .A(G125), .B(n1182), .ZN(G27) );
NAND3_X1 U889 ( .A1(n1201), .A2(n1042), .A3(n1223), .ZN(n1182) );
NOR3_X1 U890 ( .A1(n1050), .A2(n1199), .A3(n1053), .ZN(n1223) );
INV_X1 U891 ( .A(n1213), .ZN(n1199) );
NAND2_X1 U892 ( .A1(n1224), .A2(n1058), .ZN(n1213) );
NAND4_X1 U893 ( .A1(G953), .A2(G902), .A3(n1225), .A4(n1094), .ZN(n1224) );
INV_X1 U894 ( .A(G900), .ZN(n1094) );
INV_X1 U895 ( .A(n1175), .ZN(n1050) );
XNOR2_X1 U896 ( .A(n1169), .B(n1226), .ZN(G24) );
NOR2_X1 U897 ( .A1(KEYINPUT14), .A2(n1227), .ZN(n1226) );
INV_X1 U898 ( .A(G122), .ZN(n1227) );
NAND4_X1 U899 ( .A1(n1178), .A2(n1036), .A3(n1228), .A4(n1229), .ZN(n1169) );
NAND2_X1 U900 ( .A1(n1230), .A2(n1231), .ZN(n1036) );
OR2_X1 U901 ( .A1(n1045), .A2(KEYINPUT7), .ZN(n1231) );
NAND3_X1 U902 ( .A1(n1232), .A2(n1233), .A3(KEYINPUT7), .ZN(n1230) );
INV_X1 U903 ( .A(n1218), .ZN(n1232) );
XNOR2_X1 U904 ( .A(G119), .B(n1168), .ZN(G21) );
NAND4_X1 U905 ( .A1(n1178), .A2(n1033), .A3(n1217), .A4(n1218), .ZN(n1168) );
XNOR2_X1 U906 ( .A(n1233), .B(KEYINPUT39), .ZN(n1217) );
XNOR2_X1 U907 ( .A(G116), .B(n1234), .ZN(G18) );
NAND2_X1 U908 ( .A1(n1178), .A2(n1211), .ZN(n1234) );
NOR2_X1 U909 ( .A1(n1051), .A2(n1045), .ZN(n1211) );
INV_X1 U910 ( .A(n1170), .ZN(n1051) );
NOR2_X1 U911 ( .A1(n1229), .A2(n1066), .ZN(n1170) );
INV_X1 U912 ( .A(n1228), .ZN(n1066) );
AND3_X1 U913 ( .A1(n1173), .A2(n1222), .A3(n1042), .ZN(n1178) );
XNOR2_X1 U914 ( .A(G113), .B(n1235), .ZN(G15) );
NOR2_X1 U915 ( .A1(KEYINPUT0), .A2(n1236), .ZN(n1235) );
NOR4_X1 U916 ( .A1(n1237), .A2(n1045), .A3(n1238), .A4(n1239), .ZN(n1236) );
XNOR2_X1 U917 ( .A(n1173), .B(KEYINPUT2), .ZN(n1239) );
INV_X1 U918 ( .A(n1053), .ZN(n1173) );
INV_X1 U919 ( .A(n1176), .ZN(n1045) );
NOR2_X1 U920 ( .A1(n1218), .A2(n1233), .ZN(n1176) );
NAND2_X1 U921 ( .A1(n1042), .A2(n1175), .ZN(n1237) );
NOR2_X1 U922 ( .A1(n1228), .A2(n1200), .ZN(n1175) );
INV_X1 U923 ( .A(n1229), .ZN(n1200) );
NOR2_X1 U924 ( .A1(n1085), .A2(n1040), .ZN(n1042) );
XNOR2_X1 U925 ( .A(G110), .B(n1167), .ZN(G12) );
NAND3_X1 U926 ( .A1(n1201), .A2(n1171), .A3(n1033), .ZN(n1167) );
NOR2_X1 U927 ( .A1(n1228), .A2(n1229), .ZN(n1033) );
NAND3_X1 U928 ( .A1(n1240), .A2(n1241), .A3(n1074), .ZN(n1229) );
NAND2_X1 U929 ( .A1(n1071), .A2(n1072), .ZN(n1074) );
INV_X1 U930 ( .A(G475), .ZN(n1072) );
INV_X1 U931 ( .A(n1242), .ZN(n1071) );
OR2_X1 U932 ( .A1(G475), .A2(KEYINPUT48), .ZN(n1241) );
NAND3_X1 U933 ( .A1(G475), .A2(n1242), .A3(KEYINPUT48), .ZN(n1240) );
NAND2_X1 U934 ( .A1(n1126), .A2(n1243), .ZN(n1242) );
XNOR2_X1 U935 ( .A(n1244), .B(n1245), .ZN(n1126) );
XOR2_X1 U936 ( .A(n1246), .B(n1247), .Z(n1245) );
XNOR2_X1 U937 ( .A(G104), .B(n1248), .ZN(n1247) );
NOR2_X1 U938 ( .A1(KEYINPUT24), .A2(G113), .ZN(n1248) );
XNOR2_X1 U939 ( .A(G131), .B(G146), .ZN(n1246) );
XOR2_X1 U940 ( .A(n1249), .B(n1250), .Z(n1244) );
XNOR2_X1 U941 ( .A(n1100), .B(n1251), .ZN(n1250) );
XOR2_X1 U942 ( .A(n1252), .B(n1253), .Z(n1249) );
NOR2_X1 U943 ( .A1(G143), .A2(n1254), .ZN(n1253) );
XNOR2_X1 U944 ( .A(KEYINPUT4), .B(KEYINPUT30), .ZN(n1254) );
NAND2_X1 U945 ( .A1(n1255), .A2(G214), .ZN(n1252) );
XOR2_X1 U946 ( .A(n1256), .B(n1123), .Z(n1228) );
INV_X1 U947 ( .A(G478), .ZN(n1123) );
NAND2_X1 U948 ( .A1(n1257), .A2(n1120), .ZN(n1256) );
NAND2_X1 U949 ( .A1(n1258), .A2(n1259), .ZN(n1120) );
NAND2_X1 U950 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XOR2_X1 U951 ( .A(n1262), .B(KEYINPUT47), .Z(n1258) );
OR2_X1 U952 ( .A1(n1261), .A2(n1260), .ZN(n1262) );
XOR2_X1 U953 ( .A(n1263), .B(n1264), .Z(n1260) );
XOR2_X1 U954 ( .A(G107), .B(n1265), .Z(n1264) );
XOR2_X1 U955 ( .A(KEYINPUT60), .B(G116), .Z(n1265) );
XNOR2_X1 U956 ( .A(n1266), .B(n1267), .ZN(n1263) );
NOR2_X1 U957 ( .A1(KEYINPUT23), .A2(n1268), .ZN(n1267) );
XNOR2_X1 U958 ( .A(n1099), .B(n1269), .ZN(n1268) );
XOR2_X1 U959 ( .A(G143), .B(G128), .Z(n1269) );
NAND3_X1 U960 ( .A1(G234), .A2(n1025), .A3(G217), .ZN(n1261) );
XNOR2_X1 U961 ( .A(KEYINPUT20), .B(n1243), .ZN(n1257) );
NOR3_X1 U962 ( .A1(n1038), .A2(n1238), .A3(n1053), .ZN(n1171) );
NAND3_X1 U963 ( .A1(n1216), .A2(n1215), .A3(n1057), .ZN(n1053) );
NAND2_X1 U964 ( .A1(G214), .A2(n1270), .ZN(n1057) );
NAND2_X1 U965 ( .A1(n1271), .A2(n1272), .ZN(n1215) );
XNOR2_X1 U966 ( .A(KEYINPUT56), .B(n1273), .ZN(n1272) );
XNOR2_X1 U967 ( .A(KEYINPUT35), .B(n1162), .ZN(n1271) );
NAND2_X1 U968 ( .A1(n1274), .A2(n1275), .ZN(n1216) );
XNOR2_X1 U969 ( .A(n1084), .B(KEYINPUT56), .ZN(n1275) );
INV_X1 U970 ( .A(n1273), .ZN(n1084) );
NAND3_X1 U971 ( .A1(n1276), .A2(n1277), .A3(n1243), .ZN(n1273) );
OR2_X1 U972 ( .A1(n1278), .A2(n1194), .ZN(n1277) );
NAND2_X1 U973 ( .A1(n1278), .A2(n1279), .ZN(n1276) );
XNOR2_X1 U974 ( .A(n1194), .B(KEYINPUT34), .ZN(n1279) );
NOR2_X1 U975 ( .A1(n1112), .A2(n1280), .ZN(n1194) );
AND2_X1 U976 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NOR2_X1 U977 ( .A1(n1282), .A2(n1281), .ZN(n1112) );
XNOR2_X1 U978 ( .A(n1283), .B(n1251), .ZN(n1281) );
INV_X1 U979 ( .A(n1266), .ZN(n1251) );
XOR2_X1 U980 ( .A(G122), .B(KEYINPUT3), .Z(n1266) );
NAND2_X1 U981 ( .A1(KEYINPUT31), .A2(n1284), .ZN(n1283) );
XNOR2_X1 U982 ( .A(n1285), .B(n1286), .ZN(n1282) );
XOR2_X1 U983 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U984 ( .A(n1289), .B(n1290), .Z(n1285) );
XNOR2_X1 U985 ( .A(G119), .B(n1291), .ZN(n1290) );
NAND2_X1 U986 ( .A1(n1292), .A2(KEYINPUT36), .ZN(n1289) );
XNOR2_X1 U987 ( .A(G101), .B(KEYINPUT45), .ZN(n1292) );
XNOR2_X1 U988 ( .A(n1293), .B(n1191), .ZN(n1278) );
XNOR2_X1 U989 ( .A(n1294), .B(n1137), .ZN(n1191) );
NAND2_X1 U990 ( .A1(G224), .A2(n1025), .ZN(n1294) );
NAND2_X1 U991 ( .A1(KEYINPUT41), .A2(n1193), .ZN(n1293) );
XNOR2_X1 U992 ( .A(n1082), .B(KEYINPUT11), .ZN(n1274) );
INV_X1 U993 ( .A(n1162), .ZN(n1082) );
NAND2_X1 U994 ( .A1(G210), .A2(n1270), .ZN(n1162) );
NAND2_X1 U995 ( .A1(n1295), .A2(n1243), .ZN(n1270) );
XNOR2_X1 U996 ( .A(G237), .B(KEYINPUT54), .ZN(n1295) );
INV_X1 U997 ( .A(n1222), .ZN(n1238) );
NAND2_X1 U998 ( .A1(n1058), .A2(n1296), .ZN(n1222) );
NAND4_X1 U999 ( .A1(G953), .A2(G902), .A3(n1225), .A4(n1297), .ZN(n1296) );
INV_X1 U1000 ( .A(G898), .ZN(n1297) );
NAND3_X1 U1001 ( .A1(n1225), .A2(n1025), .A3(G952), .ZN(n1058) );
NAND2_X1 U1002 ( .A1(G234), .A2(G237), .ZN(n1225) );
INV_X1 U1003 ( .A(n1212), .ZN(n1038) );
NOR2_X1 U1004 ( .A1(n1041), .A2(n1040), .ZN(n1212) );
AND2_X1 U1005 ( .A1(G221), .A2(n1117), .ZN(n1040) );
INV_X1 U1006 ( .A(n1085), .ZN(n1041) );
XNOR2_X1 U1007 ( .A(n1298), .B(G469), .ZN(n1085) );
NAND2_X1 U1008 ( .A1(n1299), .A2(n1243), .ZN(n1298) );
XNOR2_X1 U1009 ( .A(n1144), .B(n1300), .ZN(n1299) );
XNOR2_X1 U1010 ( .A(n1154), .B(n1152), .ZN(n1300) );
XNOR2_X1 U1011 ( .A(G140), .B(n1284), .ZN(n1152) );
NAND2_X1 U1012 ( .A1(G227), .A2(n1025), .ZN(n1154) );
XNOR2_X1 U1013 ( .A(n1301), .B(n1302), .ZN(n1144) );
XOR2_X1 U1014 ( .A(KEYINPUT62), .B(KEYINPUT15), .Z(n1302) );
XOR2_X1 U1015 ( .A(n1303), .B(n1140), .Z(n1301) );
XNOR2_X1 U1016 ( .A(n1304), .B(n1097), .ZN(n1140) );
XNOR2_X1 U1017 ( .A(n1305), .B(n1137), .ZN(n1097) );
NAND2_X1 U1018 ( .A1(n1306), .A2(n1307), .ZN(n1303) );
OR2_X1 U1019 ( .A1(n1288), .A2(G101), .ZN(n1307) );
XOR2_X1 U1020 ( .A(n1308), .B(KEYINPUT19), .Z(n1306) );
NAND2_X1 U1021 ( .A1(G101), .A2(n1288), .ZN(n1308) );
XOR2_X1 U1022 ( .A(G104), .B(G107), .Z(n1288) );
INV_X1 U1023 ( .A(n1044), .ZN(n1201) );
NAND2_X1 U1024 ( .A1(n1309), .A2(n1218), .ZN(n1044) );
NAND3_X1 U1025 ( .A1(n1310), .A2(n1311), .A3(n1073), .ZN(n1218) );
NAND2_X1 U1026 ( .A1(n1080), .A2(n1081), .ZN(n1073) );
NAND2_X1 U1027 ( .A1(n1081), .A2(n1312), .ZN(n1311) );
OR3_X1 U1028 ( .A1(n1081), .A2(n1080), .A3(n1312), .ZN(n1310) );
INV_X1 U1029 ( .A(KEYINPUT12), .ZN(n1312) );
AND2_X1 U1030 ( .A1(n1118), .A2(n1243), .ZN(n1080) );
XOR2_X1 U1031 ( .A(n1313), .B(n1314), .Z(n1118) );
XOR2_X1 U1032 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1033 ( .A(G119), .B(n1284), .ZN(n1316) );
INV_X1 U1034 ( .A(G110), .ZN(n1284) );
XOR2_X1 U1035 ( .A(KEYINPUT5), .B(G137), .Z(n1315) );
XOR2_X1 U1036 ( .A(n1317), .B(n1100), .Z(n1313) );
XNOR2_X1 U1037 ( .A(G140), .B(n1193), .ZN(n1100) );
INV_X1 U1038 ( .A(G125), .ZN(n1193) );
XOR2_X1 U1039 ( .A(n1318), .B(n1319), .Z(n1317) );
NAND3_X1 U1040 ( .A1(G234), .A2(n1025), .A3(G221), .ZN(n1318) );
INV_X1 U1041 ( .A(G953), .ZN(n1025) );
NAND2_X1 U1042 ( .A1(n1320), .A2(n1117), .ZN(n1081) );
NAND2_X1 U1043 ( .A1(G234), .A2(n1321), .ZN(n1117) );
XNOR2_X1 U1044 ( .A(KEYINPUT8), .B(n1243), .ZN(n1321) );
XOR2_X1 U1045 ( .A(KEYINPUT43), .B(G217), .Z(n1320) );
XNOR2_X1 U1046 ( .A(KEYINPUT7), .B(n1233), .ZN(n1309) );
XOR2_X1 U1047 ( .A(n1078), .B(G472), .Z(n1233) );
NAND2_X1 U1048 ( .A1(n1322), .A2(n1243), .ZN(n1078) );
INV_X1 U1049 ( .A(G902), .ZN(n1243) );
XNOR2_X1 U1050 ( .A(n1130), .B(n1323), .ZN(n1322) );
XOR2_X1 U1051 ( .A(n1324), .B(KEYINPUT37), .Z(n1323) );
NAND2_X1 U1052 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NAND2_X1 U1053 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
NAND2_X1 U1054 ( .A1(n1138), .A2(n1329), .ZN(n1328) );
XNOR2_X1 U1055 ( .A(n1139), .B(n1330), .ZN(n1327) );
NAND2_X1 U1056 ( .A1(n1331), .A2(n1329), .ZN(n1325) );
INV_X1 U1057 ( .A(KEYINPUT25), .ZN(n1329) );
NAND2_X1 U1058 ( .A1(n1141), .A2(n1332), .ZN(n1331) );
NAND3_X1 U1059 ( .A1(n1330), .A2(n1138), .A3(n1136), .ZN(n1332) );
INV_X1 U1060 ( .A(n1139), .ZN(n1136) );
INV_X1 U1061 ( .A(n1137), .ZN(n1330) );
NAND3_X1 U1062 ( .A1(n1139), .A2(n1137), .A3(n1138), .ZN(n1141) );
XNOR2_X1 U1063 ( .A(n1305), .B(n1304), .ZN(n1138) );
OR2_X1 U1064 ( .A1(KEYINPUT29), .A2(n1099), .ZN(n1304) );
XOR2_X1 U1065 ( .A(n1206), .B(KEYINPUT32), .Z(n1099) );
INV_X1 U1066 ( .A(G134), .ZN(n1206) );
XNOR2_X1 U1067 ( .A(G131), .B(G137), .ZN(n1305) );
XOR2_X1 U1068 ( .A(G143), .B(n1319), .Z(n1137) );
XOR2_X1 U1069 ( .A(G128), .B(G146), .Z(n1319) );
XNOR2_X1 U1070 ( .A(n1333), .B(KEYINPUT52), .ZN(n1139) );
NAND2_X1 U1071 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NAND2_X1 U1072 ( .A1(n1336), .A2(n1291), .ZN(n1335) );
XOR2_X1 U1073 ( .A(n1337), .B(KEYINPUT49), .Z(n1334) );
OR2_X1 U1074 ( .A1(n1336), .A2(n1291), .ZN(n1337) );
INV_X1 U1075 ( .A(G113), .ZN(n1291) );
XOR2_X1 U1076 ( .A(n1287), .B(n1338), .Z(n1336) );
NOR2_X1 U1077 ( .A1(G119), .A2(KEYINPUT57), .ZN(n1338) );
XOR2_X1 U1078 ( .A(G116), .B(KEYINPUT38), .Z(n1287) );
XOR2_X1 U1079 ( .A(n1339), .B(n1219), .Z(n1130) );
INV_X1 U1080 ( .A(G101), .ZN(n1219) );
NAND2_X1 U1081 ( .A1(n1255), .A2(G210), .ZN(n1339) );
NOR2_X1 U1082 ( .A1(G953), .A2(G237), .ZN(n1255) );
endmodule


