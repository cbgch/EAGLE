//Key = 0100000110001101000101110011000011000011110110001111110000110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362;

XNOR2_X1 U748 ( .A(G107), .B(n1033), .ZN(G9) );
NOR2_X1 U749 ( .A1(n1034), .A2(n1035), .ZN(G75) );
NOR3_X1 U750 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NOR3_X1 U751 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1037) );
NOR3_X1 U752 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
NOR2_X1 U753 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U756 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U757 ( .A1(n1053), .A2(n1054), .ZN(n1047) );
NOR2_X1 U758 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U759 ( .A1(KEYINPUT56), .A2(n1057), .ZN(n1056) );
NOR2_X1 U760 ( .A1(n1058), .A2(n1059), .ZN(n1055) );
NOR3_X1 U761 ( .A1(n1050), .A2(n1060), .A3(n1054), .ZN(n1043) );
NOR2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(n1040) );
AND4_X1 U763 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(KEYINPUT56), .ZN(n1062) );
NAND3_X1 U764 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1036) );
NAND4_X1 U765 ( .A1(n1061), .A2(n1065), .A3(n1069), .A4(n1070), .ZN(n1068) );
NAND2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U767 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
XOR2_X1 U768 ( .A(n1054), .B(KEYINPUT12), .Z(n1075) );
NAND2_X1 U769 ( .A1(n1064), .A2(n1076), .ZN(n1071) );
INV_X1 U770 ( .A(n1042), .ZN(n1061) );
NOR3_X1 U771 ( .A1(n1077), .A2(G953), .A3(G952), .ZN(n1034) );
INV_X1 U772 ( .A(n1066), .ZN(n1077) );
NAND4_X1 U773 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1066) );
NOR4_X1 U774 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1081) );
XOR2_X1 U775 ( .A(n1086), .B(n1087), .Z(n1085) );
XNOR2_X1 U776 ( .A(n1088), .B(n1089), .ZN(n1082) );
NOR2_X1 U777 ( .A1(G475), .A2(KEYINPUT35), .ZN(n1089) );
NOR2_X1 U778 ( .A1(n1090), .A2(n1074), .ZN(n1080) );
XOR2_X1 U779 ( .A(n1091), .B(n1092), .Z(n1079) );
NOR2_X1 U780 ( .A1(n1093), .A2(KEYINPUT20), .ZN(n1092) );
XNOR2_X1 U781 ( .A(n1094), .B(n1095), .ZN(n1078) );
NOR2_X1 U782 ( .A1(n1096), .A2(KEYINPUT60), .ZN(n1095) );
NAND2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(G72) );
NAND2_X1 U784 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U785 ( .A(KEYINPUT38), .B(n1101), .ZN(n1100) );
XOR2_X1 U786 ( .A(n1102), .B(n1103), .Z(n1099) );
NAND2_X1 U787 ( .A1(n1104), .A2(n1105), .ZN(n1097) );
XNOR2_X1 U788 ( .A(n1102), .B(n1103), .ZN(n1105) );
NOR2_X1 U789 ( .A1(G953), .A2(n1106), .ZN(n1103) );
NAND2_X1 U790 ( .A1(n1107), .A2(n1108), .ZN(n1102) );
XOR2_X1 U791 ( .A(n1109), .B(n1110), .Z(n1107) );
XOR2_X1 U792 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U793 ( .A(n1113), .B(n1114), .Z(n1109) );
XOR2_X1 U794 ( .A(KEYINPUT47), .B(n1115), .Z(n1114) );
NOR2_X1 U795 ( .A1(G131), .A2(KEYINPUT9), .ZN(n1115) );
XOR2_X1 U796 ( .A(n1101), .B(KEYINPUT22), .Z(n1104) );
NAND2_X1 U797 ( .A1(n1108), .A2(n1116), .ZN(n1101) );
OR2_X1 U798 ( .A1(n1067), .A2(G227), .ZN(n1116) );
INV_X1 U799 ( .A(n1117), .ZN(n1108) );
XOR2_X1 U800 ( .A(n1118), .B(n1119), .Z(G69) );
XOR2_X1 U801 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR4_X1 U802 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1121) );
AND2_X1 U803 ( .A1(n1126), .A2(KEYINPUT28), .ZN(n1125) );
NOR2_X1 U804 ( .A1(G898), .A2(n1067), .ZN(n1124) );
NOR2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1123) );
NOR2_X1 U806 ( .A1(KEYINPUT28), .A2(n1129), .ZN(n1127) );
XNOR2_X1 U807 ( .A(n1126), .B(KEYINPUT21), .ZN(n1129) );
NOR3_X1 U808 ( .A1(n1130), .A2(KEYINPUT28), .A3(n1126), .ZN(n1122) );
NAND2_X1 U809 ( .A1(n1131), .A2(n1067), .ZN(n1120) );
NAND2_X1 U810 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XNOR2_X1 U811 ( .A(KEYINPUT13), .B(n1134), .ZN(n1133) );
NAND2_X1 U812 ( .A1(G953), .A2(n1135), .ZN(n1118) );
NAND2_X1 U813 ( .A1(G898), .A2(G224), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1136), .A2(n1137), .ZN(G66) );
NOR3_X1 U815 ( .A1(n1091), .A2(n1138), .A3(n1139), .ZN(n1137) );
AND3_X1 U816 ( .A1(n1140), .A2(n1093), .A3(n1141), .ZN(n1139) );
NOR2_X1 U817 ( .A1(n1142), .A2(n1140), .ZN(n1138) );
AND2_X1 U818 ( .A1(n1038), .A2(n1093), .ZN(n1142) );
NOR2_X1 U819 ( .A1(n1136), .A2(n1143), .ZN(G63) );
NOR2_X1 U820 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U821 ( .A(KEYINPUT31), .B(n1146), .Z(n1145) );
NOR2_X1 U822 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
AND2_X1 U823 ( .A1(n1148), .A2(n1147), .ZN(n1144) );
NAND2_X1 U824 ( .A1(n1141), .A2(G478), .ZN(n1148) );
NOR2_X1 U825 ( .A1(n1136), .A2(n1149), .ZN(G60) );
NOR3_X1 U826 ( .A1(n1088), .A2(n1150), .A3(n1151), .ZN(n1149) );
AND3_X1 U827 ( .A1(n1152), .A2(G475), .A3(n1141), .ZN(n1151) );
NOR2_X1 U828 ( .A1(n1153), .A2(n1152), .ZN(n1150) );
AND2_X1 U829 ( .A1(n1038), .A2(G475), .ZN(n1153) );
XOR2_X1 U830 ( .A(n1154), .B(n1155), .Z(G6) );
NAND4_X1 U831 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1064), .ZN(n1155) );
NOR2_X1 U832 ( .A1(n1159), .A2(n1057), .ZN(n1158) );
XOR2_X1 U833 ( .A(n1160), .B(KEYINPUT33), .Z(n1156) );
NOR2_X1 U834 ( .A1(n1136), .A2(n1161), .ZN(G57) );
XOR2_X1 U835 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U836 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(n1162) );
NAND2_X1 U838 ( .A1(KEYINPUT3), .A2(n1168), .ZN(n1167) );
XOR2_X1 U839 ( .A(n1169), .B(n1170), .Z(n1166) );
AND2_X1 U840 ( .A1(G472), .A2(n1141), .ZN(n1170) );
OR2_X1 U841 ( .A1(n1168), .A2(KEYINPUT3), .ZN(n1169) );
XNOR2_X1 U842 ( .A(n1171), .B(n1172), .ZN(n1168) );
NOR2_X1 U843 ( .A1(n1136), .A2(n1173), .ZN(G54) );
XOR2_X1 U844 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U845 ( .A(n1176), .B(n1177), .Z(n1175) );
AND2_X1 U846 ( .A1(G469), .A2(n1141), .ZN(n1176) );
XNOR2_X1 U847 ( .A(KEYINPUT37), .B(n1178), .ZN(n1174) );
NOR2_X1 U848 ( .A1(KEYINPUT6), .A2(n1179), .ZN(n1178) );
XNOR2_X1 U849 ( .A(n1180), .B(n1181), .ZN(n1179) );
NAND2_X1 U850 ( .A1(n1182), .A2(n1183), .ZN(n1180) );
XOR2_X1 U851 ( .A(KEYINPUT49), .B(n1184), .Z(n1182) );
NOR2_X1 U852 ( .A1(n1136), .A2(n1185), .ZN(G51) );
NOR3_X1 U853 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1185) );
AND2_X1 U854 ( .A1(n1189), .A2(KEYINPUT25), .ZN(n1188) );
NOR3_X1 U855 ( .A1(KEYINPUT25), .A2(n1190), .A3(n1189), .ZN(n1187) );
AND3_X1 U856 ( .A1(KEYINPUT41), .A2(n1096), .A3(n1141), .ZN(n1190) );
INV_X1 U857 ( .A(n1191), .ZN(n1141) );
NOR3_X1 U858 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1186) );
NOR2_X1 U859 ( .A1(n1194), .A2(KEYINPUT25), .ZN(n1192) );
AND2_X1 U860 ( .A1(n1189), .A2(KEYINPUT41), .ZN(n1194) );
XNOR2_X1 U861 ( .A(n1195), .B(n1196), .ZN(n1189) );
XOR2_X1 U862 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U863 ( .A(n1199), .B(G125), .Z(n1195) );
NAND2_X1 U864 ( .A1(KEYINPUT26), .A2(n1200), .ZN(n1199) );
NAND2_X1 U865 ( .A1(G902), .A2(n1038), .ZN(n1191) );
NAND3_X1 U866 ( .A1(n1132), .A2(n1134), .A3(n1106), .ZN(n1038) );
AND4_X1 U867 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1106) );
NOR4_X1 U868 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
INV_X1 U869 ( .A(n1209), .ZN(n1206) );
OR3_X1 U870 ( .A1(n1160), .A2(n1060), .A3(n1210), .ZN(n1203) );
NOR2_X1 U871 ( .A1(n1157), .A2(n1211), .ZN(n1060) );
NAND2_X1 U872 ( .A1(n1212), .A2(n1213), .ZN(n1134) );
XOR2_X1 U873 ( .A(KEYINPUT63), .B(n1051), .Z(n1213) );
AND4_X1 U874 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1132) );
NOR4_X1 U875 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1217) );
INV_X1 U876 ( .A(n1222), .ZN(n1219) );
OR2_X1 U877 ( .A1(n1033), .A2(KEYINPUT17), .ZN(n1216) );
NAND4_X1 U878 ( .A1(n1211), .A2(n1064), .A3(n1223), .A4(n1224), .ZN(n1033) );
NAND4_X1 U879 ( .A1(n1064), .A2(n1223), .A3(n1225), .A4(n1226), .ZN(n1215) );
OR2_X1 U880 ( .A1(n1159), .A2(n1157), .ZN(n1226) );
NAND2_X1 U881 ( .A1(n1159), .A2(n1227), .ZN(n1225) );
NAND2_X1 U882 ( .A1(KEYINPUT17), .A2(n1211), .ZN(n1227) );
NAND3_X1 U883 ( .A1(n1051), .A2(n1211), .A3(n1228), .ZN(n1214) );
INV_X1 U884 ( .A(n1229), .ZN(n1211) );
NOR2_X1 U885 ( .A1(n1067), .A2(G952), .ZN(n1136) );
XOR2_X1 U886 ( .A(n1230), .B(n1231), .Z(G48) );
XNOR2_X1 U887 ( .A(G146), .B(KEYINPUT5), .ZN(n1231) );
NAND4_X1 U888 ( .A1(KEYINPUT53), .A2(n1232), .A3(n1157), .A4(n1076), .ZN(n1230) );
INV_X1 U889 ( .A(n1210), .ZN(n1232) );
XOR2_X1 U890 ( .A(n1233), .B(n1202), .Z(G45) );
NAND3_X1 U891 ( .A1(n1051), .A2(n1223), .A3(n1234), .ZN(n1202) );
NOR3_X1 U892 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1234) );
XOR2_X1 U893 ( .A(n1238), .B(G140), .Z(G42) );
NAND2_X1 U894 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
OR2_X1 U895 ( .A1(n1201), .A2(KEYINPUT4), .ZN(n1240) );
NAND2_X1 U896 ( .A1(n1241), .A2(n1052), .ZN(n1201) );
NAND4_X1 U897 ( .A1(n1242), .A2(n1057), .A3(n1243), .A4(KEYINPUT4), .ZN(n1239) );
XOR2_X1 U898 ( .A(G137), .B(n1207), .Z(G39) );
NOR3_X1 U899 ( .A1(n1210), .A2(n1039), .A3(n1046), .ZN(n1207) );
XOR2_X1 U900 ( .A(n1244), .B(n1209), .Z(G36) );
NAND3_X1 U901 ( .A1(n1243), .A2(n1051), .A3(n1245), .ZN(n1209) );
NOR3_X1 U902 ( .A1(n1229), .A2(n1236), .A3(n1057), .ZN(n1245) );
INV_X1 U903 ( .A(n1246), .ZN(n1236) );
XOR2_X1 U904 ( .A(G131), .B(n1208), .Z(G33) );
AND2_X1 U905 ( .A1(n1241), .A2(n1051), .ZN(n1208) );
AND4_X1 U906 ( .A1(n1243), .A2(n1157), .A3(n1063), .A4(n1246), .ZN(n1241) );
INV_X1 U907 ( .A(n1039), .ZN(n1243) );
NAND2_X1 U908 ( .A1(n1073), .A2(n1247), .ZN(n1039) );
XOR2_X1 U909 ( .A(G128), .B(n1248), .Z(G30) );
NOR3_X1 U910 ( .A1(n1210), .A2(n1249), .A3(n1229), .ZN(n1248) );
XOR2_X1 U911 ( .A(n1160), .B(KEYINPUT45), .Z(n1249) );
NAND4_X1 U912 ( .A1(n1063), .A2(n1250), .A3(n1251), .A4(n1246), .ZN(n1210) );
XOR2_X1 U913 ( .A(n1252), .B(n1218), .Z(G3) );
AND4_X1 U914 ( .A1(n1065), .A2(n1051), .A3(n1223), .A4(n1224), .ZN(n1218) );
NAND2_X1 U915 ( .A1(KEYINPUT61), .A2(n1164), .ZN(n1252) );
INV_X1 U916 ( .A(G101), .ZN(n1164) );
XOR2_X1 U917 ( .A(n1205), .B(n1253), .Z(G27) );
NOR2_X1 U918 ( .A1(KEYINPUT42), .A2(n1254), .ZN(n1253) );
AND3_X1 U919 ( .A1(n1069), .A2(n1076), .A3(n1242), .ZN(n1205) );
AND3_X1 U920 ( .A1(n1157), .A2(n1246), .A3(n1052), .ZN(n1242) );
NAND2_X1 U921 ( .A1(n1042), .A2(n1255), .ZN(n1246) );
NAND3_X1 U922 ( .A1(G902), .A2(n1256), .A3(n1117), .ZN(n1255) );
NOR2_X1 U923 ( .A1(G900), .A2(n1067), .ZN(n1117) );
XOR2_X1 U924 ( .A(G122), .B(n1221), .Z(G24) );
AND4_X1 U925 ( .A1(n1228), .A2(n1064), .A3(n1084), .A4(n1257), .ZN(n1221) );
INV_X1 U926 ( .A(n1054), .ZN(n1064) );
NAND2_X1 U927 ( .A1(n1258), .A2(n1259), .ZN(n1054) );
XOR2_X1 U928 ( .A(n1220), .B(n1260), .Z(G21) );
NOR2_X1 U929 ( .A1(KEYINPUT16), .A2(n1261), .ZN(n1260) );
AND4_X1 U930 ( .A1(n1228), .A2(n1065), .A3(n1250), .A4(n1251), .ZN(n1220) );
XNOR2_X1 U931 ( .A(G116), .B(n1262), .ZN(G18) );
NAND3_X1 U932 ( .A1(n1263), .A2(n1051), .A3(n1264), .ZN(n1262) );
NOR3_X1 U933 ( .A1(n1050), .A2(n1159), .A3(n1229), .ZN(n1264) );
NAND2_X1 U934 ( .A1(n1237), .A2(n1084), .ZN(n1229) );
XOR2_X1 U935 ( .A(n1160), .B(KEYINPUT32), .Z(n1263) );
XNOR2_X1 U936 ( .A(G113), .B(n1265), .ZN(G15) );
NAND2_X1 U937 ( .A1(n1212), .A2(n1051), .ZN(n1265) );
AND2_X1 U938 ( .A1(n1250), .A2(n1259), .ZN(n1051) );
XOR2_X1 U939 ( .A(n1251), .B(KEYINPUT19), .Z(n1259) );
AND2_X1 U940 ( .A1(n1228), .A2(n1157), .ZN(n1212) );
NOR2_X1 U941 ( .A1(n1084), .A2(n1237), .ZN(n1157) );
INV_X1 U942 ( .A(n1235), .ZN(n1084) );
NOR3_X1 U943 ( .A1(n1160), .A2(n1159), .A3(n1050), .ZN(n1228) );
INV_X1 U944 ( .A(n1069), .ZN(n1050) );
NOR2_X1 U945 ( .A1(n1058), .A2(n1090), .ZN(n1069) );
XNOR2_X1 U946 ( .A(n1266), .B(KEYINPUT54), .ZN(n1058) );
INV_X1 U947 ( .A(n1224), .ZN(n1159) );
XOR2_X1 U948 ( .A(n1267), .B(n1222), .Z(G12) );
NAND4_X1 U949 ( .A1(n1065), .A2(n1052), .A3(n1223), .A4(n1224), .ZN(n1222) );
NAND2_X1 U950 ( .A1(n1042), .A2(n1268), .ZN(n1224) );
NAND4_X1 U951 ( .A1(G953), .A2(G902), .A3(n1256), .A4(n1269), .ZN(n1268) );
INV_X1 U952 ( .A(G898), .ZN(n1269) );
NAND3_X1 U953 ( .A1(n1256), .A2(n1067), .A3(G952), .ZN(n1042) );
NAND2_X1 U954 ( .A1(G237), .A2(G234), .ZN(n1256) );
NOR2_X1 U955 ( .A1(n1057), .A2(n1160), .ZN(n1223) );
INV_X1 U956 ( .A(n1076), .ZN(n1160) );
NOR2_X1 U957 ( .A1(n1073), .A2(n1074), .ZN(n1076) );
INV_X1 U958 ( .A(n1247), .ZN(n1074) );
NAND2_X1 U959 ( .A1(G214), .A2(n1270), .ZN(n1247) );
XOR2_X1 U960 ( .A(n1271), .B(n1096), .Z(n1073) );
INV_X1 U961 ( .A(n1193), .ZN(n1096) );
NAND2_X1 U962 ( .A1(G210), .A2(n1270), .ZN(n1193) );
NAND2_X1 U963 ( .A1(n1272), .A2(n1273), .ZN(n1270) );
INV_X1 U964 ( .A(G237), .ZN(n1272) );
XOR2_X1 U965 ( .A(n1094), .B(KEYINPUT29), .Z(n1271) );
NAND2_X1 U966 ( .A1(n1274), .A2(n1273), .ZN(n1094) );
XOR2_X1 U967 ( .A(n1275), .B(n1276), .Z(n1274) );
XNOR2_X1 U968 ( .A(n1200), .B(n1198), .ZN(n1276) );
XOR2_X1 U969 ( .A(n1128), .B(n1126), .Z(n1198) );
XNOR2_X1 U970 ( .A(n1277), .B(n1278), .ZN(n1126) );
XOR2_X1 U971 ( .A(G101), .B(n1279), .Z(n1278) );
XOR2_X1 U972 ( .A(G113), .B(G107), .Z(n1279) );
XNOR2_X1 U973 ( .A(n1280), .B(n1281), .ZN(n1277) );
NAND2_X1 U974 ( .A1(KEYINPUT43), .A2(n1154), .ZN(n1281) );
NAND3_X1 U975 ( .A1(n1282), .A2(n1283), .A3(KEYINPUT52), .ZN(n1280) );
NAND2_X1 U976 ( .A1(KEYINPUT50), .A2(n1284), .ZN(n1283) );
NAND3_X1 U977 ( .A1(G116), .A2(n1261), .A3(n1285), .ZN(n1282) );
INV_X1 U978 ( .A(KEYINPUT50), .ZN(n1285) );
INV_X1 U979 ( .A(n1130), .ZN(n1128) );
XNOR2_X1 U980 ( .A(G122), .B(n1286), .ZN(n1130) );
NOR2_X1 U981 ( .A1(G110), .A2(KEYINPUT46), .ZN(n1286) );
NAND2_X1 U982 ( .A1(G224), .A2(n1067), .ZN(n1200) );
XOR2_X1 U983 ( .A(n1287), .B(KEYINPUT2), .Z(n1275) );
NAND3_X1 U984 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n1287) );
NAND2_X1 U985 ( .A1(KEYINPUT30), .A2(n1254), .ZN(n1290) );
OR3_X1 U986 ( .A1(n1254), .A2(KEYINPUT30), .A3(n1291), .ZN(n1289) );
NAND2_X1 U987 ( .A1(n1291), .A2(n1292), .ZN(n1288) );
NAND2_X1 U988 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
INV_X1 U989 ( .A(KEYINPUT30), .ZN(n1294) );
XOR2_X1 U990 ( .A(KEYINPUT57), .B(G125), .Z(n1293) );
XOR2_X1 U991 ( .A(n1172), .B(KEYINPUT7), .Z(n1291) );
INV_X1 U992 ( .A(n1063), .ZN(n1057) );
NOR2_X1 U993 ( .A1(n1266), .A2(n1090), .ZN(n1063) );
INV_X1 U994 ( .A(n1059), .ZN(n1090) );
NAND2_X1 U995 ( .A1(G221), .A2(n1295), .ZN(n1059) );
NAND2_X1 U996 ( .A1(n1296), .A2(n1297), .ZN(n1266) );
NAND2_X1 U997 ( .A1(n1298), .A2(n1087), .ZN(n1297) );
XOR2_X1 U998 ( .A(n1086), .B(n1299), .Z(n1298) );
XNOR2_X1 U999 ( .A(KEYINPUT62), .B(KEYINPUT1), .ZN(n1299) );
NAND2_X1 U1000 ( .A1(n1300), .A2(n1301), .ZN(n1296) );
XOR2_X1 U1001 ( .A(n1086), .B(KEYINPUT51), .Z(n1301) );
NAND2_X1 U1002 ( .A1(n1302), .A2(n1273), .ZN(n1086) );
XNOR2_X1 U1003 ( .A(n1303), .B(n1177), .ZN(n1302) );
XNOR2_X1 U1004 ( .A(n1304), .B(n1305), .ZN(n1177) );
XOR2_X1 U1005 ( .A(G101), .B(n1306), .Z(n1305) );
NOR2_X1 U1006 ( .A1(KEYINPUT10), .A2(n1307), .ZN(n1306) );
XOR2_X1 U1007 ( .A(n1308), .B(n1309), .Z(n1307) );
XNOR2_X1 U1008 ( .A(G107), .B(KEYINPUT34), .ZN(n1309) );
NAND2_X1 U1009 ( .A1(KEYINPUT27), .A2(n1154), .ZN(n1308) );
INV_X1 U1010 ( .A(G104), .ZN(n1154) );
XOR2_X1 U1011 ( .A(n1310), .B(n1113), .Z(n1304) );
XOR2_X1 U1012 ( .A(G128), .B(n1311), .Z(n1113) );
NAND2_X1 U1013 ( .A1(n1312), .A2(n1313), .ZN(n1303) );
NAND2_X1 U1014 ( .A1(n1314), .A2(n1181), .ZN(n1313) );
OR2_X1 U1015 ( .A1(n1184), .A2(n1315), .ZN(n1314) );
XOR2_X1 U1016 ( .A(KEYINPUT8), .B(n1316), .Z(n1312) );
NOR3_X1 U1017 ( .A1(n1181), .A2(n1184), .A3(n1315), .ZN(n1316) );
INV_X1 U1018 ( .A(n1183), .ZN(n1315) );
NAND2_X1 U1019 ( .A1(G110), .A2(n1317), .ZN(n1183) );
NOR2_X1 U1020 ( .A1(n1317), .A2(G110), .ZN(n1184) );
NAND2_X1 U1021 ( .A1(G227), .A2(n1067), .ZN(n1181) );
INV_X1 U1022 ( .A(n1087), .ZN(n1300) );
XNOR2_X1 U1023 ( .A(G469), .B(KEYINPUT36), .ZN(n1087) );
AND2_X1 U1024 ( .A1(n1258), .A2(n1251), .ZN(n1052) );
XOR2_X1 U1025 ( .A(n1093), .B(n1091), .Z(n1251) );
NOR2_X1 U1026 ( .A1(n1140), .A2(G902), .ZN(n1091) );
XOR2_X1 U1027 ( .A(n1318), .B(n1319), .Z(n1140) );
XNOR2_X1 U1028 ( .A(n1320), .B(n1112), .ZN(n1319) );
NAND2_X1 U1029 ( .A1(G221), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1030 ( .A(n1322), .B(n1323), .Z(n1318) );
NOR2_X1 U1031 ( .A1(KEYINPUT55), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1032 ( .A(n1267), .B(n1325), .Z(n1324) );
XOR2_X1 U1033 ( .A(G128), .B(G119), .Z(n1325) );
XNOR2_X1 U1034 ( .A(G137), .B(G146), .ZN(n1322) );
AND2_X1 U1035 ( .A1(G217), .A2(n1295), .ZN(n1093) );
NAND2_X1 U1036 ( .A1(G234), .A2(n1273), .ZN(n1295) );
XOR2_X1 U1037 ( .A(KEYINPUT23), .B(n1250), .Z(n1258) );
XOR2_X1 U1038 ( .A(n1083), .B(KEYINPUT24), .Z(n1250) );
XNOR2_X1 U1039 ( .A(n1326), .B(G472), .ZN(n1083) );
NAND2_X1 U1040 ( .A1(n1327), .A2(n1273), .ZN(n1326) );
XOR2_X1 U1041 ( .A(n1165), .B(n1328), .Z(n1327) );
XNOR2_X1 U1042 ( .A(n1329), .B(n1330), .ZN(n1328) );
NOR2_X1 U1043 ( .A1(KEYINPUT0), .A2(G101), .ZN(n1330) );
NAND3_X1 U1044 ( .A1(n1331), .A2(n1332), .A3(KEYINPUT44), .ZN(n1329) );
NAND2_X1 U1045 ( .A1(n1197), .A2(n1171), .ZN(n1332) );
INV_X1 U1046 ( .A(n1172), .ZN(n1197) );
NAND2_X1 U1047 ( .A1(n1333), .A2(n1172), .ZN(n1331) );
XOR2_X1 U1048 ( .A(n1334), .B(G128), .Z(n1172) );
NAND2_X1 U1049 ( .A1(KEYINPUT48), .A2(n1311), .ZN(n1334) );
XOR2_X1 U1050 ( .A(G143), .B(G146), .Z(n1311) );
XOR2_X1 U1051 ( .A(n1171), .B(KEYINPUT59), .Z(n1333) );
XOR2_X1 U1052 ( .A(n1310), .B(n1335), .Z(n1171) );
XNOR2_X1 U1053 ( .A(G113), .B(n1284), .ZN(n1335) );
XOR2_X1 U1054 ( .A(G116), .B(n1261), .Z(n1284) );
INV_X1 U1055 ( .A(G119), .ZN(n1261) );
XOR2_X1 U1056 ( .A(n1336), .B(n1111), .Z(n1310) );
XOR2_X1 U1057 ( .A(G134), .B(G137), .Z(n1111) );
NAND2_X1 U1058 ( .A1(KEYINPUT58), .A2(n1337), .ZN(n1336) );
NAND2_X1 U1059 ( .A1(G210), .A2(n1338), .ZN(n1165) );
INV_X1 U1060 ( .A(n1046), .ZN(n1065) );
NAND2_X1 U1061 ( .A1(n1235), .A2(n1237), .ZN(n1046) );
INV_X1 U1062 ( .A(n1257), .ZN(n1237) );
XOR2_X1 U1063 ( .A(n1088), .B(G475), .Z(n1257) );
NOR2_X1 U1064 ( .A1(n1152), .A2(G902), .ZN(n1088) );
XNOR2_X1 U1065 ( .A(n1339), .B(n1340), .ZN(n1152) );
XOR2_X1 U1066 ( .A(G104), .B(n1341), .Z(n1340) );
XOR2_X1 U1067 ( .A(G122), .B(G113), .Z(n1341) );
XOR2_X1 U1068 ( .A(n1342), .B(n1343), .Z(n1339) );
NOR2_X1 U1069 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
XOR2_X1 U1070 ( .A(n1346), .B(KEYINPUT40), .Z(n1345) );
NAND2_X1 U1071 ( .A1(n1347), .A2(n1337), .ZN(n1346) );
NOR2_X1 U1072 ( .A1(n1347), .A2(n1337), .ZN(n1344) );
INV_X1 U1073 ( .A(G131), .ZN(n1337) );
XOR2_X1 U1074 ( .A(n1348), .B(n1233), .Z(n1347) );
INV_X1 U1075 ( .A(G143), .ZN(n1233) );
NAND2_X1 U1076 ( .A1(G214), .A2(n1338), .ZN(n1348) );
NOR2_X1 U1077 ( .A1(G953), .A2(G237), .ZN(n1338) );
NAND2_X1 U1078 ( .A1(KEYINPUT15), .A2(n1349), .ZN(n1342) );
XOR2_X1 U1079 ( .A(G146), .B(n1350), .Z(n1349) );
NOR3_X1 U1080 ( .A1(KEYINPUT11), .A2(n1351), .A3(n1352), .ZN(n1350) );
AND3_X1 U1081 ( .A1(KEYINPUT14), .A2(n1254), .A3(G140), .ZN(n1352) );
NOR2_X1 U1082 ( .A1(KEYINPUT14), .A2(n1112), .ZN(n1351) );
XOR2_X1 U1083 ( .A(n1317), .B(n1254), .Z(n1112) );
INV_X1 U1084 ( .A(G125), .ZN(n1254) );
INV_X1 U1085 ( .A(G140), .ZN(n1317) );
XOR2_X1 U1086 ( .A(n1353), .B(G478), .Z(n1235) );
NAND2_X1 U1087 ( .A1(n1147), .A2(n1273), .ZN(n1353) );
INV_X1 U1088 ( .A(G902), .ZN(n1273) );
XNOR2_X1 U1089 ( .A(n1354), .B(n1355), .ZN(n1147) );
XOR2_X1 U1090 ( .A(n1356), .B(n1357), .Z(n1355) );
XOR2_X1 U1091 ( .A(n1358), .B(n1359), .Z(n1357) );
NOR2_X1 U1092 ( .A1(KEYINPUT18), .A2(G116), .ZN(n1359) );
NAND2_X1 U1093 ( .A1(G217), .A2(n1321), .ZN(n1358) );
AND2_X1 U1094 ( .A1(G234), .A2(n1067), .ZN(n1321) );
INV_X1 U1095 ( .A(G953), .ZN(n1067) );
NAND2_X1 U1096 ( .A1(KEYINPUT39), .A2(n1360), .ZN(n1356) );
INV_X1 U1097 ( .A(G128), .ZN(n1360) );
XOR2_X1 U1098 ( .A(n1361), .B(n1362), .Z(n1354) );
XOR2_X1 U1099 ( .A(G122), .B(G107), .Z(n1362) );
XOR2_X1 U1100 ( .A(n1244), .B(G143), .Z(n1361) );
INV_X1 U1101 ( .A(G134), .ZN(n1244) );
INV_X1 U1102 ( .A(G110), .ZN(n1267) );
endmodule


