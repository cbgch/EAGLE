//Key = 0001010110010000101111001110000111010000001001110100110010100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301;

XOR2_X1 U715 ( .A(G107), .B(n993), .Z(G9) );
NOR2_X1 U716 ( .A1(n994), .A2(n995), .ZN(n993) );
XOR2_X1 U717 ( .A(n996), .B(KEYINPUT27), .Z(n994) );
NAND4_X1 U718 ( .A1(n997), .A2(n998), .A3(n999), .A4(n1000), .ZN(n996) );
XOR2_X1 U719 ( .A(KEYINPUT60), .B(n1001), .Z(n999) );
NOR2_X1 U720 ( .A1(n1002), .A2(n1003), .ZN(G75) );
NOR3_X1 U721 ( .A1(n1004), .A2(G953), .A3(G952), .ZN(n1003) );
NOR3_X1 U722 ( .A1(n1005), .A2(n1004), .A3(n1006), .ZN(n1002) );
AND4_X1 U723 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1004) );
NOR4_X1 U724 ( .A1(n1011), .A2(n1012), .A3(n1013), .A4(n1014), .ZN(n1010) );
XOR2_X1 U725 ( .A(n1015), .B(KEYINPUT47), .Z(n1012) );
XOR2_X1 U726 ( .A(n1016), .B(G469), .Z(n1009) );
XOR2_X1 U727 ( .A(n1017), .B(KEYINPUT29), .Z(n1007) );
NAND3_X1 U728 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1005) );
NAND4_X1 U729 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1020) );
NAND2_X1 U730 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND3_X1 U731 ( .A1(n997), .A2(n1027), .A3(n1022), .ZN(n1018) );
INV_X1 U732 ( .A(n1028), .ZN(n1022) );
NAND2_X1 U733 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NAND2_X1 U734 ( .A1(n1023), .A2(n1031), .ZN(n1030) );
NAND2_X1 U735 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND3_X1 U736 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
INV_X1 U737 ( .A(KEYINPUT26), .ZN(n1035) );
NAND2_X1 U738 ( .A1(n1037), .A2(n1038), .ZN(n1032) );
NAND3_X1 U739 ( .A1(n1039), .A2(n995), .A3(n1040), .ZN(n1038) );
NAND2_X1 U740 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
INV_X1 U741 ( .A(n1043), .ZN(n995) );
NAND2_X1 U742 ( .A1(n1008), .A2(n1044), .ZN(n1039) );
INV_X1 U743 ( .A(KEYINPUT21), .ZN(n1044) );
NAND2_X1 U744 ( .A1(n1008), .A2(n1034), .ZN(n1029) );
NAND3_X1 U745 ( .A1(n1045), .A2(n1046), .A3(n1008), .ZN(n1034) );
NAND2_X1 U746 ( .A1(n1023), .A2(n1047), .ZN(n1046) );
NAND2_X1 U747 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U748 ( .A1(KEYINPUT26), .A2(n1036), .ZN(n1049) );
XOR2_X1 U749 ( .A(KEYINPUT33), .B(n998), .Z(n1048) );
NAND2_X1 U750 ( .A1(n1037), .A2(n1050), .ZN(n1045) );
NAND2_X1 U751 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
INV_X1 U752 ( .A(n1001), .ZN(n1052) );
NAND3_X1 U753 ( .A1(n1053), .A2(n1011), .A3(KEYINPUT21), .ZN(n1051) );
XOR2_X1 U754 ( .A(n1054), .B(n1055), .Z(G72) );
NOR2_X1 U755 ( .A1(n1056), .A2(G953), .ZN(n1055) );
NAND2_X1 U756 ( .A1(n1057), .A2(n1058), .ZN(n1054) );
NAND2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
INV_X1 U758 ( .A(n1061), .ZN(n1059) );
NAND2_X1 U759 ( .A1(n1062), .A2(n1061), .ZN(n1057) );
NAND2_X1 U760 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
XOR2_X1 U761 ( .A(n1065), .B(n1066), .Z(n1063) );
XOR2_X1 U762 ( .A(n1067), .B(n1068), .Z(n1066) );
NOR2_X1 U763 ( .A1(G137), .A2(KEYINPUT14), .ZN(n1067) );
XOR2_X1 U764 ( .A(n1069), .B(n1070), .Z(n1065) );
NOR4_X1 U765 ( .A1(n1071), .A2(n1072), .A3(KEYINPUT22), .A4(n1073), .ZN(n1070) );
INV_X1 U766 ( .A(n1074), .ZN(n1073) );
NOR2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(n1072) );
INV_X1 U768 ( .A(KEYINPUT42), .ZN(n1076) );
NOR2_X1 U769 ( .A1(KEYINPUT42), .A2(G125), .ZN(n1071) );
XOR2_X1 U770 ( .A(n1077), .B(G134), .Z(n1069) );
NAND2_X1 U771 ( .A1(n1064), .A2(n1060), .ZN(n1062) );
NAND2_X1 U772 ( .A1(G953), .A2(n1078), .ZN(n1060) );
INV_X1 U773 ( .A(n1079), .ZN(n1064) );
NAND2_X1 U774 ( .A1(n1080), .A2(n1081), .ZN(G69) );
NAND3_X1 U775 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
XNOR2_X1 U776 ( .A(n1085), .B(n1086), .ZN(n1084) );
NAND2_X1 U777 ( .A1(n1019), .A2(n1087), .ZN(n1086) );
NAND2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XNOR2_X1 U779 ( .A(n1090), .B(KEYINPUT46), .ZN(n1088) );
NAND2_X1 U780 ( .A1(G953), .A2(n1091), .ZN(n1082) );
NAND3_X1 U781 ( .A1(n1092), .A2(n1093), .A3(G953), .ZN(n1080) );
NAND2_X1 U782 ( .A1(n1085), .A2(n1083), .ZN(n1093) );
INV_X1 U783 ( .A(KEYINPUT1), .ZN(n1083) );
NOR3_X1 U784 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1085) );
INV_X1 U785 ( .A(n1097), .ZN(n1095) );
NAND2_X1 U786 ( .A1(G898), .A2(G224), .ZN(n1092) );
NOR2_X1 U787 ( .A1(n1098), .A2(n1099), .ZN(G66) );
XOR2_X1 U788 ( .A(n1100), .B(n1101), .Z(n1099) );
NAND2_X1 U789 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
XOR2_X1 U790 ( .A(KEYINPUT9), .B(n1104), .Z(n1103) );
NOR2_X1 U791 ( .A1(n1098), .A2(n1105), .ZN(G63) );
XOR2_X1 U792 ( .A(n1106), .B(n1107), .Z(n1105) );
NAND2_X1 U793 ( .A1(n1102), .A2(G478), .ZN(n1106) );
NOR2_X1 U794 ( .A1(n1098), .A2(n1108), .ZN(G60) );
NOR2_X1 U795 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U796 ( .A(n1111), .B(n1112), .Z(n1110) );
NAND2_X1 U797 ( .A1(n1102), .A2(G475), .ZN(n1112) );
NAND2_X1 U798 ( .A1(KEYINPUT16), .A2(n1113), .ZN(n1111) );
NOR2_X1 U799 ( .A1(KEYINPUT16), .A2(n1113), .ZN(n1109) );
XNOR2_X1 U800 ( .A(G104), .B(n1114), .ZN(G6) );
NAND4_X1 U801 ( .A1(n1115), .A2(n1000), .A3(n1001), .A4(n1116), .ZN(n1114) );
AND2_X1 U802 ( .A1(n997), .A2(n1036), .ZN(n1116) );
XOR2_X1 U803 ( .A(KEYINPUT23), .B(n1043), .Z(n1115) );
NOR2_X1 U804 ( .A1(n1098), .A2(n1117), .ZN(G57) );
XOR2_X1 U805 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U806 ( .A1(KEYINPUT30), .A2(n1120), .ZN(n1119) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
XOR2_X1 U808 ( .A(KEYINPUT2), .B(n1123), .Z(n1122) );
AND3_X1 U809 ( .A1(n1102), .A2(n1124), .A3(G472), .ZN(n1123) );
NOR2_X1 U810 ( .A1(n1125), .A2(n1124), .ZN(n1121) );
XOR2_X1 U811 ( .A(n1126), .B(n1127), .Z(n1124) );
XOR2_X1 U812 ( .A(n1128), .B(KEYINPUT8), .Z(n1126) );
AND2_X1 U813 ( .A1(G472), .A2(n1102), .ZN(n1125) );
NOR2_X1 U814 ( .A1(n1098), .A2(n1129), .ZN(G54) );
XOR2_X1 U815 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U816 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U817 ( .A1(KEYINPUT63), .A2(n1134), .ZN(n1132) );
XOR2_X1 U818 ( .A(n1135), .B(n1136), .Z(n1130) );
NAND2_X1 U819 ( .A1(KEYINPUT18), .A2(n1137), .ZN(n1136) );
NAND2_X1 U820 ( .A1(n1102), .A2(G469), .ZN(n1135) );
INV_X1 U821 ( .A(n1138), .ZN(n1102) );
NOR2_X1 U822 ( .A1(n1098), .A2(n1139), .ZN(G51) );
XOR2_X1 U823 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U824 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR3_X1 U825 ( .A1(n1138), .A2(KEYINPUT51), .A3(n1144), .ZN(n1143) );
NAND2_X1 U826 ( .A1(G902), .A2(n1006), .ZN(n1138) );
NAND3_X1 U827 ( .A1(n1056), .A2(n1090), .A3(n1089), .ZN(n1006) );
AND3_X1 U828 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(n1089) );
NAND3_X1 U829 ( .A1(n997), .A2(n1148), .A3(n1149), .ZN(n1147) );
NAND2_X1 U830 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
NOR4_X1 U831 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1090) );
NOR2_X1 U832 ( .A1(n1156), .A2(n1157), .ZN(n1152) );
AND4_X1 U833 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1056) );
AND4_X1 U834 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1161) );
NAND2_X1 U835 ( .A1(n1166), .A2(n1167), .ZN(n1160) );
NAND2_X1 U836 ( .A1(n1168), .A2(n1026), .ZN(n1167) );
XOR2_X1 U837 ( .A(KEYINPUT52), .B(n1169), .Z(n1168) );
INV_X1 U838 ( .A(n1170), .ZN(n1166) );
NAND2_X1 U839 ( .A1(n1171), .A2(n1021), .ZN(n1158) );
XOR2_X1 U840 ( .A(n1172), .B(n1173), .Z(n1140) );
NOR2_X1 U841 ( .A1(n1019), .A2(G952), .ZN(n1098) );
XNOR2_X1 U842 ( .A(G146), .B(n1159), .ZN(G48) );
NAND3_X1 U843 ( .A1(n1036), .A2(n1043), .A3(n1171), .ZN(n1159) );
XOR2_X1 U844 ( .A(n1174), .B(n1165), .Z(G45) );
NAND4_X1 U845 ( .A1(n1175), .A2(n1043), .A3(n1013), .A4(n1176), .ZN(n1165) );
NAND2_X1 U846 ( .A1(n1177), .A2(n1178), .ZN(G42) );
NAND2_X1 U847 ( .A1(G140), .A2(n1179), .ZN(n1178) );
XOR2_X1 U848 ( .A(n1180), .B(n1181), .Z(n1177) );
NOR2_X1 U849 ( .A1(n1025), .A2(n1170), .ZN(n1181) );
INV_X1 U850 ( .A(n1169), .ZN(n1025) );
NOR2_X1 U851 ( .A1(G140), .A2(n1179), .ZN(n1180) );
INV_X1 U852 ( .A(KEYINPUT58), .ZN(n1179) );
XNOR2_X1 U853 ( .A(G137), .B(n1182), .ZN(G39) );
NAND3_X1 U854 ( .A1(n1021), .A2(n1183), .A3(n1171), .ZN(n1182) );
XOR2_X1 U855 ( .A(KEYINPUT5), .B(KEYINPUT48), .Z(n1183) );
AND2_X1 U856 ( .A1(n1008), .A2(n1037), .ZN(n1021) );
XOR2_X1 U857 ( .A(n1184), .B(n1164), .Z(G36) );
NAND3_X1 U858 ( .A1(n1008), .A2(n998), .A3(n1175), .ZN(n1164) );
AND3_X1 U859 ( .A1(n1001), .A2(n1185), .A3(n1186), .ZN(n1175) );
XOR2_X1 U860 ( .A(G131), .B(n1187), .Z(G33) );
NOR3_X1 U861 ( .A1(n1170), .A2(KEYINPUT15), .A3(n1026), .ZN(n1187) );
NAND4_X1 U862 ( .A1(n1008), .A2(n1036), .A3(n1001), .A4(n1185), .ZN(n1170) );
NOR2_X1 U863 ( .A1(n1188), .A2(n1041), .ZN(n1008) );
INV_X1 U864 ( .A(n1042), .ZN(n1188) );
XNOR2_X1 U865 ( .A(G128), .B(n1163), .ZN(G30) );
NAND3_X1 U866 ( .A1(n1043), .A2(n998), .A3(n1171), .ZN(n1163) );
AND4_X1 U867 ( .A1(n1001), .A2(n1189), .A3(n1014), .A4(n1185), .ZN(n1171) );
INV_X1 U868 ( .A(n1151), .ZN(n998) );
XOR2_X1 U869 ( .A(n1190), .B(n1145), .Z(G3) );
NAND3_X1 U870 ( .A1(n1149), .A2(n1037), .A3(n1186), .ZN(n1145) );
INV_X1 U871 ( .A(n1026), .ZN(n1186) );
XOR2_X1 U872 ( .A(n1191), .B(n1162), .Z(G27) );
NAND4_X1 U873 ( .A1(n1043), .A2(n1185), .A3(n1036), .A4(n1192), .ZN(n1162) );
AND2_X1 U874 ( .A1(n1023), .A2(n1169), .ZN(n1192) );
INV_X1 U875 ( .A(n1150), .ZN(n1036) );
NAND2_X1 U876 ( .A1(n1193), .A2(n1194), .ZN(n1185) );
NAND3_X1 U877 ( .A1(G902), .A2(n1195), .A3(n1079), .ZN(n1194) );
NOR2_X1 U878 ( .A1(G900), .A2(n1019), .ZN(n1079) );
XOR2_X1 U879 ( .A(n1028), .B(KEYINPUT12), .Z(n1193) );
XOR2_X1 U880 ( .A(n1196), .B(n1197), .Z(G24) );
XOR2_X1 U881 ( .A(KEYINPUT41), .B(G122), .Z(n1197) );
NOR3_X1 U882 ( .A1(n1156), .A2(n1198), .A3(n1157), .ZN(n1196) );
XNOR2_X1 U883 ( .A(KEYINPUT36), .B(KEYINPUT25), .ZN(n1198) );
NAND3_X1 U884 ( .A1(n1013), .A2(n1176), .A3(n997), .ZN(n1156) );
NOR2_X1 U885 ( .A1(n1014), .A2(n1189), .ZN(n997) );
XOR2_X1 U886 ( .A(G119), .B(n1153), .Z(G21) );
AND4_X1 U887 ( .A1(n1199), .A2(n1037), .A3(n1189), .A4(n1014), .ZN(n1153) );
INV_X1 U888 ( .A(n1017), .ZN(n1189) );
INV_X1 U889 ( .A(n1157), .ZN(n1199) );
XOR2_X1 U890 ( .A(G116), .B(n1154), .Z(G18) );
NOR3_X1 U891 ( .A1(n1026), .A2(n1151), .A3(n1157), .ZN(n1154) );
NAND2_X1 U892 ( .A1(n1015), .A2(n1013), .ZN(n1151) );
XOR2_X1 U893 ( .A(G113), .B(n1155), .Z(G15) );
NOR3_X1 U894 ( .A1(n1026), .A2(n1150), .A3(n1157), .ZN(n1155) );
NAND3_X1 U895 ( .A1(n1043), .A2(n1000), .A3(n1023), .ZN(n1157) );
NOR2_X1 U896 ( .A1(n1200), .A2(n1011), .ZN(n1023) );
INV_X1 U897 ( .A(n1053), .ZN(n1200) );
NAND2_X1 U898 ( .A1(n1201), .A2(n1176), .ZN(n1150) );
NAND2_X1 U899 ( .A1(n1017), .A2(n1014), .ZN(n1026) );
XNOR2_X1 U900 ( .A(G110), .B(n1146), .ZN(G12) );
NAND3_X1 U901 ( .A1(n1149), .A2(n1037), .A3(n1169), .ZN(n1146) );
NOR2_X1 U902 ( .A1(n1014), .A2(n1017), .ZN(n1169) );
XOR2_X1 U903 ( .A(n1202), .B(n1104), .Z(n1017) );
AND2_X1 U904 ( .A1(G217), .A2(n1203), .ZN(n1104) );
NAND2_X1 U905 ( .A1(n1101), .A2(n1204), .ZN(n1202) );
XOR2_X1 U906 ( .A(n1205), .B(n1206), .Z(n1101) );
XOR2_X1 U907 ( .A(n1207), .B(n1208), .Z(n1206) );
XOR2_X1 U908 ( .A(G128), .B(n1209), .Z(n1208) );
NOR2_X1 U909 ( .A1(KEYINPUT59), .A2(n1210), .ZN(n1209) );
XOR2_X1 U910 ( .A(KEYINPUT50), .B(G119), .Z(n1210) );
XOR2_X1 U911 ( .A(G146), .B(G137), .Z(n1207) );
XOR2_X1 U912 ( .A(n1211), .B(n1212), .Z(n1205) );
XOR2_X1 U913 ( .A(n1213), .B(n1214), .Z(n1212) );
NAND2_X1 U914 ( .A1(G221), .A2(n1215), .ZN(n1214) );
NAND3_X1 U915 ( .A1(n1074), .A2(n1075), .A3(KEYINPUT3), .ZN(n1213) );
XNOR2_X1 U916 ( .A(n1216), .B(G472), .ZN(n1014) );
NAND2_X1 U917 ( .A1(n1217), .A2(n1204), .ZN(n1216) );
XOR2_X1 U918 ( .A(n1218), .B(n1219), .Z(n1217) );
NOR2_X1 U919 ( .A1(KEYINPUT34), .A2(n1127), .ZN(n1219) );
XNOR2_X1 U920 ( .A(n1220), .B(n1221), .ZN(n1127) );
XNOR2_X1 U921 ( .A(n1134), .B(KEYINPUT7), .ZN(n1220) );
XOR2_X1 U922 ( .A(n1128), .B(n1222), .Z(n1218) );
NOR2_X1 U923 ( .A1(KEYINPUT39), .A2(n1223), .ZN(n1222) );
XOR2_X1 U924 ( .A(KEYINPUT31), .B(n1120), .Z(n1223) );
XOR2_X1 U925 ( .A(n1224), .B(n1190), .Z(n1120) );
NAND2_X1 U926 ( .A1(n1225), .A2(G210), .ZN(n1224) );
NAND2_X1 U927 ( .A1(n1226), .A2(n1227), .ZN(n1128) );
NAND2_X1 U928 ( .A1(G113), .A2(n1228), .ZN(n1227) );
XOR2_X1 U929 ( .A(n1229), .B(KEYINPUT13), .Z(n1226) );
OR2_X1 U930 ( .A1(n1228), .A2(G113), .ZN(n1229) );
XNOR2_X1 U931 ( .A(n1230), .B(G116), .ZN(n1228) );
NAND2_X1 U932 ( .A1(KEYINPUT56), .A2(G119), .ZN(n1230) );
NOR2_X1 U933 ( .A1(n1013), .A2(n1176), .ZN(n1037) );
INV_X1 U934 ( .A(n1015), .ZN(n1176) );
XOR2_X1 U935 ( .A(n1231), .B(G475), .Z(n1015) );
NAND2_X1 U936 ( .A1(n1113), .A2(n1204), .ZN(n1231) );
XOR2_X1 U937 ( .A(n1232), .B(n1233), .Z(n1113) );
XOR2_X1 U938 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U939 ( .A(n1236), .B(n1237), .Z(n1235) );
NOR4_X1 U940 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1237) );
AND3_X1 U941 ( .A1(KEYINPUT11), .A2(n1242), .A3(n1191), .ZN(n1241) );
NOR2_X1 U942 ( .A1(KEYINPUT11), .A2(n1074), .ZN(n1240) );
NAND2_X1 U943 ( .A1(G140), .A2(n1191), .ZN(n1074) );
INV_X1 U944 ( .A(G125), .ZN(n1191) );
AND3_X1 U945 ( .A1(KEYINPUT49), .A2(G125), .A3(G140), .ZN(n1239) );
NOR2_X1 U946 ( .A1(KEYINPUT49), .A2(n1075), .ZN(n1238) );
NAND2_X1 U947 ( .A1(G125), .A2(n1242), .ZN(n1075) );
INV_X1 U948 ( .A(G140), .ZN(n1242) );
NOR2_X1 U949 ( .A1(KEYINPUT28), .A2(n1243), .ZN(n1236) );
XOR2_X1 U950 ( .A(n1077), .B(n1244), .Z(n1243) );
NAND2_X1 U951 ( .A1(KEYINPUT35), .A2(n1245), .ZN(n1244) );
XOR2_X1 U952 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U953 ( .A(n1174), .B(KEYINPUT53), .Z(n1247) );
INV_X1 U954 ( .A(G143), .ZN(n1174) );
NAND2_X1 U955 ( .A1(n1225), .A2(G214), .ZN(n1246) );
NOR2_X1 U956 ( .A1(G953), .A2(G237), .ZN(n1225) );
NOR2_X1 U957 ( .A1(G146), .A2(KEYINPUT0), .ZN(n1234) );
XNOR2_X1 U958 ( .A(G104), .B(n1248), .ZN(n1232) );
XOR2_X1 U959 ( .A(G122), .B(G113), .Z(n1248) );
INV_X1 U960 ( .A(n1201), .ZN(n1013) );
XOR2_X1 U961 ( .A(n1249), .B(G478), .Z(n1201) );
NAND2_X1 U962 ( .A1(n1107), .A2(n1204), .ZN(n1249) );
XOR2_X1 U963 ( .A(n1250), .B(n1251), .Z(n1107) );
XOR2_X1 U964 ( .A(n1252), .B(n1253), .Z(n1251) );
AND2_X1 U965 ( .A1(G217), .A2(n1215), .ZN(n1253) );
AND2_X1 U966 ( .A1(G234), .A2(n1019), .ZN(n1215) );
NOR2_X1 U967 ( .A1(KEYINPUT62), .A2(n1254), .ZN(n1252) );
XOR2_X1 U968 ( .A(G134), .B(n1255), .Z(n1254) );
NOR2_X1 U969 ( .A1(KEYINPUT37), .A2(n1256), .ZN(n1255) );
XOR2_X1 U970 ( .A(KEYINPUT20), .B(n1257), .Z(n1256) );
XNOR2_X1 U971 ( .A(G107), .B(n1258), .ZN(n1250) );
XOR2_X1 U972 ( .A(G122), .B(G116), .Z(n1258) );
AND3_X1 U973 ( .A1(n1001), .A2(n1000), .A3(n1043), .ZN(n1149) );
NOR2_X1 U974 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
AND2_X1 U975 ( .A1(G214), .A2(n1259), .ZN(n1041) );
XNOR2_X1 U976 ( .A(n1260), .B(n1144), .ZN(n1042) );
NAND2_X1 U977 ( .A1(G210), .A2(n1259), .ZN(n1144) );
NAND2_X1 U978 ( .A1(n1261), .A2(n1204), .ZN(n1259) );
INV_X1 U979 ( .A(G237), .ZN(n1261) );
NAND3_X1 U980 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1260) );
XOR2_X1 U981 ( .A(n1265), .B(KEYINPUT38), .Z(n1264) );
OR2_X1 U982 ( .A1(n1172), .A2(n1266), .ZN(n1265) );
NAND2_X1 U983 ( .A1(n1266), .A2(n1172), .ZN(n1263) );
NAND3_X1 U984 ( .A1(n1267), .A2(n1268), .A3(n1097), .ZN(n1172) );
NAND2_X1 U985 ( .A1(n1269), .A2(n1270), .ZN(n1097) );
NAND2_X1 U986 ( .A1(n1094), .A2(n1271), .ZN(n1268) );
INV_X1 U987 ( .A(KEYINPUT61), .ZN(n1271) );
NOR2_X1 U988 ( .A1(n1270), .A2(n1269), .ZN(n1094) );
XNOR2_X1 U989 ( .A(n1272), .B(n1273), .ZN(n1270) );
XOR2_X1 U990 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U991 ( .A(n1276), .B(n1277), .ZN(n1275) );
NOR2_X1 U992 ( .A1(KEYINPUT44), .A2(n1190), .ZN(n1277) );
INV_X1 U993 ( .A(G101), .ZN(n1190) );
NOR2_X1 U994 ( .A1(KEYINPUT10), .A2(n1278), .ZN(n1276) );
XOR2_X1 U995 ( .A(KEYINPUT40), .B(G119), .Z(n1278) );
XOR2_X1 U996 ( .A(n1279), .B(n1280), .Z(n1272) );
XOR2_X1 U997 ( .A(KEYINPUT45), .B(G116), .Z(n1280) );
INV_X1 U998 ( .A(G113), .ZN(n1279) );
NAND2_X1 U999 ( .A1(KEYINPUT61), .A2(n1269), .ZN(n1267) );
XOR2_X1 U1000 ( .A(n1211), .B(n1281), .Z(n1269) );
NOR2_X1 U1001 ( .A1(G122), .A2(KEYINPUT6), .ZN(n1281) );
XNOR2_X1 U1002 ( .A(n1282), .B(n1283), .ZN(n1266) );
NOR2_X1 U1003 ( .A1(KEYINPUT57), .A2(n1142), .ZN(n1283) );
XOR2_X1 U1004 ( .A(n1221), .B(G125), .Z(n1142) );
XOR2_X1 U1005 ( .A(n1284), .B(n1257), .Z(n1221) );
XOR2_X1 U1006 ( .A(G128), .B(G143), .Z(n1257) );
NAND2_X1 U1007 ( .A1(KEYINPUT19), .A2(G146), .ZN(n1284) );
XNOR2_X1 U1008 ( .A(n1173), .B(KEYINPUT17), .ZN(n1282) );
NOR2_X1 U1009 ( .A1(n1091), .A2(G953), .ZN(n1173) );
INV_X1 U1010 ( .A(G224), .ZN(n1091) );
XOR2_X1 U1011 ( .A(n1204), .B(KEYINPUT43), .Z(n1262) );
NAND2_X1 U1012 ( .A1(n1028), .A2(n1285), .ZN(n1000) );
NAND3_X1 U1013 ( .A1(G902), .A2(n1195), .A3(n1096), .ZN(n1285) );
NOR2_X1 U1014 ( .A1(n1019), .A2(G898), .ZN(n1096) );
NAND3_X1 U1015 ( .A1(n1195), .A2(n1019), .A3(G952), .ZN(n1028) );
INV_X1 U1016 ( .A(G953), .ZN(n1019) );
NAND2_X1 U1017 ( .A1(G237), .A2(G234), .ZN(n1195) );
NOR2_X1 U1018 ( .A1(n1053), .A2(n1011), .ZN(n1001) );
AND2_X1 U1019 ( .A1(G221), .A2(n1203), .ZN(n1011) );
NAND2_X1 U1020 ( .A1(G234), .A2(n1204), .ZN(n1203) );
XOR2_X1 U1021 ( .A(n1016), .B(n1286), .Z(n1053) );
NOR2_X1 U1022 ( .A1(KEYINPUT4), .A2(n1287), .ZN(n1286) );
INV_X1 U1023 ( .A(G469), .ZN(n1287) );
NAND2_X1 U1024 ( .A1(n1288), .A2(n1204), .ZN(n1016) );
INV_X1 U1025 ( .A(G902), .ZN(n1204) );
XOR2_X1 U1026 ( .A(n1289), .B(n1290), .Z(n1288) );
INV_X1 U1027 ( .A(n1133), .ZN(n1290) );
XOR2_X1 U1028 ( .A(n1274), .B(n1291), .Z(n1133) );
XOR2_X1 U1029 ( .A(G101), .B(n1068), .Z(n1291) );
XNOR2_X1 U1030 ( .A(n1292), .B(n1293), .ZN(n1068) );
NOR2_X1 U1031 ( .A1(KEYINPUT54), .A2(n1294), .ZN(n1293) );
XOR2_X1 U1032 ( .A(G146), .B(G143), .Z(n1294) );
XNOR2_X1 U1033 ( .A(G128), .B(KEYINPUT24), .ZN(n1292) );
XNOR2_X1 U1034 ( .A(G104), .B(G107), .ZN(n1274) );
XNOR2_X1 U1035 ( .A(n1134), .B(n1137), .ZN(n1289) );
XNOR2_X1 U1036 ( .A(n1211), .B(n1295), .ZN(n1137) );
XOR2_X1 U1037 ( .A(G140), .B(n1296), .Z(n1295) );
NOR2_X1 U1038 ( .A1(G953), .A2(n1078), .ZN(n1296) );
INV_X1 U1039 ( .A(G227), .ZN(n1078) );
XNOR2_X1 U1040 ( .A(G110), .B(KEYINPUT32), .ZN(n1211) );
AND2_X1 U1041 ( .A1(n1297), .A2(n1298), .ZN(n1134) );
NAND2_X1 U1042 ( .A1(G131), .A2(n1299), .ZN(n1298) );
XOR2_X1 U1043 ( .A(G137), .B(G134), .Z(n1299) );
XOR2_X1 U1044 ( .A(n1300), .B(KEYINPUT55), .Z(n1297) );
NAND2_X1 U1045 ( .A1(n1301), .A2(n1077), .ZN(n1300) );
INV_X1 U1046 ( .A(G131), .ZN(n1077) );
XOR2_X1 U1047 ( .A(n1184), .B(G137), .Z(n1301) );
INV_X1 U1048 ( .A(G134), .ZN(n1184) );
endmodule


