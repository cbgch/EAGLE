//Key = 0001110110100011001110101101001101000010010100100111010011110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402;

XOR2_X1 U763 ( .A(G107), .B(n1061), .Z(G9) );
NOR2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(G75) );
NOR3_X1 U765 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
INV_X1 U766 ( .A(n1067), .ZN(n1066) );
NOR2_X1 U767 ( .A1(n1068), .A2(n1069), .ZN(n1065) );
NOR2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
INV_X1 U770 ( .A(KEYINPUT28), .ZN(n1073) );
NOR4_X1 U771 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1072) );
NOR2_X1 U772 ( .A1(n1078), .A2(n1077), .ZN(n1070) );
NOR2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
AND2_X1 U774 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U775 ( .A1(n1083), .A2(n1076), .ZN(n1079) );
NOR2_X1 U776 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U777 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
INV_X1 U778 ( .A(n1088), .ZN(n1087) );
NOR2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NOR3_X1 U780 ( .A1(n1075), .A2(KEYINPUT28), .A3(n1074), .ZN(n1084) );
INV_X1 U781 ( .A(n1081), .ZN(n1074) );
NAND3_X1 U782 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1064) );
NAND3_X1 U783 ( .A1(n1081), .A2(n1094), .A3(n1095), .ZN(n1093) );
INV_X1 U784 ( .A(n1077), .ZN(n1095) );
NAND2_X1 U785 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NAND3_X1 U786 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1097) );
NAND2_X1 U787 ( .A1(n1088), .A2(n1101), .ZN(n1096) );
NAND2_X1 U788 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND4_X1 U789 ( .A1(n1104), .A2(n1100), .A3(n1105), .A4(n1106), .ZN(n1103) );
INV_X1 U790 ( .A(KEYINPUT44), .ZN(n1106) );
NAND2_X1 U791 ( .A1(n1098), .A2(n1107), .ZN(n1102) );
NAND3_X1 U792 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1107) );
NAND2_X1 U793 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U794 ( .A1(KEYINPUT44), .A2(n1100), .ZN(n1108) );
NOR3_X1 U795 ( .A1(n1113), .A2(G953), .A3(G952), .ZN(n1062) );
INV_X1 U796 ( .A(n1091), .ZN(n1113) );
NAND4_X1 U797 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1091) );
NOR4_X1 U798 ( .A1(n1112), .A2(n1104), .A3(n1118), .A4(n1119), .ZN(n1117) );
XNOR2_X1 U799 ( .A(n1120), .B(n1121), .ZN(n1119) );
NOR2_X1 U800 ( .A1(G478), .A2(n1122), .ZN(n1121) );
XNOR2_X1 U801 ( .A(KEYINPUT40), .B(KEYINPUT33), .ZN(n1122) );
XOR2_X1 U802 ( .A(n1123), .B(n1124), .Z(n1118) );
XNOR2_X1 U803 ( .A(KEYINPUT18), .B(n1125), .ZN(n1124) );
NOR2_X1 U804 ( .A1(n1126), .A2(n1127), .ZN(n1116) );
XOR2_X1 U805 ( .A(n1128), .B(n1129), .Z(n1115) );
XOR2_X1 U806 ( .A(KEYINPUT37), .B(n1130), .Z(n1129) );
NAND2_X1 U807 ( .A1(KEYINPUT5), .A2(n1131), .ZN(n1128) );
XOR2_X1 U808 ( .A(n1132), .B(n1133), .Z(n1114) );
NOR2_X1 U809 ( .A1(KEYINPUT16), .A2(n1134), .ZN(n1133) );
NAND2_X1 U810 ( .A1(n1135), .A2(n1136), .ZN(G72) );
NAND2_X1 U811 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U812 ( .A(n1139), .B(n1140), .Z(n1135) );
XOR2_X1 U813 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U814 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U815 ( .A(n1145), .B(n1146), .Z(n1144) );
XNOR2_X1 U816 ( .A(n1147), .B(n1148), .ZN(n1146) );
XNOR2_X1 U817 ( .A(n1149), .B(n1150), .ZN(n1145) );
XOR2_X1 U818 ( .A(KEYINPUT38), .B(n1151), .Z(n1150) );
NOR2_X1 U819 ( .A1(G131), .A2(KEYINPUT23), .ZN(n1151) );
NOR2_X1 U820 ( .A1(G900), .A2(n1092), .ZN(n1143) );
NOR2_X1 U821 ( .A1(n1152), .A2(n1153), .ZN(n1141) );
XNOR2_X1 U822 ( .A(G953), .B(KEYINPUT58), .ZN(n1153) );
NOR2_X1 U823 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
XOR2_X1 U824 ( .A(KEYINPUT52), .B(n1156), .Z(n1155) );
OR2_X1 U825 ( .A1(n1138), .A2(n1137), .ZN(n1139) );
NAND2_X1 U826 ( .A1(G953), .A2(n1157), .ZN(n1137) );
NAND2_X1 U827 ( .A1(G900), .A2(G227), .ZN(n1157) );
INV_X1 U828 ( .A(KEYINPUT15), .ZN(n1138) );
XOR2_X1 U829 ( .A(n1158), .B(n1159), .Z(G69) );
XOR2_X1 U830 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U831 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U832 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U833 ( .A1(KEYINPUT8), .A2(n1166), .ZN(n1164) );
NOR2_X1 U834 ( .A1(n1092), .A2(n1167), .ZN(n1162) );
XNOR2_X1 U835 ( .A(KEYINPUT2), .B(n1168), .ZN(n1167) );
NAND2_X1 U836 ( .A1(n1092), .A2(n1169), .ZN(n1160) );
NAND2_X1 U837 ( .A1(G953), .A2(n1170), .ZN(n1158) );
NAND2_X1 U838 ( .A1(G898), .A2(G224), .ZN(n1170) );
NOR2_X1 U839 ( .A1(n1171), .A2(n1172), .ZN(G66) );
NOR3_X1 U840 ( .A1(n1130), .A2(n1173), .A3(n1174), .ZN(n1172) );
AND3_X1 U841 ( .A1(n1175), .A2(n1131), .A3(n1176), .ZN(n1174) );
INV_X1 U842 ( .A(n1177), .ZN(n1131) );
NOR2_X1 U843 ( .A1(n1178), .A2(n1175), .ZN(n1173) );
NOR2_X1 U844 ( .A1(n1067), .A2(n1177), .ZN(n1178) );
NOR2_X1 U845 ( .A1(n1171), .A2(n1179), .ZN(G63) );
NOR3_X1 U846 ( .A1(n1120), .A2(n1180), .A3(n1181), .ZN(n1179) );
NOR4_X1 U847 ( .A1(n1182), .A2(n1183), .A3(KEYINPUT17), .A4(n1184), .ZN(n1181) );
NOR2_X1 U848 ( .A1(n1185), .A2(n1186), .ZN(n1180) );
NOR3_X1 U849 ( .A1(n1184), .A2(KEYINPUT17), .A3(n1067), .ZN(n1185) );
NOR2_X1 U850 ( .A1(n1171), .A2(n1187), .ZN(G60) );
XOR2_X1 U851 ( .A(n1188), .B(n1189), .Z(n1187) );
NAND2_X1 U852 ( .A1(n1176), .A2(G475), .ZN(n1188) );
XOR2_X1 U853 ( .A(G104), .B(n1190), .Z(G6) );
NOR2_X1 U854 ( .A1(n1171), .A2(n1191), .ZN(G57) );
XOR2_X1 U855 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U856 ( .A(n1194), .B(n1195), .Z(n1193) );
AND2_X1 U857 ( .A1(G472), .A2(n1176), .ZN(n1195) );
NOR2_X1 U858 ( .A1(KEYINPUT29), .A2(n1196), .ZN(n1194) );
XNOR2_X1 U859 ( .A(n1197), .B(n1198), .ZN(n1196) );
XNOR2_X1 U860 ( .A(n1199), .B(n1200), .ZN(n1198) );
NOR2_X1 U861 ( .A1(KEYINPUT26), .A2(n1201), .ZN(n1199) );
NAND2_X1 U862 ( .A1(KEYINPUT7), .A2(n1202), .ZN(n1192) );
NOR2_X1 U863 ( .A1(n1171), .A2(n1203), .ZN(G54) );
XOR2_X1 U864 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U865 ( .A(n1206), .B(n1207), .Z(n1205) );
NAND3_X1 U866 ( .A1(KEYINPUT53), .A2(n1208), .A3(n1209), .ZN(n1207) );
XOR2_X1 U867 ( .A(n1210), .B(KEYINPUT55), .Z(n1209) );
NAND2_X1 U868 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
OR2_X1 U869 ( .A1(n1212), .A2(n1211), .ZN(n1208) );
XNOR2_X1 U870 ( .A(n1213), .B(KEYINPUT6), .ZN(n1212) );
NAND2_X1 U871 ( .A1(n1214), .A2(n1215), .ZN(n1206) );
NAND3_X1 U872 ( .A1(n1216), .A2(n1217), .A3(n1201), .ZN(n1215) );
NAND2_X1 U873 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
XNOR2_X1 U874 ( .A(KEYINPUT32), .B(n1220), .ZN(n1218) );
NAND2_X1 U875 ( .A1(n1221), .A2(n1222), .ZN(n1214) );
XNOR2_X1 U876 ( .A(n1223), .B(n1220), .ZN(n1222) );
OR2_X1 U877 ( .A1(n1147), .A2(KEYINPUT32), .ZN(n1223) );
XNOR2_X1 U878 ( .A(n1201), .B(KEYINPUT0), .ZN(n1221) );
NOR2_X1 U879 ( .A1(n1125), .A2(n1183), .ZN(n1204) );
NOR2_X1 U880 ( .A1(n1171), .A2(n1224), .ZN(G51) );
NOR2_X1 U881 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U882 ( .A(KEYINPUT61), .B(n1227), .Z(n1226) );
NOR2_X1 U883 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
AND2_X1 U884 ( .A1(n1229), .A2(n1228), .ZN(n1225) );
XOR2_X1 U885 ( .A(n1230), .B(n1231), .Z(n1228) );
XNOR2_X1 U886 ( .A(n1232), .B(n1233), .ZN(n1231) );
NAND3_X1 U887 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
INV_X1 U888 ( .A(n1237), .ZN(n1236) );
OR2_X1 U889 ( .A1(n1238), .A2(KEYINPUT46), .ZN(n1235) );
NAND2_X1 U890 ( .A1(n1239), .A2(KEYINPUT46), .ZN(n1234) );
OR2_X1 U891 ( .A1(n1183), .A2(n1132), .ZN(n1229) );
INV_X1 U892 ( .A(n1176), .ZN(n1183) );
NOR2_X1 U893 ( .A1(n1240), .A2(n1067), .ZN(n1176) );
NOR3_X1 U894 ( .A1(n1154), .A2(n1156), .A3(n1169), .ZN(n1067) );
NAND4_X1 U895 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1169) );
NOR4_X1 U896 ( .A1(n1061), .A2(n1245), .A3(n1246), .A4(n1190), .ZN(n1244) );
AND2_X1 U897 ( .A1(n1247), .A2(n1248), .ZN(n1190) );
INV_X1 U898 ( .A(n1249), .ZN(n1246) );
AND2_X1 U899 ( .A1(n1248), .A2(n1099), .ZN(n1061) );
AND3_X1 U900 ( .A1(n1081), .A2(n1250), .A3(n1251), .ZN(n1248) );
NAND2_X1 U901 ( .A1(KEYINPUT25), .A2(n1252), .ZN(n1243) );
NAND2_X1 U902 ( .A1(n1253), .A2(n1254), .ZN(n1242) );
NAND2_X1 U903 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
NAND2_X1 U904 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND2_X1 U905 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NAND3_X1 U906 ( .A1(n1089), .A2(n1261), .A3(n1082), .ZN(n1260) );
INV_X1 U907 ( .A(KEYINPUT25), .ZN(n1261) );
NAND2_X1 U908 ( .A1(KEYINPUT60), .A2(n1262), .ZN(n1259) );
NAND2_X1 U909 ( .A1(KEYINPUT42), .A2(n1263), .ZN(n1255) );
NAND3_X1 U910 ( .A1(n1082), .A2(n1264), .A3(n1090), .ZN(n1263) );
NAND2_X1 U911 ( .A1(n1250), .A2(n1265), .ZN(n1241) );
NAND3_X1 U912 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(n1265) );
NAND2_X1 U913 ( .A1(n1262), .A2(n1269), .ZN(n1268) );
INV_X1 U914 ( .A(KEYINPUT60), .ZN(n1269) );
NAND3_X1 U915 ( .A1(n1082), .A2(n1270), .A3(n1090), .ZN(n1267) );
INV_X1 U916 ( .A(KEYINPUT42), .ZN(n1270) );
NAND2_X1 U917 ( .A1(n1271), .A2(n1272), .ZN(n1266) );
XNOR2_X1 U918 ( .A(n1098), .B(KEYINPUT24), .ZN(n1271) );
NAND4_X1 U919 ( .A1(n1273), .A2(n1274), .A3(n1275), .A4(n1276), .ZN(n1154) );
NOR4_X1 U920 ( .A1(n1277), .A2(n1278), .A3(n1279), .A4(n1280), .ZN(n1276) );
NOR2_X1 U921 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NOR2_X1 U922 ( .A1(n1076), .A2(n1283), .ZN(n1279) );
NOR3_X1 U923 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1278) );
NAND3_X1 U924 ( .A1(n1251), .A2(n1287), .A3(n1089), .ZN(n1286) );
NAND3_X1 U925 ( .A1(n1288), .A2(n1109), .A3(n1289), .ZN(n1285) );
INV_X1 U926 ( .A(KEYINPUT13), .ZN(n1284) );
NOR2_X1 U927 ( .A1(KEYINPUT13), .A2(n1290), .ZN(n1277) );
NOR2_X1 U928 ( .A1(n1291), .A2(n1292), .ZN(n1275) );
INV_X1 U929 ( .A(n1293), .ZN(n1292) );
NOR2_X1 U930 ( .A1(n1092), .A2(G952), .ZN(n1171) );
XOR2_X1 U931 ( .A(G146), .B(n1156), .Z(G48) );
AND2_X1 U932 ( .A1(n1247), .A2(n1294), .ZN(n1156) );
XNOR2_X1 U933 ( .A(G143), .B(n1290), .ZN(G45) );
NAND4_X1 U934 ( .A1(n1089), .A2(n1295), .A3(n1289), .A4(n1287), .ZN(n1290) );
NAND2_X1 U935 ( .A1(n1296), .A2(n1297), .ZN(G42) );
NAND2_X1 U936 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
XOR2_X1 U937 ( .A(n1273), .B(KEYINPUT31), .Z(n1298) );
NAND2_X1 U938 ( .A1(n1300), .A2(G140), .ZN(n1296) );
XOR2_X1 U939 ( .A(n1273), .B(KEYINPUT48), .Z(n1300) );
NAND3_X1 U940 ( .A1(n1090), .A2(n1247), .A3(n1301), .ZN(n1273) );
XNOR2_X1 U941 ( .A(G137), .B(n1302), .ZN(G39) );
NAND2_X1 U942 ( .A1(KEYINPUT57), .A2(n1303), .ZN(n1302) );
INV_X1 U943 ( .A(n1274), .ZN(n1303) );
NAND4_X1 U944 ( .A1(n1301), .A2(n1088), .A3(n1304), .A4(n1127), .ZN(n1274) );
XNOR2_X1 U945 ( .A(G134), .B(n1305), .ZN(G36) );
NAND4_X1 U946 ( .A1(n1306), .A2(n1100), .A3(n1272), .A4(n1288), .ZN(n1305) );
INV_X1 U947 ( .A(n1281), .ZN(n1272) );
XNOR2_X1 U948 ( .A(n1251), .B(KEYINPUT51), .ZN(n1306) );
NAND2_X1 U949 ( .A1(n1307), .A2(n1308), .ZN(G33) );
OR2_X1 U950 ( .A1(n1293), .A2(G131), .ZN(n1308) );
XOR2_X1 U951 ( .A(n1309), .B(KEYINPUT1), .Z(n1307) );
NAND2_X1 U952 ( .A1(G131), .A2(n1293), .ZN(n1309) );
NAND3_X1 U953 ( .A1(n1089), .A2(n1247), .A3(n1301), .ZN(n1293) );
INV_X1 U954 ( .A(n1282), .ZN(n1301) );
NAND3_X1 U955 ( .A1(n1251), .A2(n1288), .A3(n1100), .ZN(n1282) );
INV_X1 U956 ( .A(n1069), .ZN(n1100) );
NAND2_X1 U957 ( .A1(n1111), .A2(n1310), .ZN(n1069) );
XOR2_X1 U958 ( .A(KEYINPUT20), .B(n1112), .Z(n1310) );
XOR2_X1 U959 ( .A(G128), .B(n1291), .Z(G30) );
AND2_X1 U960 ( .A1(n1294), .A2(n1099), .ZN(n1291) );
AND3_X1 U961 ( .A1(n1304), .A2(n1127), .A3(n1295), .ZN(n1294) );
AND3_X1 U962 ( .A1(n1253), .A2(n1288), .A3(n1251), .ZN(n1295) );
XOR2_X1 U963 ( .A(n1311), .B(n1252), .Z(G3) );
AND3_X1 U964 ( .A1(n1089), .A2(n1250), .A3(n1082), .ZN(n1252) );
AND2_X1 U965 ( .A1(n1088), .A2(n1251), .ZN(n1082) );
NAND2_X1 U966 ( .A1(KEYINPUT43), .A2(n1312), .ZN(n1311) );
XOR2_X1 U967 ( .A(G125), .B(n1313), .Z(G27) );
NOR2_X1 U968 ( .A1(n1314), .A2(n1283), .ZN(n1313) );
NAND4_X1 U969 ( .A1(n1090), .A2(n1247), .A3(n1253), .A4(n1288), .ZN(n1283) );
NAND2_X1 U970 ( .A1(n1077), .A2(n1315), .ZN(n1288) );
NAND4_X1 U971 ( .A1(G953), .A2(G902), .A3(n1316), .A4(n1317), .ZN(n1315) );
INV_X1 U972 ( .A(G900), .ZN(n1317) );
XNOR2_X1 U973 ( .A(n1098), .B(KEYINPUT45), .ZN(n1314) );
XNOR2_X1 U974 ( .A(G122), .B(n1249), .ZN(G24) );
NAND4_X1 U975 ( .A1(n1289), .A2(n1318), .A3(n1081), .A4(n1287), .ZN(n1249) );
NOR2_X1 U976 ( .A1(n1319), .A2(n1304), .ZN(n1081) );
XNOR2_X1 U977 ( .A(KEYINPUT27), .B(n1127), .ZN(n1319) );
XNOR2_X1 U978 ( .A(G119), .B(n1320), .ZN(G21) );
NAND3_X1 U979 ( .A1(n1262), .A2(n1250), .A3(KEYINPUT19), .ZN(n1320) );
AND4_X1 U980 ( .A1(n1088), .A2(n1098), .A3(n1304), .A4(n1127), .ZN(n1262) );
XOR2_X1 U981 ( .A(G116), .B(n1321), .Z(G18) );
NOR2_X1 U982 ( .A1(n1322), .A2(n1281), .ZN(n1321) );
NAND2_X1 U983 ( .A1(n1089), .A2(n1099), .ZN(n1281) );
NOR2_X1 U984 ( .A1(n1126), .A2(n1323), .ZN(n1099) );
XOR2_X1 U985 ( .A(G113), .B(n1245), .Z(G15) );
AND3_X1 U986 ( .A1(n1318), .A2(n1247), .A3(n1089), .ZN(n1245) );
AND2_X1 U987 ( .A1(n1324), .A2(n1127), .ZN(n1089) );
XNOR2_X1 U988 ( .A(KEYINPUT21), .B(n1304), .ZN(n1324) );
INV_X1 U989 ( .A(n1075), .ZN(n1247) );
NAND2_X1 U990 ( .A1(n1323), .A2(n1289), .ZN(n1075) );
XNOR2_X1 U991 ( .A(n1126), .B(KEYINPUT41), .ZN(n1289) );
INV_X1 U992 ( .A(n1322), .ZN(n1318) );
NAND2_X1 U993 ( .A1(n1098), .A2(n1250), .ZN(n1322) );
INV_X1 U994 ( .A(n1076), .ZN(n1098) );
NAND2_X1 U995 ( .A1(n1105), .A2(n1325), .ZN(n1076) );
XNOR2_X1 U996 ( .A(G110), .B(n1326), .ZN(G12) );
NAND4_X1 U997 ( .A1(n1327), .A2(n1090), .A3(n1088), .A4(n1250), .ZN(n1326) );
NOR2_X1 U998 ( .A1(n1109), .A2(n1257), .ZN(n1250) );
INV_X1 U999 ( .A(n1264), .ZN(n1257) );
NAND2_X1 U1000 ( .A1(n1077), .A2(n1328), .ZN(n1264) );
NAND4_X1 U1001 ( .A1(G953), .A2(G902), .A3(n1316), .A4(n1168), .ZN(n1328) );
INV_X1 U1002 ( .A(G898), .ZN(n1168) );
NAND3_X1 U1003 ( .A1(n1316), .A2(n1092), .A3(G952), .ZN(n1077) );
NAND2_X1 U1004 ( .A1(G237), .A2(G234), .ZN(n1316) );
INV_X1 U1005 ( .A(n1253), .ZN(n1109) );
NOR2_X1 U1006 ( .A1(n1111), .A2(n1112), .ZN(n1253) );
AND2_X1 U1007 ( .A1(G214), .A2(n1329), .ZN(n1112) );
XNOR2_X1 U1008 ( .A(n1134), .B(n1132), .ZN(n1111) );
NAND2_X1 U1009 ( .A1(G210), .A2(n1329), .ZN(n1132) );
NAND2_X1 U1010 ( .A1(n1240), .A2(n1330), .ZN(n1329) );
NAND2_X1 U1011 ( .A1(n1331), .A2(n1240), .ZN(n1134) );
XNOR2_X1 U1012 ( .A(n1332), .B(n1333), .ZN(n1331) );
INV_X1 U1013 ( .A(n1230), .ZN(n1333) );
XOR2_X1 U1014 ( .A(n1166), .B(n1165), .Z(n1230) );
XNOR2_X1 U1015 ( .A(n1334), .B(G122), .ZN(n1165) );
XOR2_X1 U1016 ( .A(n1335), .B(n1336), .Z(n1166) );
NOR3_X1 U1017 ( .A1(KEYINPUT39), .A2(n1337), .A3(n1338), .ZN(n1332) );
NOR3_X1 U1018 ( .A1(n1339), .A2(n1239), .A3(n1237), .ZN(n1338) );
NOR2_X1 U1019 ( .A1(n1232), .A2(n1340), .ZN(n1337) );
NOR2_X1 U1020 ( .A1(n1239), .A2(n1237), .ZN(n1340) );
NOR2_X1 U1021 ( .A1(n1341), .A2(n1238), .ZN(n1237) );
NOR2_X1 U1022 ( .A1(n1200), .A2(n1342), .ZN(n1239) );
INV_X1 U1023 ( .A(n1339), .ZN(n1232) );
NAND2_X1 U1024 ( .A1(G224), .A2(n1092), .ZN(n1339) );
NOR2_X1 U1025 ( .A1(n1287), .A2(n1126), .ZN(n1088) );
XNOR2_X1 U1026 ( .A(n1343), .B(G475), .ZN(n1126) );
NAND2_X1 U1027 ( .A1(n1189), .A2(n1240), .ZN(n1343) );
XNOR2_X1 U1028 ( .A(n1344), .B(n1345), .ZN(n1189) );
XOR2_X1 U1029 ( .A(n1149), .B(n1346), .Z(n1345) );
XOR2_X1 U1030 ( .A(G104), .B(n1347), .Z(n1346) );
NOR3_X1 U1031 ( .A1(KEYINPUT9), .A2(n1348), .A3(n1349), .ZN(n1347) );
NOR2_X1 U1032 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
XNOR2_X1 U1033 ( .A(KEYINPUT10), .B(n1352), .ZN(n1350) );
AND2_X1 U1034 ( .A1(n1352), .A2(n1351), .ZN(n1348) );
NAND3_X1 U1035 ( .A1(n1330), .A2(n1092), .A3(G214), .ZN(n1351) );
XOR2_X1 U1036 ( .A(G140), .B(n1341), .Z(n1149) );
XOR2_X1 U1037 ( .A(n1353), .B(n1354), .Z(n1344) );
XOR2_X1 U1038 ( .A(G146), .B(G131), .Z(n1354) );
XNOR2_X1 U1039 ( .A(G113), .B(G122), .ZN(n1353) );
INV_X1 U1040 ( .A(n1323), .ZN(n1287) );
XOR2_X1 U1041 ( .A(n1120), .B(n1184), .Z(n1323) );
INV_X1 U1042 ( .A(G478), .ZN(n1184) );
NOR2_X1 U1043 ( .A1(n1186), .A2(G902), .ZN(n1120) );
INV_X1 U1044 ( .A(n1182), .ZN(n1186) );
XNOR2_X1 U1045 ( .A(n1355), .B(n1356), .ZN(n1182) );
XOR2_X1 U1046 ( .A(n1357), .B(n1358), .Z(n1356) );
XOR2_X1 U1047 ( .A(G116), .B(G107), .Z(n1358) );
AND3_X1 U1048 ( .A1(G217), .A2(n1092), .A3(G234), .ZN(n1357) );
XOR2_X1 U1049 ( .A(n1359), .B(n1360), .Z(n1355) );
XNOR2_X1 U1050 ( .A(G128), .B(n1361), .ZN(n1360) );
INV_X1 U1051 ( .A(G122), .ZN(n1361) );
XNOR2_X1 U1052 ( .A(G134), .B(G143), .ZN(n1359) );
AND2_X1 U1053 ( .A1(n1304), .A2(n1362), .ZN(n1090) );
XOR2_X1 U1054 ( .A(KEYINPUT27), .B(n1127), .Z(n1362) );
XNOR2_X1 U1055 ( .A(n1363), .B(G472), .ZN(n1127) );
NAND2_X1 U1056 ( .A1(n1364), .A2(n1240), .ZN(n1363) );
XOR2_X1 U1057 ( .A(n1365), .B(n1366), .Z(n1364) );
XNOR2_X1 U1058 ( .A(n1202), .B(n1201), .ZN(n1366) );
XOR2_X1 U1059 ( .A(n1312), .B(n1367), .Z(n1202) );
AND3_X1 U1060 ( .A1(G210), .A2(n1092), .A3(n1330), .ZN(n1367) );
INV_X1 U1061 ( .A(G237), .ZN(n1330) );
INV_X1 U1062 ( .A(G101), .ZN(n1312) );
XNOR2_X1 U1063 ( .A(n1368), .B(n1369), .ZN(n1365) );
INV_X1 U1064 ( .A(n1197), .ZN(n1369) );
XNOR2_X1 U1065 ( .A(n1335), .B(n1370), .ZN(n1197) );
XOR2_X1 U1066 ( .A(KEYINPUT59), .B(KEYINPUT22), .Z(n1370) );
XNOR2_X1 U1067 ( .A(G113), .B(n1371), .ZN(n1335) );
XOR2_X1 U1068 ( .A(G119), .B(G116), .Z(n1371) );
NOR2_X1 U1069 ( .A1(KEYINPUT54), .A2(n1200), .ZN(n1368) );
INV_X1 U1070 ( .A(n1238), .ZN(n1200) );
XOR2_X1 U1071 ( .A(G128), .B(n1372), .Z(n1238) );
NOR2_X1 U1072 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
AND2_X1 U1073 ( .A1(KEYINPUT34), .A2(n1375), .ZN(n1374) );
NOR2_X1 U1074 ( .A1(KEYINPUT36), .A2(n1375), .ZN(n1373) );
XOR2_X1 U1075 ( .A(n1376), .B(n1130), .Z(n1304) );
NOR2_X1 U1076 ( .A1(n1175), .A2(G902), .ZN(n1130) );
XNOR2_X1 U1077 ( .A(n1377), .B(n1378), .ZN(n1175) );
XOR2_X1 U1078 ( .A(n1379), .B(n1380), .Z(n1378) );
XNOR2_X1 U1079 ( .A(G110), .B(n1381), .ZN(n1380) );
AND3_X1 U1080 ( .A1(G221), .A2(n1092), .A3(G234), .ZN(n1381) );
NAND2_X1 U1081 ( .A1(KEYINPUT3), .A2(n1382), .ZN(n1379) );
XNOR2_X1 U1082 ( .A(n1342), .B(n1383), .ZN(n1382) );
XNOR2_X1 U1083 ( .A(G146), .B(n1384), .ZN(n1383) );
NAND2_X1 U1084 ( .A1(KEYINPUT63), .A2(G140), .ZN(n1384) );
INV_X1 U1085 ( .A(n1341), .ZN(n1342) );
XOR2_X1 U1086 ( .A(G125), .B(KEYINPUT11), .Z(n1341) );
XOR2_X1 U1087 ( .A(n1385), .B(n1386), .Z(n1377) );
XOR2_X1 U1088 ( .A(KEYINPUT62), .B(G137), .Z(n1386) );
XNOR2_X1 U1089 ( .A(G119), .B(G128), .ZN(n1385) );
NAND2_X1 U1090 ( .A1(KEYINPUT4), .A2(n1177), .ZN(n1376) );
NAND2_X1 U1091 ( .A1(G217), .A2(n1387), .ZN(n1177) );
XNOR2_X1 U1092 ( .A(n1251), .B(KEYINPUT56), .ZN(n1327) );
NOR2_X1 U1093 ( .A1(n1105), .A2(n1104), .ZN(n1251) );
INV_X1 U1094 ( .A(n1325), .ZN(n1104) );
NAND2_X1 U1095 ( .A1(G221), .A2(n1387), .ZN(n1325) );
NAND2_X1 U1096 ( .A1(n1388), .A2(n1240), .ZN(n1387) );
XNOR2_X1 U1097 ( .A(G234), .B(KEYINPUT30), .ZN(n1388) );
XOR2_X1 U1098 ( .A(n1389), .B(n1123), .Z(n1105) );
NAND2_X1 U1099 ( .A1(n1390), .A2(n1240), .ZN(n1123) );
INV_X1 U1100 ( .A(G902), .ZN(n1240) );
XOR2_X1 U1101 ( .A(n1391), .B(n1392), .Z(n1390) );
XNOR2_X1 U1102 ( .A(n1213), .B(n1201), .ZN(n1392) );
XOR2_X1 U1103 ( .A(n1148), .B(n1393), .Z(n1201) );
NOR2_X1 U1104 ( .A1(G131), .A2(KEYINPUT35), .ZN(n1393) );
XOR2_X1 U1105 ( .A(G134), .B(G137), .Z(n1148) );
NAND2_X1 U1106 ( .A1(G227), .A2(n1092), .ZN(n1213) );
INV_X1 U1107 ( .A(G953), .ZN(n1092) );
XNOR2_X1 U1108 ( .A(n1394), .B(n1395), .ZN(n1391) );
NOR2_X1 U1109 ( .A1(KEYINPUT47), .A2(n1211), .ZN(n1395) );
XNOR2_X1 U1110 ( .A(n1334), .B(n1299), .ZN(n1211) );
INV_X1 U1111 ( .A(G140), .ZN(n1299) );
INV_X1 U1112 ( .A(G110), .ZN(n1334) );
NAND3_X1 U1113 ( .A1(n1396), .A2(n1217), .A3(KEYINPUT14), .ZN(n1394) );
NAND2_X1 U1114 ( .A1(n1147), .A2(n1220), .ZN(n1217) );
NAND2_X1 U1115 ( .A1(n1336), .A2(n1219), .ZN(n1396) );
INV_X1 U1116 ( .A(n1147), .ZN(n1219) );
XOR2_X1 U1117 ( .A(G128), .B(n1397), .Z(n1147) );
NOR2_X1 U1118 ( .A1(n1398), .A2(n1399), .ZN(n1397) );
NOR3_X1 U1119 ( .A1(n1400), .A2(G146), .A3(n1352), .ZN(n1399) );
AND2_X1 U1120 ( .A1(n1400), .A2(n1375), .ZN(n1398) );
XOR2_X1 U1121 ( .A(G146), .B(n1352), .Z(n1375) );
INV_X1 U1122 ( .A(G143), .ZN(n1352) );
INV_X1 U1123 ( .A(KEYINPUT12), .ZN(n1400) );
INV_X1 U1124 ( .A(n1220), .ZN(n1336) );
XNOR2_X1 U1125 ( .A(n1401), .B(n1402), .ZN(n1220) );
XOR2_X1 U1126 ( .A(KEYINPUT50), .B(G107), .Z(n1402) );
XNOR2_X1 U1127 ( .A(G101), .B(G104), .ZN(n1401) );
NAND2_X1 U1128 ( .A1(KEYINPUT49), .A2(n1125), .ZN(n1389) );
INV_X1 U1129 ( .A(G469), .ZN(n1125) );
endmodule


