//Key = 1111011000100010000000110111010010001111011100010001011011000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382;

XOR2_X1 U768 ( .A(n1051), .B(n1052), .Z(G9) );
XNOR2_X1 U769 ( .A(G107), .B(KEYINPUT51), .ZN(n1051) );
NOR2_X1 U770 ( .A1(n1053), .A2(n1054), .ZN(G75) );
NOR3_X1 U771 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NAND3_X1 U772 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1055) );
NAND2_X1 U773 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U774 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U775 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NAND2_X1 U776 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NAND2_X1 U777 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
OR2_X1 U778 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U779 ( .A1(n1074), .A2(n1075), .ZN(n1068) );
NAND2_X1 U780 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND3_X1 U781 ( .A1(n1070), .A2(n1078), .A3(n1074), .ZN(n1063) );
NAND2_X1 U782 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U783 ( .A1(n1067), .A2(n1081), .ZN(n1080) );
NAND2_X1 U784 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U785 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U786 ( .A1(n1065), .A2(n1086), .ZN(n1079) );
NAND2_X1 U787 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U788 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
INV_X1 U789 ( .A(n1091), .ZN(n1061) );
NOR3_X1 U790 ( .A1(n1092), .A2(G953), .A3(G952), .ZN(n1053) );
INV_X1 U791 ( .A(n1058), .ZN(n1092) );
NAND4_X1 U792 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1058) );
NOR4_X1 U793 ( .A1(n1084), .A2(n1097), .A3(n1089), .A4(n1098), .ZN(n1096) );
NOR2_X1 U794 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
INV_X1 U795 ( .A(n1101), .ZN(n1097) );
NOR2_X1 U796 ( .A1(n1102), .A2(n1103), .ZN(n1095) );
XOR2_X1 U797 ( .A(G478), .B(n1104), .Z(n1103) );
XNOR2_X1 U798 ( .A(n1105), .B(G469), .ZN(n1094) );
XNOR2_X1 U799 ( .A(n1106), .B(n1107), .ZN(n1093) );
XOR2_X1 U800 ( .A(n1108), .B(n1109), .Z(G72) );
NOR2_X1 U801 ( .A1(n1110), .A2(n1059), .ZN(n1109) );
AND2_X1 U802 ( .A1(G227), .A2(G900), .ZN(n1110) );
NAND2_X1 U803 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
NAND2_X1 U804 ( .A1(n1113), .A2(n1059), .ZN(n1112) );
XOR2_X1 U805 ( .A(n1056), .B(n1114), .Z(n1113) );
NAND3_X1 U806 ( .A1(G900), .A2(n1114), .A3(G953), .ZN(n1111) );
XNOR2_X1 U807 ( .A(n1115), .B(n1116), .ZN(n1114) );
XOR2_X1 U808 ( .A(n1117), .B(n1118), .Z(n1115) );
NOR2_X1 U809 ( .A1(KEYINPUT9), .A2(n1119), .ZN(n1118) );
NAND3_X1 U810 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1117) );
OR2_X1 U811 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U812 ( .A1(KEYINPUT12), .A2(n1125), .ZN(n1121) );
NAND2_X1 U813 ( .A1(n1126), .A2(n1124), .ZN(n1125) );
XNOR2_X1 U814 ( .A(n1123), .B(KEYINPUT56), .ZN(n1126) );
NAND2_X1 U815 ( .A1(n1127), .A2(n1128), .ZN(n1120) );
INV_X1 U816 ( .A(KEYINPUT12), .ZN(n1128) );
NAND2_X1 U817 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
OR2_X1 U818 ( .A1(n1123), .A2(KEYINPUT56), .ZN(n1130) );
NAND3_X1 U819 ( .A1(n1123), .A2(n1124), .A3(KEYINPUT56), .ZN(n1129) );
XOR2_X1 U820 ( .A(n1131), .B(n1132), .Z(n1123) );
NAND2_X1 U821 ( .A1(KEYINPUT54), .A2(n1133), .ZN(n1131) );
XOR2_X1 U822 ( .A(n1134), .B(n1135), .Z(G69) );
NOR2_X1 U823 ( .A1(n1136), .A2(n1059), .ZN(n1135) );
NOR2_X1 U824 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR3_X1 U825 ( .A1(KEYINPUT13), .A2(n1139), .A3(n1140), .ZN(n1134) );
NOR2_X1 U826 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
INV_X1 U827 ( .A(n1143), .ZN(n1142) );
NOR2_X1 U828 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
NOR2_X1 U829 ( .A1(G898), .A2(n1059), .ZN(n1144) );
NOR2_X1 U830 ( .A1(n1145), .A2(n1143), .ZN(n1139) );
XNOR2_X1 U831 ( .A(n1146), .B(n1147), .ZN(n1143) );
XOR2_X1 U832 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U833 ( .A(n1150), .B(n1151), .Z(n1146) );
XNOR2_X1 U834 ( .A(KEYINPUT46), .B(n1152), .ZN(n1151) );
NOR2_X1 U835 ( .A1(G953), .A2(n1153), .ZN(n1145) );
INV_X1 U836 ( .A(n1057), .ZN(n1153) );
NOR2_X1 U837 ( .A1(n1154), .A2(n1155), .ZN(G66) );
NOR2_X1 U838 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U839 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND2_X1 U840 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U841 ( .A1(KEYINPUT22), .A2(n1162), .ZN(n1158) );
NOR2_X1 U842 ( .A1(KEYINPUT22), .A2(n1162), .ZN(n1156) );
NOR2_X1 U843 ( .A1(n1154), .A2(n1163), .ZN(G63) );
XOR2_X1 U844 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U845 ( .A1(n1160), .A2(G478), .ZN(n1164) );
NOR2_X1 U846 ( .A1(n1154), .A2(n1166), .ZN(G60) );
XOR2_X1 U847 ( .A(n1167), .B(n1168), .Z(n1166) );
NAND2_X1 U848 ( .A1(n1160), .A2(G475), .ZN(n1167) );
XNOR2_X1 U849 ( .A(n1169), .B(n1170), .ZN(G6) );
NOR2_X1 U850 ( .A1(n1154), .A2(n1171), .ZN(G57) );
XOR2_X1 U851 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U852 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U853 ( .A(n1176), .B(n1177), .ZN(n1175) );
NAND2_X1 U854 ( .A1(KEYINPUT63), .A2(n1178), .ZN(n1176) );
XOR2_X1 U855 ( .A(n1179), .B(n1180), .Z(n1172) );
XOR2_X1 U856 ( .A(n1181), .B(n1182), .Z(n1180) );
NAND2_X1 U857 ( .A1(KEYINPUT41), .A2(n1183), .ZN(n1181) );
NAND2_X1 U858 ( .A1(n1160), .A2(G472), .ZN(n1179) );
NOR2_X1 U859 ( .A1(n1154), .A2(n1184), .ZN(G54) );
XOR2_X1 U860 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U861 ( .A(n1183), .B(n1187), .Z(n1186) );
XNOR2_X1 U862 ( .A(n1119), .B(n1188), .ZN(n1187) );
XOR2_X1 U863 ( .A(n1189), .B(n1190), .Z(n1185) );
XNOR2_X1 U864 ( .A(n1152), .B(n1191), .ZN(n1190) );
NOR2_X1 U865 ( .A1(KEYINPUT55), .A2(n1192), .ZN(n1191) );
XOR2_X1 U866 ( .A(n1193), .B(n1194), .Z(n1189) );
AND2_X1 U867 ( .A1(G469), .A2(n1160), .ZN(n1194) );
INV_X1 U868 ( .A(n1195), .ZN(n1160) );
NAND2_X1 U869 ( .A1(KEYINPUT3), .A2(n1196), .ZN(n1193) );
NOR2_X1 U870 ( .A1(n1154), .A2(n1197), .ZN(G51) );
XOR2_X1 U871 ( .A(n1198), .B(n1199), .Z(n1197) );
XNOR2_X1 U872 ( .A(n1200), .B(n1116), .ZN(n1199) );
XNOR2_X1 U873 ( .A(G125), .B(n1188), .ZN(n1116) );
OR2_X1 U874 ( .A1(n1195), .A2(n1107), .ZN(n1200) );
NAND2_X1 U875 ( .A1(G902), .A2(n1201), .ZN(n1195) );
OR2_X1 U876 ( .A1(n1057), .A2(n1056), .ZN(n1201) );
NAND4_X1 U877 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1056) );
NOR3_X1 U878 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1205) );
NOR2_X1 U879 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NOR2_X1 U880 ( .A1(n1211), .A2(n1212), .ZN(n1206) );
NOR2_X1 U881 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
NOR2_X1 U882 ( .A1(n1215), .A2(n1216), .ZN(n1213) );
NOR2_X1 U883 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
NOR2_X1 U884 ( .A1(n1076), .A2(n1219), .ZN(n1218) );
NOR2_X1 U885 ( .A1(n1220), .A2(n1077), .ZN(n1217) );
XNOR2_X1 U886 ( .A(n1073), .B(KEYINPUT48), .ZN(n1220) );
NAND4_X1 U887 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1057) );
NOR4_X1 U888 ( .A1(n1225), .A2(n1226), .A3(n1170), .A4(n1052), .ZN(n1224) );
AND3_X1 U889 ( .A1(n1073), .A2(n1070), .A3(n1227), .ZN(n1052) );
AND3_X1 U890 ( .A1(n1227), .A2(n1070), .A3(n1072), .ZN(n1170) );
NOR2_X1 U891 ( .A1(n1228), .A2(n1229), .ZN(n1223) );
NOR2_X1 U892 ( .A1(n1087), .A2(n1230), .ZN(n1229) );
XNOR2_X1 U893 ( .A(KEYINPUT25), .B(n1231), .ZN(n1230) );
XOR2_X1 U894 ( .A(n1232), .B(n1233), .Z(n1198) );
NAND2_X1 U895 ( .A1(KEYINPUT43), .A2(n1234), .ZN(n1233) );
NOR2_X1 U896 ( .A1(n1059), .A2(G952), .ZN(n1154) );
XNOR2_X1 U897 ( .A(n1207), .B(n1235), .ZN(G48) );
NAND2_X1 U898 ( .A1(KEYINPUT61), .A2(G146), .ZN(n1235) );
AND3_X1 U899 ( .A1(n1072), .A2(n1236), .A3(n1237), .ZN(n1207) );
XNOR2_X1 U900 ( .A(G143), .B(n1204), .ZN(G45) );
NAND4_X1 U901 ( .A1(n1238), .A2(n1236), .A3(n1239), .A4(n1240), .ZN(n1204) );
XOR2_X1 U902 ( .A(n1241), .B(n1242), .Z(G42) );
NOR2_X1 U903 ( .A1(G140), .A2(KEYINPUT28), .ZN(n1242) );
NAND4_X1 U904 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1241) );
XNOR2_X1 U905 ( .A(KEYINPUT7), .B(n1212), .ZN(n1246) );
XNOR2_X1 U906 ( .A(KEYINPUT35), .B(n1219), .ZN(n1245) );
XNOR2_X1 U907 ( .A(G137), .B(n1202), .ZN(G39) );
NAND3_X1 U908 ( .A1(n1237), .A2(n1074), .A3(n1067), .ZN(n1202) );
NOR3_X1 U909 ( .A1(n1247), .A2(n1248), .A3(n1216), .ZN(n1237) );
XNOR2_X1 U910 ( .A(G134), .B(n1249), .ZN(G36) );
NAND3_X1 U911 ( .A1(n1067), .A2(n1073), .A3(n1238), .ZN(n1249) );
INV_X1 U912 ( .A(n1212), .ZN(n1067) );
XNOR2_X1 U913 ( .A(n1250), .B(n1251), .ZN(G33) );
NOR2_X1 U914 ( .A1(n1252), .A2(n1212), .ZN(n1251) );
NAND2_X1 U915 ( .A1(n1090), .A2(n1253), .ZN(n1212) );
XNOR2_X1 U916 ( .A(n1214), .B(KEYINPUT4), .ZN(n1252) );
AND2_X1 U917 ( .A1(n1238), .A2(n1072), .ZN(n1214) );
NOR2_X1 U918 ( .A1(n1216), .A2(n1077), .ZN(n1238) );
INV_X1 U919 ( .A(n1254), .ZN(n1077) );
INV_X1 U920 ( .A(n1243), .ZN(n1216) );
NOR2_X1 U921 ( .A1(n1082), .A2(n1209), .ZN(n1243) );
XOR2_X1 U922 ( .A(n1255), .B(KEYINPUT36), .Z(n1082) );
XOR2_X1 U923 ( .A(n1256), .B(n1257), .Z(G30) );
NOR2_X1 U924 ( .A1(n1258), .A2(n1210), .ZN(n1257) );
NAND4_X1 U925 ( .A1(n1073), .A2(n1236), .A3(n1259), .A4(n1255), .ZN(n1210) );
NOR2_X1 U926 ( .A1(n1248), .A2(n1247), .ZN(n1259) );
XNOR2_X1 U927 ( .A(n1209), .B(KEYINPUT38), .ZN(n1258) );
INV_X1 U928 ( .A(n1260), .ZN(n1209) );
XNOR2_X1 U929 ( .A(G128), .B(KEYINPUT5), .ZN(n1256) );
XNOR2_X1 U930 ( .A(n1178), .B(n1228), .ZN(G3) );
AND3_X1 U931 ( .A1(n1074), .A2(n1227), .A3(n1254), .ZN(n1228) );
XNOR2_X1 U932 ( .A(G125), .B(n1203), .ZN(G27) );
NAND4_X1 U933 ( .A1(n1236), .A2(n1260), .A3(n1244), .A4(n1261), .ZN(n1203) );
NOR2_X1 U934 ( .A1(n1262), .A2(n1219), .ZN(n1261) );
NAND2_X1 U935 ( .A1(n1091), .A2(n1263), .ZN(n1260) );
NAND4_X1 U936 ( .A1(G902), .A2(G953), .A3(n1264), .A4(n1265), .ZN(n1263) );
INV_X1 U937 ( .A(G900), .ZN(n1265) );
XOR2_X1 U938 ( .A(n1221), .B(n1266), .Z(G24) );
XNOR2_X1 U939 ( .A(G122), .B(KEYINPUT31), .ZN(n1266) );
NAND4_X1 U940 ( .A1(n1267), .A2(n1070), .A3(n1239), .A4(n1240), .ZN(n1221) );
INV_X1 U941 ( .A(n1102), .ZN(n1070) );
NAND2_X1 U942 ( .A1(n1248), .A2(n1247), .ZN(n1102) );
XOR2_X1 U943 ( .A(G119), .B(n1268), .Z(G21) );
NOR2_X1 U944 ( .A1(n1087), .A2(n1231), .ZN(n1268) );
NAND3_X1 U945 ( .A1(n1065), .A2(n1074), .A3(n1269), .ZN(n1231) );
NOR3_X1 U946 ( .A1(n1247), .A2(n1270), .A3(n1248), .ZN(n1269) );
INV_X1 U947 ( .A(n1271), .ZN(n1247) );
INV_X1 U948 ( .A(n1262), .ZN(n1065) );
XOR2_X1 U949 ( .A(G116), .B(n1226), .Z(G18) );
AND3_X1 U950 ( .A1(n1267), .A2(n1073), .A3(n1254), .ZN(n1226) );
NOR2_X1 U951 ( .A1(n1240), .A2(n1272), .ZN(n1073) );
XOR2_X1 U952 ( .A(G113), .B(n1273), .Z(G15) );
NOR2_X1 U953 ( .A1(KEYINPUT11), .A2(n1222), .ZN(n1273) );
NAND3_X1 U954 ( .A1(n1254), .A2(n1267), .A3(n1072), .ZN(n1222) );
INV_X1 U955 ( .A(n1219), .ZN(n1072) );
NAND2_X1 U956 ( .A1(n1272), .A2(n1240), .ZN(n1219) );
INV_X1 U957 ( .A(n1239), .ZN(n1272) );
NOR3_X1 U958 ( .A1(n1087), .A2(n1270), .A3(n1262), .ZN(n1267) );
NAND2_X1 U959 ( .A1(n1085), .A2(n1274), .ZN(n1262) );
NOR2_X1 U960 ( .A1(n1271), .A2(n1248), .ZN(n1254) );
XNOR2_X1 U961 ( .A(n1152), .B(n1225), .ZN(G12) );
AND3_X1 U962 ( .A1(n1244), .A2(n1227), .A3(n1074), .ZN(n1225) );
NOR2_X1 U963 ( .A1(n1239), .A2(n1240), .ZN(n1074) );
NAND3_X1 U964 ( .A1(n1275), .A2(n1276), .A3(n1101), .ZN(n1240) );
NAND2_X1 U965 ( .A1(n1099), .A2(n1100), .ZN(n1101) );
OR3_X1 U966 ( .A1(n1100), .A2(n1099), .A3(KEYINPUT44), .ZN(n1276) );
AND2_X1 U967 ( .A1(n1168), .A2(n1277), .ZN(n1099) );
XOR2_X1 U968 ( .A(n1278), .B(n1279), .Z(n1168) );
XNOR2_X1 U969 ( .A(n1148), .B(n1280), .ZN(n1279) );
XOR2_X1 U970 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR2_X1 U971 ( .A1(KEYINPUT33), .A2(n1283), .ZN(n1282) );
XOR2_X1 U972 ( .A(G143), .B(n1284), .Z(n1283) );
NOR3_X1 U973 ( .A1(n1285), .A2(G953), .A3(n1286), .ZN(n1284) );
INV_X1 U974 ( .A(G214), .ZN(n1286) );
NAND2_X1 U975 ( .A1(n1287), .A2(n1288), .ZN(n1281) );
NAND2_X1 U976 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XNOR2_X1 U977 ( .A(n1291), .B(n1119), .ZN(n1290) );
XNOR2_X1 U978 ( .A(G146), .B(KEYINPUT26), .ZN(n1289) );
XOR2_X1 U979 ( .A(n1292), .B(KEYINPUT60), .Z(n1287) );
NAND2_X1 U980 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XNOR2_X1 U981 ( .A(G125), .B(n1119), .ZN(n1293) );
XOR2_X1 U982 ( .A(G113), .B(G122), .Z(n1148) );
XNOR2_X1 U983 ( .A(G104), .B(n1295), .ZN(n1278) );
XNOR2_X1 U984 ( .A(KEYINPUT15), .B(n1250), .ZN(n1295) );
INV_X1 U985 ( .A(G131), .ZN(n1250) );
NAND2_X1 U986 ( .A1(KEYINPUT44), .A2(n1100), .ZN(n1275) );
XOR2_X1 U987 ( .A(G475), .B(KEYINPUT1), .Z(n1100) );
XNOR2_X1 U988 ( .A(n1296), .B(G478), .ZN(n1239) );
NAND2_X1 U989 ( .A1(KEYINPUT23), .A2(n1104), .ZN(n1296) );
AND2_X1 U990 ( .A1(n1165), .A2(n1277), .ZN(n1104) );
XNOR2_X1 U991 ( .A(n1297), .B(n1298), .ZN(n1165) );
XNOR2_X1 U992 ( .A(n1299), .B(n1300), .ZN(n1298) );
NOR3_X1 U993 ( .A1(n1301), .A2(KEYINPUT49), .A3(n1302), .ZN(n1300) );
INV_X1 U994 ( .A(G217), .ZN(n1301) );
NAND2_X1 U995 ( .A1(KEYINPUT37), .A2(n1303), .ZN(n1299) );
XNOR2_X1 U996 ( .A(n1133), .B(n1304), .ZN(n1303) );
XNOR2_X1 U997 ( .A(G107), .B(n1305), .ZN(n1297) );
XOR2_X1 U998 ( .A(G122), .B(G116), .Z(n1305) );
NOR3_X1 U999 ( .A1(n1306), .A2(n1270), .A3(n1087), .ZN(n1227) );
INV_X1 U1000 ( .A(n1236), .ZN(n1087) );
NOR2_X1 U1001 ( .A1(n1090), .A2(n1089), .ZN(n1236) );
INV_X1 U1002 ( .A(n1253), .ZN(n1089) );
NAND2_X1 U1003 ( .A1(n1307), .A2(n1308), .ZN(n1253) );
XNOR2_X1 U1004 ( .A(G214), .B(KEYINPUT29), .ZN(n1307) );
XOR2_X1 U1005 ( .A(n1106), .B(n1309), .Z(n1090) );
NOR2_X1 U1006 ( .A1(KEYINPUT50), .A2(n1107), .ZN(n1309) );
NAND2_X1 U1007 ( .A1(G210), .A2(n1308), .ZN(n1107) );
NAND2_X1 U1008 ( .A1(n1310), .A2(n1277), .ZN(n1308) );
INV_X1 U1009 ( .A(G237), .ZN(n1310) );
NAND2_X1 U1010 ( .A1(n1311), .A2(n1277), .ZN(n1106) );
XOR2_X1 U1011 ( .A(n1312), .B(n1313), .Z(n1311) );
XNOR2_X1 U1012 ( .A(n1314), .B(n1188), .ZN(n1313) );
INV_X1 U1013 ( .A(n1177), .ZN(n1188) );
NOR2_X1 U1014 ( .A1(G125), .A2(n1315), .ZN(n1314) );
XOR2_X1 U1015 ( .A(KEYINPUT40), .B(KEYINPUT20), .Z(n1315) );
XNOR2_X1 U1016 ( .A(n1232), .B(n1234), .ZN(n1312) );
NOR2_X1 U1017 ( .A1(n1137), .A2(G953), .ZN(n1234) );
INV_X1 U1018 ( .A(G224), .ZN(n1137) );
NAND2_X1 U1019 ( .A1(n1316), .A2(n1317), .ZN(n1232) );
NAND2_X1 U1020 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
XNOR2_X1 U1021 ( .A(n1320), .B(n1321), .ZN(n1319) );
XNOR2_X1 U1022 ( .A(G122), .B(G110), .ZN(n1318) );
XOR2_X1 U1023 ( .A(n1322), .B(KEYINPUT59), .Z(n1316) );
NAND2_X1 U1024 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1025 ( .A(n1321), .B(n1320), .Z(n1324) );
XOR2_X1 U1026 ( .A(n1150), .B(G113), .Z(n1320) );
NAND2_X1 U1027 ( .A1(n1325), .A2(KEYINPUT6), .ZN(n1150) );
XNOR2_X1 U1028 ( .A(n1326), .B(KEYINPUT17), .ZN(n1325) );
NAND2_X1 U1029 ( .A1(KEYINPUT0), .A2(n1149), .ZN(n1321) );
XNOR2_X1 U1030 ( .A(n1178), .B(n1327), .ZN(n1149) );
NOR2_X1 U1031 ( .A1(KEYINPUT19), .A2(n1328), .ZN(n1327) );
XNOR2_X1 U1032 ( .A(G104), .B(G107), .ZN(n1328) );
XNOR2_X1 U1033 ( .A(G122), .B(n1152), .ZN(n1323) );
AND2_X1 U1034 ( .A1(n1091), .A2(n1329), .ZN(n1270) );
NAND4_X1 U1035 ( .A1(G902), .A2(G953), .A3(n1264), .A4(n1138), .ZN(n1329) );
INV_X1 U1036 ( .A(G898), .ZN(n1138) );
NAND3_X1 U1037 ( .A1(n1264), .A2(n1059), .A3(G952), .ZN(n1091) );
NAND2_X1 U1038 ( .A1(G237), .A2(G234), .ZN(n1264) );
INV_X1 U1039 ( .A(n1255), .ZN(n1306) );
NOR2_X1 U1040 ( .A1(n1085), .A2(n1084), .ZN(n1255) );
INV_X1 U1041 ( .A(n1274), .ZN(n1084) );
NAND2_X1 U1042 ( .A1(G221), .A2(n1330), .ZN(n1274) );
XOR2_X1 U1043 ( .A(G469), .B(n1331), .Z(n1085) );
NOR2_X1 U1044 ( .A1(n1105), .A2(KEYINPUT52), .ZN(n1331) );
AND2_X1 U1045 ( .A1(n1332), .A2(n1277), .ZN(n1105) );
XOR2_X1 U1046 ( .A(n1333), .B(n1334), .Z(n1332) );
XOR2_X1 U1047 ( .A(n1335), .B(n1336), .Z(n1334) );
XNOR2_X1 U1048 ( .A(G110), .B(n1337), .ZN(n1336) );
NOR2_X1 U1049 ( .A1(KEYINPUT30), .A2(n1338), .ZN(n1337) );
XNOR2_X1 U1050 ( .A(n1196), .B(n1177), .ZN(n1338) );
AND2_X1 U1051 ( .A1(n1339), .A2(n1340), .ZN(n1196) );
NAND2_X1 U1052 ( .A1(G104), .A2(n1341), .ZN(n1340) );
NAND2_X1 U1053 ( .A1(n1342), .A2(n1169), .ZN(n1339) );
INV_X1 U1054 ( .A(G104), .ZN(n1169) );
XNOR2_X1 U1055 ( .A(KEYINPUT16), .B(n1341), .ZN(n1342) );
XOR2_X1 U1056 ( .A(n1178), .B(n1343), .Z(n1341) );
XOR2_X1 U1057 ( .A(KEYINPUT8), .B(G107), .Z(n1343) );
INV_X1 U1058 ( .A(G101), .ZN(n1178) );
NAND2_X1 U1059 ( .A1(KEYINPUT53), .A2(n1192), .ZN(n1335) );
AND2_X1 U1060 ( .A1(G227), .A2(n1344), .ZN(n1192) );
XNOR2_X1 U1061 ( .A(KEYINPUT42), .B(n1059), .ZN(n1344) );
XOR2_X1 U1062 ( .A(n1183), .B(n1345), .Z(n1333) );
NOR2_X1 U1063 ( .A1(KEYINPUT58), .A2(n1119), .ZN(n1345) );
INV_X1 U1064 ( .A(n1076), .ZN(n1244) );
NAND2_X1 U1065 ( .A1(n1248), .A2(n1271), .ZN(n1076) );
XNOR2_X1 U1066 ( .A(n1346), .B(n1161), .ZN(n1271) );
AND2_X1 U1067 ( .A1(G217), .A2(n1330), .ZN(n1161) );
NAND2_X1 U1068 ( .A1(G234), .A2(n1277), .ZN(n1330) );
NAND2_X1 U1069 ( .A1(n1162), .A2(n1277), .ZN(n1346) );
XOR2_X1 U1070 ( .A(n1347), .B(n1348), .Z(n1162) );
XOR2_X1 U1071 ( .A(n1349), .B(n1350), .Z(n1348) );
XNOR2_X1 U1072 ( .A(G119), .B(n1152), .ZN(n1350) );
XNOR2_X1 U1073 ( .A(n1294), .B(G128), .ZN(n1349) );
INV_X1 U1074 ( .A(G146), .ZN(n1294) );
XOR2_X1 U1075 ( .A(n1351), .B(n1352), .Z(n1347) );
XOR2_X1 U1076 ( .A(n1353), .B(n1354), .Z(n1352) );
NAND2_X1 U1077 ( .A1(n1355), .A2(G221), .ZN(n1354) );
INV_X1 U1078 ( .A(n1302), .ZN(n1355) );
NAND2_X1 U1079 ( .A1(G234), .A2(n1059), .ZN(n1302) );
INV_X1 U1080 ( .A(G953), .ZN(n1059) );
NAND3_X1 U1081 ( .A1(n1356), .A2(n1357), .A3(n1358), .ZN(n1353) );
OR2_X1 U1082 ( .A1(n1291), .A2(n1119), .ZN(n1358) );
NAND2_X1 U1083 ( .A1(KEYINPUT24), .A2(n1359), .ZN(n1357) );
NAND2_X1 U1084 ( .A1(n1360), .A2(n1291), .ZN(n1359) );
XNOR2_X1 U1085 ( .A(KEYINPUT47), .B(n1119), .ZN(n1360) );
NAND2_X1 U1086 ( .A1(n1361), .A2(n1362), .ZN(n1356) );
INV_X1 U1087 ( .A(KEYINPUT24), .ZN(n1362) );
NAND2_X1 U1088 ( .A1(n1363), .A2(n1364), .ZN(n1361) );
OR2_X1 U1089 ( .A1(n1119), .A2(KEYINPUT47), .ZN(n1364) );
NAND3_X1 U1090 ( .A1(n1119), .A2(n1291), .A3(KEYINPUT47), .ZN(n1363) );
INV_X1 U1091 ( .A(G125), .ZN(n1291) );
XOR2_X1 U1092 ( .A(G140), .B(KEYINPUT34), .Z(n1119) );
NAND2_X1 U1093 ( .A1(KEYINPUT39), .A2(G137), .ZN(n1351) );
XOR2_X1 U1094 ( .A(n1365), .B(G472), .Z(n1248) );
NAND2_X1 U1095 ( .A1(n1366), .A2(n1277), .ZN(n1365) );
INV_X1 U1096 ( .A(G902), .ZN(n1277) );
XOR2_X1 U1097 ( .A(n1367), .B(n1368), .Z(n1366) );
XNOR2_X1 U1098 ( .A(n1183), .B(n1174), .ZN(n1368) );
XNOR2_X1 U1099 ( .A(n1369), .B(n1370), .ZN(n1174) );
XOR2_X1 U1100 ( .A(KEYINPUT62), .B(KEYINPUT14), .Z(n1370) );
XNOR2_X1 U1101 ( .A(G113), .B(n1326), .ZN(n1369) );
XOR2_X1 U1102 ( .A(G116), .B(G119), .Z(n1326) );
XOR2_X1 U1103 ( .A(n1371), .B(n1372), .Z(n1183) );
NOR3_X1 U1104 ( .A1(n1373), .A2(n1374), .A3(n1375), .ZN(n1372) );
NOR2_X1 U1105 ( .A1(G137), .A2(n1376), .ZN(n1375) );
NOR3_X1 U1106 ( .A1(n1377), .A2(KEYINPUT45), .A3(n1132), .ZN(n1374) );
INV_X1 U1107 ( .A(G137), .ZN(n1132) );
INV_X1 U1108 ( .A(n1376), .ZN(n1377) );
NOR2_X1 U1109 ( .A1(KEYINPUT21), .A2(n1133), .ZN(n1376) );
AND2_X1 U1110 ( .A1(n1133), .A2(KEYINPUT45), .ZN(n1373) );
INV_X1 U1111 ( .A(G134), .ZN(n1133) );
NAND2_X1 U1112 ( .A1(n1378), .A2(KEYINPUT27), .ZN(n1371) );
XNOR2_X1 U1113 ( .A(n1124), .B(KEYINPUT10), .ZN(n1378) );
XOR2_X1 U1114 ( .A(G131), .B(KEYINPUT32), .Z(n1124) );
XOR2_X1 U1115 ( .A(n1379), .B(n1380), .Z(n1367) );
XNOR2_X1 U1116 ( .A(G101), .B(n1381), .ZN(n1380) );
NAND2_X1 U1117 ( .A1(KEYINPUT2), .A2(n1177), .ZN(n1381) );
XOR2_X1 U1118 ( .A(G146), .B(n1304), .Z(n1177) );
XOR2_X1 U1119 ( .A(G128), .B(G143), .Z(n1304) );
NAND2_X1 U1120 ( .A1(KEYINPUT57), .A2(n1182), .ZN(n1379) );
NOR3_X1 U1121 ( .A1(n1382), .A2(G953), .A3(n1285), .ZN(n1182) );
XOR2_X1 U1122 ( .A(G237), .B(KEYINPUT18), .Z(n1285) );
INV_X1 U1123 ( .A(G210), .ZN(n1382) );
INV_X1 U1124 ( .A(G110), .ZN(n1152) );
endmodule


