//Key = 1101001000110111110111011110010111110111100100010010010101100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337;

XNOR2_X1 U752 ( .A(G107), .B(n1021), .ZN(G9) );
NOR2_X1 U753 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR4_X1 U754 ( .A1(G953), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1023) );
NOR2_X1 U755 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR2_X1 U756 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U757 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
INV_X1 U758 ( .A(n1033), .ZN(n1032) );
NOR2_X1 U759 ( .A1(n1034), .A2(n1035), .ZN(n1031) );
NOR2_X1 U760 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR2_X1 U761 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U762 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U763 ( .A1(n1042), .A2(n1043), .ZN(n1038) );
NOR3_X1 U764 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1042) );
AND2_X1 U765 ( .A1(n1047), .A2(KEYINPUT9), .ZN(n1046) );
NOR2_X1 U766 ( .A1(n1048), .A2(n1049), .ZN(n1044) );
NOR3_X1 U767 ( .A1(n1041), .A2(n1050), .A3(n1043), .ZN(n1034) );
NOR2_X1 U768 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U769 ( .A1(n1053), .A2(KEYINPUT9), .A3(n1054), .ZN(n1051) );
NOR4_X1 U770 ( .A1(n1055), .A2(n1043), .A3(n1041), .A4(n1037), .ZN(n1029) );
INV_X1 U771 ( .A(n1056), .ZN(n1037) );
INV_X1 U772 ( .A(n1047), .ZN(n1041) );
INV_X1 U773 ( .A(n1057), .ZN(n1043) );
NOR2_X1 U774 ( .A1(n1058), .A2(n1059), .ZN(n1055) );
NOR3_X1 U775 ( .A1(n1024), .A2(G953), .A3(G952), .ZN(n1022) );
AND4_X1 U776 ( .A1(n1047), .A2(n1053), .A3(n1033), .A4(n1060), .ZN(n1024) );
NOR3_X1 U777 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NOR2_X1 U778 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
INV_X1 U779 ( .A(KEYINPUT30), .ZN(n1065) );
NOR2_X1 U780 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U781 ( .A1(KEYINPUT30), .A2(n1057), .ZN(n1062) );
XOR2_X1 U782 ( .A(n1068), .B(n1069), .Z(n1061) );
XNOR2_X1 U783 ( .A(G469), .B(KEYINPUT62), .ZN(n1069) );
NAND2_X1 U784 ( .A1(KEYINPUT57), .A2(n1070), .ZN(n1068) );
XOR2_X1 U785 ( .A(n1071), .B(n1072), .Z(G72) );
NOR2_X1 U786 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U787 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NAND2_X1 U788 ( .A1(n1077), .A2(n1078), .ZN(n1071) );
NAND2_X1 U789 ( .A1(n1079), .A2(n1074), .ZN(n1078) );
XOR2_X1 U790 ( .A(n1080), .B(n1081), .Z(n1079) );
NAND3_X1 U791 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1080) );
INV_X1 U792 ( .A(n1085), .ZN(n1084) );
XOR2_X1 U793 ( .A(KEYINPUT63), .B(n1086), .Z(n1082) );
NAND3_X1 U794 ( .A1(G900), .A2(n1081), .A3(G953), .ZN(n1077) );
XNOR2_X1 U795 ( .A(n1087), .B(n1088), .ZN(n1081) );
XNOR2_X1 U796 ( .A(n1089), .B(n1090), .ZN(n1088) );
NOR2_X1 U797 ( .A1(G137), .A2(KEYINPUT8), .ZN(n1090) );
NAND2_X1 U798 ( .A1(KEYINPUT53), .A2(n1091), .ZN(n1089) );
XOR2_X1 U799 ( .A(n1092), .B(n1093), .Z(n1087) );
NOR3_X1 U800 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
NOR2_X1 U801 ( .A1(G134), .A2(n1097), .ZN(n1096) );
AND3_X1 U802 ( .A1(G134), .A2(G140), .A3(G125), .ZN(n1095) );
NOR2_X1 U803 ( .A1(G140), .A2(n1098), .ZN(n1094) );
XNOR2_X1 U804 ( .A(G134), .B(G125), .ZN(n1098) );
NAND2_X1 U805 ( .A1(n1099), .A2(n1100), .ZN(G69) );
NAND2_X1 U806 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U807 ( .A(KEYINPUT32), .B(n1103), .Z(n1099) );
NOR2_X1 U808 ( .A1(n1104), .A2(n1102), .ZN(n1103) );
NAND2_X1 U809 ( .A1(G953), .A2(n1105), .ZN(n1102) );
NAND2_X1 U810 ( .A1(G898), .A2(G224), .ZN(n1105) );
XNOR2_X1 U811 ( .A(n1101), .B(KEYINPUT24), .ZN(n1104) );
XNOR2_X1 U812 ( .A(n1106), .B(n1107), .ZN(n1101) );
NOR2_X1 U813 ( .A1(n1108), .A2(G953), .ZN(n1107) );
NOR2_X1 U814 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND3_X1 U815 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1106) );
INV_X1 U816 ( .A(n1114), .ZN(n1113) );
NAND2_X1 U817 ( .A1(G953), .A2(n1115), .ZN(n1111) );
NOR2_X1 U818 ( .A1(n1116), .A2(n1117), .ZN(G66) );
XNOR2_X1 U819 ( .A(n1118), .B(n1119), .ZN(n1117) );
NOR2_X1 U820 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U821 ( .A1(n1116), .A2(n1122), .ZN(G63) );
XOR2_X1 U822 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U823 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U824 ( .A1(n1127), .A2(n1121), .ZN(n1125) );
INV_X1 U825 ( .A(G478), .ZN(n1127) );
XNOR2_X1 U826 ( .A(KEYINPUT54), .B(KEYINPUT10), .ZN(n1123) );
NOR2_X1 U827 ( .A1(n1116), .A2(n1128), .ZN(G60) );
XNOR2_X1 U828 ( .A(n1129), .B(n1130), .ZN(n1128) );
NOR2_X1 U829 ( .A1(n1131), .A2(n1121), .ZN(n1130) );
XNOR2_X1 U830 ( .A(G104), .B(n1132), .ZN(G6) );
NOR2_X1 U831 ( .A1(n1116), .A2(n1133), .ZN(G57) );
XOR2_X1 U832 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U833 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U834 ( .A(n1138), .B(n1139), .Z(n1134) );
XOR2_X1 U835 ( .A(n1140), .B(n1141), .Z(n1138) );
NOR2_X1 U836 ( .A1(n1142), .A2(n1121), .ZN(n1141) );
NAND2_X1 U837 ( .A1(KEYINPUT26), .A2(n1143), .ZN(n1140) );
NOR2_X1 U838 ( .A1(n1116), .A2(n1144), .ZN(G54) );
XOR2_X1 U839 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U840 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U841 ( .A1(n1149), .A2(n1121), .ZN(n1147) );
XOR2_X1 U842 ( .A(n1150), .B(n1151), .Z(n1145) );
NOR2_X1 U843 ( .A1(KEYINPUT28), .A2(n1152), .ZN(n1151) );
XOR2_X1 U844 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U845 ( .A1(KEYINPUT45), .A2(n1155), .ZN(n1154) );
XNOR2_X1 U846 ( .A(KEYINPUT15), .B(n1092), .ZN(n1155) );
NAND2_X1 U847 ( .A1(n1156), .A2(KEYINPUT34), .ZN(n1150) );
XNOR2_X1 U848 ( .A(G110), .B(KEYINPUT18), .ZN(n1156) );
NOR2_X1 U849 ( .A1(n1116), .A2(n1157), .ZN(G51) );
XOR2_X1 U850 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U851 ( .A1(n1160), .A2(n1121), .ZN(n1159) );
NAND2_X1 U852 ( .A1(G902), .A2(n1026), .ZN(n1121) );
NAND3_X1 U853 ( .A1(n1161), .A2(n1086), .A3(n1162), .ZN(n1026) );
NOR3_X1 U854 ( .A1(n1085), .A2(n1163), .A3(n1110), .ZN(n1162) );
NAND3_X1 U855 ( .A1(n1132), .A2(n1021), .A3(n1164), .ZN(n1110) );
OR2_X1 U856 ( .A1(n1165), .A2(n1040), .ZN(n1164) );
NOR2_X1 U857 ( .A1(n1166), .A2(n1167), .ZN(n1040) );
NAND3_X1 U858 ( .A1(n1168), .A2(n1058), .A3(n1057), .ZN(n1021) );
NAND3_X1 U859 ( .A1(n1057), .A2(n1168), .A3(n1059), .ZN(n1132) );
INV_X1 U860 ( .A(n1083), .ZN(n1163) );
NAND2_X1 U861 ( .A1(n1169), .A2(n1059), .ZN(n1083) );
NAND3_X1 U862 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1085) );
AND4_X1 U863 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1086) );
NAND2_X1 U864 ( .A1(n1177), .A2(n1178), .ZN(n1173) );
XOR2_X1 U865 ( .A(n1109), .B(KEYINPUT38), .Z(n1161) );
NAND4_X1 U866 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1109) );
NAND3_X1 U867 ( .A1(n1059), .A2(n1166), .A3(n1183), .ZN(n1179) );
XOR2_X1 U868 ( .A(n1184), .B(n1185), .Z(n1158) );
NOR2_X1 U869 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
XOR2_X1 U870 ( .A(n1188), .B(KEYINPUT55), .Z(n1187) );
NAND2_X1 U871 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NOR2_X1 U872 ( .A1(n1189), .A2(n1190), .ZN(n1186) );
XNOR2_X1 U873 ( .A(n1191), .B(G125), .ZN(n1190) );
NAND2_X1 U874 ( .A1(KEYINPUT11), .A2(n1192), .ZN(n1191) );
NOR2_X1 U875 ( .A1(n1074), .A2(G952), .ZN(n1116) );
XOR2_X1 U876 ( .A(n1193), .B(n1194), .Z(G48) );
XOR2_X1 U877 ( .A(KEYINPUT50), .B(G146), .Z(n1194) );
NAND3_X1 U878 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1193) );
XOR2_X1 U879 ( .A(KEYINPUT59), .B(n1052), .Z(n1196) );
XOR2_X1 U880 ( .A(n1198), .B(n1199), .Z(G45) );
XNOR2_X1 U881 ( .A(KEYINPUT61), .B(n1200), .ZN(n1199) );
NAND2_X1 U882 ( .A1(KEYINPUT25), .A2(n1171), .ZN(n1198) );
NAND3_X1 U883 ( .A1(n1201), .A2(n1166), .A3(n1202), .ZN(n1171) );
AND3_X1 U884 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1202) );
XNOR2_X1 U885 ( .A(G140), .B(n1172), .ZN(G42) );
NAND3_X1 U886 ( .A1(n1167), .A2(n1059), .A3(n1178), .ZN(n1172) );
XNOR2_X1 U887 ( .A(G137), .B(n1170), .ZN(G39) );
NAND3_X1 U888 ( .A1(n1197), .A2(n1033), .A3(n1178), .ZN(n1170) );
XNOR2_X1 U889 ( .A(G134), .B(n1206), .ZN(G36) );
NAND4_X1 U890 ( .A1(n1177), .A2(n1047), .A3(n1052), .A4(n1207), .ZN(n1206) );
XNOR2_X1 U891 ( .A(KEYINPUT14), .B(n1204), .ZN(n1207) );
XOR2_X1 U892 ( .A(n1174), .B(n1208), .Z(G33) );
NAND2_X1 U893 ( .A1(KEYINPUT37), .A2(G131), .ZN(n1208) );
NAND3_X1 U894 ( .A1(n1059), .A2(n1166), .A3(n1178), .ZN(n1174) );
AND3_X1 U895 ( .A1(n1052), .A2(n1204), .A3(n1047), .ZN(n1178) );
NOR2_X1 U896 ( .A1(n1048), .A2(n1209), .ZN(n1047) );
INV_X1 U897 ( .A(n1049), .ZN(n1209) );
XNOR2_X1 U898 ( .A(n1175), .B(n1210), .ZN(G30) );
NOR2_X1 U899 ( .A1(KEYINPUT60), .A2(n1211), .ZN(n1210) );
NAND2_X1 U900 ( .A1(n1169), .A2(n1058), .ZN(n1175) );
AND3_X1 U901 ( .A1(n1201), .A2(n1204), .A3(n1197), .ZN(n1169) );
XNOR2_X1 U902 ( .A(G101), .B(n1212), .ZN(G3) );
NAND3_X1 U903 ( .A1(n1213), .A2(n1166), .A3(KEYINPUT13), .ZN(n1212) );
INV_X1 U904 ( .A(n1165), .ZN(n1213) );
XNOR2_X1 U905 ( .A(G125), .B(n1176), .ZN(G27) );
NAND3_X1 U906 ( .A1(n1056), .A2(n1195), .A3(n1167), .ZN(n1176) );
AND3_X1 U907 ( .A1(n1045), .A2(n1204), .A3(n1059), .ZN(n1195) );
NAND2_X1 U908 ( .A1(n1028), .A2(n1214), .ZN(n1204) );
NAND4_X1 U909 ( .A1(G953), .A2(G902), .A3(n1215), .A4(n1076), .ZN(n1214) );
INV_X1 U910 ( .A(G900), .ZN(n1076) );
XNOR2_X1 U911 ( .A(G122), .B(n1180), .ZN(G24) );
NAND4_X1 U912 ( .A1(n1183), .A2(n1057), .A3(n1203), .A4(n1205), .ZN(n1180) );
NOR2_X1 U913 ( .A1(n1216), .A2(n1067), .ZN(n1057) );
XNOR2_X1 U914 ( .A(G119), .B(n1181), .ZN(G21) );
NAND3_X1 U915 ( .A1(n1197), .A2(n1033), .A3(n1183), .ZN(n1181) );
XNOR2_X1 U916 ( .A(G116), .B(n1182), .ZN(G18) );
NAND2_X1 U917 ( .A1(n1183), .A2(n1177), .ZN(n1182) );
AND2_X1 U918 ( .A1(n1058), .A2(n1166), .ZN(n1177) );
NOR2_X1 U919 ( .A1(n1205), .A2(n1217), .ZN(n1058) );
AND3_X1 U920 ( .A1(n1045), .A2(n1218), .A3(n1056), .ZN(n1183) );
XNOR2_X1 U921 ( .A(G113), .B(n1219), .ZN(G15) );
NAND4_X1 U922 ( .A1(KEYINPUT20), .A2(n1056), .A3(n1220), .A4(n1221), .ZN(n1219) );
AND3_X1 U923 ( .A1(n1059), .A2(n1218), .A3(n1166), .ZN(n1221) );
NAND2_X1 U924 ( .A1(n1222), .A2(n1223), .ZN(n1166) );
NAND2_X1 U925 ( .A1(n1197), .A2(n1224), .ZN(n1223) );
AND2_X1 U926 ( .A1(n1067), .A2(n1216), .ZN(n1197) );
OR3_X1 U927 ( .A1(n1066), .A2(n1067), .A3(n1224), .ZN(n1222) );
INV_X1 U928 ( .A(KEYINPUT31), .ZN(n1224) );
AND2_X1 U929 ( .A1(n1217), .A2(n1205), .ZN(n1059) );
INV_X1 U930 ( .A(n1203), .ZN(n1217) );
XNOR2_X1 U931 ( .A(n1045), .B(KEYINPUT0), .ZN(n1220) );
NOR2_X1 U932 ( .A1(n1054), .A2(n1225), .ZN(n1056) );
INV_X1 U933 ( .A(n1053), .ZN(n1225) );
XOR2_X1 U934 ( .A(n1226), .B(n1227), .Z(G12) );
NOR2_X1 U935 ( .A1(n1165), .A2(n1228), .ZN(n1227) );
XOR2_X1 U936 ( .A(KEYINPUT35), .B(n1167), .Z(n1228) );
AND2_X1 U937 ( .A1(n1066), .A2(n1067), .ZN(n1167) );
XNOR2_X1 U938 ( .A(n1229), .B(n1230), .ZN(n1067) );
NOR2_X1 U939 ( .A1(n1231), .A2(n1120), .ZN(n1230) );
INV_X1 U940 ( .A(G217), .ZN(n1120) );
XOR2_X1 U941 ( .A(n1232), .B(KEYINPUT3), .Z(n1231) );
NAND2_X1 U942 ( .A1(n1118), .A2(n1233), .ZN(n1229) );
XNOR2_X1 U943 ( .A(n1234), .B(n1235), .ZN(n1118) );
XNOR2_X1 U944 ( .A(n1236), .B(n1137), .ZN(n1235) );
XNOR2_X1 U945 ( .A(G119), .B(n1211), .ZN(n1137) );
NAND2_X1 U946 ( .A1(KEYINPUT39), .A2(n1237), .ZN(n1236) );
XOR2_X1 U947 ( .A(n1238), .B(n1239), .Z(n1234) );
XOR2_X1 U948 ( .A(n1240), .B(n1241), .Z(n1239) );
XOR2_X1 U949 ( .A(KEYINPUT19), .B(G146), .Z(n1241) );
XOR2_X1 U950 ( .A(KEYINPUT51), .B(KEYINPUT42), .Z(n1240) );
XOR2_X1 U951 ( .A(n1242), .B(n1243), .Z(n1238) );
XOR2_X1 U952 ( .A(G140), .B(G137), .Z(n1243) );
XNOR2_X1 U953 ( .A(n1244), .B(n1245), .ZN(n1242) );
NAND3_X1 U954 ( .A1(G221), .A2(n1074), .A3(n1246), .ZN(n1244) );
XNOR2_X1 U955 ( .A(G234), .B(KEYINPUT17), .ZN(n1246) );
INV_X1 U956 ( .A(n1216), .ZN(n1066) );
XOR2_X1 U957 ( .A(n1247), .B(n1142), .Z(n1216) );
INV_X1 U958 ( .A(G472), .ZN(n1142) );
NAND2_X1 U959 ( .A1(n1248), .A2(n1233), .ZN(n1247) );
XOR2_X1 U960 ( .A(n1249), .B(n1250), .Z(n1248) );
XOR2_X1 U961 ( .A(n1136), .B(n1251), .Z(n1250) );
XOR2_X1 U962 ( .A(n1252), .B(n1253), .Z(n1136) );
NOR2_X1 U963 ( .A1(G116), .A2(KEYINPUT56), .ZN(n1253) );
XNOR2_X1 U964 ( .A(G101), .B(n1254), .ZN(n1252) );
NOR2_X1 U965 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XOR2_X1 U966 ( .A(KEYINPUT16), .B(G210), .Z(n1256) );
XOR2_X1 U967 ( .A(n1257), .B(KEYINPUT12), .Z(n1249) );
NAND3_X1 U968 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1257) );
NAND2_X1 U969 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
OR3_X1 U970 ( .A1(n1262), .A2(n1261), .A3(KEYINPUT7), .ZN(n1259) );
NAND2_X1 U971 ( .A1(n1192), .A2(n1263), .ZN(n1262) );
XOR2_X1 U972 ( .A(KEYINPUT6), .B(KEYINPUT2), .Z(n1263) );
NAND2_X1 U973 ( .A1(n1264), .A2(KEYINPUT7), .ZN(n1258) );
NAND2_X1 U974 ( .A1(n1033), .A2(n1168), .ZN(n1165) );
AND2_X1 U975 ( .A1(n1201), .A2(n1218), .ZN(n1168) );
NAND2_X1 U976 ( .A1(n1028), .A2(n1265), .ZN(n1218) );
NAND4_X1 U977 ( .A1(G953), .A2(G902), .A3(n1215), .A4(n1115), .ZN(n1265) );
INV_X1 U978 ( .A(G898), .ZN(n1115) );
NAND3_X1 U979 ( .A1(n1215), .A2(n1074), .A3(G952), .ZN(n1028) );
NAND2_X1 U980 ( .A1(G234), .A2(G237), .ZN(n1215) );
AND2_X1 U981 ( .A1(n1052), .A2(n1045), .ZN(n1201) );
AND2_X1 U982 ( .A1(n1048), .A2(n1049), .ZN(n1045) );
NAND2_X1 U983 ( .A1(G214), .A2(n1266), .ZN(n1049) );
XOR2_X1 U984 ( .A(n1267), .B(n1160), .Z(n1048) );
NAND2_X1 U985 ( .A1(G210), .A2(n1266), .ZN(n1160) );
NAND2_X1 U986 ( .A1(n1268), .A2(n1233), .ZN(n1266) );
NAND2_X1 U987 ( .A1(n1269), .A2(n1233), .ZN(n1267) );
XOR2_X1 U988 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U989 ( .A(n1189), .B(n1272), .Z(n1271) );
XNOR2_X1 U990 ( .A(KEYINPUT46), .B(n1237), .ZN(n1272) );
AND2_X1 U991 ( .A1(G224), .A2(n1074), .ZN(n1189) );
XNOR2_X1 U992 ( .A(n1184), .B(n1192), .ZN(n1270) );
INV_X1 U993 ( .A(n1264), .ZN(n1192) );
XOR2_X1 U994 ( .A(G128), .B(n1273), .Z(n1264) );
NAND3_X1 U995 ( .A1(n1274), .A2(n1275), .A3(n1112), .ZN(n1184) );
NAND3_X1 U996 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1112) );
NAND2_X1 U997 ( .A1(n1279), .A2(n1280), .ZN(n1275) );
INV_X1 U998 ( .A(KEYINPUT58), .ZN(n1280) );
XOR2_X1 U999 ( .A(n1281), .B(n1277), .Z(n1279) );
NOR2_X1 U1000 ( .A1(n1278), .A2(n1276), .ZN(n1281) );
INV_X1 U1001 ( .A(n1282), .ZN(n1278) );
NAND2_X1 U1002 ( .A1(KEYINPUT58), .A2(n1114), .ZN(n1274) );
NAND2_X1 U1003 ( .A1(n1283), .A2(n1284), .ZN(n1114) );
OR3_X1 U1004 ( .A1(n1276), .A2(n1277), .A3(n1282), .ZN(n1284) );
NAND2_X1 U1005 ( .A1(n1285), .A2(n1282), .ZN(n1283) );
XNOR2_X1 U1006 ( .A(n1286), .B(n1251), .ZN(n1282) );
XOR2_X1 U1007 ( .A(G113), .B(G119), .Z(n1251) );
XNOR2_X1 U1008 ( .A(G116), .B(KEYINPUT36), .ZN(n1286) );
XOR2_X1 U1009 ( .A(n1277), .B(n1276), .Z(n1285) );
XNOR2_X1 U1010 ( .A(n1287), .B(n1288), .ZN(n1276) );
NOR2_X1 U1011 ( .A1(KEYINPUT49), .A2(n1289), .ZN(n1288) );
XNOR2_X1 U1012 ( .A(G101), .B(KEYINPUT23), .ZN(n1289) );
XNOR2_X1 U1013 ( .A(G104), .B(G107), .ZN(n1287) );
XNOR2_X1 U1014 ( .A(G110), .B(n1290), .ZN(n1277) );
AND2_X1 U1015 ( .A1(n1054), .A2(n1053), .ZN(n1052) );
NAND2_X1 U1016 ( .A1(G221), .A2(n1232), .ZN(n1053) );
NAND2_X1 U1017 ( .A1(G234), .A2(n1233), .ZN(n1232) );
XOR2_X1 U1018 ( .A(n1070), .B(n1149), .Z(n1054) );
INV_X1 U1019 ( .A(G469), .ZN(n1149) );
NAND2_X1 U1020 ( .A1(n1291), .A2(n1233), .ZN(n1070) );
XOR2_X1 U1021 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U1022 ( .A(n1153), .B(n1148), .Z(n1293) );
XOR2_X1 U1023 ( .A(G140), .B(n1294), .Z(n1148) );
NOR2_X1 U1024 ( .A1(G953), .A2(n1075), .ZN(n1294) );
INV_X1 U1025 ( .A(G227), .ZN(n1075) );
XNOR2_X1 U1026 ( .A(n1295), .B(n1261), .ZN(n1153) );
INV_X1 U1027 ( .A(n1143), .ZN(n1261) );
XNOR2_X1 U1028 ( .A(n1296), .B(n1297), .ZN(n1143) );
XOR2_X1 U1029 ( .A(KEYINPUT48), .B(G137), .Z(n1297) );
XOR2_X1 U1030 ( .A(G134), .B(n1091), .Z(n1296) );
NAND3_X1 U1031 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1295) );
OR2_X1 U1032 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND3_X1 U1033 ( .A1(n1302), .A2(n1301), .A3(KEYINPUT1), .ZN(n1299) );
INV_X1 U1034 ( .A(G101), .ZN(n1301) );
NOR2_X1 U1035 ( .A1(KEYINPUT27), .A2(n1303), .ZN(n1302) );
NAND2_X1 U1036 ( .A1(n1303), .A2(n1304), .ZN(n1298) );
INV_X1 U1037 ( .A(KEYINPUT1), .ZN(n1304) );
NAND3_X1 U1038 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1303) );
OR2_X1 U1039 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND3_X1 U1040 ( .A1(n1309), .A2(n1308), .A3(KEYINPUT47), .ZN(n1306) );
NOR2_X1 U1041 ( .A1(G104), .A2(KEYINPUT44), .ZN(n1309) );
OR2_X1 U1042 ( .A1(n1310), .A2(KEYINPUT47), .ZN(n1305) );
XNOR2_X1 U1043 ( .A(n1311), .B(n1312), .ZN(n1292) );
NOR2_X1 U1044 ( .A1(KEYINPUT5), .A2(n1092), .ZN(n1312) );
XNOR2_X1 U1045 ( .A(n1313), .B(n1211), .ZN(n1092) );
INV_X1 U1046 ( .A(G128), .ZN(n1211) );
NAND2_X1 U1047 ( .A1(KEYINPUT40), .A2(n1273), .ZN(n1313) );
NOR2_X1 U1048 ( .A1(G110), .A2(KEYINPUT52), .ZN(n1311) );
NOR2_X1 U1049 ( .A1(n1203), .A2(n1205), .ZN(n1033) );
XOR2_X1 U1050 ( .A(n1314), .B(n1131), .Z(n1205) );
INV_X1 U1051 ( .A(G475), .ZN(n1131) );
NAND2_X1 U1052 ( .A1(n1129), .A2(n1233), .ZN(n1314) );
INV_X1 U1053 ( .A(G902), .ZN(n1233) );
XNOR2_X1 U1054 ( .A(n1315), .B(n1316), .ZN(n1129) );
XOR2_X1 U1055 ( .A(n1139), .B(n1317), .Z(n1316) );
XNOR2_X1 U1056 ( .A(n1318), .B(n1091), .ZN(n1317) );
XNOR2_X1 U1057 ( .A(G131), .B(KEYINPUT41), .ZN(n1091) );
NOR2_X1 U1058 ( .A1(n1255), .A2(n1319), .ZN(n1318) );
INV_X1 U1059 ( .A(G214), .ZN(n1319) );
NAND2_X1 U1060 ( .A1(n1320), .A2(n1074), .ZN(n1255) );
XNOR2_X1 U1061 ( .A(KEYINPUT33), .B(n1268), .ZN(n1320) );
INV_X1 U1062 ( .A(G237), .ZN(n1268) );
XOR2_X1 U1063 ( .A(G113), .B(n1273), .Z(n1139) );
XOR2_X1 U1064 ( .A(G146), .B(G143), .Z(n1273) );
XOR2_X1 U1065 ( .A(n1321), .B(n1322), .Z(n1315) );
XNOR2_X1 U1066 ( .A(KEYINPUT19), .B(n1290), .ZN(n1322) );
XNOR2_X1 U1067 ( .A(n1323), .B(n1310), .ZN(n1321) );
INV_X1 U1068 ( .A(G104), .ZN(n1310) );
NAND2_X1 U1069 ( .A1(n1324), .A2(n1097), .ZN(n1323) );
NAND2_X1 U1070 ( .A1(G140), .A2(n1237), .ZN(n1097) );
XOR2_X1 U1071 ( .A(KEYINPUT29), .B(n1325), .Z(n1324) );
NOR2_X1 U1072 ( .A1(G140), .A2(n1237), .ZN(n1325) );
INV_X1 U1073 ( .A(G125), .ZN(n1237) );
XOR2_X1 U1074 ( .A(G478), .B(n1326), .Z(n1203) );
NOR2_X1 U1075 ( .A1(G902), .A2(n1126), .ZN(n1326) );
XNOR2_X1 U1076 ( .A(n1327), .B(n1328), .ZN(n1126) );
XNOR2_X1 U1077 ( .A(n1308), .B(n1329), .ZN(n1328) );
XNOR2_X1 U1078 ( .A(n1290), .B(G116), .ZN(n1329) );
INV_X1 U1079 ( .A(G122), .ZN(n1290) );
INV_X1 U1080 ( .A(G107), .ZN(n1308) );
XOR2_X1 U1081 ( .A(n1330), .B(n1331), .Z(n1327) );
NOR2_X1 U1082 ( .A1(KEYINPUT4), .A2(n1332), .ZN(n1331) );
XOR2_X1 U1083 ( .A(G134), .B(n1333), .Z(n1332) );
NOR2_X1 U1084 ( .A1(KEYINPUT22), .A2(n1334), .ZN(n1333) );
NOR2_X1 U1085 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
XOR2_X1 U1086 ( .A(n1337), .B(KEYINPUT43), .Z(n1336) );
NAND2_X1 U1087 ( .A1(G128), .A2(n1200), .ZN(n1337) );
NOR2_X1 U1088 ( .A1(G128), .A2(n1200), .ZN(n1335) );
INV_X1 U1089 ( .A(G143), .ZN(n1200) );
NAND3_X1 U1090 ( .A1(G234), .A2(n1074), .A3(G217), .ZN(n1330) );
INV_X1 U1091 ( .A(G953), .ZN(n1074) );
NAND2_X1 U1092 ( .A1(KEYINPUT21), .A2(n1245), .ZN(n1226) );
INV_X1 U1093 ( .A(G110), .ZN(n1245) );
endmodule


