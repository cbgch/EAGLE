//Key = 1100000110011010100001110101101010011000111001011101101000011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356;

XOR2_X1 U743 ( .A(G107), .B(n1033), .Z(G9) );
NOR2_X1 U744 ( .A1(n1034), .A2(n1035), .ZN(G75) );
NOR4_X1 U745 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
NOR2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U747 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U748 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
INV_X1 U749 ( .A(n1046), .ZN(n1045) );
NOR2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(n1044) );
NOR2_X1 U751 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U754 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
XOR2_X1 U755 ( .A(KEYINPUT34), .B(n1057), .Z(n1056) );
NOR2_X1 U756 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR3_X1 U757 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1047) );
NOR3_X1 U758 ( .A1(n1054), .A2(n1063), .A3(n1064), .ZN(n1062) );
NOR2_X1 U759 ( .A1(KEYINPUT33), .A2(n1065), .ZN(n1064) );
NOR2_X1 U760 ( .A1(n1066), .A2(n1067), .ZN(n1061) );
AND2_X1 U761 ( .A1(n1068), .A2(KEYINPUT33), .ZN(n1066) );
NOR4_X1 U762 ( .A1(n1069), .A2(n1054), .A3(n1060), .A4(n1050), .ZN(n1042) );
INV_X1 U763 ( .A(n1067), .ZN(n1054) );
NOR2_X1 U764 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR2_X1 U765 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NAND4_X1 U766 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1036) );
NAND4_X1 U767 ( .A1(n1046), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1074) );
NOR3_X1 U768 ( .A1(n1081), .A2(n1082), .A3(n1041), .ZN(n1080) );
XNOR2_X1 U769 ( .A(KEYINPUT42), .B(n1060), .ZN(n1081) );
XNOR2_X1 U770 ( .A(KEYINPUT58), .B(n1083), .ZN(n1078) );
AND3_X1 U771 ( .A1(n1076), .A2(n1077), .A3(n1084), .ZN(n1034) );
NAND4_X1 U772 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1076) );
NOR4_X1 U773 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1088) );
XNOR2_X1 U774 ( .A(n1093), .B(n1094), .ZN(n1092) );
NAND2_X1 U775 ( .A1(KEYINPUT36), .A2(n1095), .ZN(n1093) );
NOR2_X1 U776 ( .A1(n1096), .A2(n1097), .ZN(n1091) );
XNOR2_X1 U777 ( .A(KEYINPUT22), .B(n1098), .ZN(n1097) );
INV_X1 U778 ( .A(n1099), .ZN(n1089) );
NOR3_X1 U779 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1087) );
NOR2_X1 U780 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U781 ( .A1(G475), .A2(n1105), .ZN(n1101) );
NOR2_X1 U782 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
AND2_X1 U783 ( .A1(n1104), .A2(KEYINPUT16), .ZN(n1107) );
NAND2_X1 U784 ( .A1(KEYINPUT28), .A2(n1108), .ZN(n1104) );
NOR2_X1 U785 ( .A1(KEYINPUT16), .A2(n1109), .ZN(n1106) );
XNOR2_X1 U786 ( .A(n1110), .B(n1111), .ZN(n1100) );
XOR2_X1 U787 ( .A(n1112), .B(n1113), .Z(G72) );
NOR2_X1 U788 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U789 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U790 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U791 ( .A(n1120), .B(G134), .Z(n1119) );
NAND2_X1 U792 ( .A1(KEYINPUT35), .A2(n1121), .ZN(n1120) );
NAND2_X1 U793 ( .A1(KEYINPUT32), .A2(n1122), .ZN(n1118) );
INV_X1 U794 ( .A(G131), .ZN(n1122) );
XNOR2_X1 U795 ( .A(n1123), .B(n1124), .ZN(n1116) );
NOR2_X1 U796 ( .A1(G900), .A2(n1077), .ZN(n1114) );
NAND2_X1 U797 ( .A1(n1125), .A2(n1126), .ZN(n1112) );
NAND2_X1 U798 ( .A1(n1039), .A2(n1077), .ZN(n1126) );
NAND2_X1 U799 ( .A1(G953), .A2(n1127), .ZN(n1125) );
NAND2_X1 U800 ( .A1(n1128), .A2(G900), .ZN(n1127) );
XNOR2_X1 U801 ( .A(G227), .B(KEYINPUT8), .ZN(n1128) );
XOR2_X1 U802 ( .A(n1129), .B(n1130), .Z(G69) );
NOR2_X1 U803 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR2_X1 U804 ( .A1(KEYINPUT41), .A2(n1133), .ZN(n1132) );
INV_X1 U805 ( .A(n1134), .ZN(n1133) );
NOR2_X1 U806 ( .A1(KEYINPUT53), .A2(n1134), .ZN(n1131) );
NAND2_X1 U807 ( .A1(n1077), .A2(n1135), .ZN(n1134) );
NAND2_X1 U808 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XNOR2_X1 U809 ( .A(KEYINPUT25), .B(n1075), .ZN(n1137) );
XOR2_X1 U810 ( .A(n1138), .B(n1139), .Z(n1129) );
NOR2_X1 U811 ( .A1(n1140), .A2(n1077), .ZN(n1139) );
AND2_X1 U812 ( .A1(G224), .A2(G898), .ZN(n1140) );
NAND2_X1 U813 ( .A1(n1141), .A2(n1142), .ZN(n1138) );
NAND2_X1 U814 ( .A1(G953), .A2(n1143), .ZN(n1142) );
XOR2_X1 U815 ( .A(n1144), .B(n1145), .Z(n1141) );
NOR2_X1 U816 ( .A1(KEYINPUT55), .A2(n1146), .ZN(n1144) );
NOR2_X1 U817 ( .A1(n1147), .A2(n1148), .ZN(G66) );
XNOR2_X1 U818 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR3_X1 U819 ( .A1(n1151), .A2(KEYINPUT17), .A3(n1095), .ZN(n1150) );
NOR2_X1 U820 ( .A1(n1147), .A2(n1152), .ZN(G63) );
XNOR2_X1 U821 ( .A(n1153), .B(n1154), .ZN(n1152) );
NOR2_X1 U822 ( .A1(n1155), .A2(n1151), .ZN(n1154) );
INV_X1 U823 ( .A(G478), .ZN(n1155) );
NOR2_X1 U824 ( .A1(n1147), .A2(n1156), .ZN(G60) );
XOR2_X1 U825 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U826 ( .A1(n1103), .A2(n1151), .ZN(n1157) );
INV_X1 U827 ( .A(G475), .ZN(n1103) );
XNOR2_X1 U828 ( .A(G104), .B(n1159), .ZN(G6) );
NOR2_X1 U829 ( .A1(n1147), .A2(n1160), .ZN(G57) );
XOR2_X1 U830 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U831 ( .A(n1163), .B(n1164), .ZN(n1161) );
NOR3_X1 U832 ( .A1(n1151), .A2(KEYINPUT6), .A3(n1165), .ZN(n1164) );
NOR2_X1 U833 ( .A1(KEYINPUT39), .A2(n1166), .ZN(n1163) );
XOR2_X1 U834 ( .A(G101), .B(n1167), .Z(n1166) );
NOR2_X1 U835 ( .A1(KEYINPUT56), .A2(n1168), .ZN(n1167) );
NOR2_X1 U836 ( .A1(n1147), .A2(n1169), .ZN(G54) );
XOR2_X1 U837 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U838 ( .A1(n1098), .A2(n1151), .ZN(n1171) );
NOR2_X1 U839 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
XOR2_X1 U840 ( .A(n1174), .B(KEYINPUT27), .Z(n1173) );
NAND2_X1 U841 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NOR2_X1 U842 ( .A1(n1176), .A2(n1175), .ZN(n1172) );
XOR2_X1 U843 ( .A(n1177), .B(n1178), .Z(n1175) );
NOR2_X1 U844 ( .A1(KEYINPUT61), .A2(n1179), .ZN(n1178) );
XNOR2_X1 U845 ( .A(G110), .B(n1180), .ZN(n1179) );
XNOR2_X1 U846 ( .A(n1181), .B(n1182), .ZN(n1176) );
NOR2_X1 U847 ( .A1(KEYINPUT44), .A2(n1183), .ZN(n1182) );
NOR3_X1 U848 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(G51) );
AND2_X1 U849 ( .A1(KEYINPUT14), .A2(n1147), .ZN(n1186) );
NOR2_X1 U850 ( .A1(n1077), .A2(G952), .ZN(n1147) );
NOR3_X1 U851 ( .A1(KEYINPUT14), .A2(n1077), .A3(n1084), .ZN(n1185) );
INV_X1 U852 ( .A(G952), .ZN(n1084) );
XOR2_X1 U853 ( .A(n1187), .B(n1188), .Z(n1184) );
XNOR2_X1 U854 ( .A(n1189), .B(n1190), .ZN(n1188) );
NAND2_X1 U855 ( .A1(n1191), .A2(KEYINPUT51), .ZN(n1189) );
XNOR2_X1 U856 ( .A(n1192), .B(n1193), .ZN(n1191) );
NAND2_X1 U857 ( .A1(KEYINPUT47), .A2(n1194), .ZN(n1192) );
INV_X1 U858 ( .A(n1195), .ZN(n1194) );
XOR2_X1 U859 ( .A(KEYINPUT11), .B(n1196), .Z(n1187) );
NOR2_X1 U860 ( .A1(n1197), .A2(n1151), .ZN(n1196) );
NAND2_X1 U861 ( .A1(n1198), .A2(n1199), .ZN(n1151) );
NAND3_X1 U862 ( .A1(n1200), .A2(n1075), .A3(n1136), .ZN(n1199) );
INV_X1 U863 ( .A(n1037), .ZN(n1136) );
NAND4_X1 U864 ( .A1(n1159), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1037) );
NOR4_X1 U865 ( .A1(n1033), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1203) );
INV_X1 U866 ( .A(n1207), .ZN(n1204) );
AND3_X1 U867 ( .A1(n1063), .A2(n1046), .A3(n1208), .ZN(n1033) );
NAND4_X1 U868 ( .A1(n1209), .A2(n1046), .A3(n1210), .A4(n1211), .ZN(n1202) );
XOR2_X1 U869 ( .A(KEYINPUT10), .B(n1212), .Z(n1210) );
NAND3_X1 U870 ( .A1(n1208), .A2(n1046), .A3(n1068), .ZN(n1159) );
NAND2_X1 U871 ( .A1(n1213), .A2(n1214), .ZN(n1075) );
XOR2_X1 U872 ( .A(KEYINPUT38), .B(n1063), .Z(n1214) );
INV_X1 U873 ( .A(n1039), .ZN(n1200) );
NAND4_X1 U874 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1039) );
NOR4_X1 U875 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1218) );
INV_X1 U876 ( .A(n1223), .ZN(n1219) );
NAND3_X1 U877 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1217) );
OR2_X1 U878 ( .A1(n1052), .A2(KEYINPUT13), .ZN(n1225) );
NAND2_X1 U879 ( .A1(KEYINPUT13), .A2(n1227), .ZN(n1224) );
NAND2_X1 U880 ( .A1(n1086), .A2(n1228), .ZN(n1227) );
NAND3_X1 U881 ( .A1(n1071), .A2(n1229), .A3(n1052), .ZN(n1215) );
NAND2_X1 U882 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND2_X1 U883 ( .A1(n1068), .A2(n1232), .ZN(n1231) );
XNOR2_X1 U884 ( .A(KEYINPUT45), .B(n1233), .ZN(n1232) );
NAND2_X1 U885 ( .A1(n1063), .A2(n1233), .ZN(n1230) );
XNOR2_X1 U886 ( .A(KEYINPUT2), .B(n1234), .ZN(n1198) );
XOR2_X1 U887 ( .A(G146), .B(n1222), .Z(G48) );
AND2_X1 U888 ( .A1(n1235), .A2(n1068), .ZN(n1222) );
NAND2_X1 U889 ( .A1(n1236), .A2(n1237), .ZN(G45) );
NAND2_X1 U890 ( .A1(n1221), .A2(n1238), .ZN(n1237) );
XOR2_X1 U891 ( .A(KEYINPUT59), .B(n1239), .Z(n1236) );
NOR2_X1 U892 ( .A1(n1221), .A2(n1238), .ZN(n1239) );
AND4_X1 U893 ( .A1(n1212), .A2(n1071), .A3(n1240), .A4(n1233), .ZN(n1221) );
XNOR2_X1 U894 ( .A(G140), .B(n1241), .ZN(G42) );
NAND2_X1 U895 ( .A1(n1052), .A2(n1226), .ZN(n1241) );
NAND2_X1 U896 ( .A1(n1242), .A2(n1243), .ZN(G39) );
NAND2_X1 U897 ( .A1(G137), .A2(n1216), .ZN(n1243) );
XOR2_X1 U898 ( .A(n1244), .B(KEYINPUT31), .Z(n1242) );
OR2_X1 U899 ( .A1(n1216), .A2(G137), .ZN(n1244) );
NAND4_X1 U900 ( .A1(n1052), .A2(n1245), .A3(n1073), .A4(n1233), .ZN(n1216) );
XNOR2_X1 U901 ( .A(G134), .B(n1246), .ZN(G36) );
NAND4_X1 U902 ( .A1(n1071), .A2(n1063), .A3(n1247), .A4(n1248), .ZN(n1246) );
NOR2_X1 U903 ( .A1(n1249), .A2(n1250), .ZN(n1247) );
XNOR2_X1 U904 ( .A(n1086), .B(KEYINPUT3), .ZN(n1250) );
INV_X1 U905 ( .A(n1060), .ZN(n1086) );
XNOR2_X1 U906 ( .A(G131), .B(n1251), .ZN(G33) );
NAND4_X1 U907 ( .A1(n1252), .A2(n1052), .A3(n1068), .A4(n1071), .ZN(n1251) );
INV_X1 U908 ( .A(n1065), .ZN(n1068) );
NOR2_X1 U909 ( .A1(n1060), .A2(n1228), .ZN(n1052) );
NAND2_X1 U910 ( .A1(n1253), .A2(n1059), .ZN(n1060) );
INV_X1 U911 ( .A(n1058), .ZN(n1253) );
XNOR2_X1 U912 ( .A(n1249), .B(KEYINPUT46), .ZN(n1252) );
XOR2_X1 U913 ( .A(n1220), .B(n1254), .Z(G30) );
NOR2_X1 U914 ( .A1(KEYINPUT43), .A2(n1255), .ZN(n1254) );
AND2_X1 U915 ( .A1(n1235), .A2(n1063), .ZN(n1220) );
AND4_X1 U916 ( .A1(n1240), .A2(n1256), .A3(n1073), .A4(n1233), .ZN(n1235) );
XNOR2_X1 U917 ( .A(G101), .B(n1201), .ZN(G3) );
NAND3_X1 U918 ( .A1(n1079), .A2(n1208), .A3(n1071), .ZN(n1201) );
NAND2_X1 U919 ( .A1(n1257), .A2(n1258), .ZN(G27) );
NAND2_X1 U920 ( .A1(G125), .A2(n1223), .ZN(n1258) );
XOR2_X1 U921 ( .A(KEYINPUT21), .B(n1259), .Z(n1257) );
NOR2_X1 U922 ( .A1(G125), .A2(n1223), .ZN(n1259) );
NAND2_X1 U923 ( .A1(n1226), .A2(n1209), .ZN(n1223) );
NOR4_X1 U924 ( .A1(n1073), .A2(n1065), .A3(n1072), .A4(n1249), .ZN(n1226) );
INV_X1 U925 ( .A(n1233), .ZN(n1249) );
NAND2_X1 U926 ( .A1(n1041), .A2(n1260), .ZN(n1233) );
NAND2_X1 U927 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
INV_X1 U928 ( .A(G900), .ZN(n1262) );
XOR2_X1 U929 ( .A(n1263), .B(n1264), .Z(G24) );
NAND2_X1 U930 ( .A1(KEYINPUT1), .A2(G122), .ZN(n1264) );
NAND4_X1 U931 ( .A1(n1212), .A2(n1209), .A3(n1046), .A4(n1265), .ZN(n1263) );
XNOR2_X1 U932 ( .A(KEYINPUT52), .B(n1211), .ZN(n1265) );
NOR2_X1 U933 ( .A1(n1073), .A2(n1256), .ZN(n1046) );
AND2_X1 U934 ( .A1(n1266), .A2(n1267), .ZN(n1212) );
XOR2_X1 U935 ( .A(G119), .B(n1206), .Z(G21) );
AND4_X1 U936 ( .A1(n1209), .A2(n1245), .A3(n1073), .A4(n1211), .ZN(n1206) );
XOR2_X1 U937 ( .A(G116), .B(n1268), .Z(G18) );
AND2_X1 U938 ( .A1(n1063), .A2(n1213), .ZN(n1268) );
INV_X1 U939 ( .A(n1269), .ZN(n1213) );
NOR2_X1 U940 ( .A1(n1267), .A2(n1270), .ZN(n1063) );
XOR2_X1 U941 ( .A(G113), .B(n1205), .Z(G15) );
NOR2_X1 U942 ( .A1(n1269), .A2(n1065), .ZN(n1205) );
NAND2_X1 U943 ( .A1(n1270), .A2(n1267), .ZN(n1065) );
NAND3_X1 U944 ( .A1(n1209), .A2(n1211), .A3(n1071), .ZN(n1269) );
NOR2_X1 U945 ( .A1(n1256), .A2(n1085), .ZN(n1071) );
INV_X1 U946 ( .A(n1072), .ZN(n1256) );
AND2_X1 U947 ( .A1(n1055), .A2(n1067), .ZN(n1209) );
NAND2_X1 U948 ( .A1(n1271), .A2(n1272), .ZN(n1067) );
OR3_X1 U949 ( .A1(n1083), .A2(n1090), .A3(KEYINPUT58), .ZN(n1272) );
INV_X1 U950 ( .A(n1082), .ZN(n1090) );
NAND2_X1 U951 ( .A1(KEYINPUT58), .A2(n1248), .ZN(n1271) );
XNOR2_X1 U952 ( .A(G110), .B(n1207), .ZN(G12) );
NAND3_X1 U953 ( .A1(n1085), .A2(n1208), .A3(n1245), .ZN(n1207) );
NOR2_X1 U954 ( .A1(n1050), .A2(n1072), .ZN(n1245) );
XNOR2_X1 U955 ( .A(n1094), .B(n1095), .ZN(n1072) );
NAND2_X1 U956 ( .A1(G217), .A2(n1273), .ZN(n1095) );
NAND2_X1 U957 ( .A1(n1274), .A2(n1234), .ZN(n1094) );
XNOR2_X1 U958 ( .A(KEYINPUT63), .B(n1275), .ZN(n1274) );
INV_X1 U959 ( .A(n1149), .ZN(n1275) );
XNOR2_X1 U960 ( .A(n1276), .B(n1277), .ZN(n1149) );
AND2_X1 U961 ( .A1(G221), .A2(n1278), .ZN(n1277) );
XNOR2_X1 U962 ( .A(n1279), .B(n1121), .ZN(n1276) );
NAND3_X1 U963 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1279) );
NAND2_X1 U964 ( .A1(KEYINPUT50), .A2(n1283), .ZN(n1282) );
NAND3_X1 U965 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1281) );
INV_X1 U966 ( .A(KEYINPUT50), .ZN(n1285) );
OR2_X1 U967 ( .A1(n1286), .A2(n1284), .ZN(n1280) );
NOR2_X1 U968 ( .A1(KEYINPUT29), .A2(n1283), .ZN(n1284) );
XNOR2_X1 U969 ( .A(n1124), .B(n1287), .ZN(n1283) );
XOR2_X1 U970 ( .A(G110), .B(n1288), .Z(n1286) );
XNOR2_X1 U971 ( .A(n1255), .B(G119), .ZN(n1288) );
INV_X1 U972 ( .A(n1079), .ZN(n1050) );
NOR2_X1 U973 ( .A1(n1267), .A2(n1266), .ZN(n1079) );
INV_X1 U974 ( .A(n1270), .ZN(n1266) );
XNOR2_X1 U975 ( .A(n1110), .B(n1289), .ZN(n1270) );
NOR2_X1 U976 ( .A1(KEYINPUT9), .A2(n1111), .ZN(n1289) );
XOR2_X1 U977 ( .A(G478), .B(KEYINPUT20), .Z(n1111) );
NAND2_X1 U978 ( .A1(n1153), .A2(n1234), .ZN(n1110) );
XNOR2_X1 U979 ( .A(n1290), .B(n1291), .ZN(n1153) );
XOR2_X1 U980 ( .A(n1292), .B(n1293), .Z(n1291) );
XNOR2_X1 U981 ( .A(n1294), .B(n1295), .ZN(n1293) );
NOR2_X1 U982 ( .A1(G122), .A2(KEYINPUT37), .ZN(n1295) );
NOR2_X1 U983 ( .A1(KEYINPUT57), .A2(n1296), .ZN(n1294) );
XNOR2_X1 U984 ( .A(G143), .B(KEYINPUT49), .ZN(n1296) );
NAND2_X1 U985 ( .A1(G217), .A2(n1278), .ZN(n1292) );
AND2_X1 U986 ( .A1(G234), .A2(n1077), .ZN(n1278) );
XOR2_X1 U987 ( .A(n1297), .B(n1298), .Z(n1290) );
XNOR2_X1 U988 ( .A(G134), .B(n1255), .ZN(n1298) );
INV_X1 U989 ( .A(G128), .ZN(n1255) );
XNOR2_X1 U990 ( .A(G116), .B(G107), .ZN(n1297) );
XNOR2_X1 U991 ( .A(n1108), .B(G475), .ZN(n1267) );
INV_X1 U992 ( .A(n1109), .ZN(n1108) );
NOR2_X1 U993 ( .A1(n1158), .A2(G902), .ZN(n1109) );
XNOR2_X1 U994 ( .A(n1299), .B(n1300), .ZN(n1158) );
XOR2_X1 U995 ( .A(n1287), .B(n1301), .Z(n1300) );
XNOR2_X1 U996 ( .A(n1302), .B(n1303), .ZN(n1301) );
NOR2_X1 U997 ( .A1(KEYINPUT19), .A2(n1124), .ZN(n1303) );
XNOR2_X1 U998 ( .A(G125), .B(n1180), .ZN(n1124) );
NAND2_X1 U999 ( .A1(KEYINPUT62), .A2(n1304), .ZN(n1302) );
XOR2_X1 U1000 ( .A(n1305), .B(n1306), .Z(n1299) );
XNOR2_X1 U1001 ( .A(G113), .B(n1307), .ZN(n1306) );
NAND2_X1 U1002 ( .A1(n1308), .A2(KEYINPUT54), .ZN(n1307) );
XNOR2_X1 U1003 ( .A(n1309), .B(n1238), .ZN(n1308) );
INV_X1 U1004 ( .A(G143), .ZN(n1238) );
NAND2_X1 U1005 ( .A1(n1310), .A2(G214), .ZN(n1309) );
XNOR2_X1 U1006 ( .A(G122), .B(G131), .ZN(n1305) );
AND2_X1 U1007 ( .A1(n1240), .A2(n1211), .ZN(n1208) );
NAND2_X1 U1008 ( .A1(n1041), .A2(n1311), .ZN(n1211) );
NAND2_X1 U1009 ( .A1(n1261), .A2(n1143), .ZN(n1311) );
INV_X1 U1010 ( .A(G898), .ZN(n1143) );
AND3_X1 U1011 ( .A1(n1312), .A2(n1313), .A3(G953), .ZN(n1261) );
XNOR2_X1 U1012 ( .A(KEYINPUT5), .B(n1234), .ZN(n1312) );
NAND3_X1 U1013 ( .A1(n1313), .A2(n1077), .A3(G952), .ZN(n1041) );
NAND2_X1 U1014 ( .A1(G237), .A2(G234), .ZN(n1313) );
AND2_X1 U1015 ( .A1(n1248), .A2(n1055), .ZN(n1240) );
AND2_X1 U1016 ( .A1(n1058), .A2(n1059), .ZN(n1055) );
NAND2_X1 U1017 ( .A1(G214), .A2(n1314), .ZN(n1059) );
XOR2_X1 U1018 ( .A(n1315), .B(n1197), .Z(n1058) );
NAND2_X1 U1019 ( .A1(G210), .A2(n1314), .ZN(n1197) );
NAND2_X1 U1020 ( .A1(n1316), .A2(n1234), .ZN(n1314) );
INV_X1 U1021 ( .A(G237), .ZN(n1316) );
NAND2_X1 U1022 ( .A1(n1317), .A2(n1234), .ZN(n1315) );
XNOR2_X1 U1023 ( .A(n1318), .B(n1319), .ZN(n1317) );
INV_X1 U1024 ( .A(n1190), .ZN(n1319) );
XOR2_X1 U1025 ( .A(n1145), .B(n1146), .Z(n1190) );
XNOR2_X1 U1026 ( .A(n1320), .B(n1321), .ZN(n1145) );
XNOR2_X1 U1027 ( .A(G122), .B(n1322), .ZN(n1321) );
INV_X1 U1028 ( .A(G110), .ZN(n1322) );
NAND2_X1 U1029 ( .A1(n1323), .A2(n1324), .ZN(n1320) );
NAND2_X1 U1030 ( .A1(G101), .A2(n1325), .ZN(n1324) );
XOR2_X1 U1031 ( .A(KEYINPUT48), .B(n1326), .Z(n1323) );
NOR2_X1 U1032 ( .A1(G101), .A2(n1325), .ZN(n1326) );
XNOR2_X1 U1033 ( .A(G107), .B(n1304), .ZN(n1325) );
INV_X1 U1034 ( .A(G104), .ZN(n1304) );
NAND2_X1 U1035 ( .A1(n1327), .A2(n1328), .ZN(n1318) );
NAND2_X1 U1036 ( .A1(n1193), .A2(n1195), .ZN(n1328) );
XOR2_X1 U1037 ( .A(KEYINPUT12), .B(n1329), .Z(n1327) );
NOR2_X1 U1038 ( .A1(n1193), .A2(n1195), .ZN(n1329) );
NAND2_X1 U1039 ( .A1(G224), .A2(n1077), .ZN(n1195) );
XOR2_X1 U1040 ( .A(n1330), .B(G125), .Z(n1193) );
INV_X1 U1041 ( .A(n1228), .ZN(n1248) );
NAND2_X1 U1042 ( .A1(n1082), .A2(n1083), .ZN(n1228) );
NAND2_X1 U1043 ( .A1(n1331), .A2(n1099), .ZN(n1083) );
NAND2_X1 U1044 ( .A1(n1096), .A2(n1098), .ZN(n1099) );
INV_X1 U1045 ( .A(G469), .ZN(n1098) );
NAND2_X1 U1046 ( .A1(G469), .A2(n1332), .ZN(n1331) );
XOR2_X1 U1047 ( .A(KEYINPUT23), .B(n1096), .Z(n1332) );
AND2_X1 U1048 ( .A1(n1333), .A2(n1234), .ZN(n1096) );
XOR2_X1 U1049 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1050 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1051 ( .A(n1177), .B(n1338), .Z(n1337) );
NOR2_X1 U1052 ( .A1(KEYINPUT4), .A2(n1183), .ZN(n1338) );
XNOR2_X1 U1053 ( .A(n1339), .B(n1340), .ZN(n1183) );
XOR2_X1 U1054 ( .A(KEYINPUT24), .B(G101), .Z(n1340) );
XOR2_X1 U1055 ( .A(n1123), .B(n1341), .Z(n1339) );
NOR2_X1 U1056 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
XOR2_X1 U1057 ( .A(KEYINPUT26), .B(n1344), .Z(n1343) );
NOR2_X1 U1058 ( .A1(G104), .A2(n1345), .ZN(n1344) );
AND2_X1 U1059 ( .A1(n1345), .A2(G104), .ZN(n1342) );
XOR2_X1 U1060 ( .A(G107), .B(KEYINPUT40), .Z(n1345) );
XOR2_X1 U1061 ( .A(n1346), .B(n1347), .Z(n1123) );
NAND2_X1 U1062 ( .A1(KEYINPUT7), .A2(G128), .ZN(n1346) );
NAND2_X1 U1063 ( .A1(G227), .A2(n1077), .ZN(n1177) );
INV_X1 U1064 ( .A(G953), .ZN(n1077) );
NAND2_X1 U1065 ( .A1(KEYINPUT0), .A2(G110), .ZN(n1336) );
XNOR2_X1 U1066 ( .A(n1181), .B(n1180), .ZN(n1334) );
XOR2_X1 U1067 ( .A(G140), .B(KEYINPUT15), .Z(n1180) );
NAND2_X1 U1068 ( .A1(G221), .A2(n1273), .ZN(n1082) );
NAND2_X1 U1069 ( .A1(G234), .A2(n1234), .ZN(n1273) );
INV_X1 U1070 ( .A(n1073), .ZN(n1085) );
XOR2_X1 U1071 ( .A(n1348), .B(n1165), .Z(n1073) );
INV_X1 U1072 ( .A(G472), .ZN(n1165) );
NAND2_X1 U1073 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
XNOR2_X1 U1074 ( .A(KEYINPUT30), .B(n1234), .ZN(n1350) );
INV_X1 U1075 ( .A(G902), .ZN(n1234) );
XOR2_X1 U1076 ( .A(n1351), .B(n1352), .Z(n1349) );
XOR2_X1 U1077 ( .A(KEYINPUT18), .B(G101), .Z(n1352) );
XOR2_X1 U1078 ( .A(n1162), .B(n1168), .Z(n1351) );
NAND2_X1 U1079 ( .A1(n1310), .A2(G210), .ZN(n1168) );
NOR2_X1 U1080 ( .A1(G953), .A2(G237), .ZN(n1310) );
XNOR2_X1 U1081 ( .A(n1330), .B(n1353), .ZN(n1162) );
XNOR2_X1 U1082 ( .A(n1146), .B(n1354), .ZN(n1353) );
INV_X1 U1083 ( .A(n1181), .ZN(n1354) );
XOR2_X1 U1084 ( .A(G131), .B(n1355), .Z(n1181) );
XNOR2_X1 U1085 ( .A(n1121), .B(G134), .ZN(n1355) );
INV_X1 U1086 ( .A(G137), .ZN(n1121) );
XOR2_X1 U1087 ( .A(G113), .B(n1356), .Z(n1146) );
XOR2_X1 U1088 ( .A(G119), .B(G116), .Z(n1356) );
XNOR2_X1 U1089 ( .A(n1347), .B(G128), .ZN(n1330) );
XOR2_X1 U1090 ( .A(G143), .B(n1287), .Z(n1347) );
XOR2_X1 U1091 ( .A(G146), .B(KEYINPUT60), .Z(n1287) );
endmodule


