//Key = 1000010100011001000101110010011101101111000100010111100110111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290;

XNOR2_X1 U717 ( .A(G107), .B(n984), .ZN(G9) );
NOR2_X1 U718 ( .A1(n985), .A2(KEYINPUT18), .ZN(n984) );
NOR2_X1 U719 ( .A1(n986), .A2(n987), .ZN(G75) );
NOR3_X1 U720 ( .A1(n988), .A2(G953), .A3(n989), .ZN(n987) );
INV_X1 U721 ( .A(n990), .ZN(n989) );
XNOR2_X1 U722 ( .A(KEYINPUT53), .B(n991), .ZN(n988) );
NOR4_X1 U723 ( .A1(n992), .A2(n993), .A3(n994), .A4(n991), .ZN(n986) );
INV_X1 U724 ( .A(G952), .ZN(n991) );
XOR2_X1 U725 ( .A(n995), .B(KEYINPUT46), .Z(n994) );
NAND2_X1 U726 ( .A1(n996), .A2(n997), .ZN(n995) );
NAND3_X1 U727 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n997) );
NAND2_X1 U728 ( .A1(n1001), .A2(n1002), .ZN(n996) );
NAND2_X1 U729 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND2_X1 U730 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND2_X1 U731 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NAND3_X1 U732 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1008) );
XNOR2_X1 U733 ( .A(n998), .B(KEYINPUT61), .ZN(n1011) );
NAND3_X1 U734 ( .A1(n998), .A2(n1012), .A3(n1013), .ZN(n1007) );
NAND2_X1 U735 ( .A1(n1014), .A2(n1000), .ZN(n1003) );
NAND4_X1 U736 ( .A1(n990), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n992) );
NAND3_X1 U737 ( .A1(n1018), .A2(n1001), .A3(n1000), .ZN(n1016) );
NAND2_X1 U738 ( .A1(n998), .A2(n1019), .ZN(n1015) );
NAND2_X1 U739 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND3_X1 U740 ( .A1(n1022), .A2(n1006), .A3(n1001), .ZN(n1021) );
NAND2_X1 U741 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND3_X1 U742 ( .A1(n1025), .A2(n1013), .A3(n1026), .ZN(n1024) );
NAND2_X1 U743 ( .A1(n1010), .A2(n1027), .ZN(n1023) );
NAND3_X1 U744 ( .A1(n1028), .A2(n1000), .A3(n1029), .ZN(n1020) );
AND3_X1 U745 ( .A1(n1010), .A2(n1006), .A3(n1013), .ZN(n1000) );
NAND4_X1 U746 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n990) );
AND4_X1 U747 ( .A1(n1034), .A2(n1035), .A3(n1010), .A4(n1001), .ZN(n1033) );
INV_X1 U748 ( .A(n1036), .ZN(n1001) );
XNOR2_X1 U749 ( .A(n1037), .B(n1038), .ZN(n1035) );
NOR2_X1 U750 ( .A1(KEYINPUT24), .A2(n1039), .ZN(n1038) );
XOR2_X1 U751 ( .A(n1040), .B(KEYINPUT33), .Z(n1039) );
NOR2_X1 U752 ( .A1(n1041), .A2(n1042), .ZN(n1032) );
AND2_X1 U753 ( .A1(n1043), .A2(KEYINPUT20), .ZN(n1042) );
NOR3_X1 U754 ( .A1(KEYINPUT20), .A2(n1044), .A3(n1043), .ZN(n1041) );
XNOR2_X1 U755 ( .A(n1045), .B(n1046), .ZN(n1031) );
XNOR2_X1 U756 ( .A(n1047), .B(KEYINPUT62), .ZN(n1030) );
XOR2_X1 U757 ( .A(n1048), .B(n1049), .Z(G72) );
NOR3_X1 U758 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
NOR2_X1 U759 ( .A1(G953), .A2(n1053), .ZN(n1052) );
NOR2_X1 U760 ( .A1(G227), .A2(n1017), .ZN(n1051) );
NAND2_X1 U761 ( .A1(n1054), .A2(n1055), .ZN(n1048) );
INV_X1 U762 ( .A(n1050), .ZN(n1055) );
XOR2_X1 U763 ( .A(n1056), .B(n1057), .Z(n1054) );
NAND2_X1 U764 ( .A1(KEYINPUT31), .A2(n1058), .ZN(n1056) );
XNOR2_X1 U765 ( .A(n1059), .B(n1060), .ZN(n1058) );
NAND2_X1 U766 ( .A1(KEYINPUT37), .A2(n1061), .ZN(n1059) );
XOR2_X1 U767 ( .A(n1062), .B(n1063), .Z(G69) );
NOR3_X1 U768 ( .A1(n1017), .A2(KEYINPUT17), .A3(n1064), .ZN(n1063) );
AND2_X1 U769 ( .A1(G224), .A2(G898), .ZN(n1064) );
XOR2_X1 U770 ( .A(n1065), .B(n1066), .Z(n1062) );
NOR2_X1 U771 ( .A1(n1067), .A2(G953), .ZN(n1066) );
NAND2_X1 U772 ( .A1(KEYINPUT43), .A2(n1068), .ZN(n1065) );
NAND2_X1 U773 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
INV_X1 U774 ( .A(n1071), .ZN(n1070) );
XOR2_X1 U775 ( .A(n1072), .B(n1073), .Z(n1069) );
NOR2_X1 U776 ( .A1(n1074), .A2(n1075), .ZN(G66) );
XOR2_X1 U777 ( .A(n1076), .B(n1077), .Z(n1075) );
XOR2_X1 U778 ( .A(KEYINPUT6), .B(n1078), .Z(n1077) );
NOR2_X1 U779 ( .A1(n1043), .A2(n1079), .ZN(n1078) );
NOR2_X1 U780 ( .A1(n1074), .A2(n1080), .ZN(G63) );
XOR2_X1 U781 ( .A(n1081), .B(n1082), .Z(n1080) );
NOR2_X1 U782 ( .A1(n1083), .A2(n1079), .ZN(n1082) );
INV_X1 U783 ( .A(G478), .ZN(n1083) );
NOR2_X1 U784 ( .A1(n1074), .A2(n1084), .ZN(G60) );
XNOR2_X1 U785 ( .A(n1085), .B(n1086), .ZN(n1084) );
NOR2_X1 U786 ( .A1(n1046), .A2(n1079), .ZN(n1086) );
INV_X1 U787 ( .A(G475), .ZN(n1046) );
XNOR2_X1 U788 ( .A(G104), .B(n1087), .ZN(G6) );
NOR2_X1 U789 ( .A1(n1088), .A2(n1089), .ZN(G57) );
XOR2_X1 U790 ( .A(n1090), .B(n1091), .Z(n1089) );
XOR2_X1 U791 ( .A(G101), .B(n1092), .Z(n1091) );
NOR2_X1 U792 ( .A1(n1037), .A2(n1079), .ZN(n1092) );
NOR2_X1 U793 ( .A1(G952), .A2(n1093), .ZN(n1088) );
XNOR2_X1 U794 ( .A(KEYINPUT22), .B(n1017), .ZN(n1093) );
NOR2_X1 U795 ( .A1(n1074), .A2(n1094), .ZN(G54) );
XOR2_X1 U796 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U797 ( .A1(n1097), .A2(n1079), .ZN(n1096) );
NOR2_X1 U798 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
XOR2_X1 U799 ( .A(n1100), .B(KEYINPUT15), .Z(n1099) );
NAND2_X1 U800 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U801 ( .A1(n1101), .A2(n1103), .ZN(n1098) );
XNOR2_X1 U802 ( .A(n1102), .B(KEYINPUT11), .ZN(n1103) );
AND2_X1 U803 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NAND2_X1 U804 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U805 ( .A(KEYINPUT63), .B(n1108), .Z(n1104) );
NOR2_X1 U806 ( .A1(n1107), .A2(n1106), .ZN(n1108) );
AND2_X1 U807 ( .A1(n1109), .A2(n1110), .ZN(n1106) );
NAND2_X1 U808 ( .A1(G140), .A2(n1111), .ZN(n1110) );
NAND2_X1 U809 ( .A1(n1112), .A2(n1113), .ZN(n1109) );
XNOR2_X1 U810 ( .A(KEYINPUT1), .B(n1111), .ZN(n1112) );
AND2_X1 U811 ( .A1(n1114), .A2(n1115), .ZN(n1101) );
NAND2_X1 U812 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XNOR2_X1 U813 ( .A(n1118), .B(n1060), .ZN(n1117) );
NAND2_X1 U814 ( .A1(n1119), .A2(n1120), .ZN(n1114) );
XNOR2_X1 U815 ( .A(n1118), .B(n1121), .ZN(n1120) );
NAND2_X1 U816 ( .A1(n1122), .A2(KEYINPUT21), .ZN(n1118) );
XNOR2_X1 U817 ( .A(n1123), .B(KEYINPUT35), .ZN(n1122) );
XOR2_X1 U818 ( .A(n1116), .B(KEYINPUT30), .Z(n1119) );
NOR2_X1 U819 ( .A1(n1074), .A2(n1124), .ZN(G51) );
XOR2_X1 U820 ( .A(n1125), .B(n1126), .Z(n1124) );
XNOR2_X1 U821 ( .A(n1127), .B(n1128), .ZN(n1126) );
XOR2_X1 U822 ( .A(n1129), .B(n1130), .Z(n1125) );
NOR2_X1 U823 ( .A1(n1131), .A2(n1079), .ZN(n1130) );
NAND2_X1 U824 ( .A1(n1132), .A2(n993), .ZN(n1079) );
NAND2_X1 U825 ( .A1(n1067), .A2(n1053), .ZN(n993) );
AND2_X1 U826 ( .A1(n1133), .A2(n1134), .ZN(n1053) );
NOR4_X1 U827 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1134) );
INV_X1 U828 ( .A(n1139), .ZN(n1138) );
NOR4_X1 U829 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1133) );
NOR3_X1 U830 ( .A1(n1144), .A2(n1145), .A3(n1036), .ZN(n1143) );
NOR3_X1 U831 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1142) );
XNOR2_X1 U832 ( .A(n1012), .B(KEYINPUT45), .ZN(n1147) );
XNOR2_X1 U833 ( .A(KEYINPUT58), .B(n1036), .ZN(n1146) );
INV_X1 U834 ( .A(n1149), .ZN(n1140) );
AND4_X1 U835 ( .A1(n1087), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1067) );
NOR4_X1 U836 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n985), .ZN(n1152) );
AND3_X1 U837 ( .A1(n1156), .A2(n998), .A3(n1027), .ZN(n985) );
NAND3_X1 U838 ( .A1(n1157), .A2(n1158), .A3(n1156), .ZN(n1151) );
NAND2_X1 U839 ( .A1(n1159), .A2(n1145), .ZN(n1158) );
NAND2_X1 U840 ( .A1(KEYINPUT9), .A2(n1014), .ZN(n1159) );
NAND3_X1 U841 ( .A1(n1160), .A2(n1161), .A3(n1013), .ZN(n1157) );
OR2_X1 U842 ( .A1(n1162), .A2(KEYINPUT9), .ZN(n1160) );
NAND3_X1 U843 ( .A1(n1156), .A2(n998), .A3(n1009), .ZN(n1087) );
INV_X1 U844 ( .A(n1163), .ZN(n1156) );
XNOR2_X1 U845 ( .A(KEYINPUT4), .B(n1164), .ZN(n1132) );
NAND2_X1 U846 ( .A1(KEYINPUT59), .A2(G125), .ZN(n1129) );
NOR2_X1 U847 ( .A1(n1017), .A2(G952), .ZN(n1074) );
XOR2_X1 U848 ( .A(n1141), .B(n1165), .Z(G48) );
NOR2_X1 U849 ( .A1(KEYINPUT57), .A2(n1166), .ZN(n1165) );
AND3_X1 U850 ( .A1(n1009), .A2(n999), .A3(n1167), .ZN(n1141) );
XNOR2_X1 U851 ( .A(G143), .B(n1149), .ZN(G45) );
NAND4_X1 U852 ( .A1(n1047), .A2(n1168), .A3(n999), .A4(n1169), .ZN(n1149) );
NOR3_X1 U853 ( .A1(n1162), .A2(n1170), .A3(n1171), .ZN(n1169) );
XNOR2_X1 U854 ( .A(n1113), .B(n1172), .ZN(G42) );
AND2_X1 U855 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U856 ( .A(G137), .B(n1175), .Z(G39) );
NOR4_X1 U857 ( .A1(KEYINPUT16), .A2(n1145), .A3(n1036), .A4(n1144), .ZN(n1175) );
XNOR2_X1 U858 ( .A(n1137), .B(n1176), .ZN(G36) );
NAND2_X1 U859 ( .A1(KEYINPUT36), .A2(G134), .ZN(n1176) );
AND4_X1 U860 ( .A1(n1174), .A2(n1014), .A3(n1027), .A4(n1168), .ZN(n1137) );
XNOR2_X1 U861 ( .A(G131), .B(n1139), .ZN(G33) );
NAND4_X1 U862 ( .A1(n1174), .A2(n1009), .A3(n1014), .A4(n1168), .ZN(n1139) );
NOR2_X1 U863 ( .A1(n1036), .A2(n1170), .ZN(n1174) );
INV_X1 U864 ( .A(n1012), .ZN(n1170) );
NAND2_X1 U865 ( .A1(n1028), .A2(n1177), .ZN(n1036) );
XOR2_X1 U866 ( .A(G128), .B(n1136), .Z(G30) );
AND3_X1 U867 ( .A1(n1027), .A2(n999), .A3(n1167), .ZN(n1136) );
INV_X1 U868 ( .A(n1144), .ZN(n1167) );
NAND4_X1 U869 ( .A1(n1012), .A2(n1178), .A3(n1168), .A4(n1179), .ZN(n1144) );
XOR2_X1 U870 ( .A(G101), .B(n1180), .Z(G3) );
NOR3_X1 U871 ( .A1(n1162), .A2(n1163), .A3(n1145), .ZN(n1180) );
XOR2_X1 U872 ( .A(G125), .B(n1135), .Z(G27) );
AND3_X1 U873 ( .A1(n1010), .A2(n999), .A3(n1173), .ZN(n1135) );
INV_X1 U874 ( .A(n1148), .ZN(n1173) );
NAND3_X1 U875 ( .A1(n1018), .A2(n1168), .A3(n1009), .ZN(n1148) );
NAND2_X1 U876 ( .A1(n1181), .A2(n1182), .ZN(n1168) );
XOR2_X1 U877 ( .A(n1183), .B(KEYINPUT32), .Z(n1181) );
NAND3_X1 U878 ( .A1(G902), .A2(n1006), .A3(n1050), .ZN(n1183) );
NOR2_X1 U879 ( .A1(G900), .A2(n1017), .ZN(n1050) );
INV_X1 U880 ( .A(n1161), .ZN(n1018) );
XNOR2_X1 U881 ( .A(G122), .B(n1184), .ZN(G24) );
NAND2_X1 U882 ( .A1(KEYINPUT51), .A2(n1155), .ZN(n1184) );
AND4_X1 U883 ( .A1(n1185), .A2(n1186), .A3(n998), .A4(n1047), .ZN(n1155) );
AND2_X1 U884 ( .A1(n1187), .A2(n1188), .ZN(n998) );
XOR2_X1 U885 ( .A(G119), .B(n1189), .Z(G21) );
NOR2_X1 U886 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U887 ( .A1(KEYINPUT3), .A2(n1192), .ZN(n1191) );
INV_X1 U888 ( .A(n1150), .ZN(n1192) );
NOR2_X1 U889 ( .A1(KEYINPUT12), .A2(n1150), .ZN(n1190) );
NAND4_X1 U890 ( .A1(n1186), .A2(n1013), .A3(n1178), .A4(n1179), .ZN(n1150) );
XNOR2_X1 U891 ( .A(n1193), .B(n1154), .ZN(G18) );
AND3_X1 U892 ( .A1(n1014), .A2(n1027), .A3(n1186), .ZN(n1154) );
NOR2_X1 U893 ( .A1(n1185), .A2(n1194), .ZN(n1027) );
INV_X1 U894 ( .A(n1047), .ZN(n1194) );
XOR2_X1 U895 ( .A(G113), .B(n1153), .Z(G15) );
AND3_X1 U896 ( .A1(n1009), .A2(n1014), .A3(n1186), .ZN(n1153) );
AND3_X1 U897 ( .A1(n999), .A2(n1195), .A3(n1010), .ZN(n1186) );
NOR2_X1 U898 ( .A1(n1196), .A2(n1026), .ZN(n1010) );
INV_X1 U899 ( .A(n1162), .ZN(n1014) );
NAND2_X1 U900 ( .A1(n1187), .A2(n1178), .ZN(n1162) );
INV_X1 U901 ( .A(n1179), .ZN(n1187) );
NOR2_X1 U902 ( .A1(n1171), .A2(n1047), .ZN(n1009) );
XOR2_X1 U903 ( .A(n1197), .B(n1198), .Z(G12) );
NOR4_X1 U904 ( .A1(KEYINPUT2), .A2(n1163), .A3(n1145), .A4(n1161), .ZN(n1198) );
NAND2_X1 U905 ( .A1(n1188), .A2(n1179), .ZN(n1161) );
NAND2_X1 U906 ( .A1(n1199), .A2(n1034), .ZN(n1179) );
NAND2_X1 U907 ( .A1(n1044), .A2(n1043), .ZN(n1034) );
OR2_X1 U908 ( .A1(n1043), .A2(n1044), .ZN(n1199) );
NOR2_X1 U909 ( .A1(n1076), .A2(n1200), .ZN(n1044) );
XNOR2_X1 U910 ( .A(n1201), .B(n1202), .ZN(n1076) );
XOR2_X1 U911 ( .A(n1057), .B(n1203), .Z(n1202) );
XOR2_X1 U912 ( .A(n1204), .B(n1205), .Z(n1203) );
AND3_X1 U913 ( .A1(G221), .A2(n1017), .A3(G234), .ZN(n1204) );
XOR2_X1 U914 ( .A(n1206), .B(n1207), .Z(n1201) );
XOR2_X1 U915 ( .A(KEYINPUT19), .B(G137), .Z(n1207) );
XNOR2_X1 U916 ( .A(n1208), .B(n1111), .ZN(n1206) );
INV_X1 U917 ( .A(G110), .ZN(n1111) );
NAND2_X1 U918 ( .A1(n1209), .A2(KEYINPUT38), .ZN(n1208) );
XNOR2_X1 U919 ( .A(G119), .B(n1210), .ZN(n1209) );
NOR2_X1 U920 ( .A1(G128), .A2(KEYINPUT8), .ZN(n1210) );
NAND2_X1 U921 ( .A1(G217), .A2(n1211), .ZN(n1043) );
XOR2_X1 U922 ( .A(n1178), .B(KEYINPUT49), .Z(n1188) );
XOR2_X1 U923 ( .A(n1040), .B(n1037), .Z(n1178) );
INV_X1 U924 ( .A(G472), .ZN(n1037) );
NAND2_X1 U925 ( .A1(n1212), .A2(n1213), .ZN(n1040) );
XOR2_X1 U926 ( .A(n1214), .B(n1090), .Z(n1212) );
XNOR2_X1 U927 ( .A(n1215), .B(n1216), .ZN(n1090) );
XOR2_X1 U928 ( .A(n1127), .B(n1217), .Z(n1216) );
XOR2_X1 U929 ( .A(n1218), .B(n1219), .Z(n1217) );
NAND2_X1 U930 ( .A1(G210), .A2(n1220), .ZN(n1219) );
NAND2_X1 U931 ( .A1(KEYINPUT26), .A2(G113), .ZN(n1218) );
XOR2_X1 U932 ( .A(n1116), .B(n1221), .Z(n1215) );
NOR2_X1 U933 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NOR3_X1 U934 ( .A1(n1224), .A2(G119), .A3(n1193), .ZN(n1223) );
INV_X1 U935 ( .A(KEYINPUT41), .ZN(n1224) );
NOR2_X1 U936 ( .A1(KEYINPUT41), .A2(n1225), .ZN(n1222) );
NOR2_X1 U937 ( .A1(KEYINPUT40), .A2(n1226), .ZN(n1214) );
XNOR2_X1 U938 ( .A(G101), .B(KEYINPUT60), .ZN(n1226) );
INV_X1 U939 ( .A(n1013), .ZN(n1145) );
NOR2_X1 U940 ( .A1(n1047), .A2(n1185), .ZN(n1013) );
INV_X1 U941 ( .A(n1171), .ZN(n1185) );
XNOR2_X1 U942 ( .A(n1045), .B(n1227), .ZN(n1171) );
NOR2_X1 U943 ( .A1(G475), .A2(KEYINPUT14), .ZN(n1227) );
NAND2_X1 U944 ( .A1(n1085), .A2(n1213), .ZN(n1045) );
XNOR2_X1 U945 ( .A(n1228), .B(n1229), .ZN(n1085) );
XOR2_X1 U946 ( .A(n1230), .B(n1231), .Z(n1229) );
NAND2_X1 U947 ( .A1(n1232), .A2(KEYINPUT34), .ZN(n1231) );
XNOR2_X1 U948 ( .A(G104), .B(n1233), .ZN(n1232) );
NAND2_X1 U949 ( .A1(n1234), .A2(n1235), .ZN(n1230) );
OR2_X1 U950 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
XOR2_X1 U951 ( .A(n1238), .B(KEYINPUT10), .Z(n1234) );
NAND2_X1 U952 ( .A1(n1237), .A2(n1236), .ZN(n1238) );
INV_X1 U953 ( .A(G131), .ZN(n1236) );
XOR2_X1 U954 ( .A(n1239), .B(n1240), .Z(n1237) );
NAND2_X1 U955 ( .A1(G214), .A2(n1220), .ZN(n1239) );
NOR2_X1 U956 ( .A1(G953), .A2(G237), .ZN(n1220) );
XOR2_X1 U957 ( .A(n1241), .B(n1057), .Z(n1228) );
XOR2_X1 U958 ( .A(G125), .B(G140), .Z(n1057) );
NAND2_X1 U959 ( .A1(KEYINPUT56), .A2(n1205), .ZN(n1241) );
XNOR2_X1 U960 ( .A(n1166), .B(KEYINPUT13), .ZN(n1205) );
XOR2_X1 U961 ( .A(G478), .B(n1242), .Z(n1047) );
NOR2_X1 U962 ( .A1(n1081), .A2(n1200), .ZN(n1242) );
INV_X1 U963 ( .A(n1213), .ZN(n1200) );
AND2_X1 U964 ( .A1(n1243), .A2(n1244), .ZN(n1081) );
NAND2_X1 U965 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND3_X1 U966 ( .A1(G217), .A2(n1017), .A3(G234), .ZN(n1246) );
XOR2_X1 U967 ( .A(KEYINPUT50), .B(n1247), .Z(n1243) );
AND4_X1 U968 ( .A1(n1017), .A2(G217), .A3(G234), .A4(n1248), .ZN(n1247) );
XNOR2_X1 U969 ( .A(KEYINPUT25), .B(n1245), .ZN(n1248) );
XNOR2_X1 U970 ( .A(n1249), .B(n1250), .ZN(n1245) );
XNOR2_X1 U971 ( .A(n1251), .B(n1252), .ZN(n1250) );
XNOR2_X1 U972 ( .A(G107), .B(n1253), .ZN(n1252) );
NOR2_X1 U973 ( .A1(G116), .A2(KEYINPUT42), .ZN(n1253) );
XNOR2_X1 U974 ( .A(G122), .B(n1254), .ZN(n1249) );
XOR2_X1 U975 ( .A(KEYINPUT55), .B(G134), .Z(n1254) );
NAND3_X1 U976 ( .A1(n999), .A2(n1195), .A3(n1012), .ZN(n1163) );
NOR2_X1 U977 ( .A1(n1025), .A2(n1026), .ZN(n1012) );
AND2_X1 U978 ( .A1(G221), .A2(n1211), .ZN(n1026) );
NAND2_X1 U979 ( .A1(G234), .A2(n1164), .ZN(n1211) );
INV_X1 U980 ( .A(n1196), .ZN(n1025) );
XOR2_X1 U981 ( .A(n1255), .B(n1097), .Z(n1196) );
INV_X1 U982 ( .A(G469), .ZN(n1097) );
NAND2_X1 U983 ( .A1(n1256), .A2(n1213), .ZN(n1255) );
XOR2_X1 U984 ( .A(n1257), .B(n1258), .Z(n1256) );
XNOR2_X1 U985 ( .A(n1259), .B(n1121), .ZN(n1258) );
INV_X1 U986 ( .A(n1060), .ZN(n1121) );
XNOR2_X1 U987 ( .A(n1260), .B(G128), .ZN(n1060) );
NAND3_X1 U988 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1260) );
NAND2_X1 U989 ( .A1(G143), .A2(n1166), .ZN(n1263) );
NAND2_X1 U990 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
INV_X1 U991 ( .A(KEYINPUT52), .ZN(n1265) );
NAND2_X1 U992 ( .A1(n1266), .A2(G146), .ZN(n1264) );
XNOR2_X1 U993 ( .A(KEYINPUT48), .B(G143), .ZN(n1266) );
NAND2_X1 U994 ( .A1(KEYINPUT52), .A2(n1267), .ZN(n1261) );
NAND2_X1 U995 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
OR3_X1 U996 ( .A1(n1166), .A2(G143), .A3(KEYINPUT48), .ZN(n1269) );
INV_X1 U997 ( .A(G146), .ZN(n1166) );
NAND2_X1 U998 ( .A1(KEYINPUT48), .A2(G143), .ZN(n1268) );
XNOR2_X1 U999 ( .A(n1116), .B(n1270), .ZN(n1259) );
INV_X1 U1000 ( .A(n1123), .ZN(n1270) );
XOR2_X1 U1001 ( .A(n1271), .B(n1272), .Z(n1123) );
XOR2_X1 U1002 ( .A(n1061), .B(KEYINPUT39), .Z(n1116) );
XNOR2_X1 U1003 ( .A(G131), .B(n1273), .ZN(n1061) );
XOR2_X1 U1004 ( .A(G137), .B(G134), .Z(n1273) );
XNOR2_X1 U1005 ( .A(n1107), .B(n1274), .ZN(n1257) );
XNOR2_X1 U1006 ( .A(n1113), .B(G110), .ZN(n1274) );
INV_X1 U1007 ( .A(G140), .ZN(n1113) );
AND2_X1 U1008 ( .A1(G227), .A2(n1017), .ZN(n1107) );
NAND2_X1 U1009 ( .A1(n1275), .A2(n1276), .ZN(n1195) );
NAND3_X1 U1010 ( .A1(G902), .A2(n1006), .A3(n1071), .ZN(n1276) );
NOR2_X1 U1011 ( .A1(n1017), .A2(G898), .ZN(n1071) );
XNOR2_X1 U1012 ( .A(KEYINPUT47), .B(n1182), .ZN(n1275) );
NAND3_X1 U1013 ( .A1(G952), .A2(n1017), .A3(n1277), .ZN(n1182) );
XOR2_X1 U1014 ( .A(n1006), .B(KEYINPUT54), .Z(n1277) );
NAND2_X1 U1015 ( .A1(G237), .A2(G234), .ZN(n1006) );
NOR2_X1 U1016 ( .A1(n1028), .A2(n1029), .ZN(n999) );
INV_X1 U1017 ( .A(n1177), .ZN(n1029) );
NAND2_X1 U1018 ( .A1(G214), .A2(n1278), .ZN(n1177) );
XNOR2_X1 U1019 ( .A(n1279), .B(n1131), .ZN(n1028) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1278), .ZN(n1131) );
NAND2_X1 U1021 ( .A1(n1280), .A2(n1164), .ZN(n1278) );
INV_X1 U1022 ( .A(G902), .ZN(n1164) );
INV_X1 U1023 ( .A(G237), .ZN(n1280) );
NAND2_X1 U1024 ( .A1(n1281), .A2(n1213), .ZN(n1279) );
XOR2_X1 U1025 ( .A(G902), .B(KEYINPUT23), .Z(n1213) );
XOR2_X1 U1026 ( .A(n1128), .B(n1282), .Z(n1281) );
XNOR2_X1 U1027 ( .A(G125), .B(n1283), .ZN(n1282) );
NOR2_X1 U1028 ( .A1(KEYINPUT28), .A2(n1284), .ZN(n1283) );
XOR2_X1 U1029 ( .A(KEYINPUT0), .B(n1127), .Z(n1284) );
XOR2_X1 U1030 ( .A(G146), .B(n1251), .Z(n1127) );
XNOR2_X1 U1031 ( .A(G128), .B(n1240), .ZN(n1251) );
INV_X1 U1032 ( .A(G143), .ZN(n1240) );
XOR2_X1 U1033 ( .A(n1072), .B(n1285), .Z(n1128) );
XOR2_X1 U1034 ( .A(n1286), .B(n1287), .Z(n1285) );
NAND2_X1 U1035 ( .A1(G224), .A2(n1017), .ZN(n1287) );
INV_X1 U1036 ( .A(G953), .ZN(n1017) );
NAND2_X1 U1037 ( .A1(KEYINPUT29), .A2(n1073), .ZN(n1286) );
XOR2_X1 U1038 ( .A(n1271), .B(n1288), .Z(n1073) );
XNOR2_X1 U1039 ( .A(n1289), .B(KEYINPUT27), .ZN(n1288) );
NAND2_X1 U1040 ( .A1(KEYINPUT5), .A2(n1272), .ZN(n1289) );
XNOR2_X1 U1041 ( .A(G101), .B(KEYINPUT44), .ZN(n1272) );
XNOR2_X1 U1042 ( .A(G104), .B(G107), .ZN(n1271) );
XOR2_X1 U1043 ( .A(n1290), .B(n1233), .Z(n1072) );
XOR2_X1 U1044 ( .A(G122), .B(G113), .Z(n1233) );
XNOR2_X1 U1045 ( .A(G110), .B(n1225), .ZN(n1290) );
XNOR2_X1 U1046 ( .A(n1193), .B(G119), .ZN(n1225) );
INV_X1 U1047 ( .A(G116), .ZN(n1193) );
XNOR2_X1 U1048 ( .A(G110), .B(KEYINPUT7), .ZN(n1197) );
endmodule


