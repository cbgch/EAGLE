//Key = 1010110110100011000101001011000011010101011001111111011001110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398;

XNOR2_X1 U768 ( .A(G107), .B(n1058), .ZN(G9) );
NOR2_X1 U769 ( .A1(n1059), .A2(n1060), .ZN(G75) );
NOR3_X1 U770 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NAND3_X1 U771 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1061) );
NAND4_X1 U772 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
NAND2_X1 U773 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U774 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U775 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND3_X1 U776 ( .A1(n1077), .A2(n1078), .A3(KEYINPUT2), .ZN(n1076) );
NAND2_X1 U777 ( .A1(n1079), .A2(n1080), .ZN(n1071) );
NAND3_X1 U778 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1080) );
OR2_X1 U779 ( .A1(n1084), .A2(KEYINPUT2), .ZN(n1083) );
NAND2_X1 U780 ( .A1(n1085), .A2(n1086), .ZN(n1081) );
XNOR2_X1 U781 ( .A(KEYINPUT32), .B(n1087), .ZN(n1086) );
NAND4_X1 U782 ( .A1(n1079), .A2(n1073), .A3(n1088), .A4(n1089), .ZN(n1064) );
NAND2_X1 U783 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U784 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
INV_X1 U785 ( .A(KEYINPUT39), .ZN(n1093) );
NAND4_X1 U786 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1067), .ZN(n1088) );
INV_X1 U787 ( .A(n1091), .ZN(n1067) );
NAND2_X1 U788 ( .A1(KEYINPUT39), .A2(n1092), .ZN(n1096) );
NAND2_X1 U789 ( .A1(n1069), .A2(n1097), .ZN(n1095) );
NAND2_X1 U790 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U791 ( .A1(n1100), .A2(n1068), .ZN(n1094) );
AND3_X1 U792 ( .A1(n1101), .A2(n1102), .A3(n1065), .ZN(n1059) );
NAND4_X1 U793 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1065) );
NOR4_X1 U794 ( .A1(n1107), .A2(n1108), .A3(n1109), .A4(n1110), .ZN(n1106) );
XOR2_X1 U795 ( .A(G478), .B(n1111), .Z(n1110) );
NOR2_X1 U796 ( .A1(KEYINPUT9), .A2(n1112), .ZN(n1111) );
NOR3_X1 U797 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1105) );
NOR2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1113) );
XNOR2_X1 U799 ( .A(KEYINPUT29), .B(n1118), .ZN(n1117) );
XNOR2_X1 U800 ( .A(G472), .B(KEYINPUT1), .ZN(n1116) );
NAND2_X1 U801 ( .A1(n1119), .A2(n1120), .ZN(n1104) );
XNOR2_X1 U802 ( .A(KEYINPUT14), .B(n1121), .ZN(n1103) );
XOR2_X1 U803 ( .A(n1122), .B(n1123), .Z(G72) );
XOR2_X1 U804 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND2_X1 U805 ( .A1(G953), .A2(n1126), .ZN(n1125) );
NAND2_X1 U806 ( .A1(G900), .A2(G227), .ZN(n1126) );
NAND2_X1 U807 ( .A1(n1127), .A2(n1128), .ZN(n1124) );
NAND2_X1 U808 ( .A1(G953), .A2(n1129), .ZN(n1128) );
XNOR2_X1 U809 ( .A(n1130), .B(n1131), .ZN(n1127) );
XNOR2_X1 U810 ( .A(n1132), .B(n1133), .ZN(n1131) );
NAND2_X1 U811 ( .A1(KEYINPUT0), .A2(n1134), .ZN(n1133) );
NAND3_X1 U812 ( .A1(n1135), .A2(n1136), .A3(KEYINPUT7), .ZN(n1132) );
NAND2_X1 U813 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U814 ( .A(KEYINPUT16), .B(n1139), .Z(n1137) );
NAND2_X1 U815 ( .A1(G137), .A2(n1140), .ZN(n1135) );
XNOR2_X1 U816 ( .A(n1139), .B(KEYINPUT30), .ZN(n1140) );
XOR2_X1 U817 ( .A(n1141), .B(n1142), .Z(n1139) );
XNOR2_X1 U818 ( .A(n1143), .B(G131), .ZN(n1142) );
NOR2_X1 U819 ( .A1(n1144), .A2(G953), .ZN(n1122) );
NAND4_X1 U820 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(G69) );
NAND3_X1 U821 ( .A1(KEYINPUT35), .A2(n1149), .A3(n1150), .ZN(n1148) );
NAND2_X1 U822 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
OR2_X1 U823 ( .A1(n1153), .A2(G224), .ZN(n1152) );
OR2_X1 U824 ( .A1(n1150), .A2(KEYINPUT35), .ZN(n1147) );
NAND3_X1 U825 ( .A1(G224), .A2(n1154), .A3(G898), .ZN(n1146) );
NAND2_X1 U826 ( .A1(KEYINPUT35), .A2(n1155), .ZN(n1154) );
OR2_X1 U827 ( .A1(n1150), .A2(n1153), .ZN(n1155) );
NAND2_X1 U828 ( .A1(n1156), .A2(n1153), .ZN(n1145) );
NAND2_X1 U829 ( .A1(n1157), .A2(KEYINPUT35), .ZN(n1156) );
XOR2_X1 U830 ( .A(n1150), .B(n1158), .Z(n1157) );
NOR2_X1 U831 ( .A1(n1159), .A2(KEYINPUT23), .ZN(n1158) );
NAND2_X1 U832 ( .A1(n1160), .A2(n1151), .ZN(n1150) );
INV_X1 U833 ( .A(n1161), .ZN(n1151) );
XNOR2_X1 U834 ( .A(n1162), .B(n1163), .ZN(n1160) );
XNOR2_X1 U835 ( .A(n1164), .B(KEYINPUT34), .ZN(n1163) );
NAND3_X1 U836 ( .A1(n1165), .A2(n1166), .A3(KEYINPUT46), .ZN(n1164) );
NAND2_X1 U837 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U838 ( .A(KEYINPUT59), .B(n1169), .Z(n1165) );
NOR2_X1 U839 ( .A1(n1167), .A2(n1168), .ZN(n1169) );
NOR2_X1 U840 ( .A1(n1170), .A2(n1171), .ZN(G66) );
NOR3_X1 U841 ( .A1(n1119), .A2(n1172), .A3(n1173), .ZN(n1171) );
NOR3_X1 U842 ( .A1(n1174), .A2(n1120), .A3(n1175), .ZN(n1173) );
NOR2_X1 U843 ( .A1(n1176), .A2(n1177), .ZN(n1172) );
NOR2_X1 U844 ( .A1(n1178), .A2(n1120), .ZN(n1176) );
NOR2_X1 U845 ( .A1(n1170), .A2(n1179), .ZN(G63) );
XOR2_X1 U846 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U847 ( .A(KEYINPUT13), .B(n1182), .Z(n1181) );
AND2_X1 U848 ( .A1(G478), .A2(n1183), .ZN(n1182) );
NOR2_X1 U849 ( .A1(n1170), .A2(n1184), .ZN(G60) );
XOR2_X1 U850 ( .A(n1185), .B(n1186), .Z(n1184) );
AND2_X1 U851 ( .A1(G475), .A2(n1183), .ZN(n1185) );
XNOR2_X1 U852 ( .A(G104), .B(n1187), .ZN(G6) );
NOR2_X1 U853 ( .A1(n1170), .A2(n1188), .ZN(G57) );
NOR2_X1 U854 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U855 ( .A(n1191), .B(KEYINPUT50), .Z(n1190) );
NAND2_X1 U856 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NOR2_X1 U857 ( .A1(n1192), .A2(n1193), .ZN(n1189) );
XNOR2_X1 U858 ( .A(n1194), .B(n1195), .ZN(n1193) );
XOR2_X1 U859 ( .A(KEYINPUT15), .B(G101), .Z(n1195) );
AND2_X1 U860 ( .A1(n1196), .A2(n1197), .ZN(n1192) );
NAND2_X1 U861 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U862 ( .A(KEYINPUT51), .B(n1200), .Z(n1199) );
XNOR2_X1 U863 ( .A(n1201), .B(n1202), .ZN(n1198) );
NAND2_X1 U864 ( .A1(n1200), .A2(n1203), .ZN(n1196) );
XNOR2_X1 U865 ( .A(n1204), .B(n1201), .ZN(n1203) );
AND2_X1 U866 ( .A1(n1183), .A2(G472), .ZN(n1200) );
NOR2_X1 U867 ( .A1(n1170), .A2(n1205), .ZN(G54) );
XOR2_X1 U868 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U869 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U870 ( .A(n1210), .B(n1211), .Z(n1209) );
XNOR2_X1 U871 ( .A(G110), .B(G140), .ZN(n1208) );
XNOR2_X1 U872 ( .A(n1212), .B(n1213), .ZN(n1206) );
XOR2_X1 U873 ( .A(n1214), .B(n1215), .Z(n1213) );
NOR2_X1 U874 ( .A1(n1141), .A2(KEYINPUT11), .ZN(n1215) );
INV_X1 U875 ( .A(n1216), .ZN(n1141) );
AND2_X1 U876 ( .A1(G469), .A2(n1183), .ZN(n1214) );
NOR2_X1 U877 ( .A1(n1170), .A2(n1217), .ZN(G51) );
XOR2_X1 U878 ( .A(n1218), .B(n1219), .Z(n1217) );
NOR2_X1 U879 ( .A1(n1220), .A2(n1175), .ZN(n1219) );
INV_X1 U880 ( .A(n1183), .ZN(n1175) );
NOR2_X1 U881 ( .A1(n1221), .A2(n1178), .ZN(n1183) );
INV_X1 U882 ( .A(n1062), .ZN(n1178) );
NAND2_X1 U883 ( .A1(n1159), .A2(n1144), .ZN(n1062) );
AND2_X1 U884 ( .A1(n1222), .A2(n1223), .ZN(n1144) );
NOR4_X1 U885 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1223) );
NOR4_X1 U886 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1222) );
NOR2_X1 U887 ( .A1(n1109), .A2(n1232), .ZN(n1231) );
INV_X1 U888 ( .A(n1233), .ZN(n1230) );
AND4_X1 U889 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1159) );
AND4_X1 U890 ( .A1(n1238), .A2(n1239), .A3(n1058), .A4(n1240), .ZN(n1237) );
NAND3_X1 U891 ( .A1(n1241), .A2(n1242), .A3(n1069), .ZN(n1058) );
OR3_X1 U892 ( .A1(n1243), .A2(n1099), .A3(n1244), .ZN(n1239) );
INV_X1 U893 ( .A(n1242), .ZN(n1099) );
XOR2_X1 U894 ( .A(KEYINPUT24), .B(n1100), .Z(n1243) );
NOR3_X1 U895 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1236) );
NOR2_X1 U896 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
INV_X1 U897 ( .A(KEYINPUT57), .ZN(n1248) );
NOR2_X1 U898 ( .A1(KEYINPUT57), .A2(n1250), .ZN(n1246) );
NAND4_X1 U899 ( .A1(n1092), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1250) );
INV_X1 U900 ( .A(n1187), .ZN(n1245) );
NAND3_X1 U901 ( .A1(n1069), .A2(n1241), .A3(n1254), .ZN(n1187) );
NAND2_X1 U902 ( .A1(n1255), .A2(KEYINPUT53), .ZN(n1218) );
XNOR2_X1 U903 ( .A(n1256), .B(n1257), .ZN(n1255) );
XOR2_X1 U904 ( .A(n1258), .B(n1259), .Z(n1256) );
AND2_X1 U905 ( .A1(n1260), .A2(n1102), .ZN(n1170) );
INV_X1 U906 ( .A(G952), .ZN(n1102) );
XNOR2_X1 U907 ( .A(G953), .B(KEYINPUT8), .ZN(n1260) );
XNOR2_X1 U908 ( .A(G146), .B(n1261), .ZN(G48) );
NAND2_X1 U909 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NAND2_X1 U910 ( .A1(KEYINPUT55), .A2(n1228), .ZN(n1263) );
OR2_X1 U911 ( .A1(KEYINPUT60), .A2(n1228), .ZN(n1262) );
AND3_X1 U912 ( .A1(n1264), .A2(n1254), .A3(n1265), .ZN(n1228) );
XNOR2_X1 U913 ( .A(G143), .B(n1233), .ZN(G45) );
NAND3_X1 U914 ( .A1(n1266), .A2(n1100), .A3(n1267), .ZN(n1233) );
NOR3_X1 U915 ( .A1(n1075), .A2(n1268), .A3(n1269), .ZN(n1267) );
XOR2_X1 U916 ( .A(n1270), .B(n1271), .Z(G42) );
NOR2_X1 U917 ( .A1(n1232), .A2(n1272), .ZN(n1271) );
XNOR2_X1 U918 ( .A(KEYINPUT45), .B(n1109), .ZN(n1272) );
NAND4_X1 U919 ( .A1(n1266), .A2(n1254), .A3(n1273), .A4(n1274), .ZN(n1232) );
XNOR2_X1 U920 ( .A(G140), .B(KEYINPUT41), .ZN(n1270) );
XNOR2_X1 U921 ( .A(n1138), .B(n1227), .ZN(G39) );
AND3_X1 U922 ( .A1(n1068), .A2(n1079), .A3(n1265), .ZN(n1227) );
XNOR2_X1 U923 ( .A(n1143), .B(n1229), .ZN(G36) );
NOR3_X1 U924 ( .A1(n1275), .A2(n1109), .A3(n1276), .ZN(n1229) );
XOR2_X1 U925 ( .A(G131), .B(n1226), .Z(G33) );
AND4_X1 U926 ( .A1(n1266), .A2(n1254), .A3(n1100), .A4(n1079), .ZN(n1226) );
INV_X1 U927 ( .A(n1109), .ZN(n1079) );
NAND2_X1 U928 ( .A1(n1077), .A2(n1277), .ZN(n1109) );
INV_X1 U929 ( .A(n1275), .ZN(n1266) );
XNOR2_X1 U930 ( .A(n1278), .B(n1225), .ZN(G30) );
AND3_X1 U931 ( .A1(n1264), .A2(n1242), .A3(n1265), .ZN(n1225) );
NOR3_X1 U932 ( .A1(n1279), .A2(n1273), .A3(n1275), .ZN(n1265) );
NAND2_X1 U933 ( .A1(n1251), .A2(n1280), .ZN(n1275) );
INV_X1 U934 ( .A(n1075), .ZN(n1264) );
XNOR2_X1 U935 ( .A(G101), .B(n1234), .ZN(G3) );
NAND3_X1 U936 ( .A1(n1068), .A2(n1241), .A3(n1100), .ZN(n1234) );
XOR2_X1 U937 ( .A(G125), .B(n1224), .Z(G27) );
AND4_X1 U938 ( .A1(n1280), .A2(n1274), .A3(n1073), .A4(n1281), .ZN(n1224) );
NOR3_X1 U939 ( .A1(n1098), .A2(n1282), .A3(n1075), .ZN(n1281) );
INV_X1 U940 ( .A(n1254), .ZN(n1098) );
NAND2_X1 U941 ( .A1(n1091), .A2(n1283), .ZN(n1280) );
NAND4_X1 U942 ( .A1(n1284), .A2(G902), .A3(G953), .A4(n1129), .ZN(n1283) );
INV_X1 U943 ( .A(G900), .ZN(n1129) );
XOR2_X1 U944 ( .A(n1285), .B(KEYINPUT18), .Z(n1284) );
XNOR2_X1 U945 ( .A(G122), .B(n1235), .ZN(G24) );
NAND4_X1 U946 ( .A1(n1286), .A2(n1069), .A3(n1287), .A4(n1107), .ZN(n1235) );
NOR2_X1 U947 ( .A1(n1282), .A2(n1274), .ZN(n1069) );
XNOR2_X1 U948 ( .A(G119), .B(n1238), .ZN(G21) );
NAND4_X1 U949 ( .A1(n1068), .A2(n1286), .A3(n1274), .A4(n1282), .ZN(n1238) );
INV_X1 U950 ( .A(n1273), .ZN(n1282) );
XOR2_X1 U951 ( .A(G116), .B(n1288), .Z(G18) );
NOR2_X1 U952 ( .A1(n1244), .A2(n1276), .ZN(n1288) );
NAND2_X1 U953 ( .A1(n1100), .A2(n1242), .ZN(n1276) );
NOR2_X1 U954 ( .A1(n1107), .A2(n1269), .ZN(n1242) );
INV_X1 U955 ( .A(n1287), .ZN(n1269) );
INV_X1 U956 ( .A(n1286), .ZN(n1244) );
NOR3_X1 U957 ( .A1(n1084), .A2(n1289), .A3(n1075), .ZN(n1286) );
XNOR2_X1 U958 ( .A(n1253), .B(KEYINPUT4), .ZN(n1075) );
XNOR2_X1 U959 ( .A(G113), .B(n1240), .ZN(G15) );
NAND3_X1 U960 ( .A1(n1254), .A2(n1100), .A3(n1290), .ZN(n1240) );
NOR3_X1 U961 ( .A1(n1253), .A2(n1289), .A3(n1084), .ZN(n1290) );
INV_X1 U962 ( .A(n1073), .ZN(n1084) );
NAND2_X1 U963 ( .A1(n1291), .A2(n1292), .ZN(n1073) );
OR2_X1 U964 ( .A1(n1082), .A2(KEYINPUT32), .ZN(n1292) );
NAND3_X1 U965 ( .A1(n1087), .A2(n1121), .A3(KEYINPUT32), .ZN(n1291) );
AND2_X1 U966 ( .A1(n1293), .A2(n1279), .ZN(n1100) );
XNOR2_X1 U967 ( .A(n1273), .B(KEYINPUT36), .ZN(n1293) );
NOR2_X1 U968 ( .A1(n1287), .A2(n1268), .ZN(n1254) );
INV_X1 U969 ( .A(n1107), .ZN(n1268) );
XNOR2_X1 U970 ( .A(n1249), .B(n1294), .ZN(G12) );
NOR2_X1 U971 ( .A1(KEYINPUT20), .A2(n1295), .ZN(n1294) );
NAND2_X1 U972 ( .A1(n1092), .A2(n1241), .ZN(n1249) );
NOR3_X1 U973 ( .A1(n1253), .A2(n1289), .A3(n1082), .ZN(n1241) );
INV_X1 U974 ( .A(n1251), .ZN(n1082) );
NOR2_X1 U975 ( .A1(n1087), .A2(n1085), .ZN(n1251) );
INV_X1 U976 ( .A(n1121), .ZN(n1085) );
NAND2_X1 U977 ( .A1(G221), .A2(n1296), .ZN(n1121) );
INV_X1 U978 ( .A(n1108), .ZN(n1087) );
XNOR2_X1 U979 ( .A(n1297), .B(G469), .ZN(n1108) );
NAND3_X1 U980 ( .A1(n1298), .A2(n1299), .A3(n1221), .ZN(n1297) );
OR3_X1 U981 ( .A1(n1300), .A2(n1301), .A3(KEYINPUT27), .ZN(n1299) );
NAND2_X1 U982 ( .A1(n1302), .A2(KEYINPUT27), .ZN(n1298) );
XOR2_X1 U983 ( .A(n1301), .B(n1300), .Z(n1302) );
XOR2_X1 U984 ( .A(n1303), .B(n1304), .Z(n1300) );
INV_X1 U985 ( .A(n1212), .ZN(n1304) );
XNOR2_X1 U986 ( .A(KEYINPUT28), .B(n1305), .ZN(n1303) );
NOR2_X1 U987 ( .A1(KEYINPUT17), .A2(n1306), .ZN(n1305) );
XNOR2_X1 U988 ( .A(n1210), .B(n1216), .ZN(n1306) );
NAND3_X1 U989 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1216) );
NAND3_X1 U990 ( .A1(G143), .A2(n1310), .A3(G128), .ZN(n1309) );
NAND2_X1 U991 ( .A1(n1311), .A2(n1312), .ZN(n1308) );
INV_X1 U992 ( .A(KEYINPUT38), .ZN(n1312) );
NAND2_X1 U993 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
NAND3_X1 U994 ( .A1(n1278), .A2(n1315), .A3(n1310), .ZN(n1314) );
NAND2_X1 U995 ( .A1(n1316), .A2(G146), .ZN(n1313) );
NAND2_X1 U996 ( .A1(n1317), .A2(KEYINPUT38), .ZN(n1307) );
XNOR2_X1 U997 ( .A(n1278), .B(n1318), .ZN(n1317) );
NOR2_X1 U998 ( .A1(G143), .A2(n1310), .ZN(n1318) );
NAND4_X1 U999 ( .A1(n1319), .A2(n1320), .A3(n1321), .A4(n1322), .ZN(n1210) );
NAND2_X1 U1000 ( .A1(KEYINPUT12), .A2(n1323), .ZN(n1322) );
NAND2_X1 U1001 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
NAND2_X1 U1002 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
OR3_X1 U1003 ( .A1(n1326), .A2(n1328), .A3(KEYINPUT12), .ZN(n1321) );
NAND3_X1 U1004 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1320) );
INV_X1 U1005 ( .A(KEYINPUT62), .ZN(n1330) );
XOR2_X1 U1006 ( .A(KEYINPUT12), .B(n1326), .Z(n1329) );
NOR2_X1 U1007 ( .A1(n1327), .A2(G101), .ZN(n1328) );
INV_X1 U1008 ( .A(KEYINPUT37), .ZN(n1327) );
NAND2_X1 U1009 ( .A1(KEYINPUT62), .A2(G101), .ZN(n1319) );
XNOR2_X1 U1010 ( .A(n1331), .B(n1211), .ZN(n1301) );
AND2_X1 U1011 ( .A1(G227), .A2(n1153), .ZN(n1211) );
NAND2_X1 U1012 ( .A1(n1332), .A2(KEYINPUT54), .ZN(n1331) );
XNOR2_X1 U1013 ( .A(G140), .B(n1333), .ZN(n1332) );
NOR2_X1 U1014 ( .A1(G110), .A2(KEYINPUT52), .ZN(n1333) );
INV_X1 U1015 ( .A(n1252), .ZN(n1289) );
NAND2_X1 U1016 ( .A1(n1091), .A2(n1334), .ZN(n1252) );
NAND3_X1 U1017 ( .A1(n1161), .A2(n1285), .A3(G902), .ZN(n1334) );
NOR2_X1 U1018 ( .A1(n1153), .A2(G898), .ZN(n1161) );
NAND3_X1 U1019 ( .A1(n1101), .A2(n1285), .A3(G952), .ZN(n1091) );
NAND2_X1 U1020 ( .A1(G237), .A2(G234), .ZN(n1285) );
INV_X1 U1021 ( .A(n1063), .ZN(n1101) );
XOR2_X1 U1022 ( .A(G953), .B(KEYINPUT31), .Z(n1063) );
OR2_X1 U1023 ( .A1(n1077), .A2(n1078), .ZN(n1253) );
INV_X1 U1024 ( .A(n1277), .ZN(n1078) );
NAND2_X1 U1025 ( .A1(G214), .A2(n1335), .ZN(n1277) );
XNOR2_X1 U1026 ( .A(n1336), .B(n1220), .ZN(n1077) );
NAND2_X1 U1027 ( .A1(G210), .A2(n1335), .ZN(n1220) );
NAND2_X1 U1028 ( .A1(n1337), .A2(n1221), .ZN(n1335) );
NAND2_X1 U1029 ( .A1(n1338), .A2(n1221), .ZN(n1336) );
XOR2_X1 U1030 ( .A(n1258), .B(n1339), .Z(n1338) );
NOR2_X1 U1031 ( .A1(KEYINPUT25), .A2(n1340), .ZN(n1339) );
XOR2_X1 U1032 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1033 ( .A(KEYINPUT19), .B(n1259), .Z(n1342) );
AND2_X1 U1034 ( .A1(n1343), .A2(n1153), .ZN(n1259) );
XNOR2_X1 U1035 ( .A(G224), .B(KEYINPUT26), .ZN(n1343) );
NAND2_X1 U1036 ( .A1(KEYINPUT10), .A2(n1257), .ZN(n1341) );
XNOR2_X1 U1037 ( .A(n1344), .B(n1130), .ZN(n1257) );
XOR2_X1 U1038 ( .A(n1345), .B(n1162), .Z(n1258) );
XOR2_X1 U1039 ( .A(G110), .B(G122), .Z(n1162) );
XNOR2_X1 U1040 ( .A(n1167), .B(n1168), .ZN(n1345) );
XNOR2_X1 U1041 ( .A(n1202), .B(KEYINPUT63), .ZN(n1168) );
AND2_X1 U1042 ( .A1(n1346), .A2(n1324), .ZN(n1167) );
NAND2_X1 U1043 ( .A1(G101), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1044 ( .A(KEYINPUT47), .B(n1347), .Z(n1346) );
NOR2_X1 U1045 ( .A1(G101), .A2(n1326), .ZN(n1347) );
XNOR2_X1 U1046 ( .A(G104), .B(n1348), .ZN(n1326) );
AND3_X1 U1047 ( .A1(n1273), .A2(n1274), .A3(n1068), .ZN(n1092) );
NOR2_X1 U1048 ( .A1(n1287), .A2(n1107), .ZN(n1068) );
XNOR2_X1 U1049 ( .A(n1349), .B(G475), .ZN(n1107) );
OR2_X1 U1050 ( .A1(n1186), .A2(G902), .ZN(n1349) );
XNOR2_X1 U1051 ( .A(n1350), .B(n1351), .ZN(n1186) );
XOR2_X1 U1052 ( .A(n1352), .B(n1353), .Z(n1351) );
XNOR2_X1 U1053 ( .A(n1354), .B(n1355), .ZN(n1353) );
NOR2_X1 U1054 ( .A1(KEYINPUT22), .A2(n1356), .ZN(n1355) );
XOR2_X1 U1055 ( .A(n1357), .B(n1358), .Z(n1356) );
XNOR2_X1 U1056 ( .A(n1315), .B(G131), .ZN(n1358) );
INV_X1 U1057 ( .A(G143), .ZN(n1315) );
NAND3_X1 U1058 ( .A1(n1337), .A2(n1153), .A3(G214), .ZN(n1357) );
INV_X1 U1059 ( .A(G104), .ZN(n1354) );
XNOR2_X1 U1060 ( .A(G113), .B(n1359), .ZN(n1350) );
XNOR2_X1 U1061 ( .A(n1310), .B(G122), .ZN(n1359) );
INV_X1 U1062 ( .A(G146), .ZN(n1310) );
XNOR2_X1 U1063 ( .A(n1112), .B(G478), .ZN(n1287) );
OR2_X1 U1064 ( .A1(n1180), .A2(G902), .ZN(n1112) );
XNOR2_X1 U1065 ( .A(n1360), .B(n1361), .ZN(n1180) );
XOR2_X1 U1066 ( .A(n1362), .B(n1363), .Z(n1361) );
XOR2_X1 U1067 ( .A(G122), .B(G116), .Z(n1363) );
XNOR2_X1 U1068 ( .A(KEYINPUT21), .B(n1143), .ZN(n1362) );
XOR2_X1 U1069 ( .A(n1364), .B(n1316), .Z(n1360) );
XNOR2_X1 U1070 ( .A(n1365), .B(n1348), .ZN(n1364) );
INV_X1 U1071 ( .A(G107), .ZN(n1348) );
NAND2_X1 U1072 ( .A1(G217), .A2(n1366), .ZN(n1365) );
INV_X1 U1073 ( .A(n1279), .ZN(n1274) );
NOR2_X1 U1074 ( .A1(n1367), .A2(n1115), .ZN(n1279) );
NOR2_X1 U1075 ( .A1(n1120), .A2(n1119), .ZN(n1115) );
AND2_X1 U1076 ( .A1(n1368), .A2(n1120), .ZN(n1367) );
NAND2_X1 U1077 ( .A1(G217), .A2(n1296), .ZN(n1120) );
NAND2_X1 U1078 ( .A1(G234), .A2(n1221), .ZN(n1296) );
XOR2_X1 U1079 ( .A(KEYINPUT56), .B(n1119), .Z(n1368) );
NOR2_X1 U1080 ( .A1(n1177), .A2(G902), .ZN(n1119) );
INV_X1 U1081 ( .A(n1174), .ZN(n1177) );
XNOR2_X1 U1082 ( .A(n1369), .B(n1370), .ZN(n1174) );
XOR2_X1 U1083 ( .A(n1371), .B(n1372), .Z(n1370) );
XNOR2_X1 U1084 ( .A(n1373), .B(n1295), .ZN(n1372) );
INV_X1 U1085 ( .A(G110), .ZN(n1295) );
NAND2_X1 U1086 ( .A1(KEYINPUT58), .A2(n1374), .ZN(n1373) );
XOR2_X1 U1087 ( .A(n1375), .B(n1352), .Z(n1374) );
XNOR2_X1 U1088 ( .A(n1134), .B(n1130), .ZN(n1352) );
XOR2_X1 U1089 ( .A(G125), .B(KEYINPUT48), .Z(n1130) );
INV_X1 U1090 ( .A(G140), .ZN(n1134) );
NOR2_X1 U1091 ( .A1(G146), .A2(KEYINPUT6), .ZN(n1375) );
NAND2_X1 U1092 ( .A1(G221), .A2(n1366), .ZN(n1371) );
AND2_X1 U1093 ( .A1(G234), .A2(n1153), .ZN(n1366) );
XNOR2_X1 U1094 ( .A(G119), .B(n1376), .ZN(n1369) );
XNOR2_X1 U1095 ( .A(n1138), .B(G128), .ZN(n1376) );
INV_X1 U1096 ( .A(G137), .ZN(n1138) );
NOR2_X1 U1097 ( .A1(n1377), .A2(n1114), .ZN(n1273) );
NOR2_X1 U1098 ( .A1(n1118), .A2(G472), .ZN(n1114) );
AND2_X1 U1099 ( .A1(n1378), .A2(n1118), .ZN(n1377) );
NAND2_X1 U1100 ( .A1(n1221), .A2(n1379), .ZN(n1118) );
NAND2_X1 U1101 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
NAND2_X1 U1102 ( .A1(n1382), .A2(n1383), .ZN(n1381) );
XOR2_X1 U1103 ( .A(n1384), .B(n1201), .Z(n1383) );
XOR2_X1 U1104 ( .A(n1194), .B(n1385), .Z(n1382) );
XOR2_X1 U1105 ( .A(n1386), .B(KEYINPUT3), .Z(n1380) );
NAND2_X1 U1106 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
XNOR2_X1 U1107 ( .A(n1194), .B(n1385), .ZN(n1388) );
NOR2_X1 U1108 ( .A1(n1389), .A2(G101), .ZN(n1385) );
INV_X1 U1109 ( .A(KEYINPUT5), .ZN(n1389) );
NAND3_X1 U1110 ( .A1(n1337), .A2(n1153), .A3(G210), .ZN(n1194) );
INV_X1 U1111 ( .A(G953), .ZN(n1153) );
INV_X1 U1112 ( .A(G237), .ZN(n1337) );
XNOR2_X1 U1113 ( .A(n1201), .B(n1384), .ZN(n1387) );
NAND2_X1 U1114 ( .A1(KEYINPUT33), .A2(n1202), .ZN(n1384) );
INV_X1 U1115 ( .A(n1204), .ZN(n1202) );
XOR2_X1 U1116 ( .A(G113), .B(n1390), .Z(n1204) );
XOR2_X1 U1117 ( .A(G119), .B(G116), .Z(n1390) );
XNOR2_X1 U1118 ( .A(n1212), .B(n1344), .ZN(n1201) );
XOR2_X1 U1119 ( .A(G146), .B(n1316), .Z(n1344) );
XNOR2_X1 U1120 ( .A(n1278), .B(G143), .ZN(n1316) );
INV_X1 U1121 ( .A(G128), .ZN(n1278) );
XNOR2_X1 U1122 ( .A(n1391), .B(KEYINPUT42), .ZN(n1212) );
NAND3_X1 U1123 ( .A1(n1392), .A2(n1393), .A3(n1394), .ZN(n1391) );
NAND2_X1 U1124 ( .A1(G131), .A2(n1395), .ZN(n1394) );
OR3_X1 U1125 ( .A1(n1395), .A2(G131), .A3(KEYINPUT43), .ZN(n1393) );
OR2_X1 U1126 ( .A1(KEYINPUT40), .A2(n1396), .ZN(n1395) );
NAND2_X1 U1127 ( .A1(KEYINPUT43), .A2(n1396), .ZN(n1392) );
XOR2_X1 U1128 ( .A(n1397), .B(n1398), .Z(n1396) );
NOR2_X1 U1129 ( .A1(KEYINPUT61), .A2(n1143), .ZN(n1398) );
INV_X1 U1130 ( .A(G134), .ZN(n1143) );
XNOR2_X1 U1131 ( .A(G137), .B(KEYINPUT44), .ZN(n1397) );
INV_X1 U1132 ( .A(G902), .ZN(n1221) );
XNOR2_X1 U1133 ( .A(G472), .B(KEYINPUT49), .ZN(n1378) );
endmodule


