//Key = 1001000111010011111100101110110011000110110111010100110011110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340;

XNOR2_X1 U723 ( .A(G107), .B(n1008), .ZN(G9) );
NOR2_X1 U724 ( .A1(n1009), .A2(n1010), .ZN(G75) );
NOR4_X1 U725 ( .A1(n1011), .A2(n1012), .A3(G953), .A4(n1013), .ZN(n1010) );
NOR2_X1 U726 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR2_X1 U727 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR3_X1 U728 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1017) );
NOR3_X1 U729 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1019) );
NOR2_X1 U730 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NOR2_X1 U731 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U732 ( .A1(KEYINPUT6), .A2(n1028), .ZN(n1026) );
NOR3_X1 U733 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1022) );
XOR2_X1 U734 ( .A(KEYINPUT29), .B(n1032), .Z(n1029) );
NOR2_X1 U735 ( .A1(n1033), .A2(n1034), .ZN(n1021) );
NOR3_X1 U736 ( .A1(n1034), .A2(n1035), .A3(n1025), .ZN(n1016) );
INV_X1 U737 ( .A(n1036), .ZN(n1025) );
NOR2_X1 U738 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U739 ( .A1(n1039), .A2(n1020), .ZN(n1038) );
NOR2_X1 U740 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U741 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U742 ( .A1(n1044), .A2(n1018), .ZN(n1037) );
NOR2_X1 U743 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U744 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND3_X1 U745 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1011) );
NAND2_X1 U746 ( .A1(KEYINPUT6), .A2(n1052), .ZN(n1050) );
NAND4_X1 U747 ( .A1(n1036), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1052) );
NOR2_X1 U748 ( .A1(n1015), .A2(n1020), .ZN(n1054) );
NOR3_X1 U749 ( .A1(n1013), .A2(G953), .A3(G952), .ZN(n1009) );
AND3_X1 U750 ( .A1(n1056), .A2(n1053), .A3(n1057), .ZN(n1013) );
NOR3_X1 U751 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
INV_X1 U752 ( .A(n1030), .ZN(n1059) );
NOR2_X1 U753 ( .A1(G469), .A2(n1061), .ZN(n1058) );
XOR2_X1 U754 ( .A(n1062), .B(KEYINPUT37), .Z(n1056) );
NAND4_X1 U755 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1062) );
XOR2_X1 U756 ( .A(n1067), .B(n1068), .Z(n1063) );
NAND2_X1 U757 ( .A1(KEYINPUT43), .A2(G478), .ZN(n1067) );
XOR2_X1 U758 ( .A(n1069), .B(n1070), .Z(G72) );
NOR2_X1 U759 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
AND2_X1 U760 ( .A1(G227), .A2(G900), .ZN(n1071) );
NOR2_X1 U761 ( .A1(KEYINPUT46), .A2(n1073), .ZN(n1069) );
XOR2_X1 U762 ( .A(n1074), .B(n1075), .Z(n1073) );
NOR2_X1 U763 ( .A1(n1051), .A2(G953), .ZN(n1075) );
NAND2_X1 U764 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NAND2_X1 U765 ( .A1(G953), .A2(n1078), .ZN(n1077) );
XOR2_X1 U766 ( .A(n1079), .B(n1080), .Z(n1076) );
XOR2_X1 U767 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND2_X1 U768 ( .A1(n1083), .A2(KEYINPUT58), .ZN(n1081) );
XOR2_X1 U769 ( .A(n1084), .B(n1085), .Z(n1083) );
NOR2_X1 U770 ( .A1(KEYINPUT21), .A2(n1086), .ZN(n1085) );
NAND2_X1 U771 ( .A1(n1087), .A2(n1088), .ZN(G69) );
NAND3_X1 U772 ( .A1(G953), .A2(n1089), .A3(n1090), .ZN(n1088) );
XOR2_X1 U773 ( .A(KEYINPUT3), .B(n1091), .Z(n1087) );
NOR2_X1 U774 ( .A1(n1092), .A2(n1090), .ZN(n1091) );
AND2_X1 U775 ( .A1(n1093), .A2(n1094), .ZN(n1090) );
NAND2_X1 U776 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U777 ( .A1(n1097), .A2(n1072), .ZN(n1096) );
INV_X1 U778 ( .A(n1098), .ZN(n1095) );
NAND2_X1 U779 ( .A1(n1099), .A2(n1098), .ZN(n1093) );
NAND3_X1 U780 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1098) );
XOR2_X1 U781 ( .A(n1103), .B(KEYINPUT4), .Z(n1102) );
NAND2_X1 U782 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
OR2_X1 U783 ( .A1(n1104), .A2(n1105), .ZN(n1101) );
XNOR2_X1 U784 ( .A(n1106), .B(n1107), .ZN(n1104) );
XNOR2_X1 U785 ( .A(G101), .B(KEYINPUT20), .ZN(n1106) );
NAND2_X1 U786 ( .A1(G953), .A2(n1108), .ZN(n1100) );
XOR2_X1 U787 ( .A(KEYINPUT54), .B(n1109), .Z(n1099) );
NOR2_X1 U788 ( .A1(n1049), .A2(G953), .ZN(n1109) );
AND2_X1 U789 ( .A1(n1089), .A2(G953), .ZN(n1092) );
NAND2_X1 U790 ( .A1(G898), .A2(G224), .ZN(n1089) );
NOR2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(G66) );
XOR2_X1 U792 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND2_X1 U793 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U794 ( .A1(n1116), .A2(KEYINPUT44), .ZN(n1112) );
XOR2_X1 U795 ( .A(n1117), .B(KEYINPUT59), .Z(n1116) );
NOR2_X1 U796 ( .A1(n1110), .A2(n1118), .ZN(G63) );
XOR2_X1 U797 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U798 ( .A(KEYINPUT27), .B(n1121), .Z(n1120) );
NOR2_X1 U799 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U800 ( .A1(n1110), .A2(n1124), .ZN(G60) );
XNOR2_X1 U801 ( .A(n1125), .B(n1126), .ZN(n1124) );
NOR2_X1 U802 ( .A1(n1127), .A2(n1123), .ZN(n1125) );
XOR2_X1 U803 ( .A(n1128), .B(n1129), .Z(G6) );
NOR2_X1 U804 ( .A1(n1110), .A2(n1130), .ZN(G57) );
XOR2_X1 U805 ( .A(n1131), .B(n1132), .Z(n1130) );
AND2_X1 U806 ( .A1(G472), .A2(n1114), .ZN(n1132) );
NOR4_X1 U807 ( .A1(n1133), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(G54) );
AND2_X1 U808 ( .A1(KEYINPUT11), .A2(n1110), .ZN(n1136) );
NOR3_X1 U809 ( .A1(KEYINPUT11), .A2(G953), .A3(G952), .ZN(n1135) );
NOR3_X1 U810 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1134) );
NOR2_X1 U811 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U812 ( .A(KEYINPUT55), .B(n1142), .Z(n1141) );
INV_X1 U813 ( .A(n1143), .ZN(n1137) );
NOR2_X1 U814 ( .A1(n1144), .A2(n1143), .ZN(n1133) );
XOR2_X1 U815 ( .A(n1145), .B(n1146), .Z(n1143) );
NOR3_X1 U816 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1146) );
AND2_X1 U817 ( .A1(n1150), .A2(KEYINPUT31), .ZN(n1149) );
NOR2_X1 U818 ( .A1(KEYINPUT31), .A2(n1151), .ZN(n1148) );
INV_X1 U819 ( .A(n1152), .ZN(n1151) );
NOR2_X1 U820 ( .A1(n1153), .A2(n1154), .ZN(n1144) );
NOR2_X1 U821 ( .A1(KEYINPUT55), .A2(n1155), .ZN(n1154) );
INV_X1 U822 ( .A(n1138), .ZN(n1155) );
NOR2_X1 U823 ( .A1(n1156), .A2(n1157), .ZN(n1138) );
NOR2_X1 U824 ( .A1(n1142), .A2(n1158), .ZN(n1153) );
NOR2_X1 U825 ( .A1(KEYINPUT55), .A2(n1157), .ZN(n1158) );
INV_X1 U826 ( .A(n1140), .ZN(n1157) );
XNOR2_X1 U827 ( .A(n1159), .B(n1160), .ZN(n1140) );
XOR2_X1 U828 ( .A(KEYINPUT47), .B(KEYINPUT38), .Z(n1160) );
INV_X1 U829 ( .A(n1156), .ZN(n1142) );
NAND3_X1 U830 ( .A1(n1161), .A2(n1162), .A3(G469), .ZN(n1156) );
NAND2_X1 U831 ( .A1(KEYINPUT0), .A2(n1123), .ZN(n1162) );
NAND2_X1 U832 ( .A1(n1163), .A2(n1164), .ZN(n1161) );
INV_X1 U833 ( .A(KEYINPUT0), .ZN(n1164) );
NAND2_X1 U834 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
NOR2_X1 U835 ( .A1(n1110), .A2(n1167), .ZN(G51) );
XOR2_X1 U836 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U837 ( .A1(n1170), .A2(n1123), .ZN(n1168) );
INV_X1 U838 ( .A(n1114), .ZN(n1123) );
NOR2_X1 U839 ( .A1(n1165), .A2(n1171), .ZN(n1114) );
INV_X1 U840 ( .A(n1166), .ZN(n1171) );
NAND2_X1 U841 ( .A1(n1051), .A2(n1172), .ZN(n1166) );
XOR2_X1 U842 ( .A(KEYINPUT34), .B(n1049), .Z(n1172) );
INV_X1 U843 ( .A(n1097), .ZN(n1049) );
NAND2_X1 U844 ( .A1(n1173), .A2(n1174), .ZN(n1097) );
AND4_X1 U845 ( .A1(n1008), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1174) );
NAND3_X1 U846 ( .A1(n1064), .A2(n1178), .A3(n1055), .ZN(n1008) );
AND4_X1 U847 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1129), .ZN(n1173) );
NAND3_X1 U848 ( .A1(n1064), .A2(n1178), .A3(n1027), .ZN(n1129) );
AND2_X1 U849 ( .A1(n1182), .A2(n1183), .ZN(n1051) );
NOR4_X1 U850 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1183) );
INV_X1 U851 ( .A(n1188), .ZN(n1185) );
AND4_X1 U852 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1182) );
NAND3_X1 U853 ( .A1(n1046), .A2(n1027), .A3(n1193), .ZN(n1192) );
XOR2_X1 U854 ( .A(n1194), .B(KEYINPUT63), .Z(n1165) );
NOR2_X1 U855 ( .A1(n1072), .A2(G952), .ZN(n1110) );
XOR2_X1 U856 ( .A(n1195), .B(n1191), .Z(G48) );
NAND4_X1 U857 ( .A1(n1048), .A2(n1027), .A3(n1196), .A4(n1197), .ZN(n1191) );
XNOR2_X1 U858 ( .A(G143), .B(n1190), .ZN(G45) );
NAND4_X1 U859 ( .A1(n1197), .A2(n1041), .A3(n1046), .A4(n1198), .ZN(n1190) );
AND3_X1 U860 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1198) );
XNOR2_X1 U861 ( .A(G140), .B(n1189), .ZN(G42) );
NAND4_X1 U862 ( .A1(n1193), .A2(n1027), .A3(n1202), .A4(n1203), .ZN(n1189) );
XOR2_X1 U863 ( .A(n1204), .B(n1187), .Z(G39) );
AND3_X1 U864 ( .A1(n1048), .A2(n1193), .A3(n1205), .ZN(n1187) );
INV_X1 U865 ( .A(n1206), .ZN(n1193) );
XOR2_X1 U866 ( .A(n1207), .B(KEYINPUT7), .Z(n1204) );
XOR2_X1 U867 ( .A(G134), .B(n1186), .Z(G36) );
NOR3_X1 U868 ( .A1(n1206), .A2(n1028), .A3(n1208), .ZN(n1186) );
INV_X1 U869 ( .A(n1055), .ZN(n1028) );
NAND3_X1 U870 ( .A1(n1197), .A2(n1201), .A3(n1053), .ZN(n1206) );
XOR2_X1 U871 ( .A(n1084), .B(n1209), .Z(G33) );
NAND4_X1 U872 ( .A1(n1053), .A2(n1197), .A3(n1027), .A4(n1210), .ZN(n1209) );
NOR2_X1 U873 ( .A1(n1208), .A2(n1211), .ZN(n1210) );
XNOR2_X1 U874 ( .A(KEYINPUT30), .B(n1201), .ZN(n1211) );
INV_X1 U875 ( .A(n1033), .ZN(n1197) );
INV_X1 U876 ( .A(n1018), .ZN(n1053) );
NAND2_X1 U877 ( .A1(n1212), .A2(n1043), .ZN(n1018) );
XOR2_X1 U878 ( .A(n1213), .B(n1188), .Z(G30) );
NAND4_X1 U879 ( .A1(n1048), .A2(n1196), .A3(n1214), .A4(n1055), .ZN(n1188) );
XNOR2_X1 U880 ( .A(G101), .B(n1181), .ZN(G3) );
NAND3_X1 U881 ( .A1(n1046), .A2(n1178), .A3(n1032), .ZN(n1181) );
XOR2_X1 U882 ( .A(G125), .B(n1184), .Z(G27) );
AND4_X1 U883 ( .A1(n1027), .A2(n1036), .A3(n1196), .A4(n1202), .ZN(n1184) );
AND3_X1 U884 ( .A1(n1203), .A2(n1201), .A3(n1041), .ZN(n1196) );
NAND2_X1 U885 ( .A1(n1015), .A2(n1215), .ZN(n1201) );
NAND4_X1 U886 ( .A1(G953), .A2(G902), .A3(n1216), .A4(n1078), .ZN(n1215) );
INV_X1 U887 ( .A(G900), .ZN(n1078) );
INV_X1 U888 ( .A(n1047), .ZN(n1203) );
XOR2_X1 U889 ( .A(n1217), .B(n1180), .Z(G24) );
NAND4_X1 U890 ( .A1(n1218), .A2(n1064), .A3(n1199), .A4(n1200), .ZN(n1180) );
INV_X1 U891 ( .A(n1020), .ZN(n1064) );
NAND2_X1 U892 ( .A1(n1047), .A2(n1202), .ZN(n1020) );
NAND2_X1 U893 ( .A1(n1219), .A2(n1220), .ZN(G21) );
OR2_X1 U894 ( .A1(n1221), .A2(G119), .ZN(n1220) );
NAND2_X1 U895 ( .A1(n1222), .A2(G119), .ZN(n1219) );
NAND2_X1 U896 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
OR2_X1 U897 ( .A1(n1179), .A2(KEYINPUT17), .ZN(n1224) );
NAND2_X1 U898 ( .A1(KEYINPUT17), .A2(n1221), .ZN(n1223) );
NAND2_X1 U899 ( .A1(KEYINPUT26), .A2(n1225), .ZN(n1221) );
INV_X1 U900 ( .A(n1179), .ZN(n1225) );
NAND3_X1 U901 ( .A1(n1048), .A2(n1205), .A3(n1218), .ZN(n1179) );
XOR2_X1 U902 ( .A(n1177), .B(n1226), .Z(G18) );
NAND2_X1 U903 ( .A1(KEYINPUT28), .A2(G116), .ZN(n1226) );
NAND3_X1 U904 ( .A1(n1046), .A2(n1055), .A3(n1218), .ZN(n1177) );
NOR2_X1 U905 ( .A1(n1200), .A2(n1227), .ZN(n1055) );
XNOR2_X1 U906 ( .A(G113), .B(n1176), .ZN(G15) );
NAND3_X1 U907 ( .A1(n1046), .A2(n1027), .A3(n1218), .ZN(n1176) );
AND2_X1 U908 ( .A1(n1036), .A2(n1228), .ZN(n1218) );
NOR2_X1 U909 ( .A1(n1031), .A2(n1229), .ZN(n1036) );
XOR2_X1 U910 ( .A(KEYINPUT19), .B(n1030), .Z(n1229) );
AND2_X1 U911 ( .A1(n1227), .A2(n1200), .ZN(n1027) );
INV_X1 U912 ( .A(n1199), .ZN(n1227) );
INV_X1 U913 ( .A(n1208), .ZN(n1046) );
NAND2_X1 U914 ( .A1(n1048), .A2(n1047), .ZN(n1208) );
XNOR2_X1 U915 ( .A(G110), .B(n1175), .ZN(G12) );
NAND3_X1 U916 ( .A1(n1178), .A2(n1202), .A3(n1205), .ZN(n1175) );
NOR2_X1 U917 ( .A1(n1034), .A2(n1047), .ZN(n1205) );
XOR2_X1 U918 ( .A(n1230), .B(n1115), .Z(n1047) );
AND2_X1 U919 ( .A1(G217), .A2(n1231), .ZN(n1115) );
NAND2_X1 U920 ( .A1(n1117), .A2(n1194), .ZN(n1230) );
XOR2_X1 U921 ( .A(n1232), .B(n1233), .Z(n1117) );
XOR2_X1 U922 ( .A(n1207), .B(n1234), .Z(n1233) );
NAND2_X1 U923 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NAND4_X1 U924 ( .A1(n1079), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1236) );
NAND2_X1 U925 ( .A1(n1240), .A2(n1195), .ZN(n1239) );
NAND2_X1 U926 ( .A1(G146), .A2(n1241), .ZN(n1238) );
NAND3_X1 U927 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1235) );
NAND2_X1 U928 ( .A1(n1079), .A2(n1237), .ZN(n1244) );
INV_X1 U929 ( .A(KEYINPUT61), .ZN(n1237) );
NAND2_X1 U930 ( .A1(n1241), .A2(n1195), .ZN(n1243) );
XOR2_X1 U931 ( .A(n1245), .B(KEYINPUT25), .Z(n1241) );
NAND2_X1 U932 ( .A1(G146), .A2(n1240), .ZN(n1242) );
XOR2_X1 U933 ( .A(n1245), .B(KEYINPUT36), .Z(n1240) );
XOR2_X1 U934 ( .A(n1246), .B(G110), .Z(n1245) );
NAND2_X1 U935 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND2_X1 U936 ( .A1(G119), .A2(n1213), .ZN(n1248) );
XOR2_X1 U937 ( .A(KEYINPUT56), .B(n1249), .Z(n1247) );
NOR2_X1 U938 ( .A1(G119), .A2(n1213), .ZN(n1249) );
INV_X1 U939 ( .A(G128), .ZN(n1213) );
INV_X1 U940 ( .A(G137), .ZN(n1207) );
NAND2_X1 U941 ( .A1(G221), .A2(n1250), .ZN(n1232) );
INV_X1 U942 ( .A(n1032), .ZN(n1034) );
NOR2_X1 U943 ( .A1(n1200), .A2(n1199), .ZN(n1032) );
XOR2_X1 U944 ( .A(n1251), .B(n1068), .Z(n1199) );
NOR2_X1 U945 ( .A1(n1119), .A2(G902), .ZN(n1068) );
XOR2_X1 U946 ( .A(n1252), .B(n1253), .Z(n1119) );
NOR2_X1 U947 ( .A1(KEYINPUT50), .A2(n1254), .ZN(n1253) );
XOR2_X1 U948 ( .A(n1255), .B(n1256), .Z(n1254) );
XOR2_X1 U949 ( .A(n1257), .B(n1258), .Z(n1256) );
XOR2_X1 U950 ( .A(n1259), .B(G107), .Z(n1257) );
NAND2_X1 U951 ( .A1(KEYINPUT32), .A2(n1260), .ZN(n1259) );
XOR2_X1 U952 ( .A(G122), .B(G116), .Z(n1260) );
XOR2_X1 U953 ( .A(n1261), .B(G134), .Z(n1255) );
XNOR2_X1 U954 ( .A(KEYINPUT49), .B(KEYINPUT35), .ZN(n1261) );
NAND2_X1 U955 ( .A1(G217), .A2(n1250), .ZN(n1252) );
AND2_X1 U956 ( .A1(G234), .A2(n1072), .ZN(n1250) );
NAND2_X1 U957 ( .A1(KEYINPUT9), .A2(n1122), .ZN(n1251) );
INV_X1 U958 ( .A(G478), .ZN(n1122) );
NAND2_X1 U959 ( .A1(n1262), .A2(n1066), .ZN(n1200) );
NAND3_X1 U960 ( .A1(n1127), .A2(n1194), .A3(n1126), .ZN(n1066) );
INV_X1 U961 ( .A(G475), .ZN(n1127) );
XNOR2_X1 U962 ( .A(KEYINPUT16), .B(n1065), .ZN(n1262) );
NAND2_X1 U963 ( .A1(G475), .A2(n1263), .ZN(n1065) );
NAND2_X1 U964 ( .A1(n1126), .A2(n1194), .ZN(n1263) );
XOR2_X1 U965 ( .A(n1264), .B(n1265), .Z(n1126) );
XNOR2_X1 U966 ( .A(n1266), .B(n1267), .ZN(n1265) );
NOR2_X1 U967 ( .A1(KEYINPUT12), .A2(n1128), .ZN(n1267) );
NAND2_X1 U968 ( .A1(n1268), .A2(KEYINPUT18), .ZN(n1266) );
XOR2_X1 U969 ( .A(n1269), .B(n1270), .Z(n1268) );
XOR2_X1 U970 ( .A(KEYINPUT40), .B(G146), .Z(n1270) );
XOR2_X1 U971 ( .A(n1271), .B(n1079), .Z(n1269) );
XOR2_X1 U972 ( .A(G140), .B(n1272), .Z(n1079) );
NAND2_X1 U973 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
NAND2_X1 U974 ( .A1(n1275), .A2(n1084), .ZN(n1274) );
XOR2_X1 U975 ( .A(KEYINPUT15), .B(n1276), .Z(n1273) );
NOR2_X1 U976 ( .A1(n1275), .A2(n1084), .ZN(n1276) );
XOR2_X1 U977 ( .A(n1277), .B(n1278), .Z(n1275) );
NOR2_X1 U978 ( .A1(n1279), .A2(G143), .ZN(n1278) );
INV_X1 U979 ( .A(KEYINPUT8), .ZN(n1279) );
NAND2_X1 U980 ( .A1(n1280), .A2(n1281), .ZN(n1277) );
XOR2_X1 U981 ( .A(KEYINPUT48), .B(G214), .Z(n1281) );
XOR2_X1 U982 ( .A(G113), .B(n1217), .Z(n1264) );
INV_X1 U983 ( .A(G122), .ZN(n1217) );
INV_X1 U984 ( .A(n1048), .ZN(n1202) );
XOR2_X1 U985 ( .A(n1282), .B(n1283), .Z(n1048) );
XOR2_X1 U986 ( .A(KEYINPUT24), .B(G472), .Z(n1283) );
NAND2_X1 U987 ( .A1(n1284), .A2(n1194), .ZN(n1282) );
XOR2_X1 U988 ( .A(KEYINPUT5), .B(n1285), .Z(n1284) );
INV_X1 U989 ( .A(n1131), .ZN(n1285) );
XOR2_X1 U990 ( .A(n1286), .B(n1287), .Z(n1131) );
XOR2_X1 U991 ( .A(n1159), .B(n1288), .Z(n1287) );
XOR2_X1 U992 ( .A(n1289), .B(G113), .Z(n1288) );
NAND2_X1 U993 ( .A1(KEYINPUT22), .A2(n1290), .ZN(n1289) );
XOR2_X1 U994 ( .A(n1291), .B(n1292), .Z(n1286) );
AND2_X1 U995 ( .A1(n1280), .A2(G210), .ZN(n1292) );
NOR2_X1 U996 ( .A1(G953), .A2(G237), .ZN(n1280) );
AND2_X1 U997 ( .A1(n1228), .A2(n1214), .ZN(n1178) );
XOR2_X1 U998 ( .A(n1033), .B(KEYINPUT33), .Z(n1214) );
NAND2_X1 U999 ( .A1(n1030), .A2(n1031), .ZN(n1033) );
NAND2_X1 U1000 ( .A1(n1293), .A2(n1294), .ZN(n1031) );
NAND2_X1 U1001 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
INV_X1 U1002 ( .A(G469), .ZN(n1296) );
XNOR2_X1 U1003 ( .A(KEYINPUT39), .B(n1061), .ZN(n1295) );
XOR2_X1 U1004 ( .A(KEYINPUT41), .B(n1060), .Z(n1293) );
AND2_X1 U1005 ( .A1(G469), .A2(n1061), .ZN(n1060) );
NAND2_X1 U1006 ( .A1(n1297), .A2(n1194), .ZN(n1061) );
XOR2_X1 U1007 ( .A(n1298), .B(n1299), .Z(n1297) );
NOR2_X1 U1008 ( .A1(n1152), .A2(n1147), .ZN(n1299) );
AND2_X1 U1009 ( .A1(n1150), .A2(n1300), .ZN(n1147) );
NOR2_X1 U1010 ( .A1(n1300), .A2(n1150), .ZN(n1152) );
XOR2_X1 U1011 ( .A(G140), .B(G110), .Z(n1150) );
NAND2_X1 U1012 ( .A1(G227), .A2(n1072), .ZN(n1300) );
NAND2_X1 U1013 ( .A1(n1301), .A2(n1302), .ZN(n1298) );
NAND2_X1 U1014 ( .A1(n1145), .A2(n1159), .ZN(n1302) );
XOR2_X1 U1015 ( .A(KEYINPUT14), .B(n1303), .Z(n1301) );
NOR2_X1 U1016 ( .A1(n1145), .A2(n1159), .ZN(n1303) );
NAND3_X1 U1017 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n1159) );
NAND2_X1 U1018 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NAND2_X1 U1019 ( .A1(KEYINPUT52), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1020 ( .A(KEYINPUT45), .B(G131), .Z(n1309) );
NAND3_X1 U1021 ( .A1(KEYINPUT52), .A2(n1086), .A3(n1084), .ZN(n1305) );
INV_X1 U1022 ( .A(n1307), .ZN(n1086) );
XOR2_X1 U1023 ( .A(G134), .B(G137), .Z(n1307) );
OR2_X1 U1024 ( .A1(n1084), .A2(KEYINPUT52), .ZN(n1304) );
INV_X1 U1025 ( .A(G131), .ZN(n1084) );
XOR2_X1 U1026 ( .A(n1310), .B(n1311), .Z(n1145) );
XOR2_X1 U1027 ( .A(KEYINPUT62), .B(G107), .Z(n1311) );
XOR2_X1 U1028 ( .A(n1291), .B(n1312), .Z(n1310) );
NOR2_X1 U1029 ( .A1(KEYINPUT60), .A2(n1128), .ZN(n1312) );
INV_X1 U1030 ( .A(G104), .ZN(n1128) );
NAND2_X1 U1031 ( .A1(G221), .A2(n1231), .ZN(n1030) );
NAND2_X1 U1032 ( .A1(n1313), .A2(n1194), .ZN(n1231) );
AND2_X1 U1033 ( .A1(n1041), .A2(n1314), .ZN(n1228) );
NAND2_X1 U1034 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND4_X1 U1035 ( .A1(G953), .A2(G902), .A3(n1216), .A4(n1108), .ZN(n1316) );
INV_X1 U1036 ( .A(G898), .ZN(n1108) );
XNOR2_X1 U1037 ( .A(KEYINPUT57), .B(n1015), .ZN(n1315) );
NAND3_X1 U1038 ( .A1(n1216), .A2(n1072), .A3(G952), .ZN(n1015) );
NAND2_X1 U1039 ( .A1(G237), .A2(n1313), .ZN(n1216) );
XOR2_X1 U1040 ( .A(G234), .B(KEYINPUT42), .Z(n1313) );
AND2_X1 U1041 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U1042 ( .A1(G214), .A2(n1317), .ZN(n1043) );
INV_X1 U1043 ( .A(n1212), .ZN(n1042) );
XNOR2_X1 U1044 ( .A(n1318), .B(n1170), .ZN(n1212) );
NAND2_X1 U1045 ( .A1(G210), .A2(n1317), .ZN(n1170) );
NAND2_X1 U1046 ( .A1(n1194), .A2(n1319), .ZN(n1317) );
INV_X1 U1047 ( .A(G237), .ZN(n1319) );
INV_X1 U1048 ( .A(G902), .ZN(n1194) );
OR2_X1 U1049 ( .A1(n1169), .A2(G902), .ZN(n1318) );
XNOR2_X1 U1050 ( .A(n1320), .B(n1321), .ZN(n1169) );
XOR2_X1 U1051 ( .A(n1107), .B(n1105), .Z(n1321) );
XOR2_X1 U1052 ( .A(G110), .B(n1322), .Z(n1105) );
XOR2_X1 U1053 ( .A(KEYINPUT53), .B(G122), .Z(n1322) );
XNOR2_X1 U1054 ( .A(n1323), .B(n1324), .ZN(n1107) );
NOR2_X1 U1055 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NOR2_X1 U1056 ( .A1(KEYINPUT1), .A2(n1327), .ZN(n1326) );
AND2_X1 U1057 ( .A1(KEYINPUT10), .A2(n1327), .ZN(n1325) );
AND3_X1 U1058 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1327) );
NAND2_X1 U1059 ( .A1(KEYINPUT2), .A2(G104), .ZN(n1330) );
OR4_X1 U1060 ( .A1(KEYINPUT13), .A2(KEYINPUT2), .A3(G104), .A4(G107), .ZN(n1329) );
NAND2_X1 U1061 ( .A1(G107), .A2(n1331), .ZN(n1328) );
OR2_X1 U1062 ( .A1(G104), .A2(KEYINPUT13), .ZN(n1331) );
NAND2_X1 U1063 ( .A1(n1332), .A2(n1333), .ZN(n1323) );
NAND2_X1 U1064 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
INV_X1 U1065 ( .A(KEYINPUT23), .ZN(n1335) );
XNOR2_X1 U1066 ( .A(G113), .B(n1290), .ZN(n1334) );
XOR2_X1 U1067 ( .A(G116), .B(G119), .Z(n1290) );
NAND2_X1 U1068 ( .A1(n1336), .A2(KEYINPUT23), .ZN(n1332) );
XNOR2_X1 U1069 ( .A(G113), .B(n1337), .ZN(n1336) );
NAND2_X1 U1070 ( .A1(G119), .A2(n1338), .ZN(n1337) );
INV_X1 U1071 ( .A(G116), .ZN(n1338) );
XOR2_X1 U1072 ( .A(n1339), .B(n1272), .Z(n1320) );
XOR2_X1 U1073 ( .A(G125), .B(KEYINPUT51), .Z(n1272) );
XOR2_X1 U1074 ( .A(n1291), .B(n1340), .Z(n1339) );
AND2_X1 U1075 ( .A1(n1072), .A2(G224), .ZN(n1340) );
INV_X1 U1076 ( .A(G953), .ZN(n1072) );
XOR2_X1 U1077 ( .A(n1082), .B(G101), .Z(n1291) );
XOR2_X1 U1078 ( .A(n1195), .B(n1258), .Z(n1082) );
XOR2_X1 U1079 ( .A(G143), .B(G128), .Z(n1258) );
INV_X1 U1080 ( .A(G146), .ZN(n1195) );
endmodule


