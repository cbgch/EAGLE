//Key = 0110010010111100001011010010111000100111100110110010000111101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413, n1414;

XOR2_X1 U765 ( .A(G107), .B(n1072), .Z(G9) );
NOR2_X1 U766 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(G75) );
NOR4_X1 U768 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1076) );
INV_X1 U769 ( .A(G952), .ZN(n1079) );
NAND4_X1 U770 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1077) );
NAND4_X1 U771 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1082) );
AND3_X1 U772 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
OR2_X1 U773 ( .A1(n1092), .A2(n1093), .ZN(n1086) );
OR3_X1 U774 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1085) );
NAND3_X1 U775 ( .A1(n1093), .A2(n1097), .A3(n1087), .ZN(n1081) );
INV_X1 U776 ( .A(n1098), .ZN(n1087) );
NAND2_X1 U777 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NAND3_X1 U778 ( .A1(n1101), .A2(n1090), .A3(n1091), .ZN(n1100) );
NAND2_X1 U779 ( .A1(n1102), .A2(n1103), .ZN(n1099) );
NAND2_X1 U780 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U781 ( .A1(n1091), .A2(n1106), .ZN(n1105) );
NAND2_X1 U782 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U783 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
INV_X1 U784 ( .A(n1111), .ZN(n1107) );
NAND2_X1 U785 ( .A1(n1090), .A2(n1112), .ZN(n1104) );
NAND2_X1 U786 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND2_X1 U787 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR3_X1 U788 ( .A1(n1117), .A2(G953), .A3(n1118), .ZN(n1075) );
INV_X1 U789 ( .A(n1083), .ZN(n1118) );
NAND4_X1 U790 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1083) );
NOR4_X1 U791 ( .A1(n1096), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1122) );
XOR2_X1 U792 ( .A(n1126), .B(n1127), .Z(n1123) );
NOR2_X1 U793 ( .A1(G472), .A2(n1128), .ZN(n1127) );
XNOR2_X1 U794 ( .A(KEYINPUT33), .B(KEYINPUT1), .ZN(n1128) );
XOR2_X1 U795 ( .A(n1129), .B(n1130), .Z(n1121) );
NOR2_X1 U796 ( .A1(KEYINPUT16), .A2(n1131), .ZN(n1130) );
XNOR2_X1 U797 ( .A(G478), .B(KEYINPUT46), .ZN(n1129) );
XOR2_X1 U798 ( .A(n1132), .B(KEYINPUT8), .Z(n1120) );
NAND3_X1 U799 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
NAND2_X1 U800 ( .A1(G469), .A2(n1136), .ZN(n1135) );
NAND2_X1 U801 ( .A1(KEYINPUT61), .A2(n1137), .ZN(n1134) );
NAND2_X1 U802 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
INV_X1 U803 ( .A(G469), .ZN(n1139) );
XNOR2_X1 U804 ( .A(KEYINPUT45), .B(n1136), .ZN(n1138) );
NAND2_X1 U805 ( .A1(n1140), .A2(n1141), .ZN(n1133) );
INV_X1 U806 ( .A(KEYINPUT61), .ZN(n1141) );
NAND2_X1 U807 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
OR3_X1 U808 ( .A1(n1136), .A2(G469), .A3(KEYINPUT45), .ZN(n1143) );
NAND2_X1 U809 ( .A1(KEYINPUT45), .A2(n1136), .ZN(n1142) );
XNOR2_X1 U810 ( .A(n1144), .B(n1145), .ZN(n1119) );
NAND2_X1 U811 ( .A1(KEYINPUT43), .A2(n1146), .ZN(n1144) );
XNOR2_X1 U812 ( .A(G952), .B(KEYINPUT40), .ZN(n1117) );
XOR2_X1 U813 ( .A(n1147), .B(n1148), .Z(G72) );
NOR2_X1 U814 ( .A1(n1149), .A2(n1084), .ZN(n1148) );
NOR2_X1 U815 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XNOR2_X1 U816 ( .A(KEYINPUT10), .B(n1152), .ZN(n1151) );
INV_X1 U817 ( .A(G227), .ZN(n1150) );
NAND2_X1 U818 ( .A1(n1153), .A2(n1154), .ZN(n1147) );
NAND2_X1 U819 ( .A1(n1155), .A2(n1084), .ZN(n1154) );
XOR2_X1 U820 ( .A(n1156), .B(n1080), .Z(n1155) );
NAND3_X1 U821 ( .A1(G900), .A2(n1156), .A3(G953), .ZN(n1153) );
XNOR2_X1 U822 ( .A(n1157), .B(n1158), .ZN(n1156) );
XOR2_X1 U823 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U824 ( .A(G134), .B(G125), .Z(n1160) );
XOR2_X1 U825 ( .A(KEYINPUT5), .B(KEYINPUT31), .Z(n1159) );
XNOR2_X1 U826 ( .A(n1161), .B(n1162), .ZN(n1157) );
XOR2_X1 U827 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U828 ( .A1(G140), .A2(KEYINPUT52), .ZN(n1163) );
XOR2_X1 U829 ( .A(n1165), .B(n1166), .Z(G69) );
NOR2_X1 U830 ( .A1(n1167), .A2(n1084), .ZN(n1166) );
AND2_X1 U831 ( .A1(G224), .A2(G898), .ZN(n1167) );
NAND2_X1 U832 ( .A1(n1168), .A2(n1169), .ZN(n1165) );
NAND2_X1 U833 ( .A1(n1170), .A2(n1084), .ZN(n1169) );
XOR2_X1 U834 ( .A(n1171), .B(n1078), .Z(n1170) );
NAND3_X1 U835 ( .A1(G898), .A2(n1171), .A3(G953), .ZN(n1168) );
XOR2_X1 U836 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U837 ( .A(n1174), .B(KEYINPUT51), .Z(n1172) );
NOR2_X1 U838 ( .A1(n1175), .A2(n1176), .ZN(G66) );
XNOR2_X1 U839 ( .A(n1177), .B(n1178), .ZN(n1176) );
NOR2_X1 U840 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NOR2_X1 U841 ( .A1(n1181), .A2(n1182), .ZN(G63) );
XOR2_X1 U842 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U843 ( .A(KEYINPUT18), .B(n1185), .Z(n1184) );
NOR2_X1 U844 ( .A1(n1186), .A2(n1180), .ZN(n1185) );
NOR2_X1 U845 ( .A1(G952), .A2(n1187), .ZN(n1181) );
XNOR2_X1 U846 ( .A(G953), .B(KEYINPUT17), .ZN(n1187) );
NOR2_X1 U847 ( .A1(n1175), .A2(n1188), .ZN(G60) );
XNOR2_X1 U848 ( .A(n1189), .B(n1190), .ZN(n1188) );
AND2_X1 U849 ( .A1(G475), .A2(n1191), .ZN(n1190) );
XNOR2_X1 U850 ( .A(G104), .B(n1192), .ZN(G6) );
NAND2_X1 U851 ( .A1(KEYINPUT60), .A2(n1193), .ZN(n1192) );
INV_X1 U852 ( .A(n1194), .ZN(n1193) );
NOR2_X1 U853 ( .A1(n1175), .A2(n1195), .ZN(G57) );
XOR2_X1 U854 ( .A(n1196), .B(n1197), .Z(n1195) );
XOR2_X1 U855 ( .A(n1198), .B(n1199), .Z(n1197) );
XNOR2_X1 U856 ( .A(n1200), .B(n1201), .ZN(n1198) );
NAND3_X1 U857 ( .A1(n1191), .A2(G472), .A3(KEYINPUT26), .ZN(n1200) );
XOR2_X1 U858 ( .A(n1202), .B(n1203), .Z(n1196) );
NOR2_X1 U859 ( .A1(KEYINPUT14), .A2(n1204), .ZN(n1203) );
XNOR2_X1 U860 ( .A(n1205), .B(n1206), .ZN(n1204) );
XNOR2_X1 U861 ( .A(G101), .B(KEYINPUT4), .ZN(n1202) );
NOR2_X1 U862 ( .A1(n1175), .A2(n1207), .ZN(G54) );
XOR2_X1 U863 ( .A(n1208), .B(n1209), .Z(n1207) );
XNOR2_X1 U864 ( .A(n1210), .B(KEYINPUT41), .ZN(n1209) );
NAND3_X1 U865 ( .A1(n1191), .A2(G469), .A3(KEYINPUT38), .ZN(n1210) );
XOR2_X1 U866 ( .A(n1211), .B(n1212), .Z(n1208) );
NOR2_X1 U867 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XOR2_X1 U868 ( .A(n1215), .B(KEYINPUT63), .Z(n1214) );
NAND2_X1 U869 ( .A1(n1206), .A2(n1216), .ZN(n1215) );
NOR2_X1 U870 ( .A1(n1175), .A2(n1217), .ZN(G51) );
XOR2_X1 U871 ( .A(n1218), .B(n1219), .Z(n1217) );
NOR2_X1 U872 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NOR2_X1 U873 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NOR2_X1 U874 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
INV_X1 U875 ( .A(KEYINPUT29), .ZN(n1225) );
NOR2_X1 U876 ( .A1(n1226), .A2(n1227), .ZN(n1224) );
XOR2_X1 U877 ( .A(KEYINPUT44), .B(n1228), .Z(n1227) );
AND2_X1 U878 ( .A1(KEYINPUT29), .A2(n1222), .ZN(n1220) );
NOR2_X1 U879 ( .A1(n1228), .A2(n1229), .ZN(n1222) );
XNOR2_X1 U880 ( .A(n1230), .B(n1231), .ZN(n1228) );
NAND2_X1 U881 ( .A1(KEYINPUT20), .A2(n1232), .ZN(n1218) );
NAND2_X1 U882 ( .A1(n1191), .A2(n1233), .ZN(n1232) );
INV_X1 U883 ( .A(n1180), .ZN(n1191) );
NAND2_X1 U884 ( .A1(G902), .A2(n1234), .ZN(n1180) );
OR2_X1 U885 ( .A1(n1078), .A2(n1080), .ZN(n1234) );
NAND2_X1 U886 ( .A1(n1235), .A2(n1236), .ZN(n1080) );
NOR4_X1 U887 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1236) );
NOR4_X1 U888 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1235) );
NOR2_X1 U889 ( .A1(n1124), .A2(n1245), .ZN(n1244) );
INV_X1 U890 ( .A(n1246), .ZN(n1243) );
INV_X1 U891 ( .A(n1247), .ZN(n1242) );
NAND4_X1 U892 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1078) );
AND4_X1 U893 ( .A1(n1252), .A2(n1253), .A3(n1194), .A4(n1254), .ZN(n1251) );
NAND3_X1 U894 ( .A1(n1255), .A2(n1090), .A3(n1095), .ZN(n1194) );
AND2_X1 U895 ( .A1(n1256), .A2(n1257), .ZN(n1250) );
NAND2_X1 U896 ( .A1(n1258), .A2(n1259), .ZN(n1248) );
XOR2_X1 U897 ( .A(n1073), .B(KEYINPUT11), .Z(n1258) );
NAND4_X1 U898 ( .A1(n1101), .A2(n1094), .A3(n1090), .A4(n1260), .ZN(n1073) );
NOR2_X1 U899 ( .A1(n1084), .A2(G952), .ZN(n1175) );
XOR2_X1 U900 ( .A(G146), .B(n1241), .Z(G48) );
AND3_X1 U901 ( .A1(n1095), .A2(n1261), .A3(n1262), .ZN(n1241) );
XNOR2_X1 U902 ( .A(G143), .B(n1246), .ZN(G45) );
NAND4_X1 U903 ( .A1(n1101), .A2(n1261), .A3(n1111), .A4(n1263), .ZN(n1246) );
AND3_X1 U904 ( .A1(n1125), .A2(n1264), .A3(n1265), .ZN(n1263) );
XOR2_X1 U905 ( .A(G140), .B(n1266), .Z(G42) );
NOR2_X1 U906 ( .A1(n1267), .A2(n1124), .ZN(n1266) );
XOR2_X1 U907 ( .A(n1245), .B(KEYINPUT35), .Z(n1267) );
NAND3_X1 U908 ( .A1(n1095), .A2(n1264), .A3(n1268), .ZN(n1245) );
XOR2_X1 U909 ( .A(n1269), .B(G137), .Z(G39) );
NAND2_X1 U910 ( .A1(KEYINPUT34), .A2(n1247), .ZN(n1269) );
NAND3_X1 U911 ( .A1(n1093), .A2(n1091), .A3(n1262), .ZN(n1247) );
XOR2_X1 U912 ( .A(G134), .B(n1240), .Z(G36) );
AND2_X1 U913 ( .A1(n1270), .A2(n1094), .ZN(n1240) );
XOR2_X1 U914 ( .A(G131), .B(n1239), .Z(G33) );
AND2_X1 U915 ( .A1(n1270), .A2(n1095), .ZN(n1239) );
AND4_X1 U916 ( .A1(n1111), .A2(n1091), .A3(n1101), .A4(n1264), .ZN(n1270) );
INV_X1 U917 ( .A(n1124), .ZN(n1091) );
NAND2_X1 U918 ( .A1(n1116), .A2(n1271), .ZN(n1124) );
XOR2_X1 U919 ( .A(G128), .B(n1238), .Z(G30) );
AND3_X1 U920 ( .A1(n1094), .A2(n1261), .A3(n1262), .ZN(n1238) );
AND4_X1 U921 ( .A1(n1101), .A2(n1272), .A3(n1110), .A4(n1264), .ZN(n1262) );
XNOR2_X1 U922 ( .A(G101), .B(n1253), .ZN(G3) );
NAND3_X1 U923 ( .A1(n1255), .A2(n1111), .A3(n1093), .ZN(n1253) );
AND3_X1 U924 ( .A1(n1101), .A2(n1260), .A3(n1259), .ZN(n1255) );
XOR2_X1 U925 ( .A(G125), .B(n1237), .Z(G27) );
AND4_X1 U926 ( .A1(n1109), .A2(n1102), .A3(n1095), .A4(n1273), .ZN(n1237) );
AND3_X1 U927 ( .A1(n1261), .A2(n1264), .A3(n1110), .ZN(n1273) );
NAND2_X1 U928 ( .A1(n1098), .A2(n1274), .ZN(n1264) );
NAND4_X1 U929 ( .A1(G953), .A2(G902), .A3(n1275), .A4(n1152), .ZN(n1274) );
INV_X1 U930 ( .A(G900), .ZN(n1152) );
INV_X1 U931 ( .A(n1276), .ZN(n1102) );
XNOR2_X1 U932 ( .A(G122), .B(n1252), .ZN(G24) );
NAND4_X1 U933 ( .A1(n1277), .A2(n1090), .A3(n1125), .A4(n1265), .ZN(n1252) );
NOR2_X1 U934 ( .A1(n1110), .A2(n1272), .ZN(n1090) );
XNOR2_X1 U935 ( .A(G119), .B(n1249), .ZN(G21) );
NAND4_X1 U936 ( .A1(n1093), .A2(n1277), .A3(n1272), .A4(n1110), .ZN(n1249) );
XNOR2_X1 U937 ( .A(n1278), .B(n1279), .ZN(G18) );
NOR2_X1 U938 ( .A1(KEYINPUT48), .A2(n1257), .ZN(n1279) );
NAND3_X1 U939 ( .A1(n1277), .A2(n1094), .A3(n1111), .ZN(n1257) );
AND2_X1 U940 ( .A1(n1280), .A2(n1265), .ZN(n1094) );
NOR3_X1 U941 ( .A1(n1113), .A2(n1281), .A3(n1276), .ZN(n1277) );
INV_X1 U942 ( .A(n1261), .ZN(n1113) );
XOR2_X1 U943 ( .A(n1259), .B(KEYINPUT0), .Z(n1261) );
XNOR2_X1 U944 ( .A(G113), .B(n1256), .ZN(G15) );
NAND3_X1 U945 ( .A1(n1095), .A2(n1111), .A3(n1282), .ZN(n1256) );
NOR3_X1 U946 ( .A1(n1276), .A2(n1281), .A3(n1074), .ZN(n1282) );
INV_X1 U947 ( .A(n1259), .ZN(n1074) );
INV_X1 U948 ( .A(n1260), .ZN(n1281) );
NAND2_X1 U949 ( .A1(n1089), .A2(n1092), .ZN(n1276) );
NOR2_X1 U950 ( .A1(n1110), .A2(n1109), .ZN(n1111) );
NOR2_X1 U951 ( .A1(n1265), .A2(n1280), .ZN(n1095) );
INV_X1 U952 ( .A(n1125), .ZN(n1280) );
XNOR2_X1 U953 ( .A(G110), .B(n1254), .ZN(G12) );
NAND4_X1 U954 ( .A1(n1268), .A2(n1093), .A3(n1259), .A4(n1260), .ZN(n1254) );
NAND2_X1 U955 ( .A1(n1098), .A2(n1283), .ZN(n1260) );
NAND4_X1 U956 ( .A1(G953), .A2(G902), .A3(n1275), .A4(n1284), .ZN(n1283) );
INV_X1 U957 ( .A(G898), .ZN(n1284) );
NAND3_X1 U958 ( .A1(n1275), .A2(n1084), .A3(G952), .ZN(n1098) );
NAND2_X1 U959 ( .A1(G237), .A2(G234), .ZN(n1275) );
NOR2_X1 U960 ( .A1(n1116), .A2(n1115), .ZN(n1259) );
INV_X1 U961 ( .A(n1271), .ZN(n1115) );
NAND2_X1 U962 ( .A1(G214), .A2(n1285), .ZN(n1271) );
XOR2_X1 U963 ( .A(n1286), .B(n1233), .Z(n1116) );
AND2_X1 U964 ( .A1(G210), .A2(n1285), .ZN(n1233) );
NAND2_X1 U965 ( .A1(n1287), .A2(n1288), .ZN(n1285) );
INV_X1 U966 ( .A(G237), .ZN(n1287) );
NAND2_X1 U967 ( .A1(n1289), .A2(n1290), .ZN(n1286) );
XOR2_X1 U968 ( .A(n1291), .B(n1292), .Z(n1289) );
XOR2_X1 U969 ( .A(n1230), .B(n1293), .Z(n1292) );
NOR2_X1 U970 ( .A1(KEYINPUT6), .A2(n1231), .ZN(n1293) );
XNOR2_X1 U971 ( .A(n1294), .B(G125), .ZN(n1231) );
INV_X1 U972 ( .A(n1205), .ZN(n1294) );
NAND2_X1 U973 ( .A1(G224), .A2(n1084), .ZN(n1230) );
NAND2_X1 U974 ( .A1(KEYINPUT37), .A2(n1229), .ZN(n1291) );
INV_X1 U975 ( .A(n1226), .ZN(n1229) );
XNOR2_X1 U976 ( .A(n1174), .B(n1295), .ZN(n1226) );
XNOR2_X1 U977 ( .A(n1296), .B(KEYINPUT50), .ZN(n1295) );
NAND2_X1 U978 ( .A1(KEYINPUT47), .A2(n1173), .ZN(n1296) );
XNOR2_X1 U979 ( .A(G110), .B(G122), .ZN(n1173) );
XOR2_X1 U980 ( .A(n1297), .B(n1298), .Z(n1174) );
XOR2_X1 U981 ( .A(n1299), .B(n1300), .Z(n1298) );
XNOR2_X1 U982 ( .A(n1278), .B(G113), .ZN(n1300) );
XNOR2_X1 U983 ( .A(KEYINPUT39), .B(n1301), .ZN(n1299) );
XNOR2_X1 U984 ( .A(n1302), .B(n1303), .ZN(n1297) );
XNOR2_X1 U985 ( .A(n1304), .B(n1305), .ZN(n1302) );
NAND2_X1 U986 ( .A1(KEYINPUT30), .A2(n1306), .ZN(n1304) );
INV_X1 U987 ( .A(G104), .ZN(n1306) );
NOR2_X1 U988 ( .A1(n1265), .A2(n1125), .ZN(n1093) );
XNOR2_X1 U989 ( .A(n1307), .B(G475), .ZN(n1125) );
NAND2_X1 U990 ( .A1(n1189), .A2(n1290), .ZN(n1307) );
XNOR2_X1 U991 ( .A(n1308), .B(n1309), .ZN(n1189) );
XOR2_X1 U992 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U993 ( .A(n1312), .B(G131), .ZN(n1311) );
NOR2_X1 U994 ( .A1(KEYINPUT22), .A2(n1313), .ZN(n1310) );
NOR2_X1 U995 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
XOR2_X1 U996 ( .A(KEYINPUT25), .B(n1316), .Z(n1315) );
AND2_X1 U997 ( .A1(n1317), .A2(G104), .ZN(n1316) );
NOR2_X1 U998 ( .A1(G104), .A2(n1317), .ZN(n1314) );
NAND3_X1 U999 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1317) );
NAND2_X1 U1000 ( .A1(G113), .A2(n1321), .ZN(n1320) );
NAND2_X1 U1001 ( .A1(KEYINPUT54), .A2(n1322), .ZN(n1319) );
NAND2_X1 U1002 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
INV_X1 U1003 ( .A(n1321), .ZN(n1324) );
XNOR2_X1 U1004 ( .A(KEYINPUT36), .B(G113), .ZN(n1323) );
NAND2_X1 U1005 ( .A1(n1325), .A2(n1326), .ZN(n1318) );
INV_X1 U1006 ( .A(KEYINPUT54), .ZN(n1326) );
NAND2_X1 U1007 ( .A1(n1327), .A2(n1328), .ZN(n1325) );
OR3_X1 U1008 ( .A1(n1321), .A2(G113), .A3(KEYINPUT36), .ZN(n1328) );
XOR2_X1 U1009 ( .A(G122), .B(KEYINPUT28), .Z(n1321) );
NAND2_X1 U1010 ( .A1(KEYINPUT36), .A2(G113), .ZN(n1327) );
XOR2_X1 U1011 ( .A(n1329), .B(n1330), .Z(n1308) );
NAND2_X1 U1012 ( .A1(n1331), .A2(G214), .ZN(n1329) );
XOR2_X1 U1013 ( .A(n1131), .B(n1332), .Z(n1265) );
XNOR2_X1 U1014 ( .A(KEYINPUT53), .B(n1186), .ZN(n1332) );
INV_X1 U1015 ( .A(G478), .ZN(n1186) );
AND2_X1 U1016 ( .A1(n1290), .A2(n1183), .ZN(n1131) );
NAND2_X1 U1017 ( .A1(n1333), .A2(n1334), .ZN(n1183) );
NAND4_X1 U1018 ( .A1(n1335), .A2(G217), .A3(n1336), .A4(G234), .ZN(n1334) );
AND2_X1 U1019 ( .A1(n1084), .A2(n1337), .ZN(n1336) );
NAND2_X1 U1020 ( .A1(n1338), .A2(n1339), .ZN(n1333) );
NAND3_X1 U1021 ( .A1(G234), .A2(n1084), .A3(G217), .ZN(n1339) );
NAND2_X1 U1022 ( .A1(n1335), .A2(n1337), .ZN(n1338) );
NAND2_X1 U1023 ( .A1(n1340), .A2(n1341), .ZN(n1337) );
XOR2_X1 U1024 ( .A(n1342), .B(n1343), .Z(n1340) );
XOR2_X1 U1025 ( .A(n1344), .B(KEYINPUT7), .Z(n1335) );
NAND2_X1 U1026 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
XNOR2_X1 U1027 ( .A(n1342), .B(n1343), .ZN(n1346) );
XOR2_X1 U1028 ( .A(G128), .B(G134), .Z(n1343) );
NAND2_X1 U1029 ( .A1(KEYINPUT13), .A2(n1312), .ZN(n1342) );
INV_X1 U1030 ( .A(G143), .ZN(n1312) );
INV_X1 U1031 ( .A(n1341), .ZN(n1345) );
NAND2_X1 U1032 ( .A1(n1347), .A2(n1348), .ZN(n1341) );
NAND2_X1 U1033 ( .A1(n1303), .A2(n1349), .ZN(n1348) );
XOR2_X1 U1034 ( .A(n1350), .B(KEYINPUT62), .Z(n1347) );
OR2_X1 U1035 ( .A1(n1349), .A2(n1303), .ZN(n1350) );
XNOR2_X1 U1036 ( .A(G122), .B(n1278), .ZN(n1349) );
AND3_X1 U1037 ( .A1(n1109), .A2(n1110), .A3(n1101), .ZN(n1268) );
NOR2_X1 U1038 ( .A1(n1089), .A2(n1096), .ZN(n1101) );
INV_X1 U1039 ( .A(n1092), .ZN(n1096) );
NAND2_X1 U1040 ( .A1(G221), .A2(n1351), .ZN(n1092) );
XOR2_X1 U1041 ( .A(n1136), .B(n1352), .Z(n1089) );
XOR2_X1 U1042 ( .A(KEYINPUT23), .B(n1353), .Z(n1352) );
NOR2_X1 U1043 ( .A1(KEYINPUT42), .A2(G469), .ZN(n1353) );
NAND2_X1 U1044 ( .A1(n1354), .A2(n1290), .ZN(n1136) );
XOR2_X1 U1045 ( .A(n1355), .B(n1211), .Z(n1354) );
XOR2_X1 U1046 ( .A(n1356), .B(n1357), .Z(n1211) );
XOR2_X1 U1047 ( .A(G140), .B(G110), .Z(n1357) );
NAND2_X1 U1048 ( .A1(G227), .A2(n1084), .ZN(n1356) );
NAND3_X1 U1049 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1355) );
NAND2_X1 U1050 ( .A1(n1213), .A2(n1361), .ZN(n1360) );
INV_X1 U1051 ( .A(KEYINPUT49), .ZN(n1361) );
NOR2_X1 U1052 ( .A1(n1216), .A2(n1206), .ZN(n1213) );
OR2_X1 U1053 ( .A1(n1362), .A2(n1363), .ZN(n1216) );
AND2_X1 U1054 ( .A1(n1364), .A2(n1161), .ZN(n1363) );
NAND3_X1 U1055 ( .A1(n1362), .A2(KEYINPUT49), .A3(n1365), .ZN(n1359) );
NAND2_X1 U1056 ( .A1(n1206), .A2(n1366), .ZN(n1358) );
NAND2_X1 U1057 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
NAND2_X1 U1058 ( .A1(n1364), .A2(n1161), .ZN(n1368) );
XNOR2_X1 U1059 ( .A(n1362), .B(KEYINPUT49), .ZN(n1367) );
NOR2_X1 U1060 ( .A1(n1161), .A2(n1364), .ZN(n1362) );
XOR2_X1 U1061 ( .A(n1369), .B(n1303), .Z(n1364) );
XNOR2_X1 U1062 ( .A(G107), .B(KEYINPUT57), .ZN(n1303) );
XNOR2_X1 U1063 ( .A(n1370), .B(n1305), .ZN(n1369) );
NAND2_X1 U1064 ( .A1(KEYINPUT56), .A2(G104), .ZN(n1370) );
XNOR2_X1 U1065 ( .A(n1371), .B(n1372), .ZN(n1161) );
NAND2_X1 U1066 ( .A1(KEYINPUT55), .A2(G128), .ZN(n1371) );
XNOR2_X1 U1067 ( .A(n1145), .B(n1146), .ZN(n1110) );
INV_X1 U1068 ( .A(n1179), .ZN(n1146) );
NAND2_X1 U1069 ( .A1(G217), .A2(n1351), .ZN(n1179) );
NAND2_X1 U1070 ( .A1(G234), .A2(n1288), .ZN(n1351) );
NAND2_X1 U1071 ( .A1(n1290), .A2(n1177), .ZN(n1145) );
NAND3_X1 U1072 ( .A1(n1373), .A2(n1374), .A3(n1375), .ZN(n1177) );
NAND2_X1 U1073 ( .A1(n1376), .A2(n1377), .ZN(n1375) );
NAND2_X1 U1074 ( .A1(n1378), .A2(n1379), .ZN(n1374) );
INV_X1 U1075 ( .A(KEYINPUT58), .ZN(n1379) );
NAND2_X1 U1076 ( .A1(n1380), .A2(n1381), .ZN(n1378) );
XNOR2_X1 U1077 ( .A(n1376), .B(KEYINPUT27), .ZN(n1380) );
NAND2_X1 U1078 ( .A1(KEYINPUT58), .A2(n1382), .ZN(n1373) );
NAND2_X1 U1079 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
OR3_X1 U1080 ( .A1(n1377), .A2(KEYINPUT27), .A3(n1376), .ZN(n1384) );
INV_X1 U1081 ( .A(n1381), .ZN(n1377) );
XNOR2_X1 U1082 ( .A(n1385), .B(G137), .ZN(n1381) );
NAND3_X1 U1083 ( .A1(G234), .A2(n1084), .A3(G221), .ZN(n1385) );
INV_X1 U1084 ( .A(G953), .ZN(n1084) );
NAND2_X1 U1085 ( .A1(KEYINPUT27), .A2(n1376), .ZN(n1383) );
XNOR2_X1 U1086 ( .A(n1386), .B(n1387), .ZN(n1376) );
XNOR2_X1 U1087 ( .A(G128), .B(n1301), .ZN(n1387) );
NAND2_X1 U1088 ( .A1(n1388), .A2(n1389), .ZN(n1386) );
NAND2_X1 U1089 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
INV_X1 U1090 ( .A(KEYINPUT19), .ZN(n1391) );
XOR2_X1 U1091 ( .A(G110), .B(n1330), .Z(n1390) );
XNOR2_X1 U1092 ( .A(n1392), .B(n1393), .ZN(n1330) );
NAND2_X1 U1093 ( .A1(KEYINPUT19), .A2(n1394), .ZN(n1388) );
XOR2_X1 U1094 ( .A(n1395), .B(G110), .Z(n1394) );
NAND2_X1 U1095 ( .A1(n1392), .A2(n1393), .ZN(n1395) );
XOR2_X1 U1096 ( .A(G125), .B(G140), .Z(n1393) );
INV_X1 U1097 ( .A(n1272), .ZN(n1109) );
XNOR2_X1 U1098 ( .A(n1126), .B(G472), .ZN(n1272) );
NAND2_X1 U1099 ( .A1(n1396), .A2(n1290), .ZN(n1126) );
XNOR2_X1 U1100 ( .A(n1288), .B(KEYINPUT2), .ZN(n1290) );
INV_X1 U1101 ( .A(G902), .ZN(n1288) );
XOR2_X1 U1102 ( .A(n1397), .B(n1398), .Z(n1396) );
XNOR2_X1 U1103 ( .A(n1365), .B(n1199), .ZN(n1398) );
XOR2_X1 U1104 ( .A(n1399), .B(n1400), .Z(n1199) );
INV_X1 U1105 ( .A(G113), .ZN(n1400) );
NAND3_X1 U1106 ( .A1(n1401), .A2(n1402), .A3(n1403), .ZN(n1399) );
NAND2_X1 U1107 ( .A1(n1404), .A2(n1301), .ZN(n1403) );
INV_X1 U1108 ( .A(G119), .ZN(n1301) );
NAND2_X1 U1109 ( .A1(n1405), .A2(n1406), .ZN(n1404) );
XNOR2_X1 U1110 ( .A(G116), .B(KEYINPUT9), .ZN(n1405) );
NAND3_X1 U1111 ( .A1(G119), .A2(n1278), .A3(n1406), .ZN(n1402) );
INV_X1 U1112 ( .A(KEYINPUT15), .ZN(n1406) );
INV_X1 U1113 ( .A(G116), .ZN(n1278) );
NAND2_X1 U1114 ( .A1(G116), .A2(KEYINPUT15), .ZN(n1401) );
INV_X1 U1115 ( .A(n1206), .ZN(n1365) );
XOR2_X1 U1116 ( .A(n1164), .B(n1407), .Z(n1206) );
NOR2_X1 U1117 ( .A1(G134), .A2(KEYINPUT59), .ZN(n1407) );
XOR2_X1 U1118 ( .A(G131), .B(G137), .Z(n1164) );
XOR2_X1 U1119 ( .A(n1408), .B(n1409), .Z(n1397) );
XNOR2_X1 U1120 ( .A(KEYINPUT24), .B(n1410), .ZN(n1409) );
NOR2_X1 U1121 ( .A1(KEYINPUT3), .A2(n1411), .ZN(n1410) );
NOR2_X1 U1122 ( .A1(n1412), .A2(n1413), .ZN(n1411) );
XOR2_X1 U1123 ( .A(KEYINPUT32), .B(n1414), .Z(n1413) );
AND2_X1 U1124 ( .A1(n1201), .A2(n1305), .ZN(n1414) );
NOR2_X1 U1125 ( .A1(n1305), .A2(n1201), .ZN(n1412) );
NAND2_X1 U1126 ( .A1(n1331), .A2(G210), .ZN(n1201) );
NOR2_X1 U1127 ( .A1(G953), .A2(G237), .ZN(n1331) );
INV_X1 U1128 ( .A(G101), .ZN(n1305) );
NAND2_X1 U1129 ( .A1(KEYINPUT12), .A2(n1205), .ZN(n1408) );
XOR2_X1 U1130 ( .A(n1372), .B(G128), .Z(n1205) );
XNOR2_X1 U1131 ( .A(G143), .B(n1392), .ZN(n1372) );
XNOR2_X1 U1132 ( .A(G146), .B(KEYINPUT21), .ZN(n1392) );
endmodule


