//Key = 0111111100110011011111011101001000010001000100111100000011001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357;

XOR2_X1 U743 ( .A(n1028), .B(G107), .Z(G9) );
NAND2_X1 U744 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND2_X1 U745 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
INV_X1 U746 ( .A(KEYINPUT16), .ZN(n1032) );
NAND3_X1 U747 ( .A1(n1033), .A2(n1034), .A3(KEYINPUT16), .ZN(n1029) );
NOR2_X1 U748 ( .A1(n1035), .A2(n1036), .ZN(G75) );
NOR4_X1 U749 ( .A1(n1037), .A2(n1038), .A3(G953), .A4(n1039), .ZN(n1036) );
AND3_X1 U750 ( .A1(KEYINPUT39), .A2(n1040), .A3(n1041), .ZN(n1038) );
OR2_X1 U751 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U753 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U754 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U755 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR3_X1 U756 ( .A1(n1052), .A2(n1034), .A3(n1053), .ZN(n1051) );
NOR2_X1 U757 ( .A1(n1054), .A2(n1055), .ZN(n1050) );
AND3_X1 U758 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1046) );
AND3_X1 U759 ( .A1(n1056), .A2(n1059), .A3(n1060), .ZN(n1042) );
NAND2_X1 U760 ( .A1(n1061), .A2(n1062), .ZN(n1037) );
XOR2_X1 U761 ( .A(n1063), .B(KEYINPUT51), .Z(n1061) );
NAND3_X1 U762 ( .A1(n1064), .A2(n1040), .A3(KEYINPUT39), .ZN(n1063) );
NAND2_X1 U763 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND3_X1 U764 ( .A1(n1060), .A2(n1067), .A3(n1056), .ZN(n1066) );
NAND2_X1 U765 ( .A1(n1068), .A2(n1069), .ZN(n1065) );
NAND2_X1 U766 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U767 ( .A1(n1056), .A2(n1072), .ZN(n1071) );
NOR2_X1 U768 ( .A1(n1054), .A2(n1034), .ZN(n1056) );
NAND2_X1 U769 ( .A1(n1060), .A2(n1073), .ZN(n1070) );
NAND2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XNOR2_X1 U772 ( .A(n1078), .B(KEYINPUT62), .ZN(n1076) );
NAND2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1074) );
NOR3_X1 U774 ( .A1(n1039), .A2(G953), .A3(G952), .ZN(n1035) );
AND4_X1 U775 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1039) );
NOR4_X1 U776 ( .A1(n1057), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1084) );
XOR2_X1 U777 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U778 ( .A1(KEYINPUT17), .A2(n1090), .ZN(n1088) );
XOR2_X1 U779 ( .A(n1091), .B(n1092), .Z(n1086) );
NAND2_X1 U780 ( .A1(KEYINPUT43), .A2(n1093), .ZN(n1091) );
NOR2_X1 U781 ( .A1(n1094), .A2(n1095), .ZN(n1083) );
XNOR2_X1 U782 ( .A(n1096), .B(n1097), .ZN(n1095) );
XNOR2_X1 U783 ( .A(n1098), .B(n1099), .ZN(n1094) );
XOR2_X1 U784 ( .A(n1100), .B(n1101), .Z(n1082) );
XNOR2_X1 U785 ( .A(G472), .B(KEYINPUT1), .ZN(n1101) );
NAND2_X1 U786 ( .A1(n1102), .A2(KEYINPUT7), .ZN(n1100) );
XOR2_X1 U787 ( .A(n1103), .B(KEYINPUT35), .Z(n1102) );
XOR2_X1 U788 ( .A(KEYINPUT14), .B(n1104), .Z(n1081) );
XOR2_X1 U789 ( .A(n1105), .B(n1106), .Z(G72) );
XOR2_X1 U790 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR3_X1 U791 ( .A1(n1109), .A2(KEYINPUT44), .A3(G953), .ZN(n1108) );
INV_X1 U792 ( .A(n1110), .ZN(n1109) );
NOR2_X1 U793 ( .A1(n1111), .A2(n1112), .ZN(n1107) );
XOR2_X1 U794 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U795 ( .A(n1115), .B(n1116), .Z(n1114) );
XNOR2_X1 U796 ( .A(G125), .B(KEYINPUT0), .ZN(n1113) );
NOR2_X1 U797 ( .A1(G900), .A2(n1117), .ZN(n1111) );
XNOR2_X1 U798 ( .A(n1118), .B(KEYINPUT50), .ZN(n1117) );
NOR2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1105) );
NOR2_X1 U800 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
XOR2_X1 U801 ( .A(n1123), .B(n1124), .Z(G69) );
XOR2_X1 U802 ( .A(n1125), .B(n1126), .Z(n1124) );
OR2_X1 U803 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U804 ( .A1(n1129), .A2(n1120), .ZN(n1125) );
NOR2_X1 U805 ( .A1(n1130), .A2(n1120), .ZN(n1123) );
AND2_X1 U806 ( .A1(G224), .A2(G898), .ZN(n1130) );
NOR2_X1 U807 ( .A1(n1131), .A2(n1132), .ZN(G66) );
NOR3_X1 U808 ( .A1(n1098), .A2(n1133), .A3(n1134), .ZN(n1132) );
NOR3_X1 U809 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1134) );
INV_X1 U810 ( .A(n1138), .ZN(n1135) );
NOR2_X1 U811 ( .A1(n1139), .A2(n1138), .ZN(n1133) );
NOR2_X1 U812 ( .A1(n1062), .A2(n1136), .ZN(n1139) );
NOR2_X1 U813 ( .A1(n1131), .A2(n1140), .ZN(G63) );
NOR3_X1 U814 ( .A1(n1092), .A2(n1141), .A3(n1142), .ZN(n1140) );
NOR3_X1 U815 ( .A1(n1143), .A2(n1093), .A3(n1137), .ZN(n1142) );
INV_X1 U816 ( .A(n1144), .ZN(n1143) );
NOR2_X1 U817 ( .A1(n1145), .A2(n1144), .ZN(n1141) );
NOR2_X1 U818 ( .A1(n1062), .A2(n1093), .ZN(n1145) );
INV_X1 U819 ( .A(G478), .ZN(n1093) );
NOR2_X1 U820 ( .A1(n1131), .A2(n1146), .ZN(G60) );
NOR3_X1 U821 ( .A1(n1089), .A2(n1147), .A3(n1148), .ZN(n1146) );
NOR3_X1 U822 ( .A1(n1149), .A2(n1090), .A3(n1137), .ZN(n1148) );
INV_X1 U823 ( .A(n1150), .ZN(n1149) );
NOR2_X1 U824 ( .A1(n1151), .A2(n1150), .ZN(n1147) );
NOR2_X1 U825 ( .A1(n1062), .A2(n1090), .ZN(n1151) );
XNOR2_X1 U826 ( .A(G104), .B(n1152), .ZN(G6) );
NAND2_X1 U827 ( .A1(n1153), .A2(n1080), .ZN(n1152) );
XOR2_X1 U828 ( .A(n1154), .B(KEYINPUT10), .Z(n1153) );
NOR2_X1 U829 ( .A1(n1155), .A2(n1156), .ZN(G57) );
XOR2_X1 U830 ( .A(KEYINPUT38), .B(n1131), .Z(n1156) );
XOR2_X1 U831 ( .A(n1157), .B(n1158), .Z(n1155) );
NOR2_X1 U832 ( .A1(n1159), .A2(n1137), .ZN(n1158) );
NOR2_X1 U833 ( .A1(n1131), .A2(n1160), .ZN(G54) );
XOR2_X1 U834 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U835 ( .A(n1115), .B(n1163), .Z(n1162) );
XOR2_X1 U836 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U837 ( .A1(n1166), .A2(n1137), .ZN(n1165) );
NAND2_X1 U838 ( .A1(G902), .A2(n1167), .ZN(n1137) );
NAND2_X1 U839 ( .A1(KEYINPUT46), .A2(n1116), .ZN(n1164) );
XNOR2_X1 U840 ( .A(n1168), .B(n1169), .ZN(n1115) );
XOR2_X1 U841 ( .A(n1170), .B(n1171), .Z(n1161) );
XOR2_X1 U842 ( .A(n1172), .B(n1173), .Z(n1171) );
XNOR2_X1 U843 ( .A(G110), .B(KEYINPUT59), .ZN(n1170) );
NOR2_X1 U844 ( .A1(n1131), .A2(n1174), .ZN(G51) );
XOR2_X1 U845 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U846 ( .A(n1177), .B(n1178), .ZN(n1176) );
XOR2_X1 U847 ( .A(n1179), .B(n1180), .Z(n1175) );
XNOR2_X1 U848 ( .A(G125), .B(n1181), .ZN(n1180) );
NAND4_X1 U849 ( .A1(n1182), .A2(G210), .A3(n1167), .A4(n1183), .ZN(n1179) );
INV_X1 U850 ( .A(n1062), .ZN(n1167) );
NOR2_X1 U851 ( .A1(n1110), .A2(n1129), .ZN(n1062) );
NAND4_X1 U852 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1129) );
NOR4_X1 U853 ( .A1(n1188), .A2(n1031), .A3(n1189), .A4(n1190), .ZN(n1187) );
AND2_X1 U854 ( .A1(n1079), .A2(n1033), .ZN(n1031) );
AND3_X1 U855 ( .A1(n1059), .A2(n1191), .A3(n1072), .ZN(n1033) );
NOR2_X1 U856 ( .A1(n1192), .A2(n1193), .ZN(n1186) );
NOR2_X1 U857 ( .A1(n1194), .A2(n1154), .ZN(n1193) );
NAND4_X1 U858 ( .A1(n1067), .A2(n1079), .A3(n1072), .A4(n1195), .ZN(n1154) );
NOR2_X1 U859 ( .A1(n1080), .A2(n1196), .ZN(n1192) );
NAND4_X1 U860 ( .A1(KEYINPUT12), .A2(n1197), .A3(n1068), .A4(n1195), .ZN(n1196) );
NAND3_X1 U861 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1185) );
INV_X1 U862 ( .A(n1201), .ZN(n1200) );
OR2_X1 U863 ( .A1(n1202), .A2(KEYINPUT60), .ZN(n1199) );
NAND2_X1 U864 ( .A1(n1203), .A2(KEYINPUT60), .ZN(n1198) );
NAND2_X1 U865 ( .A1(n1204), .A2(n1205), .ZN(n1184) );
INV_X1 U866 ( .A(KEYINPUT12), .ZN(n1205) );
NAND4_X1 U867 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1110) );
NOR3_X1 U868 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1209) );
INV_X1 U869 ( .A(n1213), .ZN(n1212) );
NOR2_X1 U870 ( .A1(n1214), .A2(n1194), .ZN(n1210) );
NOR2_X1 U871 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NOR2_X1 U872 ( .A1(n1203), .A2(n1217), .ZN(n1216) );
NOR2_X1 U873 ( .A1(n1067), .A2(n1059), .ZN(n1203) );
NOR3_X1 U874 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1215) );
XOR2_X1 U875 ( .A(KEYINPUT5), .B(n1072), .Z(n1220) );
NAND3_X1 U876 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1218) );
XNOR2_X1 U877 ( .A(G902), .B(KEYINPUT49), .ZN(n1182) );
NOR2_X1 U878 ( .A1(n1120), .A2(G952), .ZN(n1131) );
XNOR2_X1 U879 ( .A(n1224), .B(n1225), .ZN(G48) );
NOR4_X1 U880 ( .A1(KEYINPUT54), .A2(n1226), .A3(n1217), .A4(n1202), .ZN(n1225) );
XNOR2_X1 U881 ( .A(n1080), .B(KEYINPUT13), .ZN(n1226) );
XNOR2_X1 U882 ( .A(G143), .B(n1227), .ZN(G45) );
NAND3_X1 U883 ( .A1(KEYINPUT30), .A2(n1228), .A3(n1229), .ZN(n1227) );
NOR3_X1 U884 ( .A1(n1194), .A2(n1230), .A3(n1231), .ZN(n1229) );
XNOR2_X1 U885 ( .A(G140), .B(n1213), .ZN(G42) );
NAND4_X1 U886 ( .A1(n1197), .A2(n1067), .A3(n1078), .A4(n1222), .ZN(n1213) );
AND2_X1 U887 ( .A1(n1232), .A2(n1072), .ZN(n1197) );
XNOR2_X1 U888 ( .A(n1233), .B(n1211), .ZN(G39) );
NOR3_X1 U889 ( .A1(n1045), .A2(n1217), .A3(n1054), .ZN(n1211) );
INV_X1 U890 ( .A(n1078), .ZN(n1054) );
NAND2_X1 U891 ( .A1(n1234), .A2(n1235), .ZN(G36) );
NAND2_X1 U892 ( .A1(G134), .A2(n1208), .ZN(n1235) );
XOR2_X1 U893 ( .A(KEYINPUT47), .B(n1236), .Z(n1234) );
NOR2_X1 U894 ( .A1(G134), .A2(n1208), .ZN(n1236) );
NAND3_X1 U895 ( .A1(n1078), .A2(n1059), .A3(n1228), .ZN(n1208) );
XNOR2_X1 U896 ( .A(n1237), .B(n1238), .ZN(G33) );
NOR2_X1 U897 ( .A1(KEYINPUT41), .A2(n1206), .ZN(n1238) );
NAND3_X1 U898 ( .A1(n1067), .A2(n1078), .A3(n1228), .ZN(n1206) );
AND3_X1 U899 ( .A1(n1072), .A2(n1222), .A3(n1077), .ZN(n1228) );
NOR2_X1 U900 ( .A1(n1053), .A2(n1085), .ZN(n1078) );
XOR2_X1 U901 ( .A(n1239), .B(n1240), .Z(G30) );
NOR4_X1 U902 ( .A1(KEYINPUT52), .A2(n1194), .A3(n1241), .A4(n1217), .ZN(n1240) );
NAND4_X1 U903 ( .A1(n1242), .A2(n1072), .A3(n1243), .A4(n1222), .ZN(n1217) );
INV_X1 U904 ( .A(n1080), .ZN(n1194) );
XNOR2_X1 U905 ( .A(G128), .B(KEYINPUT6), .ZN(n1239) );
XNOR2_X1 U906 ( .A(n1244), .B(n1190), .ZN(G3) );
AND2_X1 U907 ( .A1(n1245), .A2(n1077), .ZN(n1190) );
XNOR2_X1 U908 ( .A(G125), .B(n1207), .ZN(G27) );
NAND4_X1 U909 ( .A1(n1060), .A2(n1067), .A3(n1246), .A4(n1232), .ZN(n1207) );
AND2_X1 U910 ( .A1(n1222), .A2(n1080), .ZN(n1246) );
NAND2_X1 U911 ( .A1(n1247), .A2(n1248), .ZN(n1222) );
NAND4_X1 U912 ( .A1(n1118), .A2(n1249), .A3(n1040), .A4(n1122), .ZN(n1248) );
INV_X1 U913 ( .A(G900), .ZN(n1122) );
XOR2_X1 U914 ( .A(G122), .B(n1189), .Z(G24) );
AND4_X1 U915 ( .A1(n1060), .A2(n1079), .A3(n1250), .A4(n1191), .ZN(n1189) );
NOR2_X1 U916 ( .A1(n1230), .A2(n1231), .ZN(n1250) );
INV_X1 U917 ( .A(n1034), .ZN(n1079) );
NAND2_X1 U918 ( .A1(n1251), .A2(n1252), .ZN(n1034) );
XOR2_X1 U919 ( .A(G119), .B(n1188), .Z(G21) );
AND4_X1 U920 ( .A1(n1191), .A2(n1243), .A3(n1242), .A4(n1253), .ZN(n1188) );
NOR2_X1 U921 ( .A1(n1045), .A2(n1049), .ZN(n1253) );
INV_X1 U922 ( .A(n1068), .ZN(n1045) );
XOR2_X1 U923 ( .A(G116), .B(n1254), .Z(G18) );
NOR2_X1 U924 ( .A1(n1241), .A2(n1201), .ZN(n1254) );
INV_X1 U925 ( .A(n1059), .ZN(n1241) );
NOR2_X1 U926 ( .A1(n1231), .A2(n1221), .ZN(n1059) );
XOR2_X1 U927 ( .A(G113), .B(n1255), .Z(G15) );
NOR2_X1 U928 ( .A1(n1202), .A2(n1201), .ZN(n1255) );
NAND3_X1 U929 ( .A1(n1077), .A2(n1191), .A3(n1060), .ZN(n1201) );
INV_X1 U930 ( .A(n1049), .ZN(n1060) );
NAND2_X1 U931 ( .A1(n1058), .A2(n1256), .ZN(n1049) );
XOR2_X1 U932 ( .A(KEYINPUT25), .B(n1057), .Z(n1256) );
INV_X1 U933 ( .A(n1219), .ZN(n1077) );
NAND2_X1 U934 ( .A1(n1242), .A2(n1252), .ZN(n1219) );
XOR2_X1 U935 ( .A(n1243), .B(KEYINPUT21), .Z(n1252) );
INV_X1 U936 ( .A(n1251), .ZN(n1242) );
INV_X1 U937 ( .A(n1067), .ZN(n1202) );
NOR2_X1 U938 ( .A1(n1230), .A2(n1223), .ZN(n1067) );
XOR2_X1 U939 ( .A(n1204), .B(n1257), .Z(G12) );
NOR2_X1 U940 ( .A1(KEYINPUT32), .A2(n1258), .ZN(n1257) );
AND2_X1 U941 ( .A1(n1245), .A2(n1232), .ZN(n1204) );
INV_X1 U942 ( .A(n1055), .ZN(n1232) );
NAND2_X1 U943 ( .A1(n1251), .A2(n1243), .ZN(n1055) );
XOR2_X1 U944 ( .A(n1098), .B(n1259), .Z(n1243) );
NOR2_X1 U945 ( .A1(KEYINPUT8), .A2(n1099), .ZN(n1259) );
NAND2_X1 U946 ( .A1(G217), .A2(n1260), .ZN(n1099) );
XOR2_X1 U947 ( .A(KEYINPUT23), .B(n1261), .Z(n1260) );
AND2_X1 U948 ( .A1(n1262), .A2(G234), .ZN(n1261) );
NOR2_X1 U949 ( .A1(n1138), .A2(G902), .ZN(n1098) );
XNOR2_X1 U950 ( .A(n1263), .B(n1264), .ZN(n1138) );
XNOR2_X1 U951 ( .A(n1258), .B(n1265), .ZN(n1264) );
XNOR2_X1 U952 ( .A(n1266), .B(G119), .ZN(n1265) );
XOR2_X1 U953 ( .A(n1267), .B(n1268), .Z(n1263) );
NOR2_X1 U954 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
NOR2_X1 U955 ( .A1(n1271), .A2(G137), .ZN(n1270) );
NOR2_X1 U956 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NOR3_X1 U957 ( .A1(n1273), .A2(n1274), .A3(n1272), .ZN(n1269) );
XNOR2_X1 U958 ( .A(G137), .B(KEYINPUT37), .ZN(n1274) );
INV_X1 U959 ( .A(G221), .ZN(n1273) );
NAND2_X1 U960 ( .A1(KEYINPUT48), .A2(n1275), .ZN(n1267) );
XNOR2_X1 U961 ( .A(G146), .B(n1276), .ZN(n1275) );
NAND2_X1 U962 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND2_X1 U963 ( .A1(G125), .A2(n1169), .ZN(n1278) );
XOR2_X1 U964 ( .A(n1279), .B(KEYINPUT26), .Z(n1277) );
OR2_X1 U965 ( .A1(n1169), .A2(G125), .ZN(n1279) );
INV_X1 U966 ( .A(G140), .ZN(n1169) );
XOR2_X1 U967 ( .A(n1280), .B(n1103), .Z(n1251) );
NAND2_X1 U968 ( .A1(n1281), .A2(n1262), .ZN(n1103) );
XOR2_X1 U969 ( .A(n1157), .B(n1282), .Z(n1281) );
XOR2_X1 U970 ( .A(KEYINPUT42), .B(KEYINPUT11), .Z(n1282) );
XOR2_X1 U971 ( .A(n1283), .B(n1284), .Z(n1157) );
XOR2_X1 U972 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U973 ( .A(KEYINPUT56), .B(n1244), .ZN(n1286) );
AND3_X1 U974 ( .A1(G210), .A2(n1120), .A3(n1287), .ZN(n1285) );
XOR2_X1 U975 ( .A(n1288), .B(n1289), .Z(n1283) );
XNOR2_X1 U976 ( .A(n1168), .B(n1290), .ZN(n1288) );
INV_X1 U977 ( .A(n1177), .ZN(n1290) );
NAND2_X1 U978 ( .A1(KEYINPUT57), .A2(n1159), .ZN(n1280) );
INV_X1 U979 ( .A(G472), .ZN(n1159) );
AND3_X1 U980 ( .A1(n1072), .A2(n1191), .A3(n1068), .ZN(n1245) );
NOR2_X1 U981 ( .A1(n1221), .A2(n1223), .ZN(n1068) );
INV_X1 U982 ( .A(n1231), .ZN(n1223) );
XOR2_X1 U983 ( .A(G478), .B(n1291), .Z(n1231) );
NOR2_X1 U984 ( .A1(n1092), .A2(KEYINPUT55), .ZN(n1291) );
NOR2_X1 U985 ( .A1(n1144), .A2(G902), .ZN(n1092) );
XNOR2_X1 U986 ( .A(n1292), .B(n1293), .ZN(n1144) );
XOR2_X1 U987 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U988 ( .A(G107), .B(n1296), .ZN(n1295) );
NOR2_X1 U989 ( .A1(KEYINPUT33), .A2(n1297), .ZN(n1296) );
XOR2_X1 U990 ( .A(G116), .B(n1298), .Z(n1297) );
XOR2_X1 U991 ( .A(KEYINPUT15), .B(G122), .Z(n1298) );
NAND2_X1 U992 ( .A1(KEYINPUT3), .A2(n1299), .ZN(n1294) );
OR2_X1 U993 ( .A1(n1136), .A2(n1272), .ZN(n1299) );
NAND2_X1 U994 ( .A1(G234), .A2(n1120), .ZN(n1272) );
INV_X1 U995 ( .A(G217), .ZN(n1136) );
XNOR2_X1 U996 ( .A(G128), .B(n1300), .ZN(n1292) );
XOR2_X1 U997 ( .A(G143), .B(G134), .Z(n1300) );
INV_X1 U998 ( .A(n1230), .ZN(n1221) );
XOR2_X1 U999 ( .A(n1089), .B(n1090), .Z(n1230) );
INV_X1 U1000 ( .A(G475), .ZN(n1090) );
NOR2_X1 U1001 ( .A1(n1150), .A2(G902), .ZN(n1089) );
XNOR2_X1 U1002 ( .A(n1301), .B(G125), .ZN(n1150) );
XOR2_X1 U1003 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U1004 ( .A(n1304), .B(n1305), .Z(n1303) );
XOR2_X1 U1005 ( .A(G122), .B(G113), .Z(n1305) );
XNOR2_X1 U1006 ( .A(KEYINPUT9), .B(n1237), .ZN(n1304) );
INV_X1 U1007 ( .A(G131), .ZN(n1237) );
XOR2_X1 U1008 ( .A(n1306), .B(n1307), .Z(n1302) );
XOR2_X1 U1009 ( .A(n1308), .B(n1309), .Z(n1307) );
NOR2_X1 U1010 ( .A1(G140), .A2(KEYINPUT34), .ZN(n1308) );
XNOR2_X1 U1011 ( .A(G104), .B(n1310), .ZN(n1306) );
AND3_X1 U1012 ( .A1(G214), .A2(n1120), .A3(n1287), .ZN(n1310) );
AND2_X1 U1013 ( .A1(n1080), .A2(n1195), .ZN(n1191) );
NAND2_X1 U1014 ( .A1(n1311), .A2(n1312), .ZN(n1195) );
NAND3_X1 U1015 ( .A1(n1249), .A2(n1040), .A3(n1128), .ZN(n1312) );
NOR2_X1 U1016 ( .A1(n1313), .A2(G898), .ZN(n1128) );
INV_X1 U1017 ( .A(n1118), .ZN(n1313) );
XOR2_X1 U1018 ( .A(G953), .B(KEYINPUT58), .Z(n1118) );
XNOR2_X1 U1019 ( .A(n1262), .B(KEYINPUT45), .ZN(n1249) );
XOR2_X1 U1020 ( .A(n1247), .B(KEYINPUT53), .Z(n1311) );
NAND3_X1 U1021 ( .A1(n1040), .A2(n1120), .A3(G952), .ZN(n1247) );
NAND2_X1 U1022 ( .A1(G237), .A2(G234), .ZN(n1040) );
NOR2_X1 U1023 ( .A1(n1314), .A2(n1085), .ZN(n1080) );
INV_X1 U1024 ( .A(n1052), .ZN(n1085) );
NAND2_X1 U1025 ( .A1(G214), .A2(n1183), .ZN(n1052) );
INV_X1 U1026 ( .A(n1053), .ZN(n1314) );
XOR2_X1 U1027 ( .A(n1315), .B(n1097), .Z(n1053) );
NAND2_X1 U1028 ( .A1(G210), .A2(n1316), .ZN(n1097) );
XNOR2_X1 U1029 ( .A(KEYINPUT18), .B(n1183), .ZN(n1316) );
NAND2_X1 U1030 ( .A1(n1287), .A2(n1262), .ZN(n1183) );
INV_X1 U1031 ( .A(G237), .ZN(n1287) );
NAND2_X1 U1032 ( .A1(KEYINPUT4), .A2(n1096), .ZN(n1315) );
AND2_X1 U1033 ( .A1(n1317), .A2(n1262), .ZN(n1096) );
XNOR2_X1 U1034 ( .A(n1178), .B(n1318), .ZN(n1317) );
XNOR2_X1 U1035 ( .A(n1181), .B(n1319), .ZN(n1318) );
NAND2_X1 U1036 ( .A1(KEYINPUT63), .A2(n1320), .ZN(n1319) );
NAND2_X1 U1037 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NAND2_X1 U1038 ( .A1(n1323), .A2(G125), .ZN(n1322) );
XOR2_X1 U1039 ( .A(KEYINPUT27), .B(n1324), .Z(n1321) );
NOR2_X1 U1040 ( .A1(G125), .A2(n1323), .ZN(n1324) );
XNOR2_X1 U1041 ( .A(KEYINPUT24), .B(n1177), .ZN(n1323) );
XOR2_X1 U1042 ( .A(n1309), .B(n1325), .Z(n1177) );
NOR2_X1 U1043 ( .A1(G128), .A2(KEYINPUT36), .ZN(n1325) );
AND2_X1 U1044 ( .A1(G224), .A2(n1120), .ZN(n1181) );
INV_X1 U1045 ( .A(G953), .ZN(n1120) );
INV_X1 U1046 ( .A(n1127), .ZN(n1178) );
XNOR2_X1 U1047 ( .A(n1326), .B(n1327), .ZN(n1127) );
XNOR2_X1 U1048 ( .A(n1328), .B(n1289), .ZN(n1327) );
XOR2_X1 U1049 ( .A(G113), .B(n1329), .Z(n1289) );
XOR2_X1 U1050 ( .A(G119), .B(G116), .Z(n1329) );
NAND2_X1 U1051 ( .A1(n1330), .A2(n1331), .ZN(n1328) );
NAND2_X1 U1052 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
NAND2_X1 U1053 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NAND2_X1 U1054 ( .A1(G101), .A2(n1336), .ZN(n1335) );
INV_X1 U1055 ( .A(KEYINPUT22), .ZN(n1334) );
NAND2_X1 U1056 ( .A1(n1337), .A2(n1244), .ZN(n1330) );
NAND2_X1 U1057 ( .A1(n1336), .A2(n1338), .ZN(n1337) );
OR2_X1 U1058 ( .A1(n1332), .A2(KEYINPUT22), .ZN(n1338) );
INV_X1 U1059 ( .A(KEYINPUT31), .ZN(n1336) );
XNOR2_X1 U1060 ( .A(G122), .B(n1339), .ZN(n1326) );
NOR2_X1 U1061 ( .A1(G110), .A2(KEYINPUT61), .ZN(n1339) );
NOR2_X1 U1062 ( .A1(n1058), .A2(n1057), .ZN(n1072) );
AND2_X1 U1063 ( .A1(G221), .A2(n1340), .ZN(n1057) );
NAND2_X1 U1064 ( .A1(G234), .A2(n1262), .ZN(n1340) );
XNOR2_X1 U1065 ( .A(n1104), .B(KEYINPUT29), .ZN(n1058) );
XOR2_X1 U1066 ( .A(n1341), .B(n1166), .Z(n1104) );
INV_X1 U1067 ( .A(G469), .ZN(n1166) );
NAND2_X1 U1068 ( .A1(n1342), .A2(n1262), .ZN(n1341) );
INV_X1 U1069 ( .A(G902), .ZN(n1262) );
XOR2_X1 U1070 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1071 ( .A(n1116), .B(n1345), .Z(n1344) );
XOR2_X1 U1072 ( .A(n1172), .B(n1346), .Z(n1345) );
NAND2_X1 U1073 ( .A1(KEYINPUT20), .A2(n1168), .ZN(n1346) );
XNOR2_X1 U1074 ( .A(G131), .B(n1347), .ZN(n1168) );
XNOR2_X1 U1075 ( .A(n1233), .B(G134), .ZN(n1347) );
INV_X1 U1076 ( .A(G137), .ZN(n1233) );
NAND3_X1 U1077 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1172) );
NAND2_X1 U1078 ( .A1(KEYINPUT28), .A2(n1332), .ZN(n1350) );
NAND3_X1 U1079 ( .A1(n1351), .A2(n1352), .A3(n1244), .ZN(n1349) );
INV_X1 U1080 ( .A(KEYINPUT28), .ZN(n1352) );
OR2_X1 U1081 ( .A1(n1244), .A2(n1351), .ZN(n1348) );
NOR2_X1 U1082 ( .A1(KEYINPUT40), .A2(n1332), .ZN(n1351) );
XNOR2_X1 U1083 ( .A(G104), .B(G107), .ZN(n1332) );
INV_X1 U1084 ( .A(G101), .ZN(n1244) );
XNOR2_X1 U1085 ( .A(n1266), .B(n1309), .ZN(n1116) );
XNOR2_X1 U1086 ( .A(G143), .B(n1224), .ZN(n1309) );
INV_X1 U1087 ( .A(G146), .ZN(n1224) );
INV_X1 U1088 ( .A(G128), .ZN(n1266) );
XNOR2_X1 U1089 ( .A(n1173), .B(n1353), .ZN(n1343) );
XOR2_X1 U1090 ( .A(n1354), .B(KEYINPUT19), .Z(n1353) );
NAND2_X1 U1091 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
NAND2_X1 U1092 ( .A1(G140), .A2(n1258), .ZN(n1356) );
XOR2_X1 U1093 ( .A(KEYINPUT2), .B(n1357), .Z(n1355) );
NOR2_X1 U1094 ( .A1(G140), .A2(n1258), .ZN(n1357) );
INV_X1 U1095 ( .A(G110), .ZN(n1258) );
NOR2_X1 U1096 ( .A1(n1121), .A2(G953), .ZN(n1173) );
INV_X1 U1097 ( .A(G227), .ZN(n1121) );
endmodule


