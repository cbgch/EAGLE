//Key = 1111000110011000111000100100011100011001010010110101100111011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;

XNOR2_X1 U740 ( .A(G107), .B(n1019), .ZN(G9) );
NOR2_X1 U741 ( .A1(n1020), .A2(n1021), .ZN(G75) );
NOR4_X1 U742 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1021) );
NOR2_X1 U743 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR3_X1 U744 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1026) );
NOR2_X1 U745 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
INV_X1 U746 ( .A(n1033), .ZN(n1032) );
NOR4_X1 U747 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1031) );
NOR2_X1 U748 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
XOR2_X1 U749 ( .A(KEYINPUT31), .B(n1040), .Z(n1039) );
AND3_X1 U750 ( .A1(KEYINPUT47), .A2(n1040), .A3(n1041), .ZN(n1035) );
NOR2_X1 U751 ( .A1(n1042), .A2(n1043), .ZN(n1034) );
XOR2_X1 U752 ( .A(KEYINPUT55), .B(n1044), .Z(n1043) );
NOR3_X1 U753 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1029) );
NOR2_X1 U754 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U755 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR3_X1 U756 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1048) );
XOR2_X1 U757 ( .A(n1051), .B(KEYINPUT6), .Z(n1053) );
NOR2_X1 U758 ( .A1(KEYINPUT47), .A2(n1055), .ZN(n1028) );
NOR3_X1 U759 ( .A1(n1051), .A2(n1047), .A3(n1056), .ZN(n1055) );
INV_X1 U760 ( .A(n1057), .ZN(n1056) );
INV_X1 U761 ( .A(n1040), .ZN(n1047) );
NAND3_X1 U762 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1022) );
NAND4_X1 U763 ( .A1(n1033), .A2(n1044), .A3(n1040), .A4(n1061), .ZN(n1060) );
NAND2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
XOR2_X1 U766 ( .A(KEYINPUT41), .B(n1066), .Z(n1062) );
NOR3_X1 U767 ( .A1(n1052), .A2(n1067), .A3(n1051), .ZN(n1033) );
NOR3_X1 U768 ( .A1(n1068), .A2(G953), .A3(G952), .ZN(n1020) );
INV_X1 U769 ( .A(n1058), .ZN(n1068) );
NAND4_X1 U770 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1058) );
NOR4_X1 U771 ( .A1(n1073), .A2(n1074), .A3(n1027), .A4(n1075), .ZN(n1072) );
XOR2_X1 U772 ( .A(KEYINPUT27), .B(n1076), .Z(n1075) );
NOR2_X1 U773 ( .A1(n1077), .A2(n1067), .ZN(n1071) );
NAND2_X1 U774 ( .A1(G478), .A2(n1078), .ZN(n1070) );
XOR2_X1 U775 ( .A(n1079), .B(n1080), .Z(G72) );
NOR2_X1 U776 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U778 ( .A(n1085), .B(KEYINPUT0), .Z(n1084) );
NOR2_X1 U779 ( .A1(n1086), .A2(n1085), .ZN(n1081) );
NAND2_X1 U780 ( .A1(n1087), .A2(n1023), .ZN(n1085) );
XOR2_X1 U781 ( .A(KEYINPUT12), .B(G953), .Z(n1087) );
INV_X1 U782 ( .A(n1083), .ZN(n1086) );
NAND2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1083) );
NAND2_X1 U784 ( .A1(G953), .A2(n1090), .ZN(n1089) );
XOR2_X1 U785 ( .A(n1091), .B(n1092), .Z(n1088) );
XNOR2_X1 U786 ( .A(n1093), .B(n1094), .ZN(n1092) );
XNOR2_X1 U787 ( .A(n1095), .B(n1096), .ZN(n1091) );
NAND2_X1 U788 ( .A1(KEYINPUT49), .A2(n1097), .ZN(n1095) );
NAND2_X1 U789 ( .A1(G953), .A2(n1098), .ZN(n1079) );
NAND2_X1 U790 ( .A1(G900), .A2(G227), .ZN(n1098) );
XOR2_X1 U791 ( .A(n1099), .B(n1100), .Z(G69) );
NOR2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR3_X1 U793 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
NOR2_X1 U794 ( .A1(G224), .A2(n1059), .ZN(n1105) );
INV_X1 U795 ( .A(n1106), .ZN(n1103) );
NOR2_X1 U796 ( .A1(KEYINPUT8), .A2(n1106), .ZN(n1101) );
NAND3_X1 U797 ( .A1(n1107), .A2(n1108), .A3(n1059), .ZN(n1106) );
NAND2_X1 U798 ( .A1(KEYINPUT50), .A2(n1109), .ZN(n1108) );
OR2_X1 U799 ( .A1(n1025), .A2(KEYINPUT50), .ZN(n1107) );
NOR2_X1 U800 ( .A1(n1104), .A2(n1110), .ZN(n1099) );
XOR2_X1 U801 ( .A(KEYINPUT52), .B(n1111), .Z(n1110) );
NOR2_X1 U802 ( .A1(n1112), .A2(n1113), .ZN(G66) );
XOR2_X1 U803 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U804 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NOR2_X1 U805 ( .A1(n1112), .A2(n1118), .ZN(G63) );
XOR2_X1 U806 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U807 ( .A(n1121), .B(KEYINPUT53), .Z(n1119) );
NAND2_X1 U808 ( .A1(n1116), .A2(G478), .ZN(n1121) );
NOR2_X1 U809 ( .A1(n1122), .A2(n1123), .ZN(G60) );
XOR2_X1 U810 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND2_X1 U811 ( .A1(n1116), .A2(G475), .ZN(n1124) );
XNOR2_X1 U812 ( .A(n1112), .B(KEYINPUT56), .ZN(n1122) );
XNOR2_X1 U813 ( .A(G104), .B(n1126), .ZN(G6) );
NOR2_X1 U814 ( .A1(n1112), .A2(n1127), .ZN(G57) );
XOR2_X1 U815 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U816 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U817 ( .A1(KEYINPUT11), .A2(n1132), .ZN(n1130) );
XOR2_X1 U818 ( .A(n1133), .B(n1134), .Z(n1128) );
NOR3_X1 U819 ( .A1(n1135), .A2(KEYINPUT48), .A3(n1136), .ZN(n1134) );
INV_X1 U820 ( .A(G472), .ZN(n1136) );
XOR2_X1 U821 ( .A(n1137), .B(G101), .Z(n1133) );
NOR2_X1 U822 ( .A1(n1112), .A2(n1138), .ZN(G54) );
XOR2_X1 U823 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U824 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U825 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
NAND2_X1 U826 ( .A1(KEYINPUT38), .A2(n1145), .ZN(n1144) );
NAND2_X1 U827 ( .A1(KEYINPUT1), .A2(n1146), .ZN(n1143) );
INV_X1 U828 ( .A(n1145), .ZN(n1146) );
NAND2_X1 U829 ( .A1(n1116), .A2(G469), .ZN(n1145) );
XNOR2_X1 U830 ( .A(n1147), .B(n1132), .ZN(n1139) );
XNOR2_X1 U831 ( .A(n1148), .B(n1149), .ZN(n1147) );
NOR2_X1 U832 ( .A1(n1150), .A2(KEYINPUT62), .ZN(n1149) );
NOR2_X1 U833 ( .A1(KEYINPUT43), .A2(n1093), .ZN(n1148) );
NOR2_X1 U834 ( .A1(n1112), .A2(n1151), .ZN(G51) );
XOR2_X1 U835 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U836 ( .A1(KEYINPUT32), .A2(n1154), .ZN(n1153) );
XOR2_X1 U837 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U838 ( .A1(KEYINPUT20), .A2(n1157), .ZN(n1155) );
XOR2_X1 U839 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U840 ( .A1(G125), .A2(KEYINPUT13), .ZN(n1158) );
NAND2_X1 U841 ( .A1(n1116), .A2(G210), .ZN(n1152) );
INV_X1 U842 ( .A(n1135), .ZN(n1116) );
NAND2_X1 U843 ( .A1(G902), .A2(n1160), .ZN(n1135) );
NAND2_X1 U844 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XNOR2_X1 U845 ( .A(KEYINPUT40), .B(n1025), .ZN(n1162) );
NAND4_X1 U846 ( .A1(n1019), .A2(n1126), .A3(n1163), .A4(n1164), .ZN(n1025) );
NOR2_X1 U847 ( .A1(n1165), .A2(n1109), .ZN(n1164) );
NAND4_X1 U848 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1109) );
NAND3_X1 U849 ( .A1(n1040), .A2(n1170), .A3(n1041), .ZN(n1126) );
NAND3_X1 U850 ( .A1(n1040), .A2(n1170), .A3(n1171), .ZN(n1019) );
INV_X1 U851 ( .A(n1023), .ZN(n1161) );
NAND4_X1 U852 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1023) );
NOR3_X1 U853 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1175) );
NOR2_X1 U854 ( .A1(n1027), .A2(n1179), .ZN(n1176) );
XNOR2_X1 U855 ( .A(KEYINPUT51), .B(n1180), .ZN(n1179) );
NAND2_X1 U856 ( .A1(n1181), .A2(n1182), .ZN(n1174) );
NAND3_X1 U857 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1182) );
OR2_X1 U858 ( .A1(n1186), .A2(KEYINPUT34), .ZN(n1185) );
OR2_X1 U859 ( .A1(n1187), .A2(n1038), .ZN(n1184) );
NAND2_X1 U860 ( .A1(n1041), .A2(n1188), .ZN(n1183) );
NAND2_X1 U861 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U862 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U863 ( .A(n1027), .B(KEYINPUT25), .Z(n1191) );
NAND2_X1 U864 ( .A1(n1193), .A2(n1194), .ZN(n1189) );
NAND2_X1 U865 ( .A1(n1195), .A2(n1196), .ZN(n1173) );
NAND2_X1 U866 ( .A1(n1197), .A2(n1198), .ZN(n1195) );
NAND3_X1 U867 ( .A1(n1199), .A2(n1050), .A3(KEYINPUT34), .ZN(n1198) );
INV_X1 U868 ( .A(n1186), .ZN(n1199) );
OR2_X1 U869 ( .A1(n1200), .A2(KEYINPUT26), .ZN(n1197) );
NAND3_X1 U870 ( .A1(KEYINPUT26), .A2(n1201), .A3(n1202), .ZN(n1172) );
INV_X1 U871 ( .A(n1200), .ZN(n1201) );
NOR2_X1 U872 ( .A1(n1059), .A2(G952), .ZN(n1112) );
XOR2_X1 U873 ( .A(G146), .B(n1178), .Z(G48) );
NOR3_X1 U874 ( .A1(n1203), .A2(n1204), .A3(n1187), .ZN(n1178) );
XOR2_X1 U875 ( .A(G143), .B(n1205), .Z(G45) );
NOR2_X1 U876 ( .A1(n1204), .A2(n1186), .ZN(n1205) );
NAND4_X1 U877 ( .A1(n1193), .A2(n1066), .A3(n1206), .A4(n1207), .ZN(n1186) );
NAND2_X1 U878 ( .A1(n1208), .A2(n1209), .ZN(G42) );
OR2_X1 U879 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U880 ( .A(n1212), .B(KEYINPUT61), .Z(n1208) );
NAND2_X1 U881 ( .A1(n1211), .A2(n1210), .ZN(n1212) );
NOR4_X1 U882 ( .A1(n1042), .A2(n1203), .A3(n1204), .A4(n1027), .ZN(n1211) );
XOR2_X1 U883 ( .A(G137), .B(n1213), .Z(G39) );
NOR3_X1 U884 ( .A1(n1180), .A2(KEYINPUT9), .A3(n1027), .ZN(n1213) );
INV_X1 U885 ( .A(n1194), .ZN(n1027) );
NAND2_X1 U886 ( .A1(n1214), .A2(n1181), .ZN(n1180) );
XOR2_X1 U887 ( .A(G134), .B(n1177), .Z(G36) );
NOR2_X1 U888 ( .A1(n1215), .A2(n1038), .ZN(n1177) );
XOR2_X1 U889 ( .A(G131), .B(n1216), .Z(G33) );
NOR2_X1 U890 ( .A1(n1217), .A2(n1215), .ZN(n1216) );
NAND3_X1 U891 ( .A1(n1193), .A2(n1194), .A3(n1181), .ZN(n1215) );
NOR2_X1 U892 ( .A1(n1218), .A2(n1064), .ZN(n1194) );
XOR2_X1 U893 ( .A(n1203), .B(KEYINPUT21), .Z(n1217) );
XOR2_X1 U894 ( .A(G128), .B(n1219), .Z(G30) );
NOR4_X1 U895 ( .A1(KEYINPUT58), .A2(n1038), .A3(n1204), .A4(n1187), .ZN(n1219) );
NAND3_X1 U896 ( .A1(n1066), .A2(n1220), .A3(n1221), .ZN(n1187) );
INV_X1 U897 ( .A(n1181), .ZN(n1204) );
NOR2_X1 U898 ( .A1(n1050), .A2(n1202), .ZN(n1181) );
NAND2_X1 U899 ( .A1(n1222), .A2(n1223), .ZN(G3) );
NAND2_X1 U900 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
XNOR2_X1 U901 ( .A(n1165), .B(KEYINPUT22), .ZN(n1224) );
NAND2_X1 U902 ( .A1(G101), .A2(n1226), .ZN(n1222) );
XNOR2_X1 U903 ( .A(n1165), .B(KEYINPUT63), .ZN(n1226) );
AND2_X1 U904 ( .A1(n1036), .A2(n1170), .ZN(n1165) );
AND2_X1 U905 ( .A1(n1044), .A2(n1193), .ZN(n1036) );
XOR2_X1 U906 ( .A(G125), .B(n1227), .Z(G27) );
NOR2_X1 U907 ( .A1(n1202), .A2(n1200), .ZN(n1227) );
NAND3_X1 U908 ( .A1(n1192), .A2(n1066), .A3(n1057), .ZN(n1200) );
NOR3_X1 U909 ( .A1(n1203), .A2(n1067), .A3(n1052), .ZN(n1057) );
INV_X1 U910 ( .A(n1196), .ZN(n1202) );
NAND2_X1 U911 ( .A1(n1051), .A2(n1228), .ZN(n1196) );
NAND4_X1 U912 ( .A1(G902), .A2(G953), .A3(n1229), .A4(n1090), .ZN(n1228) );
INV_X1 U913 ( .A(G900), .ZN(n1090) );
XOR2_X1 U914 ( .A(n1230), .B(n1166), .Z(G24) );
NAND4_X1 U915 ( .A1(n1231), .A2(n1040), .A3(n1206), .A4(n1207), .ZN(n1166) );
NOR2_X1 U916 ( .A1(n1074), .A2(n1076), .ZN(n1040) );
INV_X1 U917 ( .A(n1232), .ZN(n1076) );
XNOR2_X1 U918 ( .A(G119), .B(n1167), .ZN(G21) );
NAND2_X1 U919 ( .A1(n1231), .A2(n1214), .ZN(n1167) );
AND3_X1 U920 ( .A1(n1221), .A2(n1220), .A3(n1044), .ZN(n1214) );
XNOR2_X1 U921 ( .A(n1168), .B(n1233), .ZN(G18) );
NOR2_X1 U922 ( .A1(KEYINPUT37), .A2(n1234), .ZN(n1233) );
INV_X1 U923 ( .A(G116), .ZN(n1234) );
NAND3_X1 U924 ( .A1(n1193), .A2(n1171), .A3(n1231), .ZN(n1168) );
INV_X1 U925 ( .A(n1038), .ZN(n1171) );
NAND2_X1 U926 ( .A1(n1069), .A2(n1207), .ZN(n1038) );
XOR2_X1 U927 ( .A(n1235), .B(KEYINPUT59), .Z(n1207) );
XOR2_X1 U928 ( .A(n1236), .B(n1169), .Z(G15) );
NAND3_X1 U929 ( .A1(n1041), .A2(n1193), .A3(n1231), .ZN(n1169) );
NOR3_X1 U930 ( .A1(n1237), .A2(n1067), .A3(n1052), .ZN(n1231) );
INV_X1 U931 ( .A(n1054), .ZN(n1067) );
AND2_X1 U932 ( .A1(n1232), .A2(n1220), .ZN(n1193) );
XNOR2_X1 U933 ( .A(n1238), .B(KEYINPUT42), .ZN(n1220) );
INV_X1 U934 ( .A(n1203), .ZN(n1041) );
NAND2_X1 U935 ( .A1(n1235), .A2(n1206), .ZN(n1203) );
XNOR2_X1 U936 ( .A(n1069), .B(KEYINPUT45), .ZN(n1206) );
NAND2_X1 U937 ( .A1(n1239), .A2(n1240), .ZN(G12) );
NAND2_X1 U938 ( .A1(G110), .A2(n1163), .ZN(n1240) );
XOR2_X1 U939 ( .A(n1241), .B(KEYINPUT10), .Z(n1239) );
OR2_X1 U940 ( .A1(n1163), .A2(G110), .ZN(n1241) );
NAND3_X1 U941 ( .A1(n1044), .A2(n1170), .A3(n1192), .ZN(n1163) );
INV_X1 U942 ( .A(n1042), .ZN(n1192) );
NAND2_X1 U943 ( .A1(n1221), .A2(n1238), .ZN(n1042) );
INV_X1 U944 ( .A(n1074), .ZN(n1238) );
XNOR2_X1 U945 ( .A(n1242), .B(G472), .ZN(n1074) );
NAND2_X1 U946 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XOR2_X1 U947 ( .A(n1245), .B(n1246), .Z(n1243) );
XOR2_X1 U948 ( .A(n1137), .B(n1131), .Z(n1246) );
XNOR2_X1 U949 ( .A(n1247), .B(n1248), .ZN(n1131) );
XOR2_X1 U950 ( .A(n1249), .B(n1159), .Z(n1248) );
INV_X1 U951 ( .A(n1250), .ZN(n1159) );
NOR2_X1 U952 ( .A1(KEYINPUT15), .A2(G116), .ZN(n1249) );
XOR2_X1 U953 ( .A(n1236), .B(G119), .Z(n1247) );
INV_X1 U954 ( .A(G113), .ZN(n1236) );
NAND3_X1 U955 ( .A1(n1251), .A2(n1059), .A3(G210), .ZN(n1137) );
XOR2_X1 U956 ( .A(n1252), .B(n1253), .Z(n1245) );
NOR2_X1 U957 ( .A1(KEYINPUT14), .A2(G101), .ZN(n1253) );
NAND2_X1 U958 ( .A1(KEYINPUT60), .A2(n1132), .ZN(n1252) );
XOR2_X1 U959 ( .A(n1232), .B(KEYINPUT29), .Z(n1221) );
XOR2_X1 U960 ( .A(n1254), .B(n1117), .Z(n1232) );
AND2_X1 U961 ( .A1(G217), .A2(n1255), .ZN(n1117) );
NAND2_X1 U962 ( .A1(n1115), .A2(n1244), .ZN(n1254) );
XNOR2_X1 U963 ( .A(n1256), .B(n1257), .ZN(n1115) );
XOR2_X1 U964 ( .A(G110), .B(n1258), .Z(n1257) );
XOR2_X1 U965 ( .A(G137), .B(G119), .Z(n1258) );
XOR2_X1 U966 ( .A(n1259), .B(n1094), .Z(n1256) );
XOR2_X1 U967 ( .A(n1260), .B(n1261), .Z(n1259) );
NAND2_X1 U968 ( .A1(G221), .A2(n1262), .ZN(n1260) );
NOR2_X1 U969 ( .A1(n1237), .A2(n1050), .ZN(n1170) );
NAND2_X1 U970 ( .A1(n1263), .A2(n1052), .ZN(n1050) );
XOR2_X1 U971 ( .A(n1073), .B(KEYINPUT54), .Z(n1052) );
XNOR2_X1 U972 ( .A(n1264), .B(G469), .ZN(n1073) );
NAND2_X1 U973 ( .A1(n1265), .A2(n1244), .ZN(n1264) );
XOR2_X1 U974 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U975 ( .A(n1093), .B(n1142), .Z(n1267) );
XNOR2_X1 U976 ( .A(G143), .B(n1261), .ZN(n1093) );
XOR2_X1 U977 ( .A(G128), .B(G146), .Z(n1261) );
XOR2_X1 U978 ( .A(n1268), .B(n1150), .Z(n1266) );
AND2_X1 U979 ( .A1(n1269), .A2(n1270), .ZN(n1150) );
NAND3_X1 U980 ( .A1(n1271), .A2(G227), .A3(n1272), .ZN(n1270) );
XOR2_X1 U981 ( .A(n1210), .B(G110), .Z(n1272) );
NAND2_X1 U982 ( .A1(n1273), .A2(n1274), .ZN(n1269) );
NAND2_X1 U983 ( .A1(n1271), .A2(G227), .ZN(n1274) );
XOR2_X1 U984 ( .A(KEYINPUT5), .B(n1059), .Z(n1271) );
XOR2_X1 U985 ( .A(G140), .B(G110), .Z(n1273) );
NAND2_X1 U986 ( .A1(KEYINPUT36), .A2(n1132), .ZN(n1268) );
XOR2_X1 U987 ( .A(n1275), .B(n1096), .Z(n1132) );
XOR2_X1 U988 ( .A(G131), .B(G134), .Z(n1096) );
XOR2_X1 U989 ( .A(n1097), .B(KEYINPUT57), .Z(n1275) );
INV_X1 U990 ( .A(G137), .ZN(n1097) );
XOR2_X1 U991 ( .A(n1054), .B(KEYINPUT19), .Z(n1263) );
NAND2_X1 U992 ( .A1(G221), .A2(n1255), .ZN(n1054) );
NAND2_X1 U993 ( .A1(G234), .A2(n1244), .ZN(n1255) );
NAND2_X1 U994 ( .A1(n1066), .A2(n1276), .ZN(n1237) );
NAND2_X1 U995 ( .A1(n1277), .A2(n1051), .ZN(n1276) );
NAND3_X1 U996 ( .A1(n1229), .A2(n1059), .A3(G952), .ZN(n1051) );
NAND3_X1 U997 ( .A1(n1104), .A2(n1229), .A3(G902), .ZN(n1277) );
NAND2_X1 U998 ( .A1(G237), .A2(G234), .ZN(n1229) );
NOR2_X1 U999 ( .A1(G898), .A2(n1059), .ZN(n1104) );
NOR2_X1 U1000 ( .A1(n1065), .A2(n1064), .ZN(n1066) );
AND2_X1 U1001 ( .A1(G214), .A2(n1278), .ZN(n1064) );
NAND2_X1 U1002 ( .A1(n1244), .A2(n1251), .ZN(n1278) );
INV_X1 U1003 ( .A(n1218), .ZN(n1065) );
NAND2_X1 U1004 ( .A1(n1279), .A2(n1280), .ZN(n1218) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1281), .ZN(n1280) );
NAND2_X1 U1006 ( .A1(n1244), .A2(n1282), .ZN(n1281) );
OR2_X1 U1007 ( .A1(n1251), .A2(n1283), .ZN(n1282) );
NAND3_X1 U1008 ( .A1(n1284), .A2(n1244), .A3(n1283), .ZN(n1279) );
XOR2_X1 U1009 ( .A(n1285), .B(n1156), .Z(n1283) );
XOR2_X1 U1010 ( .A(n1111), .B(n1286), .Z(n1156) );
AND2_X1 U1011 ( .A1(n1059), .A2(G224), .ZN(n1286) );
XNOR2_X1 U1012 ( .A(n1287), .B(n1288), .ZN(n1111) );
XOR2_X1 U1013 ( .A(G110), .B(n1289), .Z(n1288) );
XOR2_X1 U1014 ( .A(G122), .B(G113), .Z(n1289) );
XOR2_X1 U1015 ( .A(n1290), .B(n1142), .Z(n1287) );
XNOR2_X1 U1016 ( .A(n1291), .B(n1292), .ZN(n1142) );
XOR2_X1 U1017 ( .A(KEYINPUT44), .B(G107), .Z(n1292) );
XOR2_X1 U1018 ( .A(G104), .B(n1225), .Z(n1291) );
INV_X1 U1019 ( .A(G101), .ZN(n1225) );
NAND2_X1 U1020 ( .A1(n1293), .A2(KEYINPUT30), .ZN(n1290) );
XOR2_X1 U1021 ( .A(n1294), .B(G116), .Z(n1293) );
NAND2_X1 U1022 ( .A1(KEYINPUT2), .A2(n1295), .ZN(n1294) );
XOR2_X1 U1023 ( .A(KEYINPUT16), .B(G119), .Z(n1295) );
NAND2_X1 U1024 ( .A1(n1296), .A2(KEYINPUT35), .ZN(n1285) );
XOR2_X1 U1025 ( .A(n1250), .B(n1297), .Z(n1296) );
NOR2_X1 U1026 ( .A1(G125), .A2(KEYINPUT33), .ZN(n1297) );
XOR2_X1 U1027 ( .A(n1298), .B(G128), .Z(n1250) );
NAND2_X1 U1028 ( .A1(KEYINPUT3), .A2(n1299), .ZN(n1298) );
XOR2_X1 U1029 ( .A(G146), .B(G143), .Z(n1299) );
NAND2_X1 U1030 ( .A1(G237), .A2(G210), .ZN(n1284) );
INV_X1 U1031 ( .A(n1045), .ZN(n1044) );
NAND2_X1 U1032 ( .A1(n1069), .A2(n1235), .ZN(n1045) );
NOR2_X1 U1033 ( .A1(n1300), .A2(n1077), .ZN(n1235) );
NOR3_X1 U1034 ( .A1(G478), .A2(G902), .A3(n1301), .ZN(n1077) );
AND2_X1 U1035 ( .A1(n1302), .A2(n1078), .ZN(n1300) );
NAND2_X1 U1036 ( .A1(n1120), .A2(n1244), .ZN(n1078) );
INV_X1 U1037 ( .A(n1301), .ZN(n1120) );
XOR2_X1 U1038 ( .A(n1303), .B(n1304), .Z(n1301) );
XOR2_X1 U1039 ( .A(G107), .B(n1305), .Z(n1304) );
XOR2_X1 U1040 ( .A(G143), .B(G128), .Z(n1305) );
XOR2_X1 U1041 ( .A(n1306), .B(n1307), .Z(n1303) );
XOR2_X1 U1042 ( .A(n1308), .B(n1309), .Z(n1307) );
NAND2_X1 U1043 ( .A1(KEYINPUT39), .A2(n1310), .ZN(n1309) );
INV_X1 U1044 ( .A(G134), .ZN(n1310) );
NAND2_X1 U1045 ( .A1(n1311), .A2(n1312), .ZN(n1308) );
NAND2_X1 U1046 ( .A1(G116), .A2(n1230), .ZN(n1312) );
XOR2_X1 U1047 ( .A(KEYINPUT7), .B(n1313), .Z(n1311) );
NOR2_X1 U1048 ( .A1(G116), .A2(n1230), .ZN(n1313) );
INV_X1 U1049 ( .A(G122), .ZN(n1230) );
NAND2_X1 U1050 ( .A1(G217), .A2(n1262), .ZN(n1306) );
AND2_X1 U1051 ( .A1(G234), .A2(n1059), .ZN(n1262) );
XNOR2_X1 U1052 ( .A(G478), .B(KEYINPUT46), .ZN(n1302) );
XOR2_X1 U1053 ( .A(n1314), .B(G475), .Z(n1069) );
NAND2_X1 U1054 ( .A1(n1315), .A2(n1244), .ZN(n1314) );
INV_X1 U1055 ( .A(G902), .ZN(n1244) );
XOR2_X1 U1056 ( .A(n1125), .B(KEYINPUT28), .Z(n1315) );
XOR2_X1 U1057 ( .A(n1316), .B(n1317), .Z(n1125) );
XOR2_X1 U1058 ( .A(G113), .B(G104), .Z(n1317) );
XNOR2_X1 U1059 ( .A(n1318), .B(n1319), .ZN(n1316) );
NOR2_X1 U1060 ( .A1(KEYINPUT24), .A2(n1320), .ZN(n1319) );
XOR2_X1 U1061 ( .A(KEYINPUT17), .B(G122), .Z(n1320) );
NOR2_X1 U1062 ( .A1(KEYINPUT23), .A2(n1321), .ZN(n1318) );
XOR2_X1 U1063 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U1064 ( .A(n1324), .B(n1325), .Z(n1323) );
NOR2_X1 U1065 ( .A1(KEYINPUT4), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1066 ( .A(n1327), .B(n1328), .Z(n1326) );
AND3_X1 U1067 ( .A1(G214), .A2(n1059), .A3(n1251), .ZN(n1328) );
INV_X1 U1068 ( .A(G237), .ZN(n1251) );
INV_X1 U1069 ( .A(G953), .ZN(n1059) );
XNOR2_X1 U1070 ( .A(G131), .B(G143), .ZN(n1327) );
INV_X1 U1071 ( .A(G146), .ZN(n1324) );
NAND2_X1 U1072 ( .A1(KEYINPUT18), .A2(n1094), .ZN(n1322) );
XNOR2_X1 U1073 ( .A(G125), .B(n1210), .ZN(n1094) );
INV_X1 U1074 ( .A(G140), .ZN(n1210) );
endmodule


