//Key = 0111100011010000100111000001001011000000010110011101000010001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372;

XOR2_X1 U749 ( .A(G107), .B(n1036), .Z(G9) );
NOR2_X1 U750 ( .A1(KEYINPUT53), .A2(n1037), .ZN(n1036) );
NOR2_X1 U751 ( .A1(n1038), .A2(n1039), .ZN(G75) );
NOR3_X1 U752 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
INV_X1 U753 ( .A(G952), .ZN(n1041) );
NAND3_X1 U754 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1040) );
NAND2_X1 U755 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U756 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND3_X1 U757 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
NAND2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NAND2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
OR2_X1 U760 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(n1053) );
NAND2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U764 ( .A1(n1059), .A2(n1065), .A3(n1055), .ZN(n1048) );
NAND2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U766 ( .A1(n1052), .A2(n1068), .ZN(n1067) );
NAND2_X1 U767 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U768 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U769 ( .A1(n1050), .A2(n1073), .ZN(n1066) );
NAND2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
INV_X1 U772 ( .A(n1078), .ZN(n1046) );
NOR3_X1 U773 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1038) );
NOR2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
INV_X1 U775 ( .A(KEYINPUT47), .ZN(n1083) );
NOR2_X1 U776 ( .A1(G953), .A2(G952), .ZN(n1082) );
NOR2_X1 U777 ( .A1(KEYINPUT47), .A2(n1084), .ZN(n1080) );
INV_X1 U778 ( .A(n1043), .ZN(n1079) );
NAND4_X1 U779 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1043) );
NOR4_X1 U780 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1088) );
XNOR2_X1 U781 ( .A(n1093), .B(n1094), .ZN(n1092) );
XNOR2_X1 U782 ( .A(G478), .B(n1095), .ZN(n1091) );
XNOR2_X1 U783 ( .A(G472), .B(n1096), .ZN(n1090) );
XOR2_X1 U784 ( .A(n1097), .B(n1098), .Z(n1089) );
XOR2_X1 U785 ( .A(n1099), .B(KEYINPUT36), .Z(n1098) );
NOR2_X1 U786 ( .A1(n1063), .A2(n1076), .ZN(n1087) );
INV_X1 U787 ( .A(n1100), .ZN(n1076) );
XNOR2_X1 U788 ( .A(n1101), .B(n1102), .ZN(n1086) );
NOR2_X1 U789 ( .A1(KEYINPUT62), .A2(n1103), .ZN(n1102) );
XNOR2_X1 U790 ( .A(KEYINPUT35), .B(n1104), .ZN(n1103) );
INV_X1 U791 ( .A(n1072), .ZN(n1085) );
XOR2_X1 U792 ( .A(n1105), .B(n1106), .Z(G72) );
XOR2_X1 U793 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U794 ( .A1(G953), .A2(n1109), .ZN(n1108) );
NOR2_X1 U795 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XNOR2_X1 U796 ( .A(n1112), .B(KEYINPUT22), .ZN(n1110) );
NAND2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1107) );
NAND2_X1 U798 ( .A1(G953), .A2(n1115), .ZN(n1114) );
XOR2_X1 U799 ( .A(n1116), .B(n1117), .Z(n1113) );
XNOR2_X1 U800 ( .A(n1118), .B(n1119), .ZN(n1117) );
XOR2_X1 U801 ( .A(n1120), .B(n1121), .Z(n1116) );
XOR2_X1 U802 ( .A(KEYINPUT50), .B(G125), .Z(n1121) );
NAND2_X1 U803 ( .A1(KEYINPUT30), .A2(n1122), .ZN(n1120) );
NAND2_X1 U804 ( .A1(n1123), .A2(n1124), .ZN(n1105) );
NAND2_X1 U805 ( .A1(G900), .A2(G227), .ZN(n1124) );
XNOR2_X1 U806 ( .A(G953), .B(KEYINPUT44), .ZN(n1123) );
NAND2_X1 U807 ( .A1(n1125), .A2(n1126), .ZN(G69) );
NAND3_X1 U808 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1126) );
XNOR2_X1 U809 ( .A(n1130), .B(n1131), .ZN(n1129) );
NAND2_X1 U810 ( .A1(G953), .A2(n1132), .ZN(n1127) );
NAND2_X1 U811 ( .A1(n1133), .A2(n1134), .ZN(n1125) );
NAND2_X1 U812 ( .A1(n1135), .A2(n1128), .ZN(n1134) );
INV_X1 U813 ( .A(KEYINPUT18), .ZN(n1128) );
NAND2_X1 U814 ( .A1(G953), .A2(n1136), .ZN(n1135) );
NAND2_X1 U815 ( .A1(G898), .A2(G224), .ZN(n1136) );
XOR2_X1 U816 ( .A(n1131), .B(n1130), .Z(n1133) );
AND2_X1 U817 ( .A1(n1137), .A2(n1044), .ZN(n1130) );
NAND3_X1 U818 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1137) );
XNOR2_X1 U819 ( .A(KEYINPUT19), .B(n1037), .ZN(n1139) );
NAND2_X1 U820 ( .A1(n1141), .A2(n1142), .ZN(n1131) );
NAND2_X1 U821 ( .A1(G953), .A2(n1143), .ZN(n1142) );
XNOR2_X1 U822 ( .A(n1144), .B(n1145), .ZN(n1141) );
NAND2_X1 U823 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
NAND2_X1 U824 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND2_X1 U825 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
OR2_X1 U826 ( .A1(n1152), .A2(KEYINPUT32), .ZN(n1151) );
NAND3_X1 U827 ( .A1(n1153), .A2(n1154), .A3(KEYINPUT32), .ZN(n1146) );
NAND2_X1 U828 ( .A1(KEYINPUT21), .A2(n1155), .ZN(n1154) );
NAND2_X1 U829 ( .A1(n1156), .A2(n1150), .ZN(n1155) );
INV_X1 U830 ( .A(n1148), .ZN(n1156) );
NAND2_X1 U831 ( .A1(n1150), .A2(n1152), .ZN(n1153) );
INV_X1 U832 ( .A(KEYINPUT21), .ZN(n1152) );
NOR2_X1 U833 ( .A1(n1084), .A2(n1157), .ZN(G66) );
XNOR2_X1 U834 ( .A(n1158), .B(n1159), .ZN(n1157) );
NOR2_X1 U835 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR3_X1 U836 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(G63) );
NOR3_X1 U837 ( .A1(n1165), .A2(G953), .A3(G952), .ZN(n1164) );
AND2_X1 U838 ( .A1(n1165), .A2(n1084), .ZN(n1163) );
INV_X1 U839 ( .A(KEYINPUT26), .ZN(n1165) );
NOR3_X1 U840 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1162) );
NOR3_X1 U841 ( .A1(n1169), .A2(n1170), .A3(n1161), .ZN(n1168) );
NOR2_X1 U842 ( .A1(n1171), .A2(n1172), .ZN(n1167) );
NOR2_X1 U843 ( .A1(n1173), .A2(n1170), .ZN(n1171) );
NOR2_X1 U844 ( .A1(n1084), .A2(n1174), .ZN(G60) );
NOR3_X1 U845 ( .A1(n1094), .A2(n1175), .A3(n1176), .ZN(n1174) );
NOR4_X1 U846 ( .A1(n1177), .A2(n1161), .A3(KEYINPUT0), .A4(n1093), .ZN(n1176) );
NOR2_X1 U847 ( .A1(n1178), .A2(n1179), .ZN(n1175) );
NOR3_X1 U848 ( .A1(n1093), .A2(KEYINPUT0), .A3(n1173), .ZN(n1179) );
INV_X1 U849 ( .A(n1042), .ZN(n1173) );
INV_X1 U850 ( .A(G475), .ZN(n1093) );
XNOR2_X1 U851 ( .A(G104), .B(n1180), .ZN(G6) );
NOR2_X1 U852 ( .A1(n1084), .A2(n1181), .ZN(G57) );
XOR2_X1 U853 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U854 ( .A(n1184), .B(n1185), .Z(n1183) );
XNOR2_X1 U855 ( .A(n1186), .B(n1187), .ZN(n1182) );
NOR3_X1 U856 ( .A1(n1161), .A2(KEYINPUT29), .A3(n1188), .ZN(n1187) );
INV_X1 U857 ( .A(G472), .ZN(n1188) );
NOR2_X1 U858 ( .A1(n1084), .A2(n1189), .ZN(G54) );
XOR2_X1 U859 ( .A(n1190), .B(n1191), .Z(n1189) );
XNOR2_X1 U860 ( .A(n1192), .B(n1193), .ZN(n1191) );
NOR2_X1 U861 ( .A1(KEYINPUT58), .A2(n1194), .ZN(n1192) );
XNOR2_X1 U862 ( .A(G110), .B(G140), .ZN(n1194) );
XOR2_X1 U863 ( .A(n1195), .B(n1196), .Z(n1190) );
NOR2_X1 U864 ( .A1(n1101), .A2(n1161), .ZN(n1196) );
NAND2_X1 U865 ( .A1(n1197), .A2(n1198), .ZN(n1195) );
NAND2_X1 U866 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U867 ( .A(KEYINPUT55), .B(n1201), .Z(n1200) );
NOR2_X1 U868 ( .A1(n1084), .A2(n1202), .ZN(G51) );
XOR2_X1 U869 ( .A(n1203), .B(n1204), .Z(n1202) );
XNOR2_X1 U870 ( .A(n1205), .B(n1206), .ZN(n1204) );
XNOR2_X1 U871 ( .A(n1207), .B(n1208), .ZN(n1203) );
XOR2_X1 U872 ( .A(KEYINPUT59), .B(n1209), .Z(n1208) );
NOR2_X1 U873 ( .A1(n1097), .A2(n1161), .ZN(n1209) );
NAND2_X1 U874 ( .A1(G902), .A2(n1042), .ZN(n1161) );
NAND4_X1 U875 ( .A1(n1140), .A2(n1138), .A3(n1210), .A4(n1112), .ZN(n1042) );
AND4_X1 U876 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1112) );
NOR2_X1 U877 ( .A1(n1215), .A2(n1111), .ZN(n1210) );
NAND4_X1 U878 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1111) );
NAND3_X1 U879 ( .A1(n1220), .A2(n1058), .A3(n1221), .ZN(n1217) );
XNOR2_X1 U880 ( .A(n1052), .B(KEYINPUT41), .ZN(n1221) );
NAND2_X1 U881 ( .A1(n1052), .A2(n1222), .ZN(n1216) );
XOR2_X1 U882 ( .A(KEYINPUT52), .B(n1223), .Z(n1222) );
INV_X1 U883 ( .A(n1037), .ZN(n1215) );
NAND3_X1 U884 ( .A1(n1058), .A2(n1050), .A3(n1224), .ZN(n1037) );
AND3_X1 U885 ( .A1(n1225), .A2(n1226), .A3(n1227), .ZN(n1138) );
NAND2_X1 U886 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND2_X1 U887 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND4_X1 U888 ( .A1(n1232), .A2(n1233), .A3(n1050), .A4(n1234), .ZN(n1231) );
NOR2_X1 U889 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XNOR2_X1 U890 ( .A(n1237), .B(KEYINPUT23), .ZN(n1230) );
AND3_X1 U891 ( .A1(n1180), .A2(n1238), .A3(n1239), .ZN(n1140) );
NAND3_X1 U892 ( .A1(n1059), .A2(n1224), .A3(n1240), .ZN(n1239) );
NAND3_X1 U893 ( .A1(n1050), .A2(n1057), .A3(n1224), .ZN(n1180) );
NOR2_X1 U894 ( .A1(n1044), .A2(G952), .ZN(n1084) );
XNOR2_X1 U895 ( .A(G146), .B(n1211), .ZN(G48) );
NAND3_X1 U896 ( .A1(n1228), .A2(n1057), .A3(n1241), .ZN(n1211) );
XNOR2_X1 U897 ( .A(n1212), .B(n1242), .ZN(G45) );
XNOR2_X1 U898 ( .A(KEYINPUT7), .B(n1243), .ZN(n1242) );
NAND2_X1 U899 ( .A1(n1220), .A2(n1244), .ZN(n1212) );
NAND2_X1 U900 ( .A1(n1245), .A2(n1246), .ZN(G42) );
NAND2_X1 U901 ( .A1(n1247), .A2(n1122), .ZN(n1246) );
NAND2_X1 U902 ( .A1(G140), .A2(n1248), .ZN(n1245) );
NAND2_X1 U903 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
NAND2_X1 U904 ( .A1(KEYINPUT13), .A2(n1251), .ZN(n1250) );
INV_X1 U905 ( .A(n1213), .ZN(n1251) );
OR2_X1 U906 ( .A1(n1247), .A2(KEYINPUT13), .ZN(n1249) );
NOR2_X1 U907 ( .A1(KEYINPUT34), .A2(n1213), .ZN(n1247) );
NAND3_X1 U908 ( .A1(n1052), .A2(n1252), .A3(n1253), .ZN(n1213) );
XNOR2_X1 U909 ( .A(G137), .B(n1214), .ZN(G39) );
NAND3_X1 U910 ( .A1(n1052), .A2(n1059), .A3(n1241), .ZN(n1214) );
XOR2_X1 U911 ( .A(G134), .B(n1254), .Z(G36) );
AND3_X1 U912 ( .A1(n1220), .A2(n1058), .A3(n1052), .ZN(n1254) );
XNOR2_X1 U913 ( .A(G131), .B(n1255), .ZN(G33) );
NAND2_X1 U914 ( .A1(n1223), .A2(n1052), .ZN(n1255) );
AND2_X1 U915 ( .A1(n1256), .A2(n1100), .ZN(n1052) );
XNOR2_X1 U916 ( .A(n1077), .B(KEYINPUT27), .ZN(n1256) );
XNOR2_X1 U917 ( .A(n1257), .B(KEYINPUT12), .ZN(n1077) );
AND2_X1 U918 ( .A1(n1220), .A2(n1057), .ZN(n1223) );
AND3_X1 U919 ( .A1(n1252), .A2(n1258), .A3(n1240), .ZN(n1220) );
XNOR2_X1 U920 ( .A(G128), .B(n1218), .ZN(G30) );
NAND3_X1 U921 ( .A1(n1228), .A2(n1058), .A3(n1241), .ZN(n1218) );
AND4_X1 U922 ( .A1(n1259), .A2(n1252), .A3(n1072), .A4(n1258), .ZN(n1241) );
XNOR2_X1 U923 ( .A(G101), .B(n1260), .ZN(G3) );
NAND3_X1 U924 ( .A1(n1224), .A2(n1261), .A3(n1240), .ZN(n1260) );
XOR2_X1 U925 ( .A(KEYINPUT45), .B(n1059), .Z(n1261) );
NAND2_X1 U926 ( .A1(n1262), .A2(n1263), .ZN(G27) );
NAND2_X1 U927 ( .A1(G125), .A2(n1219), .ZN(n1263) );
XOR2_X1 U928 ( .A(n1264), .B(KEYINPUT39), .Z(n1262) );
OR2_X1 U929 ( .A1(n1219), .A2(G125), .ZN(n1264) );
NAND3_X1 U930 ( .A1(n1228), .A2(n1055), .A3(n1253), .ZN(n1219) );
AND4_X1 U931 ( .A1(n1057), .A2(n1071), .A3(n1072), .A4(n1258), .ZN(n1253) );
NAND2_X1 U932 ( .A1(n1078), .A2(n1265), .ZN(n1258) );
NAND4_X1 U933 ( .A1(G953), .A2(G902), .A3(n1266), .A4(n1115), .ZN(n1265) );
INV_X1 U934 ( .A(G900), .ZN(n1115) );
XNOR2_X1 U935 ( .A(G122), .B(n1267), .ZN(G24) );
NAND4_X1 U936 ( .A1(n1244), .A2(n1050), .A3(n1268), .A4(n1233), .ZN(n1267) );
XNOR2_X1 U937 ( .A(KEYINPUT31), .B(n1235), .ZN(n1268) );
NOR2_X1 U938 ( .A1(n1072), .A2(n1259), .ZN(n1050) );
NOR3_X1 U939 ( .A1(n1269), .A2(n1236), .A3(n1074), .ZN(n1244) );
XNOR2_X1 U940 ( .A(G119), .B(n1270), .ZN(G21) );
NAND2_X1 U941 ( .A1(n1237), .A2(n1228), .ZN(n1270) );
AND3_X1 U942 ( .A1(n1259), .A2(n1055), .A3(n1271), .ZN(n1237) );
AND3_X1 U943 ( .A1(n1059), .A2(n1233), .A3(n1072), .ZN(n1271) );
INV_X1 U944 ( .A(n1235), .ZN(n1055) );
INV_X1 U945 ( .A(n1071), .ZN(n1259) );
XOR2_X1 U946 ( .A(n1225), .B(n1272), .Z(G18) );
NAND2_X1 U947 ( .A1(KEYINPUT11), .A2(G116), .ZN(n1272) );
NAND3_X1 U948 ( .A1(n1273), .A2(n1058), .A3(n1228), .ZN(n1225) );
INV_X1 U949 ( .A(n1074), .ZN(n1228) );
XOR2_X1 U950 ( .A(n1274), .B(KEYINPUT51), .Z(n1074) );
NOR2_X1 U951 ( .A1(n1269), .A2(n1275), .ZN(n1058) );
NAND2_X1 U952 ( .A1(n1276), .A2(n1277), .ZN(G15) );
NAND2_X1 U953 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
XOR2_X1 U954 ( .A(KEYINPUT43), .B(n1280), .Z(n1276) );
NOR2_X1 U955 ( .A1(n1278), .A2(n1279), .ZN(n1280) );
INV_X1 U956 ( .A(G113), .ZN(n1279) );
INV_X1 U957 ( .A(n1226), .ZN(n1278) );
NAND3_X1 U958 ( .A1(n1274), .A2(n1057), .A3(n1273), .ZN(n1226) );
NOR3_X1 U959 ( .A1(n1069), .A2(n1281), .A3(n1235), .ZN(n1273) );
NAND2_X1 U960 ( .A1(n1282), .A2(n1064), .ZN(n1235) );
XNOR2_X1 U961 ( .A(KEYINPUT60), .B(n1283), .ZN(n1282) );
INV_X1 U962 ( .A(n1240), .ZN(n1069) );
NOR2_X1 U963 ( .A1(n1071), .A2(n1072), .ZN(n1240) );
NAND2_X1 U964 ( .A1(n1284), .A2(n1285), .ZN(n1057) );
OR3_X1 U965 ( .A1(n1232), .A2(n1236), .A3(KEYINPUT6), .ZN(n1285) );
NAND2_X1 U966 ( .A1(KEYINPUT6), .A2(n1059), .ZN(n1284) );
INV_X1 U967 ( .A(n1286), .ZN(n1274) );
XNOR2_X1 U968 ( .A(G110), .B(n1238), .ZN(G12) );
NAND4_X1 U969 ( .A1(n1059), .A2(n1224), .A3(n1071), .A4(n1072), .ZN(n1238) );
XOR2_X1 U970 ( .A(n1287), .B(n1160), .Z(n1072) );
NAND2_X1 U971 ( .A1(G217), .A2(n1288), .ZN(n1160) );
NAND2_X1 U972 ( .A1(n1158), .A2(n1289), .ZN(n1287) );
XNOR2_X1 U973 ( .A(n1290), .B(n1291), .ZN(n1158) );
XOR2_X1 U974 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U975 ( .A(n1294), .B(G110), .Z(n1293) );
NAND2_X1 U976 ( .A1(n1295), .A2(G221), .ZN(n1294) );
XNOR2_X1 U977 ( .A(G137), .B(KEYINPUT48), .ZN(n1292) );
XNOR2_X1 U978 ( .A(n1296), .B(n1297), .ZN(n1290) );
XOR2_X1 U979 ( .A(n1298), .B(n1299), .Z(n1297) );
NOR2_X1 U980 ( .A1(G119), .A2(KEYINPUT42), .ZN(n1298) );
XNOR2_X1 U981 ( .A(n1096), .B(n1300), .ZN(n1071) );
NOR2_X1 U982 ( .A1(G472), .A2(KEYINPUT24), .ZN(n1300) );
NAND2_X1 U983 ( .A1(n1301), .A2(n1289), .ZN(n1096) );
XNOR2_X1 U984 ( .A(n1302), .B(n1303), .ZN(n1301) );
INV_X1 U985 ( .A(n1186), .ZN(n1303) );
XNOR2_X1 U986 ( .A(n1304), .B(G101), .ZN(n1186) );
NAND2_X1 U987 ( .A1(n1305), .A2(G210), .ZN(n1304) );
NOR2_X1 U988 ( .A1(KEYINPUT25), .A2(n1306), .ZN(n1302) );
XOR2_X1 U989 ( .A(n1307), .B(n1185), .Z(n1306) );
XNOR2_X1 U990 ( .A(n1308), .B(n1309), .ZN(n1185) );
XOR2_X1 U991 ( .A(KEYINPUT8), .B(KEYINPUT16), .Z(n1309) );
NOR2_X1 U992 ( .A1(KEYINPUT5), .A2(n1184), .ZN(n1307) );
XNOR2_X1 U993 ( .A(n1310), .B(n1311), .ZN(n1184) );
INV_X1 U994 ( .A(n1207), .ZN(n1311) );
NOR3_X1 U995 ( .A1(n1286), .A2(n1281), .A3(n1061), .ZN(n1224) );
INV_X1 U996 ( .A(n1252), .ZN(n1061) );
NOR2_X1 U997 ( .A1(n1064), .A2(n1312), .ZN(n1252) );
XNOR2_X1 U998 ( .A(KEYINPUT60), .B(n1063), .ZN(n1312) );
INV_X1 U999 ( .A(n1283), .ZN(n1063) );
NAND2_X1 U1000 ( .A1(G221), .A2(n1288), .ZN(n1283) );
NAND2_X1 U1001 ( .A1(G234), .A2(n1313), .ZN(n1288) );
XNOR2_X1 U1002 ( .A(KEYINPUT1), .B(n1289), .ZN(n1313) );
XOR2_X1 U1003 ( .A(n1314), .B(n1101), .Z(n1064) );
INV_X1 U1004 ( .A(G469), .ZN(n1101) );
NAND2_X1 U1005 ( .A1(KEYINPUT56), .A2(n1104), .ZN(n1314) );
NAND2_X1 U1006 ( .A1(n1315), .A2(n1289), .ZN(n1104) );
XOR2_X1 U1007 ( .A(n1316), .B(n1317), .Z(n1315) );
XOR2_X1 U1008 ( .A(n1318), .B(n1319), .Z(n1317) );
NOR2_X1 U1009 ( .A1(KEYINPUT10), .A2(n1193), .ZN(n1319) );
NAND2_X1 U1010 ( .A1(G227), .A2(n1044), .ZN(n1193) );
NOR2_X1 U1011 ( .A1(G110), .A2(KEYINPUT14), .ZN(n1318) );
XNOR2_X1 U1012 ( .A(n1320), .B(n1122), .ZN(n1316) );
INV_X1 U1013 ( .A(G140), .ZN(n1122) );
NAND2_X1 U1014 ( .A1(n1197), .A2(n1321), .ZN(n1320) );
NAND2_X1 U1015 ( .A1(n1199), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1016 ( .A(KEYINPUT57), .B(n1201), .Z(n1322) );
OR2_X1 U1017 ( .A1(n1201), .A2(n1199), .ZN(n1197) );
AND2_X1 U1018 ( .A1(n1323), .A2(n1324), .ZN(n1199) );
NAND2_X1 U1019 ( .A1(n1150), .A2(n1325), .ZN(n1324) );
INV_X1 U1020 ( .A(KEYINPUT38), .ZN(n1325) );
NAND3_X1 U1021 ( .A1(G101), .A2(n1326), .A3(KEYINPUT38), .ZN(n1323) );
XOR2_X1 U1022 ( .A(n1310), .B(n1327), .Z(n1201) );
INV_X1 U1023 ( .A(n1118), .ZN(n1327) );
XOR2_X1 U1024 ( .A(n1207), .B(KEYINPUT37), .Z(n1118) );
XNOR2_X1 U1025 ( .A(n1119), .B(KEYINPUT9), .ZN(n1310) );
XOR2_X1 U1026 ( .A(G131), .B(n1328), .Z(n1119) );
XOR2_X1 U1027 ( .A(G137), .B(G134), .Z(n1328) );
INV_X1 U1028 ( .A(n1233), .ZN(n1281) );
NAND2_X1 U1029 ( .A1(n1078), .A2(n1329), .ZN(n1233) );
NAND4_X1 U1030 ( .A1(G953), .A2(G902), .A3(n1266), .A4(n1143), .ZN(n1329) );
INV_X1 U1031 ( .A(G898), .ZN(n1143) );
NAND3_X1 U1032 ( .A1(n1266), .A2(n1044), .A3(G952), .ZN(n1078) );
NAND2_X1 U1033 ( .A1(G237), .A2(G234), .ZN(n1266) );
NAND2_X1 U1034 ( .A1(n1257), .A2(n1100), .ZN(n1286) );
NAND2_X1 U1035 ( .A1(G214), .A2(n1330), .ZN(n1100) );
XNOR2_X1 U1036 ( .A(n1331), .B(n1099), .ZN(n1257) );
NAND3_X1 U1037 ( .A1(n1332), .A2(n1333), .A3(n1289), .ZN(n1099) );
NAND2_X1 U1038 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
INV_X1 U1039 ( .A(n1206), .ZN(n1334) );
NAND2_X1 U1040 ( .A1(n1206), .A2(n1336), .ZN(n1332) );
NAND2_X1 U1041 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
NAND2_X1 U1042 ( .A1(KEYINPUT3), .A2(n1339), .ZN(n1338) );
INV_X1 U1043 ( .A(n1335), .ZN(n1339) );
NOR2_X1 U1044 ( .A1(KEYINPUT54), .A2(n1340), .ZN(n1335) );
OR2_X1 U1045 ( .A1(n1340), .A2(KEYINPUT3), .ZN(n1337) );
XOR2_X1 U1046 ( .A(n1205), .B(n1341), .Z(n1340) );
NOR2_X1 U1047 ( .A1(KEYINPUT46), .A2(n1207), .ZN(n1341) );
XOR2_X1 U1048 ( .A(G143), .B(n1299), .Z(n1207) );
XOR2_X1 U1049 ( .A(G128), .B(G146), .Z(n1299) );
XNOR2_X1 U1050 ( .A(G125), .B(n1342), .ZN(n1205) );
NOR2_X1 U1051 ( .A1(G953), .A2(n1132), .ZN(n1342) );
INV_X1 U1052 ( .A(G224), .ZN(n1132) );
XNOR2_X1 U1053 ( .A(n1343), .B(n1150), .ZN(n1206) );
XOR2_X1 U1054 ( .A(G101), .B(n1326), .Z(n1150) );
XNOR2_X1 U1055 ( .A(n1344), .B(G107), .ZN(n1326) );
INV_X1 U1056 ( .A(G104), .ZN(n1344) );
XNOR2_X1 U1057 ( .A(n1148), .B(n1145), .ZN(n1343) );
XOR2_X1 U1058 ( .A(G110), .B(n1345), .Z(n1145) );
NOR2_X1 U1059 ( .A1(KEYINPUT17), .A2(n1346), .ZN(n1345) );
XNOR2_X1 U1060 ( .A(n1308), .B(KEYINPUT2), .ZN(n1148) );
XNOR2_X1 U1061 ( .A(G113), .B(n1347), .ZN(n1308) );
XOR2_X1 U1062 ( .A(G119), .B(G116), .Z(n1347) );
NAND2_X1 U1063 ( .A1(KEYINPUT33), .A2(n1097), .ZN(n1331) );
NAND2_X1 U1064 ( .A1(G210), .A2(n1330), .ZN(n1097) );
NAND2_X1 U1065 ( .A1(n1348), .A2(n1289), .ZN(n1330) );
INV_X1 U1066 ( .A(G902), .ZN(n1289) );
INV_X1 U1067 ( .A(G237), .ZN(n1348) );
NOR2_X1 U1068 ( .A1(n1232), .A2(n1275), .ZN(n1059) );
INV_X1 U1069 ( .A(n1236), .ZN(n1275) );
XOR2_X1 U1070 ( .A(n1094), .B(n1349), .Z(n1236) );
NOR2_X1 U1071 ( .A1(G475), .A2(KEYINPUT63), .ZN(n1349) );
NOR2_X1 U1072 ( .A1(n1178), .A2(G902), .ZN(n1094) );
INV_X1 U1073 ( .A(n1177), .ZN(n1178) );
NAND2_X1 U1074 ( .A1(n1350), .A2(n1351), .ZN(n1177) );
NAND2_X1 U1075 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
XOR2_X1 U1076 ( .A(n1354), .B(KEYINPUT15), .Z(n1350) );
OR2_X1 U1077 ( .A1(n1353), .A2(n1352), .ZN(n1354) );
XNOR2_X1 U1078 ( .A(n1355), .B(n1356), .ZN(n1352) );
XNOR2_X1 U1079 ( .A(n1243), .B(n1357), .ZN(n1356) );
XOR2_X1 U1080 ( .A(KEYINPUT20), .B(G146), .Z(n1357) );
XOR2_X1 U1081 ( .A(n1358), .B(n1296), .Z(n1355) );
XOR2_X1 U1082 ( .A(G125), .B(G140), .Z(n1296) );
XOR2_X1 U1083 ( .A(n1359), .B(G131), .Z(n1358) );
NAND2_X1 U1084 ( .A1(n1305), .A2(G214), .ZN(n1359) );
NOR2_X1 U1085 ( .A1(G953), .A2(G237), .ZN(n1305) );
XNOR2_X1 U1086 ( .A(n1360), .B(n1346), .ZN(n1353) );
XNOR2_X1 U1087 ( .A(G104), .B(G113), .ZN(n1360) );
INV_X1 U1088 ( .A(n1269), .ZN(n1232) );
NAND2_X1 U1089 ( .A1(n1361), .A2(n1362), .ZN(n1269) );
NAND2_X1 U1090 ( .A1(n1363), .A2(n1170), .ZN(n1362) );
INV_X1 U1091 ( .A(G478), .ZN(n1170) );
XNOR2_X1 U1092 ( .A(KEYINPUT4), .B(n1095), .ZN(n1363) );
NAND2_X1 U1093 ( .A1(n1364), .A2(G478), .ZN(n1361) );
XNOR2_X1 U1094 ( .A(KEYINPUT40), .B(n1095), .ZN(n1364) );
INV_X1 U1095 ( .A(n1166), .ZN(n1095) );
NOR2_X1 U1096 ( .A1(n1172), .A2(G902), .ZN(n1166) );
INV_X1 U1097 ( .A(n1169), .ZN(n1172) );
XNOR2_X1 U1098 ( .A(n1365), .B(n1366), .ZN(n1169) );
XNOR2_X1 U1099 ( .A(n1346), .B(n1367), .ZN(n1366) );
XNOR2_X1 U1100 ( .A(n1368), .B(n1369), .ZN(n1367) );
NAND2_X1 U1101 ( .A1(KEYINPUT61), .A2(n1370), .ZN(n1369) );
XNOR2_X1 U1102 ( .A(n1243), .B(G128), .ZN(n1370) );
INV_X1 U1103 ( .A(G143), .ZN(n1243) );
NAND2_X1 U1104 ( .A1(KEYINPUT49), .A2(G107), .ZN(n1368) );
XOR2_X1 U1105 ( .A(G122), .B(KEYINPUT28), .Z(n1346) );
XOR2_X1 U1106 ( .A(n1371), .B(n1372), .Z(n1365) );
XOR2_X1 U1107 ( .A(G134), .B(G116), .Z(n1372) );
NAND2_X1 U1108 ( .A1(G217), .A2(n1295), .ZN(n1371) );
AND2_X1 U1109 ( .A1(G234), .A2(n1044), .ZN(n1295) );
INV_X1 U1110 ( .A(G953), .ZN(n1044) );
endmodule


