//Key = 1000011101000000010011010110001101110001010010100111011111010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356;

XNOR2_X1 U737 ( .A(n1034), .B(n1035), .ZN(G9) );
NAND4_X1 U738 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(G75) );
NAND4_X1 U739 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1038) );
NAND2_X1 U740 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NAND3_X1 U741 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
XOR2_X1 U742 ( .A(n1049), .B(G469), .Z(n1048) );
XOR2_X1 U743 ( .A(KEYINPUT22), .B(n1050), .Z(n1047) );
NAND3_X1 U744 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1044) );
NAND2_X1 U745 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NAND3_X1 U746 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1051) );
NAND4_X1 U747 ( .A1(n1059), .A2(n1060), .A3(n1053), .A4(n1061), .ZN(n1037) );
NOR2_X1 U748 ( .A1(n1055), .A2(n1054), .ZN(n1061) );
INV_X1 U749 ( .A(n1062), .ZN(n1053) );
NAND2_X1 U750 ( .A1(n1063), .A2(n1064), .ZN(n1060) );
NAND2_X1 U751 ( .A1(n1040), .A2(n1041), .ZN(n1064) );
NAND3_X1 U752 ( .A1(n1065), .A2(n1066), .A3(n1043), .ZN(n1059) );
NAND2_X1 U753 ( .A1(n1040), .A2(n1067), .ZN(n1066) );
NAND2_X1 U754 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U755 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U756 ( .A1(n1041), .A2(n1072), .ZN(n1065) );
NAND2_X1 U757 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U758 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
INV_X1 U759 ( .A(n1077), .ZN(n1073) );
XOR2_X1 U760 ( .A(n1078), .B(n1079), .Z(G72) );
NOR2_X1 U761 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XNOR2_X1 U762 ( .A(n1082), .B(KEYINPUT54), .ZN(n1081) );
XOR2_X1 U763 ( .A(n1083), .B(n1084), .Z(n1080) );
XOR2_X1 U764 ( .A(n1085), .B(n1086), .Z(n1084) );
XNOR2_X1 U765 ( .A(n1087), .B(G134), .ZN(n1086) );
NOR2_X1 U766 ( .A1(G125), .A2(KEYINPUT10), .ZN(n1085) );
XNOR2_X1 U767 ( .A(n1088), .B(n1089), .ZN(n1083) );
NAND2_X1 U768 ( .A1(n1090), .A2(n1091), .ZN(n1078) );
NAND2_X1 U769 ( .A1(n1092), .A2(n1039), .ZN(n1091) );
NAND2_X1 U770 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XNOR2_X1 U771 ( .A(KEYINPUT17), .B(n1095), .ZN(n1094) );
NAND3_X1 U772 ( .A1(KEYINPUT0), .A2(n1096), .A3(G953), .ZN(n1090) );
NAND2_X1 U773 ( .A1(G900), .A2(G227), .ZN(n1096) );
XOR2_X1 U774 ( .A(n1097), .B(n1098), .Z(G69) );
NOR2_X1 U775 ( .A1(n1099), .A2(G953), .ZN(n1098) );
NAND2_X1 U776 ( .A1(n1100), .A2(n1101), .ZN(n1097) );
NAND2_X1 U777 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND2_X1 U778 ( .A1(G953), .A2(n1104), .ZN(n1103) );
NAND2_X1 U779 ( .A1(G953), .A2(n1105), .ZN(n1100) );
NAND2_X1 U780 ( .A1(G898), .A2(n1106), .ZN(n1105) );
OR2_X1 U781 ( .A1(n1102), .A2(G224), .ZN(n1106) );
XOR2_X1 U782 ( .A(n1107), .B(n1108), .Z(n1102) );
XOR2_X1 U783 ( .A(KEYINPUT48), .B(n1109), .Z(n1108) );
XOR2_X1 U784 ( .A(n1110), .B(n1111), .Z(n1107) );
NOR2_X1 U785 ( .A1(KEYINPUT1), .A2(n1112), .ZN(n1111) );
NOR2_X1 U786 ( .A1(n1113), .A2(n1114), .ZN(G66) );
XOR2_X1 U787 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U788 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NOR2_X1 U789 ( .A1(n1113), .A2(n1119), .ZN(G63) );
NOR2_X1 U790 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U791 ( .A(n1122), .B(KEYINPUT44), .Z(n1121) );
NAND2_X1 U792 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U793 ( .A1(n1124), .A2(n1123), .ZN(n1120) );
AND2_X1 U794 ( .A1(n1125), .A2(G478), .ZN(n1123) );
NOR2_X1 U795 ( .A1(n1113), .A2(n1126), .ZN(G60) );
XOR2_X1 U796 ( .A(n1127), .B(n1128), .Z(n1126) );
AND2_X1 U797 ( .A1(G475), .A2(n1125), .ZN(n1127) );
XNOR2_X1 U798 ( .A(n1129), .B(n1130), .ZN(G6) );
NOR2_X1 U799 ( .A1(n1113), .A2(n1131), .ZN(G57) );
NOR2_X1 U800 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XOR2_X1 U801 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U802 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U803 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
XNOR2_X1 U804 ( .A(n1140), .B(n1141), .ZN(n1139) );
XNOR2_X1 U805 ( .A(KEYINPUT6), .B(KEYINPUT28), .ZN(n1141) );
XOR2_X1 U806 ( .A(n1142), .B(KEYINPUT43), .Z(n1138) );
NAND2_X1 U807 ( .A1(n1143), .A2(n1144), .ZN(n1136) );
XNOR2_X1 U808 ( .A(KEYINPUT32), .B(n1145), .ZN(n1144) );
INV_X1 U809 ( .A(n1140), .ZN(n1145) );
XOR2_X1 U810 ( .A(n1146), .B(n1147), .Z(n1140) );
AND2_X1 U811 ( .A1(G472), .A2(n1125), .ZN(n1147) );
XNOR2_X1 U812 ( .A(KEYINPUT43), .B(n1142), .ZN(n1143) );
NAND2_X1 U813 ( .A1(n1148), .A2(n1149), .ZN(n1134) );
NOR2_X1 U814 ( .A1(n1148), .A2(n1149), .ZN(n1132) );
INV_X1 U815 ( .A(KEYINPUT29), .ZN(n1149) );
NOR3_X1 U816 ( .A1(n1113), .A2(n1150), .A3(n1151), .ZN(G54) );
NOR2_X1 U817 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U818 ( .A(n1154), .B(n1155), .Z(n1152) );
OR2_X1 U819 ( .A1(n1156), .A2(KEYINPUT2), .ZN(n1154) );
NOR2_X1 U820 ( .A1(n1157), .A2(n1158), .ZN(n1150) );
XOR2_X1 U821 ( .A(n1159), .B(n1155), .Z(n1158) );
XOR2_X1 U822 ( .A(n1160), .B(n1161), .Z(n1155) );
XOR2_X1 U823 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U824 ( .A1(KEYINPUT3), .A2(n1164), .ZN(n1162) );
XOR2_X1 U825 ( .A(n1165), .B(n1166), .Z(n1160) );
AND2_X1 U826 ( .A1(G469), .A2(n1125), .ZN(n1166) );
NAND2_X1 U827 ( .A1(KEYINPUT59), .A2(n1088), .ZN(n1165) );
NAND2_X1 U828 ( .A1(n1156), .A2(n1167), .ZN(n1159) );
INV_X1 U829 ( .A(KEYINPUT2), .ZN(n1167) );
XOR2_X1 U830 ( .A(n1168), .B(n1169), .Z(n1156) );
NAND2_X1 U831 ( .A1(KEYINPUT20), .A2(n1087), .ZN(n1168) );
NOR2_X1 U832 ( .A1(n1113), .A2(n1170), .ZN(G51) );
XOR2_X1 U833 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U834 ( .A1(n1173), .A2(n1118), .ZN(n1172) );
INV_X1 U835 ( .A(n1125), .ZN(n1118) );
NOR2_X1 U836 ( .A1(n1174), .A2(n1036), .ZN(n1125) );
AND3_X1 U837 ( .A1(n1093), .A2(n1095), .A3(n1099), .ZN(n1036) );
AND2_X1 U838 ( .A1(n1175), .A2(n1176), .ZN(n1099) );
NOR4_X1 U839 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
NOR4_X1 U840 ( .A1(n1035), .A2(n1181), .A3(n1182), .A4(n1130), .ZN(n1175) );
AND3_X1 U841 ( .A1(n1183), .A2(n1041), .A3(n1184), .ZN(n1130) );
INV_X1 U842 ( .A(n1185), .ZN(n1182) );
INV_X1 U843 ( .A(n1186), .ZN(n1181) );
AND3_X1 U844 ( .A1(n1187), .A2(n1041), .A3(n1183), .ZN(n1035) );
AND4_X1 U845 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1093) );
AND3_X1 U846 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1191) );
NAND3_X1 U847 ( .A1(n1077), .A2(n1195), .A3(n1196), .ZN(n1190) );
NAND2_X1 U848 ( .A1(n1056), .A2(n1057), .ZN(n1195) );
INV_X1 U849 ( .A(n1187), .ZN(n1056) );
NAND4_X1 U850 ( .A1(n1197), .A2(n1077), .A3(n1198), .A4(n1199), .ZN(n1188) );
XNOR2_X1 U851 ( .A(KEYINPUT14), .B(n1068), .ZN(n1199) );
INV_X1 U852 ( .A(n1200), .ZN(n1068) );
NOR2_X1 U853 ( .A1(n1201), .A2(n1202), .ZN(n1171) );
XOR2_X1 U854 ( .A(KEYINPUT19), .B(n1203), .Z(n1202) );
AND2_X1 U855 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NOR2_X1 U856 ( .A1(n1205), .A2(n1204), .ZN(n1201) );
XNOR2_X1 U857 ( .A(n1206), .B(KEYINPUT26), .ZN(n1205) );
NOR2_X1 U858 ( .A1(n1039), .A2(G952), .ZN(n1113) );
XOR2_X1 U859 ( .A(n1207), .B(n1208), .Z(G48) );
XNOR2_X1 U860 ( .A(G146), .B(KEYINPUT52), .ZN(n1208) );
NAND3_X1 U861 ( .A1(n1184), .A2(n1077), .A3(n1196), .ZN(n1207) );
XNOR2_X1 U862 ( .A(G143), .B(n1209), .ZN(G45) );
NAND2_X1 U863 ( .A1(n1077), .A2(n1210), .ZN(n1209) );
XOR2_X1 U864 ( .A(KEYINPUT58), .B(n1211), .Z(n1210) );
AND2_X1 U865 ( .A1(n1198), .A2(n1212), .ZN(n1211) );
XNOR2_X1 U866 ( .A(G140), .B(n1189), .ZN(G42) );
NAND3_X1 U867 ( .A1(n1197), .A2(n1213), .A3(n1040), .ZN(n1189) );
NAND2_X1 U868 ( .A1(n1214), .A2(n1215), .ZN(G39) );
OR2_X1 U869 ( .A1(n1192), .A2(G137), .ZN(n1215) );
XOR2_X1 U870 ( .A(n1216), .B(KEYINPUT45), .Z(n1214) );
NAND2_X1 U871 ( .A1(G137), .A2(n1192), .ZN(n1216) );
NAND3_X1 U872 ( .A1(n1040), .A2(n1217), .A3(n1196), .ZN(n1192) );
XOR2_X1 U873 ( .A(n1194), .B(n1218), .Z(G36) );
NAND2_X1 U874 ( .A1(KEYINPUT51), .A2(G134), .ZN(n1218) );
NAND3_X1 U875 ( .A1(n1212), .A2(n1187), .A3(n1040), .ZN(n1194) );
NAND2_X1 U876 ( .A1(n1219), .A2(n1220), .ZN(G33) );
NAND2_X1 U877 ( .A1(G131), .A2(n1193), .ZN(n1220) );
XOR2_X1 U878 ( .A(n1221), .B(KEYINPUT4), .Z(n1219) );
OR2_X1 U879 ( .A1(n1193), .A2(G131), .ZN(n1221) );
NAND3_X1 U880 ( .A1(n1212), .A2(n1184), .A3(n1040), .ZN(n1193) );
NOR2_X1 U881 ( .A1(n1222), .A2(n1075), .ZN(n1040) );
AND2_X1 U882 ( .A1(n1197), .A2(n1200), .ZN(n1212) );
NAND3_X1 U883 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(G30) );
OR2_X1 U884 ( .A1(n1226), .A2(G128), .ZN(n1225) );
NAND2_X1 U885 ( .A1(KEYINPUT12), .A2(n1227), .ZN(n1224) );
NAND2_X1 U886 ( .A1(G128), .A2(n1228), .ZN(n1227) );
XNOR2_X1 U887 ( .A(KEYINPUT9), .B(n1226), .ZN(n1228) );
NAND2_X1 U888 ( .A1(n1229), .A2(n1230), .ZN(n1223) );
INV_X1 U889 ( .A(KEYINPUT12), .ZN(n1230) );
NAND2_X1 U890 ( .A1(n1231), .A2(n1232), .ZN(n1229) );
OR2_X1 U891 ( .A1(n1226), .A2(KEYINPUT9), .ZN(n1232) );
NAND3_X1 U892 ( .A1(G128), .A2(n1226), .A3(KEYINPUT9), .ZN(n1231) );
NAND3_X1 U893 ( .A1(n1196), .A2(n1187), .A3(n1233), .ZN(n1226) );
XNOR2_X1 U894 ( .A(n1077), .B(KEYINPUT35), .ZN(n1233) );
AND3_X1 U895 ( .A1(n1071), .A2(n1234), .A3(n1197), .ZN(n1196) );
NOR3_X1 U896 ( .A1(n1063), .A2(n1235), .A3(n1058), .ZN(n1197) );
XOR2_X1 U897 ( .A(n1180), .B(n1236), .Z(G3) );
NOR2_X1 U898 ( .A1(KEYINPUT18), .A2(n1237), .ZN(n1236) );
AND3_X1 U899 ( .A1(n1217), .A2(n1183), .A3(n1200), .ZN(n1180) );
XOR2_X1 U900 ( .A(n1095), .B(n1238), .Z(G27) );
NAND2_X1 U901 ( .A1(KEYINPUT57), .A2(G125), .ZN(n1238) );
NAND4_X1 U902 ( .A1(n1058), .A2(n1213), .A3(n1239), .A4(n1077), .ZN(n1095) );
NOR2_X1 U903 ( .A1(n1235), .A2(n1063), .ZN(n1239) );
INV_X1 U904 ( .A(n1043), .ZN(n1063) );
AND2_X1 U905 ( .A1(n1240), .A2(n1062), .ZN(n1235) );
NAND3_X1 U906 ( .A1(G902), .A2(n1241), .A3(n1082), .ZN(n1240) );
NOR2_X1 U907 ( .A1(n1039), .A2(G900), .ZN(n1082) );
AND3_X1 U908 ( .A1(n1070), .A2(n1071), .A3(n1184), .ZN(n1213) );
XOR2_X1 U909 ( .A(G122), .B(n1179), .Z(G24) );
AND3_X1 U910 ( .A1(n1041), .A2(n1198), .A3(n1242), .ZN(n1179) );
NAND2_X1 U911 ( .A1(n1243), .A2(n1244), .ZN(n1198) );
OR3_X1 U912 ( .A1(n1046), .A2(n1050), .A3(KEYINPUT37), .ZN(n1244) );
NAND2_X1 U913 ( .A1(KEYINPUT37), .A2(n1184), .ZN(n1243) );
NOR2_X1 U914 ( .A1(n1234), .A2(n1071), .ZN(n1041) );
XNOR2_X1 U915 ( .A(G119), .B(n1185), .ZN(G21) );
NAND4_X1 U916 ( .A1(n1242), .A2(n1217), .A3(n1071), .A4(n1234), .ZN(n1185) );
XOR2_X1 U917 ( .A(G116), .B(n1178), .Z(G18) );
AND3_X1 U918 ( .A1(n1242), .A2(n1187), .A3(n1200), .ZN(n1178) );
NOR2_X1 U919 ( .A1(n1245), .A2(n1050), .ZN(n1187) );
NAND2_X1 U920 ( .A1(n1246), .A2(n1247), .ZN(G15) );
NAND2_X1 U921 ( .A1(G113), .A2(n1186), .ZN(n1247) );
XOR2_X1 U922 ( .A(n1248), .B(KEYINPUT42), .Z(n1246) );
OR2_X1 U923 ( .A1(n1186), .A2(G113), .ZN(n1248) );
NAND3_X1 U924 ( .A1(n1200), .A2(n1242), .A3(n1184), .ZN(n1186) );
INV_X1 U925 ( .A(n1057), .ZN(n1184) );
NAND2_X1 U926 ( .A1(n1050), .A2(n1245), .ZN(n1057) );
AND3_X1 U927 ( .A1(n1249), .A2(n1043), .A3(n1058), .ZN(n1242) );
INV_X1 U928 ( .A(n1054), .ZN(n1058) );
NOR2_X1 U929 ( .A1(n1071), .A2(n1070), .ZN(n1200) );
NAND2_X1 U930 ( .A1(n1250), .A2(n1251), .ZN(G12) );
NAND2_X1 U931 ( .A1(n1177), .A2(n1169), .ZN(n1251) );
XOR2_X1 U932 ( .A(KEYINPUT61), .B(n1252), .Z(n1250) );
NOR2_X1 U933 ( .A1(n1177), .A2(n1169), .ZN(n1252) );
INV_X1 U934 ( .A(G110), .ZN(n1169) );
AND4_X1 U935 ( .A1(n1217), .A2(n1183), .A3(n1070), .A4(n1071), .ZN(n1177) );
XOR2_X1 U936 ( .A(n1253), .B(n1117), .Z(n1071) );
NAND2_X1 U937 ( .A1(G217), .A2(n1254), .ZN(n1117) );
OR2_X1 U938 ( .A1(n1115), .A2(G902), .ZN(n1253) );
NAND2_X1 U939 ( .A1(n1255), .A2(n1256), .ZN(n1115) );
NAND2_X1 U940 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND2_X1 U941 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
NAND2_X1 U942 ( .A1(KEYINPUT5), .A2(n1261), .ZN(n1260) );
INV_X1 U943 ( .A(KEYINPUT40), .ZN(n1259) );
NAND2_X1 U944 ( .A1(n1262), .A2(n1263), .ZN(n1255) );
NAND2_X1 U945 ( .A1(KEYINPUT5), .A2(n1264), .ZN(n1263) );
OR2_X1 U946 ( .A1(n1258), .A2(KEYINPUT40), .ZN(n1264) );
NAND2_X1 U947 ( .A1(n1265), .A2(n1266), .ZN(n1258) );
NAND3_X1 U948 ( .A1(G221), .A2(n1267), .A3(n1268), .ZN(n1266) );
XOR2_X1 U949 ( .A(KEYINPUT15), .B(G137), .Z(n1267) );
NAND2_X1 U950 ( .A1(n1269), .A2(n1270), .ZN(n1265) );
NAND2_X1 U951 ( .A1(n1268), .A2(G221), .ZN(n1270) );
XOR2_X1 U952 ( .A(KEYINPUT46), .B(G137), .Z(n1269) );
INV_X1 U953 ( .A(n1261), .ZN(n1262) );
XNOR2_X1 U954 ( .A(n1271), .B(n1272), .ZN(n1261) );
XOR2_X1 U955 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U956 ( .A(n1275), .B(G110), .ZN(n1274) );
XOR2_X1 U957 ( .A(KEYINPUT36), .B(KEYINPUT16), .Z(n1273) );
XOR2_X1 U958 ( .A(n1276), .B(n1277), .Z(n1271) );
XNOR2_X1 U959 ( .A(n1278), .B(n1279), .ZN(n1276) );
NAND2_X1 U960 ( .A1(KEYINPUT34), .A2(n1280), .ZN(n1279) );
NAND2_X1 U961 ( .A1(KEYINPUT21), .A2(G146), .ZN(n1278) );
INV_X1 U962 ( .A(n1234), .ZN(n1070) );
XNOR2_X1 U963 ( .A(n1281), .B(G472), .ZN(n1234) );
NAND2_X1 U964 ( .A1(n1282), .A2(n1174), .ZN(n1281) );
XOR2_X1 U965 ( .A(n1283), .B(n1148), .Z(n1282) );
XNOR2_X1 U966 ( .A(n1284), .B(G101), .ZN(n1148) );
NAND2_X1 U967 ( .A1(n1285), .A2(G210), .ZN(n1284) );
NOR2_X1 U968 ( .A1(KEYINPUT24), .A2(n1286), .ZN(n1283) );
XOR2_X1 U969 ( .A(n1142), .B(n1146), .Z(n1286) );
XNOR2_X1 U970 ( .A(n1164), .B(n1287), .ZN(n1146) );
XOR2_X1 U971 ( .A(n1288), .B(n1289), .Z(n1142) );
NOR2_X1 U972 ( .A1(G113), .A2(KEYINPUT11), .ZN(n1289) );
AND3_X1 U973 ( .A1(n1054), .A2(n1043), .A3(n1249), .ZN(n1183) );
AND2_X1 U974 ( .A1(n1077), .A2(n1290), .ZN(n1249) );
NAND2_X1 U975 ( .A1(n1062), .A2(n1291), .ZN(n1290) );
NAND4_X1 U976 ( .A1(G953), .A2(G902), .A3(n1241), .A4(n1292), .ZN(n1291) );
INV_X1 U977 ( .A(G898), .ZN(n1292) );
NAND3_X1 U978 ( .A1(n1241), .A2(n1039), .A3(G952), .ZN(n1062) );
NAND2_X1 U979 ( .A1(G237), .A2(G234), .ZN(n1241) );
NOR2_X1 U980 ( .A1(n1076), .A2(n1075), .ZN(n1077) );
AND2_X1 U981 ( .A1(G214), .A2(n1293), .ZN(n1075) );
INV_X1 U982 ( .A(n1222), .ZN(n1076) );
XOR2_X1 U983 ( .A(n1294), .B(n1173), .Z(n1222) );
NAND2_X1 U984 ( .A1(G210), .A2(n1293), .ZN(n1173) );
NAND2_X1 U985 ( .A1(n1174), .A2(n1295), .ZN(n1293) );
INV_X1 U986 ( .A(G237), .ZN(n1295) );
NAND2_X1 U987 ( .A1(n1296), .A2(n1174), .ZN(n1294) );
XNOR2_X1 U988 ( .A(n1204), .B(n1297), .ZN(n1296) );
XOR2_X1 U989 ( .A(n1206), .B(KEYINPUT63), .Z(n1297) );
XOR2_X1 U990 ( .A(n1110), .B(n1298), .Z(n1206) );
XOR2_X1 U991 ( .A(n1299), .B(n1112), .Z(n1298) );
XOR2_X1 U992 ( .A(G122), .B(G110), .Z(n1112) );
NOR2_X1 U993 ( .A1(n1109), .A2(KEYINPUT38), .ZN(n1299) );
AND2_X1 U994 ( .A1(n1300), .A2(n1301), .ZN(n1109) );
NAND2_X1 U995 ( .A1(G101), .A2(n1302), .ZN(n1301) );
XOR2_X1 U996 ( .A(KEYINPUT53), .B(n1303), .Z(n1300) );
NOR2_X1 U997 ( .A1(G101), .A2(n1302), .ZN(n1303) );
XNOR2_X1 U998 ( .A(n1129), .B(G107), .ZN(n1302) );
XOR2_X1 U999 ( .A(n1304), .B(n1305), .Z(n1110) );
XOR2_X1 U1000 ( .A(KEYINPUT23), .B(G113), .Z(n1305) );
NAND2_X1 U1001 ( .A1(n1306), .A2(n1307), .ZN(n1304) );
NAND2_X1 U1002 ( .A1(KEYINPUT25), .A2(n1288), .ZN(n1307) );
XNOR2_X1 U1003 ( .A(G119), .B(n1308), .ZN(n1288) );
NAND3_X1 U1004 ( .A1(n1308), .A2(n1280), .A3(n1309), .ZN(n1306) );
INV_X1 U1005 ( .A(KEYINPUT25), .ZN(n1309) );
INV_X1 U1006 ( .A(G119), .ZN(n1280) );
XOR2_X1 U1007 ( .A(G116), .B(KEYINPUT8), .Z(n1308) );
XOR2_X1 U1008 ( .A(n1310), .B(n1287), .Z(n1204) );
XNOR2_X1 U1009 ( .A(G125), .B(n1311), .ZN(n1310) );
NOR2_X1 U1010 ( .A1(G953), .A2(n1104), .ZN(n1311) );
INV_X1 U1011 ( .A(G224), .ZN(n1104) );
NAND2_X1 U1012 ( .A1(G221), .A2(n1254), .ZN(n1043) );
NAND2_X1 U1013 ( .A1(G234), .A2(n1174), .ZN(n1254) );
XNOR2_X1 U1014 ( .A(n1049), .B(n1312), .ZN(n1054) );
XOR2_X1 U1015 ( .A(KEYINPUT39), .B(n1313), .Z(n1312) );
NOR2_X1 U1016 ( .A1(KEYINPUT60), .A2(G469), .ZN(n1313) );
NAND2_X1 U1017 ( .A1(n1314), .A2(n1174), .ZN(n1049) );
INV_X1 U1018 ( .A(G902), .ZN(n1174) );
XOR2_X1 U1019 ( .A(n1164), .B(n1315), .Z(n1314) );
XNOR2_X1 U1020 ( .A(n1316), .B(n1317), .ZN(n1315) );
NOR2_X1 U1021 ( .A1(KEYINPUT27), .A2(n1318), .ZN(n1317) );
XNOR2_X1 U1022 ( .A(n1157), .B(n1319), .ZN(n1318) );
XNOR2_X1 U1023 ( .A(n1087), .B(G110), .ZN(n1319) );
INV_X1 U1024 ( .A(n1153), .ZN(n1157) );
NAND2_X1 U1025 ( .A1(G227), .A2(n1039), .ZN(n1153) );
NAND2_X1 U1026 ( .A1(KEYINPUT41), .A2(n1320), .ZN(n1316) );
XNOR2_X1 U1027 ( .A(n1287), .B(n1163), .ZN(n1320) );
XOR2_X1 U1028 ( .A(n1321), .B(n1237), .Z(n1163) );
INV_X1 U1029 ( .A(G101), .ZN(n1237) );
NAND3_X1 U1030 ( .A1(n1322), .A2(n1323), .A3(n1324), .ZN(n1321) );
NAND2_X1 U1031 ( .A1(KEYINPUT47), .A2(G107), .ZN(n1324) );
NAND3_X1 U1032 ( .A1(n1034), .A2(n1325), .A3(G104), .ZN(n1323) );
NAND2_X1 U1033 ( .A1(n1326), .A2(n1129), .ZN(n1322) );
INV_X1 U1034 ( .A(G104), .ZN(n1129) );
NAND2_X1 U1035 ( .A1(n1327), .A2(n1325), .ZN(n1326) );
INV_X1 U1036 ( .A(KEYINPUT47), .ZN(n1325) );
XNOR2_X1 U1037 ( .A(KEYINPUT31), .B(n1034), .ZN(n1327) );
INV_X1 U1038 ( .A(n1088), .ZN(n1287) );
XOR2_X1 U1039 ( .A(G128), .B(n1328), .Z(n1088) );
XOR2_X1 U1040 ( .A(n1089), .B(n1329), .Z(n1164) );
NOR2_X1 U1041 ( .A1(KEYINPUT13), .A2(n1330), .ZN(n1329) );
XNOR2_X1 U1042 ( .A(G134), .B(KEYINPUT50), .ZN(n1330) );
XOR2_X1 U1043 ( .A(G131), .B(G137), .Z(n1089) );
INV_X1 U1044 ( .A(n1055), .ZN(n1217) );
NAND2_X1 U1045 ( .A1(n1046), .A2(n1050), .ZN(n1055) );
XNOR2_X1 U1046 ( .A(n1331), .B(n1332), .ZN(n1050) );
NOR2_X1 U1047 ( .A1(G902), .A2(n1333), .ZN(n1332) );
XOR2_X1 U1048 ( .A(KEYINPUT62), .B(n1124), .Z(n1333) );
AND2_X1 U1049 ( .A1(n1334), .A2(n1335), .ZN(n1124) );
NAND2_X1 U1050 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
NAND2_X1 U1051 ( .A1(G217), .A2(n1268), .ZN(n1337) );
INV_X1 U1052 ( .A(n1338), .ZN(n1268) );
XOR2_X1 U1053 ( .A(KEYINPUT33), .B(n1339), .Z(n1334) );
NOR3_X1 U1054 ( .A1(n1340), .A2(n1336), .A3(n1338), .ZN(n1339) );
NAND2_X1 U1055 ( .A1(G234), .A2(n1039), .ZN(n1338) );
INV_X1 U1056 ( .A(G953), .ZN(n1039) );
XOR2_X1 U1057 ( .A(n1341), .B(n1342), .Z(n1336) );
XOR2_X1 U1058 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1059 ( .A(n1345), .B(n1034), .ZN(n1344) );
INV_X1 U1060 ( .A(G107), .ZN(n1034) );
NAND2_X1 U1061 ( .A1(KEYINPUT30), .A2(G143), .ZN(n1345) );
NAND2_X1 U1062 ( .A1(KEYINPUT56), .A2(n1346), .ZN(n1343) );
INV_X1 U1063 ( .A(G134), .ZN(n1346) );
XNOR2_X1 U1064 ( .A(G116), .B(n1347), .ZN(n1341) );
XNOR2_X1 U1065 ( .A(n1275), .B(G122), .ZN(n1347) );
INV_X1 U1066 ( .A(G128), .ZN(n1275) );
INV_X1 U1067 ( .A(G217), .ZN(n1340) );
XNOR2_X1 U1068 ( .A(G478), .B(KEYINPUT49), .ZN(n1331) );
INV_X1 U1069 ( .A(n1245), .ZN(n1046) );
XNOR2_X1 U1070 ( .A(n1348), .B(G475), .ZN(n1245) );
OR2_X1 U1071 ( .A1(n1128), .A2(G902), .ZN(n1348) );
XNOR2_X1 U1072 ( .A(n1349), .B(n1350), .ZN(n1128) );
XOR2_X1 U1073 ( .A(n1351), .B(n1352), .Z(n1350) );
XOR2_X1 U1074 ( .A(n1277), .B(n1328), .Z(n1352) );
XOR2_X1 U1075 ( .A(G143), .B(G146), .Z(n1328) );
XNOR2_X1 U1076 ( .A(G125), .B(n1087), .ZN(n1277) );
INV_X1 U1077 ( .A(G140), .ZN(n1087) );
XOR2_X1 U1078 ( .A(n1353), .B(n1354), .Z(n1351) );
NAND2_X1 U1079 ( .A1(KEYINPUT7), .A2(G113), .ZN(n1354) );
NAND2_X1 U1080 ( .A1(n1285), .A2(G214), .ZN(n1353) );
NOR2_X1 U1081 ( .A1(G953), .A2(G237), .ZN(n1285) );
XOR2_X1 U1082 ( .A(n1355), .B(n1356), .Z(n1349) );
XOR2_X1 U1083 ( .A(KEYINPUT55), .B(G131), .Z(n1356) );
XNOR2_X1 U1084 ( .A(G104), .B(G122), .ZN(n1355) );
endmodule


