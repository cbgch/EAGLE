//Key = 0100111100110000100010000110001010111111001000111111010101111111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411;

XOR2_X1 U761 ( .A(G107), .B(n1066), .Z(G9) );
NOR2_X1 U762 ( .A1(n1067), .A2(n1068), .ZN(G75) );
NOR4_X1 U763 ( .A1(n1069), .A2(n1070), .A3(G953), .A4(n1071), .ZN(n1068) );
NOR2_X1 U764 ( .A1(KEYINPUT26), .A2(n1072), .ZN(n1070) );
AND2_X1 U765 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U766 ( .A1(n1075), .A2(n1076), .ZN(n1069) );
NAND2_X1 U767 ( .A1(n1074), .A2(n1077), .ZN(n1076) );
NAND3_X1 U768 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
NAND2_X1 U769 ( .A1(KEYINPUT26), .A2(n1073), .ZN(n1080) );
NAND2_X1 U770 ( .A1(n1081), .A2(n1082), .ZN(n1073) );
NAND3_X1 U771 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
NAND2_X1 U772 ( .A1(n1086), .A2(n1087), .ZN(n1081) );
NAND2_X1 U773 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U774 ( .A1(n1090), .A2(n1085), .A3(n1091), .ZN(n1089) );
XOR2_X1 U775 ( .A(n1092), .B(KEYINPUT31), .Z(n1091) );
NAND2_X1 U776 ( .A1(n1083), .A2(n1093), .ZN(n1088) );
NAND2_X1 U777 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND3_X1 U778 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
INV_X1 U779 ( .A(n1099), .ZN(n1098) );
NAND2_X1 U780 ( .A1(n1100), .A2(n1101), .ZN(n1094) );
NAND3_X1 U781 ( .A1(n1102), .A2(n1083), .A3(n1085), .ZN(n1079) );
NAND2_X1 U782 ( .A1(n1086), .A2(n1103), .ZN(n1078) );
NAND2_X1 U783 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U784 ( .A1(n1083), .A2(n1106), .ZN(n1105) );
NAND2_X1 U785 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U786 ( .A1(n1109), .A2(n1100), .ZN(n1108) );
NAND2_X1 U787 ( .A1(n1097), .A2(n1110), .ZN(n1107) );
NAND2_X1 U788 ( .A1(n1085), .A2(n1111), .ZN(n1104) );
AND2_X1 U789 ( .A1(n1100), .A2(n1097), .ZN(n1085) );
INV_X1 U790 ( .A(n1112), .ZN(n1074) );
NOR3_X1 U791 ( .A1(n1071), .A2(G953), .A3(G952), .ZN(n1067) );
AND4_X1 U792 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1071) );
NOR3_X1 U793 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1116) );
NOR2_X1 U794 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
INV_X1 U795 ( .A(n1122), .ZN(n1118) );
NAND3_X1 U796 ( .A1(n1099), .A2(n1123), .A3(n1124), .ZN(n1117) );
NOR3_X1 U797 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1115) );
XOR2_X1 U798 ( .A(n1128), .B(KEYINPUT59), .Z(n1127) );
XNOR2_X1 U799 ( .A(n1129), .B(n1130), .ZN(n1126) );
NOR2_X1 U800 ( .A1(G478), .A2(KEYINPUT13), .ZN(n1130) );
XOR2_X1 U801 ( .A(n1131), .B(n1132), .Z(G72) );
XOR2_X1 U802 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U803 ( .A1(G953), .A2(n1135), .ZN(n1134) );
NAND2_X1 U804 ( .A1(G900), .A2(G227), .ZN(n1135) );
NAND2_X1 U805 ( .A1(n1136), .A2(n1137), .ZN(n1133) );
NAND2_X1 U806 ( .A1(G953), .A2(n1138), .ZN(n1137) );
XOR2_X1 U807 ( .A(n1139), .B(n1140), .Z(n1136) );
XOR2_X1 U808 ( .A(n1141), .B(n1142), .Z(n1140) );
INV_X1 U809 ( .A(n1143), .ZN(n1142) );
XOR2_X1 U810 ( .A(n1144), .B(n1145), .Z(n1139) );
NAND2_X1 U811 ( .A1(KEYINPUT61), .A2(G125), .ZN(n1145) );
AND2_X1 U812 ( .A1(n1146), .A2(n1147), .ZN(n1131) );
NAND2_X1 U813 ( .A1(n1148), .A2(n1149), .ZN(G69) );
NAND2_X1 U814 ( .A1(n1150), .A2(n1147), .ZN(n1149) );
XNOR2_X1 U815 ( .A(n1151), .B(n1152), .ZN(n1150) );
NAND2_X1 U816 ( .A1(n1153), .A2(G953), .ZN(n1148) );
NAND2_X1 U817 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U818 ( .A1(n1152), .A2(n1156), .ZN(n1155) );
INV_X1 U819 ( .A(G224), .ZN(n1156) );
NAND2_X1 U820 ( .A1(G224), .A2(n1157), .ZN(n1154) );
NAND2_X1 U821 ( .A1(G898), .A2(n1152), .ZN(n1157) );
NAND2_X1 U822 ( .A1(n1158), .A2(n1159), .ZN(n1152) );
NAND2_X1 U823 ( .A1(G953), .A2(n1160), .ZN(n1159) );
XOR2_X1 U824 ( .A(n1161), .B(n1162), .Z(n1158) );
XNOR2_X1 U825 ( .A(n1163), .B(n1164), .ZN(n1162) );
XOR2_X1 U826 ( .A(G122), .B(G110), .Z(n1161) );
NOR2_X1 U827 ( .A1(n1165), .A2(n1166), .ZN(G66) );
XOR2_X1 U828 ( .A(KEYINPUT56), .B(n1167), .Z(n1166) );
XOR2_X1 U829 ( .A(n1168), .B(n1169), .Z(n1165) );
NAND2_X1 U830 ( .A1(n1170), .A2(G217), .ZN(n1168) );
NOR2_X1 U831 ( .A1(n1167), .A2(n1171), .ZN(G63) );
NOR3_X1 U832 ( .A1(n1129), .A2(n1172), .A3(n1173), .ZN(n1171) );
AND3_X1 U833 ( .A1(n1174), .A2(G478), .A3(n1170), .ZN(n1173) );
NOR2_X1 U834 ( .A1(n1175), .A2(n1174), .ZN(n1172) );
NOR2_X1 U835 ( .A1(n1075), .A2(n1176), .ZN(n1175) );
INV_X1 U836 ( .A(G478), .ZN(n1176) );
NOR2_X1 U837 ( .A1(n1167), .A2(n1177), .ZN(G60) );
NOR2_X1 U838 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XOR2_X1 U839 ( .A(n1180), .B(KEYINPUT37), .Z(n1179) );
NAND2_X1 U840 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NOR2_X1 U841 ( .A1(n1181), .A2(n1182), .ZN(n1178) );
AND2_X1 U842 ( .A1(n1170), .A2(G475), .ZN(n1181) );
XOR2_X1 U843 ( .A(n1183), .B(n1184), .Z(G6) );
XNOR2_X1 U844 ( .A(G104), .B(KEYINPUT21), .ZN(n1184) );
NAND3_X1 U845 ( .A1(n1185), .A2(n1097), .A3(n1102), .ZN(n1183) );
NOR2_X1 U846 ( .A1(n1167), .A2(n1186), .ZN(G57) );
XOR2_X1 U847 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND2_X1 U848 ( .A1(n1170), .A2(G472), .ZN(n1187) );
NOR2_X1 U849 ( .A1(n1189), .A2(n1190), .ZN(G54) );
XOR2_X1 U850 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U851 ( .A(n1193), .B(n1143), .Z(n1192) );
XOR2_X1 U852 ( .A(n1194), .B(n1195), .Z(n1191) );
XOR2_X1 U853 ( .A(n1196), .B(n1197), .Z(n1195) );
NOR2_X1 U854 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U855 ( .A(KEYINPUT44), .B(KEYINPUT14), .Z(n1199) );
NAND2_X1 U856 ( .A1(KEYINPUT47), .A2(n1144), .ZN(n1196) );
NAND2_X1 U857 ( .A1(n1170), .A2(G469), .ZN(n1194) );
XNOR2_X1 U858 ( .A(n1167), .B(KEYINPUT42), .ZN(n1189) );
NOR2_X1 U859 ( .A1(n1167), .A2(n1200), .ZN(G51) );
XOR2_X1 U860 ( .A(n1201), .B(n1202), .Z(n1200) );
NAND2_X1 U861 ( .A1(n1170), .A2(n1203), .ZN(n1201) );
NOR2_X1 U862 ( .A1(n1204), .A2(n1075), .ZN(n1170) );
NOR2_X1 U863 ( .A1(n1146), .A2(n1151), .ZN(n1075) );
NAND3_X1 U864 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1151) );
NOR3_X1 U865 ( .A1(n1208), .A2(n1209), .A3(n1066), .ZN(n1207) );
AND3_X1 U866 ( .A1(n1097), .A2(n1084), .A3(n1185), .ZN(n1066) );
INV_X1 U867 ( .A(n1210), .ZN(n1084) );
NOR2_X1 U868 ( .A1(n1211), .A2(n1212), .ZN(n1208) );
NOR2_X1 U869 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
NOR2_X1 U870 ( .A1(n1215), .A2(n1216), .ZN(n1213) );
NAND2_X1 U871 ( .A1(n1110), .A2(n1217), .ZN(n1206) );
NAND2_X1 U872 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NAND3_X1 U873 ( .A1(n1220), .A2(n1086), .A3(n1221), .ZN(n1219) );
NOR3_X1 U874 ( .A1(n1222), .A2(KEYINPUT34), .A3(n1223), .ZN(n1221) );
XNOR2_X1 U875 ( .A(KEYINPUT1), .B(n1224), .ZN(n1218) );
NAND2_X1 U876 ( .A1(n1185), .A2(n1225), .ZN(n1205) );
NAND3_X1 U877 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1225) );
NAND2_X1 U878 ( .A1(n1229), .A2(n1097), .ZN(n1228) );
XOR2_X1 U879 ( .A(n1230), .B(KEYINPUT53), .Z(n1229) );
NAND2_X1 U880 ( .A1(n1086), .A2(n1231), .ZN(n1227) );
NAND2_X1 U881 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NAND2_X1 U882 ( .A1(KEYINPUT34), .A2(n1109), .ZN(n1233) );
NAND2_X1 U883 ( .A1(KEYINPUT32), .A2(n1101), .ZN(n1232) );
NAND3_X1 U884 ( .A1(n1101), .A2(n1234), .A3(n1235), .ZN(n1226) );
INV_X1 U885 ( .A(KEYINPUT32), .ZN(n1234) );
NAND4_X1 U886 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1146) );
NOR3_X1 U887 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1239) );
NOR3_X1 U888 ( .A1(n1223), .A2(n1243), .A3(n1244), .ZN(n1242) );
NOR2_X1 U889 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NOR3_X1 U890 ( .A1(n1216), .A2(n1247), .A3(n1248), .ZN(n1246) );
XOR2_X1 U891 ( .A(n1222), .B(KEYINPUT52), .Z(n1248) );
XOR2_X1 U892 ( .A(n1249), .B(KEYINPUT41), .Z(n1247) );
NOR3_X1 U893 ( .A1(n1250), .A2(n1249), .A3(n1230), .ZN(n1245) );
INV_X1 U894 ( .A(n1251), .ZN(n1243) );
NOR2_X1 U895 ( .A1(n1252), .A2(n1253), .ZN(n1240) );
NOR2_X1 U896 ( .A1(n1254), .A2(n1214), .ZN(n1252) );
NOR2_X1 U897 ( .A1(n1235), .A2(n1255), .ZN(n1254) );
XNOR2_X1 U898 ( .A(KEYINPUT60), .B(n1250), .ZN(n1255) );
NOR2_X1 U899 ( .A1(n1147), .A2(G952), .ZN(n1167) );
XOR2_X1 U900 ( .A(G146), .B(n1256), .Z(G48) );
NOR4_X1 U901 ( .A1(KEYINPUT23), .A2(n1230), .A3(n1257), .A4(n1250), .ZN(n1256) );
XOR2_X1 U902 ( .A(n1258), .B(n1259), .Z(G45) );
OR3_X1 U903 ( .A1(n1257), .A2(n1222), .A3(n1216), .ZN(n1259) );
XOR2_X1 U904 ( .A(n1238), .B(n1260), .Z(G42) );
XOR2_X1 U905 ( .A(n1144), .B(KEYINPUT19), .Z(n1260) );
INV_X1 U906 ( .A(G140), .ZN(n1144) );
NAND3_X1 U907 ( .A1(n1101), .A2(n1102), .A3(n1261), .ZN(n1238) );
XOR2_X1 U908 ( .A(G137), .B(n1262), .Z(G39) );
AND2_X1 U909 ( .A1(n1261), .A2(n1263), .ZN(n1262) );
NAND3_X1 U910 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(G36) );
NAND3_X1 U911 ( .A1(n1261), .A2(n1267), .A3(n1214), .ZN(n1266) );
NAND2_X1 U912 ( .A1(KEYINPUT10), .A2(n1268), .ZN(n1267) );
OR2_X1 U913 ( .A1(G134), .A2(KEYINPUT29), .ZN(n1268) );
OR2_X1 U914 ( .A1(G134), .A2(KEYINPUT10), .ZN(n1265) );
NAND3_X1 U915 ( .A1(G134), .A2(n1269), .A3(KEYINPUT10), .ZN(n1264) );
OR3_X1 U916 ( .A1(n1253), .A2(KEYINPUT29), .A3(n1270), .ZN(n1269) );
XOR2_X1 U917 ( .A(n1236), .B(n1271), .Z(G33) );
NAND2_X1 U918 ( .A1(KEYINPUT25), .A2(G131), .ZN(n1271) );
NAND3_X1 U919 ( .A1(n1261), .A2(n1102), .A3(n1109), .ZN(n1236) );
INV_X1 U920 ( .A(n1253), .ZN(n1261) );
NAND3_X1 U921 ( .A1(n1111), .A2(n1251), .A3(n1100), .ZN(n1253) );
AND2_X1 U922 ( .A1(n1272), .A2(n1099), .ZN(n1100) );
XOR2_X1 U923 ( .A(n1096), .B(KEYINPUT9), .Z(n1272) );
XOR2_X1 U924 ( .A(n1273), .B(KEYINPUT4), .Z(n1096) );
NAND2_X1 U925 ( .A1(n1274), .A2(n1275), .ZN(G30) );
NAND2_X1 U926 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XOR2_X1 U927 ( .A(n1278), .B(KEYINPUT22), .Z(n1274) );
OR2_X1 U928 ( .A1(n1277), .A2(n1276), .ZN(n1278) );
XNOR2_X1 U929 ( .A(n1279), .B(KEYINPUT8), .ZN(n1276) );
INV_X1 U930 ( .A(n1241), .ZN(n1277) );
NOR3_X1 U931 ( .A1(n1257), .A2(n1210), .A3(n1250), .ZN(n1241) );
NAND3_X1 U932 ( .A1(n1110), .A2(n1251), .A3(n1111), .ZN(n1257) );
INV_X1 U933 ( .A(n1223), .ZN(n1111) );
XNOR2_X1 U934 ( .A(G101), .B(n1280), .ZN(G3) );
NAND2_X1 U935 ( .A1(n1281), .A2(n1109), .ZN(n1280) );
XOR2_X1 U936 ( .A(n1282), .B(n1283), .Z(G27) );
NOR2_X1 U937 ( .A1(n1284), .A2(KEYINPUT17), .ZN(n1283) );
INV_X1 U938 ( .A(n1237), .ZN(n1284) );
NAND3_X1 U939 ( .A1(n1101), .A2(n1102), .A3(n1285), .ZN(n1237) );
AND3_X1 U940 ( .A1(n1083), .A2(n1251), .A3(n1110), .ZN(n1285) );
NAND2_X1 U941 ( .A1(n1112), .A2(n1286), .ZN(n1251) );
NAND4_X1 U942 ( .A1(G953), .A2(G902), .A3(n1287), .A4(n1138), .ZN(n1286) );
INV_X1 U943 ( .A(G900), .ZN(n1138) );
XOR2_X1 U944 ( .A(n1288), .B(n1289), .Z(G24) );
NOR3_X1 U945 ( .A1(n1290), .A2(n1215), .A3(n1212), .ZN(n1289) );
INV_X1 U946 ( .A(n1097), .ZN(n1215) );
NOR2_X1 U947 ( .A1(n1291), .A2(n1292), .ZN(n1097) );
XNOR2_X1 U948 ( .A(KEYINPUT51), .B(n1216), .ZN(n1290) );
NAND2_X1 U949 ( .A1(n1293), .A2(n1294), .ZN(n1216) );
XNOR2_X1 U950 ( .A(n1295), .B(KEYINPUT35), .ZN(n1293) );
NAND2_X1 U951 ( .A1(KEYINPUT16), .A2(n1296), .ZN(n1288) );
XOR2_X1 U952 ( .A(G119), .B(n1297), .Z(G21) );
NOR2_X1 U953 ( .A1(n1249), .A2(n1224), .ZN(n1297) );
NAND3_X1 U954 ( .A1(n1083), .A2(n1298), .A3(n1263), .ZN(n1224) );
NOR2_X1 U955 ( .A1(n1235), .A2(n1250), .ZN(n1263) );
NAND2_X1 U956 ( .A1(n1292), .A2(n1291), .ZN(n1250) );
INV_X1 U957 ( .A(n1113), .ZN(n1292) );
INV_X1 U958 ( .A(n1086), .ZN(n1235) );
XOR2_X1 U959 ( .A(G116), .B(n1299), .Z(G18) );
NOR2_X1 U960 ( .A1(n1212), .A2(n1270), .ZN(n1299) );
INV_X1 U961 ( .A(n1214), .ZN(n1270) );
NOR2_X1 U962 ( .A1(n1222), .A2(n1210), .ZN(n1214) );
NAND2_X1 U963 ( .A1(n1300), .A2(n1295), .ZN(n1210) );
XOR2_X1 U964 ( .A(G113), .B(n1209), .Z(G15) );
NOR3_X1 U965 ( .A1(n1222), .A2(n1230), .A3(n1212), .ZN(n1209) );
NAND3_X1 U966 ( .A1(n1110), .A2(n1298), .A3(n1083), .ZN(n1212) );
NOR2_X1 U967 ( .A1(n1301), .A2(n1090), .ZN(n1083) );
INV_X1 U968 ( .A(n1124), .ZN(n1090) );
INV_X1 U969 ( .A(n1249), .ZN(n1110) );
INV_X1 U970 ( .A(n1102), .ZN(n1230) );
NOR2_X1 U971 ( .A1(n1295), .A2(n1300), .ZN(n1102) );
INV_X1 U972 ( .A(n1294), .ZN(n1300) );
INV_X1 U973 ( .A(n1109), .ZN(n1222) );
NOR2_X1 U974 ( .A1(n1291), .A2(n1113), .ZN(n1109) );
XNOR2_X1 U975 ( .A(G110), .B(n1302), .ZN(G12) );
NAND2_X1 U976 ( .A1(n1281), .A2(n1101), .ZN(n1302) );
AND2_X1 U977 ( .A1(n1113), .A2(n1291), .ZN(n1101) );
NAND2_X1 U978 ( .A1(n1122), .A2(n1128), .ZN(n1291) );
NAND3_X1 U979 ( .A1(n1303), .A2(n1304), .A3(G217), .ZN(n1128) );
NAND2_X1 U980 ( .A1(n1169), .A2(n1204), .ZN(n1303) );
NAND3_X1 U981 ( .A1(n1305), .A2(n1204), .A3(n1169), .ZN(n1122) );
XNOR2_X1 U982 ( .A(n1306), .B(n1307), .ZN(n1169) );
XOR2_X1 U983 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U984 ( .A(n1310), .B(G140), .Z(n1309) );
NAND3_X1 U985 ( .A1(G221), .A2(n1147), .A3(n1311), .ZN(n1308) );
XNOR2_X1 U986 ( .A(G234), .B(KEYINPUT11), .ZN(n1311) );
XOR2_X1 U987 ( .A(n1312), .B(n1313), .Z(n1306) );
XNOR2_X1 U988 ( .A(n1314), .B(n1315), .ZN(n1312) );
NAND2_X1 U989 ( .A1(KEYINPUT20), .A2(n1316), .ZN(n1315) );
NAND2_X1 U990 ( .A1(n1317), .A2(KEYINPUT57), .ZN(n1314) );
XOR2_X1 U991 ( .A(n1282), .B(KEYINPUT3), .Z(n1317) );
NAND2_X1 U992 ( .A1(G217), .A2(n1318), .ZN(n1305) );
INV_X1 U993 ( .A(n1319), .ZN(n1318) );
XOR2_X1 U994 ( .A(n1320), .B(G472), .Z(n1113) );
NAND2_X1 U995 ( .A1(n1321), .A2(n1204), .ZN(n1320) );
XOR2_X1 U996 ( .A(n1188), .B(KEYINPUT15), .Z(n1321) );
XOR2_X1 U997 ( .A(n1322), .B(n1323), .Z(n1188) );
XOR2_X1 U998 ( .A(n1324), .B(n1325), .Z(n1323) );
XNOR2_X1 U999 ( .A(n1326), .B(n1327), .ZN(n1325) );
XOR2_X1 U1000 ( .A(n1328), .B(n1329), .Z(n1322) );
XNOR2_X1 U1001 ( .A(G101), .B(n1330), .ZN(n1329) );
NAND3_X1 U1002 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(n1330) );
NAND2_X1 U1003 ( .A1(n1334), .A2(n1335), .ZN(n1332) );
OR3_X1 U1004 ( .A1(n1334), .A2(n1336), .A3(n1335), .ZN(n1331) );
AND2_X1 U1005 ( .A1(n1337), .A2(n1338), .ZN(n1334) );
XOR2_X1 U1006 ( .A(KEYINPUT27), .B(G116), .Z(n1338) );
XOR2_X1 U1007 ( .A(n1310), .B(KEYINPUT33), .Z(n1337) );
NAND2_X1 U1008 ( .A1(n1339), .A2(G210), .ZN(n1328) );
AND2_X1 U1009 ( .A1(n1086), .A2(n1185), .ZN(n1281) );
NOR3_X1 U1010 ( .A1(n1249), .A2(n1220), .A3(n1223), .ZN(n1185) );
NAND2_X1 U1011 ( .A1(n1301), .A2(n1124), .ZN(n1223) );
NAND2_X1 U1012 ( .A1(G221), .A2(n1304), .ZN(n1124) );
NAND2_X1 U1013 ( .A1(n1319), .A2(n1204), .ZN(n1304) );
INV_X1 U1014 ( .A(n1092), .ZN(n1301) );
XNOR2_X1 U1015 ( .A(n1125), .B(KEYINPUT43), .ZN(n1092) );
XNOR2_X1 U1016 ( .A(n1340), .B(G469), .ZN(n1125) );
NAND2_X1 U1017 ( .A1(n1341), .A2(n1204), .ZN(n1340) );
XOR2_X1 U1018 ( .A(n1342), .B(n1343), .Z(n1341) );
XOR2_X1 U1019 ( .A(n1193), .B(n1344), .Z(n1343) );
NOR2_X1 U1020 ( .A1(KEYINPUT54), .A2(n1143), .ZN(n1344) );
XOR2_X1 U1021 ( .A(n1345), .B(G128), .Z(n1143) );
NAND3_X1 U1022 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1345) );
NAND2_X1 U1023 ( .A1(G143), .A2(n1349), .ZN(n1348) );
OR3_X1 U1024 ( .A1(n1349), .A2(n1350), .A3(G146), .ZN(n1347) );
INV_X1 U1025 ( .A(KEYINPUT62), .ZN(n1349) );
NAND2_X1 U1026 ( .A1(G146), .A2(n1350), .ZN(n1346) );
NAND2_X1 U1027 ( .A1(KEYINPUT63), .A2(n1258), .ZN(n1350) );
XOR2_X1 U1028 ( .A(n1351), .B(n1352), .Z(n1193) );
XOR2_X1 U1029 ( .A(n1324), .B(n1353), .Z(n1352) );
XOR2_X1 U1030 ( .A(n1354), .B(n1141), .Z(n1324) );
XNOR2_X1 U1031 ( .A(n1355), .B(n1356), .ZN(n1141) );
XOR2_X1 U1032 ( .A(n1316), .B(G134), .Z(n1355) );
INV_X1 U1033 ( .A(G137), .ZN(n1316) );
XNOR2_X1 U1034 ( .A(KEYINPUT58), .B(KEYINPUT45), .ZN(n1354) );
XNOR2_X1 U1035 ( .A(G101), .B(G110), .ZN(n1351) );
XOR2_X1 U1036 ( .A(n1198), .B(G140), .Z(n1342) );
NAND2_X1 U1037 ( .A1(G227), .A2(n1357), .ZN(n1198) );
XOR2_X1 U1038 ( .A(KEYINPUT39), .B(G953), .Z(n1357) );
INV_X1 U1039 ( .A(n1298), .ZN(n1220) );
NAND2_X1 U1040 ( .A1(n1358), .A2(n1112), .ZN(n1298) );
NAND3_X1 U1041 ( .A1(n1287), .A2(n1147), .A3(G952), .ZN(n1112) );
NAND4_X1 U1042 ( .A1(G953), .A2(G902), .A3(n1287), .A4(n1160), .ZN(n1358) );
INV_X1 U1043 ( .A(G898), .ZN(n1160) );
NAND2_X1 U1044 ( .A1(G237), .A2(n1319), .ZN(n1287) );
XNOR2_X1 U1045 ( .A(G234), .B(KEYINPUT36), .ZN(n1319) );
NAND2_X1 U1046 ( .A1(n1273), .A2(n1099), .ZN(n1249) );
NAND2_X1 U1047 ( .A1(G214), .A2(n1359), .ZN(n1099) );
NAND3_X1 U1048 ( .A1(n1360), .A2(n1361), .A3(n1123), .ZN(n1273) );
NAND2_X1 U1049 ( .A1(n1120), .A2(n1121), .ZN(n1123) );
INV_X1 U1050 ( .A(n1362), .ZN(n1120) );
OR2_X1 U1051 ( .A1(n1203), .A2(KEYINPUT38), .ZN(n1361) );
NAND3_X1 U1052 ( .A1(n1203), .A2(n1362), .A3(KEYINPUT38), .ZN(n1360) );
NAND2_X1 U1053 ( .A1(n1202), .A2(n1204), .ZN(n1362) );
XOR2_X1 U1054 ( .A(n1363), .B(n1364), .Z(n1202) );
XNOR2_X1 U1055 ( .A(n1313), .B(n1365), .ZN(n1364) );
XNOR2_X1 U1056 ( .A(n1327), .B(n1366), .ZN(n1365) );
NOR2_X1 U1057 ( .A1(KEYINPUT0), .A2(n1164), .ZN(n1366) );
XNOR2_X1 U1058 ( .A(n1353), .B(n1367), .ZN(n1164) );
NOR2_X1 U1059 ( .A1(G101), .A2(KEYINPUT18), .ZN(n1367) );
XNOR2_X1 U1060 ( .A(G104), .B(n1368), .ZN(n1353) );
XNOR2_X1 U1061 ( .A(n1258), .B(KEYINPUT5), .ZN(n1327) );
XOR2_X1 U1062 ( .A(G110), .B(n1326), .Z(n1313) );
XNOR2_X1 U1063 ( .A(n1279), .B(G146), .ZN(n1326) );
INV_X1 U1064 ( .A(G128), .ZN(n1279) );
XOR2_X1 U1065 ( .A(n1369), .B(n1370), .Z(n1363) );
XOR2_X1 U1066 ( .A(n1163), .B(n1371), .Z(n1370) );
NAND2_X1 U1067 ( .A1(G224), .A2(n1147), .ZN(n1371) );
NAND3_X1 U1068 ( .A1(n1372), .A2(n1373), .A3(n1333), .ZN(n1163) );
NAND2_X1 U1069 ( .A1(n1336), .A2(n1335), .ZN(n1333) );
NOR2_X1 U1070 ( .A1(n1310), .A2(G116), .ZN(n1336) );
NAND2_X1 U1071 ( .A1(n1374), .A2(n1310), .ZN(n1373) );
INV_X1 U1072 ( .A(G119), .ZN(n1310) );
XOR2_X1 U1073 ( .A(G116), .B(n1375), .Z(n1374) );
NAND3_X1 U1074 ( .A1(G116), .A2(n1375), .A3(G119), .ZN(n1372) );
XOR2_X1 U1075 ( .A(n1282), .B(G122), .Z(n1369) );
INV_X1 U1076 ( .A(G125), .ZN(n1282) );
INV_X1 U1077 ( .A(n1121), .ZN(n1203) );
NAND2_X1 U1078 ( .A1(G210), .A2(n1359), .ZN(n1121) );
NAND2_X1 U1079 ( .A1(n1376), .A2(n1204), .ZN(n1359) );
INV_X1 U1080 ( .A(G902), .ZN(n1204) );
INV_X1 U1081 ( .A(G237), .ZN(n1376) );
NOR2_X1 U1082 ( .A1(n1295), .A2(n1294), .ZN(n1086) );
XOR2_X1 U1083 ( .A(n1114), .B(KEYINPUT46), .Z(n1294) );
XOR2_X1 U1084 ( .A(n1377), .B(G475), .Z(n1114) );
OR2_X1 U1085 ( .A1(n1182), .A2(G902), .ZN(n1377) );
XOR2_X1 U1086 ( .A(n1378), .B(n1379), .Z(n1182) );
XOR2_X1 U1087 ( .A(G125), .B(n1380), .Z(n1379) );
XOR2_X1 U1088 ( .A(G146), .B(G140), .Z(n1380) );
XOR2_X1 U1089 ( .A(n1381), .B(n1382), .Z(n1378) );
NOR3_X1 U1090 ( .A1(n1383), .A2(n1384), .A3(n1385), .ZN(n1382) );
NOR2_X1 U1091 ( .A1(KEYINPUT2), .A2(n1386), .ZN(n1385) );
NOR2_X1 U1092 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
AND2_X1 U1093 ( .A1(n1356), .A2(KEYINPUT12), .ZN(n1388) );
NOR3_X1 U1094 ( .A1(KEYINPUT12), .A2(n1356), .A3(n1389), .ZN(n1387) );
NOR2_X1 U1095 ( .A1(n1390), .A2(n1391), .ZN(n1384) );
INV_X1 U1096 ( .A(KEYINPUT2), .ZN(n1391) );
NOR2_X1 U1097 ( .A1(n1389), .A2(n1392), .ZN(n1390) );
XOR2_X1 U1098 ( .A(KEYINPUT12), .B(n1356), .Z(n1392) );
AND2_X1 U1099 ( .A1(n1356), .A2(n1389), .ZN(n1383) );
XNOR2_X1 U1100 ( .A(n1258), .B(n1393), .ZN(n1389) );
AND2_X1 U1101 ( .A1(G214), .A2(n1339), .ZN(n1393) );
AND2_X1 U1102 ( .A1(n1394), .A2(n1147), .ZN(n1339) );
XOR2_X1 U1103 ( .A(KEYINPUT30), .B(G237), .Z(n1394) );
INV_X1 U1104 ( .A(G143), .ZN(n1258) );
XOR2_X1 U1105 ( .A(G131), .B(KEYINPUT7), .Z(n1356) );
NAND2_X1 U1106 ( .A1(KEYINPUT49), .A2(n1395), .ZN(n1381) );
XOR2_X1 U1107 ( .A(G104), .B(n1396), .Z(n1395) );
NOR4_X1 U1108 ( .A1(n1397), .A2(n1398), .A3(KEYINPUT24), .A4(n1399), .ZN(n1396) );
NOR2_X1 U1109 ( .A1(KEYINPUT6), .A2(n1375), .ZN(n1399) );
INV_X1 U1110 ( .A(n1335), .ZN(n1375) );
NOR2_X1 U1111 ( .A1(G122), .A2(n1400), .ZN(n1398) );
NOR2_X1 U1112 ( .A1(n1401), .A2(n1402), .ZN(n1400) );
XOR2_X1 U1113 ( .A(n1335), .B(KEYINPUT28), .Z(n1401) );
NOR3_X1 U1114 ( .A1(n1296), .A2(n1335), .A3(n1402), .ZN(n1397) );
INV_X1 U1115 ( .A(KEYINPUT6), .ZN(n1402) );
XNOR2_X1 U1116 ( .A(G113), .B(KEYINPUT50), .ZN(n1335) );
INV_X1 U1117 ( .A(G122), .ZN(n1296) );
XOR2_X1 U1118 ( .A(n1129), .B(G478), .Z(n1295) );
NOR2_X1 U1119 ( .A1(n1174), .A2(G902), .ZN(n1129) );
XOR2_X1 U1120 ( .A(n1403), .B(n1404), .Z(n1174) );
XOR2_X1 U1121 ( .A(G134), .B(n1405), .Z(n1404) );
XOR2_X1 U1122 ( .A(KEYINPUT55), .B(G143), .Z(n1405) );
XOR2_X1 U1123 ( .A(n1406), .B(n1407), .Z(n1403) );
XOR2_X1 U1124 ( .A(G128), .B(n1408), .Z(n1407) );
AND3_X1 U1125 ( .A1(G217), .A2(n1147), .A3(G234), .ZN(n1408) );
INV_X1 U1126 ( .A(G953), .ZN(n1147) );
NAND2_X1 U1127 ( .A1(n1409), .A2(KEYINPUT48), .ZN(n1406) );
XOR2_X1 U1128 ( .A(n1410), .B(n1368), .Z(n1409) );
XOR2_X1 U1129 ( .A(G107), .B(KEYINPUT40), .Z(n1368) );
XOR2_X1 U1130 ( .A(n1411), .B(G122), .Z(n1410) );
INV_X1 U1131 ( .A(G116), .ZN(n1411) );
endmodule


