//Key = 0011110111111110101010110000110010111101110000001001011001101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344;

XNOR2_X1 U749 ( .A(n1027), .B(n1028), .ZN(G9) );
NAND2_X1 U750 ( .A1(KEYINPUT32), .A2(G107), .ZN(n1028) );
NOR2_X1 U751 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR3_X1 U752 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
XOR2_X1 U753 ( .A(n1034), .B(KEYINPUT52), .Z(n1031) );
NAND3_X1 U754 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NAND4_X1 U755 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1036) );
NAND2_X1 U756 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND3_X1 U757 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1042) );
INV_X1 U758 ( .A(KEYINPUT11), .ZN(n1045) );
NAND3_X1 U759 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1040) );
NAND2_X1 U760 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND2_X1 U761 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U762 ( .A1(n1046), .A2(n1054), .ZN(n1047) );
NAND2_X1 U763 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U764 ( .A1(KEYINPUT11), .A2(n1044), .ZN(n1056) );
NAND4_X1 U765 ( .A1(n1049), .A2(n1046), .A3(n1050), .A4(n1057), .ZN(n1035) );
NAND2_X1 U766 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U767 ( .A1(n1039), .A2(n1060), .ZN(n1059) );
NAND2_X1 U768 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
OR2_X1 U769 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U770 ( .A1(n1038), .A2(n1065), .ZN(n1058) );
NAND2_X1 U771 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND3_X1 U772 ( .A1(G214), .A2(n1068), .A3(n1069), .ZN(n1067) );
NOR3_X1 U773 ( .A1(n1033), .A2(G952), .A3(n1032), .ZN(n1029) );
AND4_X1 U774 ( .A1(n1070), .A2(n1063), .A3(n1039), .A4(n1071), .ZN(n1032) );
NOR4_X1 U775 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1071) );
XNOR2_X1 U776 ( .A(KEYINPUT55), .B(n1076), .ZN(n1075) );
XNOR2_X1 U777 ( .A(G472), .B(n1077), .ZN(n1074) );
NOR2_X1 U778 ( .A1(KEYINPUT54), .A2(n1078), .ZN(n1073) );
AND2_X1 U779 ( .A1(n1079), .A2(KEYINPUT54), .ZN(n1072) );
XOR2_X1 U780 ( .A(n1080), .B(n1081), .Z(G72) );
XOR2_X1 U781 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR3_X1 U782 ( .A1(n1084), .A2(KEYINPUT43), .A3(n1085), .ZN(n1083) );
NOR2_X1 U783 ( .A1(G900), .A2(n1086), .ZN(n1085) );
XOR2_X1 U784 ( .A(n1087), .B(n1088), .Z(n1084) );
XOR2_X1 U785 ( .A(n1089), .B(n1090), .Z(n1088) );
NAND2_X1 U786 ( .A1(KEYINPUT14), .A2(n1091), .ZN(n1089) );
XOR2_X1 U787 ( .A(n1092), .B(n1093), .Z(n1087) );
NOR3_X1 U788 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
AND3_X1 U789 ( .A1(G140), .A2(G125), .A3(KEYINPUT41), .ZN(n1096) );
NOR2_X1 U790 ( .A1(G140), .A2(n1097), .ZN(n1095) );
NOR2_X1 U791 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
INV_X1 U792 ( .A(KEYINPUT41), .ZN(n1099) );
AND2_X1 U793 ( .A1(n1100), .A2(KEYINPUT58), .ZN(n1098) );
NOR2_X1 U794 ( .A1(KEYINPUT58), .A2(n1100), .ZN(n1094) );
NAND2_X1 U795 ( .A1(KEYINPUT35), .A2(n1101), .ZN(n1092) );
NAND2_X1 U796 ( .A1(n1102), .A2(n1103), .ZN(n1082) );
NAND2_X1 U797 ( .A1(G953), .A2(n1104), .ZN(n1080) );
NAND2_X1 U798 ( .A1(G900), .A2(G227), .ZN(n1104) );
XOR2_X1 U799 ( .A(n1105), .B(n1106), .Z(G69) );
XOR2_X1 U800 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U801 ( .A1(n1109), .A2(G953), .ZN(n1108) );
NOR3_X1 U802 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
NAND3_X1 U803 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1107) );
XOR2_X1 U804 ( .A(KEYINPUT40), .B(n1116), .Z(n1115) );
NOR2_X1 U805 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U806 ( .A1(n1117), .A2(n1118), .ZN(n1113) );
XNOR2_X1 U807 ( .A(n1119), .B(KEYINPUT16), .ZN(n1118) );
XOR2_X1 U808 ( .A(n1120), .B(KEYINPUT8), .Z(n1117) );
NAND2_X1 U809 ( .A1(G953), .A2(n1121), .ZN(n1105) );
NAND2_X1 U810 ( .A1(G898), .A2(G224), .ZN(n1121) );
NOR2_X1 U811 ( .A1(n1122), .A2(n1123), .ZN(G66) );
XOR2_X1 U812 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND2_X1 U813 ( .A1(n1126), .A2(n1127), .ZN(n1124) );
NOR2_X1 U814 ( .A1(n1128), .A2(n1129), .ZN(G63) );
XNOR2_X1 U815 ( .A(n1130), .B(n1131), .ZN(n1129) );
XOR2_X1 U816 ( .A(n1132), .B(KEYINPUT36), .Z(n1131) );
NAND2_X1 U817 ( .A1(n1126), .A2(G478), .ZN(n1132) );
NOR2_X1 U818 ( .A1(G952), .A2(n1133), .ZN(n1128) );
XNOR2_X1 U819 ( .A(KEYINPUT60), .B(n1102), .ZN(n1133) );
NOR2_X1 U820 ( .A1(n1122), .A2(n1134), .ZN(G60) );
XNOR2_X1 U821 ( .A(n1135), .B(n1136), .ZN(n1134) );
XOR2_X1 U822 ( .A(n1137), .B(KEYINPUT28), .Z(n1136) );
NAND2_X1 U823 ( .A1(n1126), .A2(G475), .ZN(n1137) );
XNOR2_X1 U824 ( .A(G104), .B(n1138), .ZN(G6) );
NOR3_X1 U825 ( .A1(n1122), .A2(n1139), .A3(n1140), .ZN(G57) );
NOR2_X1 U826 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NOR2_X1 U827 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NOR3_X1 U828 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(n1144) );
AND2_X1 U829 ( .A1(n1145), .A2(n1146), .ZN(n1143) );
INV_X1 U830 ( .A(KEYINPUT10), .ZN(n1145) );
NOR2_X1 U831 ( .A1(n1148), .A2(n1149), .ZN(n1139) );
NOR2_X1 U832 ( .A1(n1146), .A2(n1147), .ZN(n1148) );
INV_X1 U833 ( .A(KEYINPUT39), .ZN(n1147) );
XNOR2_X1 U834 ( .A(n1150), .B(n1151), .ZN(n1146) );
AND2_X1 U835 ( .A1(G472), .A2(n1126), .ZN(n1151) );
NAND2_X1 U836 ( .A1(KEYINPUT22), .A2(n1152), .ZN(n1150) );
XOR2_X1 U837 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U838 ( .A1(KEYINPUT62), .A2(n1155), .ZN(n1153) );
NOR2_X1 U839 ( .A1(n1122), .A2(n1156), .ZN(G54) );
XOR2_X1 U840 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U841 ( .A(n1159), .B(n1160), .ZN(n1158) );
NAND2_X1 U842 ( .A1(n1126), .A2(G469), .ZN(n1160) );
XOR2_X1 U843 ( .A(n1161), .B(n1162), .Z(n1157) );
NAND2_X1 U844 ( .A1(KEYINPUT34), .A2(n1101), .ZN(n1161) );
NOR2_X1 U845 ( .A1(n1122), .A2(n1163), .ZN(G51) );
XOR2_X1 U846 ( .A(n1164), .B(n1165), .Z(n1163) );
XNOR2_X1 U847 ( .A(n1166), .B(n1167), .ZN(n1165) );
XOR2_X1 U848 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND3_X1 U849 ( .A1(n1126), .A2(n1170), .A3(KEYINPUT57), .ZN(n1168) );
NOR2_X1 U850 ( .A1(n1171), .A2(n1037), .ZN(n1126) );
NOR4_X1 U851 ( .A1(n1172), .A2(n1110), .A3(n1103), .A4(n1112), .ZN(n1037) );
NAND4_X1 U852 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1112) );
NAND2_X1 U853 ( .A1(n1027), .A2(n1177), .ZN(n1176) );
INV_X1 U854 ( .A(KEYINPUT19), .ZN(n1177) );
NOR2_X1 U855 ( .A1(n1066), .A2(n1178), .ZN(n1027) );
NAND3_X1 U856 ( .A1(n1179), .A2(n1178), .A3(KEYINPUT19), .ZN(n1175) );
NAND4_X1 U857 ( .A1(n1180), .A2(n1078), .A3(n1050), .A4(n1181), .ZN(n1178) );
NAND2_X1 U858 ( .A1(n1182), .A2(n1183), .ZN(n1173) );
NAND2_X1 U859 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NAND2_X1 U860 ( .A1(n1186), .A2(n1044), .ZN(n1185) );
NAND2_X1 U861 ( .A1(n1046), .A2(n1187), .ZN(n1184) );
NAND4_X1 U862 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1103) );
NOR4_X1 U863 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
INV_X1 U864 ( .A(n1196), .ZN(n1195) );
AND2_X1 U865 ( .A1(n1197), .A2(n1198), .ZN(n1190) );
NAND4_X1 U866 ( .A1(n1199), .A2(n1200), .A3(n1187), .A4(n1201), .ZN(n1189) );
NOR2_X1 U867 ( .A1(n1053), .A2(n1066), .ZN(n1201) );
INV_X1 U868 ( .A(n1078), .ZN(n1053) );
NAND2_X1 U869 ( .A1(KEYINPUT7), .A2(n1202), .ZN(n1200) );
NAND2_X1 U870 ( .A1(n1203), .A2(n1204), .ZN(n1199) );
INV_X1 U871 ( .A(KEYINPUT7), .ZN(n1204) );
NAND2_X1 U872 ( .A1(n1205), .A2(n1061), .ZN(n1203) );
NAND2_X1 U873 ( .A1(n1206), .A2(n1039), .ZN(n1188) );
XNOR2_X1 U874 ( .A(n1207), .B(KEYINPUT12), .ZN(n1206) );
NAND3_X1 U875 ( .A1(n1208), .A2(n1209), .A3(n1138), .ZN(n1110) );
NAND4_X1 U876 ( .A1(n1186), .A2(n1210), .A3(n1180), .A4(n1050), .ZN(n1138) );
XOR2_X1 U877 ( .A(n1111), .B(KEYINPUT24), .Z(n1172) );
XOR2_X1 U878 ( .A(n1211), .B(n1212), .Z(n1164) );
XNOR2_X1 U879 ( .A(KEYINPUT6), .B(n1100), .ZN(n1212) );
NOR2_X1 U880 ( .A1(n1102), .A2(G952), .ZN(n1122) );
XNOR2_X1 U881 ( .A(G146), .B(n1213), .ZN(G48) );
NAND2_X1 U882 ( .A1(KEYINPUT37), .A2(n1194), .ZN(n1213) );
NOR4_X1 U883 ( .A1(n1214), .A2(n1202), .A3(n1052), .A4(n1066), .ZN(n1194) );
XOR2_X1 U884 ( .A(G143), .B(n1215), .Z(G45) );
NOR2_X1 U885 ( .A1(KEYINPUT1), .A2(n1198), .ZN(n1215) );
NAND3_X1 U886 ( .A1(n1216), .A2(n1044), .A3(n1217), .ZN(n1198) );
NOR3_X1 U887 ( .A1(n1066), .A2(n1218), .A3(n1219), .ZN(n1217) );
INV_X1 U888 ( .A(n1179), .ZN(n1066) );
XNOR2_X1 U889 ( .A(G140), .B(n1220), .ZN(G42) );
NAND2_X1 U890 ( .A1(n1207), .A2(n1039), .ZN(n1220) );
NOR3_X1 U891 ( .A1(n1052), .A2(n1055), .A3(n1202), .ZN(n1207) );
INV_X1 U892 ( .A(n1221), .ZN(n1055) );
XNOR2_X1 U893 ( .A(G137), .B(n1197), .ZN(G39) );
NAND4_X1 U894 ( .A1(n1046), .A2(n1187), .A3(n1216), .A4(n1039), .ZN(n1197) );
XNOR2_X1 U895 ( .A(G134), .B(n1222), .ZN(G36) );
NOR2_X1 U896 ( .A1(n1193), .A2(KEYINPUT47), .ZN(n1222) );
AND2_X1 U897 ( .A1(n1223), .A2(n1078), .ZN(n1193) );
XOR2_X1 U898 ( .A(G131), .B(n1192), .Z(G33) );
AND2_X1 U899 ( .A1(n1223), .A2(n1186), .ZN(n1192) );
AND3_X1 U900 ( .A1(n1044), .A2(n1039), .A3(n1216), .ZN(n1223) );
AND2_X1 U901 ( .A1(n1069), .A2(n1224), .ZN(n1039) );
NAND2_X1 U902 ( .A1(G214), .A2(n1068), .ZN(n1224) );
XNOR2_X1 U903 ( .A(G128), .B(n1225), .ZN(G30) );
NAND4_X1 U904 ( .A1(n1187), .A2(n1216), .A3(n1179), .A4(n1078), .ZN(n1225) );
INV_X1 U905 ( .A(n1202), .ZN(n1216) );
NAND2_X1 U906 ( .A1(n1180), .A2(n1205), .ZN(n1202) );
XNOR2_X1 U907 ( .A(G101), .B(n1174), .ZN(G3) );
NAND2_X1 U908 ( .A1(n1226), .A2(n1044), .ZN(n1174) );
XNOR2_X1 U909 ( .A(G125), .B(n1196), .ZN(G27) );
NAND4_X1 U910 ( .A1(n1221), .A2(n1205), .A3(n1179), .A4(n1227), .ZN(n1196) );
NOR2_X1 U911 ( .A1(n1228), .A2(n1052), .ZN(n1227) );
INV_X1 U912 ( .A(n1186), .ZN(n1052) );
NAND2_X1 U913 ( .A1(n1043), .A2(n1229), .ZN(n1205) );
OR4_X1 U914 ( .A1(n1086), .A2(n1171), .A3(n1230), .A4(G900), .ZN(n1229) );
XNOR2_X1 U915 ( .A(n1208), .B(n1231), .ZN(G24) );
NOR2_X1 U916 ( .A1(KEYINPUT30), .A2(n1232), .ZN(n1231) );
NAND4_X1 U917 ( .A1(n1182), .A2(n1050), .A3(n1233), .A4(n1234), .ZN(n1208) );
NOR2_X1 U918 ( .A1(n1235), .A2(n1236), .ZN(n1050) );
XOR2_X1 U919 ( .A(G119), .B(n1237), .Z(G21) );
NOR3_X1 U920 ( .A1(n1079), .A2(n1238), .A3(n1239), .ZN(n1237) );
XNOR2_X1 U921 ( .A(n1187), .B(KEYINPUT46), .ZN(n1238) );
INV_X1 U922 ( .A(n1046), .ZN(n1079) );
XNOR2_X1 U923 ( .A(G116), .B(n1209), .ZN(G18) );
NAND3_X1 U924 ( .A1(n1182), .A2(n1078), .A3(n1044), .ZN(n1209) );
NOR2_X1 U925 ( .A1(n1234), .A2(n1219), .ZN(n1078) );
INV_X1 U926 ( .A(n1233), .ZN(n1219) );
INV_X1 U927 ( .A(n1239), .ZN(n1182) );
NAND2_X1 U928 ( .A1(n1210), .A2(n1038), .ZN(n1239) );
XNOR2_X1 U929 ( .A(G113), .B(n1240), .ZN(G15) );
NAND4_X1 U930 ( .A1(n1241), .A2(n1186), .A3(n1044), .A4(n1210), .ZN(n1240) );
AND2_X1 U931 ( .A1(n1236), .A2(n1070), .ZN(n1044) );
NOR2_X1 U932 ( .A1(n1233), .A2(n1218), .ZN(n1186) );
INV_X1 U933 ( .A(n1234), .ZN(n1218) );
XNOR2_X1 U934 ( .A(n1038), .B(KEYINPUT53), .ZN(n1241) );
INV_X1 U935 ( .A(n1228), .ZN(n1038) );
NAND2_X1 U936 ( .A1(n1076), .A2(n1063), .ZN(n1228) );
INV_X1 U937 ( .A(n1064), .ZN(n1076) );
XNOR2_X1 U938 ( .A(n1111), .B(n1242), .ZN(G12) );
NAND2_X1 U939 ( .A1(KEYINPUT51), .A2(G110), .ZN(n1242) );
AND2_X1 U940 ( .A1(n1226), .A2(n1221), .ZN(n1111) );
NAND2_X1 U941 ( .A1(n1243), .A2(n1244), .ZN(n1221) );
OR3_X1 U942 ( .A1(n1236), .A2(n1070), .A3(KEYINPUT25), .ZN(n1244) );
INV_X1 U943 ( .A(n1235), .ZN(n1070) );
NAND2_X1 U944 ( .A1(KEYINPUT25), .A2(n1187), .ZN(n1243) );
INV_X1 U945 ( .A(n1214), .ZN(n1187) );
NAND2_X1 U946 ( .A1(n1236), .A2(n1235), .ZN(n1214) );
XNOR2_X1 U947 ( .A(n1245), .B(n1127), .ZN(n1235) );
AND2_X1 U948 ( .A1(G217), .A2(n1246), .ZN(n1127) );
NAND2_X1 U949 ( .A1(n1125), .A2(n1171), .ZN(n1245) );
XNOR2_X1 U950 ( .A(n1247), .B(n1248), .ZN(n1125) );
NOR2_X1 U951 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
NOR2_X1 U952 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XNOR2_X1 U953 ( .A(KEYINPUT56), .B(n1253), .ZN(n1252) );
NOR3_X1 U954 ( .A1(n1254), .A2(G953), .A3(n1255), .ZN(n1251) );
NOR4_X1 U955 ( .A1(G953), .A2(n1255), .A3(n1254), .A4(n1253), .ZN(n1249) );
INV_X1 U956 ( .A(G221), .ZN(n1254) );
NAND2_X1 U957 ( .A1(n1256), .A2(KEYINPUT48), .ZN(n1247) );
XOR2_X1 U958 ( .A(n1257), .B(n1258), .Z(n1256) );
XOR2_X1 U959 ( .A(G119), .B(n1259), .Z(n1258) );
XOR2_X1 U960 ( .A(G140), .B(G128), .Z(n1259) );
XNOR2_X1 U961 ( .A(n1260), .B(n1261), .ZN(n1257) );
XNOR2_X1 U962 ( .A(n1262), .B(n1263), .ZN(n1261) );
NOR2_X1 U963 ( .A1(KEYINPUT42), .A2(n1100), .ZN(n1263) );
NAND2_X1 U964 ( .A1(KEYINPUT5), .A2(n1264), .ZN(n1262) );
XOR2_X1 U965 ( .A(n1077), .B(n1265), .Z(n1236) );
NOR2_X1 U966 ( .A1(G472), .A2(KEYINPUT15), .ZN(n1265) );
NAND2_X1 U967 ( .A1(n1266), .A2(n1171), .ZN(n1077) );
XNOR2_X1 U968 ( .A(n1267), .B(n1149), .ZN(n1266) );
INV_X1 U969 ( .A(n1141), .ZN(n1149) );
XNOR2_X1 U970 ( .A(n1268), .B(G101), .ZN(n1141) );
NAND2_X1 U971 ( .A1(n1269), .A2(G210), .ZN(n1268) );
XNOR2_X1 U972 ( .A(n1155), .B(n1154), .ZN(n1267) );
XNOR2_X1 U973 ( .A(n1270), .B(n1169), .ZN(n1154) );
XOR2_X1 U974 ( .A(G113), .B(n1271), .Z(n1155) );
XOR2_X1 U975 ( .A(G119), .B(G116), .Z(n1271) );
AND3_X1 U976 ( .A1(n1210), .A2(n1180), .A3(n1046), .ZN(n1226) );
NOR2_X1 U977 ( .A1(n1233), .A2(n1234), .ZN(n1046) );
XNOR2_X1 U978 ( .A(n1272), .B(G475), .ZN(n1234) );
NAND2_X1 U979 ( .A1(n1135), .A2(n1171), .ZN(n1272) );
XNOR2_X1 U980 ( .A(n1273), .B(n1274), .ZN(n1135) );
XNOR2_X1 U981 ( .A(n1091), .B(n1275), .ZN(n1274) );
XOR2_X1 U982 ( .A(n1276), .B(n1277), .Z(n1275) );
NOR2_X1 U983 ( .A1(G122), .A2(KEYINPUT44), .ZN(n1277) );
NAND2_X1 U984 ( .A1(n1269), .A2(G214), .ZN(n1276) );
NOR2_X1 U985 ( .A1(G953), .A2(G237), .ZN(n1269) );
XOR2_X1 U986 ( .A(n1278), .B(n1279), .Z(n1273) );
XOR2_X1 U987 ( .A(G143), .B(G113), .Z(n1279) );
XNOR2_X1 U988 ( .A(G104), .B(n1280), .ZN(n1278) );
NOR2_X1 U989 ( .A1(KEYINPUT27), .A2(n1281), .ZN(n1280) );
XNOR2_X1 U990 ( .A(n1260), .B(n1282), .ZN(n1281) );
XNOR2_X1 U991 ( .A(G125), .B(n1283), .ZN(n1282) );
NOR2_X1 U992 ( .A1(G140), .A2(KEYINPUT17), .ZN(n1283) );
XNOR2_X1 U993 ( .A(n1284), .B(n1285), .ZN(n1233) );
XOR2_X1 U994 ( .A(KEYINPUT0), .B(G478), .Z(n1285) );
NAND2_X1 U995 ( .A1(n1130), .A2(n1171), .ZN(n1284) );
XNOR2_X1 U996 ( .A(n1286), .B(n1287), .ZN(n1130) );
XNOR2_X1 U997 ( .A(n1288), .B(n1289), .ZN(n1287) );
XNOR2_X1 U998 ( .A(KEYINPUT63), .B(n1290), .ZN(n1289) );
INV_X1 U999 ( .A(G134), .ZN(n1290) );
XOR2_X1 U1000 ( .A(n1291), .B(n1292), .Z(n1286) );
XOR2_X1 U1001 ( .A(n1293), .B(n1294), .Z(n1291) );
AND3_X1 U1002 ( .A1(G217), .A2(n1102), .A3(G234), .ZN(n1294) );
NAND3_X1 U1003 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1293) );
NAND2_X1 U1004 ( .A1(KEYINPUT33), .A2(G116), .ZN(n1297) );
NAND3_X1 U1005 ( .A1(n1298), .A2(n1299), .A3(n1232), .ZN(n1296) );
INV_X1 U1006 ( .A(KEYINPUT33), .ZN(n1299) );
OR2_X1 U1007 ( .A1(n1232), .A2(n1298), .ZN(n1295) );
NOR2_X1 U1008 ( .A1(G116), .A2(KEYINPUT59), .ZN(n1298) );
INV_X1 U1009 ( .A(n1061), .ZN(n1180) );
NAND2_X1 U1010 ( .A1(n1064), .A2(n1063), .ZN(n1061) );
NAND2_X1 U1011 ( .A1(G221), .A2(n1246), .ZN(n1063) );
NAND2_X1 U1012 ( .A1(G234), .A2(n1300), .ZN(n1246) );
XNOR2_X1 U1013 ( .A(n1301), .B(G469), .ZN(n1064) );
NAND2_X1 U1014 ( .A1(n1302), .A2(n1171), .ZN(n1301) );
XOR2_X1 U1015 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U1016 ( .A(n1162), .B(n1101), .ZN(n1304) );
XNOR2_X1 U1017 ( .A(n1305), .B(n1306), .ZN(n1162) );
XNOR2_X1 U1018 ( .A(G140), .B(n1264), .ZN(n1306) );
XNOR2_X1 U1019 ( .A(n1307), .B(n1270), .ZN(n1305) );
XNOR2_X1 U1020 ( .A(n1090), .B(n1091), .ZN(n1270) );
XOR2_X1 U1021 ( .A(G131), .B(KEYINPUT4), .Z(n1091) );
XOR2_X1 U1022 ( .A(G134), .B(n1308), .Z(n1090) );
XNOR2_X1 U1023 ( .A(KEYINPUT20), .B(n1253), .ZN(n1308) );
INV_X1 U1024 ( .A(G137), .ZN(n1253) );
NAND3_X1 U1025 ( .A1(n1309), .A2(n1310), .A3(n1311), .ZN(n1307) );
NAND2_X1 U1026 ( .A1(n1312), .A2(n1313), .ZN(n1310) );
INV_X1 U1027 ( .A(KEYINPUT50), .ZN(n1313) );
NAND2_X1 U1028 ( .A1(n1314), .A2(KEYINPUT50), .ZN(n1309) );
XOR2_X1 U1029 ( .A(G101), .B(n1315), .Z(n1314) );
NOR2_X1 U1030 ( .A1(G104), .A2(n1288), .ZN(n1315) );
XOR2_X1 U1031 ( .A(n1316), .B(KEYINPUT45), .Z(n1303) );
NAND2_X1 U1032 ( .A1(KEYINPUT18), .A2(n1159), .ZN(n1316) );
AND2_X1 U1033 ( .A1(G227), .A2(n1102), .ZN(n1159) );
AND2_X1 U1034 ( .A1(n1179), .A2(n1181), .ZN(n1210) );
NAND2_X1 U1035 ( .A1(n1043), .A2(n1317), .ZN(n1181) );
OR3_X1 U1036 ( .A1(n1171), .A2(n1230), .A3(n1114), .ZN(n1317) );
OR2_X1 U1037 ( .A1(n1086), .A2(G898), .ZN(n1114) );
XOR2_X1 U1038 ( .A(G953), .B(KEYINPUT13), .Z(n1086) );
INV_X1 U1039 ( .A(n1049), .ZN(n1043) );
NOR3_X1 U1040 ( .A1(n1033), .A2(n1230), .A3(n1318), .ZN(n1049) );
INV_X1 U1041 ( .A(G952), .ZN(n1318) );
NOR2_X1 U1042 ( .A1(n1319), .A2(n1255), .ZN(n1230) );
INV_X1 U1043 ( .A(G234), .ZN(n1255) );
XNOR2_X1 U1044 ( .A(G953), .B(KEYINPUT9), .ZN(n1033) );
NOR2_X1 U1045 ( .A1(n1069), .A2(n1320), .ZN(n1179) );
AND2_X1 U1046 ( .A1(G214), .A2(n1068), .ZN(n1320) );
XOR2_X1 U1047 ( .A(n1321), .B(n1170), .Z(n1069) );
AND2_X1 U1048 ( .A1(G210), .A2(n1068), .ZN(n1170) );
NAND2_X1 U1049 ( .A1(n1300), .A2(n1319), .ZN(n1068) );
INV_X1 U1050 ( .A(G237), .ZN(n1319) );
XNOR2_X1 U1051 ( .A(G902), .B(KEYINPUT21), .ZN(n1300) );
NAND2_X1 U1052 ( .A1(n1322), .A2(n1171), .ZN(n1321) );
INV_X1 U1053 ( .A(G902), .ZN(n1171) );
XNOR2_X1 U1054 ( .A(n1323), .B(n1324), .ZN(n1322) );
INV_X1 U1055 ( .A(n1166), .ZN(n1324) );
XNOR2_X1 U1056 ( .A(n1120), .B(n1325), .ZN(n1166) );
NOR2_X1 U1057 ( .A1(KEYINPUT26), .A2(n1119), .ZN(n1325) );
XNOR2_X1 U1058 ( .A(n1326), .B(n1327), .ZN(n1119) );
NOR2_X1 U1059 ( .A1(n1328), .A2(n1312), .ZN(n1327) );
NAND2_X1 U1060 ( .A1(n1329), .A2(n1330), .ZN(n1312) );
OR3_X1 U1061 ( .A1(G101), .A2(G104), .A3(G107), .ZN(n1330) );
NAND2_X1 U1062 ( .A1(n1331), .A2(G107), .ZN(n1329) );
XOR2_X1 U1063 ( .A(G104), .B(G101), .Z(n1331) );
INV_X1 U1064 ( .A(n1311), .ZN(n1328) );
NAND3_X1 U1065 ( .A1(G101), .A2(n1288), .A3(G104), .ZN(n1311) );
INV_X1 U1066 ( .A(G107), .ZN(n1288) );
XOR2_X1 U1067 ( .A(n1332), .B(G113), .Z(n1326) );
NAND2_X1 U1068 ( .A1(n1333), .A2(KEYINPUT29), .ZN(n1332) );
XNOR2_X1 U1069 ( .A(G119), .B(n1334), .ZN(n1333) );
NOR2_X1 U1070 ( .A1(G116), .A2(KEYINPUT31), .ZN(n1334) );
XNOR2_X1 U1071 ( .A(n1335), .B(n1264), .ZN(n1120) );
INV_X1 U1072 ( .A(G110), .ZN(n1264) );
NAND2_X1 U1073 ( .A1(KEYINPUT2), .A2(n1232), .ZN(n1335) );
INV_X1 U1074 ( .A(G122), .ZN(n1232) );
NAND2_X1 U1075 ( .A1(n1336), .A2(n1337), .ZN(n1323) );
NAND2_X1 U1076 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
XOR2_X1 U1077 ( .A(n1340), .B(n1169), .Z(n1339) );
XNOR2_X1 U1078 ( .A(KEYINPUT3), .B(n1211), .ZN(n1338) );
XOR2_X1 U1079 ( .A(n1341), .B(KEYINPUT61), .Z(n1336) );
NAND2_X1 U1080 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
XOR2_X1 U1081 ( .A(KEYINPUT3), .B(n1211), .Z(n1343) );
AND2_X1 U1082 ( .A1(G224), .A2(n1102), .ZN(n1211) );
INV_X1 U1083 ( .A(G953), .ZN(n1102) );
XNOR2_X1 U1084 ( .A(n1340), .B(n1169), .ZN(n1342) );
XOR2_X1 U1085 ( .A(n1101), .B(KEYINPUT23), .Z(n1169) );
XNOR2_X1 U1086 ( .A(n1292), .B(n1344), .ZN(n1101) );
INV_X1 U1087 ( .A(n1260), .ZN(n1344) );
XOR2_X1 U1088 ( .A(G146), .B(KEYINPUT49), .Z(n1260) );
XOR2_X1 U1089 ( .A(G128), .B(G143), .Z(n1292) );
NOR2_X1 U1090 ( .A1(KEYINPUT38), .A2(n1100), .ZN(n1340) );
INV_X1 U1091 ( .A(G125), .ZN(n1100) );
endmodule


