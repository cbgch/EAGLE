//Key = 0010110010101101010001001101100001100100100000011100011000110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349;

XNOR2_X1 U745 ( .A(G107), .B(n1027), .ZN(G9) );
NOR2_X1 U746 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR4_X1 U747 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1029) );
XOR2_X1 U748 ( .A(KEYINPUT40), .B(G952), .Z(n1033) );
XOR2_X1 U749 ( .A(KEYINPUT57), .B(n1034), .Z(n1032) );
NOR2_X1 U750 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U751 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U752 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U753 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U754 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR3_X1 U755 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1043) );
NOR2_X1 U756 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U757 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR3_X1 U758 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1046) );
NOR2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1045) );
XNOR2_X1 U760 ( .A(KEYINPUT47), .B(n1054), .ZN(n1056) );
NOR4_X1 U761 ( .A1(n1054), .A2(n1057), .A3(n1049), .A4(n1058), .ZN(n1041) );
NOR3_X1 U762 ( .A1(n1049), .A2(n1059), .A3(n1054), .ZN(n1037) );
NOR2_X1 U763 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U764 ( .A1(n1062), .A2(n1040), .ZN(n1061) );
NOR2_X1 U765 ( .A1(n1063), .A2(n1044), .ZN(n1060) );
NOR2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U767 ( .A1(n1066), .A2(n1067), .ZN(n1031) );
NOR3_X1 U768 ( .A1(n1068), .A2(G953), .A3(n1069), .ZN(n1028) );
INV_X1 U769 ( .A(n1066), .ZN(n1069) );
NAND4_X1 U770 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1066) );
XOR2_X1 U771 ( .A(n1074), .B(n1075), .Z(n1073) );
NAND2_X1 U772 ( .A1(KEYINPUT62), .A2(n1076), .ZN(n1075) );
XOR2_X1 U773 ( .A(n1077), .B(KEYINPUT49), .Z(n1070) );
NAND4_X1 U774 ( .A1(n1078), .A2(n1052), .A3(n1079), .A4(n1058), .ZN(n1077) );
AND2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U776 ( .A(n1082), .B(n1083), .Z(n1078) );
XNOR2_X1 U777 ( .A(G952), .B(KEYINPUT12), .ZN(n1068) );
XOR2_X1 U778 ( .A(n1084), .B(n1085), .Z(G72) );
XOR2_X1 U779 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U780 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U781 ( .A(n1090), .B(n1091), .Z(n1089) );
XNOR2_X1 U782 ( .A(n1092), .B(n1093), .ZN(n1091) );
XOR2_X1 U783 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U784 ( .A1(KEYINPUT48), .A2(G125), .ZN(n1094) );
XOR2_X1 U785 ( .A(G131), .B(n1096), .Z(n1090) );
XNOR2_X1 U786 ( .A(KEYINPUT63), .B(n1097), .ZN(n1096) );
NAND3_X1 U787 ( .A1(n1098), .A2(n1067), .A3(KEYINPUT28), .ZN(n1086) );
NAND2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U789 ( .A(n1101), .B(KEYINPUT61), .ZN(n1099) );
NAND2_X1 U790 ( .A1(G953), .A2(n1102), .ZN(n1084) );
NAND2_X1 U791 ( .A1(G900), .A2(G227), .ZN(n1102) );
XOR2_X1 U792 ( .A(n1103), .B(n1104), .Z(G69) );
XOR2_X1 U793 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U794 ( .A1(n1107), .A2(n1067), .ZN(n1106) );
NOR2_X1 U795 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND3_X1 U796 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1105) );
XOR2_X1 U797 ( .A(n1113), .B(KEYINPUT42), .Z(n1112) );
OR2_X1 U798 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U799 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
XNOR2_X1 U800 ( .A(n1116), .B(n1117), .ZN(n1114) );
XNOR2_X1 U801 ( .A(KEYINPUT37), .B(n1118), .ZN(n1116) );
NOR2_X1 U802 ( .A1(KEYINPUT1), .A2(n1119), .ZN(n1118) );
NAND2_X1 U803 ( .A1(G953), .A2(n1109), .ZN(n1110) );
NAND2_X1 U804 ( .A1(n1067), .A2(n1120), .ZN(n1103) );
NAND2_X1 U805 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U806 ( .A(n1027), .B(KEYINPUT43), .Z(n1121) );
NOR2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(G66) );
XOR2_X1 U808 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U809 ( .A1(n1074), .A2(n1127), .ZN(n1126) );
NAND2_X1 U810 ( .A1(KEYINPUT34), .A2(n1128), .ZN(n1125) );
NOR2_X1 U811 ( .A1(n1123), .A2(n1129), .ZN(G63) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND3_X1 U813 ( .A1(n1132), .A2(n1030), .A3(G478), .ZN(n1130) );
XNOR2_X1 U814 ( .A(KEYINPUT35), .B(n1133), .ZN(n1132) );
NOR2_X1 U815 ( .A1(n1123), .A2(n1134), .ZN(G60) );
XNOR2_X1 U816 ( .A(n1135), .B(n1136), .ZN(n1134) );
NOR2_X1 U817 ( .A1(n1137), .A2(n1127), .ZN(n1136) );
XNOR2_X1 U818 ( .A(G104), .B(n1138), .ZN(G6) );
NOR2_X1 U819 ( .A1(n1123), .A2(n1139), .ZN(G57) );
XOR2_X1 U820 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U821 ( .A(n1142), .B(n1143), .ZN(n1141) );
NOR2_X1 U822 ( .A1(n1144), .A2(n1127), .ZN(n1143) );
XOR2_X1 U823 ( .A(n1145), .B(n1146), .Z(n1140) );
NOR4_X1 U824 ( .A1(KEYINPUT60), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1146) );
INV_X1 U825 ( .A(n1150), .ZN(n1148) );
INV_X1 U826 ( .A(n1151), .ZN(n1147) );
XNOR2_X1 U827 ( .A(G101), .B(KEYINPUT50), .ZN(n1145) );
NOR2_X1 U828 ( .A1(n1123), .A2(n1152), .ZN(G54) );
NOR2_X1 U829 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U830 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U831 ( .A1(n1157), .A2(KEYINPUT22), .ZN(n1156) );
NOR2_X1 U832 ( .A1(n1158), .A2(n1127), .ZN(n1155) );
AND2_X1 U833 ( .A1(n1157), .A2(KEYINPUT22), .ZN(n1153) );
AND2_X1 U834 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NAND2_X1 U835 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XNOR2_X1 U836 ( .A(n1163), .B(n1164), .ZN(n1162) );
XOR2_X1 U837 ( .A(n1165), .B(KEYINPUT13), .Z(n1161) );
NAND2_X1 U838 ( .A1(n1166), .A2(n1165), .ZN(n1159) );
XOR2_X1 U839 ( .A(n1167), .B(KEYINPUT6), .Z(n1165) );
XNOR2_X1 U840 ( .A(n1163), .B(n1168), .ZN(n1166) );
NOR2_X1 U841 ( .A1(KEYINPUT0), .A2(n1169), .ZN(n1163) );
NOR2_X1 U842 ( .A1(n1123), .A2(n1170), .ZN(G51) );
XOR2_X1 U843 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U844 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U845 ( .A(KEYINPUT26), .B(n1175), .Z(n1174) );
AND2_X1 U846 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NOR2_X1 U847 ( .A1(n1176), .A2(n1177), .ZN(n1173) );
XOR2_X1 U848 ( .A(n1178), .B(n1179), .Z(n1177) );
NOR2_X1 U849 ( .A1(n1083), .A2(n1127), .ZN(n1171) );
NAND2_X1 U850 ( .A1(G902), .A2(n1030), .ZN(n1127) );
NAND4_X1 U851 ( .A1(n1180), .A2(n1101), .A3(n1122), .A4(n1027), .ZN(n1030) );
NAND3_X1 U852 ( .A1(n1050), .A2(n1181), .A3(n1182), .ZN(n1027) );
AND4_X1 U853 ( .A1(n1138), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1122) );
NOR4_X1 U854 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1185) );
NOR4_X1 U855 ( .A1(n1190), .A2(n1055), .A3(n1044), .A4(n1191), .ZN(n1189) );
XNOR2_X1 U856 ( .A(n1192), .B(KEYINPUT10), .ZN(n1190) );
INV_X1 U857 ( .A(n1193), .ZN(n1188) );
AND2_X1 U858 ( .A1(KEYINPUT5), .A2(n1194), .ZN(n1187) );
NOR4_X1 U859 ( .A1(KEYINPUT5), .A2(n1195), .A3(n1196), .A4(n1040), .ZN(n1186) );
NOR2_X1 U860 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NOR2_X1 U861 ( .A1(n1199), .A2(n1200), .ZN(n1184) );
NAND3_X1 U862 ( .A1(n1182), .A2(n1181), .A3(n1051), .ZN(n1138) );
INV_X1 U863 ( .A(n1040), .ZN(n1181) );
AND4_X1 U864 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1101) );
NAND3_X1 U865 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1201) );
XNOR2_X1 U866 ( .A(KEYINPUT45), .B(n1062), .ZN(n1205) );
XNOR2_X1 U867 ( .A(n1100), .B(KEYINPUT4), .ZN(n1180) );
AND4_X1 U868 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1100) );
NAND2_X1 U869 ( .A1(n1212), .A2(n1213), .ZN(n1210) );
XOR2_X1 U870 ( .A(n1214), .B(KEYINPUT15), .Z(n1212) );
OR2_X1 U871 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND3_X1 U872 ( .A1(n1071), .A2(n1217), .A3(n1218), .ZN(n1209) );
XNOR2_X1 U873 ( .A(KEYINPUT31), .B(n1216), .ZN(n1217) );
NAND3_X1 U874 ( .A1(n1051), .A2(n1065), .A3(n1218), .ZN(n1208) );
NOR2_X1 U875 ( .A1(n1067), .A2(G952), .ZN(n1123) );
XNOR2_X1 U876 ( .A(n1219), .B(n1220), .ZN(G48) );
NOR4_X1 U877 ( .A1(KEYINPUT51), .A2(n1221), .A3(n1055), .A4(n1215), .ZN(n1220) );
NAND2_X1 U878 ( .A1(n1222), .A2(n1051), .ZN(n1215) );
XNOR2_X1 U879 ( .A(n1223), .B(KEYINPUT46), .ZN(n1221) );
XNOR2_X1 U880 ( .A(G143), .B(n1211), .ZN(G45) );
NAND3_X1 U881 ( .A1(n1064), .A2(n1222), .A3(n1224), .ZN(n1211) );
NOR3_X1 U882 ( .A1(n1055), .A2(n1197), .A3(n1198), .ZN(n1224) );
XOR2_X1 U883 ( .A(n1225), .B(n1226), .Z(G42) );
NOR2_X1 U884 ( .A1(KEYINPUT9), .A2(n1097), .ZN(n1226) );
NOR4_X1 U885 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1225) );
NOR2_X1 U886 ( .A1(KEYINPUT54), .A2(n1231), .ZN(n1228) );
AND2_X1 U887 ( .A1(n1049), .A2(n1222), .ZN(n1231) );
NOR2_X1 U888 ( .A1(n1218), .A2(n1232), .ZN(n1227) );
INV_X1 U889 ( .A(KEYINPUT54), .ZN(n1232) );
XNOR2_X1 U890 ( .A(G137), .B(n1233), .ZN(G39) );
NAND3_X1 U891 ( .A1(n1234), .A2(n1218), .A3(KEYINPUT24), .ZN(n1233) );
XNOR2_X1 U892 ( .A(G134), .B(n1202), .ZN(G36) );
NAND3_X1 U893 ( .A1(n1218), .A2(n1050), .A3(n1064), .ZN(n1202) );
XNOR2_X1 U894 ( .A(G131), .B(n1203), .ZN(G33) );
NAND3_X1 U895 ( .A1(n1218), .A2(n1051), .A3(n1064), .ZN(n1203) );
NOR2_X1 U896 ( .A1(n1049), .A2(n1235), .ZN(n1218) );
INV_X1 U897 ( .A(n1222), .ZN(n1235) );
NAND2_X1 U898 ( .A1(n1236), .A2(n1052), .ZN(n1049) );
NAND3_X1 U899 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(G30) );
OR2_X1 U900 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NAND3_X1 U901 ( .A1(n1241), .A2(n1240), .A3(G128), .ZN(n1238) );
NAND2_X1 U902 ( .A1(n1242), .A2(n1243), .ZN(n1237) );
NAND2_X1 U903 ( .A1(n1244), .A2(n1240), .ZN(n1242) );
INV_X1 U904 ( .A(KEYINPUT44), .ZN(n1240) );
XNOR2_X1 U905 ( .A(KEYINPUT33), .B(n1241), .ZN(n1244) );
NAND2_X1 U906 ( .A1(n1207), .A2(n1222), .ZN(n1241) );
NOR2_X1 U907 ( .A1(n1062), .A2(n1245), .ZN(n1222) );
AND3_X1 U908 ( .A1(n1050), .A2(n1213), .A3(n1223), .ZN(n1207) );
INV_X1 U909 ( .A(n1216), .ZN(n1223) );
INV_X1 U910 ( .A(n1055), .ZN(n1213) );
XNOR2_X1 U911 ( .A(G101), .B(n1183), .ZN(G3) );
NAND3_X1 U912 ( .A1(n1071), .A2(n1182), .A3(n1064), .ZN(n1183) );
NAND2_X1 U913 ( .A1(n1246), .A2(n1247), .ZN(G27) );
OR2_X1 U914 ( .A1(n1204), .A2(G125), .ZN(n1247) );
XOR2_X1 U915 ( .A(n1248), .B(KEYINPUT19), .Z(n1246) );
NAND2_X1 U916 ( .A1(G125), .A2(n1204), .ZN(n1248) );
NAND4_X1 U917 ( .A1(n1051), .A2(n1065), .A3(n1249), .A4(n1250), .ZN(n1204) );
NOR2_X1 U918 ( .A1(n1245), .A2(n1055), .ZN(n1249) );
INV_X1 U919 ( .A(n1206), .ZN(n1245) );
NAND2_X1 U920 ( .A1(n1036), .A2(n1251), .ZN(n1206) );
NAND3_X1 U921 ( .A1(G902), .A2(n1252), .A3(n1088), .ZN(n1251) );
NOR2_X1 U922 ( .A1(n1067), .A2(G900), .ZN(n1088) );
XOR2_X1 U923 ( .A(n1194), .B(n1253), .Z(G24) );
NOR2_X1 U924 ( .A1(KEYINPUT55), .A2(n1254), .ZN(n1253) );
NOR4_X1 U925 ( .A1(n1195), .A2(n1040), .A3(n1198), .A4(n1197), .ZN(n1194) );
NAND2_X1 U926 ( .A1(n1255), .A2(n1072), .ZN(n1040) );
XOR2_X1 U927 ( .A(G119), .B(n1256), .Z(G21) );
NOR2_X1 U928 ( .A1(n1195), .A2(n1191), .ZN(n1256) );
INV_X1 U929 ( .A(n1234), .ZN(n1191) );
NOR2_X1 U930 ( .A1(n1216), .A2(n1054), .ZN(n1234) );
NAND2_X1 U931 ( .A1(n1257), .A2(n1258), .ZN(n1216) );
INV_X1 U932 ( .A(n1259), .ZN(n1195) );
XOR2_X1 U933 ( .A(G116), .B(n1200), .Z(G18) );
AND3_X1 U934 ( .A1(n1064), .A2(n1050), .A3(n1259), .ZN(n1200) );
NOR3_X1 U935 ( .A1(n1055), .A2(n1192), .A3(n1044), .ZN(n1259) );
INV_X1 U936 ( .A(n1250), .ZN(n1044) );
NOR2_X1 U937 ( .A1(n1260), .A2(n1197), .ZN(n1050) );
XNOR2_X1 U938 ( .A(G113), .B(n1193), .ZN(G15) );
NAND4_X1 U939 ( .A1(n1064), .A2(n1051), .A3(n1261), .A4(n1250), .ZN(n1193) );
NOR2_X1 U940 ( .A1(n1057), .A2(n1262), .ZN(n1250) );
INV_X1 U941 ( .A(n1058), .ZN(n1262) );
NOR2_X1 U942 ( .A1(n1192), .A2(n1263), .ZN(n1261) );
INV_X1 U943 ( .A(n1230), .ZN(n1051) );
NAND2_X1 U944 ( .A1(n1197), .A2(n1260), .ZN(n1230) );
AND2_X1 U945 ( .A1(n1255), .A2(n1258), .ZN(n1064) );
XNOR2_X1 U946 ( .A(G110), .B(n1264), .ZN(G12) );
NAND2_X1 U947 ( .A1(KEYINPUT2), .A2(n1199), .ZN(n1264) );
AND3_X1 U948 ( .A1(n1071), .A2(n1182), .A3(n1065), .ZN(n1199) );
INV_X1 U949 ( .A(n1229), .ZN(n1065) );
NAND2_X1 U950 ( .A1(n1072), .A2(n1257), .ZN(n1229) );
XNOR2_X1 U951 ( .A(n1255), .B(KEYINPUT36), .ZN(n1257) );
XNOR2_X1 U952 ( .A(n1076), .B(n1074), .ZN(n1255) );
NAND2_X1 U953 ( .A1(G217), .A2(n1265), .ZN(n1074) );
NAND2_X1 U954 ( .A1(n1128), .A2(n1133), .ZN(n1076) );
XNOR2_X1 U955 ( .A(n1266), .B(n1267), .ZN(n1128) );
XOR2_X1 U956 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U957 ( .A(n1270), .B(n1271), .Z(n1269) );
NOR2_X1 U958 ( .A1(G140), .A2(KEYINPUT29), .ZN(n1271) );
AND3_X1 U959 ( .A1(G221), .A2(n1067), .A3(G234), .ZN(n1270) );
XOR2_X1 U960 ( .A(G110), .B(n1272), .Z(n1268) );
NOR2_X1 U961 ( .A1(KEYINPUT23), .A2(G128), .ZN(n1272) );
XOR2_X1 U962 ( .A(n1273), .B(n1274), .Z(n1266) );
XNOR2_X1 U963 ( .A(n1219), .B(G137), .ZN(n1274) );
XNOR2_X1 U964 ( .A(G119), .B(G125), .ZN(n1273) );
INV_X1 U965 ( .A(n1258), .ZN(n1072) );
XOR2_X1 U966 ( .A(n1275), .B(n1144), .Z(n1258) );
INV_X1 U967 ( .A(G472), .ZN(n1144) );
NAND2_X1 U968 ( .A1(n1276), .A2(n1133), .ZN(n1275) );
XOR2_X1 U969 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U970 ( .A(G101), .B(n1279), .ZN(n1278) );
NAND4_X1 U971 ( .A1(n1150), .A2(n1151), .A3(n1280), .A4(n1281), .ZN(n1279) );
NAND2_X1 U972 ( .A1(n1149), .A2(n1282), .ZN(n1281) );
INV_X1 U973 ( .A(KEYINPUT11), .ZN(n1282) );
NOR2_X1 U974 ( .A1(n1283), .A2(n1092), .ZN(n1149) );
NAND2_X1 U975 ( .A1(n1283), .A2(KEYINPUT11), .ZN(n1280) );
XNOR2_X1 U976 ( .A(n1284), .B(n1285), .ZN(n1283) );
NAND3_X1 U977 ( .A1(n1092), .A2(n1169), .A3(n1286), .ZN(n1151) );
INV_X1 U978 ( .A(n1284), .ZN(n1286) );
NAND3_X1 U979 ( .A1(n1092), .A2(n1284), .A3(n1285), .ZN(n1150) );
XOR2_X1 U980 ( .A(G113), .B(n1287), .Z(n1284) );
NOR2_X1 U981 ( .A1(KEYINPUT3), .A2(n1142), .ZN(n1277) );
NAND2_X1 U982 ( .A1(n1288), .A2(G210), .ZN(n1142) );
NOR3_X1 U983 ( .A1(n1263), .A2(n1192), .A3(n1062), .ZN(n1182) );
NAND2_X1 U984 ( .A1(n1058), .A2(n1057), .ZN(n1062) );
NAND2_X1 U985 ( .A1(n1289), .A2(n1080), .ZN(n1057) );
NAND3_X1 U986 ( .A1(n1158), .A2(n1133), .A3(n1290), .ZN(n1080) );
INV_X1 U987 ( .A(G469), .ZN(n1158) );
XOR2_X1 U988 ( .A(n1081), .B(KEYINPUT20), .Z(n1289) );
NAND2_X1 U989 ( .A1(G469), .A2(n1291), .ZN(n1081) );
NAND2_X1 U990 ( .A1(n1290), .A2(n1133), .ZN(n1291) );
XOR2_X1 U991 ( .A(n1292), .B(n1167), .Z(n1290) );
XOR2_X1 U992 ( .A(n1293), .B(n1294), .Z(n1167) );
XNOR2_X1 U993 ( .A(n1097), .B(G110), .ZN(n1294) );
NAND2_X1 U994 ( .A1(G227), .A2(n1067), .ZN(n1293) );
NAND3_X1 U995 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1292) );
NAND2_X1 U996 ( .A1(n1285), .A2(n1164), .ZN(n1297) );
INV_X1 U997 ( .A(n1168), .ZN(n1164) );
INV_X1 U998 ( .A(n1169), .ZN(n1285) );
NAND2_X1 U999 ( .A1(KEYINPUT16), .A2(n1298), .ZN(n1296) );
NAND2_X1 U1000 ( .A1(n1299), .A2(n1169), .ZN(n1298) );
XNOR2_X1 U1001 ( .A(KEYINPUT25), .B(n1168), .ZN(n1299) );
NAND2_X1 U1002 ( .A1(n1300), .A2(n1301), .ZN(n1295) );
INV_X1 U1003 ( .A(KEYINPUT16), .ZN(n1301) );
NAND2_X1 U1004 ( .A1(n1302), .A2(n1303), .ZN(n1300) );
OR2_X1 U1005 ( .A1(n1168), .A2(KEYINPUT25), .ZN(n1303) );
NAND3_X1 U1006 ( .A1(n1168), .A2(n1169), .A3(KEYINPUT25), .ZN(n1302) );
XNOR2_X1 U1007 ( .A(n1095), .B(n1304), .ZN(n1169) );
NOR2_X1 U1008 ( .A1(G131), .A2(KEYINPUT41), .ZN(n1304) );
XNOR2_X1 U1009 ( .A(G134), .B(G137), .ZN(n1095) );
XNOR2_X1 U1010 ( .A(n1305), .B(n1306), .ZN(n1168) );
XNOR2_X1 U1011 ( .A(n1092), .B(n1307), .ZN(n1306) );
XNOR2_X1 U1012 ( .A(G104), .B(KEYINPUT21), .ZN(n1305) );
NAND2_X1 U1013 ( .A1(G221), .A2(n1265), .ZN(n1058) );
NAND2_X1 U1014 ( .A1(G234), .A2(n1133), .ZN(n1265) );
AND2_X1 U1015 ( .A1(n1036), .A2(n1308), .ZN(n1192) );
NAND4_X1 U1016 ( .A1(G953), .A2(G902), .A3(n1252), .A4(n1109), .ZN(n1308) );
INV_X1 U1017 ( .A(G898), .ZN(n1109) );
NAND3_X1 U1018 ( .A1(n1252), .A2(n1067), .A3(G952), .ZN(n1036) );
NAND2_X1 U1019 ( .A1(G237), .A2(G234), .ZN(n1252) );
XOR2_X1 U1020 ( .A(n1055), .B(KEYINPUT32), .Z(n1263) );
NAND2_X1 U1021 ( .A1(n1053), .A2(n1052), .ZN(n1055) );
NAND2_X1 U1022 ( .A1(G214), .A2(n1309), .ZN(n1052) );
INV_X1 U1023 ( .A(n1236), .ZN(n1053) );
XNOR2_X1 U1024 ( .A(n1083), .B(n1310), .ZN(n1236) );
NOR2_X1 U1025 ( .A1(n1082), .A2(KEYINPUT18), .ZN(n1310) );
AND2_X1 U1026 ( .A1(n1311), .A2(n1133), .ZN(n1082) );
XNOR2_X1 U1027 ( .A(n1179), .B(n1312), .ZN(n1311) );
XNOR2_X1 U1028 ( .A(n1313), .B(n1176), .ZN(n1312) );
XNOR2_X1 U1029 ( .A(n1314), .B(n1115), .ZN(n1176) );
XNOR2_X1 U1030 ( .A(n1254), .B(n1315), .ZN(n1115) );
NOR2_X1 U1031 ( .A1(G110), .A2(KEYINPUT52), .ZN(n1315) );
XNOR2_X1 U1032 ( .A(n1117), .B(n1316), .ZN(n1314) );
NOR2_X1 U1033 ( .A1(KEYINPUT7), .A2(n1317), .ZN(n1316) );
INV_X1 U1034 ( .A(n1119), .ZN(n1317) );
XOR2_X1 U1035 ( .A(n1307), .B(n1318), .Z(n1119) );
NOR2_X1 U1036 ( .A1(G104), .A2(KEYINPUT56), .ZN(n1318) );
XOR2_X1 U1037 ( .A(G101), .B(n1319), .Z(n1307) );
XOR2_X1 U1038 ( .A(KEYINPUT38), .B(G107), .Z(n1319) );
XNOR2_X1 U1039 ( .A(n1320), .B(n1287), .ZN(n1117) );
XOR2_X1 U1040 ( .A(G116), .B(G119), .Z(n1287) );
NAND2_X1 U1041 ( .A1(KEYINPUT58), .A2(n1321), .ZN(n1320) );
NAND2_X1 U1042 ( .A1(KEYINPUT17), .A2(n1178), .ZN(n1313) );
NOR2_X1 U1043 ( .A1(n1108), .A2(G953), .ZN(n1178) );
INV_X1 U1044 ( .A(G224), .ZN(n1108) );
XNOR2_X1 U1045 ( .A(G125), .B(n1092), .ZN(n1179) );
XNOR2_X1 U1046 ( .A(G146), .B(n1322), .ZN(n1092) );
NAND2_X1 U1047 ( .A1(G210), .A2(n1309), .ZN(n1083) );
NAND2_X1 U1048 ( .A1(n1323), .A2(n1133), .ZN(n1309) );
INV_X1 U1049 ( .A(G237), .ZN(n1323) );
INV_X1 U1050 ( .A(n1054), .ZN(n1071) );
NAND2_X1 U1051 ( .A1(n1197), .A2(n1198), .ZN(n1054) );
INV_X1 U1052 ( .A(n1260), .ZN(n1198) );
XOR2_X1 U1053 ( .A(n1324), .B(n1137), .Z(n1260) );
INV_X1 U1054 ( .A(G475), .ZN(n1137) );
NAND2_X1 U1055 ( .A1(n1135), .A2(n1133), .ZN(n1324) );
XNOR2_X1 U1056 ( .A(n1325), .B(n1326), .ZN(n1135) );
XOR2_X1 U1057 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1058 ( .A(G131), .B(n1321), .ZN(n1328) );
INV_X1 U1059 ( .A(G113), .ZN(n1321) );
XNOR2_X1 U1060 ( .A(n1219), .B(G143), .ZN(n1327) );
INV_X1 U1061 ( .A(G146), .ZN(n1219) );
XOR2_X1 U1062 ( .A(n1329), .B(n1330), .Z(n1325) );
XOR2_X1 U1063 ( .A(n1331), .B(n1332), .Z(n1330) );
NAND2_X1 U1064 ( .A1(KEYINPUT59), .A2(n1254), .ZN(n1332) );
INV_X1 U1065 ( .A(G122), .ZN(n1254) );
NAND3_X1 U1066 ( .A1(n1333), .A2(n1334), .A3(n1335), .ZN(n1331) );
OR2_X1 U1067 ( .A1(n1336), .A2(KEYINPUT53), .ZN(n1335) );
NAND3_X1 U1068 ( .A1(KEYINPUT53), .A2(n1336), .A3(G140), .ZN(n1334) );
INV_X1 U1069 ( .A(G125), .ZN(n1336) );
NAND2_X1 U1070 ( .A1(n1337), .A2(n1097), .ZN(n1333) );
INV_X1 U1071 ( .A(G140), .ZN(n1097) );
NAND2_X1 U1072 ( .A1(n1338), .A2(KEYINPUT53), .ZN(n1337) );
XNOR2_X1 U1073 ( .A(G125), .B(KEYINPUT30), .ZN(n1338) );
XOR2_X1 U1074 ( .A(n1339), .B(G104), .Z(n1329) );
NAND2_X1 U1075 ( .A1(n1288), .A2(G214), .ZN(n1339) );
NOR2_X1 U1076 ( .A1(G953), .A2(G237), .ZN(n1288) );
XOR2_X1 U1077 ( .A(n1340), .B(G478), .Z(n1197) );
NAND2_X1 U1078 ( .A1(n1131), .A2(n1133), .ZN(n1340) );
INV_X1 U1079 ( .A(G902), .ZN(n1133) );
XOR2_X1 U1080 ( .A(n1341), .B(n1342), .Z(n1131) );
XOR2_X1 U1081 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1082 ( .A(n1322), .B(n1345), .ZN(n1344) );
AND4_X1 U1083 ( .A1(n1346), .A2(n1067), .A3(G234), .A4(G217), .ZN(n1345) );
INV_X1 U1084 ( .A(G953), .ZN(n1067) );
INV_X1 U1085 ( .A(KEYINPUT39), .ZN(n1346) );
XNOR2_X1 U1086 ( .A(G143), .B(n1243), .ZN(n1322) );
INV_X1 U1087 ( .A(G128), .ZN(n1243) );
XOR2_X1 U1088 ( .A(n1347), .B(G107), .Z(n1343) );
NAND2_X1 U1089 ( .A1(KEYINPUT8), .A2(G122), .ZN(n1347) );
XOR2_X1 U1090 ( .A(n1348), .B(n1349), .Z(n1341) );
XOR2_X1 U1091 ( .A(G134), .B(G116), .Z(n1349) );
XNOR2_X1 U1092 ( .A(KEYINPUT27), .B(KEYINPUT14), .ZN(n1348) );
endmodule


