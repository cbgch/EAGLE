//Key = 1111011111110110001010000010111011001001111011000111001100110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420;

XNOR2_X1 U784 ( .A(n1086), .B(n1087), .ZN(G9) );
XNOR2_X1 U785 ( .A(G107), .B(KEYINPUT23), .ZN(n1087) );
NOR2_X1 U786 ( .A1(n1088), .A2(n1089), .ZN(G75) );
XOR2_X1 U787 ( .A(n1090), .B(KEYINPUT45), .Z(n1089) );
NAND3_X1 U788 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
NOR3_X1 U789 ( .A1(n1094), .A2(n1091), .A3(n1095), .ZN(n1088) );
INV_X1 U790 ( .A(G952), .ZN(n1091) );
NAND3_X1 U791 ( .A1(n1093), .A2(n1092), .A3(n1096), .ZN(n1094) );
NAND2_X1 U792 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U793 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND4_X1 U794 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1100) );
NAND2_X1 U795 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NAND2_X1 U796 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U797 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U798 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U799 ( .A1(n1113), .A2(n1114), .ZN(n1105) );
NAND2_X1 U800 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U801 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
INV_X1 U802 ( .A(n1119), .ZN(n1115) );
NAND3_X1 U803 ( .A1(n1113), .A2(n1120), .A3(n1107), .ZN(n1099) );
NAND2_X1 U804 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND3_X1 U805 ( .A1(n1123), .A2(n1124), .A3(n1101), .ZN(n1122) );
OR2_X1 U806 ( .A1(n1104), .A2(n1102), .ZN(n1124) );
OR3_X1 U807 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1123) );
NAND2_X1 U808 ( .A1(n1128), .A2(n1102), .ZN(n1121) );
INV_X1 U809 ( .A(n1129), .ZN(n1097) );
NAND4_X1 U810 ( .A1(n1130), .A2(n1107), .A3(n1131), .A4(n1132), .ZN(n1093) );
NOR4_X1 U811 ( .A1(n1133), .A2(n1127), .A3(n1134), .A4(n1111), .ZN(n1132) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
INV_X1 U813 ( .A(n1137), .ZN(n1133) );
NOR2_X1 U814 ( .A1(n1138), .A2(n1139), .ZN(n1131) );
XNOR2_X1 U815 ( .A(KEYINPUT22), .B(n1101), .ZN(n1139) );
XNOR2_X1 U816 ( .A(G472), .B(n1140), .ZN(n1138) );
XOR2_X1 U817 ( .A(n1141), .B(n1142), .Z(G72) );
NOR2_X1 U818 ( .A1(n1143), .A2(n1092), .ZN(n1142) );
AND2_X1 U819 ( .A1(G227), .A2(G900), .ZN(n1143) );
NAND2_X1 U820 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
NAND3_X1 U821 ( .A1(n1146), .A2(n1092), .A3(n1147), .ZN(n1145) );
NAND3_X1 U822 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1144) );
INV_X1 U823 ( .A(n1147), .ZN(n1150) );
NAND2_X1 U824 ( .A1(n1151), .A2(n1152), .ZN(n1147) );
NAND3_X1 U825 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1152) );
XOR2_X1 U826 ( .A(n1156), .B(n1157), .Z(n1155) );
OR2_X1 U827 ( .A1(n1158), .A2(KEYINPUT42), .ZN(n1154) );
NAND2_X1 U828 ( .A1(KEYINPUT42), .A2(n1159), .ZN(n1153) );
XOR2_X1 U829 ( .A(n1160), .B(KEYINPUT46), .Z(n1151) );
NAND3_X1 U830 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1160) );
XNOR2_X1 U831 ( .A(n1156), .B(n1157), .ZN(n1163) );
NAND2_X1 U832 ( .A1(KEYINPUT51), .A2(n1164), .ZN(n1156) );
XNOR2_X1 U833 ( .A(KEYINPUT42), .B(n1158), .ZN(n1161) );
NAND2_X1 U834 ( .A1(G953), .A2(n1165), .ZN(n1149) );
XNOR2_X1 U835 ( .A(n1166), .B(KEYINPUT33), .ZN(n1148) );
XOR2_X1 U836 ( .A(n1167), .B(n1168), .Z(G69) );
NAND2_X1 U837 ( .A1(G953), .A2(n1169), .ZN(n1168) );
NAND2_X1 U838 ( .A1(G898), .A2(G224), .ZN(n1169) );
NAND2_X1 U839 ( .A1(KEYINPUT6), .A2(n1170), .ZN(n1167) );
XOR2_X1 U840 ( .A(n1171), .B(n1172), .Z(n1170) );
NAND2_X1 U841 ( .A1(n1092), .A2(n1173), .ZN(n1172) );
NAND2_X1 U842 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NAND2_X1 U843 ( .A1(n1176), .A2(n1177), .ZN(n1171) );
NAND2_X1 U844 ( .A1(G953), .A2(n1178), .ZN(n1177) );
XOR2_X1 U845 ( .A(n1179), .B(n1180), .Z(n1176) );
NAND3_X1 U846 ( .A1(n1181), .A2(n1182), .A3(KEYINPUT63), .ZN(n1179) );
NAND2_X1 U847 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
INV_X1 U848 ( .A(KEYINPUT32), .ZN(n1184) );
NAND2_X1 U849 ( .A1(n1185), .A2(n1186), .ZN(n1183) );
NAND2_X1 U850 ( .A1(KEYINPUT32), .A2(n1187), .ZN(n1181) );
NOR2_X1 U851 ( .A1(n1188), .A2(n1189), .ZN(G66) );
XNOR2_X1 U852 ( .A(n1190), .B(n1191), .ZN(n1189) );
NOR2_X1 U853 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NOR2_X1 U854 ( .A1(n1188), .A2(n1194), .ZN(G63) );
XOR2_X1 U855 ( .A(n1195), .B(n1196), .Z(n1194) );
NAND3_X1 U856 ( .A1(n1197), .A2(G478), .A3(KEYINPUT29), .ZN(n1195) );
NOR2_X1 U857 ( .A1(n1188), .A2(n1198), .ZN(G60) );
XOR2_X1 U858 ( .A(n1199), .B(n1200), .Z(n1198) );
AND2_X1 U859 ( .A1(G475), .A2(n1197), .ZN(n1199) );
XOR2_X1 U860 ( .A(n1201), .B(n1202), .Z(G6) );
NAND2_X1 U861 ( .A1(KEYINPUT2), .A2(G104), .ZN(n1202) );
NOR2_X1 U862 ( .A1(n1188), .A2(n1203), .ZN(G57) );
XOR2_X1 U863 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U864 ( .A(KEYINPUT53), .B(n1206), .Z(n1205) );
NOR2_X1 U865 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NOR2_X1 U866 ( .A1(G101), .A2(n1209), .ZN(n1207) );
XNOR2_X1 U867 ( .A(KEYINPUT12), .B(n1210), .ZN(n1209) );
XOR2_X1 U868 ( .A(n1211), .B(n1212), .Z(n1204) );
AND2_X1 U869 ( .A1(G472), .A2(n1197), .ZN(n1212) );
NAND2_X1 U870 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
NOR2_X1 U871 ( .A1(n1188), .A2(n1215), .ZN(G54) );
XOR2_X1 U872 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U873 ( .A(n1218), .B(n1219), .Z(n1217) );
NAND2_X1 U874 ( .A1(KEYINPUT20), .A2(n1220), .ZN(n1218) );
XNOR2_X1 U875 ( .A(n1221), .B(n1222), .ZN(n1216) );
AND2_X1 U876 ( .A1(G469), .A2(n1197), .ZN(n1222) );
INV_X1 U877 ( .A(n1193), .ZN(n1197) );
NOR2_X1 U878 ( .A1(n1188), .A2(n1223), .ZN(G51) );
XOR2_X1 U879 ( .A(n1224), .B(n1225), .Z(n1223) );
NOR2_X1 U880 ( .A1(n1226), .A2(n1193), .ZN(n1225) );
NAND2_X1 U881 ( .A1(G902), .A2(n1095), .ZN(n1193) );
NAND3_X1 U882 ( .A1(n1174), .A2(n1227), .A3(n1166), .ZN(n1095) );
INV_X1 U883 ( .A(n1146), .ZN(n1166) );
NAND4_X1 U884 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1146) );
NOR4_X1 U885 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1231) );
INV_X1 U886 ( .A(n1236), .ZN(n1235) );
NOR2_X1 U887 ( .A1(n1237), .A2(n1238), .ZN(n1230) );
XNOR2_X1 U888 ( .A(KEYINPUT59), .B(n1175), .ZN(n1227) );
AND4_X1 U889 ( .A1(n1201), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1174) );
NOR4_X1 U890 ( .A1(n1086), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1241) );
INV_X1 U891 ( .A(n1245), .ZN(n1242) );
AND3_X1 U892 ( .A1(n1113), .A2(n1246), .A3(n1126), .ZN(n1086) );
NAND3_X1 U893 ( .A1(n1247), .A2(n1125), .A3(n1248), .ZN(n1240) );
NAND3_X1 U894 ( .A1(n1246), .A2(n1125), .A3(n1113), .ZN(n1201) );
NAND3_X1 U895 ( .A1(n1249), .A2(n1250), .A3(KEYINPUT10), .ZN(n1224) );
OR2_X1 U896 ( .A1(n1251), .A2(n1252), .ZN(n1249) );
NOR2_X1 U897 ( .A1(n1092), .A2(G952), .ZN(n1188) );
XOR2_X1 U898 ( .A(n1253), .B(n1238), .Z(G48) );
AND3_X1 U899 ( .A1(n1119), .A2(n1125), .A3(n1254), .ZN(n1238) );
XNOR2_X1 U900 ( .A(G146), .B(KEYINPUT50), .ZN(n1253) );
NAND3_X1 U901 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(G45) );
NAND2_X1 U902 ( .A1(KEYINPUT21), .A2(G143), .ZN(n1257) );
OR3_X1 U903 ( .A1(G143), .A2(KEYINPUT21), .A3(n1236), .ZN(n1256) );
NAND2_X1 U904 ( .A1(n1258), .A2(n1236), .ZN(n1255) );
NAND3_X1 U905 ( .A1(n1259), .A2(n1119), .A3(n1260), .ZN(n1236) );
NAND2_X1 U906 ( .A1(n1261), .A2(n1262), .ZN(n1258) );
INV_X1 U907 ( .A(KEYINPUT21), .ZN(n1262) );
XOR2_X1 U908 ( .A(KEYINPUT36), .B(G143), .Z(n1261) );
XOR2_X1 U909 ( .A(G140), .B(n1234), .Z(G42) );
AND3_X1 U910 ( .A1(n1107), .A2(n1128), .A3(n1263), .ZN(n1234) );
XOR2_X1 U911 ( .A(n1264), .B(n1237), .Z(G39) );
AND3_X1 U912 ( .A1(n1107), .A2(n1102), .A3(n1254), .ZN(n1237) );
XNOR2_X1 U913 ( .A(G137), .B(KEYINPUT62), .ZN(n1264) );
XOR2_X1 U914 ( .A(G134), .B(n1233), .Z(G36) );
AND3_X1 U915 ( .A1(n1107), .A2(n1126), .A3(n1260), .ZN(n1233) );
XOR2_X1 U916 ( .A(G131), .B(n1232), .Z(G33) );
AND3_X1 U917 ( .A1(n1107), .A2(n1125), .A3(n1260), .ZN(n1232) );
AND3_X1 U918 ( .A1(n1128), .A2(n1265), .A3(n1247), .ZN(n1260) );
NOR2_X1 U919 ( .A1(n1266), .A2(n1117), .ZN(n1107) );
XNOR2_X1 U920 ( .A(n1228), .B(n1267), .ZN(G30) );
NOR2_X1 U921 ( .A1(KEYINPUT25), .A2(n1268), .ZN(n1267) );
NAND3_X1 U922 ( .A1(n1126), .A2(n1119), .A3(n1254), .ZN(n1228) );
AND4_X1 U923 ( .A1(n1269), .A2(n1128), .A3(n1111), .A4(n1265), .ZN(n1254) );
XNOR2_X1 U924 ( .A(G101), .B(n1175), .ZN(G3) );
NAND3_X1 U925 ( .A1(n1246), .A2(n1102), .A3(n1247), .ZN(n1175) );
XNOR2_X1 U926 ( .A(G125), .B(n1229), .ZN(G27) );
NAND4_X1 U927 ( .A1(n1101), .A2(n1263), .A3(n1119), .A4(n1104), .ZN(n1229) );
AND4_X1 U928 ( .A1(n1125), .A2(n1111), .A3(n1265), .A4(n1112), .ZN(n1263) );
NAND2_X1 U929 ( .A1(n1129), .A2(n1270), .ZN(n1265) );
NAND4_X1 U930 ( .A1(G902), .A2(G953), .A3(n1271), .A4(n1165), .ZN(n1270) );
INV_X1 U931 ( .A(G900), .ZN(n1165) );
XOR2_X1 U932 ( .A(n1272), .B(n1273), .Z(G24) );
XOR2_X1 U933 ( .A(KEYINPUT17), .B(G122), .Z(n1273) );
NAND2_X1 U934 ( .A1(n1274), .A2(n1275), .ZN(n1272) );
OR2_X1 U935 ( .A1(n1239), .A2(KEYINPUT4), .ZN(n1275) );
NAND3_X1 U936 ( .A1(n1259), .A2(n1113), .A3(n1248), .ZN(n1239) );
NAND4_X1 U937 ( .A1(n1113), .A2(n1276), .A3(n1248), .A4(KEYINPUT4), .ZN(n1274) );
NOR2_X1 U938 ( .A1(n1111), .A2(n1269), .ZN(n1113) );
NAND2_X1 U939 ( .A1(n1277), .A2(n1278), .ZN(G21) );
NAND2_X1 U940 ( .A1(n1244), .A2(n1279), .ZN(n1278) );
INV_X1 U941 ( .A(n1280), .ZN(n1244) );
XOR2_X1 U942 ( .A(n1281), .B(KEYINPUT15), .Z(n1277) );
NAND2_X1 U943 ( .A1(G119), .A2(n1280), .ZN(n1281) );
NAND4_X1 U944 ( .A1(n1248), .A2(n1269), .A3(n1102), .A4(n1111), .ZN(n1280) );
INV_X1 U945 ( .A(n1112), .ZN(n1269) );
XNOR2_X1 U946 ( .A(n1282), .B(n1243), .ZN(G18) );
AND3_X1 U947 ( .A1(n1247), .A2(n1126), .A3(n1248), .ZN(n1243) );
INV_X1 U948 ( .A(n1283), .ZN(n1248) );
XOR2_X1 U949 ( .A(G113), .B(n1284), .Z(G15) );
NOR4_X1 U950 ( .A1(KEYINPUT52), .A2(n1285), .A3(n1109), .A4(n1283), .ZN(n1284) );
NAND3_X1 U951 ( .A1(n1286), .A2(n1104), .A3(n1101), .ZN(n1283) );
INV_X1 U952 ( .A(n1247), .ZN(n1109) );
NOR2_X1 U953 ( .A1(n1112), .A2(n1111), .ZN(n1247) );
INV_X1 U954 ( .A(n1125), .ZN(n1285) );
NAND2_X1 U955 ( .A1(n1287), .A2(n1288), .ZN(n1125) );
NAND3_X1 U956 ( .A1(n1130), .A2(n1289), .A3(n1290), .ZN(n1288) );
INV_X1 U957 ( .A(KEYINPUT43), .ZN(n1290) );
NAND2_X1 U958 ( .A1(KEYINPUT43), .A2(n1259), .ZN(n1287) );
INV_X1 U959 ( .A(n1276), .ZN(n1259) );
NAND2_X1 U960 ( .A1(n1291), .A2(n1289), .ZN(n1276) );
XNOR2_X1 U961 ( .A(G110), .B(n1245), .ZN(G12) );
NAND4_X1 U962 ( .A1(n1246), .A2(n1102), .A3(n1111), .A4(n1112), .ZN(n1245) );
NAND3_X1 U963 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n1112) );
NAND2_X1 U964 ( .A1(KEYINPUT48), .A2(G472), .ZN(n1294) );
NAND3_X1 U965 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1293) );
INV_X1 U966 ( .A(KEYINPUT48), .ZN(n1296) );
OR2_X1 U967 ( .A1(n1297), .A2(n1295), .ZN(n1292) );
NOR2_X1 U968 ( .A1(G472), .A2(KEYINPUT37), .ZN(n1295) );
XNOR2_X1 U969 ( .A(n1140), .B(KEYINPUT44), .ZN(n1297) );
NAND2_X1 U970 ( .A1(n1298), .A2(n1299), .ZN(n1140) );
NAND2_X1 U971 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NAND3_X1 U972 ( .A1(n1302), .A2(n1214), .A3(n1303), .ZN(n1301) );
XNOR2_X1 U973 ( .A(n1304), .B(KEYINPUT57), .ZN(n1303) );
XOR2_X1 U974 ( .A(KEYINPUT40), .B(n1305), .Z(n1302) );
NAND3_X1 U975 ( .A1(n1306), .A2(n1307), .A3(n1305), .ZN(n1300) );
NOR2_X1 U976 ( .A1(n1308), .A2(n1208), .ZN(n1305) );
NOR2_X1 U977 ( .A1(n1309), .A2(n1210), .ZN(n1208) );
INV_X1 U978 ( .A(G101), .ZN(n1309) );
XNOR2_X1 U979 ( .A(n1310), .B(KEYINPUT31), .ZN(n1308) );
NAND2_X1 U980 ( .A1(n1311), .A2(n1210), .ZN(n1310) );
NAND3_X1 U981 ( .A1(G210), .A2(n1312), .A3(n1313), .ZN(n1210) );
XNOR2_X1 U982 ( .A(G953), .B(KEYINPUT24), .ZN(n1313) );
XNOR2_X1 U983 ( .A(G101), .B(KEYINPUT35), .ZN(n1311) );
NAND3_X1 U984 ( .A1(n1214), .A2(n1213), .A3(n1314), .ZN(n1307) );
INV_X1 U985 ( .A(KEYINPUT57), .ZN(n1314) );
INV_X1 U986 ( .A(n1304), .ZN(n1213) );
NAND2_X1 U987 ( .A1(n1315), .A2(n1316), .ZN(n1214) );
NAND2_X1 U988 ( .A1(n1304), .A2(KEYINPUT57), .ZN(n1306) );
NOR2_X1 U989 ( .A1(n1316), .A2(n1315), .ZN(n1304) );
XNOR2_X1 U990 ( .A(n1317), .B(n1220), .ZN(n1315) );
NAND3_X1 U991 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1316) );
NAND2_X1 U992 ( .A1(n1321), .A2(G113), .ZN(n1320) );
OR3_X1 U993 ( .A1(n1282), .A2(G113), .A3(n1279), .ZN(n1319) );
NAND2_X1 U994 ( .A1(n1322), .A2(n1279), .ZN(n1318) );
XNOR2_X1 U995 ( .A(G113), .B(G116), .ZN(n1322) );
XOR2_X1 U996 ( .A(n1323), .B(n1192), .Z(n1111) );
NAND2_X1 U997 ( .A1(G217), .A2(n1324), .ZN(n1192) );
NAND2_X1 U998 ( .A1(n1190), .A2(n1298), .ZN(n1323) );
XNOR2_X1 U999 ( .A(n1325), .B(n1326), .ZN(n1190) );
XNOR2_X1 U1000 ( .A(n1327), .B(n1328), .ZN(n1326) );
NOR2_X1 U1001 ( .A1(KEYINPUT60), .A2(n1329), .ZN(n1328) );
XNOR2_X1 U1002 ( .A(G146), .B(n1330), .ZN(n1329) );
NAND2_X1 U1003 ( .A1(n1331), .A2(KEYINPUT61), .ZN(n1327) );
XOR2_X1 U1004 ( .A(n1332), .B(n1333), .Z(n1331) );
AND3_X1 U1005 ( .A1(G221), .A2(n1092), .A3(G234), .ZN(n1333) );
NAND2_X1 U1006 ( .A1(KEYINPUT18), .A2(n1334), .ZN(n1332) );
INV_X1 U1007 ( .A(G137), .ZN(n1334) );
XNOR2_X1 U1008 ( .A(G110), .B(n1335), .ZN(n1325) );
XNOR2_X1 U1009 ( .A(n1268), .B(G119), .ZN(n1335) );
NAND2_X1 U1010 ( .A1(n1336), .A2(n1337), .ZN(n1102) );
OR3_X1 U1011 ( .A1(n1289), .A2(n1291), .A3(KEYINPUT43), .ZN(n1337) );
NAND2_X1 U1012 ( .A1(KEYINPUT43), .A2(n1126), .ZN(n1336) );
NOR2_X1 U1013 ( .A1(n1289), .A2(n1130), .ZN(n1126) );
INV_X1 U1014 ( .A(n1291), .ZN(n1130) );
XNOR2_X1 U1015 ( .A(n1338), .B(G478), .ZN(n1291) );
NAND2_X1 U1016 ( .A1(n1196), .A2(n1298), .ZN(n1338) );
XNOR2_X1 U1017 ( .A(n1339), .B(n1340), .ZN(n1196) );
XNOR2_X1 U1018 ( .A(n1341), .B(n1342), .ZN(n1340) );
NAND2_X1 U1019 ( .A1(KEYINPUT39), .A2(n1268), .ZN(n1341) );
INV_X1 U1020 ( .A(G128), .ZN(n1268) );
XOR2_X1 U1021 ( .A(n1343), .B(n1344), .Z(n1339) );
XOR2_X1 U1022 ( .A(G143), .B(n1345), .Z(n1344) );
NOR2_X1 U1023 ( .A1(KEYINPUT16), .A2(n1346), .ZN(n1345) );
XNOR2_X1 U1024 ( .A(G107), .B(n1347), .ZN(n1346) );
NAND2_X1 U1025 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
XOR2_X1 U1026 ( .A(n1350), .B(G122), .Z(n1349) );
NAND2_X1 U1027 ( .A1(KEYINPUT11), .A2(n1282), .ZN(n1350) );
INV_X1 U1028 ( .A(G116), .ZN(n1282) );
XNOR2_X1 U1029 ( .A(KEYINPUT7), .B(KEYINPUT41), .ZN(n1348) );
NAND3_X1 U1030 ( .A1(G217), .A2(n1092), .A3(G234), .ZN(n1343) );
NAND3_X1 U1031 ( .A1(n1351), .A2(n1352), .A3(n1137), .ZN(n1289) );
NAND2_X1 U1032 ( .A1(n1135), .A2(n1136), .ZN(n1137) );
NAND2_X1 U1033 ( .A1(n1135), .A2(n1353), .ZN(n1352) );
OR3_X1 U1034 ( .A1(n1136), .A2(n1135), .A3(n1353), .ZN(n1351) );
INV_X1 U1035 ( .A(KEYINPUT54), .ZN(n1353) );
NOR2_X1 U1036 ( .A1(n1200), .A2(G902), .ZN(n1135) );
XNOR2_X1 U1037 ( .A(n1354), .B(n1355), .ZN(n1200) );
NOR2_X1 U1038 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
XOR2_X1 U1039 ( .A(KEYINPUT19), .B(n1358), .Z(n1357) );
AND2_X1 U1040 ( .A1(n1359), .A2(G104), .ZN(n1358) );
NOR2_X1 U1041 ( .A1(G104), .A2(n1359), .ZN(n1356) );
XOR2_X1 U1042 ( .A(G122), .B(G113), .Z(n1359) );
NAND2_X1 U1043 ( .A1(KEYINPUT30), .A2(n1360), .ZN(n1354) );
XOR2_X1 U1044 ( .A(n1361), .B(n1362), .Z(n1360) );
XOR2_X1 U1045 ( .A(n1363), .B(n1364), .Z(n1362) );
NOR3_X1 U1046 ( .A1(n1365), .A2(G953), .A3(n1366), .ZN(n1364) );
XNOR2_X1 U1047 ( .A(G237), .B(KEYINPUT55), .ZN(n1366) );
INV_X1 U1048 ( .A(G214), .ZN(n1365) );
NAND3_X1 U1049 ( .A1(n1367), .A2(n1368), .A3(KEYINPUT5), .ZN(n1363) );
NAND3_X1 U1050 ( .A1(n1369), .A2(n1370), .A3(n1371), .ZN(n1368) );
XNOR2_X1 U1051 ( .A(KEYINPUT34), .B(G146), .ZN(n1371) );
NAND2_X1 U1052 ( .A1(n1159), .A2(n1372), .ZN(n1370) );
INV_X1 U1053 ( .A(n1330), .ZN(n1159) );
NAND2_X1 U1054 ( .A1(KEYINPUT27), .A2(n1373), .ZN(n1369) );
NAND3_X1 U1055 ( .A1(n1374), .A2(n1375), .A3(n1376), .ZN(n1367) );
XNOR2_X1 U1056 ( .A(KEYINPUT34), .B(n1377), .ZN(n1376) );
NAND2_X1 U1057 ( .A1(KEYINPUT27), .A2(n1162), .ZN(n1375) );
NAND2_X1 U1058 ( .A1(n1330), .A2(n1372), .ZN(n1374) );
INV_X1 U1059 ( .A(KEYINPUT27), .ZN(n1372) );
NAND2_X1 U1060 ( .A1(n1162), .A2(n1158), .ZN(n1330) );
NAND2_X1 U1061 ( .A1(G140), .A2(n1378), .ZN(n1158) );
INV_X1 U1062 ( .A(n1373), .ZN(n1162) );
NOR2_X1 U1063 ( .A1(n1378), .A2(G140), .ZN(n1373) );
XNOR2_X1 U1064 ( .A(G131), .B(n1379), .ZN(n1361) );
XOR2_X1 U1065 ( .A(KEYINPUT38), .B(G143), .Z(n1379) );
XOR2_X1 U1066 ( .A(G475), .B(KEYINPUT26), .Z(n1136) );
AND2_X1 U1067 ( .A1(n1286), .A2(n1128), .ZN(n1246) );
NOR2_X1 U1068 ( .A1(n1101), .A2(n1127), .ZN(n1128) );
INV_X1 U1069 ( .A(n1104), .ZN(n1127) );
NAND2_X1 U1070 ( .A1(G221), .A2(n1324), .ZN(n1104) );
NAND2_X1 U1071 ( .A1(G234), .A2(n1298), .ZN(n1324) );
XOR2_X1 U1072 ( .A(n1380), .B(G469), .Z(n1101) );
NAND4_X1 U1073 ( .A1(n1381), .A2(n1298), .A3(n1382), .A4(n1383), .ZN(n1380) );
NAND4_X1 U1074 ( .A1(n1384), .A2(KEYINPUT58), .A3(KEYINPUT3), .A4(n1385), .ZN(n1383) );
XNOR2_X1 U1075 ( .A(n1221), .B(n1164), .ZN(n1384) );
INV_X1 U1076 ( .A(n1220), .ZN(n1164) );
OR2_X1 U1077 ( .A1(n1385), .A2(KEYINPUT3), .ZN(n1382) );
NAND2_X1 U1078 ( .A1(n1386), .A2(n1387), .ZN(n1381) );
NAND2_X1 U1079 ( .A1(KEYINPUT58), .A2(n1385), .ZN(n1387) );
XOR2_X1 U1080 ( .A(n1219), .B(KEYINPUT49), .Z(n1385) );
XOR2_X1 U1081 ( .A(n1388), .B(n1389), .Z(n1219) );
XNOR2_X1 U1082 ( .A(G140), .B(n1390), .ZN(n1389) );
NAND2_X1 U1083 ( .A1(G227), .A2(n1092), .ZN(n1388) );
XNOR2_X1 U1084 ( .A(n1221), .B(n1220), .ZN(n1386) );
XOR2_X1 U1085 ( .A(n1391), .B(n1392), .Z(n1220) );
INV_X1 U1086 ( .A(n1342), .ZN(n1392) );
XOR2_X1 U1087 ( .A(G134), .B(KEYINPUT47), .Z(n1342) );
XNOR2_X1 U1088 ( .A(G131), .B(G137), .ZN(n1391) );
NAND2_X1 U1089 ( .A1(n1393), .A2(n1394), .ZN(n1221) );
NAND2_X1 U1090 ( .A1(n1395), .A2(n1396), .ZN(n1394) );
XNOR2_X1 U1091 ( .A(G107), .B(n1397), .ZN(n1396) );
NAND2_X1 U1092 ( .A1(n1398), .A2(n1399), .ZN(n1393) );
XOR2_X1 U1093 ( .A(KEYINPUT0), .B(n1395), .Z(n1399) );
XNOR2_X1 U1094 ( .A(n1157), .B(G101), .ZN(n1395) );
NAND2_X1 U1095 ( .A1(n1400), .A2(n1401), .ZN(n1157) );
NAND2_X1 U1096 ( .A1(n1402), .A2(G146), .ZN(n1401) );
NAND2_X1 U1097 ( .A1(n1403), .A2(n1377), .ZN(n1400) );
XNOR2_X1 U1098 ( .A(n1402), .B(KEYINPUT56), .ZN(n1403) );
XOR2_X1 U1099 ( .A(n1397), .B(G107), .Z(n1398) );
NAND2_X1 U1100 ( .A1(KEYINPUT9), .A2(n1404), .ZN(n1397) );
INV_X1 U1101 ( .A(G104), .ZN(n1404) );
AND2_X1 U1102 ( .A1(n1119), .A2(n1405), .ZN(n1286) );
NAND2_X1 U1103 ( .A1(n1129), .A2(n1406), .ZN(n1405) );
NAND4_X1 U1104 ( .A1(G902), .A2(G953), .A3(n1271), .A4(n1178), .ZN(n1406) );
INV_X1 U1105 ( .A(G898), .ZN(n1178) );
NAND3_X1 U1106 ( .A1(n1271), .A2(n1092), .A3(G952), .ZN(n1129) );
NAND2_X1 U1107 ( .A1(G234), .A2(G237), .ZN(n1271) );
NOR2_X1 U1108 ( .A1(n1118), .A2(n1117), .ZN(n1119) );
AND2_X1 U1109 ( .A1(G214), .A2(n1407), .ZN(n1117) );
INV_X1 U1110 ( .A(n1266), .ZN(n1118) );
XOR2_X1 U1111 ( .A(n1408), .B(n1226), .Z(n1266) );
NAND2_X1 U1112 ( .A1(G210), .A2(n1407), .ZN(n1226) );
NAND2_X1 U1113 ( .A1(n1298), .A2(n1312), .ZN(n1407) );
INV_X1 U1114 ( .A(G237), .ZN(n1312) );
NAND2_X1 U1115 ( .A1(n1409), .A2(n1298), .ZN(n1408) );
INV_X1 U1116 ( .A(G902), .ZN(n1298) );
XOR2_X1 U1117 ( .A(n1410), .B(KEYINPUT8), .Z(n1409) );
NAND2_X1 U1118 ( .A1(n1411), .A2(n1250), .ZN(n1410) );
NAND2_X1 U1119 ( .A1(n1252), .A2(n1251), .ZN(n1250) );
XOR2_X1 U1120 ( .A(KEYINPUT28), .B(n1412), .Z(n1411) );
NOR2_X1 U1121 ( .A1(n1252), .A2(n1251), .ZN(n1412) );
XNOR2_X1 U1122 ( .A(n1413), .B(n1414), .ZN(n1251) );
XNOR2_X1 U1123 ( .A(KEYINPUT1), .B(n1378), .ZN(n1414) );
INV_X1 U1124 ( .A(G125), .ZN(n1378) );
XNOR2_X1 U1125 ( .A(n1317), .B(n1415), .ZN(n1413) );
AND2_X1 U1126 ( .A1(n1092), .A2(G224), .ZN(n1415) );
INV_X1 U1127 ( .A(G953), .ZN(n1092) );
XNOR2_X1 U1128 ( .A(n1377), .B(n1402), .ZN(n1317) );
XOR2_X1 U1129 ( .A(G128), .B(G143), .Z(n1402) );
INV_X1 U1130 ( .A(G146), .ZN(n1377) );
XOR2_X1 U1131 ( .A(n1187), .B(n1180), .Z(n1252) );
XNOR2_X1 U1132 ( .A(n1390), .B(G122), .ZN(n1180) );
INV_X1 U1133 ( .A(G110), .ZN(n1390) );
XNOR2_X1 U1134 ( .A(n1185), .B(n1186), .ZN(n1187) );
XOR2_X1 U1135 ( .A(n1416), .B(n1417), .Z(n1186) );
XOR2_X1 U1136 ( .A(KEYINPUT14), .B(G107), .Z(n1417) );
XNOR2_X1 U1137 ( .A(G104), .B(G101), .ZN(n1416) );
XOR2_X1 U1138 ( .A(n1418), .B(G113), .Z(n1185) );
NAND2_X1 U1139 ( .A1(n1419), .A2(n1420), .ZN(n1418) );
NAND2_X1 U1140 ( .A1(G116), .A2(n1279), .ZN(n1420) );
XOR2_X1 U1141 ( .A(KEYINPUT13), .B(n1321), .Z(n1419) );
NOR2_X1 U1142 ( .A1(n1279), .A2(G116), .ZN(n1321) );
INV_X1 U1143 ( .A(G119), .ZN(n1279) );
endmodule


