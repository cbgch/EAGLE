//Key = 0000110110011100110110011001111111111010001110110100000001110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;

XNOR2_X1 U787 ( .A(G107), .B(n1093), .ZN(G9) );
NOR2_X1 U788 ( .A1(n1094), .A2(n1095), .ZN(G75) );
XOR2_X1 U789 ( .A(n1096), .B(KEYINPUT34), .Z(n1095) );
NAND4_X1 U790 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
NOR4_X1 U791 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1100) );
INV_X1 U792 ( .A(G952), .ZN(n1103) );
NOR2_X1 U793 ( .A1(n1105), .A2(n1106), .ZN(n1102) );
NOR3_X1 U794 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1101) );
NOR2_X1 U795 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NOR2_X1 U796 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NOR2_X1 U797 ( .A1(n1114), .A2(n1115), .ZN(n1110) );
NOR2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
AND2_X1 U799 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U800 ( .A1(n1120), .A2(n1121), .ZN(n1116) );
NOR2_X1 U801 ( .A1(n1122), .A2(n1123), .ZN(n1099) );
XOR2_X1 U802 ( .A(KEYINPUT43), .B(n1124), .Z(n1123) );
NOR2_X1 U803 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR2_X1 U804 ( .A1(n1127), .A2(n1106), .ZN(n1126) );
OR3_X1 U805 ( .A1(n1113), .A2(n1115), .A3(n1107), .ZN(n1106) );
INV_X1 U806 ( .A(n1128), .ZN(n1127) );
NOR3_X1 U807 ( .A1(n1107), .A2(n1129), .A3(n1109), .ZN(n1125) );
NOR2_X1 U808 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U809 ( .A1(n1132), .A2(n1115), .ZN(n1131) );
INV_X1 U810 ( .A(n1133), .ZN(n1115) );
NOR2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
AND2_X1 U812 ( .A1(n1136), .A2(n1119), .ZN(n1135) );
NOR3_X1 U813 ( .A1(n1137), .A2(n1121), .A3(n1138), .ZN(n1134) );
INV_X1 U814 ( .A(n1139), .ZN(n1121) );
NOR3_X1 U815 ( .A1(n1140), .A2(n1141), .A3(n1113), .ZN(n1130) );
NAND2_X1 U816 ( .A1(n1119), .A2(n1139), .ZN(n1113) );
NOR2_X1 U817 ( .A1(n1142), .A2(n1104), .ZN(n1094) );
NAND2_X1 U818 ( .A1(n1143), .A2(n1144), .ZN(n1104) );
NAND4_X1 U819 ( .A1(n1145), .A2(n1133), .A3(n1146), .A4(n1147), .ZN(n1144) );
NOR4_X1 U820 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1147) );
NOR2_X1 U821 ( .A1(n1152), .A2(n1153), .ZN(n1150) );
XNOR2_X1 U822 ( .A(G472), .B(KEYINPUT54), .ZN(n1153) );
INV_X1 U823 ( .A(n1154), .ZN(n1152) );
XNOR2_X1 U824 ( .A(G952), .B(KEYINPUT23), .ZN(n1142) );
XOR2_X1 U825 ( .A(n1155), .B(n1156), .Z(G72) );
XOR2_X1 U826 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U827 ( .A1(n1159), .A2(n1143), .ZN(n1158) );
AND2_X1 U828 ( .A1(G227), .A2(G900), .ZN(n1159) );
NAND2_X1 U829 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NAND2_X1 U830 ( .A1(G953), .A2(n1162), .ZN(n1161) );
XOR2_X1 U831 ( .A(n1163), .B(n1164), .Z(n1160) );
XOR2_X1 U832 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND2_X1 U833 ( .A1(KEYINPUT42), .A2(n1167), .ZN(n1165) );
XNOR2_X1 U834 ( .A(n1168), .B(n1169), .ZN(n1167) );
XNOR2_X1 U835 ( .A(n1170), .B(n1171), .ZN(n1169) );
NAND2_X1 U836 ( .A1(KEYINPUT5), .A2(G137), .ZN(n1170) );
XOR2_X1 U837 ( .A(n1172), .B(n1173), .Z(n1163) );
XNOR2_X1 U838 ( .A(G140), .B(KEYINPUT41), .ZN(n1173) );
NAND2_X1 U839 ( .A1(KEYINPUT28), .A2(n1174), .ZN(n1172) );
NAND2_X1 U840 ( .A1(n1143), .A2(n1122), .ZN(n1155) );
NAND2_X1 U841 ( .A1(n1175), .A2(n1176), .ZN(G69) );
NAND2_X1 U842 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NAND2_X1 U843 ( .A1(G953), .A2(n1179), .ZN(n1178) );
NAND3_X1 U844 ( .A1(G953), .A2(n1180), .A3(n1181), .ZN(n1175) );
INV_X1 U845 ( .A(n1177), .ZN(n1181) );
XNOR2_X1 U846 ( .A(n1182), .B(n1183), .ZN(n1177) );
NOR2_X1 U847 ( .A1(n1184), .A2(G953), .ZN(n1183) );
AND3_X1 U848 ( .A1(n1098), .A2(n1185), .A3(n1186), .ZN(n1184) );
NAND4_X1 U849 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1182) );
NAND3_X1 U850 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1190) );
NAND2_X1 U851 ( .A1(n1194), .A2(n1195), .ZN(n1189) );
XNOR2_X1 U852 ( .A(n1192), .B(n1196), .ZN(n1194) );
NAND2_X1 U853 ( .A1(KEYINPUT44), .A2(n1197), .ZN(n1192) );
NAND2_X1 U854 ( .A1(KEYINPUT44), .A2(n1198), .ZN(n1188) );
INV_X1 U855 ( .A(n1199), .ZN(n1198) );
NAND2_X1 U856 ( .A1(G953), .A2(n1200), .ZN(n1187) );
NAND2_X1 U857 ( .A1(G898), .A2(G224), .ZN(n1180) );
NOR2_X1 U858 ( .A1(n1201), .A2(n1202), .ZN(G66) );
XNOR2_X1 U859 ( .A(n1203), .B(n1204), .ZN(n1202) );
NOR2_X1 U860 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NOR2_X1 U861 ( .A1(n1201), .A2(n1207), .ZN(G63) );
XOR2_X1 U862 ( .A(n1208), .B(n1209), .Z(n1207) );
XNOR2_X1 U863 ( .A(KEYINPUT62), .B(n1210), .ZN(n1208) );
NOR3_X1 U864 ( .A1(n1206), .A2(KEYINPUT55), .A3(n1211), .ZN(n1210) );
NOR2_X1 U865 ( .A1(n1201), .A2(n1212), .ZN(G60) );
XNOR2_X1 U866 ( .A(n1213), .B(n1214), .ZN(n1212) );
AND2_X1 U867 ( .A1(G475), .A2(n1215), .ZN(n1214) );
XNOR2_X1 U868 ( .A(G104), .B(n1185), .ZN(G6) );
NOR2_X1 U869 ( .A1(n1201), .A2(n1216), .ZN(G57) );
XOR2_X1 U870 ( .A(n1217), .B(n1218), .Z(n1216) );
XOR2_X1 U871 ( .A(n1219), .B(n1220), .Z(n1217) );
AND2_X1 U872 ( .A1(G472), .A2(n1215), .ZN(n1220) );
NAND3_X1 U873 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1219) );
INV_X1 U874 ( .A(n1224), .ZN(n1223) );
NAND2_X1 U875 ( .A1(n1225), .A2(n1226), .ZN(n1222) );
INV_X1 U876 ( .A(KEYINPUT33), .ZN(n1226) );
XNOR2_X1 U877 ( .A(n1227), .B(n1228), .ZN(n1225) );
AND2_X1 U878 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
NAND2_X1 U879 ( .A1(KEYINPUT33), .A2(n1231), .ZN(n1221) );
NOR2_X1 U880 ( .A1(n1201), .A2(n1232), .ZN(G54) );
XOR2_X1 U881 ( .A(n1233), .B(n1234), .Z(n1232) );
AND2_X1 U882 ( .A1(G469), .A2(n1215), .ZN(n1233) );
NOR2_X1 U883 ( .A1(n1201), .A2(n1235), .ZN(G51) );
XOR2_X1 U884 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U885 ( .A(n1238), .B(n1239), .Z(n1237) );
NOR2_X1 U886 ( .A1(KEYINPUT52), .A2(n1240), .ZN(n1239) );
XNOR2_X1 U887 ( .A(n1241), .B(n1242), .ZN(n1240) );
XOR2_X1 U888 ( .A(KEYINPUT27), .B(n1243), .Z(n1242) );
NAND3_X1 U889 ( .A1(G210), .A2(n1244), .A3(n1215), .ZN(n1236) );
INV_X1 U890 ( .A(n1206), .ZN(n1215) );
NAND2_X1 U891 ( .A1(n1245), .A2(n1246), .ZN(n1206) );
NAND3_X1 U892 ( .A1(n1097), .A2(n1098), .A3(n1247), .ZN(n1246) );
INV_X1 U893 ( .A(n1122), .ZN(n1247) );
NAND2_X1 U894 ( .A1(n1248), .A2(n1249), .ZN(n1122) );
NOR4_X1 U895 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1249) );
AND4_X1 U896 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1248) );
OR3_X1 U897 ( .A1(n1258), .A2(n1259), .A3(n1112), .ZN(n1257) );
XNOR2_X1 U898 ( .A(n1260), .B(KEYINPUT9), .ZN(n1259) );
AND4_X1 U899 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1098) );
NAND2_X1 U900 ( .A1(n1265), .A2(n1266), .ZN(n1261) );
XNOR2_X1 U901 ( .A(KEYINPUT14), .B(n1105), .ZN(n1266) );
XOR2_X1 U902 ( .A(n1267), .B(KEYINPUT16), .Z(n1097) );
NAND2_X1 U903 ( .A1(n1268), .A2(n1186), .ZN(n1267) );
AND4_X1 U904 ( .A1(n1269), .A2(n1093), .A3(n1270), .A4(n1271), .ZN(n1186) );
NAND2_X1 U905 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
INV_X1 U906 ( .A(KEYINPUT39), .ZN(n1273) );
NAND4_X1 U907 ( .A1(n1274), .A2(n1109), .A3(n1136), .A4(KEYINPUT39), .ZN(n1270) );
INV_X1 U908 ( .A(n1146), .ZN(n1109) );
NAND3_X1 U909 ( .A1(n1139), .A2(n1274), .A3(n1128), .ZN(n1093) );
XOR2_X1 U910 ( .A(n1185), .B(KEYINPUT40), .Z(n1268) );
NAND3_X1 U911 ( .A1(n1139), .A2(n1274), .A3(n1275), .ZN(n1185) );
XNOR2_X1 U912 ( .A(G902), .B(KEYINPUT12), .ZN(n1245) );
XOR2_X1 U913 ( .A(KEYINPUT61), .B(n1276), .Z(n1244) );
NOR2_X1 U914 ( .A1(n1143), .A2(G952), .ZN(n1201) );
XNOR2_X1 U915 ( .A(n1277), .B(n1253), .ZN(G48) );
AND3_X1 U916 ( .A1(n1275), .A2(n1278), .A3(n1279), .ZN(n1253) );
XNOR2_X1 U917 ( .A(n1280), .B(n1281), .ZN(G45) );
NOR4_X1 U918 ( .A1(KEYINPUT50), .A2(n1120), .A3(n1258), .A4(n1282), .ZN(n1281) );
XNOR2_X1 U919 ( .A(KEYINPUT35), .B(n1112), .ZN(n1282) );
NAND4_X1 U920 ( .A1(n1118), .A2(n1283), .A3(n1284), .A4(n1285), .ZN(n1258) );
XNOR2_X1 U921 ( .A(G140), .B(n1256), .ZN(G42) );
NAND3_X1 U922 ( .A1(n1133), .A2(n1260), .A3(n1286), .ZN(n1256) );
XNOR2_X1 U923 ( .A(n1252), .B(n1287), .ZN(G39) );
NAND2_X1 U924 ( .A1(KEYINPUT31), .A2(G137), .ZN(n1287) );
AND3_X1 U925 ( .A1(n1146), .A2(n1133), .A3(n1279), .ZN(n1252) );
XOR2_X1 U926 ( .A(G134), .B(n1251), .Z(G36) );
AND2_X1 U927 ( .A1(n1288), .A2(n1128), .ZN(n1251) );
XNOR2_X1 U928 ( .A(G131), .B(n1289), .ZN(G33) );
NAND2_X1 U929 ( .A1(KEYINPUT29), .A2(n1250), .ZN(n1289) );
AND2_X1 U930 ( .A1(n1275), .A2(n1288), .ZN(n1250) );
AND4_X1 U931 ( .A1(n1118), .A2(n1133), .A3(n1260), .A4(n1285), .ZN(n1288) );
NOR2_X1 U932 ( .A1(n1141), .A2(n1290), .ZN(n1133) );
NAND2_X1 U933 ( .A1(n1291), .A2(n1292), .ZN(G30) );
NAND2_X1 U934 ( .A1(G128), .A2(n1255), .ZN(n1292) );
XOR2_X1 U935 ( .A(KEYINPUT17), .B(n1293), .Z(n1291) );
NOR2_X1 U936 ( .A1(G128), .A2(n1255), .ZN(n1293) );
NAND3_X1 U937 ( .A1(n1128), .A2(n1278), .A3(n1279), .ZN(n1255) );
AND4_X1 U938 ( .A1(n1260), .A2(n1151), .A3(n1285), .A4(n1294), .ZN(n1279) );
XNOR2_X1 U939 ( .A(n1269), .B(n1295), .ZN(G3) );
NOR2_X1 U940 ( .A1(KEYINPUT37), .A2(n1296), .ZN(n1295) );
NAND3_X1 U941 ( .A1(n1146), .A2(n1274), .A3(n1118), .ZN(n1269) );
XNOR2_X1 U942 ( .A(n1174), .B(n1297), .ZN(G27) );
NOR2_X1 U943 ( .A1(KEYINPUT0), .A2(n1254), .ZN(n1297) );
NAND3_X1 U944 ( .A1(n1286), .A2(n1278), .A3(n1119), .ZN(n1254) );
AND3_X1 U945 ( .A1(n1275), .A2(n1285), .A3(n1136), .ZN(n1286) );
NAND2_X1 U946 ( .A1(n1107), .A2(n1298), .ZN(n1285) );
NAND4_X1 U947 ( .A1(G953), .A2(G902), .A3(n1299), .A4(n1162), .ZN(n1298) );
INV_X1 U948 ( .A(G900), .ZN(n1162) );
XNOR2_X1 U949 ( .A(G122), .B(n1262), .ZN(G24) );
NAND4_X1 U950 ( .A1(n1300), .A2(n1139), .A3(n1283), .A4(n1284), .ZN(n1262) );
NOR2_X1 U951 ( .A1(n1294), .A2(n1151), .ZN(n1139) );
XNOR2_X1 U952 ( .A(G119), .B(n1263), .ZN(G21) );
NAND4_X1 U953 ( .A1(n1300), .A2(n1146), .A3(n1151), .A4(n1294), .ZN(n1263) );
INV_X1 U954 ( .A(n1301), .ZN(n1294) );
XNOR2_X1 U955 ( .A(G116), .B(n1264), .ZN(G18) );
NAND2_X1 U956 ( .A1(n1265), .A2(n1128), .ZN(n1264) );
NOR2_X1 U957 ( .A1(n1284), .A2(n1302), .ZN(n1128) );
XNOR2_X1 U958 ( .A(G113), .B(n1303), .ZN(G15) );
NAND2_X1 U959 ( .A1(n1265), .A2(n1275), .ZN(n1303) );
INV_X1 U960 ( .A(n1105), .ZN(n1275) );
NAND2_X1 U961 ( .A1(n1302), .A2(n1284), .ZN(n1105) );
INV_X1 U962 ( .A(n1283), .ZN(n1302) );
AND2_X1 U963 ( .A1(n1300), .A2(n1118), .ZN(n1265) );
NOR2_X1 U964 ( .A1(n1151), .A2(n1301), .ZN(n1118) );
AND2_X1 U965 ( .A1(n1119), .A2(n1304), .ZN(n1300) );
NOR2_X1 U966 ( .A1(n1138), .A2(n1149), .ZN(n1119) );
INV_X1 U967 ( .A(n1137), .ZN(n1149) );
XNOR2_X1 U968 ( .A(n1305), .B(n1272), .ZN(G12) );
AND3_X1 U969 ( .A1(n1146), .A2(n1274), .A3(n1136), .ZN(n1272) );
AND2_X1 U970 ( .A1(n1301), .A2(n1151), .ZN(n1136) );
XOR2_X1 U971 ( .A(n1306), .B(n1205), .Z(n1151) );
NAND2_X1 U972 ( .A1(G217), .A2(n1307), .ZN(n1205) );
NAND2_X1 U973 ( .A1(n1203), .A2(n1308), .ZN(n1306) );
XNOR2_X1 U974 ( .A(n1309), .B(n1310), .ZN(n1203) );
XNOR2_X1 U975 ( .A(n1174), .B(n1311), .ZN(n1310) );
XNOR2_X1 U976 ( .A(n1277), .B(G140), .ZN(n1311) );
INV_X1 U977 ( .A(G125), .ZN(n1174) );
XOR2_X1 U978 ( .A(n1312), .B(n1313), .Z(n1309) );
NOR3_X1 U979 ( .A1(n1314), .A2(KEYINPUT26), .A3(n1315), .ZN(n1313) );
NOR2_X1 U980 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XOR2_X1 U981 ( .A(KEYINPUT10), .B(n1318), .Z(n1314) );
AND2_X1 U982 ( .A1(n1316), .A2(n1317), .ZN(n1318) );
INV_X1 U983 ( .A(G137), .ZN(n1317) );
NAND3_X1 U984 ( .A1(n1319), .A2(n1143), .A3(G221), .ZN(n1316) );
XOR2_X1 U985 ( .A(KEYINPUT1), .B(G234), .Z(n1319) );
NAND3_X1 U986 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1312) );
NAND2_X1 U987 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
OR3_X1 U988 ( .A1(n1324), .A2(n1323), .A3(n1305), .ZN(n1321) );
INV_X1 U989 ( .A(KEYINPUT7), .ZN(n1324) );
NAND2_X1 U990 ( .A1(n1325), .A2(n1305), .ZN(n1320) );
NAND2_X1 U991 ( .A1(n1326), .A2(KEYINPUT7), .ZN(n1325) );
XNOR2_X1 U992 ( .A(n1323), .B(KEYINPUT60), .ZN(n1326) );
XNOR2_X1 U993 ( .A(n1327), .B(n1328), .ZN(n1323) );
NAND2_X1 U994 ( .A1(KEYINPUT38), .A2(n1329), .ZN(n1327) );
NOR2_X1 U995 ( .A1(n1330), .A2(n1148), .ZN(n1301) );
NOR2_X1 U996 ( .A1(n1154), .A2(G472), .ZN(n1148) );
AND2_X1 U997 ( .A1(G472), .A2(n1154), .ZN(n1330) );
NAND2_X1 U998 ( .A1(n1331), .A2(n1308), .ZN(n1154) );
XOR2_X1 U999 ( .A(n1332), .B(n1218), .Z(n1331) );
XNOR2_X1 U1000 ( .A(n1296), .B(n1333), .ZN(n1218) );
NOR2_X1 U1001 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
INV_X1 U1002 ( .A(G210), .ZN(n1335) );
NOR2_X1 U1003 ( .A1(n1224), .A2(n1231), .ZN(n1332) );
NAND2_X1 U1004 ( .A1(n1336), .A2(n1337), .ZN(n1231) );
NAND2_X1 U1005 ( .A1(n1338), .A2(n1230), .ZN(n1337) );
XOR2_X1 U1006 ( .A(n1228), .B(n1229), .Z(n1338) );
NAND3_X1 U1007 ( .A1(n1229), .A2(n1228), .A3(n1339), .ZN(n1336) );
NOR3_X1 U1008 ( .A1(n1228), .A2(n1230), .A3(n1229), .ZN(n1224) );
XNOR2_X1 U1009 ( .A(n1340), .B(n1341), .ZN(n1228) );
XOR2_X1 U1010 ( .A(n1342), .B(G116), .Z(n1340) );
NAND2_X1 U1011 ( .A1(KEYINPUT4), .A2(n1328), .ZN(n1342) );
AND2_X1 U1012 ( .A1(n1260), .A2(n1304), .ZN(n1274) );
AND2_X1 U1013 ( .A1(n1278), .A2(n1343), .ZN(n1304) );
NAND2_X1 U1014 ( .A1(n1107), .A2(n1344), .ZN(n1343) );
NAND4_X1 U1015 ( .A1(G953), .A2(G902), .A3(n1299), .A4(n1200), .ZN(n1344) );
INV_X1 U1016 ( .A(G898), .ZN(n1200) );
NAND3_X1 U1017 ( .A1(n1299), .A2(n1143), .A3(G952), .ZN(n1107) );
NAND2_X1 U1018 ( .A1(G234), .A2(G237), .ZN(n1299) );
INV_X1 U1019 ( .A(n1112), .ZN(n1278) );
NAND2_X1 U1020 ( .A1(n1141), .A2(n1140), .ZN(n1112) );
INV_X1 U1021 ( .A(n1290), .ZN(n1140) );
NOR2_X1 U1022 ( .A1(n1345), .A2(n1276), .ZN(n1290) );
NOR2_X1 U1023 ( .A1(G902), .A2(G237), .ZN(n1276) );
NAND3_X1 U1024 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1141) );
NAND2_X1 U1025 ( .A1(G902), .A2(G210), .ZN(n1348) );
NAND3_X1 U1026 ( .A1(n1349), .A2(n1308), .A3(n1350), .ZN(n1347) );
OR2_X1 U1027 ( .A1(n1350), .A2(n1349), .ZN(n1346) );
XNOR2_X1 U1028 ( .A(n1351), .B(n1352), .ZN(n1349) );
XNOR2_X1 U1029 ( .A(KEYINPUT6), .B(n1238), .ZN(n1352) );
NAND3_X1 U1030 ( .A1(n1353), .A2(n1354), .A3(n1199), .ZN(n1238) );
NAND3_X1 U1031 ( .A1(n1196), .A2(n1197), .A3(n1193), .ZN(n1199) );
NAND2_X1 U1032 ( .A1(n1355), .A2(n1191), .ZN(n1354) );
XNOR2_X1 U1033 ( .A(n1195), .B(n1197), .ZN(n1355) );
OR3_X1 U1034 ( .A1(n1193), .A2(n1197), .A3(n1191), .ZN(n1353) );
INV_X1 U1035 ( .A(n1196), .ZN(n1191) );
XNOR2_X1 U1036 ( .A(G110), .B(n1356), .ZN(n1196) );
XOR2_X1 U1037 ( .A(n1357), .B(n1296), .Z(n1197) );
INV_X1 U1038 ( .A(G101), .ZN(n1296) );
NAND2_X1 U1039 ( .A1(KEYINPUT32), .A2(n1358), .ZN(n1357) );
XNOR2_X1 U1040 ( .A(n1359), .B(n1360), .ZN(n1358) );
INV_X1 U1041 ( .A(n1195), .ZN(n1193) );
XNOR2_X1 U1042 ( .A(n1361), .B(n1328), .ZN(n1195) );
XOR2_X1 U1043 ( .A(G119), .B(KEYINPUT2), .Z(n1328) );
XNOR2_X1 U1044 ( .A(n1362), .B(n1363), .ZN(n1361) );
NOR2_X1 U1045 ( .A1(KEYINPUT15), .A2(n1364), .ZN(n1363) );
NOR2_X1 U1046 ( .A1(G116), .A2(KEYINPUT18), .ZN(n1362) );
NAND2_X1 U1047 ( .A1(KEYINPUT36), .A2(n1365), .ZN(n1351) );
XNOR2_X1 U1048 ( .A(n1243), .B(n1366), .ZN(n1365) );
NAND2_X1 U1049 ( .A1(KEYINPUT20), .A2(n1367), .ZN(n1366) );
XOR2_X1 U1050 ( .A(KEYINPUT51), .B(n1241), .Z(n1367) );
XOR2_X1 U1051 ( .A(G125), .B(n1229), .Z(n1241) );
XOR2_X1 U1052 ( .A(n1368), .B(n1369), .Z(n1229) );
NOR2_X1 U1053 ( .A1(G128), .A2(KEYINPUT25), .ZN(n1369) );
NOR2_X1 U1054 ( .A1(n1179), .A2(G953), .ZN(n1243) );
INV_X1 U1055 ( .A(G224), .ZN(n1179) );
NAND2_X1 U1056 ( .A1(G210), .A2(G237), .ZN(n1350) );
INV_X1 U1057 ( .A(n1120), .ZN(n1260) );
NAND2_X1 U1058 ( .A1(n1138), .A2(n1137), .ZN(n1120) );
NAND2_X1 U1059 ( .A1(G221), .A2(n1307), .ZN(n1137) );
NAND2_X1 U1060 ( .A1(G234), .A2(n1308), .ZN(n1307) );
XNOR2_X1 U1061 ( .A(n1145), .B(KEYINPUT53), .ZN(n1138) );
XOR2_X1 U1062 ( .A(n1370), .B(G469), .Z(n1145) );
OR2_X1 U1063 ( .A1(n1234), .A2(G902), .ZN(n1370) );
XNOR2_X1 U1064 ( .A(n1371), .B(n1372), .ZN(n1234) );
XNOR2_X1 U1065 ( .A(n1230), .B(n1373), .ZN(n1372) );
XOR2_X1 U1066 ( .A(n1374), .B(n1166), .Z(n1373) );
XOR2_X1 U1067 ( .A(n1375), .B(n1376), .Z(n1166) );
XNOR2_X1 U1068 ( .A(n1280), .B(G128), .ZN(n1376) );
NAND2_X1 U1069 ( .A1(KEYINPUT24), .A2(n1277), .ZN(n1375) );
NAND2_X1 U1070 ( .A1(G227), .A2(n1143), .ZN(n1374) );
INV_X1 U1071 ( .A(n1339), .ZN(n1230) );
XOR2_X1 U1072 ( .A(n1377), .B(n1378), .Z(n1339) );
INV_X1 U1073 ( .A(n1168), .ZN(n1378) );
XOR2_X1 U1074 ( .A(G134), .B(KEYINPUT49), .Z(n1168) );
XNOR2_X1 U1075 ( .A(n1379), .B(n1380), .ZN(n1377) );
NOR2_X1 U1076 ( .A1(G137), .A2(KEYINPUT56), .ZN(n1380) );
NOR2_X1 U1077 ( .A1(KEYINPUT22), .A2(n1381), .ZN(n1379) );
XNOR2_X1 U1078 ( .A(KEYINPUT59), .B(n1171), .ZN(n1381) );
INV_X1 U1079 ( .A(G131), .ZN(n1171) );
XOR2_X1 U1080 ( .A(n1382), .B(n1383), .Z(n1371) );
XNOR2_X1 U1081 ( .A(G101), .B(n1384), .ZN(n1383) );
NAND3_X1 U1082 ( .A1(n1385), .A2(n1386), .A3(n1387), .ZN(n1384) );
NAND2_X1 U1083 ( .A1(n1360), .A2(n1388), .ZN(n1387) );
INV_X1 U1084 ( .A(KEYINPUT57), .ZN(n1388) );
NAND3_X1 U1085 ( .A1(KEYINPUT57), .A2(n1389), .A3(n1359), .ZN(n1386) );
OR2_X1 U1086 ( .A1(n1359), .A2(n1389), .ZN(n1385) );
NOR2_X1 U1087 ( .A1(n1390), .A2(n1360), .ZN(n1389) );
XOR2_X1 U1088 ( .A(G104), .B(KEYINPUT21), .Z(n1360) );
INV_X1 U1089 ( .A(KEYINPUT19), .ZN(n1390) );
XNOR2_X1 U1090 ( .A(G110), .B(G140), .ZN(n1382) );
NOR2_X1 U1091 ( .A1(n1283), .A2(n1284), .ZN(n1146) );
XNOR2_X1 U1092 ( .A(n1391), .B(G475), .ZN(n1284) );
NAND2_X1 U1093 ( .A1(n1213), .A2(n1308), .ZN(n1391) );
XNOR2_X1 U1094 ( .A(n1392), .B(n1393), .ZN(n1213) );
XOR2_X1 U1095 ( .A(n1394), .B(n1395), .Z(n1393) );
XOR2_X1 U1096 ( .A(n1396), .B(n1368), .Z(n1395) );
XNOR2_X1 U1097 ( .A(G143), .B(n1277), .ZN(n1368) );
INV_X1 U1098 ( .A(G146), .ZN(n1277) );
NAND2_X1 U1099 ( .A1(n1397), .A2(KEYINPUT13), .ZN(n1396) );
XNOR2_X1 U1100 ( .A(G125), .B(n1398), .ZN(n1397) );
NOR2_X1 U1101 ( .A1(G140), .A2(KEYINPUT48), .ZN(n1398) );
NAND2_X1 U1102 ( .A1(n1399), .A2(n1400), .ZN(n1394) );
NAND2_X1 U1103 ( .A1(n1401), .A2(n1356), .ZN(n1400) );
XNOR2_X1 U1104 ( .A(n1364), .B(KEYINPUT46), .ZN(n1401) );
NAND2_X1 U1105 ( .A1(n1402), .A2(G122), .ZN(n1399) );
XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1341), .ZN(n1402) );
INV_X1 U1107 ( .A(n1364), .ZN(n1341) );
XOR2_X1 U1108 ( .A(G113), .B(KEYINPUT63), .Z(n1364) );
XOR2_X1 U1109 ( .A(n1403), .B(n1404), .Z(n1392) );
NOR2_X1 U1110 ( .A1(n1334), .A2(n1345), .ZN(n1404) );
INV_X1 U1111 ( .A(G214), .ZN(n1345) );
NAND2_X1 U1112 ( .A1(n1405), .A2(n1143), .ZN(n1334) );
XOR2_X1 U1113 ( .A(KEYINPUT47), .B(G237), .Z(n1405) );
XNOR2_X1 U1114 ( .A(G104), .B(G131), .ZN(n1403) );
XOR2_X1 U1115 ( .A(n1406), .B(n1211), .Z(n1283) );
INV_X1 U1116 ( .A(G478), .ZN(n1211) );
NAND2_X1 U1117 ( .A1(n1407), .A2(n1308), .ZN(n1406) );
INV_X1 U1118 ( .A(G902), .ZN(n1308) );
XNOR2_X1 U1119 ( .A(n1209), .B(KEYINPUT45), .ZN(n1407) );
XNOR2_X1 U1120 ( .A(n1408), .B(n1409), .ZN(n1209) );
XOR2_X1 U1121 ( .A(n1410), .B(n1411), .Z(n1409) );
NAND3_X1 U1122 ( .A1(G217), .A2(n1143), .A3(G234), .ZN(n1411) );
INV_X1 U1123 ( .A(G953), .ZN(n1143) );
NAND2_X1 U1124 ( .A1(n1412), .A2(n1413), .ZN(n1410) );
NAND2_X1 U1125 ( .A1(G116), .A2(n1356), .ZN(n1413) );
XOR2_X1 U1126 ( .A(n1414), .B(KEYINPUT3), .Z(n1412) );
OR2_X1 U1127 ( .A1(n1356), .A2(G116), .ZN(n1414) );
INV_X1 U1128 ( .A(G122), .ZN(n1356) );
XNOR2_X1 U1129 ( .A(n1415), .B(n1359), .ZN(n1408) );
INV_X1 U1130 ( .A(G107), .ZN(n1359) );
NAND2_X1 U1131 ( .A1(n1416), .A2(KEYINPUT11), .ZN(n1415) );
XOR2_X1 U1132 ( .A(n1417), .B(G134), .Z(n1416) );
NAND3_X1 U1133 ( .A1(n1418), .A2(n1419), .A3(n1420), .ZN(n1417) );
OR2_X1 U1134 ( .A1(n1329), .A2(KEYINPUT30), .ZN(n1420) );
NAND3_X1 U1135 ( .A1(KEYINPUT30), .A2(n1329), .A3(G143), .ZN(n1419) );
NAND2_X1 U1136 ( .A1(n1421), .A2(n1280), .ZN(n1418) );
INV_X1 U1137 ( .A(G143), .ZN(n1280) );
NAND2_X1 U1138 ( .A1(KEYINPUT30), .A2(n1422), .ZN(n1421) );
XNOR2_X1 U1139 ( .A(KEYINPUT8), .B(n1329), .ZN(n1422) );
INV_X1 U1140 ( .A(G128), .ZN(n1329) );
INV_X1 U1141 ( .A(G110), .ZN(n1305) );
endmodule


