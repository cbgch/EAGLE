//Key = 0010101100100111011110100010110100100110001110001001100111100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;

XOR2_X1 U719 ( .A(G107), .B(n997), .Z(G9) );
NAND4_X1 U720 ( .A1(n998), .A2(n999), .A3(n1000), .A4(n1001), .ZN(G75) );
NAND4_X1 U721 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n1000) );
NOR4_X1 U722 ( .A1(n1006), .A2(n1007), .A3(n1008), .A4(n1009), .ZN(n1005) );
XOR2_X1 U723 ( .A(n1010), .B(n1011), .Z(n1008) );
NAND2_X1 U724 ( .A1(KEYINPUT55), .A2(n1012), .ZN(n1010) );
NOR2_X1 U725 ( .A1(n1013), .A2(n1014), .ZN(n1004) );
NOR2_X1 U726 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
INV_X1 U727 ( .A(KEYINPUT62), .ZN(n1016) );
NOR3_X1 U728 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1015) );
NOR2_X1 U729 ( .A1(KEYINPUT62), .A2(n1020), .ZN(n1013) );
NAND2_X1 U730 ( .A1(n1021), .A2(n1022), .ZN(n999) );
NAND2_X1 U731 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND4_X1 U732 ( .A1(n1025), .A2(n1002), .A3(n1020), .A4(n1026), .ZN(n1024) );
NAND2_X1 U733 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U734 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND2_X1 U735 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
OR2_X1 U736 ( .A1(n1033), .A2(n1009), .ZN(n1032) );
NAND2_X1 U737 ( .A1(n1034), .A2(n1035), .ZN(n1027) );
NAND2_X1 U738 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U739 ( .A1(n1003), .A2(n1006), .ZN(n1037) );
NAND3_X1 U740 ( .A1(n1034), .A2(n1038), .A3(n1029), .ZN(n1023) );
NAND2_X1 U741 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U742 ( .A1(n1002), .A2(n1041), .ZN(n1040) );
NAND2_X1 U743 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U744 ( .A1(n1025), .A2(n1044), .ZN(n1043) );
NAND2_X1 U745 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U746 ( .A1(n1007), .A2(n1020), .ZN(n1042) );
NAND2_X1 U747 ( .A1(n1020), .A2(n1047), .ZN(n1039) );
INV_X1 U748 ( .A(n1048), .ZN(n1021) );
XOR2_X1 U749 ( .A(n1049), .B(n1050), .Z(G72) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U751 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
XOR2_X1 U752 ( .A(n1056), .B(KEYINPUT51), .Z(n1055) );
NOR2_X1 U753 ( .A1(G900), .A2(n1001), .ZN(n1054) );
XNOR2_X1 U754 ( .A(n1057), .B(n1058), .ZN(n1053) );
NOR2_X1 U755 ( .A1(n1059), .A2(n1056), .ZN(n1051) );
NAND2_X1 U756 ( .A1(n1060), .A2(n1001), .ZN(n1056) );
XOR2_X1 U757 ( .A(n1061), .B(KEYINPUT59), .Z(n1060) );
XOR2_X1 U758 ( .A(n1058), .B(n1057), .Z(n1059) );
AND2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1058) );
NAND2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U761 ( .A1(n1066), .A2(n1067), .ZN(n1062) );
INV_X1 U762 ( .A(n1064), .ZN(n1067) );
XNOR2_X1 U763 ( .A(KEYINPUT36), .B(n1065), .ZN(n1066) );
NAND3_X1 U764 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1065) );
NAND2_X1 U765 ( .A1(KEYINPUT0), .A2(G131), .ZN(n1070) );
NAND3_X1 U766 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1069) );
INV_X1 U767 ( .A(KEYINPUT0), .ZN(n1072) );
OR2_X1 U768 ( .A1(n1073), .A2(n1071), .ZN(n1068) );
AND2_X1 U769 ( .A1(KEYINPUT43), .A2(n1074), .ZN(n1071) );
XOR2_X1 U770 ( .A(G137), .B(n1075), .Z(n1073) );
NAND2_X1 U771 ( .A1(G953), .A2(n1076), .ZN(n1049) );
NAND2_X1 U772 ( .A1(G900), .A2(G227), .ZN(n1076) );
XOR2_X1 U773 ( .A(n1077), .B(n1078), .Z(G69) );
XOR2_X1 U774 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U775 ( .A1(n1081), .A2(n1001), .ZN(n1080) );
NOR2_X1 U776 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U777 ( .A1(n1084), .A2(n1085), .ZN(n1079) );
NAND2_X1 U778 ( .A1(G953), .A2(n1083), .ZN(n1085) );
XOR2_X1 U779 ( .A(n1086), .B(n1087), .Z(n1084) );
NAND2_X1 U780 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
OR2_X1 U781 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U782 ( .A(n1092), .B(KEYINPUT5), .Z(n1088) );
NAND2_X1 U783 ( .A1(n1091), .A2(n1090), .ZN(n1092) );
NAND2_X1 U784 ( .A1(n1001), .A2(n1093), .ZN(n1077) );
NOR3_X1 U785 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(G66) );
NOR3_X1 U786 ( .A1(n1097), .A2(G952), .A3(n1098), .ZN(n1096) );
INV_X1 U787 ( .A(KEYINPUT50), .ZN(n1097) );
NOR2_X1 U788 ( .A1(KEYINPUT50), .A2(n1099), .ZN(n1095) );
INV_X1 U789 ( .A(n1100), .ZN(n1099) );
XOR2_X1 U790 ( .A(n1101), .B(n1102), .Z(n1094) );
NAND3_X1 U791 ( .A1(n1103), .A2(n1011), .A3(KEYINPUT13), .ZN(n1101) );
NOR2_X1 U792 ( .A1(n1104), .A2(n1105), .ZN(G63) );
XNOR2_X1 U793 ( .A(n1100), .B(KEYINPUT57), .ZN(n1105) );
XOR2_X1 U794 ( .A(n1106), .B(n1107), .Z(n1104) );
NAND2_X1 U795 ( .A1(KEYINPUT18), .A2(n1108), .ZN(n1106) );
NAND2_X1 U796 ( .A1(n1103), .A2(G478), .ZN(n1108) );
NOR2_X1 U797 ( .A1(n1100), .A2(n1109), .ZN(G60) );
XOR2_X1 U798 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U799 ( .A1(KEYINPUT47), .A2(n1112), .ZN(n1111) );
NOR2_X1 U800 ( .A1(n1019), .A2(n1113), .ZN(n1110) );
INV_X1 U801 ( .A(G475), .ZN(n1019) );
XOR2_X1 U802 ( .A(n1114), .B(n1115), .Z(G6) );
NAND2_X1 U803 ( .A1(KEYINPUT52), .A2(G104), .ZN(n1115) );
NOR2_X1 U804 ( .A1(n1100), .A2(n1116), .ZN(G57) );
XOR2_X1 U805 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U806 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U807 ( .A1(KEYINPUT20), .A2(n1121), .ZN(n1119) );
NAND2_X1 U808 ( .A1(n1103), .A2(G472), .ZN(n1121) );
XOR2_X1 U809 ( .A(n1122), .B(n1123), .Z(n1117) );
NOR2_X1 U810 ( .A1(KEYINPUT45), .A2(n1124), .ZN(n1123) );
XOR2_X1 U811 ( .A(n1125), .B(KEYINPUT9), .Z(n1122) );
NOR2_X1 U812 ( .A1(n1100), .A2(n1126), .ZN(G54) );
XOR2_X1 U813 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND2_X1 U814 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U815 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U816 ( .A(n1133), .B(KEYINPUT49), .Z(n1129) );
OR2_X1 U817 ( .A1(n1132), .A2(n1131), .ZN(n1133) );
AND2_X1 U818 ( .A1(n1134), .A2(n1135), .ZN(n1131) );
NAND2_X1 U819 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U820 ( .A1(n1138), .A2(n1139), .ZN(n1136) );
NAND3_X1 U821 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1134) );
INV_X1 U822 ( .A(n1137), .ZN(n1140) );
NAND2_X1 U823 ( .A1(G140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U824 ( .A(n1142), .B(KEYINPUT33), .Z(n1138) );
OR2_X1 U825 ( .A1(n1141), .A2(G140), .ZN(n1142) );
NAND2_X1 U826 ( .A1(n1103), .A2(G469), .ZN(n1127) );
NOR2_X1 U827 ( .A1(n1100), .A2(n1143), .ZN(G51) );
XOR2_X1 U828 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U829 ( .A(n1146), .B(n1147), .Z(n1145) );
XNOR2_X1 U830 ( .A(KEYINPUT24), .B(n1148), .ZN(n1147) );
XOR2_X1 U831 ( .A(n1149), .B(n1150), .Z(n1144) );
XOR2_X1 U832 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U833 ( .A1(KEYINPUT56), .A2(n1153), .ZN(n1152) );
INV_X1 U834 ( .A(n1154), .ZN(n1153) );
NAND3_X1 U835 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1151) );
NAND2_X1 U836 ( .A1(KEYINPUT6), .A2(n1113), .ZN(n1156) );
INV_X1 U837 ( .A(n1103), .ZN(n1113) );
NOR2_X1 U838 ( .A1(n1158), .A2(n998), .ZN(n1103) );
NAND2_X1 U839 ( .A1(n1159), .A2(n1160), .ZN(n1155) );
INV_X1 U840 ( .A(KEYINPUT6), .ZN(n1160) );
NAND2_X1 U841 ( .A1(n998), .A2(G902), .ZN(n1159) );
NOR2_X1 U842 ( .A1(n1093), .A2(n1061), .ZN(n998) );
NAND4_X1 U843 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1061) );
NOR4_X1 U844 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
NOR2_X1 U845 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
INV_X1 U846 ( .A(KEYINPUT28), .ZN(n1170) );
NOR2_X1 U847 ( .A1(n1171), .A2(n1172), .ZN(n1167) );
NOR2_X1 U848 ( .A1(n1173), .A2(n1174), .ZN(n1166) );
NOR4_X1 U849 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1036), .ZN(n1165) );
NOR2_X1 U850 ( .A1(n1047), .A2(n1178), .ZN(n1176) );
NOR3_X1 U851 ( .A1(n1179), .A2(KEYINPUT28), .A3(n1046), .ZN(n1178) );
NOR2_X1 U852 ( .A1(n1180), .A2(n1181), .ZN(n1175) );
AND4_X1 U853 ( .A1(n1174), .A2(n1031), .A3(n1017), .A4(n1182), .ZN(n1180) );
INV_X1 U854 ( .A(KEYINPUT31), .ZN(n1174) );
NOR3_X1 U855 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1163) );
INV_X1 U856 ( .A(n1186), .ZN(n1183) );
NAND4_X1 U857 ( .A1(n1114), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1093) );
NOR4_X1 U858 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
NOR2_X1 U859 ( .A1(n997), .A2(n1194), .ZN(n1188) );
NOR3_X1 U860 ( .A1(n1031), .A2(n1195), .A3(n1196), .ZN(n1194) );
AND3_X1 U861 ( .A1(n1197), .A2(n1198), .A3(n1034), .ZN(n997) );
NAND3_X1 U862 ( .A1(n1034), .A2(n1197), .A3(n1199), .ZN(n1114) );
INV_X1 U863 ( .A(n1195), .ZN(n1197) );
NOR2_X1 U864 ( .A1(n1200), .A2(G952), .ZN(n1100) );
INV_X1 U865 ( .A(n1098), .ZN(n1200) );
XNOR2_X1 U866 ( .A(n1001), .B(KEYINPUT40), .ZN(n1098) );
XOR2_X1 U867 ( .A(n1161), .B(n1201), .Z(G48) );
NAND2_X1 U868 ( .A1(KEYINPUT15), .A2(G146), .ZN(n1201) );
NAND3_X1 U869 ( .A1(n1199), .A2(n1202), .A3(n1203), .ZN(n1161) );
XNOR2_X1 U870 ( .A(G143), .B(n1173), .ZN(G45) );
NAND4_X1 U871 ( .A1(n1204), .A2(n1202), .A3(n1182), .A4(n1017), .ZN(n1173) );
XNOR2_X1 U872 ( .A(n1205), .B(n1162), .ZN(G42) );
NAND3_X1 U873 ( .A1(n1029), .A2(n1047), .A3(n1206), .ZN(n1162) );
XNOR2_X1 U874 ( .A(G140), .B(KEYINPUT42), .ZN(n1205) );
XNOR2_X1 U875 ( .A(n1207), .B(n1185), .ZN(G39) );
AND3_X1 U876 ( .A1(n1029), .A2(n1020), .A3(n1203), .ZN(n1185) );
INV_X1 U877 ( .A(n1196), .ZN(n1020) );
XOR2_X1 U878 ( .A(G134), .B(n1208), .Z(G36) );
NOR2_X1 U879 ( .A1(n1171), .A2(n1209), .ZN(n1208) );
XNOR2_X1 U880 ( .A(KEYINPUT14), .B(n1172), .ZN(n1209) );
NAND2_X1 U881 ( .A1(n1204), .A2(n1198), .ZN(n1172) );
XOR2_X1 U882 ( .A(n1210), .B(n1184), .Z(G33) );
AND3_X1 U883 ( .A1(n1204), .A2(n1199), .A3(n1029), .ZN(n1184) );
INV_X1 U884 ( .A(n1171), .ZN(n1029) );
NAND2_X1 U885 ( .A1(n1003), .A2(n1211), .ZN(n1171) );
INV_X1 U886 ( .A(n1212), .ZN(n1003) );
INV_X1 U887 ( .A(n1045), .ZN(n1199) );
NOR3_X1 U888 ( .A1(n1181), .A2(n1177), .A3(n1031), .ZN(n1204) );
NAND2_X1 U889 ( .A1(KEYINPUT61), .A2(n1074), .ZN(n1210) );
INV_X1 U890 ( .A(G131), .ZN(n1074) );
XNOR2_X1 U891 ( .A(n1169), .B(n1213), .ZN(G30) );
NOR2_X1 U892 ( .A1(KEYINPUT60), .A2(n1214), .ZN(n1213) );
NAND3_X1 U893 ( .A1(n1198), .A2(n1202), .A3(n1203), .ZN(n1169) );
NOR3_X1 U894 ( .A1(n1181), .A2(n1177), .A3(n1179), .ZN(n1203) );
INV_X1 U895 ( .A(n1047), .ZN(n1181) );
INV_X1 U896 ( .A(n1046), .ZN(n1198) );
XNOR2_X1 U897 ( .A(n1124), .B(n1215), .ZN(G3) );
NOR4_X1 U898 ( .A1(KEYINPUT27), .A2(n1195), .A3(n1196), .A4(n1031), .ZN(n1215) );
XNOR2_X1 U899 ( .A(G125), .B(n1186), .ZN(G27) );
NAND4_X1 U900 ( .A1(n1002), .A2(n1206), .A3(n1025), .A4(n1202), .ZN(n1186) );
NOR4_X1 U901 ( .A1(n1033), .A2(n1045), .A3(n1009), .A4(n1177), .ZN(n1206) );
AND2_X1 U902 ( .A1(n1216), .A2(n1048), .ZN(n1177) );
NAND4_X1 U903 ( .A1(G953), .A2(G902), .A3(n1217), .A4(n1218), .ZN(n1216) );
INV_X1 U904 ( .A(G900), .ZN(n1218) );
XNOR2_X1 U905 ( .A(G122), .B(n1187), .ZN(G24) );
NAND4_X1 U906 ( .A1(n1219), .A2(n1034), .A3(n1182), .A4(n1017), .ZN(n1187) );
NOR2_X1 U907 ( .A1(n1009), .A2(n1220), .ZN(n1034) );
INV_X1 U908 ( .A(n1221), .ZN(n1219) );
XOR2_X1 U909 ( .A(G119), .B(n1193), .Z(G21) );
NOR3_X1 U910 ( .A1(n1221), .A2(n1196), .A3(n1179), .ZN(n1193) );
NAND2_X1 U911 ( .A1(n1220), .A2(n1009), .ZN(n1179) );
INV_X1 U912 ( .A(n1033), .ZN(n1220) );
XOR2_X1 U913 ( .A(n1192), .B(n1222), .Z(G18) );
NOR2_X1 U914 ( .A1(KEYINPUT53), .A2(n1223), .ZN(n1222) );
NOR3_X1 U915 ( .A1(n1031), .A2(n1046), .A3(n1221), .ZN(n1192) );
NAND2_X1 U916 ( .A1(n1224), .A2(n1017), .ZN(n1046) );
XOR2_X1 U917 ( .A(G113), .B(n1191), .Z(G15) );
NOR3_X1 U918 ( .A1(n1031), .A2(n1045), .A3(n1221), .ZN(n1191) );
NAND4_X1 U919 ( .A1(n1025), .A2(n1002), .A3(n1202), .A4(n1225), .ZN(n1221) );
XNOR2_X1 U920 ( .A(n1007), .B(KEYINPUT12), .ZN(n1025) );
NAND2_X1 U921 ( .A1(n1226), .A2(n1182), .ZN(n1045) );
XNOR2_X1 U922 ( .A(n1224), .B(KEYINPUT41), .ZN(n1182) );
NAND2_X1 U923 ( .A1(n1033), .A2(n1009), .ZN(n1031) );
XNOR2_X1 U924 ( .A(n1190), .B(n1227), .ZN(G12) );
NAND2_X1 U925 ( .A1(KEYINPUT44), .A2(G110), .ZN(n1227) );
NOR4_X1 U926 ( .A1(n1033), .A2(n1196), .A3(n1009), .A4(n1195), .ZN(n1190) );
NAND3_X1 U927 ( .A1(n1202), .A2(n1225), .A3(n1047), .ZN(n1195) );
NOR2_X1 U928 ( .A1(n1002), .A2(n1007), .ZN(n1047) );
AND2_X1 U929 ( .A1(G221), .A2(n1228), .ZN(n1007) );
XOR2_X1 U930 ( .A(n1229), .B(G469), .Z(n1002) );
NAND2_X1 U931 ( .A1(n1230), .A2(n1158), .ZN(n1229) );
XOR2_X1 U932 ( .A(n1231), .B(n1232), .Z(n1230) );
XNOR2_X1 U933 ( .A(n1233), .B(n1137), .ZN(n1232) );
NAND2_X1 U934 ( .A1(n1234), .A2(n1001), .ZN(n1137) );
XNOR2_X1 U935 ( .A(G227), .B(KEYINPUT58), .ZN(n1234) );
NAND2_X1 U936 ( .A1(KEYINPUT29), .A2(n1132), .ZN(n1233) );
XNOR2_X1 U937 ( .A(n1235), .B(n1236), .ZN(n1132) );
XNOR2_X1 U938 ( .A(n1237), .B(n1238), .ZN(n1236) );
XNOR2_X1 U939 ( .A(n1064), .B(n1239), .ZN(n1235) );
XOR2_X1 U940 ( .A(n1240), .B(n1214), .Z(n1064) );
NAND3_X1 U941 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1240) );
NAND2_X1 U942 ( .A1(G146), .A2(n1244), .ZN(n1243) );
NAND2_X1 U943 ( .A1(KEYINPUT54), .A2(n1245), .ZN(n1242) );
NAND2_X1 U944 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XNOR2_X1 U945 ( .A(KEYINPUT39), .B(n1244), .ZN(n1246) );
NAND2_X1 U946 ( .A1(n1248), .A2(n1249), .ZN(n1241) );
INV_X1 U947 ( .A(KEYINPUT54), .ZN(n1249) );
NAND2_X1 U948 ( .A1(n1250), .A2(n1251), .ZN(n1248) );
NAND2_X1 U949 ( .A1(KEYINPUT39), .A2(n1244), .ZN(n1251) );
OR3_X1 U950 ( .A1(G146), .A2(KEYINPUT39), .A3(n1244), .ZN(n1250) );
XNOR2_X1 U951 ( .A(G110), .B(G140), .ZN(n1231) );
NAND2_X1 U952 ( .A1(n1048), .A2(n1252), .ZN(n1225) );
NAND4_X1 U953 ( .A1(G953), .A2(G902), .A3(n1217), .A4(n1083), .ZN(n1252) );
INV_X1 U954 ( .A(G898), .ZN(n1083) );
NAND3_X1 U955 ( .A1(n1217), .A2(n1001), .A3(G952), .ZN(n1048) );
NAND2_X1 U956 ( .A1(G237), .A2(G234), .ZN(n1217) );
INV_X1 U957 ( .A(n1036), .ZN(n1202) );
NAND2_X1 U958 ( .A1(n1211), .A2(n1212), .ZN(n1036) );
XNOR2_X1 U959 ( .A(n1253), .B(n1157), .ZN(n1212) );
AND2_X1 U960 ( .A1(G210), .A2(n1254), .ZN(n1157) );
NAND2_X1 U961 ( .A1(n1255), .A2(n1158), .ZN(n1253) );
XOR2_X1 U962 ( .A(n1256), .B(n1257), .Z(n1255) );
NOR2_X1 U963 ( .A1(KEYINPUT32), .A2(n1154), .ZN(n1257) );
XNOR2_X1 U964 ( .A(n1258), .B(n1259), .ZN(n1154) );
XNOR2_X1 U965 ( .A(KEYINPUT23), .B(n1091), .ZN(n1259) );
XNOR2_X1 U966 ( .A(n1090), .B(n1087), .ZN(n1258) );
XNOR2_X1 U967 ( .A(G122), .B(n1141), .ZN(n1087) );
INV_X1 U968 ( .A(G110), .ZN(n1141) );
XNOR2_X1 U969 ( .A(n1260), .B(n1238), .ZN(n1090) );
XNOR2_X1 U970 ( .A(n1124), .B(n1261), .ZN(n1238) );
XOR2_X1 U971 ( .A(KEYINPUT1), .B(G107), .Z(n1261) );
INV_X1 U972 ( .A(G101), .ZN(n1124) );
NAND2_X1 U973 ( .A1(KEYINPUT48), .A2(n1237), .ZN(n1260) );
INV_X1 U974 ( .A(G104), .ZN(n1237) );
NOR3_X1 U975 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1256) );
AND2_X1 U976 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NOR3_X1 U977 ( .A1(n1266), .A2(KEYINPUT3), .A3(n1265), .ZN(n1263) );
OR2_X1 U978 ( .A1(KEYINPUT35), .A2(n1267), .ZN(n1265) );
XNOR2_X1 U979 ( .A(n1268), .B(n1269), .ZN(n1266) );
XNOR2_X1 U980 ( .A(KEYINPUT10), .B(n1148), .ZN(n1269) );
INV_X1 U981 ( .A(G125), .ZN(n1148) );
NAND2_X1 U982 ( .A1(KEYINPUT17), .A2(n1149), .ZN(n1268) );
AND2_X1 U983 ( .A1(n1267), .A2(KEYINPUT3), .ZN(n1262) );
XOR2_X1 U984 ( .A(n1146), .B(KEYINPUT11), .Z(n1267) );
NOR2_X1 U985 ( .A1(n1082), .A2(G953), .ZN(n1146) );
INV_X1 U986 ( .A(G224), .ZN(n1082) );
XNOR2_X1 U987 ( .A(n1006), .B(KEYINPUT8), .ZN(n1211) );
AND2_X1 U988 ( .A1(G214), .A2(n1254), .ZN(n1006) );
NAND2_X1 U989 ( .A1(n1270), .A2(n1158), .ZN(n1254) );
INV_X1 U990 ( .A(G237), .ZN(n1270) );
XNOR2_X1 U991 ( .A(n1271), .B(G472), .ZN(n1009) );
NAND2_X1 U992 ( .A1(n1272), .A2(n1158), .ZN(n1271) );
XOR2_X1 U993 ( .A(n1120), .B(n1273), .Z(n1272) );
XNOR2_X1 U994 ( .A(G101), .B(n1125), .ZN(n1273) );
NAND2_X1 U995 ( .A1(G210), .A2(n1274), .ZN(n1125) );
XNOR2_X1 U996 ( .A(n1239), .B(n1275), .ZN(n1120) );
XOR2_X1 U997 ( .A(n1091), .B(n1149), .Z(n1275) );
XNOR2_X1 U998 ( .A(n1276), .B(n1214), .ZN(n1149) );
NAND2_X1 U999 ( .A1(n1277), .A2(KEYINPUT26), .ZN(n1276) );
XNOR2_X1 U1000 ( .A(n1278), .B(n1244), .ZN(n1277) );
NAND2_X1 U1001 ( .A1(KEYINPUT37), .A2(n1247), .ZN(n1278) );
INV_X1 U1002 ( .A(G146), .ZN(n1247) );
XNOR2_X1 U1003 ( .A(G113), .B(n1279), .ZN(n1091) );
XNOR2_X1 U1004 ( .A(G119), .B(n1223), .ZN(n1279) );
XNOR2_X1 U1005 ( .A(n1280), .B(n1281), .ZN(n1239) );
NOR2_X1 U1006 ( .A1(KEYINPUT16), .A2(n1075), .ZN(n1281) );
XOR2_X1 U1007 ( .A(G134), .B(KEYINPUT46), .Z(n1075) );
XNOR2_X1 U1008 ( .A(G137), .B(G131), .ZN(n1280) );
NAND2_X1 U1009 ( .A1(n1226), .A2(n1224), .ZN(n1196) );
XNOR2_X1 U1010 ( .A(n1018), .B(G475), .ZN(n1224) );
AND2_X1 U1011 ( .A1(n1282), .A2(n1112), .ZN(n1018) );
XNOR2_X1 U1012 ( .A(n1283), .B(n1284), .ZN(n1112) );
XOR2_X1 U1013 ( .A(KEYINPUT38), .B(n1285), .Z(n1284) );
NOR2_X1 U1014 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U1015 ( .A(n1288), .B(KEYINPUT4), .Z(n1287) );
NAND2_X1 U1016 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XNOR2_X1 U1017 ( .A(G131), .B(KEYINPUT22), .ZN(n1289) );
NOR2_X1 U1018 ( .A1(G131), .A2(n1290), .ZN(n1286) );
XNOR2_X1 U1019 ( .A(n1291), .B(n1244), .ZN(n1290) );
NAND2_X1 U1020 ( .A1(G214), .A2(n1274), .ZN(n1291) );
NOR2_X1 U1021 ( .A1(G953), .A2(G237), .ZN(n1274) );
XOR2_X1 U1022 ( .A(n1292), .B(n1293), .Z(n1283) );
NAND2_X1 U1023 ( .A1(n1294), .A2(n1295), .ZN(n1292) );
OR2_X1 U1024 ( .A1(n1296), .A2(G104), .ZN(n1295) );
XOR2_X1 U1025 ( .A(n1297), .B(KEYINPUT30), .Z(n1294) );
NAND2_X1 U1026 ( .A1(G104), .A2(n1296), .ZN(n1297) );
XOR2_X1 U1027 ( .A(G113), .B(G122), .Z(n1296) );
XNOR2_X1 U1028 ( .A(KEYINPUT7), .B(n1158), .ZN(n1282) );
INV_X1 U1029 ( .A(n1017), .ZN(n1226) );
XNOR2_X1 U1030 ( .A(n1298), .B(G478), .ZN(n1017) );
OR2_X1 U1031 ( .A1(n1107), .A2(G902), .ZN(n1298) );
XNOR2_X1 U1032 ( .A(n1299), .B(n1300), .ZN(n1107) );
XNOR2_X1 U1033 ( .A(n1214), .B(n1301), .ZN(n1300) );
XNOR2_X1 U1034 ( .A(n1244), .B(G134), .ZN(n1301) );
INV_X1 U1035 ( .A(G143), .ZN(n1244) );
XOR2_X1 U1036 ( .A(n1302), .B(n1303), .Z(n1299) );
AND2_X1 U1037 ( .A1(n1304), .A2(G217), .ZN(n1303) );
NAND2_X1 U1038 ( .A1(KEYINPUT19), .A2(n1305), .ZN(n1302) );
XOR2_X1 U1039 ( .A(G107), .B(n1306), .Z(n1305) );
NOR2_X1 U1040 ( .A1(KEYINPUT63), .A2(n1307), .ZN(n1306) );
XNOR2_X1 U1041 ( .A(G122), .B(n1223), .ZN(n1307) );
INV_X1 U1042 ( .A(G116), .ZN(n1223) );
XNOR2_X1 U1043 ( .A(n1308), .B(n1309), .ZN(n1033) );
XOR2_X1 U1044 ( .A(KEYINPUT21), .B(n1011), .Z(n1309) );
AND2_X1 U1045 ( .A1(G217), .A2(n1228), .ZN(n1011) );
NAND2_X1 U1046 ( .A1(G234), .A2(n1158), .ZN(n1228) );
NAND2_X1 U1047 ( .A1(KEYINPUT34), .A2(n1012), .ZN(n1308) );
NAND2_X1 U1048 ( .A1(n1102), .A2(n1158), .ZN(n1012) );
INV_X1 U1049 ( .A(G902), .ZN(n1158) );
XOR2_X1 U1050 ( .A(n1310), .B(n1311), .Z(n1102) );
XNOR2_X1 U1051 ( .A(KEYINPUT2), .B(n1207), .ZN(n1311) );
INV_X1 U1052 ( .A(G137), .ZN(n1207) );
XOR2_X1 U1053 ( .A(n1312), .B(n1313), .Z(n1310) );
NOR2_X1 U1054 ( .A1(KEYINPUT25), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1055 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1056 ( .A(n1214), .B(G119), .ZN(n1316) );
INV_X1 U1057 ( .A(G128), .ZN(n1214) );
XNOR2_X1 U1058 ( .A(n1293), .B(G110), .ZN(n1315) );
XOR2_X1 U1059 ( .A(G146), .B(n1057), .Z(n1293) );
XOR2_X1 U1060 ( .A(G125), .B(G140), .Z(n1057) );
NAND2_X1 U1061 ( .A1(G221), .A2(n1304), .ZN(n1312) );
AND2_X1 U1062 ( .A1(G234), .A2(n1001), .ZN(n1304) );
INV_X1 U1063 ( .A(G953), .ZN(n1001) );
endmodule


