//Key = 0000100010000000010001110000100101011110011111110011100100001010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
n1467, n1468, n1469;

XNOR2_X1 U809 ( .A(n1117), .B(n1118), .ZN(G9) );
NOR4_X1 U810 ( .A1(KEYINPUT58), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1118) );
NOR2_X1 U811 ( .A1(n1122), .A2(n1123), .ZN(G75) );
NOR4_X1 U812 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1123) );
NOR2_X1 U813 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NOR2_X1 U814 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
NOR4_X1 U815 ( .A1(n1132), .A2(n1133), .A3(n1119), .A4(n1134), .ZN(n1131) );
NOR2_X1 U816 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NOR2_X1 U817 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR3_X1 U818 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1138) );
NOR2_X1 U819 ( .A1(n1142), .A2(n1143), .ZN(n1137) );
NOR2_X1 U820 ( .A1(n1144), .A2(n1145), .ZN(n1132) );
NOR2_X1 U821 ( .A1(n1146), .A2(n1139), .ZN(n1144) );
NOR4_X1 U822 ( .A1(n1135), .A2(n1147), .A3(n1146), .A4(n1139), .ZN(n1130) );
NOR3_X1 U823 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1147) );
NOR2_X1 U824 ( .A1(n1151), .A2(n1134), .ZN(n1150) );
NOR2_X1 U825 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NOR3_X1 U826 ( .A1(n1154), .A2(n1119), .A3(n1155), .ZN(n1149) );
NOR2_X1 U827 ( .A1(n1156), .A2(n1157), .ZN(n1148) );
XNOR2_X1 U828 ( .A(n1158), .B(KEYINPUT0), .ZN(n1156) );
NAND3_X1 U829 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1124) );
NOR3_X1 U830 ( .A1(n1162), .A2(G953), .A3(G952), .ZN(n1122) );
INV_X1 U831 ( .A(n1159), .ZN(n1162) );
NAND4_X1 U832 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1159) );
NOR4_X1 U833 ( .A1(n1167), .A2(n1168), .A3(n1135), .A4(n1169), .ZN(n1166) );
NOR2_X1 U834 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NOR2_X1 U835 ( .A1(G478), .A2(n1172), .ZN(n1171) );
NOR2_X1 U836 ( .A1(n1173), .A2(KEYINPUT53), .ZN(n1172) );
NOR2_X1 U837 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NOR2_X1 U838 ( .A1(n1176), .A2(n1177), .ZN(n1170) );
INV_X1 U839 ( .A(n1174), .ZN(n1177) );
NOR2_X1 U840 ( .A1(n1178), .A2(n1175), .ZN(n1176) );
INV_X1 U841 ( .A(KEYINPUT37), .ZN(n1175) );
NOR2_X1 U842 ( .A1(KEYINPUT53), .A2(n1179), .ZN(n1178) );
INV_X1 U843 ( .A(n1180), .ZN(n1168) );
NOR2_X1 U844 ( .A1(n1134), .A2(n1181), .ZN(n1165) );
XNOR2_X1 U845 ( .A(G469), .B(n1182), .ZN(n1164) );
NAND2_X1 U846 ( .A1(KEYINPUT42), .A2(n1183), .ZN(n1182) );
NAND2_X1 U847 ( .A1(n1184), .A2(n1185), .ZN(G72) );
NAND4_X1 U848 ( .A1(G953), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1185) );
NAND2_X1 U849 ( .A1(n1189), .A2(n1190), .ZN(n1184) );
NAND2_X1 U850 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NAND3_X1 U851 ( .A1(n1193), .A2(n1186), .A3(G953), .ZN(n1192) );
NAND2_X1 U852 ( .A1(n1188), .A2(n1194), .ZN(n1193) );
INV_X1 U853 ( .A(KEYINPUT18), .ZN(n1188) );
NAND2_X1 U854 ( .A1(n1194), .A2(n1195), .ZN(n1191) );
NAND2_X1 U855 ( .A1(G953), .A2(n1186), .ZN(n1195) );
NAND2_X1 U856 ( .A1(G900), .A2(G227), .ZN(n1186) );
INV_X1 U857 ( .A(KEYINPUT20), .ZN(n1194) );
NAND2_X1 U858 ( .A1(n1196), .A2(n1187), .ZN(n1189) );
NAND3_X1 U859 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1187) );
XOR2_X1 U860 ( .A(n1200), .B(n1201), .Z(n1199) );
NAND2_X1 U861 ( .A1(G953), .A2(n1202), .ZN(n1198) );
NAND2_X1 U862 ( .A1(n1203), .A2(n1160), .ZN(n1197) );
NAND3_X1 U863 ( .A1(n1203), .A2(n1160), .A3(n1204), .ZN(n1196) );
XNOR2_X1 U864 ( .A(n1201), .B(n1200), .ZN(n1204) );
NOR2_X1 U865 ( .A1(KEYINPUT3), .A2(n1205), .ZN(n1200) );
XOR2_X1 U866 ( .A(n1206), .B(n1207), .Z(n1205) );
XNOR2_X1 U867 ( .A(G131), .B(n1208), .ZN(n1206) );
XNOR2_X1 U868 ( .A(n1209), .B(KEYINPUT45), .ZN(n1201) );
NAND4_X1 U869 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1209) );
OR2_X1 U870 ( .A1(n1214), .A2(KEYINPUT19), .ZN(n1213) );
NAND2_X1 U871 ( .A1(KEYINPUT19), .A2(G125), .ZN(n1212) );
OR2_X1 U872 ( .A1(G140), .A2(KEYINPUT31), .ZN(n1211) );
NAND2_X1 U873 ( .A1(KEYINPUT31), .A2(n1215), .ZN(n1210) );
NAND2_X1 U874 ( .A1(n1216), .A2(n1217), .ZN(n1203) );
XNOR2_X1 U875 ( .A(n1218), .B(KEYINPUT30), .ZN(n1216) );
NAND2_X1 U876 ( .A1(n1219), .A2(n1220), .ZN(G69) );
NAND2_X1 U877 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NAND2_X1 U878 ( .A1(G953), .A2(n1223), .ZN(n1222) );
NAND3_X1 U879 ( .A1(n1224), .A2(n1225), .A3(G953), .ZN(n1219) );
NAND2_X1 U880 ( .A1(G898), .A2(G224), .ZN(n1225) );
XOR2_X1 U881 ( .A(KEYINPUT43), .B(n1221), .Z(n1224) );
XNOR2_X1 U882 ( .A(n1226), .B(n1227), .ZN(n1221) );
NOR2_X1 U883 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
XOR2_X1 U884 ( .A(n1230), .B(n1231), .Z(n1229) );
NOR2_X1 U885 ( .A1(KEYINPUT63), .A2(n1232), .ZN(n1230) );
NOR2_X1 U886 ( .A1(G898), .A2(n1160), .ZN(n1228) );
NAND2_X1 U887 ( .A1(n1160), .A2(n1233), .ZN(n1226) );
NAND3_X1 U888 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
NOR2_X1 U889 ( .A1(n1237), .A2(n1238), .ZN(G66) );
XNOR2_X1 U890 ( .A(n1239), .B(n1240), .ZN(n1238) );
AND2_X1 U891 ( .A1(G217), .A2(n1241), .ZN(n1239) );
NOR2_X1 U892 ( .A1(n1237), .A2(n1242), .ZN(G63) );
NOR3_X1 U893 ( .A1(n1174), .A2(n1243), .A3(n1244), .ZN(n1242) );
AND3_X1 U894 ( .A1(n1245), .A2(G478), .A3(n1241), .ZN(n1244) );
NOR2_X1 U895 ( .A1(n1246), .A2(n1245), .ZN(n1243) );
NOR2_X1 U896 ( .A1(n1247), .A2(n1179), .ZN(n1246) );
NOR2_X1 U897 ( .A1(n1237), .A2(n1248), .ZN(G60) );
XOR2_X1 U898 ( .A(n1249), .B(n1250), .Z(n1248) );
NAND2_X1 U899 ( .A1(KEYINPUT62), .A2(n1251), .ZN(n1250) );
NAND2_X1 U900 ( .A1(n1241), .A2(G475), .ZN(n1249) );
XNOR2_X1 U901 ( .A(n1252), .B(n1253), .ZN(G6) );
NOR2_X1 U902 ( .A1(n1237), .A2(n1254), .ZN(G57) );
XOR2_X1 U903 ( .A(n1255), .B(n1256), .Z(n1254) );
XOR2_X1 U904 ( .A(n1257), .B(n1258), .Z(n1256) );
NAND2_X1 U905 ( .A1(n1241), .A2(G472), .ZN(n1257) );
XOR2_X1 U906 ( .A(n1259), .B(n1260), .Z(n1255) );
NOR2_X1 U907 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U908 ( .A(n1263), .B(KEYINPUT50), .Z(n1262) );
NAND3_X1 U909 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1263) );
NAND2_X1 U910 ( .A1(n1267), .A2(n1268), .ZN(n1264) );
XNOR2_X1 U911 ( .A(KEYINPUT25), .B(n1269), .ZN(n1268) );
NOR2_X1 U912 ( .A1(n1270), .A2(n1266), .ZN(n1261) );
NOR3_X1 U913 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1270) );
NOR3_X1 U914 ( .A1(n1269), .A2(KEYINPUT25), .A3(n1274), .ZN(n1273) );
AND2_X1 U915 ( .A1(n1269), .A2(KEYINPUT25), .ZN(n1272) );
NOR2_X1 U916 ( .A1(n1275), .A2(n1276), .ZN(G54) );
XOR2_X1 U917 ( .A(KEYINPUT14), .B(n1277), .Z(n1276) );
NOR2_X1 U918 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NOR2_X1 U919 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
XOR2_X1 U920 ( .A(n1282), .B(KEYINPUT13), .Z(n1281) );
AND2_X1 U921 ( .A1(n1282), .A2(n1280), .ZN(n1278) );
XNOR2_X1 U922 ( .A(n1283), .B(n1284), .ZN(n1280) );
XNOR2_X1 U923 ( .A(n1285), .B(n1286), .ZN(n1283) );
NOR2_X1 U924 ( .A1(KEYINPUT9), .A2(n1287), .ZN(n1286) );
XOR2_X1 U925 ( .A(n1269), .B(n1288), .Z(n1287) );
NOR2_X1 U926 ( .A1(KEYINPUT48), .A2(n1289), .ZN(n1285) );
XNOR2_X1 U927 ( .A(G110), .B(G140), .ZN(n1289) );
NAND2_X1 U928 ( .A1(n1241), .A2(G469), .ZN(n1282) );
NOR2_X1 U929 ( .A1(G952), .A2(n1290), .ZN(n1275) );
XNOR2_X1 U930 ( .A(KEYINPUT17), .B(n1160), .ZN(n1290) );
NOR2_X1 U931 ( .A1(n1291), .A2(n1292), .ZN(G51) );
XOR2_X1 U932 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U933 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U934 ( .A(n1297), .B(n1298), .Z(n1293) );
NOR2_X1 U935 ( .A1(KEYINPUT6), .A2(n1267), .ZN(n1298) );
INV_X1 U936 ( .A(n1274), .ZN(n1267) );
NAND2_X1 U937 ( .A1(n1241), .A2(n1299), .ZN(n1297) );
NOR2_X1 U938 ( .A1(n1300), .A2(n1247), .ZN(n1241) );
AND3_X1 U939 ( .A1(n1301), .A2(n1161), .A3(n1217), .ZN(n1247) );
INV_X1 U940 ( .A(n1127), .ZN(n1217) );
NAND4_X1 U941 ( .A1(n1302), .A2(n1303), .A3(n1304), .A4(n1305), .ZN(n1127) );
AND4_X1 U942 ( .A1(n1306), .A2(n1307), .A3(n1308), .A4(n1309), .ZN(n1305) );
NOR2_X1 U943 ( .A1(n1310), .A2(n1311), .ZN(n1304) );
NOR2_X1 U944 ( .A1(KEYINPUT26), .A2(n1312), .ZN(n1311) );
NOR2_X1 U945 ( .A1(n1157), .A2(n1313), .ZN(n1310) );
NAND4_X1 U946 ( .A1(n1314), .A2(n1142), .A3(KEYINPUT26), .A4(n1134), .ZN(n1303) );
NAND4_X1 U947 ( .A1(n1141), .A2(n1315), .A3(n1316), .A4(n1317), .ZN(n1302) );
XOR2_X1 U948 ( .A(KEYINPUT27), .B(n1153), .Z(n1315) );
XNOR2_X1 U949 ( .A(KEYINPUT56), .B(n1125), .ZN(n1301) );
NAND3_X1 U950 ( .A1(n1318), .A2(n1236), .A3(n1319), .ZN(n1125) );
XNOR2_X1 U951 ( .A(n1234), .B(KEYINPUT60), .ZN(n1319) );
NOR4_X1 U952 ( .A1(n1320), .A2(n1321), .A3(n1322), .A4(n1323), .ZN(n1234) );
AND4_X1 U953 ( .A1(n1324), .A2(n1325), .A3(n1181), .A4(n1326), .ZN(n1320) );
XNOR2_X1 U954 ( .A(n1142), .B(KEYINPUT46), .ZN(n1324) );
NOR3_X1 U955 ( .A1(n1253), .A2(n1327), .A3(n1328), .ZN(n1236) );
NOR3_X1 U956 ( .A1(n1120), .A2(n1119), .A3(n1121), .ZN(n1328) );
AND3_X1 U957 ( .A1(n1329), .A2(n1158), .A3(n1140), .ZN(n1253) );
XOR2_X1 U958 ( .A(n1235), .B(KEYINPUT61), .Z(n1318) );
XNOR2_X1 U959 ( .A(n1237), .B(KEYINPUT36), .ZN(n1291) );
NOR2_X1 U960 ( .A1(n1160), .A2(G952), .ZN(n1237) );
XNOR2_X1 U961 ( .A(G146), .B(n1308), .ZN(G48) );
NAND3_X1 U962 ( .A1(n1140), .A2(n1330), .A3(n1314), .ZN(n1308) );
NAND3_X1 U963 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(G45) );
OR2_X1 U964 ( .A1(n1218), .A2(KEYINPUT35), .ZN(n1333) );
NAND3_X1 U965 ( .A1(KEYINPUT35), .A2(n1218), .A3(n1334), .ZN(n1332) );
NAND2_X1 U966 ( .A1(G143), .A2(n1335), .ZN(n1331) );
NAND2_X1 U967 ( .A1(n1336), .A2(KEYINPUT35), .ZN(n1335) );
XNOR2_X1 U968 ( .A(n1218), .B(KEYINPUT47), .ZN(n1336) );
INV_X1 U969 ( .A(n1161), .ZN(n1218) );
NAND3_X1 U970 ( .A1(n1153), .A2(n1316), .A3(n1337), .ZN(n1161) );
NOR3_X1 U971 ( .A1(n1157), .A2(n1163), .A3(n1338), .ZN(n1337) );
XNOR2_X1 U972 ( .A(n1339), .B(n1340), .ZN(G42) );
NOR2_X1 U973 ( .A1(KEYINPUT7), .A2(n1309), .ZN(n1340) );
NAND4_X1 U974 ( .A1(n1140), .A2(n1152), .A3(n1316), .A4(n1317), .ZN(n1309) );
XNOR2_X1 U975 ( .A(G137), .B(n1312), .ZN(G39) );
NAND3_X1 U976 ( .A1(n1142), .A2(n1317), .A3(n1314), .ZN(n1312) );
XNOR2_X1 U977 ( .A(G134), .B(n1341), .ZN(G36) );
NAND2_X1 U978 ( .A1(n1342), .A2(n1317), .ZN(n1341) );
XOR2_X1 U979 ( .A(n1343), .B(KEYINPUT41), .Z(n1342) );
NAND3_X1 U980 ( .A1(n1316), .A2(n1141), .A3(n1153), .ZN(n1343) );
XNOR2_X1 U981 ( .A(G131), .B(n1307), .ZN(G33) );
NAND4_X1 U982 ( .A1(n1140), .A2(n1153), .A3(n1316), .A4(n1317), .ZN(n1307) );
INV_X1 U983 ( .A(n1134), .ZN(n1317) );
NAND2_X1 U984 ( .A1(n1344), .A2(n1154), .ZN(n1134) );
INV_X1 U985 ( .A(n1155), .ZN(n1344) );
XNOR2_X1 U986 ( .A(G128), .B(n1306), .ZN(G30) );
NAND3_X1 U987 ( .A1(n1141), .A2(n1330), .A3(n1314), .ZN(n1306) );
AND3_X1 U988 ( .A1(n1181), .A2(n1326), .A3(n1316), .ZN(n1314) );
NOR3_X1 U989 ( .A1(n1135), .A2(n1143), .A3(n1345), .ZN(n1316) );
XNOR2_X1 U990 ( .A(G101), .B(n1235), .ZN(G3) );
NAND3_X1 U991 ( .A1(n1153), .A2(n1329), .A3(n1142), .ZN(n1235) );
INV_X1 U992 ( .A(n1146), .ZN(n1142) );
INV_X1 U993 ( .A(n1121), .ZN(n1329) );
XOR2_X1 U994 ( .A(n1346), .B(n1347), .Z(G27) );
XNOR2_X1 U995 ( .A(KEYINPUT51), .B(n1348), .ZN(n1347) );
NAND2_X1 U996 ( .A1(n1349), .A2(n1330), .ZN(n1346) );
XOR2_X1 U997 ( .A(n1313), .B(KEYINPUT21), .Z(n1349) );
NAND3_X1 U998 ( .A1(n1143), .A2(n1140), .A3(n1350), .ZN(n1313) );
NOR3_X1 U999 ( .A1(n1351), .A2(n1135), .A3(n1345), .ZN(n1350) );
AND2_X1 U1000 ( .A1(n1129), .A2(n1352), .ZN(n1345) );
NAND4_X1 U1001 ( .A1(G953), .A2(G902), .A3(n1353), .A4(n1202), .ZN(n1352) );
INV_X1 U1002 ( .A(G900), .ZN(n1202) );
INV_X1 U1003 ( .A(n1145), .ZN(n1135) );
XOR2_X1 U1004 ( .A(G122), .B(n1321), .Z(G24) );
NOR4_X1 U1005 ( .A1(n1354), .A2(n1119), .A3(n1338), .A4(n1163), .ZN(n1321) );
INV_X1 U1006 ( .A(n1158), .ZN(n1119) );
NOR2_X1 U1007 ( .A1(n1326), .A2(n1181), .ZN(n1158) );
XOR2_X1 U1008 ( .A(G119), .B(n1355), .Z(G21) );
NOR4_X1 U1009 ( .A1(n1356), .A2(n1357), .A3(n1146), .A4(n1354), .ZN(n1355) );
XNOR2_X1 U1010 ( .A(n1358), .B(n1322), .ZN(G18) );
AND3_X1 U1011 ( .A1(n1153), .A2(n1141), .A3(n1325), .ZN(n1322) );
INV_X1 U1012 ( .A(n1120), .ZN(n1141) );
NAND2_X1 U1013 ( .A1(n1163), .A2(n1359), .ZN(n1120) );
XOR2_X1 U1014 ( .A(G113), .B(n1323), .Z(G15) );
AND3_X1 U1015 ( .A1(n1140), .A2(n1153), .A3(n1325), .ZN(n1323) );
INV_X1 U1016 ( .A(n1354), .ZN(n1325) );
NAND3_X1 U1017 ( .A1(n1360), .A2(n1145), .A3(n1143), .ZN(n1354) );
INV_X1 U1018 ( .A(n1139), .ZN(n1143) );
NOR2_X1 U1019 ( .A1(n1326), .A2(n1357), .ZN(n1153) );
INV_X1 U1020 ( .A(n1181), .ZN(n1357) );
NOR2_X1 U1021 ( .A1(n1359), .A2(n1163), .ZN(n1140) );
XNOR2_X1 U1022 ( .A(n1361), .B(n1327), .ZN(G12) );
NOR3_X1 U1023 ( .A1(n1351), .A2(n1121), .A3(n1146), .ZN(n1327) );
NAND2_X1 U1024 ( .A1(n1338), .A2(n1163), .ZN(n1146) );
XOR2_X1 U1025 ( .A(n1362), .B(G475), .Z(n1163) );
OR2_X1 U1026 ( .A1(n1251), .A2(G902), .ZN(n1362) );
XNOR2_X1 U1027 ( .A(n1363), .B(n1364), .ZN(n1251) );
XNOR2_X1 U1028 ( .A(G113), .B(n1252), .ZN(n1364) );
INV_X1 U1029 ( .A(G104), .ZN(n1252) );
XOR2_X1 U1030 ( .A(n1365), .B(n1366), .Z(n1363) );
NAND3_X1 U1031 ( .A1(n1367), .A2(n1368), .A3(n1369), .ZN(n1365) );
NAND2_X1 U1032 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
NAND2_X1 U1033 ( .A1(KEYINPUT11), .A2(n1372), .ZN(n1368) );
NAND2_X1 U1034 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
XNOR2_X1 U1035 ( .A(n1371), .B(KEYINPUT59), .ZN(n1373) );
NAND2_X1 U1036 ( .A1(n1375), .A2(n1376), .ZN(n1367) );
INV_X1 U1037 ( .A(KEYINPUT11), .ZN(n1376) );
NAND2_X1 U1038 ( .A1(n1377), .A2(n1378), .ZN(n1375) );
OR3_X1 U1039 ( .A1(n1370), .A2(n1371), .A3(KEYINPUT59), .ZN(n1378) );
INV_X1 U1040 ( .A(n1374), .ZN(n1370) );
XNOR2_X1 U1041 ( .A(n1379), .B(n1380), .ZN(n1374) );
AND3_X1 U1042 ( .A1(G214), .A2(n1160), .A3(n1381), .ZN(n1380) );
XNOR2_X1 U1043 ( .A(G131), .B(G143), .ZN(n1379) );
NAND2_X1 U1044 ( .A1(KEYINPUT59), .A2(n1371), .ZN(n1377) );
XNOR2_X1 U1045 ( .A(n1382), .B(n1383), .ZN(n1371) );
NOR2_X1 U1046 ( .A1(G146), .A2(KEYINPUT15), .ZN(n1383) );
NAND3_X1 U1047 ( .A1(n1384), .A2(n1385), .A3(n1386), .ZN(n1382) );
OR2_X1 U1048 ( .A1(n1348), .A2(KEYINPUT33), .ZN(n1385) );
NAND2_X1 U1049 ( .A1(n1387), .A2(KEYINPUT33), .ZN(n1384) );
INV_X1 U1050 ( .A(n1359), .ZN(n1338) );
XNOR2_X1 U1051 ( .A(n1174), .B(n1179), .ZN(n1359) );
INV_X1 U1052 ( .A(G478), .ZN(n1179) );
NOR2_X1 U1053 ( .A1(n1245), .A2(G902), .ZN(n1174) );
XNOR2_X1 U1054 ( .A(n1388), .B(n1389), .ZN(n1245) );
XOR2_X1 U1055 ( .A(n1390), .B(n1391), .Z(n1389) );
XNOR2_X1 U1056 ( .A(G134), .B(n1392), .ZN(n1391) );
XNOR2_X1 U1057 ( .A(KEYINPUT57), .B(n1334), .ZN(n1390) );
XOR2_X1 U1058 ( .A(n1393), .B(n1394), .Z(n1388) );
XNOR2_X1 U1059 ( .A(n1358), .B(G107), .ZN(n1394) );
XOR2_X1 U1060 ( .A(n1395), .B(n1366), .Z(n1393) );
NAND2_X1 U1061 ( .A1(G217), .A2(n1396), .ZN(n1395) );
NAND3_X1 U1062 ( .A1(n1145), .A2(n1139), .A3(n1360), .ZN(n1121) );
AND2_X1 U1063 ( .A1(n1330), .A2(n1397), .ZN(n1360) );
NAND2_X1 U1064 ( .A1(n1129), .A2(n1398), .ZN(n1397) );
NAND4_X1 U1065 ( .A1(G953), .A2(G902), .A3(n1353), .A4(n1399), .ZN(n1398) );
INV_X1 U1066 ( .A(G898), .ZN(n1399) );
NAND3_X1 U1067 ( .A1(n1353), .A2(n1160), .A3(G952), .ZN(n1129) );
NAND2_X1 U1068 ( .A1(G237), .A2(n1400), .ZN(n1353) );
XOR2_X1 U1069 ( .A(KEYINPUT49), .B(G234), .Z(n1400) );
INV_X1 U1070 ( .A(n1157), .ZN(n1330) );
NAND2_X1 U1071 ( .A1(n1155), .A2(n1154), .ZN(n1157) );
NAND2_X1 U1072 ( .A1(G214), .A2(n1401), .ZN(n1154) );
XNOR2_X1 U1073 ( .A(n1402), .B(n1299), .ZN(n1155) );
AND2_X1 U1074 ( .A1(G210), .A2(n1401), .ZN(n1299) );
NAND2_X1 U1075 ( .A1(n1381), .A2(n1300), .ZN(n1401) );
NAND2_X1 U1076 ( .A1(n1403), .A2(n1300), .ZN(n1402) );
XOR2_X1 U1077 ( .A(n1404), .B(n1296), .Z(n1403) );
XNOR2_X1 U1078 ( .A(n1348), .B(n1405), .ZN(n1296) );
NOR2_X1 U1079 ( .A1(G953), .A2(n1223), .ZN(n1405) );
INV_X1 U1080 ( .A(G224), .ZN(n1223) );
XNOR2_X1 U1081 ( .A(n1274), .B(n1406), .ZN(n1404) );
NOR2_X1 U1082 ( .A1(KEYINPUT54), .A2(n1295), .ZN(n1406) );
XOR2_X1 U1083 ( .A(n1231), .B(n1232), .Z(n1295) );
XNOR2_X1 U1084 ( .A(G110), .B(n1366), .ZN(n1232) );
XOR2_X1 U1085 ( .A(G122), .B(KEYINPUT52), .Z(n1366) );
XNOR2_X1 U1086 ( .A(n1407), .B(n1408), .ZN(n1231) );
XOR2_X1 U1087 ( .A(KEYINPUT22), .B(G113), .Z(n1408) );
XNOR2_X1 U1088 ( .A(n1409), .B(n1117), .ZN(n1407) );
NAND3_X1 U1089 ( .A1(n1410), .A2(n1411), .A3(n1412), .ZN(n1409) );
NAND2_X1 U1090 ( .A1(n1413), .A2(n1414), .ZN(n1412) );
OR3_X1 U1091 ( .A1(n1414), .A2(G116), .A3(G119), .ZN(n1411) );
NAND2_X1 U1092 ( .A1(G119), .A2(n1415), .ZN(n1410) );
XNOR2_X1 U1093 ( .A(n1414), .B(n1358), .ZN(n1415) );
NAND2_X1 U1094 ( .A1(n1416), .A2(n1417), .ZN(n1139) );
NAND2_X1 U1095 ( .A1(G469), .A2(n1183), .ZN(n1417) );
XOR2_X1 U1096 ( .A(n1418), .B(KEYINPUT10), .Z(n1416) );
OR2_X1 U1097 ( .A1(n1183), .A2(G469), .ZN(n1418) );
NAND3_X1 U1098 ( .A1(n1419), .A2(n1420), .A3(n1300), .ZN(n1183) );
NAND2_X1 U1099 ( .A1(n1421), .A2(n1422), .ZN(n1420) );
XOR2_X1 U1100 ( .A(n1423), .B(n1424), .Z(n1421) );
OR3_X1 U1101 ( .A1(n1423), .A2(n1424), .A3(n1422), .ZN(n1419) );
INV_X1 U1102 ( .A(KEYINPUT32), .ZN(n1422) );
XOR2_X1 U1103 ( .A(n1425), .B(n1426), .Z(n1424) );
NOR2_X1 U1104 ( .A1(KEYINPUT40), .A2(n1284), .ZN(n1426) );
NAND2_X1 U1105 ( .A1(G227), .A2(n1160), .ZN(n1284) );
XNOR2_X1 U1106 ( .A(n1427), .B(n1339), .ZN(n1425) );
NAND2_X1 U1107 ( .A1(KEYINPUT38), .A2(n1361), .ZN(n1427) );
NAND2_X1 U1108 ( .A1(n1428), .A2(n1429), .ZN(n1423) );
NAND2_X1 U1109 ( .A1(n1288), .A2(n1269), .ZN(n1429) );
XOR2_X1 U1110 ( .A(KEYINPUT4), .B(n1430), .Z(n1428) );
NOR2_X1 U1111 ( .A1(n1288), .A2(n1269), .ZN(n1430) );
XOR2_X1 U1112 ( .A(n1431), .B(n1207), .Z(n1288) );
XNOR2_X1 U1113 ( .A(n1392), .B(n1432), .ZN(n1207) );
NOR2_X1 U1114 ( .A1(n1433), .A2(n1434), .ZN(n1432) );
NOR2_X1 U1115 ( .A1(KEYINPUT34), .A2(n1435), .ZN(n1434) );
AND2_X1 U1116 ( .A1(KEYINPUT24), .A2(n1435), .ZN(n1433) );
NAND2_X1 U1117 ( .A1(n1436), .A2(n1437), .ZN(n1431) );
NAND2_X1 U1118 ( .A1(G107), .A2(n1414), .ZN(n1437) );
NAND2_X1 U1119 ( .A1(n1438), .A2(n1117), .ZN(n1436) );
INV_X1 U1120 ( .A(G107), .ZN(n1117) );
XOR2_X1 U1121 ( .A(n1414), .B(KEYINPUT23), .Z(n1438) );
XNOR2_X1 U1122 ( .A(G104), .B(n1258), .ZN(n1414) );
NAND2_X1 U1123 ( .A1(G221), .A2(n1439), .ZN(n1145) );
INV_X1 U1124 ( .A(n1152), .ZN(n1351) );
NOR2_X1 U1125 ( .A1(n1181), .A2(n1356), .ZN(n1152) );
INV_X1 U1126 ( .A(n1326), .ZN(n1356) );
NAND2_X1 U1127 ( .A1(n1440), .A2(n1180), .ZN(n1326) );
NAND3_X1 U1128 ( .A1(n1441), .A2(n1300), .A3(n1240), .ZN(n1180) );
XNOR2_X1 U1129 ( .A(n1167), .B(KEYINPUT39), .ZN(n1440) );
NOR2_X1 U1130 ( .A1(n1441), .A2(n1442), .ZN(n1167) );
AND2_X1 U1131 ( .A1(n1240), .A2(n1300), .ZN(n1442) );
XOR2_X1 U1132 ( .A(n1443), .B(n1444), .Z(n1240) );
XOR2_X1 U1133 ( .A(n1445), .B(n1446), .Z(n1444) );
XOR2_X1 U1134 ( .A(n1447), .B(n1448), .Z(n1446) );
NOR2_X1 U1135 ( .A1(G119), .A2(KEYINPUT1), .ZN(n1448) );
NAND3_X1 U1136 ( .A1(n1449), .A2(n1450), .A3(n1214), .ZN(n1447) );
INV_X1 U1137 ( .A(n1387), .ZN(n1214) );
NOR2_X1 U1138 ( .A1(G125), .A2(G140), .ZN(n1387) );
NAND2_X1 U1139 ( .A1(KEYINPUT29), .A2(n1339), .ZN(n1450) );
OR2_X1 U1140 ( .A1(n1386), .A2(KEYINPUT29), .ZN(n1449) );
INV_X1 U1141 ( .A(n1215), .ZN(n1386) );
NOR2_X1 U1142 ( .A1(n1339), .A2(n1348), .ZN(n1215) );
INV_X1 U1143 ( .A(G125), .ZN(n1348) );
INV_X1 U1144 ( .A(G140), .ZN(n1339) );
NAND2_X1 U1145 ( .A1(n1396), .A2(G221), .ZN(n1445) );
AND2_X1 U1146 ( .A1(G234), .A2(n1160), .ZN(n1396) );
XOR2_X1 U1147 ( .A(n1451), .B(n1452), .Z(n1443) );
XNOR2_X1 U1148 ( .A(n1392), .B(G110), .ZN(n1452) );
XNOR2_X1 U1149 ( .A(G137), .B(G146), .ZN(n1451) );
NAND2_X1 U1150 ( .A1(G217), .A2(n1439), .ZN(n1441) );
NAND2_X1 U1151 ( .A1(G234), .A2(n1300), .ZN(n1439) );
XNOR2_X1 U1152 ( .A(n1453), .B(G472), .ZN(n1181) );
NAND2_X1 U1153 ( .A1(n1454), .A2(n1300), .ZN(n1453) );
INV_X1 U1154 ( .A(G902), .ZN(n1300) );
XOR2_X1 U1155 ( .A(n1455), .B(n1456), .Z(n1454) );
XNOR2_X1 U1156 ( .A(n1266), .B(n1258), .ZN(n1456) );
XOR2_X1 U1157 ( .A(G101), .B(KEYINPUT44), .Z(n1258) );
XNOR2_X1 U1158 ( .A(G113), .B(n1457), .ZN(n1266) );
NOR2_X1 U1159 ( .A1(n1413), .A2(n1458), .ZN(n1457) );
XOR2_X1 U1160 ( .A(n1459), .B(KEYINPUT28), .Z(n1458) );
NAND2_X1 U1161 ( .A1(n1460), .A2(n1358), .ZN(n1459) );
XOR2_X1 U1162 ( .A(KEYINPUT5), .B(G119), .Z(n1460) );
NOR2_X1 U1163 ( .A1(n1358), .A2(G119), .ZN(n1413) );
INV_X1 U1164 ( .A(G116), .ZN(n1358) );
XNOR2_X1 U1165 ( .A(n1461), .B(n1462), .ZN(n1455) );
NOR2_X1 U1166 ( .A1(KEYINPUT2), .A2(n1259), .ZN(n1462) );
NAND3_X1 U1167 ( .A1(n1381), .A2(n1160), .A3(G210), .ZN(n1259) );
INV_X1 U1168 ( .A(G953), .ZN(n1160) );
INV_X1 U1169 ( .A(G237), .ZN(n1381) );
NOR2_X1 U1170 ( .A1(KEYINPUT16), .A2(n1463), .ZN(n1461) );
NOR2_X1 U1171 ( .A1(n1464), .A2(n1271), .ZN(n1463) );
INV_X1 U1172 ( .A(n1265), .ZN(n1271) );
NAND2_X1 U1173 ( .A1(n1274), .A2(n1269), .ZN(n1265) );
NOR2_X1 U1174 ( .A1(n1274), .A2(n1269), .ZN(n1464) );
NAND2_X1 U1175 ( .A1(n1465), .A2(n1466), .ZN(n1269) );
NAND2_X1 U1176 ( .A1(G131), .A2(n1208), .ZN(n1466) );
XOR2_X1 U1177 ( .A(KEYINPUT8), .B(n1467), .Z(n1465) );
NOR2_X1 U1178 ( .A1(G131), .A2(n1208), .ZN(n1467) );
XOR2_X1 U1179 ( .A(G134), .B(G137), .Z(n1208) );
XNOR2_X1 U1180 ( .A(n1468), .B(n1435), .ZN(n1274) );
XNOR2_X1 U1181 ( .A(n1334), .B(G146), .ZN(n1435) );
INV_X1 U1182 ( .A(G143), .ZN(n1334) );
NAND2_X1 U1183 ( .A1(n1469), .A2(n1392), .ZN(n1468) );
INV_X1 U1184 ( .A(G128), .ZN(n1392) );
XOR2_X1 U1185 ( .A(KEYINPUT55), .B(KEYINPUT12), .Z(n1469) );
INV_X1 U1186 ( .A(G110), .ZN(n1361) );
endmodule


