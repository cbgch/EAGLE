//Key = 0111101011000011100010101000010100011000001110111011100001000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309;

XNOR2_X1 U719 ( .A(G107), .B(n989), .ZN(G9) );
NOR2_X1 U720 ( .A1(n990), .A2(n991), .ZN(G75) );
NOR4_X1 U721 ( .A1(G953), .A2(n992), .A3(n993), .A4(n994), .ZN(n991) );
NOR2_X1 U722 ( .A1(n995), .A2(n996), .ZN(n993) );
NOR2_X1 U723 ( .A1(n997), .A2(n998), .ZN(n995) );
NOR3_X1 U724 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n998) );
NOR3_X1 U725 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(n1001) );
NOR2_X1 U726 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NOR2_X1 U727 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR2_X1 U728 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U729 ( .A1(n1011), .A2(n1012), .ZN(n1003) );
NOR2_X1 U730 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
NOR2_X1 U731 ( .A1(n1015), .A2(n1016), .ZN(n1000) );
NOR3_X1 U732 ( .A1(n1006), .A2(n1017), .A3(n1018), .ZN(n1016) );
NOR2_X1 U733 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
XNOR2_X1 U734 ( .A(n1021), .B(KEYINPUT46), .ZN(n1020) );
NOR2_X1 U735 ( .A1(n1022), .A2(n1023), .ZN(n1017) );
NOR2_X1 U736 ( .A1(n1024), .A2(n1012), .ZN(n1022) );
INV_X1 U737 ( .A(n1025), .ZN(n999) );
NOR4_X1 U738 ( .A1(n1026), .A2(n1006), .A3(n1002), .A4(n1012), .ZN(n997) );
NOR2_X1 U739 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NOR3_X1 U740 ( .A1(n992), .A2(G953), .A3(G952), .ZN(n990) );
AND4_X1 U741 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n992) );
NOR4_X1 U742 ( .A1(n1033), .A2(n1034), .A3(n1002), .A4(n1035), .ZN(n1032) );
XNOR2_X1 U743 ( .A(KEYINPUT30), .B(n1036), .ZN(n1035) );
INV_X1 U744 ( .A(n1015), .ZN(n1002) );
NOR3_X1 U745 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1031) );
INV_X1 U746 ( .A(n1040), .ZN(n1037) );
NAND2_X1 U747 ( .A1(n1041), .A2(n1042), .ZN(n1029) );
XNOR2_X1 U748 ( .A(KEYINPUT37), .B(n1043), .ZN(n1041) );
XOR2_X1 U749 ( .A(n1044), .B(n1045), .Z(G72) );
NOR2_X1 U750 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
XOR2_X1 U751 ( .A(n1048), .B(n1049), .Z(n1047) );
XNOR2_X1 U752 ( .A(n1050), .B(n1051), .ZN(n1049) );
XNOR2_X1 U753 ( .A(KEYINPUT4), .B(n1052), .ZN(n1048) );
NOR2_X1 U754 ( .A1(KEYINPUT12), .A2(n1053), .ZN(n1052) );
XNOR2_X1 U755 ( .A(G131), .B(n1054), .ZN(n1053) );
NOR2_X1 U756 ( .A1(KEYINPUT56), .A2(n1055), .ZN(n1054) );
NOR2_X1 U757 ( .A1(G900), .A2(n1056), .ZN(n1046) );
XNOR2_X1 U758 ( .A(G953), .B(KEYINPUT38), .ZN(n1056) );
NAND2_X1 U759 ( .A1(n1057), .A2(n1058), .ZN(n1044) );
NAND2_X1 U760 ( .A1(G953), .A2(n1059), .ZN(n1058) );
NAND2_X1 U761 ( .A1(G900), .A2(G227), .ZN(n1059) );
XOR2_X1 U762 ( .A(n1060), .B(n1061), .Z(G69) );
NOR3_X1 U763 ( .A1(n1062), .A2(KEYINPUT27), .A3(n1063), .ZN(n1061) );
AND2_X1 U764 ( .A1(G224), .A2(G898), .ZN(n1063) );
NAND2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1060) );
NAND3_X1 U766 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
NAND2_X1 U767 ( .A1(G953), .A2(n1069), .ZN(n1067) );
OR2_X1 U768 ( .A1(n1068), .A2(n1066), .ZN(n1064) );
NAND2_X1 U769 ( .A1(n1062), .A2(n1070), .ZN(n1068) );
NAND2_X1 U770 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XNOR2_X1 U771 ( .A(n1073), .B(KEYINPUT31), .ZN(n1071) );
NOR2_X1 U772 ( .A1(n1074), .A2(n1075), .ZN(G66) );
XOR2_X1 U773 ( .A(n1076), .B(n1077), .Z(n1075) );
NAND3_X1 U774 ( .A1(n1078), .A2(n994), .A3(n1079), .ZN(n1076) );
XNOR2_X1 U775 ( .A(G902), .B(KEYINPUT3), .ZN(n1079) );
NOR2_X1 U776 ( .A1(n1074), .A2(n1080), .ZN(G63) );
XOR2_X1 U777 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND3_X1 U778 ( .A1(G902), .A2(n994), .A3(G478), .ZN(n1081) );
NOR2_X1 U779 ( .A1(n1074), .A2(n1083), .ZN(G60) );
NOR2_X1 U780 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XOR2_X1 U781 ( .A(KEYINPUT11), .B(n1086), .Z(n1085) );
NOR2_X1 U782 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
AND2_X1 U783 ( .A1(n1088), .A2(n1087), .ZN(n1084) );
NAND3_X1 U784 ( .A1(G475), .A2(n994), .A3(n1089), .ZN(n1088) );
XNOR2_X1 U785 ( .A(G902), .B(KEYINPUT8), .ZN(n1089) );
XNOR2_X1 U786 ( .A(G104), .B(n1090), .ZN(G6) );
NOR2_X1 U787 ( .A1(n1074), .A2(n1091), .ZN(G57) );
XOR2_X1 U788 ( .A(n1092), .B(n1093), .Z(n1091) );
XOR2_X1 U789 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U790 ( .A1(G101), .A2(KEYINPUT61), .ZN(n1094) );
XOR2_X1 U791 ( .A(n1096), .B(n1097), .Z(n1092) );
XOR2_X1 U792 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U793 ( .A1(KEYINPUT41), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U794 ( .A(n1101), .B(n1102), .ZN(n1100) );
NAND3_X1 U795 ( .A1(G472), .A2(n994), .A3(n1103), .ZN(n1096) );
XNOR2_X1 U796 ( .A(G902), .B(KEYINPUT6), .ZN(n1103) );
NOR2_X1 U797 ( .A1(n1062), .A2(G952), .ZN(n1074) );
NOR2_X1 U798 ( .A1(n1104), .A2(n1105), .ZN(G54) );
XOR2_X1 U799 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U800 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U801 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
OR2_X1 U802 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND4_X1 U803 ( .A1(n1114), .A2(n1062), .A3(G227), .A4(n1112), .ZN(n1110) );
INV_X1 U804 ( .A(KEYINPUT57), .ZN(n1112) );
NAND2_X1 U805 ( .A1(n1115), .A2(n1116), .ZN(n1108) );
NAND2_X1 U806 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U807 ( .A(n1119), .B(KEYINPUT49), .Z(n1115) );
NAND2_X1 U808 ( .A1(n1120), .A2(n1051), .ZN(n1119) );
XOR2_X1 U809 ( .A(n1121), .B(n1122), .Z(n1106) );
NOR2_X1 U810 ( .A1(KEYINPUT5), .A2(n1123), .ZN(n1122) );
XNOR2_X1 U811 ( .A(n1102), .B(KEYINPUT47), .ZN(n1123) );
XOR2_X1 U812 ( .A(n1124), .B(KEYINPUT20), .Z(n1121) );
NAND3_X1 U813 ( .A1(G902), .A2(n994), .A3(G469), .ZN(n1124) );
NOR2_X1 U814 ( .A1(G952), .A2(n1125), .ZN(n1104) );
XNOR2_X1 U815 ( .A(G953), .B(KEYINPUT19), .ZN(n1125) );
NOR2_X1 U816 ( .A1(n1126), .A2(n1127), .ZN(G51) );
XOR2_X1 U817 ( .A(n1128), .B(n1066), .Z(n1127) );
XOR2_X1 U818 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U819 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U820 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U821 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NOR2_X1 U822 ( .A1(n1135), .A2(n1136), .ZN(n1131) );
INV_X1 U823 ( .A(KEYINPUT53), .ZN(n1136) );
XOR2_X1 U824 ( .A(n1137), .B(n1138), .Z(n1135) );
XNOR2_X1 U825 ( .A(n1139), .B(KEYINPUT17), .ZN(n1137) );
NAND3_X1 U826 ( .A1(n1140), .A2(n994), .A3(G902), .ZN(n1129) );
NAND3_X1 U827 ( .A1(n1057), .A2(n1072), .A3(n1073), .ZN(n994) );
AND4_X1 U828 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1073) );
AND4_X1 U829 ( .A1(n1090), .A2(n1145), .A3(n989), .A4(n1146), .ZN(n1072) );
NAND3_X1 U830 ( .A1(n1027), .A2(n1147), .A3(n1148), .ZN(n989) );
NAND3_X1 U831 ( .A1(n1148), .A2(n1147), .A3(n1028), .ZN(n1090) );
AND4_X1 U832 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1057) );
NOR4_X1 U833 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1152) );
NOR3_X1 U834 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1156) );
NOR3_X1 U835 ( .A1(n1160), .A2(n1161), .A3(n1012), .ZN(n1155) );
NOR2_X1 U836 ( .A1(n1162), .A2(n1163), .ZN(n1151) );
INV_X1 U837 ( .A(n1164), .ZN(n1150) );
XNOR2_X1 U838 ( .A(KEYINPUT60), .B(n1165), .ZN(n1140) );
NOR2_X1 U839 ( .A1(G952), .A2(n1166), .ZN(n1126) );
XNOR2_X1 U840 ( .A(KEYINPUT36), .B(n1062), .ZN(n1166) );
XNOR2_X1 U841 ( .A(G146), .B(n1167), .ZN(G48) );
NAND4_X1 U842 ( .A1(KEYINPUT2), .A2(n1168), .A3(n1028), .A4(n1008), .ZN(n1167) );
XNOR2_X1 U843 ( .A(n1154), .B(n1169), .ZN(G45) );
NOR2_X1 U844 ( .A1(G143), .A2(KEYINPUT18), .ZN(n1169) );
NOR4_X1 U845 ( .A1(n1160), .A2(n1158), .A3(n1170), .A4(n1171), .ZN(n1154) );
XOR2_X1 U846 ( .A(G140), .B(n1153), .Z(G42) );
AND4_X1 U847 ( .A1(n1021), .A2(n1172), .A3(n1036), .A4(n1028), .ZN(n1153) );
XNOR2_X1 U848 ( .A(G137), .B(n1149), .ZN(G39) );
NAND3_X1 U849 ( .A1(n1168), .A2(n1025), .A3(n1021), .ZN(n1149) );
INV_X1 U850 ( .A(n1157), .ZN(n1168) );
XOR2_X1 U851 ( .A(G134), .B(n1173), .Z(G36) );
NOR3_X1 U852 ( .A1(n1160), .A2(n1174), .A3(n1161), .ZN(n1173) );
XNOR2_X1 U853 ( .A(n1021), .B(KEYINPUT25), .ZN(n1174) );
XNOR2_X1 U854 ( .A(n1175), .B(n1164), .ZN(G33) );
NOR3_X1 U855 ( .A1(n1012), .A2(n1159), .A3(n1160), .ZN(n1164) );
NAND4_X1 U856 ( .A1(n1014), .A2(n1024), .A3(n1176), .A4(n1023), .ZN(n1160) );
INV_X1 U857 ( .A(n1028), .ZN(n1159) );
INV_X1 U858 ( .A(n1021), .ZN(n1012) );
NOR2_X1 U859 ( .A1(n1009), .A2(n1039), .ZN(n1021) );
INV_X1 U860 ( .A(n1177), .ZN(n1009) );
XOR2_X1 U861 ( .A(G128), .B(n1163), .Z(G30) );
NOR3_X1 U862 ( .A1(n1161), .A2(n1158), .A3(n1157), .ZN(n1163) );
NAND2_X1 U863 ( .A1(n1172), .A2(n1178), .ZN(n1157) );
AND4_X1 U864 ( .A1(n1024), .A2(n1176), .A3(n1179), .A4(n1023), .ZN(n1172) );
INV_X1 U865 ( .A(n1008), .ZN(n1158) );
INV_X1 U866 ( .A(n1027), .ZN(n1161) );
NAND3_X1 U867 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(G3) );
NAND2_X1 U868 ( .A1(G101), .A2(n1145), .ZN(n1182) );
NAND2_X1 U869 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
INV_X1 U870 ( .A(KEYINPUT22), .ZN(n1184) );
NAND2_X1 U871 ( .A1(n1185), .A2(n1186), .ZN(n1183) );
XNOR2_X1 U872 ( .A(KEYINPUT15), .B(n1187), .ZN(n1185) );
NAND2_X1 U873 ( .A1(KEYINPUT22), .A2(n1188), .ZN(n1180) );
NAND2_X1 U874 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
OR2_X1 U875 ( .A1(n1187), .A2(KEYINPUT15), .ZN(n1190) );
NAND3_X1 U876 ( .A1(n1187), .A2(n1186), .A3(KEYINPUT15), .ZN(n1189) );
INV_X1 U877 ( .A(G101), .ZN(n1186) );
INV_X1 U878 ( .A(n1145), .ZN(n1187) );
NAND3_X1 U879 ( .A1(n1014), .A2(n1148), .A3(n1025), .ZN(n1145) );
XNOR2_X1 U880 ( .A(G125), .B(n1191), .ZN(G27) );
NAND2_X1 U881 ( .A1(KEYINPUT43), .A2(n1162), .ZN(n1191) );
AND4_X1 U882 ( .A1(n1013), .A2(n1028), .A3(n1192), .A4(n1015), .ZN(n1162) );
AND2_X1 U883 ( .A1(n1176), .A2(n1008), .ZN(n1192) );
NAND2_X1 U884 ( .A1(n996), .A2(n1193), .ZN(n1176) );
NAND4_X1 U885 ( .A1(G953), .A2(G902), .A3(n1194), .A4(n1195), .ZN(n1193) );
INV_X1 U886 ( .A(G900), .ZN(n1195) );
XNOR2_X1 U887 ( .A(n1141), .B(n1196), .ZN(G24) );
NOR2_X1 U888 ( .A1(KEYINPUT26), .A2(n1197), .ZN(n1196) );
NAND4_X1 U889 ( .A1(n1198), .A2(n1147), .A3(n1033), .A4(n1199), .ZN(n1141) );
INV_X1 U890 ( .A(n1006), .ZN(n1147) );
NAND2_X1 U891 ( .A1(n1200), .A2(n1201), .ZN(n1006) );
XNOR2_X1 U892 ( .A(KEYINPUT52), .B(n1036), .ZN(n1201) );
XNOR2_X1 U893 ( .A(G119), .B(n1142), .ZN(G21) );
NAND4_X1 U894 ( .A1(n1025), .A2(n1198), .A3(n1178), .A4(n1179), .ZN(n1142) );
XNOR2_X1 U895 ( .A(G116), .B(n1143), .ZN(G18) );
NAND3_X1 U896 ( .A1(n1014), .A2(n1027), .A3(n1198), .ZN(n1143) );
NOR2_X1 U897 ( .A1(n1199), .A2(n1170), .ZN(n1027) );
INV_X1 U898 ( .A(n1033), .ZN(n1170) );
XNOR2_X1 U899 ( .A(G113), .B(n1144), .ZN(G15) );
NAND3_X1 U900 ( .A1(n1198), .A2(n1014), .A3(n1028), .ZN(n1144) );
NOR2_X1 U901 ( .A1(n1033), .A2(n1171), .ZN(n1028) );
INV_X1 U902 ( .A(n1199), .ZN(n1171) );
NOR2_X1 U903 ( .A1(n1179), .A2(n1036), .ZN(n1014) );
INV_X1 U904 ( .A(n1178), .ZN(n1036) );
AND3_X1 U905 ( .A1(n1008), .A2(n1202), .A3(n1015), .ZN(n1198) );
NOR2_X1 U906 ( .A1(n1024), .A2(n1019), .ZN(n1015) );
INV_X1 U907 ( .A(n1023), .ZN(n1019) );
XNOR2_X1 U908 ( .A(G110), .B(n1146), .ZN(G12) );
NAND3_X1 U909 ( .A1(n1025), .A2(n1148), .A3(n1013), .ZN(n1146) );
NOR2_X1 U910 ( .A1(n1178), .A2(n1200), .ZN(n1013) );
INV_X1 U911 ( .A(n1179), .ZN(n1200) );
NAND3_X1 U912 ( .A1(n1203), .A2(n1204), .A3(n1040), .ZN(n1179) );
NAND3_X1 U913 ( .A1(n1205), .A2(n1206), .A3(n1077), .ZN(n1040) );
NAND2_X1 U914 ( .A1(KEYINPUT28), .A2(n1206), .ZN(n1204) );
OR2_X1 U915 ( .A1(n1030), .A2(KEYINPUT28), .ZN(n1203) );
NAND2_X1 U916 ( .A1(n1078), .A2(n1207), .ZN(n1030) );
NAND2_X1 U917 ( .A1(n1077), .A2(n1205), .ZN(n1207) );
AND2_X1 U918 ( .A1(n1208), .A2(n1209), .ZN(n1077) );
NAND2_X1 U919 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND2_X1 U920 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
OR2_X1 U921 ( .A1(n1214), .A2(KEYINPUT33), .ZN(n1212) );
XNOR2_X1 U922 ( .A(n1215), .B(n1216), .ZN(n1210) );
NAND2_X1 U923 ( .A1(n1214), .A2(n1217), .ZN(n1208) );
NAND2_X1 U924 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
INV_X1 U925 ( .A(KEYINPUT33), .ZN(n1219) );
NAND2_X1 U926 ( .A1(n1220), .A2(n1213), .ZN(n1218) );
INV_X1 U927 ( .A(KEYINPUT45), .ZN(n1213) );
XNOR2_X1 U928 ( .A(n1215), .B(n1221), .ZN(n1220) );
NAND2_X1 U929 ( .A1(n1222), .A2(n1223), .ZN(n1215) );
NAND2_X1 U930 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
XOR2_X1 U931 ( .A(KEYINPUT9), .B(n1226), .Z(n1222) );
NOR2_X1 U932 ( .A1(n1225), .A2(n1224), .ZN(n1226) );
XOR2_X1 U933 ( .A(KEYINPUT23), .B(G110), .Z(n1224) );
XOR2_X1 U934 ( .A(G119), .B(G128), .Z(n1225) );
XOR2_X1 U935 ( .A(n1227), .B(G137), .Z(n1214) );
NAND2_X1 U936 ( .A1(n1228), .A2(G221), .ZN(n1227) );
INV_X1 U937 ( .A(n1206), .ZN(n1078) );
NAND2_X1 U938 ( .A1(G217), .A2(n1229), .ZN(n1206) );
XNOR2_X1 U939 ( .A(n1230), .B(G472), .ZN(n1178) );
NAND2_X1 U940 ( .A1(n1231), .A2(n1205), .ZN(n1230) );
XOR2_X1 U941 ( .A(n1232), .B(n1233), .Z(n1231) );
XNOR2_X1 U942 ( .A(n1234), .B(n1102), .ZN(n1233) );
INV_X1 U943 ( .A(n1235), .ZN(n1234) );
XOR2_X1 U944 ( .A(n1236), .B(n1237), .Z(n1232) );
XOR2_X1 U945 ( .A(KEYINPUT29), .B(n1099), .Z(n1237) );
NOR3_X1 U946 ( .A1(G237), .A2(G953), .A3(n1165), .ZN(n1099) );
INV_X1 U947 ( .A(G210), .ZN(n1165) );
NOR2_X1 U948 ( .A1(KEYINPUT40), .A2(n1139), .ZN(n1236) );
AND4_X1 U949 ( .A1(n1008), .A2(n1024), .A3(n1202), .A4(n1023), .ZN(n1148) );
NAND2_X1 U950 ( .A1(G221), .A2(n1229), .ZN(n1023) );
NAND2_X1 U951 ( .A1(G234), .A2(n1238), .ZN(n1229) );
NAND2_X1 U952 ( .A1(n1239), .A2(n1240), .ZN(n1202) );
NAND4_X1 U953 ( .A1(G902), .A2(n1241), .A3(n1194), .A4(n1069), .ZN(n1240) );
INV_X1 U954 ( .A(G898), .ZN(n1069) );
XNOR2_X1 U955 ( .A(KEYINPUT0), .B(n1062), .ZN(n1241) );
XOR2_X1 U956 ( .A(n996), .B(KEYINPUT39), .Z(n1239) );
NAND3_X1 U957 ( .A1(n1194), .A2(n1062), .A3(G952), .ZN(n996) );
NAND2_X1 U958 ( .A1(G237), .A2(G234), .ZN(n1194) );
XNOR2_X1 U959 ( .A(n1242), .B(G469), .ZN(n1024) );
NAND3_X1 U960 ( .A1(n1243), .A2(n1244), .A3(n1205), .ZN(n1242) );
NAND2_X1 U961 ( .A1(KEYINPUT63), .A2(n1245), .ZN(n1244) );
XNOR2_X1 U962 ( .A(n1113), .B(n1246), .ZN(n1245) );
NOR2_X1 U963 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
INV_X1 U964 ( .A(KEYINPUT48), .ZN(n1247) );
OR3_X1 U965 ( .A1(n1249), .A2(n1248), .A3(KEYINPUT63), .ZN(n1243) );
XOR2_X1 U966 ( .A(n1250), .B(n1251), .Z(n1248) );
INV_X1 U967 ( .A(n1102), .ZN(n1251) );
XOR2_X1 U968 ( .A(G131), .B(n1055), .Z(n1102) );
XOR2_X1 U969 ( .A(G134), .B(G137), .Z(n1055) );
NAND2_X1 U970 ( .A1(n1252), .A2(n1253), .ZN(n1250) );
NAND2_X1 U971 ( .A1(n1051), .A2(n1254), .ZN(n1253) );
NAND2_X1 U972 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
NAND2_X1 U973 ( .A1(KEYINPUT14), .A2(n1117), .ZN(n1256) );
INV_X1 U974 ( .A(n1118), .ZN(n1051) );
NAND2_X1 U975 ( .A1(n1120), .A2(n1257), .ZN(n1252) );
NAND2_X1 U976 ( .A1(KEYINPUT14), .A2(n1258), .ZN(n1257) );
NAND2_X1 U977 ( .A1(n1118), .A2(n1255), .ZN(n1258) );
INV_X1 U978 ( .A(KEYINPUT13), .ZN(n1255) );
XOR2_X1 U979 ( .A(G128), .B(n1259), .Z(n1118) );
NOR2_X1 U980 ( .A1(KEYINPUT10), .A2(n1260), .ZN(n1259) );
INV_X1 U981 ( .A(n1117), .ZN(n1120) );
XNOR2_X1 U982 ( .A(n1261), .B(n1262), .ZN(n1117) );
NOR2_X1 U983 ( .A1(G101), .A2(KEYINPUT62), .ZN(n1262) );
NAND2_X1 U984 ( .A1(n1263), .A2(n1264), .ZN(n1261) );
NAND2_X1 U985 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NAND2_X1 U986 ( .A1(KEYINPUT44), .A2(n1267), .ZN(n1265) );
NAND2_X1 U987 ( .A1(KEYINPUT1), .A2(n1268), .ZN(n1267) );
INV_X1 U988 ( .A(G107), .ZN(n1268) );
NAND2_X1 U989 ( .A1(G107), .A2(n1269), .ZN(n1263) );
NAND2_X1 U990 ( .A1(KEYINPUT1), .A2(n1270), .ZN(n1269) );
NAND2_X1 U991 ( .A1(KEYINPUT44), .A2(G104), .ZN(n1270) );
XNOR2_X1 U992 ( .A(KEYINPUT48), .B(n1113), .ZN(n1249) );
XOR2_X1 U993 ( .A(n1271), .B(n1114), .Z(n1113) );
XNOR2_X1 U994 ( .A(G140), .B(G110), .ZN(n1114) );
NAND2_X1 U995 ( .A1(G227), .A2(n1062), .ZN(n1271) );
NOR2_X1 U996 ( .A1(n1039), .A2(n1177), .ZN(n1008) );
NOR2_X1 U997 ( .A1(n1272), .A2(n1038), .ZN(n1177) );
NOR2_X1 U998 ( .A1(n1042), .A2(n1273), .ZN(n1038) );
AND2_X1 U999 ( .A1(n1274), .A2(n1042), .ZN(n1272) );
NAND2_X1 U1000 ( .A1(n1275), .A2(n1205), .ZN(n1042) );
XOR2_X1 U1001 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U1002 ( .A(n1066), .B(n1138), .ZN(n1277) );
XNOR2_X1 U1003 ( .A(n1278), .B(n1279), .ZN(n1066) );
XNOR2_X1 U1004 ( .A(n1266), .B(n1280), .ZN(n1279) );
XNOR2_X1 U1005 ( .A(n1197), .B(G107), .ZN(n1280) );
XNOR2_X1 U1006 ( .A(n1235), .B(n1281), .ZN(n1278) );
NOR2_X1 U1007 ( .A1(G110), .A2(KEYINPUT7), .ZN(n1281) );
XOR2_X1 U1008 ( .A(G101), .B(n1095), .Z(n1235) );
XNOR2_X1 U1009 ( .A(n1282), .B(n1283), .ZN(n1095) );
XNOR2_X1 U1010 ( .A(G113), .B(G119), .ZN(n1282) );
XOR2_X1 U1011 ( .A(n1133), .B(n1284), .Z(n1276) );
NOR2_X1 U1012 ( .A1(KEYINPUT34), .A2(n1101), .ZN(n1284) );
INV_X1 U1013 ( .A(n1139), .ZN(n1101) );
XOR2_X1 U1014 ( .A(G128), .B(n1260), .Z(n1139) );
XOR2_X1 U1015 ( .A(G146), .B(G143), .Z(n1260) );
NAND2_X1 U1016 ( .A1(G224), .A2(n1062), .ZN(n1133) );
XNOR2_X1 U1017 ( .A(n1273), .B(KEYINPUT50), .ZN(n1274) );
INV_X1 U1018 ( .A(n1043), .ZN(n1273) );
NAND2_X1 U1019 ( .A1(n1285), .A2(n1286), .ZN(n1043) );
XNOR2_X1 U1020 ( .A(G210), .B(KEYINPUT16), .ZN(n1285) );
INV_X1 U1021 ( .A(n1010), .ZN(n1039) );
NAND2_X1 U1022 ( .A1(G214), .A2(n1286), .ZN(n1010) );
NAND2_X1 U1023 ( .A1(n1287), .A2(n1238), .ZN(n1286) );
NOR2_X1 U1024 ( .A1(n1033), .A2(n1199), .ZN(n1025) );
XOR2_X1 U1025 ( .A(n1034), .B(KEYINPUT58), .Z(n1199) );
XNOR2_X1 U1026 ( .A(n1288), .B(G475), .ZN(n1034) );
NAND2_X1 U1027 ( .A1(n1087), .A2(n1205), .ZN(n1288) );
XNOR2_X1 U1028 ( .A(n1289), .B(n1290), .ZN(n1087) );
XNOR2_X1 U1029 ( .A(n1266), .B(n1291), .ZN(n1290) );
XNOR2_X1 U1030 ( .A(KEYINPUT24), .B(n1175), .ZN(n1291) );
INV_X1 U1031 ( .A(G131), .ZN(n1175) );
INV_X1 U1032 ( .A(G104), .ZN(n1266) );
XOR2_X1 U1033 ( .A(n1292), .B(n1293), .Z(n1289) );
NOR2_X1 U1034 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
AND4_X1 U1035 ( .A1(n1296), .A2(G214), .A3(n1062), .A4(n1287), .ZN(n1295) );
NOR2_X1 U1036 ( .A1(n1297), .A2(n1296), .ZN(n1294) );
XOR2_X1 U1037 ( .A(G143), .B(KEYINPUT59), .Z(n1296) );
AND3_X1 U1038 ( .A1(G214), .A2(n1062), .A3(n1287), .ZN(n1297) );
INV_X1 U1039 ( .A(G237), .ZN(n1287) );
XNOR2_X1 U1040 ( .A(n1298), .B(n1216), .ZN(n1292) );
INV_X1 U1041 ( .A(n1221), .ZN(n1216) );
XNOR2_X1 U1042 ( .A(n1050), .B(G146), .ZN(n1221) );
XNOR2_X1 U1043 ( .A(G140), .B(n1138), .ZN(n1050) );
XOR2_X1 U1044 ( .A(G125), .B(KEYINPUT42), .Z(n1138) );
NAND2_X1 U1045 ( .A1(KEYINPUT35), .A2(n1299), .ZN(n1298) );
XNOR2_X1 U1046 ( .A(n1197), .B(G113), .ZN(n1299) );
XNOR2_X1 U1047 ( .A(n1300), .B(G478), .ZN(n1033) );
NAND2_X1 U1048 ( .A1(n1082), .A2(n1205), .ZN(n1300) );
XNOR2_X1 U1049 ( .A(n1238), .B(KEYINPUT51), .ZN(n1205) );
INV_X1 U1050 ( .A(G902), .ZN(n1238) );
XNOR2_X1 U1051 ( .A(n1301), .B(n1302), .ZN(n1082) );
XOR2_X1 U1052 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U1053 ( .A(n1197), .B(n1305), .ZN(n1304) );
NOR2_X1 U1054 ( .A1(KEYINPUT32), .A2(n1306), .ZN(n1305) );
XOR2_X1 U1055 ( .A(G134), .B(n1307), .Z(n1306) );
NOR2_X1 U1056 ( .A1(KEYINPUT55), .A2(n1308), .ZN(n1307) );
XNOR2_X1 U1057 ( .A(G128), .B(G143), .ZN(n1308) );
INV_X1 U1058 ( .A(G122), .ZN(n1197) );
AND2_X1 U1059 ( .A1(n1228), .A2(G217), .ZN(n1303) );
AND2_X1 U1060 ( .A1(G234), .A2(n1062), .ZN(n1228) );
INV_X1 U1061 ( .A(G953), .ZN(n1062) );
XNOR2_X1 U1062 ( .A(n1283), .B(n1309), .ZN(n1301) );
NOR2_X1 U1063 ( .A1(G107), .A2(KEYINPUT21), .ZN(n1309) );
XOR2_X1 U1064 ( .A(G116), .B(KEYINPUT54), .Z(n1283) );
endmodule


