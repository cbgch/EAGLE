//Key = 0010110111001101110101100101100000011110010010000000010000011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343;

XOR2_X1 U738 ( .A(G107), .B(n1023), .Z(G9) );
NOR2_X1 U739 ( .A1(n1024), .A2(n1025), .ZN(G75) );
NOR3_X1 U740 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NAND3_X1 U741 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1026) );
NAND2_X1 U742 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U743 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND3_X1 U744 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NAND2_X1 U745 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NAND3_X1 U746 ( .A1(n1041), .A2(n1042), .A3(KEYINPUT43), .ZN(n1039) );
NAND4_X1 U747 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1036) );
NAND2_X1 U748 ( .A1(n1041), .A2(n1047), .ZN(n1045) );
NAND2_X1 U749 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U750 ( .A1(n1042), .A2(n1050), .ZN(n1048) );
INV_X1 U751 ( .A(KEYINPUT43), .ZN(n1050) );
INV_X1 U752 ( .A(n1051), .ZN(n1044) );
NAND3_X1 U753 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1043) );
NAND3_X1 U754 ( .A1(n1041), .A2(n1055), .A3(n1053), .ZN(n1034) );
NAND2_X1 U755 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U756 ( .A1(n1038), .A2(n1058), .ZN(n1057) );
OR2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U758 ( .A1(n1046), .A2(n1061), .ZN(n1056) );
NAND2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
INV_X1 U761 ( .A(n1066), .ZN(n1032) );
NOR3_X1 U762 ( .A1(n1067), .A2(G953), .A3(G952), .ZN(n1024) );
INV_X1 U763 ( .A(n1029), .ZN(n1067) );
NAND4_X1 U764 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1029) );
NOR4_X1 U765 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1071) );
XNOR2_X1 U766 ( .A(G469), .B(n1076), .ZN(n1075) );
NAND2_X1 U767 ( .A1(KEYINPUT27), .A2(n1077), .ZN(n1076) );
XNOR2_X1 U768 ( .A(KEYINPUT46), .B(n1078), .ZN(n1077) );
XOR2_X1 U769 ( .A(n1079), .B(n1080), .Z(n1072) );
XOR2_X1 U770 ( .A(KEYINPUT14), .B(n1081), .Z(n1080) );
NOR2_X1 U771 ( .A1(KEYINPUT54), .A2(n1082), .ZN(n1081) );
NOR3_X1 U772 ( .A1(n1054), .A2(n1083), .A3(n1064), .ZN(n1070) );
NAND2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1069) );
XNOR2_X1 U774 ( .A(KEYINPUT58), .B(n1086), .ZN(n1084) );
XOR2_X1 U775 ( .A(n1087), .B(n1088), .Z(n1068) );
NAND2_X1 U776 ( .A1(KEYINPUT35), .A2(n1089), .ZN(n1088) );
NAND2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(G72) );
NAND2_X1 U778 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U779 ( .A(KEYINPUT5), .B(n1094), .Z(n1090) );
NOR2_X1 U780 ( .A1(n1095), .A2(n1092), .ZN(n1094) );
NAND2_X1 U781 ( .A1(G953), .A2(n1096), .ZN(n1092) );
NAND2_X1 U782 ( .A1(G227), .A2(n1097), .ZN(n1096) );
XNOR2_X1 U783 ( .A(KEYINPUT39), .B(n1098), .ZN(n1097) );
XOR2_X1 U784 ( .A(n1093), .B(KEYINPUT29), .Z(n1095) );
NAND2_X1 U785 ( .A1(n1099), .A2(n1100), .ZN(n1093) );
NAND2_X1 U786 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U787 ( .A(KEYINPUT38), .B(n1103), .Z(n1099) );
NOR2_X1 U788 ( .A1(n1101), .A2(n1102), .ZN(n1103) );
NAND2_X1 U789 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NAND2_X1 U790 ( .A1(G953), .A2(n1098), .ZN(n1105) );
XNOR2_X1 U791 ( .A(n1106), .B(n1107), .ZN(n1104) );
XOR2_X1 U792 ( .A(n1108), .B(n1109), .Z(n1107) );
AND2_X1 U793 ( .A1(n1110), .A2(n1028), .ZN(n1101) );
XNOR2_X1 U794 ( .A(KEYINPUT59), .B(n1030), .ZN(n1110) );
XOR2_X1 U795 ( .A(n1111), .B(n1112), .Z(G69) );
NOR3_X1 U796 ( .A1(n1113), .A2(KEYINPUT42), .A3(n1114), .ZN(n1112) );
NOR3_X1 U797 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
AND2_X1 U798 ( .A1(n1030), .A2(n1027), .ZN(n1117) );
NOR2_X1 U799 ( .A1(G898), .A2(n1030), .ZN(n1116) );
XOR2_X1 U800 ( .A(KEYINPUT30), .B(n1118), .Z(n1113) );
AND3_X1 U801 ( .A1(n1115), .A2(n1030), .A3(n1027), .ZN(n1118) );
NAND2_X1 U802 ( .A1(G953), .A2(n1119), .ZN(n1111) );
NAND2_X1 U803 ( .A1(G898), .A2(G224), .ZN(n1119) );
NOR2_X1 U804 ( .A1(n1120), .A2(n1121), .ZN(G66) );
XOR2_X1 U805 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U806 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
NOR2_X1 U807 ( .A1(n1120), .A2(n1126), .ZN(G63) );
NOR2_X1 U808 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U809 ( .A(KEYINPUT45), .B(n1129), .Z(n1128) );
AND2_X1 U810 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U811 ( .A1(n1131), .A2(n1130), .ZN(n1127) );
XOR2_X1 U812 ( .A(n1132), .B(KEYINPUT2), .Z(n1130) );
NOR2_X1 U813 ( .A1(n1125), .A2(n1086), .ZN(n1131) );
NOR2_X1 U814 ( .A1(n1120), .A2(n1133), .ZN(G60) );
XOR2_X1 U815 ( .A(n1134), .B(n1135), .Z(n1133) );
AND2_X1 U816 ( .A1(G475), .A2(n1136), .ZN(n1134) );
XOR2_X1 U817 ( .A(G104), .B(n1137), .Z(G6) );
NOR3_X1 U818 ( .A1(n1049), .A2(n1138), .A3(n1040), .ZN(n1137) );
NOR3_X1 U819 ( .A1(n1120), .A2(n1139), .A3(n1140), .ZN(G57) );
NOR2_X1 U820 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
INV_X1 U821 ( .A(n1143), .ZN(n1142) );
NOR2_X1 U822 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
AND2_X1 U823 ( .A1(KEYINPUT56), .A2(n1146), .ZN(n1145) );
NOR3_X1 U824 ( .A1(KEYINPUT56), .A2(n1146), .A3(n1147), .ZN(n1144) );
NOR2_X1 U825 ( .A1(n1148), .A2(n1143), .ZN(n1139) );
XOR2_X1 U826 ( .A(n1149), .B(n1150), .Z(n1143) );
NOR2_X1 U827 ( .A1(n1089), .A2(n1125), .ZN(n1150) );
NOR2_X1 U828 ( .A1(n1146), .A2(n1147), .ZN(n1148) );
INV_X1 U829 ( .A(KEYINPUT7), .ZN(n1147) );
XOR2_X1 U830 ( .A(n1151), .B(n1152), .Z(n1146) );
NOR2_X1 U831 ( .A1(n1120), .A2(n1153), .ZN(G54) );
XOR2_X1 U832 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U833 ( .A(n1108), .B(n1156), .Z(n1155) );
XOR2_X1 U834 ( .A(n1157), .B(n1158), .Z(n1154) );
XNOR2_X1 U835 ( .A(G140), .B(n1159), .ZN(n1157) );
NOR2_X1 U836 ( .A1(n1160), .A2(n1125), .ZN(n1159) );
NOR2_X1 U837 ( .A1(n1120), .A2(n1161), .ZN(G51) );
XOR2_X1 U838 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U839 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND3_X1 U840 ( .A1(n1136), .A2(n1082), .A3(KEYINPUT22), .ZN(n1164) );
INV_X1 U841 ( .A(n1125), .ZN(n1136) );
NAND2_X1 U842 ( .A1(G902), .A2(n1166), .ZN(n1125) );
OR2_X1 U843 ( .A1(n1028), .A2(n1027), .ZN(n1166) );
NAND4_X1 U844 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1027) );
NOR4_X1 U845 ( .A1(n1171), .A2(n1172), .A3(n1023), .A4(n1173), .ZN(n1170) );
INV_X1 U846 ( .A(n1174), .ZN(n1173) );
AND3_X1 U847 ( .A1(n1046), .A2(n1175), .A3(n1042), .ZN(n1023) );
NAND2_X1 U848 ( .A1(n1176), .A2(n1177), .ZN(n1169) );
NAND2_X1 U849 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XOR2_X1 U850 ( .A(n1180), .B(KEYINPUT61), .Z(n1178) );
NAND3_X1 U851 ( .A1(n1059), .A2(n1181), .A3(n1051), .ZN(n1180) );
NAND3_X1 U852 ( .A1(n1182), .A2(n1175), .A3(n1183), .ZN(n1168) );
XNOR2_X1 U853 ( .A(n1046), .B(KEYINPUT25), .ZN(n1183) );
INV_X1 U854 ( .A(n1138), .ZN(n1175) );
NAND3_X1 U855 ( .A1(n1053), .A2(n1184), .A3(n1185), .ZN(n1167) );
NAND4_X1 U856 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1028) );
NOR4_X1 U857 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
INV_X1 U858 ( .A(n1194), .ZN(n1190) );
NAND3_X1 U859 ( .A1(n1195), .A2(n1196), .A3(n1184), .ZN(n1188) );
NAND2_X1 U860 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NAND2_X1 U861 ( .A1(n1199), .A2(n1182), .ZN(n1198) );
XNOR2_X1 U862 ( .A(n1200), .B(KEYINPUT28), .ZN(n1199) );
NAND2_X1 U863 ( .A1(n1053), .A2(n1038), .ZN(n1197) );
INV_X1 U864 ( .A(n1201), .ZN(n1053) );
XNOR2_X1 U865 ( .A(n1202), .B(n1203), .ZN(n1162) );
NAND2_X1 U866 ( .A1(KEYINPUT53), .A2(n1204), .ZN(n1203) );
NOR2_X1 U867 ( .A1(n1030), .A2(G952), .ZN(n1120) );
XNOR2_X1 U868 ( .A(G146), .B(n1205), .ZN(G48) );
NAND4_X1 U869 ( .A1(n1182), .A2(n1184), .A3(n1195), .A4(n1200), .ZN(n1205) );
XNOR2_X1 U870 ( .A(G143), .B(n1186), .ZN(G45) );
NAND3_X1 U871 ( .A1(n1059), .A2(n1195), .A3(n1206), .ZN(n1186) );
NOR3_X1 U872 ( .A1(n1062), .A2(n1207), .A3(n1208), .ZN(n1206) );
XNOR2_X1 U873 ( .A(G140), .B(n1209), .ZN(G42) );
NAND2_X1 U874 ( .A1(KEYINPUT19), .A2(n1192), .ZN(n1209) );
AND4_X1 U875 ( .A1(n1182), .A2(n1060), .A3(n1038), .A4(n1195), .ZN(n1192) );
XOR2_X1 U876 ( .A(n1210), .B(n1211), .Z(G39) );
XNOR2_X1 U877 ( .A(G137), .B(KEYINPUT55), .ZN(n1211) );
NAND4_X1 U878 ( .A1(n1212), .A2(n1051), .A3(n1038), .A4(n1184), .ZN(n1210) );
XNOR2_X1 U879 ( .A(n1213), .B(KEYINPUT18), .ZN(n1212) );
XOR2_X1 U880 ( .A(n1191), .B(n1214), .Z(G36) );
NOR2_X1 U881 ( .A1(KEYINPUT1), .A2(n1215), .ZN(n1214) );
XNOR2_X1 U882 ( .A(G134), .B(KEYINPUT50), .ZN(n1215) );
AND4_X1 U883 ( .A1(n1059), .A2(n1038), .A3(n1195), .A4(n1042), .ZN(n1191) );
XNOR2_X1 U884 ( .A(G131), .B(n1187), .ZN(G33) );
NAND4_X1 U885 ( .A1(n1182), .A2(n1059), .A3(n1038), .A4(n1195), .ZN(n1187) );
NOR2_X1 U886 ( .A1(n1216), .A2(n1064), .ZN(n1038) );
XNOR2_X1 U887 ( .A(G128), .B(n1194), .ZN(G30) );
NAND4_X1 U888 ( .A1(n1184), .A2(n1195), .A3(n1042), .A4(n1200), .ZN(n1194) );
NOR3_X1 U889 ( .A1(n1213), .A2(n1054), .A3(n1217), .ZN(n1195) );
XNOR2_X1 U890 ( .A(n1152), .B(n1218), .ZN(G3) );
NOR3_X1 U891 ( .A1(n1219), .A2(n1138), .A3(n1201), .ZN(n1218) );
NAND4_X1 U892 ( .A1(n1176), .A2(n1220), .A3(n1181), .A4(n1221), .ZN(n1138) );
XOR2_X1 U893 ( .A(KEYINPUT21), .B(n1059), .Z(n1219) );
NAND2_X1 U894 ( .A1(n1222), .A2(n1223), .ZN(G27) );
NAND2_X1 U895 ( .A1(n1224), .A2(n1204), .ZN(n1223) );
NAND2_X1 U896 ( .A1(G125), .A2(n1225), .ZN(n1222) );
NAND2_X1 U897 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
NAND2_X1 U898 ( .A1(KEYINPUT49), .A2(n1193), .ZN(n1227) );
INV_X1 U899 ( .A(n1228), .ZN(n1193) );
OR2_X1 U900 ( .A1(n1224), .A2(KEYINPUT49), .ZN(n1226) );
NOR2_X1 U901 ( .A1(KEYINPUT48), .A2(n1228), .ZN(n1224) );
NAND3_X1 U902 ( .A1(n1041), .A2(n1182), .A3(n1229), .ZN(n1228) );
NOR3_X1 U903 ( .A1(n1230), .A2(n1213), .A3(n1062), .ZN(n1229) );
INV_X1 U904 ( .A(n1200), .ZN(n1062) );
AND2_X1 U905 ( .A1(n1066), .A2(n1231), .ZN(n1213) );
NAND2_X1 U906 ( .A1(n1232), .A2(n1098), .ZN(n1231) );
INV_X1 U907 ( .A(G900), .ZN(n1098) );
XOR2_X1 U908 ( .A(n1233), .B(n1172), .Z(G24) );
NOR4_X1 U909 ( .A1(n1234), .A2(n1040), .A3(n1208), .A4(n1207), .ZN(n1172) );
INV_X1 U910 ( .A(n1046), .ZN(n1040) );
NOR2_X1 U911 ( .A1(n1074), .A2(n1235), .ZN(n1046) );
NAND2_X1 U912 ( .A1(KEYINPUT41), .A2(n1236), .ZN(n1233) );
XOR2_X1 U913 ( .A(G119), .B(n1237), .Z(G21) );
NOR3_X1 U914 ( .A1(n1234), .A2(n1238), .A3(n1201), .ZN(n1237) );
XNOR2_X1 U915 ( .A(n1184), .B(KEYINPUT62), .ZN(n1238) );
AND2_X1 U916 ( .A1(n1235), .A2(n1074), .ZN(n1184) );
XNOR2_X1 U917 ( .A(G116), .B(n1239), .ZN(G18) );
NAND2_X1 U918 ( .A1(KEYINPUT60), .A2(n1171), .ZN(n1239) );
AND3_X1 U919 ( .A1(n1059), .A2(n1042), .A3(n1185), .ZN(n1171) );
INV_X1 U920 ( .A(n1234), .ZN(n1185) );
NAND3_X1 U921 ( .A1(n1200), .A2(n1181), .A3(n1041), .ZN(n1234) );
XOR2_X1 U922 ( .A(n1176), .B(KEYINPUT51), .Z(n1200) );
NOR2_X1 U923 ( .A1(n1073), .A2(n1207), .ZN(n1042) );
XNOR2_X1 U924 ( .A(G113), .B(n1174), .ZN(G15) );
NAND3_X1 U925 ( .A1(n1041), .A2(n1182), .A3(n1240), .ZN(n1174) );
AND3_X1 U926 ( .A1(n1059), .A2(n1181), .A3(n1176), .ZN(n1240) );
NOR2_X1 U927 ( .A1(n1074), .A2(n1241), .ZN(n1059) );
INV_X1 U928 ( .A(n1049), .ZN(n1182) );
NAND2_X1 U929 ( .A1(n1207), .A2(n1073), .ZN(n1049) );
AND2_X1 U930 ( .A1(n1052), .A2(n1221), .ZN(n1041) );
XNOR2_X1 U931 ( .A(n1220), .B(KEYINPUT20), .ZN(n1052) );
XNOR2_X1 U932 ( .A(G110), .B(n1242), .ZN(G12) );
NAND3_X1 U933 ( .A1(KEYINPUT15), .A2(n1176), .A3(n1243), .ZN(n1242) );
XOR2_X1 U934 ( .A(n1179), .B(KEYINPUT8), .Z(n1243) );
NAND3_X1 U935 ( .A1(n1060), .A2(n1181), .A3(n1051), .ZN(n1179) );
NOR3_X1 U936 ( .A1(n1217), .A2(n1054), .A3(n1201), .ZN(n1051) );
NAND2_X1 U937 ( .A1(n1207), .A2(n1208), .ZN(n1201) );
INV_X1 U938 ( .A(n1073), .ZN(n1208) );
XNOR2_X1 U939 ( .A(n1244), .B(G475), .ZN(n1073) );
OR2_X1 U940 ( .A1(n1135), .A2(G902), .ZN(n1244) );
XNOR2_X1 U941 ( .A(n1245), .B(n1246), .ZN(n1135) );
XNOR2_X1 U942 ( .A(n1247), .B(n1248), .ZN(n1246) );
XNOR2_X1 U943 ( .A(n1249), .B(n1250), .ZN(n1245) );
NAND2_X1 U944 ( .A1(n1251), .A2(n1252), .ZN(n1249) );
NAND2_X1 U945 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
XOR2_X1 U946 ( .A(n1255), .B(KEYINPUT6), .Z(n1251) );
OR2_X1 U947 ( .A1(n1254), .A2(n1253), .ZN(n1255) );
XOR2_X1 U948 ( .A(n1256), .B(n1257), .Z(n1253) );
NAND2_X1 U949 ( .A1(G214), .A2(n1258), .ZN(n1256) );
INV_X1 U950 ( .A(G131), .ZN(n1254) );
NOR2_X1 U951 ( .A1(n1259), .A2(n1083), .ZN(n1207) );
NOR2_X1 U952 ( .A1(n1085), .A2(G478), .ZN(n1083) );
XNOR2_X1 U953 ( .A(KEYINPUT37), .B(n1260), .ZN(n1259) );
NOR2_X1 U954 ( .A1(n1086), .A2(n1261), .ZN(n1260) );
XNOR2_X1 U955 ( .A(KEYINPUT34), .B(n1085), .ZN(n1261) );
NAND2_X1 U956 ( .A1(n1132), .A2(n1262), .ZN(n1085) );
XNOR2_X1 U957 ( .A(n1263), .B(n1264), .ZN(n1132) );
NOR2_X1 U958 ( .A1(n1265), .A2(KEYINPUT10), .ZN(n1264) );
AND2_X1 U959 ( .A1(n1266), .A2(G217), .ZN(n1265) );
XOR2_X1 U960 ( .A(n1267), .B(n1268), .Z(n1263) );
NOR2_X1 U961 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
XOR2_X1 U962 ( .A(KEYINPUT11), .B(n1271), .Z(n1270) );
NOR2_X1 U963 ( .A1(G134), .A2(n1272), .ZN(n1271) );
AND2_X1 U964 ( .A1(n1272), .A2(G134), .ZN(n1269) );
NAND2_X1 U965 ( .A1(n1273), .A2(KEYINPUT4), .ZN(n1267) );
XOR2_X1 U966 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U967 ( .A(n1276), .B(G107), .ZN(n1275) );
XNOR2_X1 U968 ( .A(G122), .B(KEYINPUT32), .ZN(n1274) );
INV_X1 U969 ( .A(G478), .ZN(n1086) );
INV_X1 U970 ( .A(n1221), .ZN(n1054) );
NAND2_X1 U971 ( .A1(G221), .A2(n1277), .ZN(n1221) );
NAND2_X1 U972 ( .A1(G234), .A2(n1262), .ZN(n1277) );
INV_X1 U973 ( .A(n1220), .ZN(n1217) );
XOR2_X1 U974 ( .A(n1078), .B(n1160), .Z(n1220) );
INV_X1 U975 ( .A(G469), .ZN(n1160) );
NAND2_X1 U976 ( .A1(n1278), .A2(n1262), .ZN(n1078) );
XOR2_X1 U977 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U978 ( .A(n1281), .B(n1282), .Z(n1280) );
XNOR2_X1 U979 ( .A(G101), .B(KEYINPUT24), .ZN(n1282) );
NAND2_X1 U980 ( .A1(n1283), .A2(KEYINPUT17), .ZN(n1281) );
XNOR2_X1 U981 ( .A(G110), .B(G140), .ZN(n1283) );
XOR2_X1 U982 ( .A(n1284), .B(n1158), .Z(n1279) );
XNOR2_X1 U983 ( .A(n1285), .B(n1286), .ZN(n1158) );
XOR2_X1 U984 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U985 ( .A(KEYINPUT23), .B(G104), .Z(n1288) );
NOR2_X1 U986 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
INV_X1 U987 ( .A(G227), .ZN(n1290) );
XOR2_X1 U988 ( .A(n1291), .B(n1292), .Z(n1285) );
NOR2_X1 U989 ( .A1(G107), .A2(KEYINPUT31), .ZN(n1292) );
NAND2_X1 U990 ( .A1(KEYINPUT63), .A2(n1108), .ZN(n1284) );
XOR2_X1 U991 ( .A(n1293), .B(n1294), .Z(n1108) );
NOR2_X1 U992 ( .A1(KEYINPUT33), .A2(n1257), .ZN(n1294) );
XNOR2_X1 U993 ( .A(n1295), .B(n1250), .ZN(n1293) );
NAND2_X1 U994 ( .A1(KEYINPUT44), .A2(n1296), .ZN(n1295) );
NAND2_X1 U995 ( .A1(n1066), .A2(n1297), .ZN(n1181) );
NAND2_X1 U996 ( .A1(n1232), .A2(n1298), .ZN(n1297) );
XOR2_X1 U997 ( .A(KEYINPUT16), .B(G898), .Z(n1298) );
AND3_X1 U998 ( .A1(n1299), .A2(n1300), .A3(G953), .ZN(n1232) );
XNOR2_X1 U999 ( .A(KEYINPUT3), .B(n1262), .ZN(n1299) );
NAND3_X1 U1000 ( .A1(n1300), .A2(n1030), .A3(G952), .ZN(n1066) );
INV_X1 U1001 ( .A(G953), .ZN(n1030) );
NAND2_X1 U1002 ( .A1(G237), .A2(G234), .ZN(n1300) );
INV_X1 U1003 ( .A(n1230), .ZN(n1060) );
NAND2_X1 U1004 ( .A1(n1241), .A2(n1074), .ZN(n1230) );
NAND3_X1 U1005 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1074) );
NAND2_X1 U1006 ( .A1(n1304), .A2(n1123), .ZN(n1303) );
OR3_X1 U1007 ( .A1(n1123), .A2(n1304), .A3(G902), .ZN(n1302) );
NOR2_X1 U1008 ( .A1(n1124), .A2(G234), .ZN(n1304) );
INV_X1 U1009 ( .A(G217), .ZN(n1124) );
XNOR2_X1 U1010 ( .A(n1305), .B(n1306), .ZN(n1123) );
XOR2_X1 U1011 ( .A(n1307), .B(n1308), .Z(n1306) );
XOR2_X1 U1012 ( .A(n1309), .B(n1310), .Z(n1308) );
NOR2_X1 U1013 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U1014 ( .A(KEYINPUT26), .B(n1313), .Z(n1312) );
NOR2_X1 U1015 ( .A1(G146), .A2(n1106), .ZN(n1313) );
NOR2_X1 U1016 ( .A1(n1248), .A2(n1250), .ZN(n1311) );
INV_X1 U1017 ( .A(n1106), .ZN(n1248) );
XOR2_X1 U1018 ( .A(G125), .B(G140), .Z(n1106) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1266), .ZN(n1309) );
NOR2_X1 U1020 ( .A1(n1314), .A2(n1289), .ZN(n1266) );
INV_X1 U1021 ( .A(G234), .ZN(n1314) );
NAND2_X1 U1022 ( .A1(KEYINPUT13), .A2(n1296), .ZN(n1307) );
INV_X1 U1023 ( .A(G128), .ZN(n1296) );
XNOR2_X1 U1024 ( .A(G110), .B(n1315), .ZN(n1305) );
XOR2_X1 U1025 ( .A(G137), .B(G119), .Z(n1315) );
NAND2_X1 U1026 ( .A1(G902), .A2(G217), .ZN(n1301) );
INV_X1 U1027 ( .A(n1235), .ZN(n1241) );
XOR2_X1 U1028 ( .A(n1087), .B(n1089), .Z(n1235) );
INV_X1 U1029 ( .A(G472), .ZN(n1089) );
NAND2_X1 U1030 ( .A1(n1316), .A2(n1262), .ZN(n1087) );
XNOR2_X1 U1031 ( .A(n1317), .B(n1318), .ZN(n1316) );
INV_X1 U1032 ( .A(n1149), .ZN(n1318) );
XNOR2_X1 U1033 ( .A(n1319), .B(n1320), .ZN(n1149) );
XOR2_X1 U1034 ( .A(n1291), .B(n1321), .Z(n1319) );
NOR2_X1 U1035 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XOR2_X1 U1036 ( .A(n1324), .B(KEYINPUT36), .Z(n1323) );
NAND2_X1 U1037 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1038 ( .A(n1327), .B(KEYINPUT40), .Z(n1325) );
NOR2_X1 U1039 ( .A1(n1326), .A2(n1327), .ZN(n1322) );
NAND2_X1 U1040 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NAND2_X1 U1041 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
OR3_X1 U1042 ( .A1(n1276), .A2(G119), .A3(n1331), .ZN(n1328) );
INV_X1 U1043 ( .A(KEYINPUT47), .ZN(n1331) );
INV_X1 U1044 ( .A(G116), .ZN(n1276) );
INV_X1 U1045 ( .A(G113), .ZN(n1326) );
XNOR2_X1 U1046 ( .A(n1109), .B(KEYINPUT9), .ZN(n1291) );
XOR2_X1 U1047 ( .A(G131), .B(n1332), .Z(n1109) );
XOR2_X1 U1048 ( .A(G137), .B(G134), .Z(n1332) );
XNOR2_X1 U1049 ( .A(G101), .B(n1333), .ZN(n1317) );
NOR2_X1 U1050 ( .A1(KEYINPUT57), .A2(n1151), .ZN(n1333) );
NAND2_X1 U1051 ( .A1(G210), .A2(n1258), .ZN(n1151) );
NOR2_X1 U1052 ( .A1(n1289), .A2(G237), .ZN(n1258) );
NOR2_X1 U1053 ( .A1(n1065), .A2(n1064), .ZN(n1176) );
AND2_X1 U1054 ( .A1(G214), .A2(n1334), .ZN(n1064) );
INV_X1 U1055 ( .A(n1216), .ZN(n1065) );
XNOR2_X1 U1056 ( .A(n1079), .B(n1082), .ZN(n1216) );
AND2_X1 U1057 ( .A1(G210), .A2(n1334), .ZN(n1082) );
NAND2_X1 U1058 ( .A1(n1335), .A2(n1262), .ZN(n1334) );
INV_X1 U1059 ( .A(G237), .ZN(n1335) );
NAND2_X1 U1060 ( .A1(n1336), .A2(n1262), .ZN(n1079) );
INV_X1 U1061 ( .A(G902), .ZN(n1262) );
XOR2_X1 U1062 ( .A(n1165), .B(n1337), .Z(n1336) );
XNOR2_X1 U1063 ( .A(n1338), .B(n1204), .ZN(n1337) );
INV_X1 U1064 ( .A(G125), .ZN(n1204) );
NAND2_X1 U1065 ( .A1(KEYINPUT12), .A2(n1202), .ZN(n1338) );
NOR2_X1 U1066 ( .A1(n1339), .A2(n1289), .ZN(n1202) );
XOR2_X1 U1067 ( .A(G953), .B(KEYINPUT0), .Z(n1289) );
INV_X1 U1068 ( .A(G224), .ZN(n1339) );
XNOR2_X1 U1069 ( .A(n1115), .B(n1320), .ZN(n1165) );
XNOR2_X1 U1070 ( .A(n1250), .B(n1272), .ZN(n1320) );
XNOR2_X1 U1071 ( .A(G128), .B(n1257), .ZN(n1272) );
INV_X1 U1072 ( .A(G143), .ZN(n1257) );
INV_X1 U1073 ( .A(G146), .ZN(n1250) );
XNOR2_X1 U1074 ( .A(n1340), .B(n1341), .ZN(n1115) );
XOR2_X1 U1075 ( .A(G107), .B(n1342), .Z(n1341) );
NOR2_X1 U1076 ( .A1(KEYINPUT52), .A2(n1330), .ZN(n1342) );
XNOR2_X1 U1077 ( .A(G116), .B(G119), .ZN(n1330) );
XNOR2_X1 U1078 ( .A(n1247), .B(n1156), .ZN(n1340) );
XNOR2_X1 U1079 ( .A(n1152), .B(G110), .ZN(n1156) );
INV_X1 U1080 ( .A(G101), .ZN(n1152) );
XOR2_X1 U1081 ( .A(G104), .B(n1343), .Z(n1247) );
XNOR2_X1 U1082 ( .A(n1236), .B(G113), .ZN(n1343) );
INV_X1 U1083 ( .A(G122), .ZN(n1236) );
endmodule


