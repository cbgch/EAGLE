//Key = 0011001000101101110101000110001100101001010101010010010100101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417;

XNOR2_X1 U770 ( .A(G107), .B(n1067), .ZN(G9) );
NAND4_X1 U771 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(G75) );
NAND3_X1 U772 ( .A1(n1072), .A2(n1073), .A3(G952), .ZN(n1071) );
NAND2_X1 U773 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NAND4_X1 U774 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1075) );
NAND2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NAND2_X1 U776 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U777 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
INV_X1 U779 ( .A(n1088), .ZN(n1084) );
NAND2_X1 U780 ( .A1(n1089), .A2(n1090), .ZN(n1080) );
NAND2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U782 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND3_X1 U783 ( .A1(n1082), .A2(n1095), .A3(n1089), .ZN(n1074) );
NAND2_X1 U784 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U785 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U786 ( .A(KEYINPUT42), .B(n1076), .Z(n1099) );
NAND3_X1 U787 ( .A1(n1100), .A2(n1101), .A3(n1077), .ZN(n1096) );
OR2_X1 U788 ( .A1(n1079), .A2(n1076), .ZN(n1101) );
OR3_X1 U789 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1100) );
NOR2_X1 U790 ( .A1(G953), .A2(n1105), .ZN(n1070) );
NOR4_X1 U791 ( .A1(n1106), .A2(n1107), .A3(n1104), .A4(n1108), .ZN(n1105) );
NOR2_X1 U792 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U793 ( .A(n1111), .B(KEYINPUT35), .Z(n1110) );
NOR2_X1 U794 ( .A1(G902), .A2(n1112), .ZN(n1109) );
NAND3_X1 U795 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1107) );
NAND4_X1 U796 ( .A1(n1116), .A2(n1117), .A3(n1089), .A4(n1118), .ZN(n1106) );
NOR2_X1 U797 ( .A1(n1094), .A2(n1119), .ZN(n1118) );
NAND2_X1 U798 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
XOR2_X1 U799 ( .A(n1122), .B(KEYINPUT13), .Z(n1120) );
NAND2_X1 U800 ( .A1(n1123), .A2(n1124), .ZN(n1116) );
XOR2_X1 U801 ( .A(n1122), .B(KEYINPUT14), .Z(n1123) );
XOR2_X1 U802 ( .A(n1125), .B(n1126), .Z(G72) );
NOR2_X1 U803 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U804 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
XOR2_X1 U805 ( .A(n1131), .B(n1132), .Z(n1125) );
NOR2_X1 U806 ( .A1(n1068), .A2(G953), .ZN(n1132) );
NAND2_X1 U807 ( .A1(KEYINPUT26), .A2(n1133), .ZN(n1131) );
NAND2_X1 U808 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND2_X1 U809 ( .A1(n1136), .A2(G953), .ZN(n1135) );
XOR2_X1 U810 ( .A(n1130), .B(KEYINPUT32), .Z(n1136) );
XOR2_X1 U811 ( .A(n1137), .B(n1138), .Z(n1134) );
XOR2_X1 U812 ( .A(n1139), .B(G125), .Z(n1138) );
NAND3_X1 U813 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
OR2_X1 U814 ( .A1(n1143), .A2(KEYINPUT21), .ZN(n1142) );
NAND3_X1 U815 ( .A1(KEYINPUT21), .A2(n1144), .A3(n1145), .ZN(n1141) );
OR2_X1 U816 ( .A1(n1145), .A2(n1144), .ZN(n1140) );
NOR2_X1 U817 ( .A1(KEYINPUT5), .A2(n1146), .ZN(n1144) );
XOR2_X1 U818 ( .A(n1147), .B(KEYINPUT40), .Z(n1137) );
NAND2_X1 U819 ( .A1(n1148), .A2(n1149), .ZN(G69) );
NAND2_X1 U820 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND3_X1 U821 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1150) );
XNOR2_X1 U822 ( .A(KEYINPUT6), .B(n1069), .ZN(n1154) );
OR2_X1 U823 ( .A1(n1128), .A2(G224), .ZN(n1152) );
NAND2_X1 U824 ( .A1(n1155), .A2(n1156), .ZN(n1148) );
NAND2_X1 U825 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
OR2_X1 U826 ( .A1(n1069), .A2(KEYINPUT6), .ZN(n1158) );
NAND2_X1 U827 ( .A1(KEYINPUT6), .A2(n1159), .ZN(n1157) );
NAND2_X1 U828 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U829 ( .A1(n1069), .A2(n1128), .ZN(n1161) );
NAND2_X1 U830 ( .A1(G953), .A2(G224), .ZN(n1160) );
INV_X1 U831 ( .A(n1151), .ZN(n1155) );
NAND3_X1 U832 ( .A1(n1162), .A2(n1163), .A3(n1153), .ZN(n1151) );
INV_X1 U833 ( .A(n1164), .ZN(n1153) );
NAND2_X1 U834 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
INV_X1 U835 ( .A(n1167), .ZN(n1166) );
NAND2_X1 U836 ( .A1(n1168), .A2(n1169), .ZN(n1165) );
OR2_X1 U837 ( .A1(n1170), .A2(KEYINPUT7), .ZN(n1169) );
NAND2_X1 U838 ( .A1(KEYINPUT7), .A2(n1171), .ZN(n1168) );
INV_X1 U839 ( .A(n1172), .ZN(n1171) );
NAND2_X1 U840 ( .A1(n1167), .A2(n1170), .ZN(n1162) );
NOR2_X1 U841 ( .A1(KEYINPUT54), .A2(n1172), .ZN(n1170) );
XOR2_X1 U842 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U843 ( .A(n1175), .B(KEYINPUT51), .Z(n1173) );
NOR2_X1 U844 ( .A1(n1176), .A2(n1177), .ZN(G66) );
XNOR2_X1 U845 ( .A(n1178), .B(n1179), .ZN(n1177) );
NOR3_X1 U846 ( .A1(n1180), .A2(KEYINPUT52), .A3(n1181), .ZN(n1179) );
XOR2_X1 U847 ( .A(KEYINPUT19), .B(G217), .Z(n1180) );
NOR2_X1 U848 ( .A1(n1176), .A2(n1182), .ZN(G63) );
XOR2_X1 U849 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND3_X1 U850 ( .A1(n1185), .A2(G478), .A3(KEYINPUT30), .ZN(n1183) );
NOR2_X1 U851 ( .A1(n1176), .A2(n1186), .ZN(G60) );
XOR2_X1 U852 ( .A(n1112), .B(n1187), .Z(n1186) );
NOR2_X1 U853 ( .A1(n1111), .A2(n1181), .ZN(n1187) );
NAND3_X1 U854 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(G6) );
OR2_X1 U855 ( .A1(n1191), .A2(KEYINPUT58), .ZN(n1190) );
NAND3_X1 U856 ( .A1(KEYINPUT58), .A2(n1191), .A3(G104), .ZN(n1189) );
NAND2_X1 U857 ( .A1(n1192), .A2(n1193), .ZN(n1188) );
NAND2_X1 U858 ( .A1(n1194), .A2(KEYINPUT58), .ZN(n1192) );
XOR2_X1 U859 ( .A(n1191), .B(KEYINPUT38), .Z(n1194) );
NOR2_X1 U860 ( .A1(n1176), .A2(n1195), .ZN(G57) );
XNOR2_X1 U861 ( .A(n1196), .B(n1197), .ZN(n1195) );
XOR2_X1 U862 ( .A(n1198), .B(n1199), .Z(n1196) );
AND2_X1 U863 ( .A1(G472), .A2(n1185), .ZN(n1199) );
NAND2_X1 U864 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
NAND2_X1 U865 ( .A1(n1202), .A2(n1203), .ZN(n1200) );
XNOR2_X1 U866 ( .A(n1204), .B(KEYINPUT62), .ZN(n1202) );
NOR2_X1 U867 ( .A1(n1176), .A2(n1205), .ZN(G54) );
XOR2_X1 U868 ( .A(n1206), .B(n1207), .Z(n1205) );
AND2_X1 U869 ( .A1(G469), .A2(n1185), .ZN(n1207) );
NOR2_X1 U870 ( .A1(n1208), .A2(n1209), .ZN(n1206) );
XOR2_X1 U871 ( .A(n1210), .B(KEYINPUT17), .Z(n1209) );
NAND2_X1 U872 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NOR2_X1 U873 ( .A1(n1212), .A2(n1211), .ZN(n1208) );
XOR2_X1 U874 ( .A(n1213), .B(n1203), .Z(n1211) );
XOR2_X1 U875 ( .A(n1146), .B(n1214), .Z(n1213) );
NOR2_X1 U876 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
AND2_X1 U877 ( .A1(KEYINPUT31), .A2(n1217), .ZN(n1216) );
NOR2_X1 U878 ( .A1(KEYINPUT16), .A2(n1217), .ZN(n1215) );
XNOR2_X1 U879 ( .A(n1218), .B(n1219), .ZN(n1212) );
NAND2_X1 U880 ( .A1(KEYINPUT12), .A2(n1220), .ZN(n1218) );
NOR2_X1 U881 ( .A1(n1176), .A2(n1221), .ZN(G51) );
NOR3_X1 U882 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1221) );
NOR3_X1 U883 ( .A1(n1225), .A2(n1181), .A3(n1226), .ZN(n1224) );
INV_X1 U884 ( .A(n1185), .ZN(n1181) );
NOR2_X1 U885 ( .A1(n1227), .A2(n1228), .ZN(n1185) );
NOR2_X1 U886 ( .A1(n1229), .A2(n1230), .ZN(n1223) );
INV_X1 U887 ( .A(n1225), .ZN(n1230) );
NOR2_X1 U888 ( .A1(n1228), .A2(n1226), .ZN(n1229) );
NAND2_X1 U889 ( .A1(KEYINPUT41), .A2(n1124), .ZN(n1226) );
INV_X1 U890 ( .A(n1121), .ZN(n1124) );
AND2_X1 U891 ( .A1(n1069), .A2(n1231), .ZN(n1228) );
XOR2_X1 U892 ( .A(KEYINPUT1), .B(n1068), .Z(n1231) );
AND4_X1 U893 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1068) );
NOR4_X1 U894 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235) );
INV_X1 U895 ( .A(n1240), .ZN(n1236) );
NAND4_X1 U896 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1234) );
NOR2_X1 U897 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND2_X1 U898 ( .A1(n1247), .A2(n1248), .ZN(n1242) );
NAND2_X1 U899 ( .A1(n1249), .A2(n1250), .ZN(n1241) );
NAND2_X1 U900 ( .A1(n1077), .A2(n1079), .ZN(n1250) );
INV_X1 U901 ( .A(n1251), .ZN(n1077) );
AND4_X1 U902 ( .A1(n1252), .A2(n1191), .A3(n1253), .A4(n1254), .ZN(n1069) );
AND4_X1 U903 ( .A1(n1067), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1254) );
NAND3_X1 U904 ( .A1(n1102), .A2(n1082), .A3(n1258), .ZN(n1067) );
AND2_X1 U905 ( .A1(n1259), .A2(n1260), .ZN(n1253) );
NAND3_X1 U906 ( .A1(n1258), .A2(n1082), .A3(n1103), .ZN(n1191) );
NAND3_X1 U907 ( .A1(n1103), .A2(n1261), .A3(n1262), .ZN(n1252) );
XOR2_X1 U908 ( .A(KEYINPUT29), .B(n1243), .Z(n1261) );
NOR2_X1 U909 ( .A1(n1128), .A2(G952), .ZN(n1176) );
XNOR2_X1 U910 ( .A(G146), .B(n1232), .ZN(G48) );
NAND3_X1 U911 ( .A1(n1263), .A2(n1103), .A3(n1264), .ZN(n1232) );
INV_X1 U912 ( .A(n1265), .ZN(n1103) );
XOR2_X1 U913 ( .A(n1266), .B(n1267), .Z(G45) );
XOR2_X1 U914 ( .A(KEYINPUT53), .B(G143), .Z(n1267) );
NAND3_X1 U915 ( .A1(n1243), .A2(n1263), .A3(n1268), .ZN(n1266) );
XNOR2_X1 U916 ( .A(n1269), .B(KEYINPUT3), .ZN(n1268) );
XOR2_X1 U917 ( .A(n1147), .B(n1233), .Z(G42) );
NAND2_X1 U918 ( .A1(n1270), .A2(n1271), .ZN(n1233) );
XOR2_X1 U919 ( .A(G137), .B(n1239), .Z(G39) );
AND3_X1 U920 ( .A1(n1270), .A2(n1264), .A3(n1076), .ZN(n1239) );
XNOR2_X1 U921 ( .A(G134), .B(n1272), .ZN(G36) );
NAND3_X1 U922 ( .A1(n1270), .A2(n1102), .A3(n1273), .ZN(n1272) );
XOR2_X1 U923 ( .A(n1091), .B(KEYINPUT34), .Z(n1273) );
XOR2_X1 U924 ( .A(G131), .B(n1238), .Z(G33) );
AND2_X1 U925 ( .A1(n1270), .A2(n1274), .ZN(n1238) );
NOR3_X1 U926 ( .A1(n1251), .A2(n1104), .A3(n1246), .ZN(n1270) );
INV_X1 U927 ( .A(n1079), .ZN(n1104) );
NAND2_X1 U928 ( .A1(n1275), .A2(n1276), .ZN(G30) );
NAND2_X1 U929 ( .A1(n1237), .A2(n1277), .ZN(n1276) );
XOR2_X1 U930 ( .A(KEYINPUT2), .B(n1278), .Z(n1275) );
NOR2_X1 U931 ( .A1(n1237), .A2(n1277), .ZN(n1278) );
AND3_X1 U932 ( .A1(n1263), .A2(n1102), .A3(n1264), .ZN(n1237) );
NOR2_X1 U933 ( .A1(n1246), .A2(n1248), .ZN(n1263) );
NAND2_X1 U934 ( .A1(n1279), .A2(n1088), .ZN(n1246) );
XOR2_X1 U935 ( .A(n1260), .B(n1280), .Z(G3) );
XOR2_X1 U936 ( .A(KEYINPUT39), .B(G101), .Z(n1280) );
NAND3_X1 U937 ( .A1(n1243), .A2(n1258), .A3(n1076), .ZN(n1260) );
XOR2_X1 U938 ( .A(n1281), .B(n1240), .Z(G27) );
NAND4_X1 U939 ( .A1(n1089), .A2(n1279), .A3(n1271), .A4(n1098), .ZN(n1240) );
NOR3_X1 U940 ( .A1(n1282), .A2(n1283), .A3(n1265), .ZN(n1271) );
AND3_X1 U941 ( .A1(n1284), .A2(n1285), .A3(n1073), .ZN(n1279) );
OR2_X1 U942 ( .A1(G952), .A2(G953), .ZN(n1285) );
NAND2_X1 U943 ( .A1(G953), .A2(n1286), .ZN(n1284) );
NAND2_X1 U944 ( .A1(G902), .A2(n1130), .ZN(n1286) );
INV_X1 U945 ( .A(G900), .ZN(n1130) );
XOR2_X1 U946 ( .A(n1287), .B(n1259), .Z(G24) );
NAND3_X1 U947 ( .A1(n1262), .A2(n1082), .A3(n1269), .ZN(n1259) );
NOR2_X1 U948 ( .A1(n1245), .A2(n1249), .ZN(n1269) );
INV_X1 U949 ( .A(n1247), .ZN(n1249) );
NOR2_X1 U950 ( .A1(n1094), .A2(n1282), .ZN(n1082) );
NAND2_X1 U951 ( .A1(n1288), .A2(n1289), .ZN(G21) );
NAND2_X1 U952 ( .A1(G119), .A2(n1257), .ZN(n1289) );
XOR2_X1 U953 ( .A(n1290), .B(KEYINPUT20), .Z(n1288) );
OR2_X1 U954 ( .A1(n1257), .A2(G119), .ZN(n1290) );
NAND3_X1 U955 ( .A1(n1076), .A2(n1264), .A3(n1262), .ZN(n1257) );
NOR2_X1 U956 ( .A1(n1093), .A2(n1283), .ZN(n1264) );
XNOR2_X1 U957 ( .A(G116), .B(n1256), .ZN(G18) );
NAND3_X1 U958 ( .A1(n1243), .A2(n1102), .A3(n1262), .ZN(n1256) );
NOR2_X1 U959 ( .A1(n1247), .A2(n1245), .ZN(n1102) );
INV_X1 U960 ( .A(n1091), .ZN(n1243) );
XOR2_X1 U961 ( .A(G113), .B(n1291), .Z(G15) );
AND2_X1 U962 ( .A1(n1274), .A2(n1262), .ZN(n1291) );
AND2_X1 U963 ( .A1(n1089), .A2(n1292), .ZN(n1262) );
NOR2_X1 U964 ( .A1(n1293), .A2(n1086), .ZN(n1089) );
INV_X1 U965 ( .A(n1087), .ZN(n1293) );
NOR2_X1 U966 ( .A1(n1091), .A2(n1265), .ZN(n1274) );
NAND2_X1 U967 ( .A1(n1245), .A2(n1247), .ZN(n1265) );
INV_X1 U968 ( .A(n1294), .ZN(n1245) );
NAND2_X1 U969 ( .A1(n1283), .A2(n1282), .ZN(n1091) );
INV_X1 U970 ( .A(n1093), .ZN(n1282) );
INV_X1 U971 ( .A(n1094), .ZN(n1283) );
XOR2_X1 U972 ( .A(n1295), .B(n1255), .Z(G12) );
NAND4_X1 U973 ( .A1(n1076), .A2(n1258), .A3(n1093), .A4(n1094), .ZN(n1255) );
NAND3_X1 U974 ( .A1(n1296), .A2(n1297), .A3(n1298), .ZN(n1094) );
NAND2_X1 U975 ( .A1(G217), .A2(G902), .ZN(n1298) );
NAND3_X1 U976 ( .A1(n1178), .A2(n1227), .A3(n1299), .ZN(n1297) );
OR2_X1 U977 ( .A1(n1299), .A2(n1178), .ZN(n1296) );
AND3_X1 U978 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1178) );
NAND2_X1 U979 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
INV_X1 U980 ( .A(KEYINPUT63), .ZN(n1304) );
NAND3_X1 U981 ( .A1(KEYINPUT63), .A2(n1305), .A3(n1306), .ZN(n1301) );
OR2_X1 U982 ( .A1(n1306), .A2(n1305), .ZN(n1300) );
NOR2_X1 U983 ( .A1(KEYINPUT28), .A2(n1303), .ZN(n1305) );
XOR2_X1 U984 ( .A(n1307), .B(n1308), .Z(n1303) );
NOR3_X1 U985 ( .A1(n1309), .A2(n1310), .A3(n1311), .ZN(n1308) );
NOR2_X1 U986 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
INV_X1 U987 ( .A(KEYINPUT50), .ZN(n1312) );
NOR3_X1 U988 ( .A1(KEYINPUT50), .A2(G140), .A3(G125), .ZN(n1310) );
XOR2_X1 U989 ( .A(KEYINPUT9), .B(n1314), .Z(n1309) );
NOR2_X1 U990 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XOR2_X1 U991 ( .A(KEYINPUT49), .B(G125), .Z(n1316) );
XOR2_X1 U992 ( .A(n1147), .B(KEYINPUT44), .Z(n1315) );
XNOR2_X1 U993 ( .A(n1317), .B(n1318), .ZN(n1307) );
NOR2_X1 U994 ( .A1(KEYINPUT18), .A2(G146), .ZN(n1318) );
NOR3_X1 U995 ( .A1(n1319), .A2(KEYINPUT59), .A3(n1320), .ZN(n1317) );
NOR2_X1 U996 ( .A1(G110), .A2(n1321), .ZN(n1320) );
XOR2_X1 U997 ( .A(G128), .B(G119), .Z(n1321) );
XOR2_X1 U998 ( .A(KEYINPUT57), .B(n1322), .Z(n1319) );
NOR2_X1 U999 ( .A1(n1323), .A2(n1295), .ZN(n1322) );
XOR2_X1 U1000 ( .A(G119), .B(n1277), .Z(n1323) );
INV_X1 U1001 ( .A(G128), .ZN(n1277) );
XNOR2_X1 U1002 ( .A(n1324), .B(G137), .ZN(n1306) );
NAND2_X1 U1003 ( .A1(n1325), .A2(G221), .ZN(n1324) );
NAND2_X1 U1004 ( .A1(G217), .A2(n1326), .ZN(n1299) );
XNOR2_X1 U1005 ( .A(n1119), .B(KEYINPUT4), .ZN(n1093) );
XNOR2_X1 U1006 ( .A(n1327), .B(G472), .ZN(n1119) );
NAND4_X1 U1007 ( .A1(n1328), .A2(n1227), .A3(n1329), .A4(n1330), .ZN(n1327) );
NAND3_X1 U1008 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(n1330) );
INV_X1 U1009 ( .A(KEYINPUT0), .ZN(n1332) );
OR2_X1 U1010 ( .A1(n1333), .A2(n1331), .ZN(n1329) );
AND3_X1 U1011 ( .A1(n1334), .A2(n1335), .A3(n1201), .ZN(n1331) );
NAND2_X1 U1012 ( .A1(n1145), .A2(n1204), .ZN(n1201) );
OR3_X1 U1013 ( .A1(n1145), .A2(n1204), .A3(KEYINPUT27), .ZN(n1335) );
NAND2_X1 U1014 ( .A1(KEYINPUT27), .A2(n1204), .ZN(n1334) );
XOR2_X1 U1015 ( .A(n1336), .B(n1337), .Z(n1204) );
XOR2_X1 U1016 ( .A(KEYINPUT8), .B(n1174), .Z(n1337) );
NOR2_X1 U1017 ( .A1(KEYINPUT56), .A2(n1197), .ZN(n1333) );
NAND2_X1 U1018 ( .A1(KEYINPUT0), .A2(n1197), .ZN(n1328) );
XOR2_X1 U1019 ( .A(n1338), .B(G101), .Z(n1197) );
NAND2_X1 U1020 ( .A1(n1339), .A2(G210), .ZN(n1338) );
AND2_X1 U1021 ( .A1(n1292), .A2(n1088), .ZN(n1258) );
NOR2_X1 U1022 ( .A1(n1087), .A2(n1086), .ZN(n1088) );
AND2_X1 U1023 ( .A1(G221), .A2(n1340), .ZN(n1086) );
NAND2_X1 U1024 ( .A1(G234), .A2(n1227), .ZN(n1340) );
XOR2_X1 U1025 ( .A(n1341), .B(G469), .Z(n1087) );
NAND2_X1 U1026 ( .A1(n1342), .A2(n1227), .ZN(n1341) );
XOR2_X1 U1027 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1028 ( .A(n1345), .B(n1220), .ZN(n1344) );
XOR2_X1 U1029 ( .A(n1295), .B(n1147), .Z(n1220) );
NAND2_X1 U1030 ( .A1(n1346), .A2(KEYINPUT45), .ZN(n1345) );
XOR2_X1 U1031 ( .A(n1347), .B(n1143), .Z(n1346) );
INV_X1 U1032 ( .A(n1146), .ZN(n1143) );
XOR2_X1 U1033 ( .A(n1348), .B(n1349), .Z(n1146) );
XNOR2_X1 U1034 ( .A(KEYINPUT25), .B(n1350), .ZN(n1348) );
NOR2_X1 U1035 ( .A1(G143), .A2(KEYINPUT22), .ZN(n1350) );
XNOR2_X1 U1036 ( .A(n1351), .B(n1217), .ZN(n1347) );
XOR2_X1 U1037 ( .A(G101), .B(n1352), .Z(n1217) );
NAND2_X1 U1038 ( .A1(KEYINPUT36), .A2(n1203), .ZN(n1351) );
INV_X1 U1039 ( .A(n1145), .ZN(n1203) );
XNOR2_X1 U1040 ( .A(G131), .B(n1353), .ZN(n1145) );
XOR2_X1 U1041 ( .A(G137), .B(G134), .Z(n1353) );
XNOR2_X1 U1042 ( .A(n1219), .B(KEYINPUT33), .ZN(n1343) );
NOR2_X1 U1043 ( .A1(n1129), .A2(G953), .ZN(n1219) );
INV_X1 U1044 ( .A(G227), .ZN(n1129) );
AND3_X1 U1045 ( .A1(n1354), .A2(n1073), .A3(n1098), .ZN(n1292) );
INV_X1 U1046 ( .A(n1248), .ZN(n1098) );
NAND2_X1 U1047 ( .A1(n1251), .A2(n1079), .ZN(n1248) );
NAND2_X1 U1048 ( .A1(G214), .A2(n1355), .ZN(n1079) );
XOR2_X1 U1049 ( .A(n1356), .B(n1222), .Z(n1251) );
INV_X1 U1050 ( .A(n1122), .ZN(n1222) );
NAND2_X1 U1051 ( .A1(n1225), .A2(n1227), .ZN(n1122) );
XOR2_X1 U1052 ( .A(n1357), .B(n1358), .Z(n1225) );
XOR2_X1 U1053 ( .A(n1359), .B(n1360), .Z(n1358) );
XOR2_X1 U1054 ( .A(n1175), .B(G125), .Z(n1360) );
NAND2_X1 U1055 ( .A1(n1361), .A2(n1362), .ZN(n1175) );
NAND2_X1 U1056 ( .A1(n1352), .A2(n1363), .ZN(n1362) );
NAND2_X1 U1057 ( .A1(G101), .A2(n1364), .ZN(n1363) );
OR2_X1 U1058 ( .A1(n1365), .A2(KEYINPUT11), .ZN(n1364) );
NAND3_X1 U1059 ( .A1(n1366), .A2(n1367), .A3(n1365), .ZN(n1361) );
INV_X1 U1060 ( .A(KEYINPUT23), .ZN(n1365) );
OR2_X1 U1061 ( .A1(G101), .A2(KEYINPUT11), .ZN(n1367) );
NAND2_X1 U1062 ( .A1(G101), .A2(n1368), .ZN(n1366) );
OR2_X1 U1063 ( .A1(n1352), .A2(KEYINPUT11), .ZN(n1368) );
XNOR2_X1 U1064 ( .A(G107), .B(G104), .ZN(n1352) );
NAND2_X1 U1065 ( .A1(G224), .A2(n1128), .ZN(n1359) );
XOR2_X1 U1066 ( .A(n1369), .B(n1167), .Z(n1357) );
XNOR2_X1 U1067 ( .A(n1295), .B(G122), .ZN(n1167) );
XOR2_X1 U1068 ( .A(n1370), .B(n1336), .Z(n1369) );
XNOR2_X1 U1069 ( .A(n1371), .B(n1349), .ZN(n1336) );
XOR2_X1 U1070 ( .A(G146), .B(G128), .Z(n1349) );
INV_X1 U1071 ( .A(G143), .ZN(n1371) );
NAND2_X1 U1072 ( .A1(KEYINPUT10), .A2(n1174), .ZN(n1370) );
XOR2_X1 U1073 ( .A(n1372), .B(n1373), .Z(n1174) );
XNOR2_X1 U1074 ( .A(G116), .B(G119), .ZN(n1372) );
NAND2_X1 U1075 ( .A1(KEYINPUT15), .A2(n1121), .ZN(n1356) );
NAND2_X1 U1076 ( .A1(G210), .A2(n1355), .ZN(n1121) );
NAND2_X1 U1077 ( .A1(n1374), .A2(n1227), .ZN(n1355) );
INV_X1 U1078 ( .A(G237), .ZN(n1374) );
NAND2_X1 U1079 ( .A1(G234), .A2(n1375), .ZN(n1073) );
XOR2_X1 U1080 ( .A(KEYINPUT24), .B(G237), .Z(n1375) );
NAND2_X1 U1081 ( .A1(n1376), .A2(n1377), .ZN(n1354) );
NAND2_X1 U1082 ( .A1(G902), .A2(n1164), .ZN(n1377) );
NOR2_X1 U1083 ( .A1(G898), .A2(n1128), .ZN(n1164) );
NAND2_X1 U1084 ( .A1(G952), .A2(n1128), .ZN(n1376) );
INV_X1 U1085 ( .A(G953), .ZN(n1128) );
NOR2_X1 U1086 ( .A1(n1294), .A2(n1247), .ZN(n1076) );
NAND2_X1 U1087 ( .A1(n1115), .A2(n1378), .ZN(n1247) );
NAND2_X1 U1088 ( .A1(G475), .A2(n1379), .ZN(n1378) );
NAND2_X1 U1089 ( .A1(n1380), .A2(n1227), .ZN(n1379) );
NAND3_X1 U1090 ( .A1(n1111), .A2(n1227), .A3(n1380), .ZN(n1115) );
INV_X1 U1091 ( .A(n1112), .ZN(n1380) );
XOR2_X1 U1092 ( .A(n1381), .B(n1382), .Z(n1112) );
XOR2_X1 U1093 ( .A(n1383), .B(n1384), .Z(n1382) );
XOR2_X1 U1094 ( .A(n1385), .B(n1386), .Z(n1384) );
AND2_X1 U1095 ( .A1(G214), .A2(n1339), .ZN(n1386) );
NOR2_X1 U1096 ( .A1(G953), .A2(G237), .ZN(n1339) );
NAND3_X1 U1097 ( .A1(n1387), .A2(n1388), .A3(n1389), .ZN(n1385) );
NAND2_X1 U1098 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
NAND3_X1 U1099 ( .A1(n1392), .A2(n1393), .A3(n1394), .ZN(n1391) );
NAND2_X1 U1100 ( .A1(KEYINPUT46), .A2(n1395), .ZN(n1394) );
OR2_X1 U1101 ( .A1(G122), .A2(KEYINPUT55), .ZN(n1393) );
NAND2_X1 U1102 ( .A1(KEYINPUT55), .A2(n1396), .ZN(n1392) );
NAND2_X1 U1103 ( .A1(n1287), .A2(n1397), .ZN(n1396) );
NAND2_X1 U1104 ( .A1(KEYINPUT37), .A2(n1398), .ZN(n1397) );
INV_X1 U1105 ( .A(n1373), .ZN(n1390) );
NAND4_X1 U1106 ( .A1(n1287), .A2(n1395), .A3(n1373), .A4(n1398), .ZN(n1388) );
INV_X1 U1107 ( .A(KEYINPUT46), .ZN(n1398) );
INV_X1 U1108 ( .A(KEYINPUT37), .ZN(n1395) );
NAND2_X1 U1109 ( .A1(KEYINPUT46), .A2(n1399), .ZN(n1387) );
NAND2_X1 U1110 ( .A1(n1287), .A2(n1400), .ZN(n1399) );
NAND2_X1 U1111 ( .A1(KEYINPUT37), .A2(n1373), .ZN(n1400) );
XNOR2_X1 U1112 ( .A(G113), .B(KEYINPUT60), .ZN(n1373) );
INV_X1 U1113 ( .A(G122), .ZN(n1287) );
NAND2_X1 U1114 ( .A1(n1401), .A2(n1313), .ZN(n1383) );
NAND2_X1 U1115 ( .A1(G125), .A2(n1147), .ZN(n1313) );
INV_X1 U1116 ( .A(G140), .ZN(n1147) );
XOR2_X1 U1117 ( .A(n1402), .B(KEYINPUT48), .Z(n1401) );
NAND2_X1 U1118 ( .A1(G140), .A2(n1281), .ZN(n1402) );
INV_X1 U1119 ( .A(G125), .ZN(n1281) );
XOR2_X1 U1120 ( .A(n1403), .B(n1404), .Z(n1381) );
XOR2_X1 U1121 ( .A(G146), .B(G143), .Z(n1404) );
XOR2_X1 U1122 ( .A(G131), .B(n1193), .Z(n1403) );
INV_X1 U1123 ( .A(G104), .ZN(n1193) );
INV_X1 U1124 ( .A(G475), .ZN(n1111) );
NAND3_X1 U1125 ( .A1(n1405), .A2(n1406), .A3(n1113), .ZN(n1294) );
NAND3_X1 U1126 ( .A1(n1184), .A2(n1227), .A3(n1407), .ZN(n1113) );
NAND2_X1 U1127 ( .A1(n1408), .A2(KEYINPUT43), .ZN(n1406) );
INV_X1 U1128 ( .A(n1114), .ZN(n1408) );
NAND2_X1 U1129 ( .A1(n1409), .A2(n1410), .ZN(n1114) );
NAND2_X1 U1130 ( .A1(n1184), .A2(n1227), .ZN(n1410) );
INV_X1 U1131 ( .A(G902), .ZN(n1227) );
XNOR2_X1 U1132 ( .A(n1411), .B(n1412), .ZN(n1184) );
XOR2_X1 U1133 ( .A(n1413), .B(n1414), .Z(n1412) );
XOR2_X1 U1134 ( .A(G128), .B(G122), .Z(n1414) );
XOR2_X1 U1135 ( .A(G143), .B(G134), .Z(n1413) );
XOR2_X1 U1136 ( .A(n1415), .B(n1416), .Z(n1411) );
XOR2_X1 U1137 ( .A(G116), .B(G107), .Z(n1416) );
NAND2_X1 U1138 ( .A1(n1417), .A2(n1325), .ZN(n1415) );
NOR2_X1 U1139 ( .A1(n1326), .A2(G953), .ZN(n1325) );
INV_X1 U1140 ( .A(G234), .ZN(n1326) );
XNOR2_X1 U1141 ( .A(G217), .B(KEYINPUT47), .ZN(n1417) );
OR2_X1 U1142 ( .A1(n1409), .A2(KEYINPUT43), .ZN(n1405) );
INV_X1 U1143 ( .A(n1407), .ZN(n1409) );
XNOR2_X1 U1144 ( .A(G478), .B(KEYINPUT61), .ZN(n1407) );
INV_X1 U1145 ( .A(G110), .ZN(n1295) );
endmodule


