//Key = 1011010010111010100110001101001001100100110101110000000111100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
n1445, n1446;

XNOR2_X1 U805 ( .A(G107), .B(n1105), .ZN(G9) );
NOR2_X1 U806 ( .A1(n1106), .A2(n1107), .ZN(G75) );
NOR3_X1 U807 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1107) );
NOR2_X1 U808 ( .A1(n1111), .A2(n1112), .ZN(n1109) );
NOR2_X1 U809 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR2_X1 U810 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U811 ( .A1(n1117), .A2(n1118), .ZN(n1115) );
NOR2_X1 U812 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NOR2_X1 U813 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
NOR2_X1 U814 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U815 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NOR2_X1 U816 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
NOR2_X1 U817 ( .A1(n1129), .A2(n1130), .ZN(n1121) );
NOR2_X1 U818 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
NOR3_X1 U819 ( .A1(n1130), .A2(n1133), .A3(n1124), .ZN(n1117) );
NOR2_X1 U820 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NOR3_X1 U821 ( .A1(n1136), .A2(n1130), .A3(n1120), .ZN(n1113) );
INV_X1 U822 ( .A(n1137), .ZN(n1120) );
NAND3_X1 U823 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1136) );
NAND3_X1 U824 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1108) );
NAND4_X1 U825 ( .A1(n1144), .A2(n1137), .A3(n1145), .A4(n1146), .ZN(n1143) );
NOR3_X1 U826 ( .A1(n1130), .A2(n1147), .A3(n1124), .ZN(n1146) );
XOR2_X1 U827 ( .A(n1139), .B(KEYINPUT20), .Z(n1145) );
INV_X1 U828 ( .A(n1112), .ZN(n1144) );
NOR3_X1 U829 ( .A1(n1148), .A2(G953), .A3(G952), .ZN(n1106) );
INV_X1 U830 ( .A(n1141), .ZN(n1148) );
NAND4_X1 U831 ( .A1(n1139), .A2(n1128), .A3(n1149), .A4(n1150), .ZN(n1141) );
NOR3_X1 U832 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
XOR2_X1 U833 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U834 ( .A1(n1156), .A2(KEYINPUT28), .ZN(n1155) );
INV_X1 U835 ( .A(n1157), .ZN(n1156) );
NOR2_X1 U836 ( .A1(n1158), .A2(n1159), .ZN(n1152) );
NOR2_X1 U837 ( .A1(G902), .A2(n1160), .ZN(n1158) );
NAND3_X1 U838 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1151) );
XNOR2_X1 U839 ( .A(G475), .B(n1164), .ZN(n1163) );
NAND2_X1 U840 ( .A1(KEYINPUT10), .A2(n1165), .ZN(n1164) );
OR2_X1 U841 ( .A1(n1140), .A2(KEYINPUT44), .ZN(n1162) );
NAND2_X1 U842 ( .A1(KEYINPUT44), .A2(n1166), .ZN(n1161) );
NAND2_X1 U843 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NOR3_X1 U844 ( .A1(n1169), .A2(n1170), .A3(n1171), .ZN(n1149) );
XOR2_X1 U845 ( .A(n1172), .B(n1173), .Z(G72) );
XOR2_X1 U846 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U847 ( .A1(n1176), .A2(n1142), .ZN(n1175) );
NOR2_X1 U848 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XNOR2_X1 U849 ( .A(G227), .B(KEYINPUT29), .ZN(n1177) );
NAND2_X1 U850 ( .A1(n1179), .A2(n1180), .ZN(n1174) );
NAND2_X1 U851 ( .A1(G953), .A2(n1178), .ZN(n1180) );
XOR2_X1 U852 ( .A(n1181), .B(n1182), .Z(n1179) );
XOR2_X1 U853 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U854 ( .A1(G140), .A2(KEYINPUT22), .ZN(n1184) );
NAND2_X1 U855 ( .A1(n1185), .A2(n1186), .ZN(n1183) );
OR2_X1 U856 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U857 ( .A(n1189), .B(KEYINPUT50), .Z(n1185) );
NAND2_X1 U858 ( .A1(n1187), .A2(n1188), .ZN(n1189) );
XNOR2_X1 U859 ( .A(n1190), .B(G131), .ZN(n1187) );
NAND2_X1 U860 ( .A1(KEYINPUT2), .A2(n1191), .ZN(n1190) );
NAND2_X1 U861 ( .A1(n1142), .A2(n1192), .ZN(n1172) );
NAND2_X1 U862 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NAND2_X1 U863 ( .A1(n1195), .A2(n1196), .ZN(G69) );
NAND2_X1 U864 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
OR2_X1 U865 ( .A1(n1142), .A2(G224), .ZN(n1198) );
NAND3_X1 U866 ( .A1(G953), .A2(n1199), .A3(n1200), .ZN(n1195) );
INV_X1 U867 ( .A(n1197), .ZN(n1200) );
XNOR2_X1 U868 ( .A(n1201), .B(n1202), .ZN(n1197) );
NOR2_X1 U869 ( .A1(G953), .A2(n1203), .ZN(n1202) );
NOR2_X1 U870 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
XNOR2_X1 U871 ( .A(KEYINPUT62), .B(n1105), .ZN(n1205) );
NAND2_X1 U872 ( .A1(n1206), .A2(n1207), .ZN(n1201) );
NAND2_X1 U873 ( .A1(G953), .A2(n1208), .ZN(n1207) );
XOR2_X1 U874 ( .A(n1209), .B(n1210), .Z(n1206) );
NAND2_X1 U875 ( .A1(KEYINPUT0), .A2(n1211), .ZN(n1209) );
NAND2_X1 U876 ( .A1(G898), .A2(G224), .ZN(n1199) );
NOR2_X1 U877 ( .A1(n1212), .A2(n1213), .ZN(G66) );
XOR2_X1 U878 ( .A(KEYINPUT39), .B(n1214), .Z(n1213) );
XNOR2_X1 U879 ( .A(n1215), .B(n1216), .ZN(n1212) );
NOR2_X1 U880 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NOR2_X1 U881 ( .A1(n1214), .A2(n1219), .ZN(G63) );
XOR2_X1 U882 ( .A(n1220), .B(n1160), .Z(n1219) );
NOR2_X1 U883 ( .A1(n1159), .A2(n1218), .ZN(n1220) );
NOR2_X1 U884 ( .A1(n1214), .A2(n1221), .ZN(G60) );
NOR3_X1 U885 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1221) );
NOR3_X1 U886 ( .A1(n1225), .A2(n1226), .A3(n1218), .ZN(n1224) );
INV_X1 U887 ( .A(n1227), .ZN(n1225) );
NOR2_X1 U888 ( .A1(n1228), .A2(n1227), .ZN(n1223) );
AND2_X1 U889 ( .A1(n1110), .A2(G475), .ZN(n1228) );
NAND2_X1 U890 ( .A1(n1229), .A2(n1230), .ZN(G6) );
OR2_X1 U891 ( .A1(n1231), .A2(G104), .ZN(n1230) );
XOR2_X1 U892 ( .A(n1232), .B(KEYINPUT4), .Z(n1229) );
NAND2_X1 U893 ( .A1(G104), .A2(n1231), .ZN(n1232) );
NOR3_X1 U894 ( .A1(n1214), .A2(n1233), .A3(n1234), .ZN(G57) );
NOR2_X1 U895 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XOR2_X1 U896 ( .A(n1237), .B(n1238), .Z(n1236) );
AND3_X1 U897 ( .A1(n1235), .A2(n1239), .A3(n1240), .ZN(n1233) );
XNOR2_X1 U898 ( .A(n1241), .B(n1242), .ZN(n1235) );
NOR2_X1 U899 ( .A1(n1243), .A2(n1218), .ZN(n1242) );
NOR2_X1 U900 ( .A1(n1214), .A2(n1244), .ZN(G54) );
XOR2_X1 U901 ( .A(n1245), .B(n1246), .Z(n1244) );
XOR2_X1 U902 ( .A(n1247), .B(n1248), .Z(n1246) );
NOR3_X1 U903 ( .A1(n1249), .A2(KEYINPUT15), .A3(n1250), .ZN(n1248) );
NOR2_X1 U904 ( .A1(n1211), .A2(n1188), .ZN(n1250) );
XOR2_X1 U905 ( .A(KEYINPUT48), .B(n1251), .Z(n1249) );
NOR2_X1 U906 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NOR2_X1 U907 ( .A1(n1254), .A2(n1218), .ZN(n1247) );
NOR2_X1 U908 ( .A1(n1142), .A2(G952), .ZN(n1214) );
NOR2_X1 U909 ( .A1(n1255), .A2(n1256), .ZN(G51) );
XOR2_X1 U910 ( .A(n1257), .B(n1258), .Z(n1256) );
XNOR2_X1 U911 ( .A(n1259), .B(n1181), .ZN(n1258) );
XNOR2_X1 U912 ( .A(n1260), .B(n1261), .ZN(n1257) );
NOR2_X1 U913 ( .A1(n1157), .A2(n1218), .ZN(n1261) );
NAND2_X1 U914 ( .A1(G902), .A2(n1110), .ZN(n1218) );
NAND4_X1 U915 ( .A1(n1193), .A2(n1262), .A3(n1263), .A4(n1105), .ZN(n1110) );
NAND3_X1 U916 ( .A1(n1134), .A2(n1264), .A3(n1140), .ZN(n1105) );
XNOR2_X1 U917 ( .A(KEYINPUT61), .B(n1194), .ZN(n1263) );
NAND2_X1 U918 ( .A1(n1265), .A2(n1266), .ZN(n1194) );
XNOR2_X1 U919 ( .A(n1131), .B(KEYINPUT41), .ZN(n1265) );
INV_X1 U920 ( .A(n1204), .ZN(n1262) );
NAND4_X1 U921 ( .A1(n1267), .A2(n1231), .A3(n1268), .A4(n1269), .ZN(n1204) );
NOR4_X1 U922 ( .A1(n1270), .A2(n1271), .A3(n1272), .A4(n1273), .ZN(n1269) );
NAND4_X1 U923 ( .A1(n1274), .A2(n1137), .A3(n1275), .A4(n1132), .ZN(n1268) );
XNOR2_X1 U924 ( .A(n1126), .B(KEYINPUT25), .ZN(n1274) );
NAND3_X1 U925 ( .A1(n1140), .A2(n1264), .A3(n1135), .ZN(n1231) );
NAND3_X1 U926 ( .A1(n1140), .A2(n1276), .A3(n1277), .ZN(n1267) );
XNOR2_X1 U927 ( .A(KEYINPUT52), .B(n1278), .ZN(n1276) );
AND4_X1 U928 ( .A1(n1279), .A2(n1280), .A3(n1281), .A4(n1282), .ZN(n1193) );
AND4_X1 U929 ( .A1(n1283), .A2(n1284), .A3(n1285), .A4(n1286), .ZN(n1282) );
NAND3_X1 U930 ( .A1(n1287), .A2(n1134), .A3(n1288), .ZN(n1281) );
XNOR2_X1 U931 ( .A(n1289), .B(KEYINPUT16), .ZN(n1288) );
NAND3_X1 U932 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1280) );
XNOR2_X1 U933 ( .A(KEYINPUT26), .B(n1130), .ZN(n1291) );
INV_X1 U934 ( .A(n1293), .ZN(n1290) );
NAND3_X1 U935 ( .A1(n1289), .A2(n1135), .A3(n1287), .ZN(n1279) );
NOR2_X1 U936 ( .A1(n1294), .A2(n1142), .ZN(n1255) );
XNOR2_X1 U937 ( .A(G952), .B(KEYINPUT47), .ZN(n1294) );
XOR2_X1 U938 ( .A(n1295), .B(n1296), .Z(G48) );
NOR2_X1 U939 ( .A1(KEYINPUT35), .A2(n1297), .ZN(n1296) );
NOR4_X1 U940 ( .A1(n1293), .A2(n1298), .A3(n1299), .A4(n1300), .ZN(n1295) );
XNOR2_X1 U941 ( .A(KEYINPUT33), .B(n1301), .ZN(n1300) );
XNOR2_X1 U942 ( .A(KEYINPUT46), .B(n1302), .ZN(n1299) );
XNOR2_X1 U943 ( .A(G143), .B(n1285), .ZN(G45) );
NAND3_X1 U944 ( .A1(n1287), .A2(n1132), .A3(n1303), .ZN(n1285) );
INV_X1 U945 ( .A(n1278), .ZN(n1303) );
XOR2_X1 U946 ( .A(G140), .B(n1304), .Z(G42) );
AND2_X1 U947 ( .A1(n1266), .A2(n1131), .ZN(n1304) );
XOR2_X1 U948 ( .A(n1284), .B(n1305), .Z(G39) );
XNOR2_X1 U949 ( .A(G137), .B(KEYINPUT36), .ZN(n1305) );
NAND3_X1 U950 ( .A1(n1289), .A2(n1306), .A3(n1137), .ZN(n1284) );
XNOR2_X1 U951 ( .A(G134), .B(n1307), .ZN(G36) );
NAND2_X1 U952 ( .A1(n1292), .A2(n1306), .ZN(n1307) );
NAND2_X1 U953 ( .A1(n1308), .A2(n1309), .ZN(G33) );
NAND2_X1 U954 ( .A1(G131), .A2(n1283), .ZN(n1309) );
XOR2_X1 U955 ( .A(KEYINPUT57), .B(n1310), .Z(n1308) );
NOR2_X1 U956 ( .A1(G131), .A2(n1283), .ZN(n1310) );
NAND2_X1 U957 ( .A1(n1266), .A2(n1132), .ZN(n1283) );
AND2_X1 U958 ( .A1(n1135), .A2(n1306), .ZN(n1266) );
NOR2_X1 U959 ( .A1(n1130), .A2(n1293), .ZN(n1306) );
NAND2_X1 U960 ( .A1(n1311), .A2(n1128), .ZN(n1130) );
INV_X1 U961 ( .A(n1127), .ZN(n1311) );
XOR2_X1 U962 ( .A(n1312), .B(n1313), .Z(G30) );
XOR2_X1 U963 ( .A(KEYINPUT19), .B(G128), .Z(n1313) );
NAND3_X1 U964 ( .A1(n1289), .A2(n1134), .A3(n1287), .ZN(n1312) );
NOR2_X1 U965 ( .A1(n1293), .A2(n1302), .ZN(n1287) );
NAND3_X1 U966 ( .A1(n1138), .A2(n1139), .A3(n1314), .ZN(n1293) );
XNOR2_X1 U967 ( .A(G101), .B(n1315), .ZN(G3) );
NAND3_X1 U968 ( .A1(n1264), .A2(n1132), .A3(n1137), .ZN(n1315) );
XOR2_X1 U969 ( .A(n1316), .B(G125), .Z(G27) );
NAND2_X1 U970 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
OR2_X1 U971 ( .A1(n1286), .A2(KEYINPUT7), .ZN(n1318) );
NAND2_X1 U972 ( .A1(n1319), .A2(n1320), .ZN(n1286) );
NAND3_X1 U973 ( .A1(n1320), .A2(n1116), .A3(KEYINPUT7), .ZN(n1317) );
AND4_X1 U974 ( .A1(n1131), .A2(n1135), .A3(n1126), .A4(n1314), .ZN(n1320) );
NAND2_X1 U975 ( .A1(n1112), .A2(n1321), .ZN(n1314) );
NAND4_X1 U976 ( .A1(G902), .A2(G953), .A3(n1322), .A4(n1178), .ZN(n1321) );
INV_X1 U977 ( .A(G900), .ZN(n1178) );
XNOR2_X1 U978 ( .A(G122), .B(n1323), .ZN(G24) );
NAND3_X1 U979 ( .A1(n1324), .A2(n1319), .A3(n1325), .ZN(n1323) );
NOR3_X1 U980 ( .A1(n1278), .A2(n1326), .A3(n1124), .ZN(n1325) );
INV_X1 U981 ( .A(n1140), .ZN(n1124) );
NOR2_X1 U982 ( .A1(n1327), .A2(n1168), .ZN(n1140) );
NAND2_X1 U983 ( .A1(n1328), .A2(n1329), .ZN(n1278) );
INV_X1 U984 ( .A(n1116), .ZN(n1319) );
XNOR2_X1 U985 ( .A(n1126), .B(KEYINPUT43), .ZN(n1324) );
XOR2_X1 U986 ( .A(n1273), .B(n1330), .Z(G21) );
NOR2_X1 U987 ( .A1(KEYINPUT32), .A2(n1331), .ZN(n1330) );
AND3_X1 U988 ( .A1(n1137), .A2(n1289), .A3(n1277), .ZN(n1273) );
INV_X1 U989 ( .A(n1301), .ZN(n1289) );
XNOR2_X1 U990 ( .A(n1332), .B(n1272), .ZN(G18) );
AND2_X1 U991 ( .A1(n1277), .A2(n1292), .ZN(n1272) );
AND2_X1 U992 ( .A1(n1134), .A2(n1132), .ZN(n1292) );
NOR2_X1 U993 ( .A1(n1329), .A2(n1333), .ZN(n1134) );
XNOR2_X1 U994 ( .A(G113), .B(n1334), .ZN(G15) );
NAND2_X1 U995 ( .A1(n1271), .A2(n1335), .ZN(n1334) );
XOR2_X1 U996 ( .A(KEYINPUT37), .B(KEYINPUT13), .Z(n1335) );
AND3_X1 U997 ( .A1(n1135), .A2(n1132), .A3(n1277), .ZN(n1271) );
NOR3_X1 U998 ( .A1(n1302), .A2(n1326), .A3(n1116), .ZN(n1277) );
NAND2_X1 U999 ( .A1(n1336), .A2(n1139), .ZN(n1116) );
INV_X1 U1000 ( .A(n1147), .ZN(n1336) );
XOR2_X1 U1001 ( .A(n1138), .B(KEYINPUT21), .Z(n1147) );
INV_X1 U1002 ( .A(n1337), .ZN(n1326) );
NAND2_X1 U1003 ( .A1(n1338), .A2(n1339), .ZN(n1132) );
OR2_X1 U1004 ( .A1(n1301), .A2(KEYINPUT58), .ZN(n1339) );
NAND2_X1 U1005 ( .A1(n1168), .A2(n1327), .ZN(n1301) );
NAND3_X1 U1006 ( .A1(n1168), .A2(n1167), .A3(KEYINPUT58), .ZN(n1338) );
INV_X1 U1007 ( .A(n1298), .ZN(n1135) );
NAND2_X1 U1008 ( .A1(n1333), .A2(n1329), .ZN(n1298) );
XOR2_X1 U1009 ( .A(n1270), .B(n1340), .Z(G12) );
NOR2_X1 U1010 ( .A1(KEYINPUT49), .A2(n1341), .ZN(n1340) );
AND3_X1 U1011 ( .A1(n1137), .A2(n1264), .A3(n1131), .ZN(n1270) );
NOR2_X1 U1012 ( .A1(n1168), .A2(n1167), .ZN(n1131) );
INV_X1 U1013 ( .A(n1327), .ZN(n1167) );
XOR2_X1 U1014 ( .A(n1342), .B(n1217), .Z(n1327) );
NAND2_X1 U1015 ( .A1(G217), .A2(n1343), .ZN(n1217) );
NAND2_X1 U1016 ( .A1(n1215), .A2(n1344), .ZN(n1342) );
XNOR2_X1 U1017 ( .A(n1345), .B(n1346), .ZN(n1215) );
XNOR2_X1 U1018 ( .A(n1347), .B(n1348), .ZN(n1346) );
NAND3_X1 U1019 ( .A1(n1349), .A2(n1350), .A3(G221), .ZN(n1347) );
XOR2_X1 U1020 ( .A(n1351), .B(n1352), .Z(n1345) );
NOR2_X1 U1021 ( .A1(KEYINPUT23), .A2(n1353), .ZN(n1352) );
XNOR2_X1 U1022 ( .A(G137), .B(G128), .ZN(n1351) );
XOR2_X1 U1023 ( .A(n1354), .B(n1243), .Z(n1168) );
INV_X1 U1024 ( .A(G472), .ZN(n1243) );
NAND3_X1 U1025 ( .A1(n1355), .A2(n1344), .A3(n1356), .ZN(n1354) );
NAND3_X1 U1026 ( .A1(n1241), .A2(n1357), .A3(KEYINPUT8), .ZN(n1356) );
NAND3_X1 U1027 ( .A1(n1358), .A2(n1359), .A3(n1239), .ZN(n1357) );
NAND2_X1 U1028 ( .A1(n1238), .A2(n1360), .ZN(n1359) );
NAND2_X1 U1029 ( .A1(n1361), .A2(KEYINPUT56), .ZN(n1358) );
NAND4_X1 U1030 ( .A1(n1362), .A2(n1240), .A3(n1363), .A4(n1364), .ZN(n1355) );
OR2_X1 U1031 ( .A1(n1239), .A2(n1360), .ZN(n1364) );
INV_X1 U1032 ( .A(KEYINPUT56), .ZN(n1360) );
NAND2_X1 U1033 ( .A1(n1237), .A2(n1238), .ZN(n1239) );
OR2_X1 U1034 ( .A1(n1238), .A2(KEYINPUT56), .ZN(n1363) );
INV_X1 U1035 ( .A(n1361), .ZN(n1240) );
NOR2_X1 U1036 ( .A1(n1238), .A2(n1237), .ZN(n1361) );
XNOR2_X1 U1037 ( .A(n1365), .B(n1366), .ZN(n1237) );
XOR2_X1 U1038 ( .A(G101), .B(n1367), .Z(n1238) );
NOR3_X1 U1039 ( .A1(n1368), .A2(G237), .A3(n1369), .ZN(n1367) );
INV_X1 U1040 ( .A(G210), .ZN(n1369) );
XOR2_X1 U1041 ( .A(KEYINPUT40), .B(n1350), .Z(n1368) );
NAND2_X1 U1042 ( .A1(KEYINPUT8), .A2(n1241), .ZN(n1362) );
AND2_X1 U1043 ( .A1(n1370), .A2(n1371), .ZN(n1241) );
NAND2_X1 U1044 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
XNOR2_X1 U1045 ( .A(n1331), .B(n1374), .ZN(n1372) );
XOR2_X1 U1046 ( .A(n1375), .B(KEYINPUT17), .Z(n1370) );
NAND2_X1 U1047 ( .A1(n1376), .A2(G113), .ZN(n1375) );
XNOR2_X1 U1048 ( .A(G119), .B(n1374), .ZN(n1376) );
NOR2_X1 U1049 ( .A1(KEYINPUT60), .A2(G116), .ZN(n1374) );
AND2_X1 U1050 ( .A1(n1126), .A2(n1275), .ZN(n1264) );
AND3_X1 U1051 ( .A1(n1139), .A2(n1337), .A3(n1138), .ZN(n1275) );
NAND2_X1 U1052 ( .A1(n1377), .A2(n1378), .ZN(n1138) );
INV_X1 U1053 ( .A(n1169), .ZN(n1378) );
NOR2_X1 U1054 ( .A1(n1379), .A2(n1380), .ZN(n1169) );
XNOR2_X1 U1055 ( .A(n1171), .B(KEYINPUT9), .ZN(n1377) );
AND2_X1 U1056 ( .A1(n1380), .A2(n1379), .ZN(n1171) );
NAND2_X1 U1057 ( .A1(n1381), .A2(n1344), .ZN(n1379) );
XOR2_X1 U1058 ( .A(n1382), .B(n1383), .Z(n1381) );
XNOR2_X1 U1059 ( .A(KEYINPUT14), .B(n1252), .ZN(n1383) );
XNOR2_X1 U1060 ( .A(n1245), .B(n1253), .ZN(n1382) );
INV_X1 U1061 ( .A(n1188), .ZN(n1253) );
XNOR2_X1 U1062 ( .A(n1384), .B(G128), .ZN(n1188) );
NAND2_X1 U1063 ( .A1(KEYINPUT34), .A2(n1385), .ZN(n1384) );
XOR2_X1 U1064 ( .A(n1386), .B(n1387), .Z(n1385) );
XOR2_X1 U1065 ( .A(KEYINPUT51), .B(G143), .Z(n1387) );
NOR2_X1 U1066 ( .A1(KEYINPUT38), .A2(n1297), .ZN(n1386) );
XOR2_X1 U1067 ( .A(n1388), .B(n1389), .Z(n1245) );
XNOR2_X1 U1068 ( .A(G140), .B(n1341), .ZN(n1389) );
INV_X1 U1069 ( .A(G110), .ZN(n1341) );
XNOR2_X1 U1070 ( .A(n1390), .B(n1391), .ZN(n1388) );
INV_X1 U1071 ( .A(n1365), .ZN(n1391) );
XNOR2_X1 U1072 ( .A(n1392), .B(n1191), .ZN(n1365) );
XOR2_X1 U1073 ( .A(G134), .B(G137), .Z(n1191) );
XNOR2_X1 U1074 ( .A(G131), .B(KEYINPUT18), .ZN(n1392) );
NAND2_X1 U1075 ( .A1(G227), .A2(n1350), .ZN(n1390) );
XNOR2_X1 U1076 ( .A(n1254), .B(KEYINPUT59), .ZN(n1380) );
INV_X1 U1077 ( .A(G469), .ZN(n1254) );
NAND2_X1 U1078 ( .A1(n1112), .A2(n1393), .ZN(n1337) );
NAND4_X1 U1079 ( .A1(G902), .A2(G953), .A3(n1322), .A4(n1208), .ZN(n1393) );
INV_X1 U1080 ( .A(G898), .ZN(n1208) );
NAND3_X1 U1081 ( .A1(n1322), .A2(n1142), .A3(G952), .ZN(n1112) );
NAND2_X1 U1082 ( .A1(G237), .A2(G234), .ZN(n1322) );
NAND2_X1 U1083 ( .A1(G221), .A2(n1343), .ZN(n1139) );
NAND2_X1 U1084 ( .A1(G234), .A2(n1344), .ZN(n1343) );
INV_X1 U1085 ( .A(n1302), .ZN(n1126) );
NAND2_X1 U1086 ( .A1(n1127), .A2(n1128), .ZN(n1302) );
NAND2_X1 U1087 ( .A1(G214), .A2(n1394), .ZN(n1128) );
XOR2_X1 U1088 ( .A(KEYINPUT55), .B(n1395), .Z(n1394) );
NOR2_X1 U1089 ( .A1(G237), .A2(G902), .ZN(n1395) );
XOR2_X1 U1090 ( .A(n1396), .B(n1157), .Z(n1127) );
NAND2_X1 U1091 ( .A1(G210), .A2(n1397), .ZN(n1157) );
NAND2_X1 U1092 ( .A1(n1398), .A2(n1344), .ZN(n1397) );
XOR2_X1 U1093 ( .A(n1154), .B(KEYINPUT53), .Z(n1396) );
NAND2_X1 U1094 ( .A1(n1399), .A2(n1344), .ZN(n1154) );
INV_X1 U1095 ( .A(G902), .ZN(n1344) );
XOR2_X1 U1096 ( .A(n1259), .B(n1400), .Z(n1399) );
XNOR2_X1 U1097 ( .A(n1401), .B(n1402), .ZN(n1400) );
INV_X1 U1098 ( .A(n1260), .ZN(n1402) );
XNOR2_X1 U1099 ( .A(n1403), .B(n1366), .ZN(n1260) );
XNOR2_X1 U1100 ( .A(n1404), .B(n1405), .ZN(n1366) );
XOR2_X1 U1101 ( .A(G143), .B(n1406), .Z(n1405) );
NOR2_X1 U1102 ( .A1(G128), .A2(KEYINPUT54), .ZN(n1406) );
NAND2_X1 U1103 ( .A1(KEYINPUT30), .A2(n1297), .ZN(n1404) );
NAND2_X1 U1104 ( .A1(G224), .A2(n1350), .ZN(n1403) );
NOR2_X1 U1105 ( .A1(KEYINPUT63), .A2(n1181), .ZN(n1401) );
NAND2_X1 U1106 ( .A1(n1407), .A2(n1408), .ZN(n1259) );
NAND2_X1 U1107 ( .A1(n1210), .A2(n1252), .ZN(n1408) );
INV_X1 U1108 ( .A(n1211), .ZN(n1252) );
XNOR2_X1 U1109 ( .A(n1409), .B(n1410), .ZN(n1210) );
XNOR2_X1 U1110 ( .A(n1411), .B(G119), .ZN(n1410) );
XNOR2_X1 U1111 ( .A(G110), .B(n1412), .ZN(n1409) );
NAND2_X1 U1112 ( .A1(n1413), .A2(n1211), .ZN(n1407) );
XOR2_X1 U1113 ( .A(G101), .B(n1414), .Z(n1211) );
XOR2_X1 U1114 ( .A(G107), .B(G104), .Z(n1414) );
XOR2_X1 U1115 ( .A(n1415), .B(n1412), .Z(n1413) );
XNOR2_X1 U1116 ( .A(n1373), .B(G116), .ZN(n1412) );
INV_X1 U1117 ( .A(G113), .ZN(n1373) );
XNOR2_X1 U1118 ( .A(G122), .B(n1348), .ZN(n1415) );
XNOR2_X1 U1119 ( .A(G110), .B(n1331), .ZN(n1348) );
INV_X1 U1120 ( .A(G119), .ZN(n1331) );
NOR2_X1 U1121 ( .A1(n1328), .A2(n1329), .ZN(n1137) );
NAND2_X1 U1122 ( .A1(n1416), .A2(n1417), .ZN(n1329) );
NAND2_X1 U1123 ( .A1(n1418), .A2(n1226), .ZN(n1417) );
XOR2_X1 U1124 ( .A(KEYINPUT24), .B(n1419), .Z(n1416) );
NOR2_X1 U1125 ( .A1(n1226), .A2(n1418), .ZN(n1419) );
XNOR2_X1 U1126 ( .A(KEYINPUT1), .B(n1165), .ZN(n1418) );
INV_X1 U1127 ( .A(n1222), .ZN(n1165) );
NOR2_X1 U1128 ( .A1(n1227), .A2(G902), .ZN(n1222) );
XNOR2_X1 U1129 ( .A(n1420), .B(n1421), .ZN(n1227) );
XOR2_X1 U1130 ( .A(n1422), .B(n1423), .Z(n1421) );
XNOR2_X1 U1131 ( .A(n1411), .B(G113), .ZN(n1423) );
XOR2_X1 U1132 ( .A(G143), .B(G131), .Z(n1422) );
XNOR2_X1 U1133 ( .A(n1353), .B(n1424), .ZN(n1420) );
XNOR2_X1 U1134 ( .A(G104), .B(n1425), .ZN(n1424) );
NAND4_X1 U1135 ( .A1(KEYINPUT5), .A2(G214), .A3(n1350), .A4(n1398), .ZN(n1425) );
INV_X1 U1136 ( .A(G237), .ZN(n1398) );
XNOR2_X1 U1137 ( .A(n1426), .B(n1427), .ZN(n1353) );
XNOR2_X1 U1138 ( .A(KEYINPUT27), .B(n1297), .ZN(n1427) );
INV_X1 U1139 ( .A(G146), .ZN(n1297) );
XOR2_X1 U1140 ( .A(G140), .B(n1181), .Z(n1426) );
XNOR2_X1 U1141 ( .A(G125), .B(KEYINPUT6), .ZN(n1181) );
INV_X1 U1142 ( .A(G475), .ZN(n1226) );
INV_X1 U1143 ( .A(n1333), .ZN(n1328) );
NOR2_X1 U1144 ( .A1(n1428), .A2(n1170), .ZN(n1333) );
NOR3_X1 U1145 ( .A1(G478), .A2(G902), .A3(n1160), .ZN(n1170) );
AND2_X1 U1146 ( .A1(n1429), .A2(n1430), .ZN(n1428) );
OR2_X1 U1147 ( .A1(n1160), .A2(G902), .ZN(n1430) );
XNOR2_X1 U1148 ( .A(n1431), .B(n1432), .ZN(n1160) );
XOR2_X1 U1149 ( .A(G107), .B(n1433), .Z(n1432) );
XOR2_X1 U1150 ( .A(G134), .B(G128), .Z(n1433) );
XOR2_X1 U1151 ( .A(n1434), .B(n1435), .Z(n1431) );
XOR2_X1 U1152 ( .A(n1436), .B(n1437), .Z(n1435) );
NAND3_X1 U1153 ( .A1(n1438), .A2(n1439), .A3(n1440), .ZN(n1437) );
NAND2_X1 U1154 ( .A1(G116), .A2(n1411), .ZN(n1440) );
INV_X1 U1155 ( .A(G122), .ZN(n1411) );
NAND2_X1 U1156 ( .A1(KEYINPUT42), .A2(n1441), .ZN(n1439) );
NAND2_X1 U1157 ( .A1(G122), .A2(n1442), .ZN(n1441) );
XNOR2_X1 U1158 ( .A(KEYINPUT12), .B(n1332), .ZN(n1442) );
NAND2_X1 U1159 ( .A1(n1443), .A2(n1444), .ZN(n1438) );
INV_X1 U1160 ( .A(KEYINPUT42), .ZN(n1444) );
NAND2_X1 U1161 ( .A1(n1445), .A2(n1446), .ZN(n1443) );
NAND3_X1 U1162 ( .A1(KEYINPUT12), .A2(G122), .A3(n1332), .ZN(n1446) );
OR2_X1 U1163 ( .A1(n1332), .A2(KEYINPUT12), .ZN(n1445) );
INV_X1 U1164 ( .A(G116), .ZN(n1332) );
NAND3_X1 U1165 ( .A1(G217), .A2(n1350), .A3(n1349), .ZN(n1436) );
XNOR2_X1 U1166 ( .A(G234), .B(KEYINPUT45), .ZN(n1349) );
XNOR2_X1 U1167 ( .A(n1142), .B(KEYINPUT11), .ZN(n1350) );
INV_X1 U1168 ( .A(G953), .ZN(n1142) );
NAND2_X1 U1169 ( .A1(KEYINPUT3), .A2(G143), .ZN(n1434) );
XNOR2_X1 U1170 ( .A(KEYINPUT31), .B(n1159), .ZN(n1429) );
INV_X1 U1171 ( .A(G478), .ZN(n1159) );
endmodule


