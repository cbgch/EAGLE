//Key = 1100011110001001001000110111101011011111011111110100101101000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303;

XNOR2_X1 U713 ( .A(G107), .B(n989), .ZN(G9) );
NOR2_X1 U714 ( .A1(n990), .A2(n991), .ZN(G75) );
NOR3_X1 U715 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
NAND3_X1 U716 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n992) );
NAND2_X1 U717 ( .A1(n998), .A2(n999), .ZN(n997) );
NAND2_X1 U718 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NAND4_X1 U719 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n1001) );
NAND2_X1 U720 ( .A1(n1006), .A2(n1007), .ZN(n1000) );
NAND2_X1 U721 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND3_X1 U722 ( .A1(n1010), .A2(n1011), .A3(n1004), .ZN(n1009) );
NAND3_X1 U723 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1010) );
NAND2_X1 U724 ( .A1(n1003), .A2(n1015), .ZN(n1014) );
NAND3_X1 U725 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1013) );
XNOR2_X1 U726 ( .A(n1003), .B(KEYINPUT38), .ZN(n1018) );
NAND2_X1 U727 ( .A1(n1002), .A2(n1019), .ZN(n1012) );
NAND2_X1 U728 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND4_X1 U729 ( .A1(n1002), .A2(n1003), .A3(n1022), .A4(n1023), .ZN(n1008) );
NAND2_X1 U730 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
OR3_X1 U731 ( .A1(n1026), .A2(n1027), .A3(n1024), .ZN(n1022) );
INV_X1 U732 ( .A(n1028), .ZN(n998) );
NOR3_X1 U733 ( .A1(n1029), .A2(G953), .A3(n1030), .ZN(n990) );
INV_X1 U734 ( .A(n995), .ZN(n1030) );
NAND4_X1 U735 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n995) );
NOR4_X1 U736 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1034) );
XNOR2_X1 U737 ( .A(n1039), .B(n1040), .ZN(n1038) );
XNOR2_X1 U738 ( .A(n1041), .B(n1042), .ZN(n1037) );
XNOR2_X1 U739 ( .A(G475), .B(KEYINPUT48), .ZN(n1042) );
XNOR2_X1 U740 ( .A(n1043), .B(n1044), .ZN(n1036) );
XNOR2_X1 U741 ( .A(n1045), .B(KEYINPUT49), .ZN(n1043) );
XOR2_X1 U742 ( .A(n1046), .B(n1047), .Z(n1035) );
NAND2_X1 U743 ( .A1(KEYINPUT15), .A2(n1048), .ZN(n1046) );
NOR3_X1 U744 ( .A1(n1024), .A2(n1049), .A3(n1017), .ZN(n1033) );
NAND2_X1 U745 ( .A1(G472), .A2(n1050), .ZN(n1032) );
XOR2_X1 U746 ( .A(n1051), .B(n1052), .Z(n1031) );
NOR2_X1 U747 ( .A1(G469), .A2(KEYINPUT34), .ZN(n1052) );
XNOR2_X1 U748 ( .A(KEYINPUT24), .B(n993), .ZN(n1029) );
XOR2_X1 U749 ( .A(n1053), .B(n1054), .Z(G72) );
NOR2_X1 U750 ( .A1(KEYINPUT56), .A2(n1055), .ZN(n1054) );
XOR2_X1 U751 ( .A(n1056), .B(n1057), .Z(n1055) );
NAND3_X1 U752 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
INV_X1 U753 ( .A(n1061), .ZN(n1060) );
NAND2_X1 U754 ( .A1(n1062), .A2(n1063), .ZN(n1059) );
NAND2_X1 U755 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
OR2_X1 U756 ( .A1(n1066), .A2(KEYINPUT17), .ZN(n1065) );
NAND2_X1 U757 ( .A1(KEYINPUT17), .A2(n1067), .ZN(n1064) );
NAND2_X1 U758 ( .A1(n1068), .A2(n1066), .ZN(n1058) );
NOR2_X1 U759 ( .A1(KEYINPUT16), .A2(n1069), .ZN(n1066) );
INV_X1 U760 ( .A(n1067), .ZN(n1069) );
XOR2_X1 U761 ( .A(n1070), .B(n1071), .Z(n1067) );
XOR2_X1 U762 ( .A(G128), .B(n1072), .Z(n1071) );
XOR2_X1 U763 ( .A(KEYINPUT29), .B(G131), .Z(n1072) );
XOR2_X1 U764 ( .A(n1073), .B(n1074), .Z(n1070) );
INV_X1 U765 ( .A(n1063), .ZN(n1068) );
NAND2_X1 U766 ( .A1(n1075), .A2(n996), .ZN(n1056) );
NAND2_X1 U767 ( .A1(G953), .A2(n1076), .ZN(n1053) );
NAND2_X1 U768 ( .A1(G900), .A2(G227), .ZN(n1076) );
XOR2_X1 U769 ( .A(n1077), .B(n1078), .Z(G69) );
XOR2_X1 U770 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U771 ( .A1(n1081), .A2(n996), .ZN(n1080) );
AND2_X1 U772 ( .A1(G224), .A2(G898), .ZN(n1081) );
NAND2_X1 U773 ( .A1(n1082), .A2(n1083), .ZN(n1079) );
NAND2_X1 U774 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XOR2_X1 U775 ( .A(n1086), .B(n1087), .Z(n1082) );
XNOR2_X1 U776 ( .A(n1088), .B(n1089), .ZN(n1087) );
XOR2_X1 U777 ( .A(KEYINPUT50), .B(KEYINPUT4), .Z(n1086) );
NAND2_X1 U778 ( .A1(n996), .A2(n1090), .ZN(n1077) );
NOR2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(G66) );
NOR3_X1 U780 ( .A1(n1045), .A2(n1093), .A3(n1094), .ZN(n1092) );
NOR3_X1 U781 ( .A1(n1095), .A2(n1044), .A3(n1096), .ZN(n1094) );
INV_X1 U782 ( .A(n1097), .ZN(n1095) );
NOR2_X1 U783 ( .A1(n1098), .A2(n1097), .ZN(n1093) );
NOR2_X1 U784 ( .A1(n1099), .A2(n1044), .ZN(n1098) );
NOR2_X1 U785 ( .A1(n1091), .A2(n1100), .ZN(G63) );
NOR3_X1 U786 ( .A1(n1047), .A2(n1101), .A3(n1102), .ZN(n1100) );
NOR3_X1 U787 ( .A1(n1103), .A2(n1048), .A3(n1096), .ZN(n1102) );
INV_X1 U788 ( .A(n1104), .ZN(n1096) );
NOR2_X1 U789 ( .A1(n1105), .A2(n1106), .ZN(n1101) );
NOR2_X1 U790 ( .A1(n1099), .A2(n1048), .ZN(n1106) );
NOR2_X1 U791 ( .A1(n1091), .A2(n1107), .ZN(G60) );
NOR3_X1 U792 ( .A1(n1041), .A2(n1108), .A3(n1109), .ZN(n1107) );
AND3_X1 U793 ( .A1(n1110), .A2(G475), .A3(n1104), .ZN(n1109) );
NOR2_X1 U794 ( .A1(n1111), .A2(n1110), .ZN(n1108) );
AND2_X1 U795 ( .A1(n994), .A2(G475), .ZN(n1111) );
INV_X1 U796 ( .A(n1099), .ZN(n994) );
XNOR2_X1 U797 ( .A(G104), .B(n1112), .ZN(G6) );
NOR3_X1 U798 ( .A1(n1091), .A2(n1113), .A3(n1114), .ZN(G57) );
NOR3_X1 U799 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
NOR2_X1 U800 ( .A1(KEYINPUT21), .A2(n1118), .ZN(n1116) );
INV_X1 U801 ( .A(KEYINPUT19), .ZN(n1118) );
INV_X1 U802 ( .A(n1119), .ZN(n1115) );
NOR2_X1 U803 ( .A1(n1120), .A2(n1119), .ZN(n1113) );
NAND3_X1 U804 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1119) );
NAND2_X1 U805 ( .A1(KEYINPUT58), .A2(n1124), .ZN(n1123) );
NAND2_X1 U806 ( .A1(n1125), .A2(n1126), .ZN(n1122) );
NAND3_X1 U807 ( .A1(G472), .A2(n1127), .A3(n1104), .ZN(n1126) );
INV_X1 U808 ( .A(KEYINPUT40), .ZN(n1127) );
OR4_X1 U809 ( .A1(KEYINPUT40), .A2(KEYINPUT58), .A3(n1124), .A4(n1125), .ZN(n1121) );
XOR2_X1 U810 ( .A(n1128), .B(n1129), .Z(n1125) );
NAND2_X1 U811 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
NAND2_X1 U812 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
INV_X1 U813 ( .A(KEYINPUT3), .ZN(n1133) );
NAND3_X1 U814 ( .A1(n1134), .A2(n1135), .A3(KEYINPUT3), .ZN(n1130) );
NAND2_X1 U815 ( .A1(n1104), .A2(G472), .ZN(n1124) );
NOR2_X1 U816 ( .A1(KEYINPUT19), .A2(n1136), .ZN(n1120) );
XNOR2_X1 U817 ( .A(n1137), .B(KEYINPUT21), .ZN(n1136) );
NOR2_X1 U818 ( .A1(n1091), .A2(n1138), .ZN(G54) );
XOR2_X1 U819 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U820 ( .A(KEYINPUT46), .B(n1141), .Z(n1140) );
AND2_X1 U821 ( .A1(G469), .A2(n1104), .ZN(n1141) );
NOR2_X1 U822 ( .A1(n1091), .A2(n1142), .ZN(G51) );
XOR2_X1 U823 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR3_X1 U824 ( .A1(KEYINPUT51), .A2(n1145), .A3(n1146), .ZN(n1144) );
NOR2_X1 U825 ( .A1(n1135), .A2(n1147), .ZN(n1146) );
XOR2_X1 U826 ( .A(KEYINPUT44), .B(n1148), .Z(n1147) );
NOR2_X1 U827 ( .A1(n1149), .A2(n1148), .ZN(n1145) );
INV_X1 U828 ( .A(n1135), .ZN(n1149) );
NAND2_X1 U829 ( .A1(n1104), .A2(n1039), .ZN(n1143) );
NOR2_X1 U830 ( .A1(n1150), .A2(n1099), .ZN(n1104) );
NOR2_X1 U831 ( .A1(n1090), .A2(n1075), .ZN(n1099) );
NAND4_X1 U832 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1075) );
NOR4_X1 U833 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1154) );
OR2_X1 U834 ( .A1(n1159), .A2(n1160), .ZN(n1153) );
NAND3_X1 U835 ( .A1(n1026), .A2(n1161), .A3(n1162), .ZN(n1152) );
NAND2_X1 U836 ( .A1(n1163), .A2(n1164), .ZN(n1151) );
NAND2_X1 U837 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NAND2_X1 U838 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND2_X1 U839 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND3_X1 U840 ( .A1(n1171), .A2(n1159), .A3(n1002), .ZN(n1170) );
INV_X1 U841 ( .A(KEYINPUT35), .ZN(n1159) );
NAND2_X1 U842 ( .A1(n1172), .A2(n1015), .ZN(n1169) );
NAND2_X1 U843 ( .A1(n1162), .A2(n1027), .ZN(n1165) );
NAND4_X1 U844 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1090) );
AND4_X1 U845 ( .A1(n989), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1176) );
NAND3_X1 U846 ( .A1(n1161), .A2(n1180), .A3(n1004), .ZN(n989) );
NOR3_X1 U847 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1175) );
NOR2_X1 U848 ( .A1(n1184), .A2(n1112), .ZN(n1183) );
NAND3_X1 U849 ( .A1(n1004), .A2(n1180), .A3(n1163), .ZN(n1112) );
INV_X1 U850 ( .A(KEYINPUT43), .ZN(n1184) );
NOR4_X1 U851 ( .A1(KEYINPUT43), .A2(n1185), .A3(n1025), .A4(n1020), .ZN(n1182) );
INV_X1 U852 ( .A(n1004), .ZN(n1025) );
NAND3_X1 U853 ( .A1(n1186), .A2(n1187), .A3(n1015), .ZN(n1185) );
INV_X1 U854 ( .A(n1005), .ZN(n1186) );
INV_X1 U855 ( .A(n1188), .ZN(n1181) );
AND2_X1 U856 ( .A1(G953), .A2(n1189), .ZN(n1091) );
XNOR2_X1 U857 ( .A(KEYINPUT41), .B(n993), .ZN(n1189) );
INV_X1 U858 ( .A(G952), .ZN(n993) );
XNOR2_X1 U859 ( .A(G146), .B(n1190), .ZN(G48) );
NAND4_X1 U860 ( .A1(KEYINPUT45), .A2(n1167), .A3(n1191), .A4(n1172), .ZN(n1190) );
NOR2_X1 U861 ( .A1(n1192), .A2(n1020), .ZN(n1191) );
INV_X1 U862 ( .A(n1163), .ZN(n1020) );
XNOR2_X1 U863 ( .A(n1015), .B(KEYINPUT31), .ZN(n1192) );
XOR2_X1 U864 ( .A(G143), .B(n1158), .Z(G45) );
AND4_X1 U865 ( .A1(n1167), .A2(n1026), .A3(n1193), .A4(n1194), .ZN(n1158) );
AND2_X1 U866 ( .A1(n1195), .A2(n1015), .ZN(n1193) );
XNOR2_X1 U867 ( .A(G140), .B(n1196), .ZN(G42) );
NAND4_X1 U868 ( .A1(KEYINPUT12), .A2(n1162), .A3(n1163), .A4(n1027), .ZN(n1196) );
XOR2_X1 U869 ( .A(n1197), .B(n1157), .Z(G39) );
AND3_X1 U870 ( .A1(n1172), .A2(n1003), .A3(n1162), .ZN(n1157) );
NAND2_X1 U871 ( .A1(KEYINPUT6), .A2(n1198), .ZN(n1197) );
INV_X1 U872 ( .A(G137), .ZN(n1198) );
XOR2_X1 U873 ( .A(G134), .B(n1199), .Z(G36) );
NOR3_X1 U874 ( .A1(n1200), .A2(n1021), .A3(n1201), .ZN(n1199) );
XOR2_X1 U875 ( .A(KEYINPUT62), .B(n1026), .Z(n1200) );
XOR2_X1 U876 ( .A(G131), .B(n1156), .Z(G33) );
AND3_X1 U877 ( .A1(n1163), .A2(n1026), .A3(n1162), .ZN(n1156) );
INV_X1 U878 ( .A(n1201), .ZN(n1162) );
NAND4_X1 U879 ( .A1(n1006), .A2(n1015), .A3(n1202), .A4(n1011), .ZN(n1201) );
XNOR2_X1 U880 ( .A(n1155), .B(n1203), .ZN(G30) );
NAND2_X1 U881 ( .A1(KEYINPUT47), .A2(G128), .ZN(n1203) );
AND4_X1 U882 ( .A1(n1167), .A2(n1172), .A3(n1161), .A4(n1015), .ZN(n1155) );
XNOR2_X1 U883 ( .A(G101), .B(n1188), .ZN(G3) );
NAND3_X1 U884 ( .A1(n1003), .A2(n1180), .A3(n1026), .ZN(n1188) );
XOR2_X1 U885 ( .A(n1160), .B(n1204), .Z(G27) );
NAND2_X1 U886 ( .A1(KEYINPUT57), .A2(G125), .ZN(n1204) );
NAND4_X1 U887 ( .A1(n1167), .A2(n1163), .A3(n1002), .A4(n1027), .ZN(n1160) );
AND2_X1 U888 ( .A1(n1005), .A2(n1202), .ZN(n1167) );
NAND2_X1 U889 ( .A1(n1028), .A2(n1205), .ZN(n1202) );
NAND3_X1 U890 ( .A1(G902), .A2(n1206), .A3(n1061), .ZN(n1205) );
NOR2_X1 U891 ( .A1(n1207), .A2(G900), .ZN(n1061) );
INV_X1 U892 ( .A(n1084), .ZN(n1207) );
XNOR2_X1 U893 ( .A(G122), .B(n1173), .ZN(G24) );
NAND4_X1 U894 ( .A1(n1194), .A2(n1208), .A3(n1004), .A4(n1195), .ZN(n1173) );
NOR2_X1 U895 ( .A1(n1209), .A2(n1210), .ZN(n1004) );
XNOR2_X1 U896 ( .A(G119), .B(n1174), .ZN(G21) );
NAND3_X1 U897 ( .A1(n1208), .A2(n1003), .A3(n1172), .ZN(n1174) );
AND2_X1 U898 ( .A1(n1210), .A2(n1209), .ZN(n1172) );
INV_X1 U899 ( .A(n1211), .ZN(n1209) );
XOR2_X1 U900 ( .A(n1179), .B(n1212), .Z(G18) );
NAND2_X1 U901 ( .A1(n1213), .A2(KEYINPUT32), .ZN(n1212) );
XNOR2_X1 U902 ( .A(G116), .B(KEYINPUT1), .ZN(n1213) );
NAND3_X1 U903 ( .A1(n1026), .A2(n1161), .A3(n1208), .ZN(n1179) );
INV_X1 U904 ( .A(n1021), .ZN(n1161) );
NAND2_X1 U905 ( .A1(n1214), .A2(n1215), .ZN(n1021) );
XNOR2_X1 U906 ( .A(n1195), .B(KEYINPUT25), .ZN(n1214) );
XNOR2_X1 U907 ( .A(G113), .B(n1178), .ZN(G15) );
NAND3_X1 U908 ( .A1(n1163), .A2(n1026), .A3(n1208), .ZN(n1178) );
AND3_X1 U909 ( .A1(n1005), .A2(n1187), .A3(n1002), .ZN(n1208) );
NOR2_X1 U910 ( .A1(n1216), .A2(n1217), .ZN(n1002) );
INV_X1 U911 ( .A(n1016), .ZN(n1216) );
NOR2_X1 U912 ( .A1(n1210), .A2(n1211), .ZN(n1026) );
NOR2_X1 U913 ( .A1(n1215), .A2(n1195), .ZN(n1163) );
XNOR2_X1 U914 ( .A(G110), .B(n1177), .ZN(G12) );
NAND3_X1 U915 ( .A1(n1027), .A2(n1180), .A3(n1003), .ZN(n1177) );
NOR2_X1 U916 ( .A1(n1195), .A2(n1194), .ZN(n1003) );
INV_X1 U917 ( .A(n1215), .ZN(n1194) );
XOR2_X1 U918 ( .A(n1041), .B(n1218), .Z(n1215) );
NOR2_X1 U919 ( .A1(G475), .A2(KEYINPUT59), .ZN(n1218) );
NOR2_X1 U920 ( .A1(n1110), .A2(G902), .ZN(n1041) );
XOR2_X1 U921 ( .A(n1219), .B(n1220), .Z(n1110) );
XOR2_X1 U922 ( .A(n1221), .B(n1222), .Z(n1220) );
XOR2_X1 U923 ( .A(G113), .B(G104), .Z(n1222) );
XOR2_X1 U924 ( .A(G131), .B(G122), .Z(n1221) );
XNOR2_X1 U925 ( .A(n1223), .B(n1063), .ZN(n1219) );
XOR2_X1 U926 ( .A(n1224), .B(n1225), .Z(n1223) );
NAND2_X1 U927 ( .A1(G214), .A2(n1226), .ZN(n1224) );
XNOR2_X1 U928 ( .A(n1047), .B(n1048), .ZN(n1195) );
INV_X1 U929 ( .A(G478), .ZN(n1048) );
NOR2_X1 U930 ( .A1(n1105), .A2(G902), .ZN(n1047) );
INV_X1 U931 ( .A(n1103), .ZN(n1105) );
NAND2_X1 U932 ( .A1(n1227), .A2(n1228), .ZN(n1103) );
NAND4_X1 U933 ( .A1(n1229), .A2(G217), .A3(n1230), .A4(G234), .ZN(n1228) );
AND2_X1 U934 ( .A1(n996), .A2(n1231), .ZN(n1230) );
NAND2_X1 U935 ( .A1(n1232), .A2(n1233), .ZN(n1227) );
NAND3_X1 U936 ( .A1(G234), .A2(n996), .A3(G217), .ZN(n1233) );
NAND2_X1 U937 ( .A1(n1229), .A2(n1231), .ZN(n1232) );
NAND2_X1 U938 ( .A1(n1234), .A2(n1235), .ZN(n1231) );
XOR2_X1 U939 ( .A(KEYINPUT13), .B(n1236), .Z(n1235) );
XOR2_X1 U940 ( .A(n1237), .B(KEYINPUT53), .Z(n1229) );
OR2_X1 U941 ( .A1(n1236), .A2(n1234), .ZN(n1237) );
XNOR2_X1 U942 ( .A(G107), .B(n1238), .ZN(n1234) );
XOR2_X1 U943 ( .A(G122), .B(G116), .Z(n1238) );
XNOR2_X1 U944 ( .A(n1239), .B(n1240), .ZN(n1236) );
XNOR2_X1 U945 ( .A(G134), .B(KEYINPUT10), .ZN(n1239) );
AND3_X1 U946 ( .A1(n1005), .A2(n1187), .A3(n1015), .ZN(n1180) );
NOR2_X1 U947 ( .A1(n1016), .A2(n1217), .ZN(n1015) );
XNOR2_X1 U948 ( .A(n1017), .B(KEYINPUT30), .ZN(n1217) );
AND2_X1 U949 ( .A1(G221), .A2(n1241), .ZN(n1017) );
XOR2_X1 U950 ( .A(n1242), .B(G469), .Z(n1016) );
NAND2_X1 U951 ( .A1(KEYINPUT18), .A2(n1051), .ZN(n1242) );
AND2_X1 U952 ( .A1(n1243), .A2(n1150), .ZN(n1051) );
XOR2_X1 U953 ( .A(n1139), .B(KEYINPUT2), .Z(n1243) );
XOR2_X1 U954 ( .A(n1244), .B(n1245), .Z(n1139) );
XOR2_X1 U955 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U956 ( .A(n1248), .B(n1249), .Z(n1247) );
NAND2_X1 U957 ( .A1(n1250), .A2(n1251), .ZN(n1248) );
NAND2_X1 U958 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
XNOR2_X1 U959 ( .A(n1254), .B(KEYINPUT54), .ZN(n1252) );
NAND2_X1 U960 ( .A1(n1255), .A2(G101), .ZN(n1250) );
XOR2_X1 U961 ( .A(KEYINPUT28), .B(n1254), .Z(n1255) );
XNOR2_X1 U962 ( .A(n1134), .B(n1256), .ZN(n1246) );
AND2_X1 U963 ( .A1(n996), .A2(G227), .ZN(n1256) );
XOR2_X1 U964 ( .A(n1257), .B(n1258), .Z(n1244) );
XOR2_X1 U965 ( .A(KEYINPUT60), .B(KEYINPUT14), .Z(n1258) );
XOR2_X1 U966 ( .A(n1073), .B(G140), .Z(n1257) );
NAND2_X1 U967 ( .A1(KEYINPUT7), .A2(n1225), .ZN(n1073) );
XOR2_X1 U968 ( .A(G143), .B(G146), .Z(n1225) );
NAND2_X1 U969 ( .A1(n1259), .A2(n1028), .ZN(n1187) );
NAND3_X1 U970 ( .A1(n1206), .A2(n996), .A3(G952), .ZN(n1028) );
XOR2_X1 U971 ( .A(KEYINPUT23), .B(n1260), .Z(n1259) );
AND4_X1 U972 ( .A1(n1085), .A2(n1206), .A3(G902), .A4(n1084), .ZN(n1260) );
XNOR2_X1 U973 ( .A(G953), .B(KEYINPUT33), .ZN(n1084) );
NAND2_X1 U974 ( .A1(G237), .A2(G234), .ZN(n1206) );
INV_X1 U975 ( .A(G898), .ZN(n1085) );
NOR2_X1 U976 ( .A1(n1006), .A2(n1024), .ZN(n1005) );
INV_X1 U977 ( .A(n1011), .ZN(n1024) );
NAND2_X1 U978 ( .A1(G214), .A2(n1261), .ZN(n1011) );
AND3_X1 U979 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1006) );
NAND2_X1 U980 ( .A1(n1265), .A2(n1040), .ZN(n1264) );
NAND2_X1 U981 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
INV_X1 U982 ( .A(KEYINPUT11), .ZN(n1267) );
XNOR2_X1 U983 ( .A(KEYINPUT36), .B(n1268), .ZN(n1266) );
OR3_X1 U984 ( .A1(n1040), .A2(n1039), .A3(KEYINPUT11), .ZN(n1263) );
NAND2_X1 U985 ( .A1(n1269), .A2(n1150), .ZN(n1040) );
XNOR2_X1 U986 ( .A(n1148), .B(n1270), .ZN(n1269) );
XNOR2_X1 U987 ( .A(n1135), .B(KEYINPUT52), .ZN(n1270) );
XNOR2_X1 U988 ( .A(n1271), .B(n1272), .ZN(n1148) );
XNOR2_X1 U989 ( .A(G125), .B(n1273), .ZN(n1272) );
XNOR2_X1 U990 ( .A(KEYINPUT61), .B(KEYINPUT20), .ZN(n1273) );
XOR2_X1 U991 ( .A(n1088), .B(n1274), .Z(n1271) );
XOR2_X1 U992 ( .A(n1275), .B(n1276), .Z(n1274) );
NAND2_X1 U993 ( .A1(KEYINPUT0), .A2(n1089), .ZN(n1276) );
XOR2_X1 U994 ( .A(G110), .B(n1277), .Z(n1089) );
XOR2_X1 U995 ( .A(KEYINPUT26), .B(G122), .Z(n1277) );
NAND2_X1 U996 ( .A1(G224), .A2(n996), .ZN(n1275) );
XOR2_X1 U997 ( .A(n1278), .B(n1279), .Z(n1088) );
XOR2_X1 U998 ( .A(KEYINPUT5), .B(n1280), .Z(n1279) );
XOR2_X1 U999 ( .A(KEYINPUT9), .B(KEYINPUT63), .Z(n1280) );
XNOR2_X1 U1000 ( .A(n1281), .B(n1129), .ZN(n1278) );
XNOR2_X1 U1001 ( .A(G101), .B(n1254), .ZN(n1281) );
XOR2_X1 U1002 ( .A(G104), .B(G107), .Z(n1254) );
NAND2_X1 U1003 ( .A1(KEYINPUT11), .A2(n1039), .ZN(n1262) );
INV_X1 U1004 ( .A(n1268), .ZN(n1039) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1261), .ZN(n1268) );
NAND2_X1 U1006 ( .A1(n1282), .A2(n1150), .ZN(n1261) );
INV_X1 U1007 ( .A(G237), .ZN(n1282) );
INV_X1 U1008 ( .A(n1171), .ZN(n1027) );
NAND2_X1 U1009 ( .A1(n1211), .A2(n1210), .ZN(n1171) );
XOR2_X1 U1010 ( .A(n1283), .B(n1044), .Z(n1210) );
NAND2_X1 U1011 ( .A1(G217), .A2(n1241), .ZN(n1044) );
NAND2_X1 U1012 ( .A1(G234), .A2(n1150), .ZN(n1241) );
NAND2_X1 U1013 ( .A1(KEYINPUT55), .A2(n1045), .ZN(n1283) );
NOR2_X1 U1014 ( .A1(n1097), .A2(G902), .ZN(n1045) );
XNOR2_X1 U1015 ( .A(n1284), .B(n1285), .ZN(n1097) );
XOR2_X1 U1016 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U1017 ( .A(G137), .B(G146), .ZN(n1287) );
NAND2_X1 U1018 ( .A1(KEYINPUT37), .A2(n1288), .ZN(n1286) );
XNOR2_X1 U1019 ( .A(n1289), .B(n1063), .ZN(n1284) );
XNOR2_X1 U1020 ( .A(G125), .B(G140), .ZN(n1063) );
XOR2_X1 U1021 ( .A(n1290), .B(n1249), .Z(n1289) );
XNOR2_X1 U1022 ( .A(n1291), .B(G128), .ZN(n1249) );
INV_X1 U1023 ( .A(G110), .ZN(n1291) );
NAND3_X1 U1024 ( .A1(G234), .A2(n996), .A3(G221), .ZN(n1290) );
INV_X1 U1025 ( .A(G953), .ZN(n996) );
NOR2_X1 U1026 ( .A1(n1292), .A2(n1049), .ZN(n1211) );
NOR2_X1 U1027 ( .A1(n1050), .A2(G472), .ZN(n1049) );
AND2_X1 U1028 ( .A1(n1293), .A2(n1050), .ZN(n1292) );
NAND2_X1 U1029 ( .A1(n1294), .A2(n1150), .ZN(n1050) );
INV_X1 U1030 ( .A(G902), .ZN(n1150) );
XNOR2_X1 U1031 ( .A(n1295), .B(n1132), .ZN(n1294) );
XOR2_X1 U1032 ( .A(n1135), .B(n1134), .Z(n1132) );
XNOR2_X1 U1033 ( .A(n1296), .B(G131), .ZN(n1134) );
NAND2_X1 U1034 ( .A1(KEYINPUT27), .A2(n1074), .ZN(n1296) );
XOR2_X1 U1035 ( .A(G134), .B(G137), .Z(n1074) );
XOR2_X1 U1036 ( .A(G146), .B(n1240), .Z(n1135) );
XOR2_X1 U1037 ( .A(G143), .B(G128), .Z(n1240) );
NAND2_X1 U1038 ( .A1(n1297), .A2(n1298), .ZN(n1295) );
NAND2_X1 U1039 ( .A1(n1299), .A2(n1129), .ZN(n1298) );
INV_X1 U1040 ( .A(n1300), .ZN(n1129) );
XNOR2_X1 U1041 ( .A(n1137), .B(KEYINPUT22), .ZN(n1299) );
NAND2_X1 U1042 ( .A1(n1301), .A2(n1300), .ZN(n1297) );
XNOR2_X1 U1043 ( .A(n1302), .B(n1288), .ZN(n1300) );
XOR2_X1 U1044 ( .A(G119), .B(KEYINPUT42), .Z(n1288) );
XNOR2_X1 U1045 ( .A(G113), .B(G116), .ZN(n1302) );
XNOR2_X1 U1046 ( .A(KEYINPUT39), .B(n1117), .ZN(n1301) );
INV_X1 U1047 ( .A(n1137), .ZN(n1117) );
XOR2_X1 U1048 ( .A(n1303), .B(n1253), .Z(n1137) );
INV_X1 U1049 ( .A(G101), .ZN(n1253) );
NAND2_X1 U1050 ( .A1(G210), .A2(n1226), .ZN(n1303) );
NOR2_X1 U1051 ( .A1(G953), .A2(G237), .ZN(n1226) );
XNOR2_X1 U1052 ( .A(G472), .B(KEYINPUT8), .ZN(n1293) );
endmodule


