//Key = 0101110100111101010110010010100001111111100001000010001010011101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361;

XNOR2_X1 U745 ( .A(G107), .B(n1042), .ZN(G9) );
NOR2_X1 U746 ( .A1(n1043), .A2(n1044), .ZN(G75) );
NOR3_X1 U747 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NOR2_X1 U748 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U749 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
XOR2_X1 U750 ( .A(n1052), .B(KEYINPUT39), .Z(n1051) );
NAND4_X1 U751 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
AND4_X1 U752 ( .A1(n1056), .A2(n1054), .A3(n1057), .A4(n1053), .ZN(n1050) );
NAND3_X1 U753 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1045) );
NAND3_X1 U754 ( .A1(n1061), .A2(n1062), .A3(n1053), .ZN(n1060) );
INV_X1 U755 ( .A(n1063), .ZN(n1053) );
NAND2_X1 U756 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND2_X1 U757 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U758 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND3_X1 U759 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
XNOR2_X1 U760 ( .A(KEYINPUT49), .B(n1073), .ZN(n1071) );
NAND2_X1 U761 ( .A1(n1074), .A2(n1056), .ZN(n1068) );
NAND2_X1 U762 ( .A1(n1054), .A2(n1075), .ZN(n1064) );
NAND3_X1 U763 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NAND2_X1 U764 ( .A1(n1066), .A2(n1079), .ZN(n1078) );
NAND2_X1 U765 ( .A1(n1056), .A2(n1080), .ZN(n1077) );
NAND2_X1 U766 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U767 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U768 ( .A1(n1085), .A2(n1086), .ZN(n1076) );
XNOR2_X1 U769 ( .A(n1066), .B(KEYINPUT34), .ZN(n1085) );
NOR3_X1 U770 ( .A1(n1087), .A2(G953), .A3(G952), .ZN(n1043) );
INV_X1 U771 ( .A(n1058), .ZN(n1087) );
NAND4_X1 U772 ( .A1(n1088), .A2(n1054), .A3(n1089), .A4(n1090), .ZN(n1058) );
NOR4_X1 U773 ( .A1(n1083), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1090) );
XNOR2_X1 U774 ( .A(n1094), .B(n1095), .ZN(n1091) );
NAND2_X1 U775 ( .A1(KEYINPUT63), .A2(n1096), .ZN(n1094) );
XOR2_X1 U776 ( .A(n1097), .B(n1098), .Z(n1089) );
NOR2_X1 U777 ( .A1(KEYINPUT47), .A2(n1099), .ZN(n1098) );
XOR2_X1 U778 ( .A(n1100), .B(n1101), .Z(G72) );
NOR2_X1 U779 ( .A1(n1102), .A2(n1059), .ZN(n1101) );
AND2_X1 U780 ( .A1(G227), .A2(G900), .ZN(n1102) );
NAND2_X1 U781 ( .A1(n1103), .A2(n1104), .ZN(n1100) );
NAND3_X1 U782 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1104) );
INV_X1 U783 ( .A(n1108), .ZN(n1106) );
OR2_X1 U784 ( .A1(n1105), .A2(n1107), .ZN(n1103) );
XOR2_X1 U785 ( .A(n1109), .B(n1110), .Z(n1107) );
XOR2_X1 U786 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U787 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U788 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XNOR2_X1 U789 ( .A(n1117), .B(KEYINPUT13), .ZN(n1116) );
NOR2_X1 U790 ( .A1(G134), .A2(n1118), .ZN(n1113) );
XOR2_X1 U791 ( .A(KEYINPUT1), .B(n1117), .Z(n1118) );
NOR2_X1 U792 ( .A1(G131), .A2(KEYINPUT51), .ZN(n1111) );
XOR2_X1 U793 ( .A(n1119), .B(G137), .Z(n1109) );
NAND2_X1 U794 ( .A1(n1120), .A2(KEYINPUT61), .ZN(n1119) );
XNOR2_X1 U795 ( .A(n1121), .B(KEYINPUT54), .ZN(n1120) );
NAND2_X1 U796 ( .A1(n1059), .A2(n1122), .ZN(n1105) );
NAND2_X1 U797 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U798 ( .A(n1125), .B(n1126), .Z(G69) );
NAND2_X1 U799 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U800 ( .A1(n1129), .A2(n1059), .ZN(n1128) );
XNOR2_X1 U801 ( .A(n1130), .B(n1131), .ZN(n1129) );
NAND3_X1 U802 ( .A1(n1131), .A2(G898), .A3(G953), .ZN(n1127) );
NOR2_X1 U803 ( .A1(KEYINPUT18), .A2(n1132), .ZN(n1131) );
XOR2_X1 U804 ( .A(n1133), .B(n1134), .Z(n1132) );
XNOR2_X1 U805 ( .A(n1135), .B(n1136), .ZN(n1134) );
XOR2_X1 U806 ( .A(n1137), .B(n1138), .Z(n1133) );
XOR2_X1 U807 ( .A(KEYINPUT27), .B(G110), .Z(n1138) );
NAND2_X1 U808 ( .A1(KEYINPUT17), .A2(n1139), .ZN(n1125) );
NAND2_X1 U809 ( .A1(G953), .A2(n1140), .ZN(n1139) );
NAND2_X1 U810 ( .A1(G898), .A2(G224), .ZN(n1140) );
NOR2_X1 U811 ( .A1(n1141), .A2(n1142), .ZN(G66) );
NOR2_X1 U812 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U813 ( .A(n1145), .B(KEYINPUT5), .Z(n1144) );
NAND2_X1 U814 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
OR3_X1 U815 ( .A1(n1148), .A2(KEYINPUT42), .A3(n1149), .ZN(n1147) );
NOR4_X1 U816 ( .A1(KEYINPUT42), .A2(n1148), .A3(n1149), .A4(n1146), .ZN(n1143) );
NOR2_X1 U817 ( .A1(n1141), .A2(n1150), .ZN(G63) );
XOR2_X1 U818 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U819 ( .A1(n1153), .A2(G478), .ZN(n1151) );
NOR2_X1 U820 ( .A1(n1141), .A2(n1154), .ZN(G60) );
XOR2_X1 U821 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND2_X1 U822 ( .A1(n1153), .A2(G475), .ZN(n1155) );
XNOR2_X1 U823 ( .A(G104), .B(n1157), .ZN(G6) );
NAND2_X1 U824 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U825 ( .A1(KEYINPUT26), .A2(n1160), .ZN(n1159) );
NAND2_X1 U826 ( .A1(KEYINPUT8), .A2(n1161), .ZN(n1158) );
NOR2_X1 U827 ( .A1(n1141), .A2(n1162), .ZN(G57) );
XOR2_X1 U828 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U829 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U830 ( .A(n1167), .B(n1168), .Z(n1163) );
XNOR2_X1 U831 ( .A(G101), .B(n1169), .ZN(n1168) );
NAND2_X1 U832 ( .A1(n1153), .A2(G472), .ZN(n1169) );
NAND2_X1 U833 ( .A1(KEYINPUT50), .A2(n1170), .ZN(n1167) );
NOR2_X1 U834 ( .A1(n1171), .A2(n1172), .ZN(G54) );
XOR2_X1 U835 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U836 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U837 ( .A(n1177), .B(n1178), .ZN(n1176) );
NOR2_X1 U838 ( .A1(KEYINPUT53), .A2(n1179), .ZN(n1178) );
NOR2_X1 U839 ( .A1(KEYINPUT6), .A2(n1180), .ZN(n1177) );
XNOR2_X1 U840 ( .A(n1181), .B(n1182), .ZN(n1180) );
XOR2_X1 U841 ( .A(KEYINPUT19), .B(n1183), .Z(n1182) );
XNOR2_X1 U842 ( .A(n1184), .B(n1185), .ZN(n1173) );
NAND2_X1 U843 ( .A1(n1153), .A2(G469), .ZN(n1184) );
NOR2_X1 U844 ( .A1(n1186), .A2(n1059), .ZN(n1171) );
XNOR2_X1 U845 ( .A(G952), .B(KEYINPUT12), .ZN(n1186) );
NOR3_X1 U846 ( .A1(n1141), .A2(n1187), .A3(n1188), .ZN(G51) );
NOR2_X1 U847 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U848 ( .A(n1191), .B(n1192), .Z(n1190) );
AND2_X1 U849 ( .A1(n1193), .A2(KEYINPUT15), .ZN(n1192) );
INV_X1 U850 ( .A(KEYINPUT23), .ZN(n1189) );
NOR2_X1 U851 ( .A1(KEYINPUT23), .A2(n1194), .ZN(n1187) );
XOR2_X1 U852 ( .A(n1191), .B(n1195), .Z(n1194) );
NOR2_X1 U853 ( .A1(n1193), .A2(n1196), .ZN(n1195) );
INV_X1 U854 ( .A(KEYINPUT15), .ZN(n1196) );
XOR2_X1 U855 ( .A(n1197), .B(n1198), .Z(n1191) );
XOR2_X1 U856 ( .A(n1199), .B(n1200), .Z(n1197) );
NAND2_X1 U857 ( .A1(n1201), .A2(n1153), .ZN(n1199) );
INV_X1 U858 ( .A(n1149), .ZN(n1153) );
NAND2_X1 U859 ( .A1(G902), .A2(n1047), .ZN(n1149) );
NAND3_X1 U860 ( .A1(n1123), .A2(n1202), .A3(n1130), .ZN(n1047) );
AND4_X1 U861 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1130) );
AND4_X1 U862 ( .A1(n1207), .A2(n1208), .A3(n1042), .A4(n1209), .ZN(n1206) );
NAND4_X1 U863 ( .A1(n1055), .A2(n1210), .A3(n1211), .A4(n1074), .ZN(n1042) );
NOR2_X1 U864 ( .A1(n1212), .A2(n1073), .ZN(n1211) );
NOR2_X1 U865 ( .A1(n1161), .A2(n1213), .ZN(n1205) );
NOR2_X1 U866 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U867 ( .A(n1216), .B(KEYINPUT0), .Z(n1214) );
INV_X1 U868 ( .A(n1160), .ZN(n1161) );
NAND3_X1 U869 ( .A1(n1074), .A2(n1056), .A3(n1217), .ZN(n1160) );
XOR2_X1 U870 ( .A(KEYINPUT41), .B(n1124), .Z(n1202) );
AND3_X1 U871 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1124) );
NOR4_X1 U872 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1220) );
NOR2_X1 U873 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
INV_X1 U874 ( .A(KEYINPUT11), .ZN(n1225) );
NOR4_X1 U875 ( .A1(KEYINPUT11), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1223) );
NAND2_X1 U876 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND3_X1 U877 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1227) );
NOR3_X1 U878 ( .A1(n1049), .A2(n1235), .A3(n1236), .ZN(n1222) );
NOR3_X1 U879 ( .A1(n1066), .A2(n1237), .A3(n1238), .ZN(n1221) );
NAND2_X1 U880 ( .A1(n1239), .A2(n1238), .ZN(n1218) );
INV_X1 U881 ( .A(KEYINPUT62), .ZN(n1238) );
AND4_X1 U882 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1123) );
XNOR2_X1 U883 ( .A(G210), .B(KEYINPUT45), .ZN(n1201) );
NOR2_X1 U884 ( .A1(n1059), .A2(G952), .ZN(n1141) );
XNOR2_X1 U885 ( .A(G146), .B(n1219), .ZN(G48) );
NAND3_X1 U886 ( .A1(n1234), .A2(n1057), .A3(n1244), .ZN(n1219) );
XNOR2_X1 U887 ( .A(G143), .B(n1226), .ZN(G45) );
NAND4_X1 U888 ( .A1(n1234), .A2(n1245), .A3(n1230), .A4(n1231), .ZN(n1226) );
XOR2_X1 U889 ( .A(n1239), .B(n1246), .Z(G42) );
NOR2_X1 U890 ( .A1(KEYINPUT29), .A2(n1247), .ZN(n1246) );
NOR2_X1 U891 ( .A1(n1237), .A2(n1049), .ZN(n1239) );
NAND4_X1 U892 ( .A1(n1086), .A2(n1057), .A3(n1074), .A4(n1232), .ZN(n1237) );
XOR2_X1 U893 ( .A(G137), .B(n1248), .Z(G39) );
NOR4_X1 U894 ( .A1(KEYINPUT9), .A2(n1235), .A3(n1236), .A4(n1049), .ZN(n1248) );
XNOR2_X1 U895 ( .A(n1249), .B(n1115), .ZN(G36) );
INV_X1 U896 ( .A(G134), .ZN(n1115) );
NAND2_X1 U897 ( .A1(KEYINPUT36), .A2(n1240), .ZN(n1249) );
NAND3_X1 U898 ( .A1(n1245), .A2(n1055), .A3(n1066), .ZN(n1240) );
XNOR2_X1 U899 ( .A(G131), .B(n1250), .ZN(G33) );
NAND2_X1 U900 ( .A1(KEYINPUT38), .A2(n1251), .ZN(n1250) );
INV_X1 U901 ( .A(n1241), .ZN(n1251) );
NAND3_X1 U902 ( .A1(n1245), .A2(n1057), .A3(n1066), .ZN(n1241) );
INV_X1 U903 ( .A(n1049), .ZN(n1066) );
NAND2_X1 U904 ( .A1(n1084), .A2(n1252), .ZN(n1049) );
INV_X1 U905 ( .A(n1083), .ZN(n1252) );
AND3_X1 U906 ( .A1(n1074), .A2(n1232), .A3(n1079), .ZN(n1245) );
XNOR2_X1 U907 ( .A(G128), .B(n1242), .ZN(G30) );
NAND3_X1 U908 ( .A1(n1234), .A2(n1055), .A3(n1244), .ZN(n1242) );
INV_X1 U909 ( .A(n1236), .ZN(n1244) );
NAND4_X1 U910 ( .A1(n1253), .A2(n1074), .A3(n1254), .A4(n1232), .ZN(n1236) );
XOR2_X1 U911 ( .A(n1208), .B(n1255), .Z(G3) );
XNOR2_X1 U912 ( .A(G101), .B(KEYINPUT22), .ZN(n1255) );
NAND3_X1 U913 ( .A1(n1079), .A2(n1210), .A3(n1256), .ZN(n1208) );
NOR3_X1 U914 ( .A1(n1233), .A2(n1212), .A3(n1235), .ZN(n1256) );
INV_X1 U915 ( .A(n1061), .ZN(n1235) );
INV_X1 U916 ( .A(n1257), .ZN(n1212) );
INV_X1 U917 ( .A(n1074), .ZN(n1233) );
XNOR2_X1 U918 ( .A(G125), .B(n1243), .ZN(G27) );
NAND3_X1 U919 ( .A1(n1086), .A2(n1057), .A3(n1258), .ZN(n1243) );
AND3_X1 U920 ( .A1(n1234), .A2(n1232), .A3(n1054), .ZN(n1258) );
NAND2_X1 U921 ( .A1(n1063), .A2(n1259), .ZN(n1232) );
NAND3_X1 U922 ( .A1(G902), .A2(n1260), .A3(n1108), .ZN(n1259) );
NOR2_X1 U923 ( .A1(n1059), .A2(G900), .ZN(n1108) );
XNOR2_X1 U924 ( .A(n1207), .B(n1261), .ZN(G24) );
NOR2_X1 U925 ( .A1(KEYINPUT30), .A2(n1262), .ZN(n1261) );
NAND4_X1 U926 ( .A1(n1263), .A2(n1056), .A3(n1230), .A4(n1231), .ZN(n1207) );
INV_X1 U927 ( .A(n1073), .ZN(n1056) );
NAND2_X1 U928 ( .A1(n1264), .A2(n1088), .ZN(n1073) );
XOR2_X1 U929 ( .A(G119), .B(n1265), .Z(G21) );
NOR2_X1 U930 ( .A1(KEYINPUT58), .A2(n1203), .ZN(n1265) );
NAND4_X1 U931 ( .A1(n1253), .A2(n1263), .A3(n1061), .A4(n1254), .ZN(n1203) );
XNOR2_X1 U932 ( .A(G116), .B(n1204), .ZN(G18) );
NAND3_X1 U933 ( .A1(n1263), .A2(n1055), .A3(n1079), .ZN(n1204) );
NOR2_X1 U934 ( .A1(n1230), .A2(n1266), .ZN(n1055) );
AND3_X1 U935 ( .A1(n1054), .A2(n1257), .A3(n1234), .ZN(n1263) );
INV_X1 U936 ( .A(n1081), .ZN(n1234) );
XOR2_X1 U937 ( .A(n1210), .B(KEYINPUT37), .Z(n1081) );
XNOR2_X1 U938 ( .A(G113), .B(n1209), .ZN(G15) );
NAND3_X1 U939 ( .A1(n1079), .A2(n1054), .A3(n1217), .ZN(n1209) );
AND3_X1 U940 ( .A1(n1210), .A2(n1257), .A3(n1057), .ZN(n1217) );
NOR2_X1 U941 ( .A1(n1267), .A2(n1072), .ZN(n1054) );
INV_X1 U942 ( .A(n1228), .ZN(n1079) );
NAND2_X1 U943 ( .A1(n1088), .A2(n1253), .ZN(n1228) );
INV_X1 U944 ( .A(n1254), .ZN(n1088) );
XOR2_X1 U945 ( .A(G110), .B(n1268), .Z(G12) );
NOR2_X1 U946 ( .A1(n1215), .A2(n1216), .ZN(n1268) );
NAND4_X1 U947 ( .A1(n1086), .A2(n1074), .A3(n1061), .A4(n1257), .ZN(n1216) );
NAND2_X1 U948 ( .A1(n1063), .A2(n1269), .ZN(n1257) );
NAND4_X1 U949 ( .A1(G953), .A2(G902), .A3(n1260), .A4(n1270), .ZN(n1269) );
INV_X1 U950 ( .A(G898), .ZN(n1270) );
NAND3_X1 U951 ( .A1(n1260), .A2(n1059), .A3(G952), .ZN(n1063) );
NAND2_X1 U952 ( .A1(G237), .A2(G234), .ZN(n1260) );
NAND2_X1 U953 ( .A1(n1271), .A2(n1272), .ZN(n1061) );
OR3_X1 U954 ( .A1(n1230), .A2(n1231), .A3(KEYINPUT32), .ZN(n1272) );
NAND2_X1 U955 ( .A1(KEYINPUT32), .A2(n1057), .ZN(n1271) );
AND2_X1 U956 ( .A1(n1266), .A2(n1230), .ZN(n1057) );
XOR2_X1 U957 ( .A(n1095), .B(n1096), .Z(n1230) );
XNOR2_X1 U958 ( .A(G475), .B(KEYINPUT24), .ZN(n1096) );
NAND2_X1 U959 ( .A1(n1156), .A2(n1273), .ZN(n1095) );
XOR2_X1 U960 ( .A(n1274), .B(n1275), .Z(n1156) );
XOR2_X1 U961 ( .A(n1276), .B(n1277), .Z(n1275) );
NOR3_X1 U962 ( .A1(n1278), .A2(G953), .A3(G237), .ZN(n1276) );
XOR2_X1 U963 ( .A(n1279), .B(n1280), .Z(n1274) );
NOR2_X1 U964 ( .A1(KEYINPUT57), .A2(n1281), .ZN(n1280) );
XOR2_X1 U965 ( .A(n1282), .B(n1283), .Z(n1281) );
NOR2_X1 U966 ( .A1(KEYINPUT14), .A2(G104), .ZN(n1283) );
XNOR2_X1 U967 ( .A(G113), .B(G122), .ZN(n1282) );
XNOR2_X1 U968 ( .A(G143), .B(G131), .ZN(n1279) );
INV_X1 U969 ( .A(n1231), .ZN(n1266) );
XOR2_X1 U970 ( .A(n1097), .B(n1099), .Z(n1231) );
INV_X1 U971 ( .A(G478), .ZN(n1099) );
NAND2_X1 U972 ( .A1(n1152), .A2(n1273), .ZN(n1097) );
XNOR2_X1 U973 ( .A(n1284), .B(n1285), .ZN(n1152) );
XNOR2_X1 U974 ( .A(n1286), .B(n1136), .ZN(n1285) );
XNOR2_X1 U975 ( .A(G116), .B(n1262), .ZN(n1136) );
NAND2_X1 U976 ( .A1(G217), .A2(n1287), .ZN(n1286) );
XOR2_X1 U977 ( .A(n1288), .B(n1289), .Z(n1284) );
NOR2_X1 U978 ( .A1(KEYINPUT52), .A2(n1290), .ZN(n1289) );
XNOR2_X1 U979 ( .A(G107), .B(G134), .ZN(n1288) );
NOR2_X1 U980 ( .A1(n1070), .A2(n1072), .ZN(n1074) );
AND2_X1 U981 ( .A1(G221), .A2(n1291), .ZN(n1072) );
OR2_X1 U982 ( .A1(n1292), .A2(G902), .ZN(n1291) );
INV_X1 U983 ( .A(n1267), .ZN(n1070) );
XNOR2_X1 U984 ( .A(n1293), .B(G469), .ZN(n1267) );
NAND2_X1 U985 ( .A1(n1294), .A2(n1273), .ZN(n1293) );
XOR2_X1 U986 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U987 ( .A(n1183), .B(n1297), .ZN(n1296) );
XNOR2_X1 U988 ( .A(KEYINPUT46), .B(n1298), .ZN(n1297) );
NOR2_X1 U989 ( .A1(KEYINPUT16), .A2(n1299), .ZN(n1298) );
XNOR2_X1 U990 ( .A(KEYINPUT28), .B(n1300), .ZN(n1299) );
INV_X1 U991 ( .A(n1181), .ZN(n1300) );
XOR2_X1 U992 ( .A(G140), .B(G110), .Z(n1181) );
AND2_X1 U993 ( .A1(G227), .A2(n1059), .ZN(n1183) );
XNOR2_X1 U994 ( .A(n1301), .B(n1179), .ZN(n1295) );
XOR2_X1 U995 ( .A(n1135), .B(KEYINPUT56), .Z(n1179) );
XNOR2_X1 U996 ( .A(n1175), .B(n1185), .ZN(n1301) );
INV_X1 U997 ( .A(n1121), .ZN(n1185) );
XNOR2_X1 U998 ( .A(n1302), .B(n1303), .ZN(n1121) );
XOR2_X1 U999 ( .A(G128), .B(n1304), .Z(n1303) );
NOR2_X1 U1000 ( .A1(G146), .A2(KEYINPUT2), .ZN(n1304) );
XNOR2_X1 U1001 ( .A(G143), .B(KEYINPUT10), .ZN(n1302) );
AND2_X1 U1002 ( .A1(n1264), .A2(n1254), .ZN(n1086) );
XNOR2_X1 U1003 ( .A(n1305), .B(n1306), .ZN(n1254) );
NOR2_X1 U1004 ( .A1(n1307), .A2(n1148), .ZN(n1306) );
INV_X1 U1005 ( .A(G217), .ZN(n1148) );
NOR2_X1 U1006 ( .A1(G902), .A2(n1292), .ZN(n1307) );
NAND2_X1 U1007 ( .A1(n1146), .A2(n1273), .ZN(n1305) );
XNOR2_X1 U1008 ( .A(n1308), .B(n1309), .ZN(n1146) );
XOR2_X1 U1009 ( .A(G119), .B(n1310), .Z(n1309) );
XOR2_X1 U1010 ( .A(G137), .B(G128), .Z(n1310) );
XOR2_X1 U1011 ( .A(n1311), .B(n1277), .Z(n1308) );
XNOR2_X1 U1012 ( .A(n1312), .B(n1117), .ZN(n1277) );
XNOR2_X1 U1013 ( .A(G125), .B(n1247), .ZN(n1117) );
INV_X1 U1014 ( .A(G140), .ZN(n1247) );
XOR2_X1 U1015 ( .A(n1313), .B(G110), .Z(n1311) );
NAND2_X1 U1016 ( .A1(G221), .A2(n1287), .ZN(n1313) );
NOR2_X1 U1017 ( .A1(n1292), .A2(G953), .ZN(n1287) );
INV_X1 U1018 ( .A(G234), .ZN(n1292) );
XOR2_X1 U1019 ( .A(n1253), .B(KEYINPUT20), .Z(n1264) );
XNOR2_X1 U1020 ( .A(n1092), .B(KEYINPUT35), .ZN(n1253) );
XNOR2_X1 U1021 ( .A(n1314), .B(n1315), .ZN(n1092) );
XOR2_X1 U1022 ( .A(KEYINPUT44), .B(G472), .Z(n1315) );
NAND2_X1 U1023 ( .A1(n1316), .A2(n1273), .ZN(n1314) );
XOR2_X1 U1024 ( .A(n1317), .B(n1318), .Z(n1316) );
XNOR2_X1 U1025 ( .A(n1319), .B(n1166), .ZN(n1318) );
XNOR2_X1 U1026 ( .A(n1320), .B(n1137), .ZN(n1166) );
NAND2_X1 U1027 ( .A1(KEYINPUT3), .A2(n1321), .ZN(n1320) );
INV_X1 U1028 ( .A(G116), .ZN(n1321) );
NAND2_X1 U1029 ( .A1(KEYINPUT40), .A2(n1322), .ZN(n1319) );
XOR2_X1 U1030 ( .A(KEYINPUT21), .B(n1170), .Z(n1322) );
NOR3_X1 U1031 ( .A1(G237), .A2(G953), .A3(n1323), .ZN(n1170) );
XNOR2_X1 U1032 ( .A(n1324), .B(n1325), .ZN(n1317) );
NOR2_X1 U1033 ( .A1(KEYINPUT25), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1034 ( .A(KEYINPUT60), .B(n1165), .Z(n1326) );
XNOR2_X1 U1035 ( .A(n1175), .B(n1200), .ZN(n1165) );
NAND3_X1 U1036 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1175) );
NAND2_X1 U1037 ( .A1(G131), .A2(n1330), .ZN(n1329) );
NAND2_X1 U1038 ( .A1(KEYINPUT31), .A2(n1331), .ZN(n1328) );
NAND2_X1 U1039 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
INV_X1 U1040 ( .A(G131), .ZN(n1333) );
XNOR2_X1 U1041 ( .A(n1334), .B(n1330), .ZN(n1332) );
NAND2_X1 U1042 ( .A1(n1335), .A2(n1336), .ZN(n1327) );
INV_X1 U1043 ( .A(KEYINPUT31), .ZN(n1336) );
NAND2_X1 U1044 ( .A1(n1337), .A2(n1338), .ZN(n1335) );
NAND2_X1 U1045 ( .A1(n1330), .A2(n1334), .ZN(n1338) );
OR3_X1 U1046 ( .A1(n1330), .A2(G131), .A3(n1334), .ZN(n1337) );
INV_X1 U1047 ( .A(KEYINPUT4), .ZN(n1334) );
XOR2_X1 U1048 ( .A(G134), .B(G137), .Z(n1330) );
INV_X1 U1049 ( .A(G101), .ZN(n1324) );
INV_X1 U1050 ( .A(n1210), .ZN(n1215) );
NOR2_X1 U1051 ( .A1(n1084), .A2(n1083), .ZN(n1210) );
NOR2_X1 U1052 ( .A1(n1278), .A2(n1339), .ZN(n1083) );
INV_X1 U1053 ( .A(G214), .ZN(n1278) );
XNOR2_X1 U1054 ( .A(n1093), .B(KEYINPUT43), .ZN(n1084) );
XNOR2_X1 U1055 ( .A(n1340), .B(n1341), .ZN(n1093) );
NOR2_X1 U1056 ( .A1(n1339), .A2(n1323), .ZN(n1341) );
INV_X1 U1057 ( .A(G210), .ZN(n1323) );
NOR2_X1 U1058 ( .A1(G902), .A2(G237), .ZN(n1339) );
NAND2_X1 U1059 ( .A1(n1342), .A2(n1273), .ZN(n1340) );
XOR2_X1 U1060 ( .A(G902), .B(KEYINPUT7), .Z(n1273) );
XOR2_X1 U1061 ( .A(n1193), .B(n1343), .Z(n1342) );
NAND2_X1 U1062 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
OR2_X1 U1063 ( .A1(n1198), .A2(n1200), .ZN(n1345) );
NAND2_X1 U1064 ( .A1(n1346), .A2(n1200), .ZN(n1344) );
XOR2_X1 U1065 ( .A(n1347), .B(n1290), .Z(n1200) );
XNOR2_X1 U1066 ( .A(G128), .B(G143), .ZN(n1290) );
NAND2_X1 U1067 ( .A1(KEYINPUT59), .A2(n1312), .ZN(n1347) );
INV_X1 U1068 ( .A(G146), .ZN(n1312) );
XOR2_X1 U1069 ( .A(KEYINPUT48), .B(n1198), .Z(n1346) );
XOR2_X1 U1070 ( .A(G125), .B(n1348), .Z(n1198) );
AND2_X1 U1071 ( .A1(n1059), .A2(G224), .ZN(n1348) );
INV_X1 U1072 ( .A(G953), .ZN(n1059) );
NAND2_X1 U1073 ( .A1(n1349), .A2(n1350), .ZN(n1193) );
NAND2_X1 U1074 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
XNOR2_X1 U1075 ( .A(n1353), .B(n1354), .ZN(n1352) );
XNOR2_X1 U1076 ( .A(n1262), .B(G110), .ZN(n1351) );
INV_X1 U1077 ( .A(G122), .ZN(n1262) );
XOR2_X1 U1078 ( .A(n1355), .B(KEYINPUT55), .Z(n1349) );
NAND2_X1 U1079 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
XNOR2_X1 U1080 ( .A(n1353), .B(n1135), .ZN(n1357) );
INV_X1 U1081 ( .A(n1354), .ZN(n1135) );
XOR2_X1 U1082 ( .A(G101), .B(n1358), .Z(n1354) );
XNOR2_X1 U1083 ( .A(n1359), .B(G104), .ZN(n1358) );
INV_X1 U1084 ( .A(G107), .ZN(n1359) );
NAND2_X1 U1085 ( .A1(n1360), .A2(KEYINPUT33), .ZN(n1353) );
XNOR2_X1 U1086 ( .A(G116), .B(n1137), .ZN(n1360) );
XNOR2_X1 U1087 ( .A(n1361), .B(G119), .ZN(n1137) );
INV_X1 U1088 ( .A(G113), .ZN(n1361) );
XNOR2_X1 U1089 ( .A(G122), .B(G110), .ZN(n1356) );
endmodule


