//Key = 0111110111100010010111100101000111111100110101000000000001110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389;

XNOR2_X1 U760 ( .A(G107), .B(n1056), .ZN(G9) );
NOR2_X1 U761 ( .A1(n1057), .A2(n1058), .ZN(G75) );
NOR4_X1 U762 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1058) );
NOR3_X1 U763 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1061) );
NOR3_X1 U764 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1064) );
AND3_X1 U765 ( .A1(n1069), .A2(n1070), .A3(KEYINPUT56), .ZN(n1068) );
NOR2_X1 U766 ( .A1(n1071), .A2(n1069), .ZN(n1067) );
NOR3_X1 U767 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
NOR2_X1 U768 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U769 ( .A1(KEYINPUT56), .A2(n1077), .ZN(n1073) );
NOR2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1072) );
NOR4_X1 U771 ( .A1(n1080), .A2(n1081), .A3(n1079), .A4(n1082), .ZN(n1066) );
INV_X1 U772 ( .A(n1083), .ZN(n1079) );
XOR2_X1 U773 ( .A(n1069), .B(KEYINPUT47), .Z(n1080) );
NAND3_X1 U774 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1059) );
NAND3_X1 U775 ( .A1(n1087), .A2(n1083), .A3(n1088), .ZN(n1086) );
NOR3_X1 U776 ( .A1(n1076), .A2(n1089), .A3(n1090), .ZN(n1088) );
NOR2_X1 U777 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR2_X1 U778 ( .A1(n1093), .A2(n1063), .ZN(n1092) );
NOR2_X1 U779 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NOR2_X1 U780 ( .A1(n1096), .A2(n1097), .ZN(n1089) );
XOR2_X1 U781 ( .A(KEYINPUT28), .B(n1098), .Z(n1097) );
NOR2_X1 U782 ( .A1(n1099), .A2(n1100), .ZN(n1096) );
NOR2_X1 U783 ( .A1(n1101), .A2(n1065), .ZN(n1099) );
INV_X1 U784 ( .A(n1102), .ZN(n1076) );
INV_X1 U785 ( .A(n1069), .ZN(n1087) );
NOR3_X1 U786 ( .A1(n1103), .A2(G953), .A3(G952), .ZN(n1057) );
INV_X1 U787 ( .A(n1084), .ZN(n1103) );
NAND4_X1 U788 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1084) );
NOR4_X1 U789 ( .A1(n1108), .A2(n1109), .A3(n1110), .A4(n1111), .ZN(n1107) );
XNOR2_X1 U790 ( .A(G475), .B(n1112), .ZN(n1111) );
XOR2_X1 U791 ( .A(n1113), .B(n1114), .Z(n1110) );
NOR2_X1 U792 ( .A1(n1115), .A2(n1116), .ZN(n1109) );
INV_X1 U793 ( .A(KEYINPUT46), .ZN(n1116) );
NOR3_X1 U794 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1115) );
AND2_X1 U795 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
INV_X1 U796 ( .A(G469), .ZN(n1117) );
NOR2_X1 U797 ( .A1(KEYINPUT46), .A2(n1091), .ZN(n1108) );
NOR2_X1 U798 ( .A1(n1122), .A2(n1123), .ZN(n1106) );
XOR2_X1 U799 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND2_X1 U800 ( .A1(KEYINPUT37), .A2(n1126), .ZN(n1124) );
INV_X1 U801 ( .A(n1081), .ZN(n1122) );
NAND2_X1 U802 ( .A1(n1127), .A2(n1128), .ZN(G72) );
NAND3_X1 U803 ( .A1(G953), .A2(n1129), .A3(n1130), .ZN(n1128) );
XOR2_X1 U804 ( .A(KEYINPUT57), .B(n1131), .Z(n1127) );
NOR2_X1 U805 ( .A1(n1132), .A2(n1130), .ZN(n1131) );
AND2_X1 U806 ( .A1(n1133), .A2(n1134), .ZN(n1130) );
NAND3_X1 U807 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1134) );
NAND2_X1 U808 ( .A1(G953), .A2(n1138), .ZN(n1136) );
XOR2_X1 U809 ( .A(n1139), .B(n1140), .Z(n1135) );
NAND2_X1 U810 ( .A1(n1141), .A2(n1142), .ZN(n1133) );
INV_X1 U811 ( .A(n1137), .ZN(n1142) );
NAND2_X1 U812 ( .A1(n1085), .A2(n1143), .ZN(n1137) );
NAND4_X1 U813 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1143) );
NOR2_X1 U814 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XNOR2_X1 U815 ( .A(n1139), .B(n1140), .ZN(n1141) );
XNOR2_X1 U816 ( .A(n1150), .B(G125), .ZN(n1140) );
NAND2_X1 U817 ( .A1(KEYINPUT19), .A2(n1151), .ZN(n1150) );
NAND2_X1 U818 ( .A1(n1152), .A2(KEYINPUT1), .ZN(n1139) );
XOR2_X1 U819 ( .A(n1153), .B(KEYINPUT6), .Z(n1152) );
AND2_X1 U820 ( .A1(n1129), .A2(G953), .ZN(n1132) );
NAND2_X1 U821 ( .A1(G900), .A2(G227), .ZN(n1129) );
XOR2_X1 U822 ( .A(n1154), .B(n1155), .Z(G69) );
XOR2_X1 U823 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U824 ( .A1(G953), .A2(n1158), .ZN(n1157) );
NAND2_X1 U825 ( .A1(G898), .A2(G224), .ZN(n1158) );
NAND3_X1 U826 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1156) );
NAND2_X1 U827 ( .A1(G953), .A2(n1162), .ZN(n1161) );
NAND2_X1 U828 ( .A1(KEYINPUT12), .A2(n1163), .ZN(n1160) );
NAND2_X1 U829 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U830 ( .A1(n1166), .A2(n1167), .ZN(n1159) );
INV_X1 U831 ( .A(KEYINPUT12), .ZN(n1167) );
NOR2_X1 U832 ( .A1(n1168), .A2(G953), .ZN(n1154) );
NOR2_X1 U833 ( .A1(n1169), .A2(n1170), .ZN(G66) );
XOR2_X1 U834 ( .A(n1171), .B(n1172), .Z(n1170) );
XNOR2_X1 U835 ( .A(n1173), .B(KEYINPUT15), .ZN(n1172) );
NAND3_X1 U836 ( .A1(n1174), .A2(G217), .A3(KEYINPUT61), .ZN(n1173) );
NOR2_X1 U837 ( .A1(n1169), .A2(n1175), .ZN(G63) );
XOR2_X1 U838 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U839 ( .A1(n1126), .A2(n1178), .ZN(n1177) );
INV_X1 U840 ( .A(G478), .ZN(n1126) );
NAND2_X1 U841 ( .A1(KEYINPUT14), .A2(n1179), .ZN(n1176) );
XNOR2_X1 U842 ( .A(KEYINPUT33), .B(n1180), .ZN(n1179) );
NOR2_X1 U843 ( .A1(n1169), .A2(n1181), .ZN(G60) );
XOR2_X1 U844 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U845 ( .A(KEYINPUT45), .B(n1184), .Z(n1183) );
AND2_X1 U846 ( .A1(G475), .A2(n1174), .ZN(n1184) );
XNOR2_X1 U847 ( .A(G104), .B(n1185), .ZN(G6) );
NOR2_X1 U848 ( .A1(n1169), .A2(n1186), .ZN(G57) );
XOR2_X1 U849 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U850 ( .A(n1189), .B(n1190), .Z(n1188) );
NAND3_X1 U851 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1189) );
NAND2_X1 U852 ( .A1(KEYINPUT42), .A2(n1194), .ZN(n1193) );
OR3_X1 U853 ( .A1(n1195), .A2(KEYINPUT42), .A3(n1196), .ZN(n1192) );
NAND2_X1 U854 ( .A1(n1195), .A2(n1196), .ZN(n1191) );
NAND2_X1 U855 ( .A1(KEYINPUT40), .A2(n1197), .ZN(n1195) );
INV_X1 U856 ( .A(n1194), .ZN(n1197) );
XNOR2_X1 U857 ( .A(G101), .B(KEYINPUT3), .ZN(n1194) );
XOR2_X1 U858 ( .A(n1198), .B(n1199), .Z(n1187) );
NOR3_X1 U859 ( .A1(n1178), .A2(KEYINPUT55), .A3(n1200), .ZN(n1199) );
INV_X1 U860 ( .A(G472), .ZN(n1200) );
NAND2_X1 U861 ( .A1(n1201), .A2(n1202), .ZN(n1198) );
NAND2_X1 U862 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
XOR2_X1 U863 ( .A(KEYINPUT4), .B(n1205), .Z(n1201) );
NOR2_X1 U864 ( .A1(n1203), .A2(n1204), .ZN(n1205) );
INV_X1 U865 ( .A(n1206), .ZN(n1203) );
NOR2_X1 U866 ( .A1(n1169), .A2(n1207), .ZN(G54) );
XOR2_X1 U867 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U868 ( .A(n1210), .B(n1211), .Z(n1209) );
NAND2_X1 U869 ( .A1(n1212), .A2(n1213), .ZN(n1210) );
OR2_X1 U870 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U871 ( .A(n1216), .B(KEYINPUT52), .Z(n1212) );
NAND2_X1 U872 ( .A1(n1215), .A2(n1214), .ZN(n1216) );
XNOR2_X1 U873 ( .A(n1217), .B(n1218), .ZN(n1214) );
XOR2_X1 U874 ( .A(n1219), .B(n1220), .Z(n1208) );
NAND3_X1 U875 ( .A1(n1174), .A2(G469), .A3(KEYINPUT5), .ZN(n1219) );
INV_X1 U876 ( .A(n1178), .ZN(n1174) );
NOR2_X1 U877 ( .A1(n1169), .A2(n1221), .ZN(G51) );
XOR2_X1 U878 ( .A(n1222), .B(n1223), .Z(n1221) );
XOR2_X1 U879 ( .A(n1224), .B(n1225), .Z(n1223) );
NAND2_X1 U880 ( .A1(KEYINPUT41), .A2(G125), .ZN(n1224) );
XOR2_X1 U881 ( .A(n1206), .B(n1226), .Z(n1222) );
NOR2_X1 U882 ( .A1(n1227), .A2(n1178), .ZN(n1226) );
NAND2_X1 U883 ( .A1(G902), .A2(n1228), .ZN(n1178) );
NAND2_X1 U884 ( .A1(n1229), .A2(n1168), .ZN(n1228) );
INV_X1 U885 ( .A(n1062), .ZN(n1168) );
NAND4_X1 U886 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1062) );
AND4_X1 U887 ( .A1(n1234), .A2(n1056), .A3(n1185), .A4(n1235), .ZN(n1233) );
NAND3_X1 U888 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1185) );
NAND3_X1 U889 ( .A1(n1236), .A2(n1239), .A3(n1237), .ZN(n1056) );
NOR2_X1 U890 ( .A1(n1240), .A2(n1241), .ZN(n1232) );
NOR4_X1 U891 ( .A1(n1242), .A2(n1243), .A3(n1075), .A4(n1244), .ZN(n1241) );
NOR2_X1 U892 ( .A1(n1245), .A2(n1246), .ZN(n1243) );
INV_X1 U893 ( .A(KEYINPUT13), .ZN(n1246) );
NOR3_X1 U894 ( .A1(n1065), .A2(n1247), .A3(n1248), .ZN(n1245) );
NOR2_X1 U895 ( .A1(KEYINPUT13), .A2(n1249), .ZN(n1242) );
INV_X1 U896 ( .A(n1250), .ZN(n1240) );
XOR2_X1 U897 ( .A(n1060), .B(KEYINPUT20), .Z(n1229) );
NAND4_X1 U898 ( .A1(n1146), .A2(n1144), .A3(n1251), .A4(n1252), .ZN(n1060) );
NOR2_X1 U899 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
XOR2_X1 U900 ( .A(n1145), .B(KEYINPUT17), .Z(n1254) );
XOR2_X1 U901 ( .A(n1149), .B(KEYINPUT23), .Z(n1253) );
NAND4_X1 U902 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1149) );
NAND3_X1 U903 ( .A1(n1259), .A2(n1247), .A3(n1091), .ZN(n1255) );
INV_X1 U904 ( .A(n1065), .ZN(n1091) );
NOR2_X1 U905 ( .A1(n1085), .A2(G952), .ZN(n1169) );
XOR2_X1 U906 ( .A(G146), .B(n1148), .Z(G48) );
INV_X1 U907 ( .A(n1251), .ZN(n1148) );
NAND3_X1 U908 ( .A1(n1260), .A2(n1247), .A3(n1238), .ZN(n1251) );
XOR2_X1 U909 ( .A(n1261), .B(G143), .Z(G45) );
NAND2_X1 U910 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
OR2_X1 U911 ( .A1(n1145), .A2(KEYINPUT16), .ZN(n1263) );
NAND2_X1 U912 ( .A1(n1264), .A2(n1247), .ZN(n1145) );
NAND3_X1 U913 ( .A1(n1264), .A2(n1078), .A3(KEYINPUT16), .ZN(n1262) );
AND3_X1 U914 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1264) );
XOR2_X1 U915 ( .A(n1146), .B(n1268), .Z(G42) );
XOR2_X1 U916 ( .A(KEYINPUT62), .B(G140), .Z(n1268) );
NAND3_X1 U917 ( .A1(n1102), .A2(n1269), .A3(n1259), .ZN(n1146) );
XNOR2_X1 U918 ( .A(G137), .B(n1144), .ZN(G39) );
NAND3_X1 U919 ( .A1(n1260), .A2(n1102), .A3(n1083), .ZN(n1144) );
XNOR2_X1 U920 ( .A(G134), .B(n1256), .ZN(G36) );
NAND3_X1 U921 ( .A1(n1102), .A2(n1239), .A3(n1267), .ZN(n1256) );
XOR2_X1 U922 ( .A(n1257), .B(n1270), .Z(G33) );
XOR2_X1 U923 ( .A(KEYINPUT22), .B(G131), .Z(n1270) );
NAND2_X1 U924 ( .A1(n1070), .A2(n1267), .ZN(n1257) );
AND2_X1 U925 ( .A1(n1271), .A2(n1272), .ZN(n1267) );
INV_X1 U926 ( .A(n1077), .ZN(n1070) );
NAND2_X1 U927 ( .A1(n1238), .A2(n1102), .ZN(n1077) );
NOR2_X1 U928 ( .A1(n1082), .A2(n1273), .ZN(n1102) );
INV_X1 U929 ( .A(n1274), .ZN(n1273) );
XNOR2_X1 U930 ( .A(n1104), .B(KEYINPUT39), .ZN(n1082) );
XOR2_X1 U931 ( .A(n1258), .B(n1275), .Z(G30) );
NOR2_X1 U932 ( .A1(G128), .A2(KEYINPUT30), .ZN(n1275) );
NAND3_X1 U933 ( .A1(n1239), .A2(n1247), .A3(n1260), .ZN(n1258) );
AND4_X1 U934 ( .A1(n1269), .A2(n1101), .A3(n1100), .A4(n1272), .ZN(n1260) );
NAND2_X1 U935 ( .A1(n1276), .A2(n1277), .ZN(G3) );
NAND2_X1 U936 ( .A1(G101), .A2(n1250), .ZN(n1277) );
XOR2_X1 U937 ( .A(n1278), .B(KEYINPUT24), .Z(n1276) );
OR2_X1 U938 ( .A1(n1250), .A2(G101), .ZN(n1278) );
NAND4_X1 U939 ( .A1(n1271), .A2(n1083), .A3(n1247), .A4(n1279), .ZN(n1250) );
AND2_X1 U940 ( .A1(n1098), .A2(n1269), .ZN(n1271) );
XOR2_X1 U941 ( .A(n1280), .B(n1281), .Z(G27) );
NAND2_X1 U942 ( .A1(KEYINPUT43), .A2(G125), .ZN(n1281) );
NAND3_X1 U943 ( .A1(n1259), .A2(n1247), .A3(n1282), .ZN(n1280) );
XOR2_X1 U944 ( .A(n1065), .B(KEYINPUT36), .Z(n1282) );
AND4_X1 U945 ( .A1(n1105), .A2(n1238), .A3(n1101), .A4(n1272), .ZN(n1259) );
NAND2_X1 U946 ( .A1(n1069), .A2(n1283), .ZN(n1272) );
NAND4_X1 U947 ( .A1(G953), .A2(G902), .A3(n1284), .A4(n1138), .ZN(n1283) );
INV_X1 U948 ( .A(G900), .ZN(n1138) );
XOR2_X1 U949 ( .A(n1285), .B(n1230), .Z(G24) );
NAND4_X1 U950 ( .A1(n1286), .A2(n1249), .A3(n1265), .A4(n1266), .ZN(n1230) );
INV_X1 U951 ( .A(n1063), .ZN(n1286) );
NAND2_X1 U952 ( .A1(n1236), .A2(n1105), .ZN(n1063) );
XNOR2_X1 U953 ( .A(G119), .B(n1231), .ZN(G21) );
NAND4_X1 U954 ( .A1(n1249), .A2(n1083), .A3(n1101), .A4(n1100), .ZN(n1231) );
NAND2_X1 U955 ( .A1(n1287), .A2(n1288), .ZN(G18) );
OR2_X1 U956 ( .A1(n1289), .A2(G116), .ZN(n1288) );
XOR2_X1 U957 ( .A(n1290), .B(KEYINPUT60), .Z(n1287) );
NAND2_X1 U958 ( .A1(G116), .A2(n1289), .ZN(n1290) );
NAND3_X1 U959 ( .A1(n1098), .A2(n1239), .A3(n1249), .ZN(n1289) );
INV_X1 U960 ( .A(n1075), .ZN(n1239) );
NAND2_X1 U961 ( .A1(n1291), .A2(n1266), .ZN(n1075) );
XNOR2_X1 U962 ( .A(G113), .B(n1235), .ZN(G15) );
NAND3_X1 U963 ( .A1(n1098), .A2(n1238), .A3(n1249), .ZN(n1235) );
NOR3_X1 U964 ( .A1(n1078), .A2(n1248), .A3(n1065), .ZN(n1249) );
NAND2_X1 U965 ( .A1(n1094), .A2(n1095), .ZN(n1065) );
INV_X1 U966 ( .A(n1279), .ZN(n1248) );
NOR2_X1 U967 ( .A1(n1291), .A2(n1266), .ZN(n1238) );
INV_X1 U968 ( .A(n1265), .ZN(n1291) );
INV_X1 U969 ( .A(n1244), .ZN(n1098) );
NAND2_X1 U970 ( .A1(n1236), .A2(n1100), .ZN(n1244) );
INV_X1 U971 ( .A(n1105), .ZN(n1100) );
XNOR2_X1 U972 ( .A(G110), .B(n1234), .ZN(G12) );
NAND3_X1 U973 ( .A1(n1237), .A2(n1101), .A3(n1083), .ZN(n1234) );
NOR2_X1 U974 ( .A1(n1266), .A2(n1265), .ZN(n1083) );
XNOR2_X1 U975 ( .A(G475), .B(n1292), .ZN(n1265) );
NOR2_X1 U976 ( .A1(KEYINPUT26), .A2(n1293), .ZN(n1292) );
XOR2_X1 U977 ( .A(n1112), .B(KEYINPUT35), .Z(n1293) );
NAND2_X1 U978 ( .A1(n1182), .A2(n1120), .ZN(n1112) );
XOR2_X1 U979 ( .A(n1294), .B(n1295), .Z(n1182) );
XOR2_X1 U980 ( .A(G104), .B(n1296), .Z(n1295) );
NOR2_X1 U981 ( .A1(KEYINPUT54), .A2(n1297), .ZN(n1296) );
NOR2_X1 U982 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
XOR2_X1 U983 ( .A(KEYINPUT29), .B(n1300), .Z(n1299) );
AND2_X1 U984 ( .A1(n1285), .A2(G113), .ZN(n1300) );
NOR2_X1 U985 ( .A1(G113), .A2(n1285), .ZN(n1298) );
NAND2_X1 U986 ( .A1(n1301), .A2(KEYINPUT27), .ZN(n1294) );
XOR2_X1 U987 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U988 ( .A(G146), .B(G131), .Z(n1303) );
XNOR2_X1 U989 ( .A(n1304), .B(n1305), .ZN(n1302) );
NAND3_X1 U990 ( .A1(n1306), .A2(n1307), .A3(KEYINPUT21), .ZN(n1305) );
NAND2_X1 U991 ( .A1(G125), .A2(n1151), .ZN(n1307) );
XOR2_X1 U992 ( .A(KEYINPUT59), .B(n1308), .Z(n1306) );
NOR2_X1 U993 ( .A1(G125), .A2(n1151), .ZN(n1308) );
NAND2_X1 U994 ( .A1(n1309), .A2(KEYINPUT2), .ZN(n1304) );
XOR2_X1 U995 ( .A(n1310), .B(G143), .Z(n1309) );
NAND2_X1 U996 ( .A1(n1311), .A2(G214), .ZN(n1310) );
XOR2_X1 U997 ( .A(n1125), .B(G478), .Z(n1266) );
AND2_X1 U998 ( .A1(n1120), .A2(n1180), .ZN(n1125) );
NAND2_X1 U999 ( .A1(n1312), .A2(n1313), .ZN(n1180) );
NAND2_X1 U1000 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
XOR2_X1 U1001 ( .A(n1316), .B(n1317), .Z(n1312) );
AND2_X1 U1002 ( .A1(n1318), .A2(G217), .ZN(n1317) );
OR2_X1 U1003 ( .A1(n1315), .A2(n1314), .ZN(n1316) );
XNOR2_X1 U1004 ( .A(n1319), .B(n1320), .ZN(n1314) );
XOR2_X1 U1005 ( .A(G116), .B(n1321), .Z(n1320) );
XOR2_X1 U1006 ( .A(KEYINPUT53), .B(G134), .Z(n1321) );
XOR2_X1 U1007 ( .A(n1322), .B(n1323), .Z(n1319) );
XOR2_X1 U1008 ( .A(n1324), .B(G107), .Z(n1322) );
NAND2_X1 U1009 ( .A1(KEYINPUT9), .A2(n1285), .ZN(n1324) );
INV_X1 U1010 ( .A(G122), .ZN(n1285) );
INV_X1 U1011 ( .A(KEYINPUT10), .ZN(n1315) );
INV_X1 U1012 ( .A(n1236), .ZN(n1101) );
XOR2_X1 U1013 ( .A(n1325), .B(n1326), .Z(n1236) );
XNOR2_X1 U1014 ( .A(KEYINPUT25), .B(n1113), .ZN(n1326) );
NAND2_X1 U1015 ( .A1(G217), .A2(n1327), .ZN(n1113) );
NAND2_X1 U1016 ( .A1(KEYINPUT58), .A2(n1114), .ZN(n1325) );
OR2_X1 U1017 ( .A1(n1171), .A2(G902), .ZN(n1114) );
XNOR2_X1 U1018 ( .A(n1328), .B(n1329), .ZN(n1171) );
XNOR2_X1 U1019 ( .A(n1330), .B(n1331), .ZN(n1329) );
NOR2_X1 U1020 ( .A1(G137), .A2(KEYINPUT38), .ZN(n1331) );
NAND2_X1 U1021 ( .A1(n1332), .A2(KEYINPUT31), .ZN(n1330) );
XOR2_X1 U1022 ( .A(n1333), .B(n1334), .Z(n1332) );
XOR2_X1 U1023 ( .A(G119), .B(G110), .Z(n1334) );
NAND3_X1 U1024 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1333) );
OR2_X1 U1025 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
NAND3_X1 U1026 ( .A1(n1338), .A2(n1340), .A3(n1341), .ZN(n1336) );
NAND2_X1 U1027 ( .A1(n1342), .A2(G146), .ZN(n1335) );
XOR2_X1 U1028 ( .A(n1340), .B(n1338), .Z(n1342) );
NAND2_X1 U1029 ( .A1(KEYINPUT63), .A2(n1343), .ZN(n1338) );
XOR2_X1 U1030 ( .A(n1151), .B(n1344), .Z(n1343) );
NAND2_X1 U1031 ( .A1(KEYINPUT8), .A2(n1345), .ZN(n1344) );
NAND2_X1 U1032 ( .A1(n1318), .A2(G221), .ZN(n1328) );
AND2_X1 U1033 ( .A1(G234), .A2(n1085), .ZN(n1318) );
AND4_X1 U1034 ( .A1(n1247), .A2(n1269), .A3(n1105), .A4(n1279), .ZN(n1237) );
NAND2_X1 U1035 ( .A1(n1069), .A2(n1346), .ZN(n1279) );
NAND4_X1 U1036 ( .A1(G953), .A2(G902), .A3(n1284), .A4(n1162), .ZN(n1346) );
INV_X1 U1037 ( .A(G898), .ZN(n1162) );
NAND3_X1 U1038 ( .A1(n1284), .A2(n1085), .A3(G952), .ZN(n1069) );
NAND2_X1 U1039 ( .A1(G237), .A2(G234), .ZN(n1284) );
XOR2_X1 U1040 ( .A(n1347), .B(G472), .Z(n1105) );
NAND2_X1 U1041 ( .A1(n1348), .A2(n1120), .ZN(n1347) );
XOR2_X1 U1042 ( .A(n1349), .B(n1350), .Z(n1348) );
XOR2_X1 U1043 ( .A(n1206), .B(n1351), .Z(n1350) );
XNOR2_X1 U1044 ( .A(G101), .B(KEYINPUT7), .ZN(n1351) );
XOR2_X1 U1045 ( .A(n1352), .B(n1190), .Z(n1349) );
XOR2_X1 U1046 ( .A(n1204), .B(n1196), .Z(n1352) );
NAND2_X1 U1047 ( .A1(n1311), .A2(G210), .ZN(n1196) );
NOR2_X1 U1048 ( .A1(G953), .A2(G237), .ZN(n1311) );
NOR2_X1 U1049 ( .A1(n1094), .A2(n1118), .ZN(n1269) );
INV_X1 U1050 ( .A(n1095), .ZN(n1118) );
NAND2_X1 U1051 ( .A1(G221), .A2(n1327), .ZN(n1095) );
NAND2_X1 U1052 ( .A1(G234), .A2(n1120), .ZN(n1327) );
XOR2_X1 U1053 ( .A(n1353), .B(G469), .Z(n1094) );
NAND2_X1 U1054 ( .A1(n1121), .A2(n1120), .ZN(n1353) );
XNOR2_X1 U1055 ( .A(n1354), .B(n1355), .ZN(n1121) );
XOR2_X1 U1056 ( .A(n1220), .B(n1356), .Z(n1355) );
NOR2_X1 U1057 ( .A1(KEYINPUT49), .A2(n1218), .ZN(n1356) );
XNOR2_X1 U1058 ( .A(n1357), .B(n1358), .ZN(n1218) );
NOR2_X1 U1059 ( .A1(G107), .A2(KEYINPUT44), .ZN(n1358) );
XNOR2_X1 U1060 ( .A(G104), .B(G101), .ZN(n1357) );
AND2_X1 U1061 ( .A1(G227), .A2(n1085), .ZN(n1220) );
XOR2_X1 U1062 ( .A(n1153), .B(n1359), .Z(n1354) );
NOR2_X1 U1063 ( .A1(KEYINPUT50), .A2(n1211), .ZN(n1359) );
XOR2_X1 U1064 ( .A(G110), .B(n1151), .Z(n1211) );
INV_X1 U1065 ( .A(G140), .ZN(n1151) );
XOR2_X1 U1066 ( .A(n1217), .B(n1204), .Z(n1153) );
INV_X1 U1067 ( .A(n1215), .ZN(n1204) );
XNOR2_X1 U1068 ( .A(G131), .B(n1360), .ZN(n1215) );
XOR2_X1 U1069 ( .A(G137), .B(G134), .Z(n1360) );
XOR2_X1 U1070 ( .A(n1341), .B(n1323), .Z(n1217) );
INV_X1 U1071 ( .A(n1078), .ZN(n1247) );
NAND2_X1 U1072 ( .A1(n1361), .A2(n1274), .ZN(n1078) );
XOR2_X1 U1073 ( .A(n1081), .B(KEYINPUT18), .Z(n1274) );
NAND2_X1 U1074 ( .A1(G214), .A2(n1362), .ZN(n1081) );
XOR2_X1 U1075 ( .A(n1104), .B(KEYINPUT32), .Z(n1361) );
XNOR2_X1 U1076 ( .A(n1363), .B(n1227), .ZN(n1104) );
NAND2_X1 U1077 ( .A1(G210), .A2(n1362), .ZN(n1227) );
NAND2_X1 U1078 ( .A1(n1364), .A2(n1120), .ZN(n1362) );
INV_X1 U1079 ( .A(G237), .ZN(n1364) );
NAND2_X1 U1080 ( .A1(n1365), .A2(n1120), .ZN(n1363) );
INV_X1 U1081 ( .A(G902), .ZN(n1120) );
XOR2_X1 U1082 ( .A(n1366), .B(n1367), .Z(n1365) );
XOR2_X1 U1083 ( .A(n1345), .B(n1206), .Z(n1367) );
NAND3_X1 U1084 ( .A1(n1368), .A2(n1369), .A3(n1370), .ZN(n1206) );
OR2_X1 U1085 ( .A1(n1371), .A2(n1339), .ZN(n1370) );
NAND2_X1 U1086 ( .A1(n1372), .A2(n1373), .ZN(n1369) );
INV_X1 U1087 ( .A(KEYINPUT34), .ZN(n1373) );
NAND3_X1 U1088 ( .A1(n1374), .A2(n1375), .A3(n1339), .ZN(n1372) );
NAND2_X1 U1089 ( .A1(G128), .A2(n1341), .ZN(n1339) );
NAND3_X1 U1090 ( .A1(G146), .A2(n1340), .A3(n1371), .ZN(n1375) );
NAND2_X1 U1091 ( .A1(G143), .A2(G128), .ZN(n1374) );
NAND2_X1 U1092 ( .A1(KEYINPUT34), .A2(n1376), .ZN(n1368) );
NAND2_X1 U1093 ( .A1(n1377), .A2(n1378), .ZN(n1376) );
NAND3_X1 U1094 ( .A1(n1340), .A2(n1371), .A3(n1341), .ZN(n1378) );
INV_X1 U1095 ( .A(G146), .ZN(n1341) );
INV_X1 U1096 ( .A(G143), .ZN(n1371) );
INV_X1 U1097 ( .A(G128), .ZN(n1340) );
NAND2_X1 U1098 ( .A1(n1323), .A2(G146), .ZN(n1377) );
XOR2_X1 U1099 ( .A(G143), .B(G128), .Z(n1323) );
INV_X1 U1100 ( .A(G125), .ZN(n1345) );
INV_X1 U1101 ( .A(n1225), .ZN(n1366) );
XOR2_X1 U1102 ( .A(n1379), .B(n1166), .Z(n1225) );
XNOR2_X1 U1103 ( .A(n1165), .B(n1164), .ZN(n1166) );
XOR2_X1 U1104 ( .A(n1380), .B(n1381), .Z(n1164) );
XOR2_X1 U1105 ( .A(KEYINPUT51), .B(KEYINPUT48), .Z(n1381) );
XNOR2_X1 U1106 ( .A(n1190), .B(n1382), .ZN(n1380) );
NOR2_X1 U1107 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
XOR2_X1 U1108 ( .A(KEYINPUT11), .B(n1385), .Z(n1384) );
NOR2_X1 U1109 ( .A1(G101), .A2(n1386), .ZN(n1385) );
NOR2_X1 U1110 ( .A1(n1387), .A2(n1388), .ZN(n1383) );
XNOR2_X1 U1111 ( .A(G101), .B(KEYINPUT0), .ZN(n1388) );
INV_X1 U1112 ( .A(n1386), .ZN(n1387) );
XOR2_X1 U1113 ( .A(G104), .B(G107), .Z(n1386) );
XOR2_X1 U1114 ( .A(G113), .B(n1389), .Z(n1190) );
XOR2_X1 U1115 ( .A(G119), .B(G116), .Z(n1389) );
XOR2_X1 U1116 ( .A(G110), .B(G122), .Z(n1165) );
NAND2_X1 U1117 ( .A1(G224), .A2(n1085), .ZN(n1379) );
INV_X1 U1118 ( .A(G953), .ZN(n1085) );
endmodule


