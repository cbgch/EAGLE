//Key = 0100000001000101001000011011001010110001010100100111111110101101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327;

XNOR2_X1 U728 ( .A(G107), .B(n1003), .ZN(G9) );
NAND4_X1 U729 ( .A1(n1004), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(G75) );
NOR2_X1 U730 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NOR4_X1 U731 ( .A1(n1010), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1008) );
NAND3_X1 U732 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1011) );
NAND4_X1 U733 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1010) );
NOR3_X1 U734 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
AND3_X1 U735 ( .A1(KEYINPUT52), .A2(n1024), .A3(G475), .ZN(n1023) );
NOR2_X1 U736 ( .A1(KEYINPUT52), .A2(G475), .ZN(n1022) );
XNOR2_X1 U737 ( .A(G478), .B(n1025), .ZN(n1021) );
XNOR2_X1 U738 ( .A(G472), .B(n1026), .ZN(n1019) );
NOR2_X1 U739 ( .A1(KEYINPUT29), .A2(n1027), .ZN(n1026) );
XNOR2_X1 U740 ( .A(n1028), .B(n1029), .ZN(n1018) );
NOR2_X1 U741 ( .A1(n1030), .A2(KEYINPUT28), .ZN(n1029) );
INV_X1 U742 ( .A(n1031), .ZN(n1030) );
XOR2_X1 U743 ( .A(n1032), .B(n1033), .Z(n1017) );
XOR2_X1 U744 ( .A(KEYINPUT60), .B(KEYINPUT46), .Z(n1033) );
XOR2_X1 U745 ( .A(n1034), .B(n1035), .Z(n1032) );
NAND3_X1 U746 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1006) );
INV_X1 U747 ( .A(n1039), .ZN(n1038) );
NAND2_X1 U748 ( .A1(n1040), .A2(n1041), .ZN(n1037) );
NAND3_X1 U749 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
NAND2_X1 U750 ( .A1(n1045), .A2(n1046), .ZN(n1040) );
NAND3_X1 U751 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND2_X1 U752 ( .A1(n1042), .A2(n1050), .ZN(n1049) );
NAND2_X1 U753 ( .A1(n1044), .A2(n1051), .ZN(n1048) );
NAND2_X1 U754 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U755 ( .A1(n1013), .A2(n1054), .ZN(n1053) );
NAND2_X1 U756 ( .A1(n1055), .A2(n1056), .ZN(n1047) );
XNOR2_X1 U757 ( .A(KEYINPUT59), .B(n1057), .ZN(n1056) );
NAND4_X1 U758 ( .A1(n1045), .A2(n1058), .A3(n1042), .A4(n1059), .ZN(n1004) );
NOR2_X1 U759 ( .A1(n1060), .A2(n1039), .ZN(n1059) );
NAND2_X1 U760 ( .A1(n1061), .A2(n1062), .ZN(n1058) );
NAND2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
XNOR2_X1 U762 ( .A(KEYINPUT22), .B(n1065), .ZN(n1064) );
NAND2_X1 U763 ( .A1(n1066), .A2(n1067), .ZN(G72) );
NAND2_X1 U764 ( .A1(n1068), .A2(n1005), .ZN(n1067) );
XNOR2_X1 U765 ( .A(n1069), .B(n1070), .ZN(n1068) );
NAND2_X1 U766 ( .A1(n1071), .A2(G953), .ZN(n1066) );
NAND2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1074), .ZN(n1073) );
INV_X1 U769 ( .A(G227), .ZN(n1074) );
NAND2_X1 U770 ( .A1(G227), .A2(n1075), .ZN(n1072) );
NAND2_X1 U771 ( .A1(G900), .A2(n1070), .ZN(n1075) );
NAND2_X1 U772 ( .A1(n1076), .A2(n1077), .ZN(n1070) );
NAND2_X1 U773 ( .A1(G953), .A2(n1078), .ZN(n1077) );
XOR2_X1 U774 ( .A(n1079), .B(n1080), .Z(n1076) );
XNOR2_X1 U775 ( .A(n1081), .B(n1082), .ZN(n1080) );
INV_X1 U776 ( .A(n1083), .ZN(n1082) );
XOR2_X1 U777 ( .A(n1084), .B(n1085), .Z(n1079) );
XOR2_X1 U778 ( .A(n1086), .B(KEYINPUT8), .Z(n1084) );
NAND3_X1 U779 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
OR2_X1 U780 ( .A1(n1090), .A2(KEYINPUT49), .ZN(n1089) );
NAND3_X1 U781 ( .A1(KEYINPUT49), .A2(n1090), .A3(G134), .ZN(n1088) );
NAND2_X1 U782 ( .A1(n1091), .A2(n1092), .ZN(n1087) );
NAND2_X1 U783 ( .A1(KEYINPUT49), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U784 ( .A(KEYINPUT53), .B(n1090), .ZN(n1093) );
XOR2_X1 U785 ( .A(n1094), .B(n1095), .Z(G69) );
NOR2_X1 U786 ( .A1(n1096), .A2(n1005), .ZN(n1095) );
NOR2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1094) );
NAND2_X1 U789 ( .A1(n1101), .A2(n1005), .ZN(n1100) );
XNOR2_X1 U790 ( .A(n1102), .B(n1103), .ZN(n1101) );
NOR3_X1 U791 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1103) );
XOR2_X1 U792 ( .A(n1107), .B(KEYINPUT57), .Z(n1106) );
NAND3_X1 U793 ( .A1(G898), .A2(n1102), .A3(G953), .ZN(n1099) );
XOR2_X1 U794 ( .A(n1108), .B(n1109), .Z(n1102) );
NOR2_X1 U795 ( .A1(n1110), .A2(n1111), .ZN(G66) );
XOR2_X1 U796 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND3_X1 U797 ( .A1(n1114), .A2(n1035), .A3(KEYINPUT51), .ZN(n1112) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(G63) );
XNOR2_X1 U799 ( .A(n1117), .B(n1118), .ZN(n1116) );
NOR2_X1 U800 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NOR2_X1 U801 ( .A1(G952), .A2(n1121), .ZN(n1115) );
XNOR2_X1 U802 ( .A(G953), .B(KEYINPUT38), .ZN(n1121) );
NOR3_X1 U803 ( .A1(n1110), .A2(n1122), .A3(n1123), .ZN(G60) );
NOR2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U805 ( .A(n1126), .B(KEYINPUT41), .Z(n1125) );
NOR2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(n1122) );
XOR2_X1 U807 ( .A(n1126), .B(KEYINPUT37), .Z(n1128) );
NAND2_X1 U808 ( .A1(n1114), .A2(G475), .ZN(n1126) );
INV_X1 U809 ( .A(n1120), .ZN(n1114) );
XOR2_X1 U810 ( .A(G104), .B(n1105), .Z(G6) );
NOR2_X1 U811 ( .A1(n1110), .A2(n1129), .ZN(G57) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1129) );
XNOR2_X1 U813 ( .A(G101), .B(n1132), .ZN(n1130) );
NOR2_X1 U814 ( .A1(n1133), .A2(n1120), .ZN(n1132) );
NOR3_X1 U815 ( .A1(n1110), .A2(n1134), .A3(n1135), .ZN(G54) );
NOR2_X1 U816 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
INV_X1 U817 ( .A(n1138), .ZN(n1137) );
NOR2_X1 U818 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
NOR2_X1 U819 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NOR2_X1 U820 ( .A1(n1143), .A2(n1144), .ZN(n1139) );
NOR2_X1 U821 ( .A1(n1138), .A2(n1145), .ZN(n1134) );
NOR2_X1 U822 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NOR2_X1 U823 ( .A1(n1144), .A2(n1141), .ZN(n1147) );
INV_X1 U824 ( .A(n1143), .ZN(n1141) );
XOR2_X1 U825 ( .A(KEYINPUT45), .B(n1148), .Z(n1144) );
NOR2_X1 U826 ( .A1(n1143), .A2(n1142), .ZN(n1146) );
XNOR2_X1 U827 ( .A(KEYINPUT2), .B(n1148), .ZN(n1142) );
NOR2_X1 U828 ( .A1(n1120), .A2(n1149), .ZN(n1148) );
XNOR2_X1 U829 ( .A(n1150), .B(n1151), .ZN(n1143) );
XNOR2_X1 U830 ( .A(n1152), .B(n1092), .ZN(n1150) );
INV_X1 U831 ( .A(G134), .ZN(n1092) );
NAND3_X1 U832 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1152) );
NAND2_X1 U833 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
OR3_X1 U834 ( .A1(n1157), .A2(n1156), .A3(n1158), .ZN(n1154) );
INV_X1 U835 ( .A(KEYINPUT35), .ZN(n1157) );
NAND2_X1 U836 ( .A1(n1158), .A2(n1159), .ZN(n1153) );
NAND2_X1 U837 ( .A1(KEYINPUT35), .A2(n1160), .ZN(n1159) );
XOR2_X1 U838 ( .A(KEYINPUT63), .B(n1156), .Z(n1160) );
XNOR2_X1 U839 ( .A(n1083), .B(n1161), .ZN(n1158) );
XOR2_X1 U840 ( .A(G128), .B(n1162), .Z(n1083) );
NOR2_X1 U841 ( .A1(n1110), .A2(n1163), .ZN(G51) );
XOR2_X1 U842 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U843 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U844 ( .A(n1168), .B(n1169), .Z(n1164) );
NOR2_X1 U845 ( .A1(G125), .A2(KEYINPUT36), .ZN(n1169) );
NOR2_X1 U846 ( .A1(n1031), .A2(n1120), .ZN(n1168) );
NAND2_X1 U847 ( .A1(G902), .A2(n1009), .ZN(n1120) );
OR4_X1 U848 ( .A1(n1069), .A2(n1107), .A3(n1104), .A4(n1105), .ZN(n1009) );
AND2_X1 U849 ( .A1(n1055), .A2(n1170), .ZN(n1105) );
NAND2_X1 U850 ( .A1(n1003), .A2(n1171), .ZN(n1104) );
NAND2_X1 U851 ( .A1(n1172), .A2(n1043), .ZN(n1171) );
NAND2_X1 U852 ( .A1(n1173), .A2(n1174), .ZN(n1043) );
NAND2_X1 U853 ( .A1(n1050), .A2(n1170), .ZN(n1003) );
AND3_X1 U854 ( .A1(n1045), .A2(n1175), .A3(n1176), .ZN(n1170) );
NAND4_X1 U855 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1107) );
NAND4_X1 U856 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1069) );
NOR4_X1 U857 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1184) );
INV_X1 U858 ( .A(n1189), .ZN(n1187) );
NAND2_X1 U859 ( .A1(n1042), .A2(n1190), .ZN(n1183) );
NAND2_X1 U860 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NOR2_X1 U861 ( .A1(n1005), .A2(G952), .ZN(n1110) );
XNOR2_X1 U862 ( .A(G146), .B(n1181), .ZN(G48) );
NAND3_X1 U863 ( .A1(n1055), .A2(n1176), .A3(n1193), .ZN(n1181) );
XNOR2_X1 U864 ( .A(G143), .B(n1182), .ZN(G45) );
NAND3_X1 U865 ( .A1(n1194), .A2(n1176), .A3(n1195), .ZN(n1182) );
NOR3_X1 U866 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1195) );
XOR2_X1 U867 ( .A(n1188), .B(n1199), .Z(G42) );
NOR2_X1 U868 ( .A1(KEYINPUT33), .A2(n1200), .ZN(n1199) );
AND3_X1 U869 ( .A1(n1055), .A2(n1201), .A3(n1202), .ZN(n1188) );
XOR2_X1 U870 ( .A(n1203), .B(n1204), .Z(G39) );
NAND2_X1 U871 ( .A1(KEYINPUT56), .A2(n1205), .ZN(n1204) );
XNOR2_X1 U872 ( .A(KEYINPUT62), .B(n1090), .ZN(n1205) );
NAND2_X1 U873 ( .A1(n1206), .A2(n1042), .ZN(n1203) );
INV_X1 U874 ( .A(n1057), .ZN(n1042) );
XOR2_X1 U875 ( .A(n1192), .B(KEYINPUT32), .Z(n1206) );
NAND3_X1 U876 ( .A1(n1193), .A2(n1207), .A3(n1044), .ZN(n1192) );
XNOR2_X1 U877 ( .A(G134), .B(n1189), .ZN(G36) );
NAND3_X1 U878 ( .A1(n1202), .A2(n1050), .A3(n1194), .ZN(n1189) );
NOR3_X1 U879 ( .A1(n1062), .A2(n1197), .A3(n1057), .ZN(n1202) );
INV_X1 U880 ( .A(n1208), .ZN(n1197) );
XNOR2_X1 U881 ( .A(n1209), .B(n1210), .ZN(G33) );
NOR2_X1 U882 ( .A1(n1211), .A2(n1057), .ZN(n1210) );
NAND2_X1 U883 ( .A1(n1054), .A2(n1212), .ZN(n1057) );
XOR2_X1 U884 ( .A(n1191), .B(KEYINPUT6), .Z(n1211) );
NAND4_X1 U885 ( .A1(n1194), .A2(n1055), .A3(n1207), .A4(n1208), .ZN(n1191) );
INV_X1 U886 ( .A(n1062), .ZN(n1207) );
XOR2_X1 U887 ( .A(n1186), .B(n1213), .Z(G30) );
NOR2_X1 U888 ( .A1(KEYINPUT7), .A2(n1214), .ZN(n1213) );
AND3_X1 U889 ( .A1(n1050), .A2(n1176), .A3(n1193), .ZN(n1186) );
AND3_X1 U890 ( .A1(n1215), .A2(n1208), .A3(n1216), .ZN(n1193) );
XOR2_X1 U891 ( .A(n1217), .B(n1218), .Z(G3) );
NOR2_X1 U892 ( .A1(KEYINPUT14), .A2(n1219), .ZN(n1218) );
NOR4_X1 U893 ( .A1(n1220), .A2(n1221), .A3(n1173), .A4(n1060), .ZN(n1217) );
INV_X1 U894 ( .A(n1044), .ZN(n1060) );
INV_X1 U895 ( .A(n1194), .ZN(n1173) );
INV_X1 U896 ( .A(n1176), .ZN(n1221) );
XOR2_X1 U897 ( .A(n1175), .B(KEYINPUT15), .Z(n1220) );
XOR2_X1 U898 ( .A(G125), .B(n1185), .Z(G27) );
AND3_X1 U899 ( .A1(n1055), .A2(n1201), .A3(n1222), .ZN(n1185) );
AND3_X1 U900 ( .A1(n1036), .A2(n1208), .A3(n1223), .ZN(n1222) );
NAND2_X1 U901 ( .A1(n1039), .A2(n1224), .ZN(n1208) );
NAND4_X1 U902 ( .A1(G953), .A2(G902), .A3(n1225), .A4(n1078), .ZN(n1224) );
INV_X1 U903 ( .A(G900), .ZN(n1078) );
XNOR2_X1 U904 ( .A(G122), .B(n1177), .ZN(G24) );
NAND4_X1 U905 ( .A1(n1226), .A2(n1045), .A3(n1227), .A4(n1228), .ZN(n1177) );
NOR2_X1 U906 ( .A1(n1215), .A2(n1229), .ZN(n1045) );
XOR2_X1 U907 ( .A(n1230), .B(G119), .Z(G21) );
NAND2_X1 U908 ( .A1(KEYINPUT30), .A2(n1180), .ZN(n1230) );
NAND4_X1 U909 ( .A1(n1226), .A2(n1044), .A3(n1216), .A4(n1215), .ZN(n1180) );
XNOR2_X1 U910 ( .A(G116), .B(n1178), .ZN(G18) );
NAND3_X1 U911 ( .A1(n1194), .A2(n1050), .A3(n1226), .ZN(n1178) );
NOR2_X1 U912 ( .A1(n1231), .A2(n1196), .ZN(n1050) );
XNOR2_X1 U913 ( .A(G113), .B(n1179), .ZN(G15) );
NAND3_X1 U914 ( .A1(n1194), .A2(n1055), .A3(n1226), .ZN(n1179) );
AND3_X1 U915 ( .A1(n1223), .A2(n1175), .A3(n1036), .ZN(n1226) );
NOR2_X1 U916 ( .A1(n1065), .A2(n1063), .ZN(n1036) );
INV_X1 U917 ( .A(n1016), .ZN(n1063) );
NOR2_X1 U918 ( .A1(n1198), .A2(n1227), .ZN(n1055) );
INV_X1 U919 ( .A(n1228), .ZN(n1198) );
XNOR2_X1 U920 ( .A(n1231), .B(KEYINPUT58), .ZN(n1228) );
NOR2_X1 U921 ( .A1(n1229), .A2(n1232), .ZN(n1194) );
INV_X1 U922 ( .A(n1233), .ZN(n1229) );
XNOR2_X1 U923 ( .A(n1234), .B(n1235), .ZN(G12) );
NAND2_X1 U924 ( .A1(KEYINPUT43), .A2(n1236), .ZN(n1234) );
NAND2_X1 U925 ( .A1(n1172), .A2(n1201), .ZN(n1236) );
INV_X1 U926 ( .A(n1174), .ZN(n1201) );
NAND2_X1 U927 ( .A1(n1232), .A2(n1216), .ZN(n1174) );
XNOR2_X1 U928 ( .A(n1233), .B(KEYINPUT16), .ZN(n1216) );
XNOR2_X1 U929 ( .A(n1034), .B(n1237), .ZN(n1233) );
NOR2_X1 U930 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NOR2_X1 U931 ( .A1(KEYINPUT54), .A2(n1035), .ZN(n1239) );
AND2_X1 U932 ( .A1(KEYINPUT1), .A2(n1035), .ZN(n1238) );
AND2_X1 U933 ( .A1(G217), .A2(n1240), .ZN(n1035) );
NAND2_X1 U934 ( .A1(n1113), .A2(n1241), .ZN(n1034) );
XNOR2_X1 U935 ( .A(n1242), .B(n1243), .ZN(n1113) );
XOR2_X1 U936 ( .A(n1244), .B(n1245), .Z(n1243) );
XNOR2_X1 U937 ( .A(n1246), .B(n1235), .ZN(n1245) );
INV_X1 U938 ( .A(G110), .ZN(n1235) );
NAND2_X1 U939 ( .A1(G221), .A2(n1247), .ZN(n1246) );
NAND2_X1 U940 ( .A1(n1248), .A2(n1249), .ZN(n1244) );
NAND2_X1 U941 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
XNOR2_X1 U942 ( .A(n1252), .B(KEYINPUT20), .ZN(n1250) );
NAND2_X1 U943 ( .A1(n1253), .A2(G146), .ZN(n1248) );
XNOR2_X1 U944 ( .A(KEYINPUT42), .B(n1254), .ZN(n1253) );
INV_X1 U945 ( .A(n1252), .ZN(n1254) );
XOR2_X1 U946 ( .A(G140), .B(n1255), .Z(n1252) );
NOR2_X1 U947 ( .A1(KEYINPUT19), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U948 ( .A(G125), .B(KEYINPUT47), .ZN(n1256) );
XNOR2_X1 U949 ( .A(G119), .B(n1257), .ZN(n1242) );
XNOR2_X1 U950 ( .A(n1090), .B(G128), .ZN(n1257) );
INV_X1 U951 ( .A(n1215), .ZN(n1232) );
XOR2_X1 U952 ( .A(n1027), .B(n1133), .Z(n1215) );
INV_X1 U953 ( .A(G472), .ZN(n1133) );
NAND2_X1 U954 ( .A1(n1258), .A2(n1241), .ZN(n1027) );
XNOR2_X1 U955 ( .A(n1131), .B(n1259), .ZN(n1258) );
XOR2_X1 U956 ( .A(KEYINPUT44), .B(n1260), .Z(n1259) );
NOR2_X1 U957 ( .A1(G101), .A2(KEYINPUT31), .ZN(n1260) );
XNOR2_X1 U958 ( .A(n1261), .B(n1262), .ZN(n1131) );
XOR2_X1 U959 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U960 ( .A(G113), .B(n1265), .Z(n1264) );
NOR2_X1 U961 ( .A1(KEYINPUT11), .A2(n1266), .ZN(n1265) );
XNOR2_X1 U962 ( .A(G116), .B(G119), .ZN(n1266) );
AND3_X1 U963 ( .A1(G210), .A2(n1005), .A3(n1267), .ZN(n1263) );
XOR2_X1 U964 ( .A(n1268), .B(n1269), .Z(n1261) );
XNOR2_X1 U965 ( .A(n1151), .B(n1270), .ZN(n1268) );
AND3_X1 U966 ( .A1(n1176), .A2(n1175), .A3(n1044), .ZN(n1172) );
NOR2_X1 U967 ( .A1(n1231), .A2(n1227), .ZN(n1044) );
INV_X1 U968 ( .A(n1196), .ZN(n1227) );
NAND3_X1 U969 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1196) );
OR2_X1 U970 ( .A1(n1119), .A2(KEYINPUT9), .ZN(n1273) );
INV_X1 U971 ( .A(G478), .ZN(n1119) );
NAND3_X1 U972 ( .A1(KEYINPUT9), .A2(n1274), .A3(n1025), .ZN(n1272) );
OR2_X1 U973 ( .A1(n1025), .A2(n1274), .ZN(n1271) );
NOR2_X1 U974 ( .A1(G478), .A2(KEYINPUT48), .ZN(n1274) );
NAND2_X1 U975 ( .A1(n1118), .A2(n1241), .ZN(n1025) );
XOR2_X1 U976 ( .A(n1275), .B(n1276), .Z(n1118) );
XOR2_X1 U977 ( .A(G116), .B(n1277), .Z(n1276) );
XOR2_X1 U978 ( .A(KEYINPUT24), .B(G122), .Z(n1277) );
XOR2_X1 U979 ( .A(n1278), .B(n1279), .Z(n1275) );
XOR2_X1 U980 ( .A(n1280), .B(G107), .Z(n1278) );
NAND2_X1 U981 ( .A1(G217), .A2(n1247), .ZN(n1280) );
AND2_X1 U982 ( .A1(G234), .A2(n1005), .ZN(n1247) );
NAND2_X1 U983 ( .A1(n1014), .A2(n1281), .ZN(n1231) );
NAND2_X1 U984 ( .A1(G475), .A2(n1024), .ZN(n1281) );
OR2_X1 U985 ( .A1(n1024), .A2(G475), .ZN(n1014) );
NAND2_X1 U986 ( .A1(n1124), .A2(n1241), .ZN(n1024) );
INV_X1 U987 ( .A(n1127), .ZN(n1124) );
XNOR2_X1 U988 ( .A(n1282), .B(n1283), .ZN(n1127) );
XOR2_X1 U989 ( .A(n1284), .B(n1285), .Z(n1283) );
NOR2_X1 U990 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U991 ( .A(n1288), .B(KEYINPUT61), .Z(n1287) );
NAND2_X1 U992 ( .A1(G104), .A2(n1289), .ZN(n1288) );
NOR2_X1 U993 ( .A1(G104), .A2(n1289), .ZN(n1286) );
XOR2_X1 U994 ( .A(G122), .B(G113), .Z(n1289) );
AND3_X1 U995 ( .A1(G214), .A2(n1005), .A3(n1267), .ZN(n1284) );
XOR2_X1 U996 ( .A(n1290), .B(n1085), .Z(n1282) );
XNOR2_X1 U997 ( .A(n1209), .B(G143), .ZN(n1085) );
INV_X1 U998 ( .A(G131), .ZN(n1209) );
NAND2_X1 U999 ( .A1(KEYINPUT23), .A2(n1291), .ZN(n1290) );
XNOR2_X1 U1000 ( .A(n1292), .B(n1081), .ZN(n1291) );
XNOR2_X1 U1001 ( .A(G125), .B(n1200), .ZN(n1081) );
NAND2_X1 U1002 ( .A1(KEYINPUT39), .A2(n1251), .ZN(n1292) );
NAND2_X1 U1003 ( .A1(n1039), .A2(n1293), .ZN(n1175) );
NAND4_X1 U1004 ( .A1(G953), .A2(G902), .A3(n1225), .A4(n1098), .ZN(n1293) );
INV_X1 U1005 ( .A(G898), .ZN(n1098) );
NAND3_X1 U1006 ( .A1(n1225), .A2(n1005), .A3(G952), .ZN(n1039) );
NAND2_X1 U1007 ( .A1(G237), .A2(G234), .ZN(n1225) );
NOR2_X1 U1008 ( .A1(n1062), .A2(n1052), .ZN(n1176) );
INV_X1 U1009 ( .A(n1223), .ZN(n1052) );
NOR2_X1 U1010 ( .A1(n1054), .A2(n1013), .ZN(n1223) );
INV_X1 U1011 ( .A(n1212), .ZN(n1013) );
NAND2_X1 U1012 ( .A1(G214), .A2(n1294), .ZN(n1212) );
XOR2_X1 U1013 ( .A(n1028), .B(n1295), .Z(n1054) );
NOR2_X1 U1014 ( .A1(KEYINPUT25), .A2(n1031), .ZN(n1295) );
NAND2_X1 U1015 ( .A1(G210), .A2(n1294), .ZN(n1031) );
NAND2_X1 U1016 ( .A1(n1267), .A2(n1296), .ZN(n1294) );
INV_X1 U1017 ( .A(G237), .ZN(n1267) );
NAND2_X1 U1018 ( .A1(n1297), .A2(n1241), .ZN(n1028) );
XOR2_X1 U1019 ( .A(n1298), .B(n1166), .Z(n1297) );
XNOR2_X1 U1020 ( .A(n1299), .B(n1109), .ZN(n1166) );
XNOR2_X1 U1021 ( .A(n1300), .B(n1301), .ZN(n1109) );
XNOR2_X1 U1022 ( .A(G110), .B(n1302), .ZN(n1301) );
NAND3_X1 U1023 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(n1302) );
NAND2_X1 U1024 ( .A1(KEYINPUT10), .A2(G101), .ZN(n1305) );
OR3_X1 U1025 ( .A1(n1306), .A2(KEYINPUT10), .A3(n1307), .ZN(n1304) );
NAND2_X1 U1026 ( .A1(n1307), .A2(n1306), .ZN(n1303) );
NAND2_X1 U1027 ( .A1(n1308), .A2(n1219), .ZN(n1306) );
XNOR2_X1 U1028 ( .A(KEYINPUT40), .B(KEYINPUT4), .ZN(n1308) );
XNOR2_X1 U1029 ( .A(G122), .B(KEYINPUT13), .ZN(n1300) );
NAND2_X1 U1030 ( .A1(KEYINPUT18), .A2(n1108), .ZN(n1299) );
XNOR2_X1 U1031 ( .A(n1309), .B(n1310), .ZN(n1108) );
NOR2_X1 U1032 ( .A1(KEYINPUT5), .A2(G116), .ZN(n1310) );
XNOR2_X1 U1033 ( .A(G113), .B(G119), .ZN(n1309) );
NOR2_X1 U1034 ( .A1(KEYINPUT3), .A2(n1311), .ZN(n1298) );
XNOR2_X1 U1035 ( .A(n1167), .B(G125), .ZN(n1311) );
XNOR2_X1 U1036 ( .A(n1312), .B(n1270), .ZN(n1167) );
XNOR2_X1 U1037 ( .A(n1313), .B(n1314), .ZN(n1270) );
NOR2_X1 U1038 ( .A1(G146), .A2(KEYINPUT17), .ZN(n1314) );
XNOR2_X1 U1039 ( .A(G143), .B(KEYINPUT0), .ZN(n1313) );
XNOR2_X1 U1040 ( .A(G128), .B(n1315), .ZN(n1312) );
NOR2_X1 U1041 ( .A1(G953), .A2(n1097), .ZN(n1315) );
INV_X1 U1042 ( .A(G224), .ZN(n1097) );
NAND2_X1 U1043 ( .A1(n1016), .A2(n1065), .ZN(n1062) );
NAND2_X1 U1044 ( .A1(n1316), .A2(n1015), .ZN(n1065) );
NAND2_X1 U1045 ( .A1(n1317), .A2(n1149), .ZN(n1015) );
XNOR2_X1 U1046 ( .A(n1012), .B(KEYINPUT12), .ZN(n1316) );
NOR2_X1 U1047 ( .A1(n1149), .A2(n1317), .ZN(n1012) );
AND2_X1 U1048 ( .A1(n1318), .A2(n1241), .ZN(n1317) );
XNOR2_X1 U1049 ( .A(n1296), .B(KEYINPUT34), .ZN(n1241) );
XNOR2_X1 U1050 ( .A(n1319), .B(n1138), .ZN(n1318) );
XNOR2_X1 U1051 ( .A(n1320), .B(n1321), .ZN(n1138) );
XNOR2_X1 U1052 ( .A(n1200), .B(G110), .ZN(n1321) );
INV_X1 U1053 ( .A(G140), .ZN(n1200) );
NAND2_X1 U1054 ( .A1(G227), .A2(n1005), .ZN(n1320) );
INV_X1 U1055 ( .A(G953), .ZN(n1005) );
NAND2_X1 U1056 ( .A1(n1322), .A2(KEYINPUT55), .ZN(n1319) );
XOR2_X1 U1057 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1058 ( .A(n1151), .B(n1279), .Z(n1324) );
XNOR2_X1 U1059 ( .A(n1161), .B(n1269), .ZN(n1279) );
XNOR2_X1 U1060 ( .A(n1214), .B(G134), .ZN(n1269) );
INV_X1 U1061 ( .A(G128), .ZN(n1214) );
INV_X1 U1062 ( .A(G143), .ZN(n1161) );
XOR2_X1 U1063 ( .A(G131), .B(n1325), .Z(n1151) );
XNOR2_X1 U1064 ( .A(KEYINPUT50), .B(n1090), .ZN(n1325) );
INV_X1 U1065 ( .A(G137), .ZN(n1090) );
XNOR2_X1 U1066 ( .A(n1156), .B(n1162), .ZN(n1323) );
XNOR2_X1 U1067 ( .A(n1251), .B(KEYINPUT26), .ZN(n1162) );
INV_X1 U1068 ( .A(G146), .ZN(n1251) );
XOR2_X1 U1069 ( .A(n1326), .B(n1307), .Z(n1156) );
XNOR2_X1 U1070 ( .A(G107), .B(G104), .ZN(n1307) );
NAND2_X1 U1071 ( .A1(KEYINPUT27), .A2(n1219), .ZN(n1326) );
INV_X1 U1072 ( .A(G101), .ZN(n1219) );
INV_X1 U1073 ( .A(G469), .ZN(n1149) );
NAND2_X1 U1074 ( .A1(n1327), .A2(G221), .ZN(n1016) );
XOR2_X1 U1075 ( .A(n1240), .B(KEYINPUT21), .Z(n1327) );
NAND2_X1 U1076 ( .A1(G234), .A2(n1296), .ZN(n1240) );
INV_X1 U1077 ( .A(G902), .ZN(n1296) );
endmodule


