//Key = 1111111011100100101111011111110001101100111010100101011001010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;

XNOR2_X1 U756 ( .A(G107), .B(n1051), .ZN(G9) );
NOR2_X1 U757 ( .A1(n1052), .A2(n1053), .ZN(G75) );
NOR4_X1 U758 ( .A1(n1054), .A2(n1055), .A3(G953), .A4(n1056), .ZN(n1053) );
NOR2_X1 U759 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U760 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U761 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
INV_X1 U762 ( .A(n1063), .ZN(n1062) );
NOR3_X1 U763 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1061) );
NOR3_X1 U764 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
XNOR2_X1 U765 ( .A(n1070), .B(KEYINPUT48), .ZN(n1068) );
NOR4_X1 U766 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1065) );
NOR2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(n1064) );
INV_X1 U768 ( .A(n1077), .ZN(n1075) );
NOR4_X1 U769 ( .A1(n1071), .A2(n1078), .A3(n1076), .A4(n1079), .ZN(n1059) );
NAND3_X1 U770 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1054) );
XOR2_X1 U771 ( .A(n1083), .B(KEYINPUT46), .Z(n1082) );
NAND2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND4_X1 U773 ( .A1(n1063), .A2(n1070), .A3(n1086), .A4(n1087), .ZN(n1085) );
NOR2_X1 U774 ( .A1(n1067), .A2(n1058), .ZN(n1087) );
NAND3_X1 U775 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1084) );
INV_X1 U776 ( .A(n1058), .ZN(n1090) );
NAND2_X1 U777 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
NAND2_X1 U778 ( .A1(n1070), .A2(n1093), .ZN(n1092) );
NAND2_X1 U779 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U780 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(n1094) );
XNOR2_X1 U782 ( .A(n1063), .B(KEYINPUT49), .ZN(n1098) );
NAND3_X1 U783 ( .A1(n1063), .A2(n1100), .A3(n1096), .ZN(n1091) );
NOR3_X1 U784 ( .A1(n1056), .A2(G953), .A3(G952), .ZN(n1052) );
AND4_X1 U785 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1056) );
NOR4_X1 U786 ( .A1(n1071), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1104) );
XNOR2_X1 U787 ( .A(KEYINPUT50), .B(n1108), .ZN(n1107) );
XNOR2_X1 U788 ( .A(n1109), .B(n1110), .ZN(n1106) );
XNOR2_X1 U789 ( .A(n1111), .B(n1112), .ZN(n1105) );
NAND2_X1 U790 ( .A1(KEYINPUT10), .A2(n1113), .ZN(n1111) );
INV_X1 U791 ( .A(n1070), .ZN(n1071) );
AND3_X1 U792 ( .A1(n1079), .A2(n1073), .A3(n1114), .ZN(n1103) );
NAND2_X1 U793 ( .A1(n1115), .A2(n1116), .ZN(n1101) );
NAND3_X1 U794 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(G72) );
XOR2_X1 U795 ( .A(n1120), .B(KEYINPUT7), .Z(n1119) );
NAND2_X1 U796 ( .A1(G953), .A2(n1121), .ZN(n1120) );
NAND2_X1 U797 ( .A1(G900), .A2(n1122), .ZN(n1121) );
OR2_X1 U798 ( .A1(n1123), .A2(G227), .ZN(n1122) );
NAND2_X1 U799 ( .A1(n1124), .A2(n1125), .ZN(n1118) );
XNOR2_X1 U800 ( .A(n1081), .B(n1123), .ZN(n1124) );
NAND4_X1 U801 ( .A1(G227), .A2(n1123), .A3(G900), .A4(G953), .ZN(n1117) );
XNOR2_X1 U802 ( .A(n1126), .B(n1127), .ZN(n1123) );
NAND2_X1 U803 ( .A1(n1128), .A2(KEYINPUT16), .ZN(n1126) );
XOR2_X1 U804 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U805 ( .A1(KEYINPUT14), .A2(n1131), .ZN(n1130) );
XNOR2_X1 U806 ( .A(n1132), .B(n1133), .ZN(n1129) );
NAND2_X1 U807 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
NAND2_X1 U808 ( .A1(G134), .A2(n1136), .ZN(n1135) );
NAND2_X1 U809 ( .A1(KEYINPUT40), .A2(n1137), .ZN(n1136) );
NAND2_X1 U810 ( .A1(G137), .A2(n1138), .ZN(n1137) );
NAND2_X1 U811 ( .A1(n1139), .A2(n1140), .ZN(n1134) );
NAND2_X1 U812 ( .A1(n1138), .A2(n1141), .ZN(n1139) );
NAND2_X1 U813 ( .A1(KEYINPUT40), .A2(n1142), .ZN(n1141) );
INV_X1 U814 ( .A(KEYINPUT62), .ZN(n1138) );
XOR2_X1 U815 ( .A(n1143), .B(n1144), .Z(G69) );
NOR2_X1 U816 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NOR2_X1 U817 ( .A1(G224), .A2(n1125), .ZN(n1145) );
NAND2_X1 U818 ( .A1(KEYINPUT59), .A2(n1147), .ZN(n1143) );
XOR2_X1 U819 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U820 ( .A1(n1080), .A2(G953), .ZN(n1149) );
NOR2_X1 U821 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
XOR2_X1 U822 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U823 ( .A(KEYINPUT41), .B(n1154), .Z(n1153) );
XNOR2_X1 U824 ( .A(n1146), .B(KEYINPUT6), .ZN(n1150) );
NOR2_X1 U825 ( .A1(n1155), .A2(n1156), .ZN(G66) );
XNOR2_X1 U826 ( .A(n1157), .B(n1158), .ZN(n1156) );
NOR2_X1 U827 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U828 ( .A1(n1161), .A2(n1162), .ZN(G63) );
XOR2_X1 U829 ( .A(KEYINPUT32), .B(n1155), .Z(n1162) );
NOR3_X1 U830 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1161) );
NOR3_X1 U831 ( .A1(n1166), .A2(n1167), .A3(n1160), .ZN(n1165) );
NOR2_X1 U832 ( .A1(n1168), .A2(n1169), .ZN(n1164) );
NOR2_X1 U833 ( .A1(n1170), .A2(n1167), .ZN(n1169) );
XNOR2_X1 U834 ( .A(G478), .B(KEYINPUT17), .ZN(n1167) );
NOR2_X1 U835 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U836 ( .A1(n1155), .A2(n1173), .ZN(G60) );
XNOR2_X1 U837 ( .A(n1174), .B(n1175), .ZN(n1173) );
NOR2_X1 U838 ( .A1(n1176), .A2(n1160), .ZN(n1175) );
XNOR2_X1 U839 ( .A(G104), .B(n1177), .ZN(G6) );
NOR2_X1 U840 ( .A1(n1155), .A2(n1178), .ZN(G57) );
XOR2_X1 U841 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U842 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U843 ( .A1(KEYINPUT63), .A2(n1183), .ZN(n1181) );
XOR2_X1 U844 ( .A(n1184), .B(n1185), .Z(n1179) );
NOR2_X1 U845 ( .A1(n1186), .A2(n1160), .ZN(n1185) );
NAND2_X1 U846 ( .A1(n1187), .A2(n1188), .ZN(n1184) );
OR2_X1 U847 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U848 ( .A(n1191), .B(KEYINPUT47), .Z(n1187) );
NAND2_X1 U849 ( .A1(n1190), .A2(n1189), .ZN(n1191) );
NOR2_X1 U850 ( .A1(n1155), .A2(n1192), .ZN(G54) );
XOR2_X1 U851 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U852 ( .A(n1195), .B(n1196), .Z(n1194) );
NOR2_X1 U853 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
XOR2_X1 U854 ( .A(n1199), .B(KEYINPUT13), .Z(n1198) );
NAND2_X1 U855 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NOR2_X1 U856 ( .A1(n1202), .A2(n1203), .ZN(n1195) );
NOR2_X1 U857 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
INV_X1 U858 ( .A(n1206), .ZN(n1202) );
NOR2_X1 U859 ( .A1(n1207), .A2(n1160), .ZN(n1193) );
NOR2_X1 U860 ( .A1(n1155), .A2(n1208), .ZN(G51) );
XNOR2_X1 U861 ( .A(n1209), .B(n1210), .ZN(n1208) );
XOR2_X1 U862 ( .A(n1211), .B(n1212), .Z(n1210) );
NOR2_X1 U863 ( .A1(n1110), .A2(n1160), .ZN(n1211) );
NAND2_X1 U864 ( .A1(G902), .A2(n1213), .ZN(n1160) );
NAND2_X1 U865 ( .A1(n1080), .A2(n1081), .ZN(n1213) );
INV_X1 U866 ( .A(n1171), .ZN(n1081) );
NAND4_X1 U867 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1171) );
NOR4_X1 U868 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1217) );
NOR2_X1 U869 ( .A1(n1222), .A2(n1223), .ZN(n1216) );
NOR2_X1 U870 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
XNOR2_X1 U871 ( .A(KEYINPUT2), .B(n1067), .ZN(n1225) );
NOR2_X1 U872 ( .A1(n1226), .A2(n1227), .ZN(n1222) );
XNOR2_X1 U873 ( .A(n1228), .B(KEYINPUT12), .ZN(n1226) );
NAND2_X1 U874 ( .A1(n1229), .A2(n1230), .ZN(n1214) );
XNOR2_X1 U875 ( .A(KEYINPUT52), .B(n1227), .ZN(n1230) );
INV_X1 U876 ( .A(n1172), .ZN(n1080) );
NAND2_X1 U877 ( .A1(n1231), .A2(n1232), .ZN(n1172) );
AND4_X1 U878 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1232) );
AND4_X1 U879 ( .A1(n1177), .A2(n1237), .A3(n1051), .A4(n1238), .ZN(n1231) );
NAND3_X1 U880 ( .A1(n1239), .A2(n1070), .A3(n1240), .ZN(n1051) );
OR3_X1 U881 ( .A1(n1241), .A2(n1072), .A3(n1242), .ZN(n1237) );
XNOR2_X1 U882 ( .A(n1243), .B(KEYINPUT42), .ZN(n1241) );
NAND3_X1 U883 ( .A1(n1240), .A2(n1070), .A3(n1086), .ZN(n1177) );
NOR2_X1 U884 ( .A1(n1125), .A2(G952), .ZN(n1155) );
XNOR2_X1 U885 ( .A(G146), .B(n1244), .ZN(G48) );
NAND3_X1 U886 ( .A1(n1228), .A2(n1099), .A3(KEYINPUT20), .ZN(n1244) );
AND3_X1 U887 ( .A1(n1086), .A2(n1245), .A3(n1246), .ZN(n1228) );
XNOR2_X1 U888 ( .A(G143), .B(n1215), .ZN(G45) );
NAND4_X1 U889 ( .A1(n1100), .A2(n1247), .A3(n1099), .A4(n1248), .ZN(n1215) );
NOR2_X1 U890 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
XOR2_X1 U891 ( .A(G140), .B(n1251), .Z(G42) );
NOR2_X1 U892 ( .A1(n1067), .A2(n1224), .ZN(n1251) );
NAND3_X1 U893 ( .A1(n1086), .A2(n1077), .A3(n1246), .ZN(n1224) );
INV_X1 U894 ( .A(n1096), .ZN(n1067) );
NAND2_X1 U895 ( .A1(n1252), .A2(n1253), .ZN(G39) );
OR2_X1 U896 ( .A1(n1254), .A2(G137), .ZN(n1253) );
NAND2_X1 U897 ( .A1(n1255), .A2(G137), .ZN(n1252) );
NAND2_X1 U898 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND2_X1 U899 ( .A1(n1221), .A2(n1258), .ZN(n1257) );
INV_X1 U900 ( .A(KEYINPUT33), .ZN(n1258) );
NAND2_X1 U901 ( .A1(KEYINPUT33), .A2(n1254), .ZN(n1256) );
NAND2_X1 U902 ( .A1(KEYINPUT28), .A2(n1221), .ZN(n1254) );
NOR3_X1 U903 ( .A1(n1249), .A2(n1243), .A3(n1076), .ZN(n1221) );
NAND2_X1 U904 ( .A1(n1096), .A2(n1088), .ZN(n1076) );
XNOR2_X1 U905 ( .A(n1142), .B(n1220), .ZN(G36) );
AND2_X1 U906 ( .A1(n1259), .A2(n1239), .ZN(n1220) );
INV_X1 U907 ( .A(G134), .ZN(n1142) );
NAND3_X1 U908 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(G33) );
OR2_X1 U909 ( .A1(n1219), .A2(KEYINPUT5), .ZN(n1262) );
NAND3_X1 U910 ( .A1(KEYINPUT5), .A2(n1219), .A3(n1133), .ZN(n1261) );
NAND2_X1 U911 ( .A1(G131), .A2(n1263), .ZN(n1260) );
NAND2_X1 U912 ( .A1(n1264), .A2(KEYINPUT5), .ZN(n1263) );
XNOR2_X1 U913 ( .A(n1219), .B(KEYINPUT29), .ZN(n1264) );
AND2_X1 U914 ( .A1(n1259), .A2(n1086), .ZN(n1219) );
AND3_X1 U915 ( .A1(n1096), .A2(n1100), .A3(n1246), .ZN(n1259) );
INV_X1 U916 ( .A(n1249), .ZN(n1246) );
NOR2_X1 U917 ( .A1(n1074), .A2(n1265), .ZN(n1096) );
XOR2_X1 U918 ( .A(KEYINPUT61), .B(n1073), .Z(n1265) );
XOR2_X1 U919 ( .A(G128), .B(n1266), .Z(G30) );
AND2_X1 U920 ( .A1(n1099), .A2(n1229), .ZN(n1266) );
NOR3_X1 U921 ( .A1(n1069), .A2(n1243), .A3(n1249), .ZN(n1229) );
NAND2_X1 U922 ( .A1(n1097), .A2(n1267), .ZN(n1249) );
INV_X1 U923 ( .A(n1239), .ZN(n1069) );
XNOR2_X1 U924 ( .A(G101), .B(n1238), .ZN(G3) );
NAND3_X1 U925 ( .A1(n1240), .A2(n1100), .A3(n1088), .ZN(n1238) );
XOR2_X1 U926 ( .A(G125), .B(n1218), .Z(G27) );
AND4_X1 U927 ( .A1(n1086), .A2(n1063), .A3(n1268), .A4(n1077), .ZN(n1218) );
AND2_X1 U928 ( .A1(n1267), .A2(n1099), .ZN(n1268) );
NAND2_X1 U929 ( .A1(n1269), .A2(n1058), .ZN(n1267) );
NAND4_X1 U930 ( .A1(G902), .A2(G953), .A3(n1270), .A4(n1271), .ZN(n1269) );
INV_X1 U931 ( .A(G900), .ZN(n1271) );
XNOR2_X1 U932 ( .A(G122), .B(n1236), .ZN(G24) );
NAND4_X1 U933 ( .A1(n1272), .A2(n1070), .A3(n1273), .A4(n1247), .ZN(n1236) );
XOR2_X1 U934 ( .A(G119), .B(n1274), .Z(G21) );
NOR3_X1 U935 ( .A1(n1242), .A2(n1243), .A3(n1072), .ZN(n1274) );
INV_X1 U936 ( .A(n1088), .ZN(n1072) );
INV_X1 U937 ( .A(n1245), .ZN(n1243) );
XNOR2_X1 U938 ( .A(G116), .B(n1235), .ZN(G18) );
NAND3_X1 U939 ( .A1(n1239), .A2(n1100), .A3(n1272), .ZN(n1235) );
NOR2_X1 U940 ( .A1(n1247), .A2(n1250), .ZN(n1239) );
XOR2_X1 U941 ( .A(n1234), .B(n1275), .Z(G15) );
NOR2_X1 U942 ( .A1(G113), .A2(KEYINPUT30), .ZN(n1275) );
NAND3_X1 U943 ( .A1(n1086), .A2(n1100), .A3(n1272), .ZN(n1234) );
INV_X1 U944 ( .A(n1242), .ZN(n1272) );
NAND2_X1 U945 ( .A1(n1063), .A2(n1276), .ZN(n1242) );
NOR2_X1 U946 ( .A1(n1078), .A2(n1277), .ZN(n1063) );
INV_X1 U947 ( .A(n1079), .ZN(n1277) );
NAND2_X1 U948 ( .A1(n1278), .A2(n1279), .ZN(n1100) );
NAND2_X1 U949 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
INV_X1 U950 ( .A(KEYINPUT15), .ZN(n1281) );
NAND2_X1 U951 ( .A1(n1282), .A2(n1283), .ZN(n1280) );
NAND3_X1 U952 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1283) );
NAND2_X1 U953 ( .A1(KEYINPUT60), .A2(n1070), .ZN(n1282) );
NOR2_X1 U954 ( .A1(n1287), .A2(n1284), .ZN(n1070) );
NAND2_X1 U955 ( .A1(KEYINPUT15), .A2(n1245), .ZN(n1278) );
NAND2_X1 U956 ( .A1(n1288), .A2(n1289), .ZN(n1245) );
NAND3_X1 U957 ( .A1(n1284), .A2(n1287), .A3(n1286), .ZN(n1289) );
INV_X1 U958 ( .A(KEYINPUT60), .ZN(n1286) );
NAND2_X1 U959 ( .A1(KEYINPUT60), .A2(n1077), .ZN(n1288) );
NOR2_X1 U960 ( .A1(n1273), .A2(n1290), .ZN(n1086) );
INV_X1 U961 ( .A(n1247), .ZN(n1290) );
XNOR2_X1 U962 ( .A(n1291), .B(n1233), .ZN(G12) );
NAND3_X1 U963 ( .A1(n1077), .A2(n1240), .A3(n1088), .ZN(n1233) );
NOR2_X1 U964 ( .A1(n1247), .A2(n1273), .ZN(n1088) );
INV_X1 U965 ( .A(n1250), .ZN(n1273) );
XOR2_X1 U966 ( .A(n1292), .B(n1113), .Z(n1250) );
INV_X1 U967 ( .A(n1163), .ZN(n1113) );
NOR2_X1 U968 ( .A1(n1168), .A2(G902), .ZN(n1163) );
INV_X1 U969 ( .A(n1166), .ZN(n1168) );
NAND2_X1 U970 ( .A1(n1293), .A2(n1294), .ZN(n1166) );
NAND3_X1 U971 ( .A1(n1295), .A2(n1296), .A3(G217), .ZN(n1294) );
INV_X1 U972 ( .A(n1297), .ZN(n1295) );
XOR2_X1 U973 ( .A(n1298), .B(KEYINPUT45), .Z(n1293) );
NAND2_X1 U974 ( .A1(n1297), .A2(n1299), .ZN(n1298) );
NAND2_X1 U975 ( .A1(G217), .A2(n1296), .ZN(n1299) );
XNOR2_X1 U976 ( .A(n1300), .B(n1301), .ZN(n1297) );
XOR2_X1 U977 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U978 ( .A(G107), .B(n1304), .ZN(n1303) );
NOR2_X1 U979 ( .A1(G128), .A2(KEYINPUT58), .ZN(n1304) );
XNOR2_X1 U980 ( .A(G134), .B(n1305), .ZN(n1300) );
XNOR2_X1 U981 ( .A(KEYINPUT8), .B(n1306), .ZN(n1305) );
INV_X1 U982 ( .A(G143), .ZN(n1306) );
NAND2_X1 U983 ( .A1(KEYINPUT57), .A2(n1112), .ZN(n1292) );
XOR2_X1 U984 ( .A(G478), .B(KEYINPUT53), .Z(n1112) );
NAND3_X1 U985 ( .A1(n1307), .A2(n1308), .A3(n1114), .ZN(n1247) );
OR2_X1 U986 ( .A1(n1116), .A2(n1115), .ZN(n1114) );
OR2_X1 U987 ( .A1(n1115), .A2(KEYINPUT54), .ZN(n1308) );
NAND3_X1 U988 ( .A1(n1115), .A2(n1116), .A3(KEYINPUT54), .ZN(n1307) );
NAND2_X1 U989 ( .A1(n1174), .A2(n1309), .ZN(n1116) );
XNOR2_X1 U990 ( .A(n1310), .B(n1311), .ZN(n1174) );
XOR2_X1 U991 ( .A(G104), .B(n1312), .Z(n1311) );
XNOR2_X1 U992 ( .A(n1133), .B(G122), .ZN(n1312) );
INV_X1 U993 ( .A(G131), .ZN(n1133) );
XOR2_X1 U994 ( .A(n1313), .B(n1314), .Z(n1310) );
XOR2_X1 U995 ( .A(n1315), .B(n1316), .Z(n1314) );
NAND2_X1 U996 ( .A1(KEYINPUT51), .A2(n1317), .ZN(n1316) );
INV_X1 U997 ( .A(G113), .ZN(n1317) );
NAND3_X1 U998 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1315) );
NAND2_X1 U999 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
INV_X1 U1000 ( .A(KEYINPUT4), .ZN(n1322) );
NAND3_X1 U1001 ( .A1(KEYINPUT4), .A2(n1323), .A3(n1324), .ZN(n1319) );
OR2_X1 U1002 ( .A1(n1324), .A2(n1323), .ZN(n1318) );
AND2_X1 U1003 ( .A1(n1325), .A2(G214), .ZN(n1323) );
NOR2_X1 U1004 ( .A1(KEYINPUT43), .A2(n1321), .ZN(n1324) );
XNOR2_X1 U1005 ( .A(G143), .B(KEYINPUT36), .ZN(n1321) );
NAND2_X1 U1006 ( .A1(n1326), .A2(n1327), .ZN(n1313) );
NAND2_X1 U1007 ( .A1(G146), .A2(n1127), .ZN(n1327) );
XOR2_X1 U1008 ( .A(n1328), .B(KEYINPUT31), .Z(n1326) );
OR2_X1 U1009 ( .A1(n1127), .A2(G146), .ZN(n1328) );
XNOR2_X1 U1010 ( .A(G140), .B(n1329), .ZN(n1127) );
XOR2_X1 U1011 ( .A(n1176), .B(KEYINPUT3), .Z(n1115) );
INV_X1 U1012 ( .A(G475), .ZN(n1176) );
AND2_X1 U1013 ( .A1(n1276), .A2(n1097), .ZN(n1240) );
AND2_X1 U1014 ( .A1(n1078), .A2(n1079), .ZN(n1097) );
NAND2_X1 U1015 ( .A1(G221), .A2(n1330), .ZN(n1079) );
NAND2_X1 U1016 ( .A1(n1102), .A2(n1108), .ZN(n1078) );
NAND2_X1 U1017 ( .A1(G469), .A2(n1331), .ZN(n1108) );
NAND2_X1 U1018 ( .A1(n1332), .A2(n1309), .ZN(n1331) );
NAND3_X1 U1019 ( .A1(n1207), .A2(n1309), .A3(n1332), .ZN(n1102) );
XOR2_X1 U1020 ( .A(n1333), .B(n1334), .Z(n1332) );
XOR2_X1 U1021 ( .A(n1335), .B(KEYINPUT11), .Z(n1334) );
XNOR2_X1 U1022 ( .A(KEYINPUT39), .B(KEYINPUT34), .ZN(n1335) );
NAND3_X1 U1023 ( .A1(n1336), .A2(n1337), .A3(n1338), .ZN(n1333) );
NAND2_X1 U1024 ( .A1(n1197), .A2(n1339), .ZN(n1338) );
NOR2_X1 U1025 ( .A1(n1201), .A2(n1200), .ZN(n1197) );
OR3_X1 U1026 ( .A1(n1339), .A2(n1340), .A3(n1201), .ZN(n1337) );
INV_X1 U1027 ( .A(n1200), .ZN(n1340) );
NAND2_X1 U1028 ( .A1(n1341), .A2(n1201), .ZN(n1336) );
XNOR2_X1 U1029 ( .A(n1200), .B(n1339), .ZN(n1341) );
NAND3_X1 U1030 ( .A1(n1342), .A2(n1343), .A3(n1206), .ZN(n1339) );
NAND2_X1 U1031 ( .A1(n1204), .A2(n1205), .ZN(n1206) );
NAND2_X1 U1032 ( .A1(KEYINPUT22), .A2(n1205), .ZN(n1343) );
OR3_X1 U1033 ( .A1(n1204), .A2(KEYINPUT22), .A3(n1205), .ZN(n1342) );
XOR2_X1 U1034 ( .A(n1344), .B(G140), .Z(n1205) );
AND2_X1 U1035 ( .A1(G227), .A2(n1125), .ZN(n1204) );
XOR2_X1 U1036 ( .A(n1345), .B(n1346), .Z(n1200) );
XNOR2_X1 U1037 ( .A(G101), .B(n1131), .ZN(n1345) );
XNOR2_X1 U1038 ( .A(n1347), .B(n1348), .ZN(n1131) );
NOR2_X1 U1039 ( .A1(G143), .A2(KEYINPUT38), .ZN(n1348) );
INV_X1 U1040 ( .A(G469), .ZN(n1207) );
AND2_X1 U1041 ( .A1(n1099), .A2(n1349), .ZN(n1276) );
NAND2_X1 U1042 ( .A1(n1058), .A2(n1350), .ZN(n1349) );
NAND3_X1 U1043 ( .A1(n1146), .A2(n1270), .A3(G902), .ZN(n1350) );
NOR2_X1 U1044 ( .A1(G898), .A2(n1125), .ZN(n1146) );
NAND3_X1 U1045 ( .A1(n1270), .A2(n1125), .A3(G952), .ZN(n1058) );
NAND2_X1 U1046 ( .A1(G237), .A2(G234), .ZN(n1270) );
INV_X1 U1047 ( .A(n1227), .ZN(n1099) );
NAND2_X1 U1048 ( .A1(n1074), .A2(n1073), .ZN(n1227) );
NAND2_X1 U1049 ( .A1(G214), .A2(n1351), .ZN(n1073) );
NAND2_X1 U1050 ( .A1(n1352), .A2(n1353), .ZN(n1074) );
OR2_X1 U1051 ( .A1(n1110), .A2(n1109), .ZN(n1353) );
NAND2_X1 U1052 ( .A1(n1354), .A2(n1109), .ZN(n1352) );
AND2_X1 U1053 ( .A1(n1355), .A2(n1309), .ZN(n1109) );
XNOR2_X1 U1054 ( .A(n1356), .B(n1357), .ZN(n1355) );
INV_X1 U1055 ( .A(n1209), .ZN(n1357) );
XNOR2_X1 U1056 ( .A(n1358), .B(n1359), .ZN(n1209) );
XOR2_X1 U1057 ( .A(KEYINPUT9), .B(n1360), .Z(n1359) );
AND2_X1 U1058 ( .A1(n1125), .A2(G224), .ZN(n1360) );
XNOR2_X1 U1059 ( .A(n1152), .B(n1361), .ZN(n1358) );
XNOR2_X1 U1060 ( .A(n1362), .B(n1363), .ZN(n1152) );
XOR2_X1 U1061 ( .A(n1364), .B(n1302), .Z(n1363) );
XNOR2_X1 U1062 ( .A(G122), .B(G116), .ZN(n1302) );
NAND2_X1 U1063 ( .A1(KEYINPUT44), .A2(G113), .ZN(n1364) );
XOR2_X1 U1064 ( .A(n1365), .B(n1366), .Z(n1362) );
XNOR2_X1 U1065 ( .A(KEYINPUT37), .B(n1190), .ZN(n1366) );
INV_X1 U1066 ( .A(G101), .ZN(n1190) );
NAND2_X1 U1067 ( .A1(KEYINPUT26), .A2(n1346), .ZN(n1365) );
XOR2_X1 U1068 ( .A(G104), .B(G107), .Z(n1346) );
NAND2_X1 U1069 ( .A1(KEYINPUT23), .A2(n1367), .ZN(n1356) );
XOR2_X1 U1070 ( .A(KEYINPUT0), .B(n1212), .Z(n1367) );
XNOR2_X1 U1071 ( .A(KEYINPUT1), .B(n1110), .ZN(n1354) );
NAND2_X1 U1072 ( .A1(G210), .A2(n1351), .ZN(n1110) );
NAND2_X1 U1073 ( .A1(n1309), .A2(n1368), .ZN(n1351) );
NOR2_X1 U1074 ( .A1(n1284), .A2(n1285), .ZN(n1077) );
INV_X1 U1075 ( .A(n1287), .ZN(n1285) );
XOR2_X1 U1076 ( .A(n1369), .B(n1159), .Z(n1287) );
NAND2_X1 U1077 ( .A1(G217), .A2(n1330), .ZN(n1159) );
NAND2_X1 U1078 ( .A1(G234), .A2(n1309), .ZN(n1330) );
NAND2_X1 U1079 ( .A1(n1157), .A2(n1309), .ZN(n1369) );
XNOR2_X1 U1080 ( .A(n1370), .B(n1371), .ZN(n1157) );
XOR2_X1 U1081 ( .A(n1361), .B(n1372), .Z(n1371) );
XOR2_X1 U1082 ( .A(n1373), .B(n1374), .Z(n1372) );
NAND2_X1 U1083 ( .A1(KEYINPUT21), .A2(n1375), .ZN(n1374) );
INV_X1 U1084 ( .A(G146), .ZN(n1375) );
NAND2_X1 U1085 ( .A1(n1296), .A2(G221), .ZN(n1373) );
AND2_X1 U1086 ( .A1(G234), .A2(n1125), .ZN(n1296) );
XNOR2_X1 U1087 ( .A(n1329), .B(n1154), .ZN(n1361) );
XNOR2_X1 U1088 ( .A(n1344), .B(G119), .ZN(n1154) );
XNOR2_X1 U1089 ( .A(G125), .B(KEYINPUT55), .ZN(n1329) );
XOR2_X1 U1090 ( .A(n1376), .B(n1377), .Z(n1370) );
XOR2_X1 U1091 ( .A(KEYINPUT27), .B(G140), .Z(n1377) );
XNOR2_X1 U1092 ( .A(G128), .B(G137), .ZN(n1376) );
XOR2_X1 U1093 ( .A(n1378), .B(n1186), .Z(n1284) );
INV_X1 U1094 ( .A(G472), .ZN(n1186) );
NAND2_X1 U1095 ( .A1(n1379), .A2(n1309), .ZN(n1378) );
INV_X1 U1096 ( .A(G902), .ZN(n1309) );
XOR2_X1 U1097 ( .A(n1380), .B(n1381), .Z(n1379) );
XNOR2_X1 U1098 ( .A(n1183), .B(n1182), .ZN(n1381) );
XNOR2_X1 U1099 ( .A(n1382), .B(n1201), .ZN(n1182) );
XOR2_X1 U1100 ( .A(G131), .B(n1383), .Z(n1201) );
XNOR2_X1 U1101 ( .A(n1140), .B(G134), .ZN(n1383) );
INV_X1 U1102 ( .A(G137), .ZN(n1140) );
NAND2_X1 U1103 ( .A1(n1384), .A2(n1385), .ZN(n1382) );
NAND2_X1 U1104 ( .A1(n1386), .A2(G113), .ZN(n1385) );
XOR2_X1 U1105 ( .A(KEYINPUT25), .B(n1387), .Z(n1384) );
NOR2_X1 U1106 ( .A1(G113), .A2(n1386), .ZN(n1387) );
XNOR2_X1 U1107 ( .A(G116), .B(n1388), .ZN(n1386) );
NOR2_X1 U1108 ( .A1(G119), .A2(KEYINPUT35), .ZN(n1388) );
XNOR2_X1 U1109 ( .A(n1212), .B(KEYINPUT56), .ZN(n1183) );
XNOR2_X1 U1110 ( .A(G143), .B(n1347), .ZN(n1212) );
XNOR2_X1 U1111 ( .A(G128), .B(G146), .ZN(n1347) );
XNOR2_X1 U1112 ( .A(n1389), .B(n1189), .ZN(n1380) );
NAND2_X1 U1113 ( .A1(n1325), .A2(G210), .ZN(n1189) );
AND2_X1 U1114 ( .A1(n1390), .A2(n1125), .ZN(n1325) );
INV_X1 U1115 ( .A(G953), .ZN(n1125) );
XNOR2_X1 U1116 ( .A(KEYINPUT18), .B(n1368), .ZN(n1390) );
INV_X1 U1117 ( .A(G237), .ZN(n1368) );
XNOR2_X1 U1118 ( .A(G101), .B(KEYINPUT19), .ZN(n1389) );
NAND2_X1 U1119 ( .A1(KEYINPUT24), .A2(n1344), .ZN(n1291) );
INV_X1 U1120 ( .A(G110), .ZN(n1344) );
endmodule


