//Key = 0101110110011001011101010101100000010110001100011011010000010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347;

XNOR2_X1 U733 ( .A(G107), .B(n1011), .ZN(G9) );
NOR2_X1 U734 ( .A1(n1012), .A2(n1013), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1014), .A2(n1015), .A3(G953), .A4(n1016), .ZN(n1013) );
NOR3_X1 U736 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1015) );
XOR2_X1 U737 ( .A(n1020), .B(KEYINPUT2), .Z(n1018) );
NAND4_X1 U738 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1014) );
NAND4_X1 U739 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
INV_X1 U740 ( .A(KEYINPUT42), .ZN(n1026) );
NAND3_X1 U741 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1023) );
NAND2_X1 U742 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NAND3_X1 U743 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NAND2_X1 U744 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NAND2_X1 U745 ( .A1(n1039), .A2(n1040), .ZN(n1032) );
NAND3_X1 U746 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NAND2_X1 U747 ( .A1(n1034), .A2(n1044), .ZN(n1043) );
NAND2_X1 U748 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U749 ( .A1(KEYINPUT42), .A2(n1025), .ZN(n1046) );
NAND2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND3_X1 U751 ( .A1(n1049), .A2(n1050), .A3(n1036), .ZN(n1041) );
OR2_X1 U752 ( .A1(n1020), .A2(n1051), .ZN(n1022) );
NAND2_X1 U753 ( .A1(n1027), .A2(n1036), .ZN(n1020) );
AND3_X1 U754 ( .A1(n1034), .A2(n1039), .A3(n1029), .ZN(n1027) );
INV_X1 U755 ( .A(n1052), .ZN(n1029) );
NOR3_X1 U756 ( .A1(n1016), .A2(G953), .A3(G952), .ZN(n1012) );
AND4_X1 U757 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1016) );
NOR4_X1 U758 ( .A1(n1057), .A2(n1058), .A3(n1047), .A4(n1059), .ZN(n1056) );
XNOR2_X1 U759 ( .A(n1060), .B(n1061), .ZN(n1059) );
NAND2_X1 U760 ( .A1(KEYINPUT23), .A2(n1062), .ZN(n1060) );
NOR2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1057) );
XOR2_X1 U762 ( .A(n1065), .B(KEYINPUT7), .Z(n1063) );
NOR2_X1 U763 ( .A1(n1028), .A2(n1066), .ZN(n1055) );
XNOR2_X1 U764 ( .A(n1067), .B(n1068), .ZN(n1054) );
XOR2_X1 U765 ( .A(n1069), .B(n1070), .Z(n1053) );
NOR2_X1 U766 ( .A1(KEYINPUT39), .A2(n1071), .ZN(n1070) );
NAND3_X1 U767 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(G72) );
NAND2_X1 U768 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U769 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XNOR2_X1 U770 ( .A(n1079), .B(n1080), .ZN(n1075) );
NOR2_X1 U771 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
INV_X1 U772 ( .A(KEYINPUT43), .ZN(n1082) );
NAND2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(n1073) );
NAND2_X1 U774 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
OR4_X1 U775 ( .A1(n1081), .A2(n1087), .A3(n1088), .A4(KEYINPUT60), .ZN(n1086) );
INV_X1 U776 ( .A(n1079), .ZN(n1083) );
NAND4_X1 U777 ( .A1(n1085), .A2(n1077), .A3(n1089), .A4(n1079), .ZN(n1072) );
NAND2_X1 U778 ( .A1(G953), .A2(n1090), .ZN(n1079) );
NAND2_X1 U779 ( .A1(G900), .A2(G227), .ZN(n1090) );
NOR2_X1 U780 ( .A1(n1088), .A2(n1091), .ZN(n1089) );
NOR2_X1 U781 ( .A1(KEYINPUT60), .A2(n1081), .ZN(n1091) );
INV_X1 U782 ( .A(n1078), .ZN(n1088) );
NAND2_X1 U783 ( .A1(n1092), .A2(n1093), .ZN(n1078) );
XOR2_X1 U784 ( .A(n1094), .B(KEYINPUT14), .Z(n1092) );
INV_X1 U785 ( .A(n1087), .ZN(n1077) );
XOR2_X1 U786 ( .A(n1095), .B(KEYINPUT28), .Z(n1087) );
AND2_X1 U787 ( .A1(KEYINPUT43), .A2(n1096), .ZN(n1085) );
NAND2_X1 U788 ( .A1(KEYINPUT60), .A2(n1081), .ZN(n1096) );
NAND2_X1 U789 ( .A1(n1097), .A2(n1098), .ZN(n1081) );
NAND2_X1 U790 ( .A1(G953), .A2(n1099), .ZN(n1098) );
XNOR2_X1 U791 ( .A(n1100), .B(n1101), .ZN(n1097) );
XOR2_X1 U792 ( .A(n1102), .B(n1103), .Z(n1100) );
NAND3_X1 U793 ( .A1(n1104), .A2(n1105), .A3(KEYINPUT37), .ZN(n1102) );
NAND2_X1 U794 ( .A1(n1106), .A2(G131), .ZN(n1105) );
XNOR2_X1 U795 ( .A(n1107), .B(G137), .ZN(n1106) );
NAND2_X1 U796 ( .A1(n1108), .A2(n1109), .ZN(n1104) );
NAND3_X1 U797 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
INV_X1 U798 ( .A(n1113), .ZN(n1112) );
NAND2_X1 U799 ( .A1(G137), .A2(n1114), .ZN(n1111) );
NAND2_X1 U800 ( .A1(n1107), .A2(n1115), .ZN(n1110) );
NOR2_X1 U801 ( .A1(n1114), .A2(n1116), .ZN(n1107) );
INV_X1 U802 ( .A(KEYINPUT50), .ZN(n1114) );
XNOR2_X1 U803 ( .A(G131), .B(n1117), .ZN(n1108) );
XNOR2_X1 U804 ( .A(KEYINPUT31), .B(KEYINPUT21), .ZN(n1117) );
XOR2_X1 U805 ( .A(n1118), .B(n1119), .Z(G69) );
XOR2_X1 U806 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U807 ( .A1(G953), .A2(n1122), .ZN(n1121) );
NAND2_X1 U808 ( .A1(G898), .A2(G224), .ZN(n1122) );
NAND2_X1 U809 ( .A1(n1123), .A2(n1124), .ZN(n1120) );
NAND2_X1 U810 ( .A1(G953), .A2(n1125), .ZN(n1124) );
XOR2_X1 U811 ( .A(n1126), .B(n1127), .Z(n1123) );
NAND2_X1 U812 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
XOR2_X1 U813 ( .A(n1130), .B(KEYINPUT61), .Z(n1128) );
NOR2_X1 U814 ( .A1(n1131), .A2(G953), .ZN(n1118) );
NOR2_X1 U815 ( .A1(n1132), .A2(n1133), .ZN(G66) );
XNOR2_X1 U816 ( .A(n1134), .B(n1135), .ZN(n1133) );
NOR3_X1 U817 ( .A1(n1136), .A2(KEYINPUT0), .A3(n1137), .ZN(n1134) );
INV_X1 U818 ( .A(n1138), .ZN(n1136) );
NOR2_X1 U819 ( .A1(n1132), .A2(n1139), .ZN(G63) );
XOR2_X1 U820 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U821 ( .A1(n1138), .A2(G478), .ZN(n1141) );
NOR2_X1 U822 ( .A1(n1132), .A2(n1142), .ZN(G60) );
XOR2_X1 U823 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U824 ( .A1(KEYINPUT45), .A2(n1145), .ZN(n1144) );
XNOR2_X1 U825 ( .A(n1146), .B(n1147), .ZN(n1145) );
NAND3_X1 U826 ( .A1(n1148), .A2(n1149), .A3(G475), .ZN(n1143) );
XNOR2_X1 U827 ( .A(KEYINPUT13), .B(n1150), .ZN(n1148) );
XOR2_X1 U828 ( .A(G104), .B(n1151), .Z(G6) );
NOR2_X1 U829 ( .A1(n1132), .A2(n1152), .ZN(G57) );
XOR2_X1 U830 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U831 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U832 ( .A(n1157), .B(KEYINPUT18), .Z(n1156) );
NAND2_X1 U833 ( .A1(n1138), .A2(G472), .ZN(n1155) );
XOR2_X1 U834 ( .A(n1158), .B(n1159), .Z(n1153) );
NOR2_X1 U835 ( .A1(n1132), .A2(n1160), .ZN(G54) );
XNOR2_X1 U836 ( .A(n1161), .B(n1162), .ZN(n1160) );
XOR2_X1 U837 ( .A(n1163), .B(n1164), .Z(n1162) );
NAND3_X1 U838 ( .A1(n1138), .A2(G469), .A3(KEYINPUT12), .ZN(n1164) );
NAND4_X1 U839 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1163) );
NAND2_X1 U840 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
INV_X1 U841 ( .A(KEYINPUT47), .ZN(n1170) );
XNOR2_X1 U842 ( .A(n1171), .B(n1103), .ZN(n1169) );
NAND2_X1 U843 ( .A1(n1172), .A2(KEYINPUT47), .ZN(n1167) );
INV_X1 U844 ( .A(n1173), .ZN(n1166) );
NOR2_X1 U845 ( .A1(n1132), .A2(n1174), .ZN(G51) );
XOR2_X1 U846 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U847 ( .A1(KEYINPUT57), .A2(n1177), .ZN(n1176) );
XOR2_X1 U848 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U849 ( .A(n1180), .B(KEYINPUT35), .Z(n1178) );
NAND3_X1 U850 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
NAND2_X1 U851 ( .A1(n1101), .A2(n1184), .ZN(n1183) );
NAND2_X1 U852 ( .A1(KEYINPUT44), .A2(n1185), .ZN(n1182) );
NAND2_X1 U853 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
XNOR2_X1 U854 ( .A(KEYINPUT9), .B(n1101), .ZN(n1187) );
NAND2_X1 U855 ( .A1(n1188), .A2(n1189), .ZN(n1181) );
INV_X1 U856 ( .A(KEYINPUT44), .ZN(n1189) );
NAND2_X1 U857 ( .A1(n1190), .A2(n1191), .ZN(n1188) );
OR3_X1 U858 ( .A1(n1184), .A2(n1101), .A3(KEYINPUT9), .ZN(n1191) );
NAND2_X1 U859 ( .A1(KEYINPUT9), .A2(n1101), .ZN(n1190) );
NAND2_X1 U860 ( .A1(n1138), .A2(n1192), .ZN(n1175) );
NOR2_X1 U861 ( .A1(n1150), .A2(n1021), .ZN(n1138) );
INV_X1 U862 ( .A(n1149), .ZN(n1021) );
NAND3_X1 U863 ( .A1(n1093), .A2(n1094), .A3(n1131), .ZN(n1149) );
AND4_X1 U864 ( .A1(n1193), .A2(n1011), .A3(n1194), .A4(n1195), .ZN(n1131) );
NOR4_X1 U865 ( .A1(n1196), .A2(n1151), .A3(n1197), .A4(n1198), .ZN(n1195) );
NOR3_X1 U866 ( .A1(n1042), .A2(n1199), .A3(n1038), .ZN(n1197) );
AND3_X1 U867 ( .A1(n1034), .A2(n1200), .A3(n1201), .ZN(n1151) );
AND2_X1 U868 ( .A1(n1202), .A2(n1203), .ZN(n1194) );
NAND3_X1 U869 ( .A1(n1034), .A2(n1200), .A3(n1204), .ZN(n1011) );
NAND3_X1 U870 ( .A1(n1205), .A2(n1031), .A3(n1206), .ZN(n1094) );
XNOR2_X1 U871 ( .A(n1025), .B(KEYINPUT11), .ZN(n1206) );
AND4_X1 U872 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1093) );
AND3_X1 U873 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1210) );
NAND2_X1 U874 ( .A1(n1214), .A2(n1215), .ZN(n1209) );
NAND2_X1 U875 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
XOR2_X1 U876 ( .A(n1218), .B(KEYINPUT30), .Z(n1216) );
NOR2_X1 U877 ( .A1(n1095), .A2(G952), .ZN(n1132) );
XOR2_X1 U878 ( .A(G146), .B(n1219), .Z(G48) );
NOR2_X1 U879 ( .A1(n1051), .A2(n1218), .ZN(n1219) );
NAND3_X1 U880 ( .A1(n1201), .A2(n1050), .A3(n1220), .ZN(n1218) );
XOR2_X1 U881 ( .A(G143), .B(n1221), .Z(G45) );
NOR2_X1 U882 ( .A1(KEYINPUT40), .A2(n1207), .ZN(n1221) );
NAND4_X1 U883 ( .A1(n1222), .A2(n1223), .A3(n1214), .A4(n1066), .ZN(n1207) );
XOR2_X1 U884 ( .A(n1224), .B(n1225), .Z(G42) );
XOR2_X1 U885 ( .A(KEYINPUT52), .B(G140), .Z(n1225) );
NOR2_X1 U886 ( .A1(n1226), .A2(n1227), .ZN(n1224) );
NOR2_X1 U887 ( .A1(KEYINPUT49), .A2(n1228), .ZN(n1227) );
INV_X1 U888 ( .A(n1229), .ZN(n1228) );
NOR2_X1 U889 ( .A1(KEYINPUT63), .A2(n1229), .ZN(n1226) );
NAND3_X1 U890 ( .A1(n1031), .A2(n1025), .A3(n1205), .ZN(n1229) );
XOR2_X1 U891 ( .A(n1208), .B(n1230), .Z(G39) );
XNOR2_X1 U892 ( .A(KEYINPUT27), .B(n1115), .ZN(n1230) );
NAND4_X1 U893 ( .A1(n1220), .A2(n1031), .A3(n1039), .A4(n1050), .ZN(n1208) );
XNOR2_X1 U894 ( .A(G134), .B(n1211), .ZN(G36) );
NAND3_X1 U895 ( .A1(n1031), .A2(n1204), .A3(n1223), .ZN(n1211) );
XNOR2_X1 U896 ( .A(G131), .B(n1213), .ZN(G33) );
NAND3_X1 U897 ( .A1(n1201), .A2(n1031), .A3(n1223), .ZN(n1213) );
AND2_X1 U898 ( .A1(n1220), .A2(n1231), .ZN(n1223) );
INV_X1 U899 ( .A(n1028), .ZN(n1031) );
NAND2_X1 U900 ( .A1(n1232), .A2(n1017), .ZN(n1028) );
INV_X1 U901 ( .A(n1019), .ZN(n1232) );
XOR2_X1 U902 ( .A(n1233), .B(n1234), .Z(G30) );
NAND2_X1 U903 ( .A1(KEYINPUT4), .A2(G128), .ZN(n1234) );
NAND2_X1 U904 ( .A1(n1235), .A2(n1214), .ZN(n1233) );
XOR2_X1 U905 ( .A(n1217), .B(KEYINPUT51), .Z(n1235) );
NAND3_X1 U906 ( .A1(n1204), .A2(n1050), .A3(n1220), .ZN(n1217) );
AND3_X1 U907 ( .A1(n1025), .A2(n1236), .A3(n1237), .ZN(n1220) );
XOR2_X1 U908 ( .A(G101), .B(n1196), .Z(G3) );
AND4_X1 U909 ( .A1(n1237), .A2(n1200), .A3(n1231), .A4(n1039), .ZN(n1196) );
XNOR2_X1 U910 ( .A(G125), .B(n1212), .ZN(G27) );
NAND3_X1 U911 ( .A1(n1036), .A2(n1214), .A3(n1205), .ZN(n1212) );
AND4_X1 U912 ( .A1(n1201), .A2(n1049), .A3(n1050), .A4(n1236), .ZN(n1205) );
NAND2_X1 U913 ( .A1(n1052), .A2(n1238), .ZN(n1236) );
NAND2_X1 U914 ( .A1(n1239), .A2(n1099), .ZN(n1238) );
INV_X1 U915 ( .A(G900), .ZN(n1099) );
XNOR2_X1 U916 ( .A(G122), .B(n1203), .ZN(G24) );
NAND4_X1 U917 ( .A1(n1240), .A2(n1066), .A3(n1034), .A4(n1241), .ZN(n1203) );
NOR2_X1 U918 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NOR2_X1 U919 ( .A1(n1050), .A2(n1237), .ZN(n1034) );
XOR2_X1 U920 ( .A(n1244), .B(G119), .Z(G21) );
NAND2_X1 U921 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND2_X1 U922 ( .A1(n1198), .A2(n1247), .ZN(n1246) );
INV_X1 U923 ( .A(KEYINPUT20), .ZN(n1247) );
AND2_X1 U924 ( .A1(n1248), .A2(n1240), .ZN(n1198) );
NAND4_X1 U925 ( .A1(n1249), .A2(n1051), .A3(n1248), .A4(KEYINPUT20), .ZN(n1245) );
AND4_X1 U926 ( .A1(n1237), .A2(n1036), .A3(n1039), .A4(n1050), .ZN(n1248) );
XNOR2_X1 U927 ( .A(G116), .B(n1250), .ZN(G18) );
NOR2_X1 U928 ( .A1(KEYINPUT55), .A2(n1251), .ZN(n1250) );
NOR4_X1 U929 ( .A1(n1252), .A2(n1051), .A3(n1038), .A4(n1042), .ZN(n1251) );
INV_X1 U930 ( .A(n1204), .ZN(n1038) );
NOR2_X1 U931 ( .A1(n1222), .A2(n1253), .ZN(n1204) );
INV_X1 U932 ( .A(n1066), .ZN(n1253) );
XOR2_X1 U933 ( .A(n1249), .B(KEYINPUT59), .Z(n1252) );
XNOR2_X1 U934 ( .A(G113), .B(n1202), .ZN(G15) );
OR3_X1 U935 ( .A1(n1037), .A2(n1199), .A3(n1042), .ZN(n1202) );
NAND3_X1 U936 ( .A1(n1231), .A2(n1237), .A3(n1036), .ZN(n1042) );
INV_X1 U937 ( .A(n1242), .ZN(n1036) );
NAND2_X1 U938 ( .A1(n1048), .A2(n1254), .ZN(n1242) );
INV_X1 U939 ( .A(n1049), .ZN(n1237) );
INV_X1 U940 ( .A(n1050), .ZN(n1231) );
INV_X1 U941 ( .A(n1201), .ZN(n1037) );
XNOR2_X1 U942 ( .A(G110), .B(n1193), .ZN(G12) );
NAND4_X1 U943 ( .A1(n1200), .A2(n1039), .A3(n1049), .A4(n1050), .ZN(n1193) );
XOR2_X1 U944 ( .A(n1071), .B(n1069), .Z(n1050) );
NAND2_X1 U945 ( .A1(n1255), .A2(n1256), .ZN(n1069) );
XNOR2_X1 U946 ( .A(KEYINPUT16), .B(n1137), .ZN(n1255) );
INV_X1 U947 ( .A(G217), .ZN(n1137) );
NAND2_X1 U948 ( .A1(n1135), .A2(n1257), .ZN(n1071) );
XOR2_X1 U949 ( .A(n1258), .B(n1259), .Z(n1135) );
XNOR2_X1 U950 ( .A(n1260), .B(n1261), .ZN(n1259) );
XOR2_X1 U951 ( .A(KEYINPUT62), .B(G119), .Z(n1261) );
XOR2_X1 U952 ( .A(n1262), .B(n1263), .Z(n1258) );
XOR2_X1 U953 ( .A(n1264), .B(n1265), .Z(n1262) );
NOR2_X1 U954 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XOR2_X1 U955 ( .A(n1268), .B(n1269), .Z(n1267) );
NOR2_X1 U956 ( .A1(G137), .A2(KEYINPUT22), .ZN(n1269) );
AND3_X1 U957 ( .A1(G221), .A2(n1095), .A3(G234), .ZN(n1268) );
XNOR2_X1 U958 ( .A(KEYINPUT6), .B(KEYINPUT53), .ZN(n1266) );
NAND2_X1 U959 ( .A1(n1270), .A2(KEYINPUT5), .ZN(n1264) );
XNOR2_X1 U960 ( .A(G146), .B(n1271), .ZN(n1270) );
XOR2_X1 U961 ( .A(n1272), .B(n1067), .Z(n1049) );
NAND2_X1 U962 ( .A1(n1273), .A2(n1257), .ZN(n1067) );
XOR2_X1 U963 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U964 ( .A(KEYINPUT34), .B(G101), .Z(n1275) );
XNOR2_X1 U965 ( .A(n1276), .B(n1157), .ZN(n1274) );
NAND2_X1 U966 ( .A1(G210), .A2(n1277), .ZN(n1157) );
NAND2_X1 U967 ( .A1(n1278), .A2(n1279), .ZN(n1276) );
NAND2_X1 U968 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
XOR2_X1 U969 ( .A(n1159), .B(n1282), .Z(n1280) );
OR3_X1 U970 ( .A1(n1159), .A2(n1282), .A3(n1281), .ZN(n1278) );
INV_X1 U971 ( .A(KEYINPUT56), .ZN(n1281) );
XOR2_X1 U972 ( .A(n1283), .B(n1284), .Z(n1159) );
NOR2_X1 U973 ( .A1(KEYINPUT54), .A2(G116), .ZN(n1284) );
XNOR2_X1 U974 ( .A(G113), .B(G119), .ZN(n1283) );
NAND2_X1 U975 ( .A1(KEYINPUT15), .A2(n1068), .ZN(n1272) );
INV_X1 U976 ( .A(G472), .ZN(n1068) );
NAND2_X1 U977 ( .A1(n1285), .A2(n1286), .ZN(n1039) );
OR3_X1 U978 ( .A1(n1222), .A2(n1066), .A3(KEYINPUT58), .ZN(n1286) );
INV_X1 U979 ( .A(n1243), .ZN(n1222) );
NAND2_X1 U980 ( .A1(KEYINPUT58), .A2(n1201), .ZN(n1285) );
NOR2_X1 U981 ( .A1(n1243), .A2(n1066), .ZN(n1201) );
XNOR2_X1 U982 ( .A(n1287), .B(G478), .ZN(n1066) );
NAND2_X1 U983 ( .A1(n1257), .A2(n1140), .ZN(n1287) );
NAND2_X1 U984 ( .A1(n1288), .A2(n1289), .ZN(n1140) );
NAND2_X1 U985 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
XOR2_X1 U986 ( .A(n1292), .B(KEYINPUT29), .Z(n1288) );
OR2_X1 U987 ( .A1(n1291), .A2(n1290), .ZN(n1292) );
XOR2_X1 U988 ( .A(n1293), .B(n1294), .Z(n1290) );
XOR2_X1 U989 ( .A(n1263), .B(n1295), .Z(n1294) );
XNOR2_X1 U990 ( .A(n1296), .B(G107), .ZN(n1295) );
XNOR2_X1 U991 ( .A(G122), .B(n1297), .ZN(n1293) );
XNOR2_X1 U992 ( .A(G143), .B(n1116), .ZN(n1297) );
INV_X1 U993 ( .A(G134), .ZN(n1116) );
NAND3_X1 U994 ( .A1(G234), .A2(G217), .A3(n1298), .ZN(n1291) );
XNOR2_X1 U995 ( .A(G953), .B(KEYINPUT10), .ZN(n1298) );
XOR2_X1 U996 ( .A(n1299), .B(n1062), .Z(n1243) );
INV_X1 U997 ( .A(G475), .ZN(n1062) );
NAND2_X1 U998 ( .A1(KEYINPUT25), .A2(n1061), .ZN(n1299) );
NAND2_X1 U999 ( .A1(n1300), .A2(n1257), .ZN(n1061) );
XNOR2_X1 U1000 ( .A(n1146), .B(n1301), .ZN(n1300) );
INV_X1 U1001 ( .A(n1147), .ZN(n1301) );
XNOR2_X1 U1002 ( .A(n1302), .B(n1303), .ZN(n1147) );
XOR2_X1 U1003 ( .A(KEYINPUT38), .B(G131), .Z(n1303) );
XNOR2_X1 U1004 ( .A(G113), .B(G122), .ZN(n1302) );
XOR2_X1 U1005 ( .A(n1304), .B(n1305), .Z(n1146) );
XOR2_X1 U1006 ( .A(n1306), .B(n1271), .Z(n1305) );
XOR2_X1 U1007 ( .A(G125), .B(n1103), .Z(n1271) );
XOR2_X1 U1008 ( .A(n1307), .B(G104), .Z(n1304) );
NAND2_X1 U1009 ( .A1(G214), .A2(n1277), .ZN(n1307) );
NOR2_X1 U1010 ( .A1(G953), .A2(G237), .ZN(n1277) );
AND2_X1 U1011 ( .A1(n1240), .A2(n1025), .ZN(n1200) );
NOR2_X1 U1012 ( .A1(n1048), .A2(n1047), .ZN(n1025) );
INV_X1 U1013 ( .A(n1254), .ZN(n1047) );
NAND2_X1 U1014 ( .A1(n1308), .A2(n1256), .ZN(n1254) );
NAND2_X1 U1015 ( .A1(G234), .A2(n1150), .ZN(n1256) );
XNOR2_X1 U1016 ( .A(G221), .B(KEYINPUT19), .ZN(n1308) );
NOR2_X1 U1017 ( .A1(n1309), .A2(n1058), .ZN(n1048) );
NOR2_X1 U1018 ( .A1(n1065), .A2(G469), .ZN(n1058) );
AND2_X1 U1019 ( .A1(n1310), .A2(n1065), .ZN(n1309) );
NAND2_X1 U1020 ( .A1(n1311), .A2(n1257), .ZN(n1065) );
XNOR2_X1 U1021 ( .A(n1312), .B(n1313), .ZN(n1311) );
INV_X1 U1022 ( .A(n1161), .ZN(n1313) );
XNOR2_X1 U1023 ( .A(n1314), .B(n1158), .ZN(n1161) );
XOR2_X1 U1024 ( .A(G101), .B(n1282), .Z(n1158) );
XOR2_X1 U1025 ( .A(n1315), .B(n1316), .Z(n1282) );
XOR2_X1 U1026 ( .A(G131), .B(n1317), .Z(n1316) );
NOR2_X1 U1027 ( .A1(n1113), .A2(n1318), .ZN(n1317) );
XOR2_X1 U1028 ( .A(n1319), .B(KEYINPUT17), .Z(n1318) );
NAND2_X1 U1029 ( .A1(G134), .A2(n1320), .ZN(n1319) );
XNOR2_X1 U1030 ( .A(KEYINPUT48), .B(n1115), .ZN(n1320) );
NOR2_X1 U1031 ( .A1(n1115), .A2(G134), .ZN(n1113) );
INV_X1 U1032 ( .A(G137), .ZN(n1115) );
XNOR2_X1 U1033 ( .A(G107), .B(n1321), .ZN(n1314) );
NOR2_X1 U1034 ( .A1(G104), .A2(KEYINPUT32), .ZN(n1321) );
NOR3_X1 U1035 ( .A1(n1172), .A2(n1173), .A3(n1322), .ZN(n1312) );
INV_X1 U1036 ( .A(n1165), .ZN(n1322) );
NAND3_X1 U1037 ( .A1(G110), .A2(n1103), .A3(n1171), .ZN(n1165) );
NOR3_X1 U1038 ( .A1(n1103), .A2(n1171), .A3(n1260), .ZN(n1173) );
INV_X1 U1039 ( .A(n1323), .ZN(n1171) );
AND2_X1 U1040 ( .A1(n1324), .A2(n1260), .ZN(n1172) );
XNOR2_X1 U1041 ( .A(n1323), .B(n1103), .ZN(n1324) );
XOR2_X1 U1042 ( .A(G140), .B(KEYINPUT33), .Z(n1103) );
NAND2_X1 U1043 ( .A1(G227), .A2(n1095), .ZN(n1323) );
XNOR2_X1 U1044 ( .A(KEYINPUT24), .B(n1064), .ZN(n1310) );
INV_X1 U1045 ( .A(G469), .ZN(n1064) );
INV_X1 U1046 ( .A(n1199), .ZN(n1240) );
NAND2_X1 U1047 ( .A1(n1214), .A2(n1249), .ZN(n1199) );
NAND2_X1 U1048 ( .A1(n1052), .A2(n1325), .ZN(n1249) );
NAND2_X1 U1049 ( .A1(n1239), .A2(n1125), .ZN(n1325) );
INV_X1 U1050 ( .A(G898), .ZN(n1125) );
AND3_X1 U1051 ( .A1(n1326), .A2(n1327), .A3(G953), .ZN(n1239) );
XNOR2_X1 U1052 ( .A(KEYINPUT26), .B(n1150), .ZN(n1326) );
NAND3_X1 U1053 ( .A1(n1327), .A2(n1095), .A3(G952), .ZN(n1052) );
NAND2_X1 U1054 ( .A1(G237), .A2(G234), .ZN(n1327) );
INV_X1 U1055 ( .A(n1051), .ZN(n1214) );
NAND2_X1 U1056 ( .A1(n1019), .A2(n1017), .ZN(n1051) );
NAND2_X1 U1057 ( .A1(G214), .A2(n1328), .ZN(n1017) );
XNOR2_X1 U1058 ( .A(n1329), .B(n1192), .ZN(n1019) );
AND2_X1 U1059 ( .A1(G210), .A2(n1328), .ZN(n1192) );
NAND2_X1 U1060 ( .A1(n1330), .A2(n1150), .ZN(n1328) );
INV_X1 U1061 ( .A(G237), .ZN(n1330) );
NAND2_X1 U1062 ( .A1(n1331), .A2(n1257), .ZN(n1329) );
XNOR2_X1 U1063 ( .A(n1150), .B(KEYINPUT3), .ZN(n1257) );
INV_X1 U1064 ( .A(G902), .ZN(n1150) );
XOR2_X1 U1065 ( .A(n1332), .B(n1333), .Z(n1331) );
XNOR2_X1 U1066 ( .A(n1179), .B(n1101), .ZN(n1333) );
XNOR2_X1 U1067 ( .A(G125), .B(n1315), .ZN(n1101) );
XOR2_X1 U1068 ( .A(n1306), .B(n1263), .Z(n1315) );
XOR2_X1 U1069 ( .A(G128), .B(KEYINPUT1), .Z(n1263) );
XOR2_X1 U1070 ( .A(G143), .B(G146), .Z(n1306) );
XNOR2_X1 U1071 ( .A(n1334), .B(n1127), .ZN(n1179) );
XNOR2_X1 U1072 ( .A(G122), .B(n1260), .ZN(n1127) );
INV_X1 U1073 ( .A(G110), .ZN(n1260) );
NAND2_X1 U1074 ( .A1(n1335), .A2(n1129), .ZN(n1334) );
NAND3_X1 U1075 ( .A1(n1336), .A2(n1337), .A3(n1338), .ZN(n1129) );
XOR2_X1 U1076 ( .A(n1130), .B(KEYINPUT46), .Z(n1335) );
NAND2_X1 U1077 ( .A1(n1339), .A2(n1340), .ZN(n1130) );
NAND2_X1 U1078 ( .A1(n1336), .A2(n1337), .ZN(n1340) );
NAND2_X1 U1079 ( .A1(n1341), .A2(n1342), .ZN(n1337) );
XNOR2_X1 U1080 ( .A(KEYINPUT36), .B(n1343), .ZN(n1342) );
INV_X1 U1081 ( .A(G113), .ZN(n1343) );
XNOR2_X1 U1082 ( .A(G119), .B(n1296), .ZN(n1341) );
INV_X1 U1083 ( .A(G116), .ZN(n1296) );
XNOR2_X1 U1084 ( .A(KEYINPUT8), .B(n1344), .ZN(n1336) );
NAND2_X1 U1085 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
XNOR2_X1 U1086 ( .A(KEYINPUT36), .B(G113), .ZN(n1346) );
XNOR2_X1 U1087 ( .A(G116), .B(G119), .ZN(n1345) );
INV_X1 U1088 ( .A(n1338), .ZN(n1339) );
XOR2_X1 U1089 ( .A(G101), .B(n1347), .Z(n1338) );
XOR2_X1 U1090 ( .A(G107), .B(G104), .Z(n1347) );
XNOR2_X1 U1091 ( .A(n1186), .B(KEYINPUT41), .ZN(n1332) );
INV_X1 U1092 ( .A(n1184), .ZN(n1186) );
NAND2_X1 U1093 ( .A1(G224), .A2(n1095), .ZN(n1184) );
INV_X1 U1094 ( .A(G953), .ZN(n1095) );
endmodule


