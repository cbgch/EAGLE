//Key = 1100010111111011010101101111000010111100111011010011110111011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366;

XOR2_X1 U753 ( .A(n1033), .B(n1034), .Z(G9) );
XOR2_X1 U754 ( .A(KEYINPUT23), .B(G107), .Z(n1034) );
NOR2_X1 U755 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U756 ( .A1(n1037), .A2(n1038), .ZN(G75) );
NOR2_X1 U757 ( .A1(G952), .A2(n1039), .ZN(n1038) );
NOR4_X1 U758 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1037) );
NAND3_X1 U759 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1040) );
INV_X1 U760 ( .A(n1039), .ZN(n1046) );
NAND2_X1 U761 ( .A1(n1047), .A2(n1048), .ZN(n1039) );
NAND4_X1 U762 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
NOR3_X1 U763 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
INV_X1 U764 ( .A(n1056), .ZN(n1054) );
XOR2_X1 U765 ( .A(KEYINPUT37), .B(n1057), .Z(n1053) );
NOR2_X1 U766 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U767 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
INV_X1 U768 ( .A(G478), .ZN(n1061) );
NOR2_X1 U769 ( .A1(G902), .A2(n1062), .ZN(n1060) );
NAND3_X1 U770 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1045) );
NAND2_X1 U771 ( .A1(n1066), .A2(n1036), .ZN(n1064) );
XOR2_X1 U772 ( .A(KEYINPUT59), .B(n1067), .Z(n1066) );
NOR2_X1 U773 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U774 ( .A1(n1070), .A2(n1071), .ZN(n1044) );
NAND3_X1 U775 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
NAND2_X1 U776 ( .A1(KEYINPUT18), .A2(n1075), .ZN(n1074) );
NAND2_X1 U777 ( .A1(n1065), .A2(n1076), .ZN(n1075) );
AND3_X1 U778 ( .A1(n1077), .A2(n1056), .A3(n1078), .ZN(n1065) );
NAND4_X1 U779 ( .A1(n1077), .A2(n1056), .A3(n1079), .A4(n1080), .ZN(n1073) );
NAND2_X1 U780 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
OR2_X1 U781 ( .A1(n1083), .A2(KEYINPUT11), .ZN(n1081) );
NAND3_X1 U782 ( .A1(n1084), .A2(n1085), .A3(n1078), .ZN(n1079) );
NAND2_X1 U783 ( .A1(KEYINPUT11), .A2(n1086), .ZN(n1085) );
OR2_X1 U784 ( .A1(n1087), .A2(KEYINPUT18), .ZN(n1084) );
NAND3_X1 U785 ( .A1(n1063), .A2(n1088), .A3(n1078), .ZN(n1072) );
INV_X1 U786 ( .A(n1082), .ZN(n1078) );
NAND2_X1 U787 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U788 ( .A1(n1056), .A2(n1091), .ZN(n1090) );
NAND2_X1 U789 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U790 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U791 ( .A1(n1077), .A2(n1096), .ZN(n1089) );
NAND2_X1 U792 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U793 ( .A(n1099), .B(n1100), .Z(G72) );
NOR2_X1 U794 ( .A1(n1101), .A2(n1047), .ZN(n1100) );
XOR2_X1 U795 ( .A(n1102), .B(KEYINPUT17), .Z(n1101) );
NAND2_X1 U796 ( .A1(G900), .A2(G227), .ZN(n1102) );
NAND2_X1 U797 ( .A1(n1103), .A2(n1104), .ZN(n1099) );
NAND2_X1 U798 ( .A1(n1105), .A2(n1047), .ZN(n1104) );
XOR2_X1 U799 ( .A(n1041), .B(n1106), .Z(n1105) );
NAND3_X1 U800 ( .A1(n1106), .A2(G900), .A3(G953), .ZN(n1103) );
AND2_X1 U801 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U802 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U803 ( .A(KEYINPUT52), .B(n1111), .Z(n1107) );
NOR2_X1 U804 ( .A1(n1109), .A2(n1110), .ZN(n1111) );
XOR2_X1 U805 ( .A(n1112), .B(n1113), .Z(n1110) );
XOR2_X1 U806 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U807 ( .A1(n1116), .A2(n1117), .ZN(n1112) );
NAND2_X1 U808 ( .A1(KEYINPUT9), .A2(n1118), .ZN(n1117) );
OR3_X1 U809 ( .A1(n1119), .A2(G137), .A3(KEYINPUT9), .ZN(n1116) );
AND2_X1 U810 ( .A1(n1120), .A2(n1121), .ZN(n1109) );
OR2_X1 U811 ( .A1(n1122), .A2(G125), .ZN(n1121) );
NAND2_X1 U812 ( .A1(n1123), .A2(n1122), .ZN(n1120) );
XOR2_X1 U813 ( .A(KEYINPUT38), .B(G125), .Z(n1123) );
XOR2_X1 U814 ( .A(n1124), .B(n1125), .Z(G69) );
NOR2_X1 U815 ( .A1(n1126), .A2(n1047), .ZN(n1125) );
AND2_X1 U816 ( .A1(G224), .A2(G898), .ZN(n1126) );
NAND2_X1 U817 ( .A1(n1127), .A2(n1128), .ZN(n1124) );
NAND2_X1 U818 ( .A1(n1129), .A2(n1047), .ZN(n1128) );
XOR2_X1 U819 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U820 ( .A1(n1132), .A2(n1133), .ZN(n1130) );
INV_X1 U821 ( .A(n1043), .ZN(n1133) );
XOR2_X1 U822 ( .A(n1042), .B(KEYINPUT8), .Z(n1132) );
NAND3_X1 U823 ( .A1(G898), .A2(n1131), .A3(G953), .ZN(n1127) );
NOR2_X1 U824 ( .A1(n1134), .A2(n1135), .ZN(G66) );
XNOR2_X1 U825 ( .A(n1136), .B(n1137), .ZN(n1135) );
XOR2_X1 U826 ( .A(n1138), .B(KEYINPUT4), .Z(n1136) );
NAND2_X1 U827 ( .A1(n1139), .A2(G217), .ZN(n1138) );
NOR2_X1 U828 ( .A1(n1134), .A2(n1140), .ZN(G63) );
XOR2_X1 U829 ( .A(n1141), .B(n1062), .Z(n1140) );
XOR2_X1 U830 ( .A(n1142), .B(KEYINPUT47), .Z(n1141) );
NAND2_X1 U831 ( .A1(n1139), .A2(G478), .ZN(n1142) );
NOR2_X1 U832 ( .A1(n1134), .A2(n1143), .ZN(G60) );
XOR2_X1 U833 ( .A(n1144), .B(n1145), .Z(n1143) );
NAND3_X1 U834 ( .A1(n1139), .A2(G475), .A3(n1146), .ZN(n1145) );
XNOR2_X1 U835 ( .A(KEYINPUT61), .B(KEYINPUT20), .ZN(n1146) );
NAND3_X1 U836 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(G6) );
NAND2_X1 U837 ( .A1(G104), .A2(n1150), .ZN(n1149) );
NAND2_X1 U838 ( .A1(n1151), .A2(KEYINPUT32), .ZN(n1150) );
XOR2_X1 U839 ( .A(n1152), .B(KEYINPUT35), .Z(n1151) );
NAND3_X1 U840 ( .A1(KEYINPUT32), .A2(n1153), .A3(n1154), .ZN(n1148) );
OR2_X1 U841 ( .A1(n1154), .A2(KEYINPUT32), .ZN(n1147) );
INV_X1 U842 ( .A(n1152), .ZN(n1154) );
NOR2_X1 U843 ( .A1(n1134), .A2(n1155), .ZN(G57) );
XOR2_X1 U844 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U845 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR3_X1 U846 ( .A1(n1160), .A2(KEYINPUT49), .A3(n1161), .ZN(n1158) );
INV_X1 U847 ( .A(G472), .ZN(n1161) );
XNOR2_X1 U848 ( .A(n1162), .B(n1163), .ZN(n1156) );
NOR2_X1 U849 ( .A1(n1134), .A2(n1164), .ZN(G54) );
XOR2_X1 U850 ( .A(n1165), .B(n1166), .Z(n1164) );
XNOR2_X1 U851 ( .A(n1167), .B(n1168), .ZN(n1166) );
XNOR2_X1 U852 ( .A(n1169), .B(n1170), .ZN(n1168) );
NAND2_X1 U853 ( .A1(n1139), .A2(G469), .ZN(n1169) );
XOR2_X1 U854 ( .A(n1171), .B(n1172), .Z(n1165) );
XOR2_X1 U855 ( .A(G140), .B(G110), .Z(n1172) );
NOR2_X1 U856 ( .A1(KEYINPUT30), .A2(n1173), .ZN(n1171) );
NOR2_X1 U857 ( .A1(n1134), .A2(n1174), .ZN(G51) );
XOR2_X1 U858 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U859 ( .A(n1177), .B(n1131), .Z(n1176) );
NAND2_X1 U860 ( .A1(n1139), .A2(n1178), .ZN(n1177) );
INV_X1 U861 ( .A(n1160), .ZN(n1139) );
NAND2_X1 U862 ( .A1(G902), .A2(n1179), .ZN(n1160) );
OR3_X1 U863 ( .A1(n1043), .A2(n1042), .A3(n1041), .ZN(n1179) );
NAND4_X1 U864 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1041) );
AND4_X1 U865 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1183) );
NOR3_X1 U866 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1182) );
NOR3_X1 U867 ( .A1(n1191), .A2(n1192), .A3(n1036), .ZN(n1190) );
INV_X1 U868 ( .A(KEYINPUT63), .ZN(n1191) );
NOR2_X1 U869 ( .A1(KEYINPUT63), .A2(n1193), .ZN(n1189) );
NOR3_X1 U870 ( .A1(n1194), .A2(n1083), .A3(n1195), .ZN(n1188) );
XOR2_X1 U871 ( .A(KEYINPUT57), .B(n1196), .Z(n1194) );
NAND4_X1 U872 ( .A1(n1197), .A2(n1198), .A3(n1070), .A4(n1199), .ZN(n1180) );
NOR2_X1 U873 ( .A1(n1087), .A2(n1098), .ZN(n1199) );
OR2_X1 U874 ( .A1(n1200), .A2(KEYINPUT29), .ZN(n1198) );
NAND2_X1 U875 ( .A1(KEYINPUT29), .A2(n1201), .ZN(n1197) );
NAND2_X1 U876 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NAND4_X1 U877 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1152), .ZN(n1042) );
NAND3_X1 U878 ( .A1(n1076), .A2(n1056), .A3(n1207), .ZN(n1152) );
NAND3_X1 U879 ( .A1(n1063), .A2(n1208), .A3(n1207), .ZN(n1205) );
NAND2_X1 U880 ( .A1(n1209), .A2(n1196), .ZN(n1204) );
XOR2_X1 U881 ( .A(n1035), .B(KEYINPUT41), .Z(n1209) );
NAND4_X1 U882 ( .A1(n1203), .A2(n1056), .A3(n1086), .A4(n1210), .ZN(n1035) );
NAND4_X1 U883 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1043) );
XOR2_X1 U884 ( .A(n1215), .B(KEYINPUT44), .Z(n1175) );
NAND3_X1 U885 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
OR2_X1 U886 ( .A1(n1219), .A2(KEYINPUT36), .ZN(n1217) );
NAND3_X1 U887 ( .A1(n1219), .A2(n1220), .A3(KEYINPUT36), .ZN(n1216) );
NOR2_X1 U888 ( .A1(n1047), .A2(G952), .ZN(n1134) );
XOR2_X1 U889 ( .A(n1193), .B(n1221), .Z(G48) );
NAND2_X1 U890 ( .A1(KEYINPUT1), .A2(G146), .ZN(n1221) );
NAND2_X1 U891 ( .A1(n1192), .A2(n1196), .ZN(n1193) );
NOR2_X1 U892 ( .A1(n1195), .A2(n1087), .ZN(n1192) );
XNOR2_X1 U893 ( .A(G143), .B(n1181), .ZN(G45) );
NAND3_X1 U894 ( .A1(n1200), .A2(n1222), .A3(n1223), .ZN(n1181) );
NOR3_X1 U895 ( .A1(n1036), .A2(n1224), .A3(n1225), .ZN(n1223) );
NAND2_X1 U896 ( .A1(n1226), .A2(n1227), .ZN(G42) );
NAND2_X1 U897 ( .A1(n1228), .A2(n1122), .ZN(n1227) );
NAND2_X1 U898 ( .A1(n1229), .A2(G140), .ZN(n1226) );
NAND2_X1 U899 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND2_X1 U900 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
OR2_X1 U901 ( .A1(n1233), .A2(n1228), .ZN(n1230) );
NOR2_X1 U902 ( .A1(KEYINPUT2), .A2(n1187), .ZN(n1228) );
INV_X1 U903 ( .A(n1232), .ZN(n1187) );
NOR2_X1 U904 ( .A1(n1234), .A2(n1097), .ZN(n1232) );
INV_X1 U905 ( .A(KEYINPUT14), .ZN(n1233) );
XNOR2_X1 U906 ( .A(n1186), .B(n1235), .ZN(G39) );
XOR2_X1 U907 ( .A(KEYINPUT16), .B(G137), .Z(n1235) );
OR3_X1 U908 ( .A1(n1236), .A2(n1055), .A3(n1195), .ZN(n1186) );
XOR2_X1 U909 ( .A(n1185), .B(n1237), .Z(G36) );
XOR2_X1 U910 ( .A(KEYINPUT15), .B(G134), .Z(n1237) );
NAND4_X1 U911 ( .A1(n1200), .A2(n1070), .A3(n1222), .A4(n1086), .ZN(n1185) );
XOR2_X1 U912 ( .A(G131), .B(n1238), .Z(G33) );
NOR2_X1 U913 ( .A1(n1098), .A2(n1234), .ZN(n1238) );
NAND3_X1 U914 ( .A1(n1070), .A2(n1076), .A3(n1200), .ZN(n1234) );
INV_X1 U915 ( .A(n1055), .ZN(n1070) );
NAND2_X1 U916 ( .A1(n1239), .A2(n1069), .ZN(n1055) );
XOR2_X1 U917 ( .A(G128), .B(n1240), .Z(G30) );
NOR3_X1 U918 ( .A1(n1195), .A2(n1241), .A3(n1036), .ZN(n1240) );
XOR2_X1 U919 ( .A(n1083), .B(KEYINPUT46), .Z(n1241) );
NAND3_X1 U920 ( .A1(n1200), .A2(n1242), .A3(n1243), .ZN(n1195) );
NOR2_X1 U921 ( .A1(n1092), .A2(n1202), .ZN(n1200) );
INV_X1 U922 ( .A(n1203), .ZN(n1092) );
XOR2_X1 U923 ( .A(n1206), .B(n1244), .Z(G3) );
NAND2_X1 U924 ( .A1(KEYINPUT24), .A2(G101), .ZN(n1244) );
NAND3_X1 U925 ( .A1(n1063), .A2(n1222), .A3(n1207), .ZN(n1206) );
INV_X1 U926 ( .A(n1245), .ZN(n1207) );
XNOR2_X1 U927 ( .A(G125), .B(n1184), .ZN(G27) );
NAND4_X1 U928 ( .A1(n1208), .A2(n1076), .A3(n1246), .A4(n1077), .ZN(n1184) );
NOR2_X1 U929 ( .A1(n1202), .A2(n1036), .ZN(n1246) );
AND2_X1 U930 ( .A1(n1247), .A2(n1082), .ZN(n1202) );
NAND4_X1 U931 ( .A1(G953), .A2(G902), .A3(n1248), .A4(n1249), .ZN(n1247) );
INV_X1 U932 ( .A(G900), .ZN(n1249) );
XOR2_X1 U933 ( .A(n1250), .B(G122), .Z(G24) );
NAND2_X1 U934 ( .A1(KEYINPUT22), .A2(n1214), .ZN(n1250) );
NAND4_X1 U935 ( .A1(n1251), .A2(n1056), .A3(n1252), .A4(n1253), .ZN(n1214) );
NOR2_X1 U936 ( .A1(n1254), .A2(n1242), .ZN(n1056) );
XOR2_X1 U937 ( .A(n1255), .B(n1256), .Z(G21) );
NAND2_X1 U938 ( .A1(KEYINPUT0), .A2(n1257), .ZN(n1256) );
INV_X1 U939 ( .A(n1211), .ZN(n1257) );
NAND4_X1 U940 ( .A1(n1251), .A2(n1063), .A3(n1243), .A4(n1242), .ZN(n1211) );
XOR2_X1 U941 ( .A(n1254), .B(KEYINPUT54), .Z(n1243) );
NAND2_X1 U942 ( .A1(n1258), .A2(n1259), .ZN(G18) );
NAND2_X1 U943 ( .A1(G116), .A2(n1212), .ZN(n1259) );
XOR2_X1 U944 ( .A(n1260), .B(KEYINPUT6), .Z(n1258) );
OR2_X1 U945 ( .A1(n1212), .A2(G116), .ZN(n1260) );
NAND3_X1 U946 ( .A1(n1222), .A2(n1086), .A3(n1251), .ZN(n1212) );
INV_X1 U947 ( .A(n1083), .ZN(n1086) );
NAND2_X1 U948 ( .A1(n1051), .A2(n1253), .ZN(n1083) );
XNOR2_X1 U949 ( .A(G113), .B(n1213), .ZN(G15) );
NAND3_X1 U950 ( .A1(n1222), .A2(n1076), .A3(n1251), .ZN(n1213) );
AND3_X1 U951 ( .A1(n1196), .A2(n1210), .A3(n1077), .ZN(n1251) );
AND2_X1 U952 ( .A1(n1095), .A2(n1050), .ZN(n1077) );
INV_X1 U953 ( .A(n1087), .ZN(n1076) );
NAND2_X1 U954 ( .A1(n1224), .A2(n1252), .ZN(n1087) );
INV_X1 U955 ( .A(n1225), .ZN(n1252) );
XOR2_X1 U956 ( .A(n1051), .B(KEYINPUT33), .Z(n1225) );
INV_X1 U957 ( .A(n1098), .ZN(n1222) );
NAND2_X1 U958 ( .A1(n1261), .A2(n1242), .ZN(n1098) );
XOR2_X1 U959 ( .A(G110), .B(n1262), .Z(G12) );
NOR3_X1 U960 ( .A1(n1263), .A2(n1097), .A3(n1245), .ZN(n1262) );
NAND3_X1 U961 ( .A1(n1203), .A2(n1210), .A3(n1196), .ZN(n1245) );
INV_X1 U962 ( .A(n1036), .ZN(n1196) );
NAND2_X1 U963 ( .A1(n1264), .A2(n1069), .ZN(n1036) );
NAND2_X1 U964 ( .A1(G214), .A2(n1265), .ZN(n1069) );
XOR2_X1 U965 ( .A(KEYINPUT58), .B(n1068), .Z(n1264) );
INV_X1 U966 ( .A(n1239), .ZN(n1068) );
XOR2_X1 U967 ( .A(n1266), .B(n1178), .Z(n1239) );
AND2_X1 U968 ( .A1(G210), .A2(n1265), .ZN(n1178) );
NAND2_X1 U969 ( .A1(n1267), .A2(n1268), .ZN(n1265) );
INV_X1 U970 ( .A(G237), .ZN(n1267) );
NAND2_X1 U971 ( .A1(n1269), .A2(n1268), .ZN(n1266) );
XOR2_X1 U972 ( .A(n1131), .B(n1270), .Z(n1269) );
XOR2_X1 U973 ( .A(n1271), .B(KEYINPUT19), .Z(n1270) );
NAND2_X1 U974 ( .A1(n1218), .A2(n1272), .ZN(n1271) );
NAND2_X1 U975 ( .A1(n1219), .A2(n1220), .ZN(n1272) );
OR2_X1 U976 ( .A1(n1220), .A2(n1219), .ZN(n1218) );
XOR2_X1 U977 ( .A(G125), .B(n1273), .Z(n1219) );
NAND2_X1 U978 ( .A1(G224), .A2(n1047), .ZN(n1220) );
XOR2_X1 U979 ( .A(n1274), .B(n1275), .Z(n1131) );
XOR2_X1 U980 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U981 ( .A(n1278), .B(n1279), .Z(n1274) );
NOR2_X1 U982 ( .A1(KEYINPUT3), .A2(n1280), .ZN(n1279) );
INV_X1 U983 ( .A(n1281), .ZN(n1280) );
XNOR2_X1 U984 ( .A(G101), .B(G122), .ZN(n1278) );
NAND2_X1 U985 ( .A1(n1082), .A2(n1282), .ZN(n1210) );
NAND4_X1 U986 ( .A1(G953), .A2(G902), .A3(n1248), .A4(n1283), .ZN(n1282) );
INV_X1 U987 ( .A(G898), .ZN(n1283) );
NAND3_X1 U988 ( .A1(n1248), .A2(n1047), .A3(G952), .ZN(n1082) );
NAND2_X1 U989 ( .A1(G237), .A2(G234), .ZN(n1248) );
NOR2_X1 U990 ( .A1(n1095), .A2(n1094), .ZN(n1203) );
INV_X1 U991 ( .A(n1050), .ZN(n1094) );
NAND2_X1 U992 ( .A1(n1284), .A2(n1285), .ZN(n1050) );
NAND2_X1 U993 ( .A1(G234), .A2(n1268), .ZN(n1285) );
XOR2_X1 U994 ( .A(KEYINPUT39), .B(G221), .Z(n1284) );
XNOR2_X1 U995 ( .A(n1049), .B(KEYINPUT51), .ZN(n1095) );
XOR2_X1 U996 ( .A(n1286), .B(G469), .Z(n1049) );
NAND2_X1 U997 ( .A1(n1287), .A2(n1268), .ZN(n1286) );
XOR2_X1 U998 ( .A(n1170), .B(n1288), .Z(n1287) );
XOR2_X1 U999 ( .A(n1289), .B(n1290), .Z(n1288) );
NOR2_X1 U1000 ( .A1(KEYINPUT13), .A2(n1167), .ZN(n1290) );
XOR2_X1 U1001 ( .A(n1115), .B(n1291), .Z(n1167) );
NOR2_X1 U1002 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XOR2_X1 U1003 ( .A(n1294), .B(KEYINPUT12), .Z(n1293) );
NAND2_X1 U1004 ( .A1(G101), .A2(n1281), .ZN(n1294) );
NOR2_X1 U1005 ( .A1(G101), .A2(n1281), .ZN(n1292) );
XOR2_X1 U1006 ( .A(G107), .B(G104), .Z(n1281) );
XOR2_X1 U1007 ( .A(n1295), .B(KEYINPUT45), .Z(n1115) );
NAND3_X1 U1008 ( .A1(n1296), .A2(n1297), .A3(n1298), .ZN(n1295) );
NAND2_X1 U1009 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
NAND2_X1 U1010 ( .A1(KEYINPUT7), .A2(n1301), .ZN(n1300) );
XOR2_X1 U1011 ( .A(KEYINPUT10), .B(G128), .Z(n1301) );
NAND3_X1 U1012 ( .A1(KEYINPUT7), .A2(n1302), .A3(n1303), .ZN(n1297) );
INV_X1 U1013 ( .A(n1299), .ZN(n1302) );
OR2_X1 U1014 ( .A1(n1303), .A2(KEYINPUT7), .ZN(n1296) );
INV_X1 U1015 ( .A(G128), .ZN(n1303) );
NOR2_X1 U1016 ( .A1(n1304), .A2(n1305), .ZN(n1289) );
XOR2_X1 U1017 ( .A(KEYINPUT62), .B(n1306), .Z(n1305) );
NOR2_X1 U1018 ( .A1(n1173), .A2(n1307), .ZN(n1306) );
AND2_X1 U1019 ( .A1(n1307), .A2(n1173), .ZN(n1304) );
NAND2_X1 U1020 ( .A1(G227), .A2(n1047), .ZN(n1173) );
NAND2_X1 U1021 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND2_X1 U1022 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
XOR2_X1 U1023 ( .A(KEYINPUT34), .B(n1312), .Z(n1308) );
NOR2_X1 U1024 ( .A1(n1310), .A2(n1311), .ZN(n1312) );
XOR2_X1 U1025 ( .A(KEYINPUT26), .B(n1122), .Z(n1310) );
INV_X1 U1026 ( .A(G140), .ZN(n1122) );
INV_X1 U1027 ( .A(n1208), .ZN(n1097) );
NOR2_X1 U1028 ( .A1(n1242), .A2(n1261), .ZN(n1208) );
INV_X1 U1029 ( .A(n1254), .ZN(n1261) );
NAND3_X1 U1030 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1254) );
NAND2_X1 U1031 ( .A1(n1316), .A2(n1137), .ZN(n1315) );
OR3_X1 U1032 ( .A1(n1137), .A2(n1316), .A3(G902), .ZN(n1314) );
NOR2_X1 U1033 ( .A1(n1317), .A2(G234), .ZN(n1316) );
INV_X1 U1034 ( .A(G217), .ZN(n1317) );
XOR2_X1 U1035 ( .A(n1318), .B(n1319), .Z(n1137) );
XNOR2_X1 U1036 ( .A(n1277), .B(n1320), .ZN(n1319) );
XNOR2_X1 U1037 ( .A(n1321), .B(n1322), .ZN(n1320) );
XOR2_X1 U1038 ( .A(n1255), .B(n1311), .Z(n1277) );
INV_X1 U1039 ( .A(G110), .ZN(n1311) );
INV_X1 U1040 ( .A(G119), .ZN(n1255) );
XOR2_X1 U1041 ( .A(n1323), .B(n1324), .Z(n1318) );
XOR2_X1 U1042 ( .A(KEYINPUT56), .B(KEYINPUT21), .Z(n1324) );
XOR2_X1 U1043 ( .A(n1325), .B(G137), .Z(n1323) );
NAND3_X1 U1044 ( .A1(G221), .A2(n1047), .A3(n1326), .ZN(n1325) );
XNOR2_X1 U1045 ( .A(G234), .B(KEYINPUT40), .ZN(n1326) );
NAND2_X1 U1046 ( .A1(G902), .A2(G217), .ZN(n1313) );
XNOR2_X1 U1047 ( .A(n1327), .B(G472), .ZN(n1242) );
NAND2_X1 U1048 ( .A1(n1328), .A2(n1268), .ZN(n1327) );
XOR2_X1 U1049 ( .A(n1329), .B(n1159), .Z(n1328) );
XOR2_X1 U1050 ( .A(G119), .B(n1276), .Z(n1159) );
XNOR2_X1 U1051 ( .A(G113), .B(n1330), .ZN(n1276) );
XNOR2_X1 U1052 ( .A(n1331), .B(n1332), .ZN(n1329) );
NOR2_X1 U1053 ( .A1(KEYINPUT48), .A2(n1162), .ZN(n1332) );
XOR2_X1 U1054 ( .A(n1273), .B(n1170), .Z(n1162) );
XOR2_X1 U1055 ( .A(n1114), .B(n1118), .Z(n1170) );
XOR2_X1 U1056 ( .A(G137), .B(n1119), .Z(n1118) );
XOR2_X1 U1057 ( .A(G143), .B(n1321), .Z(n1273) );
XOR2_X1 U1058 ( .A(G146), .B(G128), .Z(n1321) );
NOR2_X1 U1059 ( .A1(KEYINPUT31), .A2(n1333), .ZN(n1331) );
XOR2_X1 U1060 ( .A(KEYINPUT53), .B(n1163), .Z(n1333) );
XNOR2_X1 U1061 ( .A(n1334), .B(G101), .ZN(n1163) );
NAND2_X1 U1062 ( .A1(n1335), .A2(G210), .ZN(n1334) );
XOR2_X1 U1063 ( .A(KEYINPUT50), .B(n1063), .Z(n1263) );
INV_X1 U1064 ( .A(n1236), .ZN(n1063) );
NAND2_X1 U1065 ( .A1(n1224), .A2(n1051), .ZN(n1236) );
XNOR2_X1 U1066 ( .A(G475), .B(n1336), .ZN(n1051) );
AND2_X1 U1067 ( .A1(n1144), .A2(n1268), .ZN(n1336) );
INV_X1 U1068 ( .A(G902), .ZN(n1268) );
NAND2_X1 U1069 ( .A1(n1337), .A2(n1338), .ZN(n1144) );
NAND2_X1 U1070 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
XOR2_X1 U1071 ( .A(KEYINPUT5), .B(n1341), .Z(n1337) );
NOR2_X1 U1072 ( .A1(n1339), .A2(n1340), .ZN(n1341) );
XOR2_X1 U1073 ( .A(n1153), .B(n1342), .Z(n1340) );
XOR2_X1 U1074 ( .A(G122), .B(G113), .Z(n1342) );
INV_X1 U1075 ( .A(G104), .ZN(n1153) );
XOR2_X1 U1076 ( .A(n1343), .B(n1344), .Z(n1339) );
XOR2_X1 U1077 ( .A(n1322), .B(n1299), .Z(n1344) );
XOR2_X1 U1078 ( .A(G146), .B(G143), .Z(n1299) );
XOR2_X1 U1079 ( .A(G125), .B(G140), .Z(n1322) );
XOR2_X1 U1080 ( .A(n1345), .B(n1346), .Z(n1343) );
XNOR2_X1 U1081 ( .A(n1347), .B(KEYINPUT43), .ZN(n1346) );
NAND3_X1 U1082 ( .A1(n1335), .A2(G214), .A3(KEYINPUT55), .ZN(n1347) );
NOR2_X1 U1083 ( .A1(G953), .A2(G237), .ZN(n1335) );
NAND2_X1 U1084 ( .A1(KEYINPUT60), .A2(n1114), .ZN(n1345) );
INV_X1 U1085 ( .A(G131), .ZN(n1114) );
INV_X1 U1086 ( .A(n1253), .ZN(n1224) );
NAND2_X1 U1087 ( .A1(n1348), .A2(n1349), .ZN(n1253) );
NAND2_X1 U1088 ( .A1(G478), .A2(n1350), .ZN(n1349) );
OR2_X1 U1089 ( .A1(n1062), .A2(G902), .ZN(n1350) );
XNOR2_X1 U1090 ( .A(n1058), .B(KEYINPUT28), .ZN(n1348) );
NOR3_X1 U1091 ( .A1(G478), .A2(G902), .A3(n1062), .ZN(n1058) );
XNOR2_X1 U1092 ( .A(n1351), .B(n1352), .ZN(n1062) );
XOR2_X1 U1093 ( .A(n1353), .B(n1354), .Z(n1352) );
NAND2_X1 U1094 ( .A1(KEYINPUT42), .A2(n1330), .ZN(n1354) );
INV_X1 U1095 ( .A(G116), .ZN(n1330) );
NAND3_X1 U1096 ( .A1(n1355), .A2(n1356), .A3(n1357), .ZN(n1353) );
OR2_X1 U1097 ( .A1(n1358), .A2(G134), .ZN(n1357) );
NAND2_X1 U1098 ( .A1(n1359), .A2(n1360), .ZN(n1356) );
INV_X1 U1099 ( .A(KEYINPUT27), .ZN(n1360) );
NAND2_X1 U1100 ( .A1(n1361), .A2(n1358), .ZN(n1359) );
XOR2_X1 U1101 ( .A(KEYINPUT25), .B(n1119), .Z(n1361) );
INV_X1 U1102 ( .A(G134), .ZN(n1119) );
NAND2_X1 U1103 ( .A1(KEYINPUT27), .A2(n1362), .ZN(n1355) );
NAND2_X1 U1104 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
OR2_X1 U1105 ( .A1(G134), .A2(KEYINPUT25), .ZN(n1364) );
NAND3_X1 U1106 ( .A1(G134), .A2(n1358), .A3(KEYINPUT25), .ZN(n1363) );
XOR2_X1 U1107 ( .A(G143), .B(G128), .Z(n1358) );
XOR2_X1 U1108 ( .A(n1365), .B(n1366), .Z(n1351) );
XOR2_X1 U1109 ( .A(G122), .B(G107), .Z(n1366) );
NAND3_X1 U1110 ( .A1(G234), .A2(n1047), .A3(G217), .ZN(n1365) );
INV_X1 U1111 ( .A(G953), .ZN(n1047) );
endmodule


