//Key = 0111110001101101010010111110001010111000000101111101111000110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426;

XNOR2_X1 U778 ( .A(G107), .B(n1079), .ZN(G9) );
NAND3_X1 U779 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(G75) );
NAND2_X1 U780 ( .A1(G952), .A2(n1083), .ZN(n1082) );
NAND4_X1 U781 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1083) );
NOR2_X1 U782 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR2_X1 U783 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
INV_X1 U784 ( .A(KEYINPUT29), .ZN(n1091) );
NOR3_X1 U785 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1090) );
NOR3_X1 U786 ( .A1(n1095), .A2(n1096), .A3(n1094), .ZN(n1088) );
NOR2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NOR2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR2_X1 U790 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NOR2_X1 U792 ( .A1(n1107), .A2(n1108), .ZN(n1101) );
NOR2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
NOR2_X1 U794 ( .A1(KEYINPUT29), .A2(n1093), .ZN(n1110) );
NOR3_X1 U795 ( .A1(n1111), .A2(KEYINPUT60), .A3(n1112), .ZN(n1109) );
NOR3_X1 U796 ( .A1(n1104), .A2(n1113), .A3(n1108), .ZN(n1097) );
NOR2_X1 U797 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1085) );
NAND3_X1 U799 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1117) );
NAND2_X1 U800 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U801 ( .A1(KEYINPUT60), .A2(n1123), .ZN(n1119) );
NAND2_X1 U802 ( .A1(n1124), .A2(n1125), .ZN(n1118) );
INV_X1 U803 ( .A(KEYINPUT57), .ZN(n1125) );
NAND3_X1 U804 ( .A1(KEYINPUT57), .A2(n1124), .A3(n1126), .ZN(n1084) );
INV_X1 U805 ( .A(n1116), .ZN(n1126) );
NOR2_X1 U806 ( .A1(n1092), .A2(n1104), .ZN(n1116) );
OR3_X1 U807 ( .A1(n1100), .A2(n1108), .A3(n1095), .ZN(n1092) );
XNOR2_X1 U808 ( .A(n1127), .B(KEYINPUT62), .ZN(n1095) );
INV_X1 U809 ( .A(n1128), .ZN(n1108) );
INV_X1 U810 ( .A(n1129), .ZN(n1100) );
NAND4_X1 U811 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1080) );
NOR4_X1 U812 ( .A1(n1121), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n1133) );
NOR2_X1 U813 ( .A1(KEYINPUT58), .A2(n1137), .ZN(n1136) );
NOR2_X1 U814 ( .A1(n1138), .A2(G472), .ZN(n1137) );
NOR2_X1 U815 ( .A1(KEYINPUT30), .A2(n1139), .ZN(n1138) );
XNOR2_X1 U816 ( .A(n1140), .B(n1141), .ZN(n1135) );
NAND2_X1 U817 ( .A1(KEYINPUT53), .A2(n1142), .ZN(n1140) );
XOR2_X1 U818 ( .A(n1143), .B(n1144), .Z(n1134) );
NAND2_X1 U819 ( .A1(KEYINPUT4), .A2(n1145), .ZN(n1143) );
NOR3_X1 U820 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1132) );
NOR2_X1 U821 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR3_X1 U822 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
NOR2_X1 U823 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
INV_X1 U824 ( .A(KEYINPUT17), .ZN(n1155) );
NOR2_X1 U825 ( .A1(n1156), .A2(G472), .ZN(n1154) );
NOR2_X1 U826 ( .A1(KEYINPUT30), .A2(n1157), .ZN(n1156) );
NOR2_X1 U827 ( .A1(KEYINPUT17), .A2(G472), .ZN(n1152) );
NOR2_X1 U828 ( .A1(KEYINPUT58), .A2(n1158), .ZN(n1151) );
INV_X1 U829 ( .A(n1139), .ZN(n1149) );
NOR4_X1 U830 ( .A1(n1139), .A2(n1157), .A3(G472), .A4(n1158), .ZN(n1147) );
INV_X1 U831 ( .A(KEYINPUT30), .ZN(n1158) );
INV_X1 U832 ( .A(KEYINPUT58), .ZN(n1157) );
XOR2_X1 U833 ( .A(G478), .B(n1159), .Z(n1146) );
XOR2_X1 U834 ( .A(n1160), .B(n1161), .Z(G72) );
XOR2_X1 U835 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U836 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XOR2_X1 U837 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1167) );
XNOR2_X1 U839 ( .A(n1170), .B(n1171), .ZN(n1166) );
NOR2_X1 U840 ( .A1(KEYINPUT40), .A2(n1172), .ZN(n1171) );
XOR2_X1 U841 ( .A(n1173), .B(G134), .Z(n1172) );
NAND2_X1 U842 ( .A1(n1081), .A2(n1174), .ZN(n1162) );
NAND4_X1 U843 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1174) );
NAND2_X1 U844 ( .A1(G953), .A2(n1179), .ZN(n1160) );
NAND2_X1 U845 ( .A1(G900), .A2(G227), .ZN(n1179) );
XOR2_X1 U846 ( .A(n1180), .B(n1181), .Z(G69) );
XOR2_X1 U847 ( .A(n1182), .B(n1183), .Z(n1181) );
NAND3_X1 U848 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1183) );
NAND2_X1 U849 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND2_X1 U850 ( .A1(n1189), .A2(n1190), .ZN(n1185) );
NAND2_X1 U851 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NAND2_X1 U852 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
INV_X1 U853 ( .A(KEYINPUT5), .ZN(n1194) );
XOR2_X1 U854 ( .A(n1195), .B(KEYINPUT14), .Z(n1191) );
INV_X1 U855 ( .A(n1196), .ZN(n1189) );
NAND3_X1 U856 ( .A1(KEYINPUT5), .A2(n1193), .A3(n1196), .ZN(n1184) );
XOR2_X1 U857 ( .A(n1195), .B(KEYINPUT37), .Z(n1193) );
XOR2_X1 U858 ( .A(n1197), .B(n1198), .Z(n1195) );
NAND2_X1 U859 ( .A1(KEYINPUT15), .A2(n1199), .ZN(n1197) );
NAND2_X1 U860 ( .A1(n1200), .A2(n1081), .ZN(n1182) );
XNOR2_X1 U861 ( .A(n1201), .B(KEYINPUT7), .ZN(n1200) );
NOR2_X1 U862 ( .A1(n1202), .A2(n1081), .ZN(n1180) );
NOR2_X1 U863 ( .A1(n1203), .A2(n1188), .ZN(n1202) );
NOR2_X1 U864 ( .A1(n1204), .A2(n1205), .ZN(G66) );
XOR2_X1 U865 ( .A(n1206), .B(n1207), .Z(n1205) );
NOR2_X1 U866 ( .A1(KEYINPUT11), .A2(n1208), .ZN(n1207) );
NAND2_X1 U867 ( .A1(n1209), .A2(G217), .ZN(n1206) );
NOR2_X1 U868 ( .A1(n1204), .A2(n1210), .ZN(G63) );
NOR3_X1 U869 ( .A1(n1211), .A2(n1159), .A3(n1212), .ZN(n1210) );
NOR2_X1 U870 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NOR2_X1 U871 ( .A1(n1086), .A2(n1215), .ZN(n1213) );
XOR2_X1 U872 ( .A(KEYINPUT50), .B(n1216), .Z(n1211) );
AND3_X1 U873 ( .A1(n1209), .A2(n1214), .A3(G478), .ZN(n1216) );
NOR2_X1 U874 ( .A1(n1204), .A2(n1217), .ZN(G60) );
XOR2_X1 U875 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U876 ( .A(n1220), .B(KEYINPUT24), .Z(n1218) );
NAND2_X1 U877 ( .A1(n1209), .A2(G475), .ZN(n1220) );
XOR2_X1 U878 ( .A(n1221), .B(n1222), .Z(G6) );
NOR2_X1 U879 ( .A1(n1223), .A2(n1224), .ZN(G57) );
XOR2_X1 U880 ( .A(KEYINPUT19), .B(n1204), .Z(n1224) );
XOR2_X1 U881 ( .A(n1225), .B(n1226), .Z(n1223) );
NOR2_X1 U882 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NOR2_X1 U883 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NOR2_X1 U884 ( .A1(n1231), .A2(n1232), .ZN(n1229) );
NOR3_X1 U885 ( .A1(n1233), .A2(n1231), .A3(n1232), .ZN(n1227) );
XNOR2_X1 U886 ( .A(KEYINPUT31), .B(n1230), .ZN(n1233) );
XOR2_X1 U887 ( .A(n1234), .B(n1235), .Z(n1230) );
NAND2_X1 U888 ( .A1(KEYINPUT35), .A2(n1198), .ZN(n1234) );
NAND2_X1 U889 ( .A1(KEYINPUT26), .A2(n1236), .ZN(n1225) );
NOR2_X1 U890 ( .A1(n1204), .A2(n1237), .ZN(G54) );
XOR2_X1 U891 ( .A(n1238), .B(n1239), .Z(n1237) );
NAND2_X1 U892 ( .A1(n1209), .A2(G469), .ZN(n1239) );
NAND3_X1 U893 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1238) );
NAND2_X1 U894 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
NAND2_X1 U895 ( .A1(KEYINPUT45), .A2(n1245), .ZN(n1244) );
XOR2_X1 U896 ( .A(KEYINPUT41), .B(n1246), .Z(n1245) );
INV_X1 U897 ( .A(n1247), .ZN(n1243) );
NAND3_X1 U898 ( .A1(KEYINPUT45), .A2(n1247), .A3(n1246), .ZN(n1241) );
OR2_X1 U899 ( .A1(n1246), .A2(KEYINPUT45), .ZN(n1240) );
XNOR2_X1 U900 ( .A(n1248), .B(n1249), .ZN(n1246) );
NAND2_X1 U901 ( .A1(KEYINPUT54), .A2(n1250), .ZN(n1248) );
NOR2_X1 U902 ( .A1(n1204), .A2(n1251), .ZN(G51) );
XOR2_X1 U903 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U904 ( .A(n1254), .B(n1255), .Z(n1253) );
OR2_X1 U905 ( .A1(n1232), .A2(n1142), .ZN(n1254) );
INV_X1 U906 ( .A(n1209), .ZN(n1232) );
NOR2_X1 U907 ( .A1(n1256), .A2(n1086), .ZN(n1209) );
AND3_X1 U908 ( .A1(n1201), .A2(n1257), .A3(n1258), .ZN(n1086) );
AND3_X1 U909 ( .A1(n1176), .A2(n1178), .A3(n1177), .ZN(n1258) );
NAND2_X1 U910 ( .A1(n1123), .A2(n1259), .ZN(n1176) );
NAND2_X1 U911 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND3_X1 U912 ( .A1(n1115), .A2(n1106), .A3(n1262), .ZN(n1261) );
XNOR2_X1 U913 ( .A(KEYINPUT59), .B(n1263), .ZN(n1260) );
XOR2_X1 U914 ( .A(KEYINPUT44), .B(n1175), .Z(n1257) );
AND4_X1 U915 ( .A1(n1264), .A2(n1265), .A3(n1266), .A4(n1267), .ZN(n1175) );
NAND2_X1 U916 ( .A1(n1268), .A2(n1269), .ZN(n1264) );
XNOR2_X1 U917 ( .A(n1124), .B(KEYINPUT34), .ZN(n1268) );
AND2_X1 U918 ( .A1(n1270), .A2(n1271), .ZN(n1201) );
AND4_X1 U919 ( .A1(n1079), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1271) );
NAND3_X1 U920 ( .A1(n1114), .A2(n1128), .A3(n1275), .ZN(n1079) );
AND4_X1 U921 ( .A1(n1276), .A2(n1277), .A3(n1278), .A4(n1222), .ZN(n1270) );
NAND3_X1 U922 ( .A1(n1275), .A2(n1128), .A3(n1115), .ZN(n1222) );
XOR2_X1 U923 ( .A(n1279), .B(n1280), .Z(n1252) );
XOR2_X1 U924 ( .A(G125), .B(n1281), .Z(n1280) );
NOR2_X1 U925 ( .A1(KEYINPUT8), .A2(n1282), .ZN(n1279) );
AND2_X1 U926 ( .A1(G953), .A2(n1283), .ZN(n1204) );
XOR2_X1 U927 ( .A(KEYINPUT2), .B(G952), .Z(n1283) );
XNOR2_X1 U928 ( .A(n1284), .B(n1177), .ZN(G48) );
NAND3_X1 U929 ( .A1(n1115), .A2(n1124), .A3(n1285), .ZN(n1177) );
NAND2_X1 U930 ( .A1(KEYINPUT13), .A2(n1286), .ZN(n1284) );
INV_X1 U931 ( .A(G146), .ZN(n1286) );
XOR2_X1 U932 ( .A(n1287), .B(n1178), .Z(G45) );
NAND4_X1 U933 ( .A1(n1124), .A2(n1288), .A3(n1289), .A4(n1290), .ZN(n1178) );
NOR2_X1 U934 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
NAND3_X1 U935 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(G42) );
OR2_X1 U936 ( .A1(n1296), .A2(G140), .ZN(n1295) );
NAND2_X1 U937 ( .A1(KEYINPUT42), .A2(n1297), .ZN(n1294) );
NAND2_X1 U938 ( .A1(G140), .A2(n1298), .ZN(n1297) );
XNOR2_X1 U939 ( .A(KEYINPUT61), .B(n1296), .ZN(n1298) );
NAND2_X1 U940 ( .A1(n1299), .A2(n1300), .ZN(n1293) );
INV_X1 U941 ( .A(KEYINPUT42), .ZN(n1300) );
NAND2_X1 U942 ( .A1(n1301), .A2(n1302), .ZN(n1299) );
NAND3_X1 U943 ( .A1(KEYINPUT61), .A2(G140), .A3(n1296), .ZN(n1302) );
OR2_X1 U944 ( .A1(n1296), .A2(KEYINPUT61), .ZN(n1301) );
NAND4_X1 U945 ( .A1(n1303), .A2(n1123), .A3(n1262), .A4(n1115), .ZN(n1296) );
INV_X1 U946 ( .A(n1094), .ZN(n1123) );
XNOR2_X1 U947 ( .A(n1106), .B(KEYINPUT3), .ZN(n1303) );
XOR2_X1 U948 ( .A(G137), .B(n1304), .Z(G39) );
NOR2_X1 U949 ( .A1(n1263), .A2(n1094), .ZN(n1304) );
NAND2_X1 U950 ( .A1(n1285), .A2(n1129), .ZN(n1263) );
NAND2_X1 U951 ( .A1(n1305), .A2(n1306), .ZN(G36) );
OR2_X1 U952 ( .A1(n1265), .A2(G134), .ZN(n1306) );
XOR2_X1 U953 ( .A(n1307), .B(KEYINPUT55), .Z(n1305) );
NAND2_X1 U954 ( .A1(G134), .A2(n1265), .ZN(n1307) );
NAND2_X1 U955 ( .A1(n1308), .A2(n1114), .ZN(n1265) );
XNOR2_X1 U956 ( .A(G131), .B(n1266), .ZN(G33) );
NAND2_X1 U957 ( .A1(n1308), .A2(n1115), .ZN(n1266) );
NOR3_X1 U958 ( .A1(n1292), .A2(n1291), .A3(n1094), .ZN(n1308) );
NAND2_X1 U959 ( .A1(n1122), .A2(n1309), .ZN(n1094) );
XNOR2_X1 U960 ( .A(n1267), .B(n1310), .ZN(G30) );
NOR2_X1 U961 ( .A1(KEYINPUT18), .A2(n1311), .ZN(n1310) );
INV_X1 U962 ( .A(G128), .ZN(n1311) );
NAND3_X1 U963 ( .A1(n1114), .A2(n1124), .A3(n1285), .ZN(n1267) );
AND3_X1 U964 ( .A1(n1312), .A2(n1313), .A3(n1262), .ZN(n1285) );
INV_X1 U965 ( .A(n1292), .ZN(n1262) );
NAND2_X1 U966 ( .A1(n1314), .A2(n1315), .ZN(n1292) );
XOR2_X1 U967 ( .A(n1316), .B(n1278), .Z(G3) );
NAND3_X1 U968 ( .A1(n1129), .A2(n1275), .A3(n1105), .ZN(n1278) );
NAND3_X1 U969 ( .A1(n1317), .A2(n1318), .A3(n1319), .ZN(G27) );
NAND3_X1 U970 ( .A1(n1124), .A2(n1320), .A3(n1269), .ZN(n1319) );
NAND2_X1 U971 ( .A1(KEYINPUT25), .A2(n1321), .ZN(n1320) );
NAND2_X1 U972 ( .A1(KEYINPUT22), .A2(n1322), .ZN(n1321) );
OR2_X1 U973 ( .A1(G125), .A2(KEYINPUT25), .ZN(n1318) );
NAND3_X1 U974 ( .A1(G125), .A2(n1323), .A3(KEYINPUT25), .ZN(n1317) );
NAND3_X1 U975 ( .A1(n1269), .A2(n1124), .A3(KEYINPUT22), .ZN(n1323) );
AND4_X1 U976 ( .A1(n1115), .A2(n1130), .A3(n1106), .A4(n1315), .ZN(n1269) );
NAND2_X1 U977 ( .A1(n1324), .A2(n1325), .ZN(n1315) );
NAND3_X1 U978 ( .A1(G902), .A2(n1127), .A3(n1164), .ZN(n1325) );
NOR2_X1 U979 ( .A1(n1326), .A2(G900), .ZN(n1164) );
INV_X1 U980 ( .A(n1187), .ZN(n1326) );
INV_X1 U981 ( .A(n1327), .ZN(n1115) );
XOR2_X1 U982 ( .A(n1277), .B(n1328), .Z(G24) );
XOR2_X1 U983 ( .A(KEYINPUT46), .B(G122), .Z(n1328) );
NAND4_X1 U984 ( .A1(n1289), .A2(n1329), .A3(n1128), .A4(n1288), .ZN(n1277) );
NAND2_X1 U985 ( .A1(n1330), .A2(n1331), .ZN(n1128) );
OR3_X1 U986 ( .A1(n1313), .A2(n1312), .A3(KEYINPUT33), .ZN(n1331) );
NAND2_X1 U987 ( .A1(KEYINPUT33), .A2(n1106), .ZN(n1330) );
XNOR2_X1 U988 ( .A(G119), .B(n1276), .ZN(G21) );
NAND4_X1 U989 ( .A1(n1329), .A2(n1129), .A3(n1312), .A4(n1313), .ZN(n1276) );
XNOR2_X1 U990 ( .A(G116), .B(n1274), .ZN(G18) );
NAND3_X1 U991 ( .A1(n1105), .A2(n1114), .A3(n1329), .ZN(n1274) );
AND3_X1 U992 ( .A1(n1124), .A2(n1332), .A3(n1130), .ZN(n1329) );
NOR2_X1 U993 ( .A1(n1288), .A2(n1333), .ZN(n1114) );
INV_X1 U994 ( .A(n1291), .ZN(n1105) );
XNOR2_X1 U995 ( .A(G113), .B(n1273), .ZN(G15) );
NAND4_X1 U996 ( .A1(n1334), .A2(n1332), .A3(n1130), .A4(n1335), .ZN(n1273) );
NOR2_X1 U997 ( .A1(n1327), .A2(n1291), .ZN(n1335) );
NAND2_X1 U998 ( .A1(n1336), .A2(n1312), .ZN(n1291) );
XOR2_X1 U999 ( .A(KEYINPUT33), .B(n1131), .Z(n1336) );
NAND2_X1 U1000 ( .A1(n1333), .A2(n1288), .ZN(n1327) );
INV_X1 U1001 ( .A(n1104), .ZN(n1130) );
NAND2_X1 U1002 ( .A1(n1337), .A2(n1111), .ZN(n1104) );
XOR2_X1 U1003 ( .A(n1250), .B(n1272), .Z(G12) );
NAND3_X1 U1004 ( .A1(n1275), .A2(n1106), .A3(n1129), .ZN(n1272) );
NOR2_X1 U1005 ( .A1(n1288), .A2(n1289), .ZN(n1129) );
INV_X1 U1006 ( .A(n1333), .ZN(n1289) );
NAND2_X1 U1007 ( .A1(n1338), .A2(n1339), .ZN(n1333) );
NAND2_X1 U1008 ( .A1(n1340), .A2(n1215), .ZN(n1339) );
INV_X1 U1009 ( .A(G478), .ZN(n1215) );
XNOR2_X1 U1010 ( .A(n1159), .B(KEYINPUT38), .ZN(n1340) );
NAND2_X1 U1011 ( .A1(n1341), .A2(G478), .ZN(n1338) );
XNOR2_X1 U1012 ( .A(n1159), .B(KEYINPUT32), .ZN(n1341) );
NOR2_X1 U1013 ( .A1(n1214), .A2(G902), .ZN(n1159) );
XNOR2_X1 U1014 ( .A(n1342), .B(n1343), .ZN(n1214) );
XOR2_X1 U1015 ( .A(n1344), .B(n1345), .Z(n1343) );
XOR2_X1 U1016 ( .A(G122), .B(G116), .Z(n1345) );
XOR2_X1 U1017 ( .A(G143), .B(G134), .Z(n1344) );
XOR2_X1 U1018 ( .A(n1346), .B(n1347), .Z(n1342) );
XOR2_X1 U1019 ( .A(n1348), .B(G107), .Z(n1346) );
NAND3_X1 U1020 ( .A1(G234), .A2(n1081), .A3(G217), .ZN(n1348) );
NAND2_X1 U1021 ( .A1(n1349), .A2(n1350), .ZN(n1288) );
OR2_X1 U1022 ( .A1(n1145), .A2(n1144), .ZN(n1350) );
XOR2_X1 U1023 ( .A(n1351), .B(KEYINPUT21), .Z(n1349) );
NAND2_X1 U1024 ( .A1(n1144), .A2(n1145), .ZN(n1351) );
INV_X1 U1025 ( .A(G475), .ZN(n1145) );
NOR2_X1 U1026 ( .A1(n1219), .A2(G902), .ZN(n1144) );
XNOR2_X1 U1027 ( .A(n1352), .B(n1353), .ZN(n1219) );
XOR2_X1 U1028 ( .A(n1354), .B(n1355), .Z(n1353) );
XOR2_X1 U1029 ( .A(n1356), .B(n1357), .Z(n1355) );
NAND2_X1 U1030 ( .A1(n1358), .A2(G214), .ZN(n1356) );
XOR2_X1 U1031 ( .A(n1359), .B(n1360), .Z(n1352) );
XOR2_X1 U1032 ( .A(G122), .B(G113), .Z(n1360) );
XOR2_X1 U1033 ( .A(n1361), .B(G104), .Z(n1359) );
NAND2_X1 U1034 ( .A1(n1362), .A2(KEYINPUT48), .ZN(n1361) );
XNOR2_X1 U1035 ( .A(n1170), .B(KEYINPUT47), .ZN(n1362) );
NOR2_X1 U1036 ( .A1(n1312), .A2(n1131), .ZN(n1106) );
INV_X1 U1037 ( .A(n1313), .ZN(n1131) );
NAND3_X1 U1038 ( .A1(n1363), .A2(n1364), .A3(n1365), .ZN(n1313) );
NAND2_X1 U1039 ( .A1(n1366), .A2(n1208), .ZN(n1365) );
OR3_X1 U1040 ( .A1(n1208), .A2(n1366), .A3(G902), .ZN(n1364) );
NOR2_X1 U1041 ( .A1(n1367), .A2(G234), .ZN(n1366) );
INV_X1 U1042 ( .A(G217), .ZN(n1367) );
XNOR2_X1 U1043 ( .A(n1368), .B(n1369), .ZN(n1208) );
XOR2_X1 U1044 ( .A(n1173), .B(n1370), .Z(n1369) );
NAND3_X1 U1045 ( .A1(G234), .A2(n1081), .A3(G221), .ZN(n1370) );
NAND2_X1 U1046 ( .A1(n1371), .A2(n1372), .ZN(n1368) );
NAND2_X1 U1047 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
XOR2_X1 U1048 ( .A(KEYINPUT36), .B(n1375), .Z(n1371) );
NOR2_X1 U1049 ( .A1(n1374), .A2(n1373), .ZN(n1375) );
XOR2_X1 U1050 ( .A(G146), .B(n1170), .Z(n1373) );
XOR2_X1 U1051 ( .A(G140), .B(G125), .Z(n1170) );
XNOR2_X1 U1052 ( .A(n1376), .B(n1377), .ZN(n1374) );
XOR2_X1 U1053 ( .A(G119), .B(G110), .Z(n1377) );
NAND2_X1 U1054 ( .A1(KEYINPUT9), .A2(n1347), .ZN(n1376) );
NAND2_X1 U1055 ( .A1(G217), .A2(G902), .ZN(n1363) );
XOR2_X1 U1056 ( .A(n1139), .B(n1231), .Z(n1312) );
INV_X1 U1057 ( .A(G472), .ZN(n1231) );
NAND2_X1 U1058 ( .A1(n1378), .A2(n1256), .ZN(n1139) );
XNOR2_X1 U1059 ( .A(n1236), .B(n1379), .ZN(n1378) );
XOR2_X1 U1060 ( .A(n1380), .B(n1198), .Z(n1379) );
NAND2_X1 U1061 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
NAND2_X1 U1062 ( .A1(n1169), .A2(n1383), .ZN(n1382) );
NAND2_X1 U1063 ( .A1(n1384), .A2(n1282), .ZN(n1381) );
XNOR2_X1 U1064 ( .A(KEYINPUT39), .B(n1383), .ZN(n1384) );
AND2_X1 U1065 ( .A1(n1385), .A2(n1386), .ZN(n1236) );
NAND2_X1 U1066 ( .A1(n1387), .A2(n1316), .ZN(n1386) );
NAND2_X1 U1067 ( .A1(n1358), .A2(G210), .ZN(n1387) );
NAND3_X1 U1068 ( .A1(n1358), .A2(G210), .A3(G101), .ZN(n1385) );
NOR2_X1 U1069 ( .A1(G953), .A2(G237), .ZN(n1358) );
AND3_X1 U1070 ( .A1(n1334), .A2(n1332), .A3(n1314), .ZN(n1275) );
INV_X1 U1071 ( .A(n1093), .ZN(n1314) );
NAND2_X1 U1072 ( .A1(n1112), .A2(n1111), .ZN(n1093) );
NAND2_X1 U1073 ( .A1(G221), .A2(n1388), .ZN(n1111) );
NAND2_X1 U1074 ( .A1(G234), .A2(n1256), .ZN(n1388) );
INV_X1 U1075 ( .A(n1337), .ZN(n1112) );
XOR2_X1 U1076 ( .A(n1389), .B(G469), .Z(n1337) );
NAND2_X1 U1077 ( .A1(n1390), .A2(n1256), .ZN(n1389) );
XOR2_X1 U1078 ( .A(n1249), .B(n1391), .Z(n1390) );
XOR2_X1 U1079 ( .A(n1392), .B(n1247), .Z(n1391) );
XNOR2_X1 U1080 ( .A(n1235), .B(n1393), .ZN(n1247) );
XOR2_X1 U1081 ( .A(n1394), .B(n1395), .Z(n1393) );
NAND2_X1 U1082 ( .A1(KEYINPUT63), .A2(n1221), .ZN(n1394) );
XNOR2_X1 U1083 ( .A(n1383), .B(n1169), .ZN(n1235) );
INV_X1 U1084 ( .A(n1282), .ZN(n1169) );
NAND2_X1 U1085 ( .A1(n1396), .A2(n1397), .ZN(n1383) );
NAND2_X1 U1086 ( .A1(n1398), .A2(n1168), .ZN(n1397) );
XOR2_X1 U1087 ( .A(n1399), .B(G134), .Z(n1398) );
XOR2_X1 U1088 ( .A(n1400), .B(KEYINPUT56), .Z(n1396) );
NAND2_X1 U1089 ( .A1(n1401), .A2(n1357), .ZN(n1400) );
INV_X1 U1090 ( .A(n1168), .ZN(n1357) );
XNOR2_X1 U1091 ( .A(G131), .B(KEYINPUT52), .ZN(n1168) );
XNOR2_X1 U1092 ( .A(G134), .B(n1399), .ZN(n1401) );
NAND2_X1 U1093 ( .A1(KEYINPUT20), .A2(n1173), .ZN(n1399) );
INV_X1 U1094 ( .A(G137), .ZN(n1173) );
NAND2_X1 U1095 ( .A1(KEYINPUT43), .A2(n1250), .ZN(n1392) );
XOR2_X1 U1096 ( .A(G140), .B(n1402), .Z(n1249) );
AND2_X1 U1097 ( .A1(n1081), .A2(G227), .ZN(n1402) );
NAND2_X1 U1098 ( .A1(n1324), .A2(n1403), .ZN(n1332) );
NAND4_X1 U1099 ( .A1(G902), .A2(n1187), .A3(n1127), .A4(n1188), .ZN(n1403) );
INV_X1 U1100 ( .A(G898), .ZN(n1188) );
XOR2_X1 U1101 ( .A(G953), .B(KEYINPUT6), .Z(n1187) );
NAND3_X1 U1102 ( .A1(n1127), .A2(n1081), .A3(G952), .ZN(n1324) );
INV_X1 U1103 ( .A(G953), .ZN(n1081) );
NAND2_X1 U1104 ( .A1(G237), .A2(G234), .ZN(n1127) );
XOR2_X1 U1105 ( .A(n1124), .B(KEYINPUT16), .Z(n1334) );
NOR2_X1 U1106 ( .A1(n1404), .A2(n1122), .ZN(n1124) );
XOR2_X1 U1107 ( .A(n1405), .B(n1142), .Z(n1122) );
NAND2_X1 U1108 ( .A1(G210), .A2(n1406), .ZN(n1142) );
XOR2_X1 U1109 ( .A(n1141), .B(KEYINPUT23), .Z(n1405) );
NAND3_X1 U1110 ( .A1(n1407), .A2(n1256), .A3(n1408), .ZN(n1141) );
XOR2_X1 U1111 ( .A(KEYINPUT1), .B(n1409), .Z(n1408) );
NOR2_X1 U1112 ( .A1(n1410), .A2(n1411), .ZN(n1409) );
NAND2_X1 U1113 ( .A1(n1410), .A2(n1411), .ZN(n1407) );
XNOR2_X1 U1114 ( .A(KEYINPUT51), .B(n1255), .ZN(n1411) );
XNOR2_X1 U1115 ( .A(n1412), .B(n1199), .ZN(n1255) );
XNOR2_X1 U1116 ( .A(n1395), .B(n1221), .ZN(n1199) );
INV_X1 U1117 ( .A(G104), .ZN(n1221) );
XOR2_X1 U1118 ( .A(n1316), .B(n1413), .Z(n1395) );
XOR2_X1 U1119 ( .A(KEYINPUT49), .B(G107), .Z(n1413) );
INV_X1 U1120 ( .A(G101), .ZN(n1316) );
XOR2_X1 U1121 ( .A(n1196), .B(n1198), .Z(n1412) );
XOR2_X1 U1122 ( .A(G113), .B(n1414), .Z(n1198) );
XOR2_X1 U1123 ( .A(G119), .B(G116), .Z(n1414) );
NAND2_X1 U1124 ( .A1(n1415), .A2(n1416), .ZN(n1196) );
NAND2_X1 U1125 ( .A1(G122), .A2(n1250), .ZN(n1416) );
XOR2_X1 U1126 ( .A(n1417), .B(KEYINPUT28), .Z(n1415) );
NAND2_X1 U1127 ( .A1(G110), .A2(n1418), .ZN(n1417) );
INV_X1 U1128 ( .A(G122), .ZN(n1418) );
AND2_X1 U1129 ( .A1(n1419), .A2(n1420), .ZN(n1410) );
NAND2_X1 U1130 ( .A1(n1421), .A2(n1422), .ZN(n1420) );
XOR2_X1 U1131 ( .A(G125), .B(n1423), .Z(n1422) );
XNOR2_X1 U1132 ( .A(KEYINPUT10), .B(n1281), .ZN(n1421) );
NAND2_X1 U1133 ( .A1(n1424), .A2(n1425), .ZN(n1419) );
XOR2_X1 U1134 ( .A(KEYINPUT10), .B(n1281), .Z(n1425) );
NOR2_X1 U1135 ( .A1(n1203), .A2(G953), .ZN(n1281) );
INV_X1 U1136 ( .A(G224), .ZN(n1203) );
XOR2_X1 U1137 ( .A(n1322), .B(n1423), .Z(n1424) );
NOR2_X1 U1138 ( .A1(KEYINPUT27), .A2(n1282), .ZN(n1423) );
XOR2_X1 U1139 ( .A(n1354), .B(n1347), .Z(n1282) );
XOR2_X1 U1140 ( .A(G128), .B(KEYINPUT12), .Z(n1347) );
XOR2_X1 U1141 ( .A(n1287), .B(G146), .Z(n1354) );
INV_X1 U1142 ( .A(G143), .ZN(n1287) );
INV_X1 U1143 ( .A(G125), .ZN(n1322) );
XOR2_X1 U1144 ( .A(n1121), .B(KEYINPUT0), .Z(n1404) );
INV_X1 U1145 ( .A(n1309), .ZN(n1121) );
NAND2_X1 U1146 ( .A1(G214), .A2(n1406), .ZN(n1309) );
NAND2_X1 U1147 ( .A1(n1426), .A2(n1256), .ZN(n1406) );
INV_X1 U1148 ( .A(G902), .ZN(n1256) );
INV_X1 U1149 ( .A(G237), .ZN(n1426) );
INV_X1 U1150 ( .A(G110), .ZN(n1250) );
endmodule


