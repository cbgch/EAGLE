//Key = 0100110010001001110010101100010010101000110010011111101100010110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420;

XNOR2_X1 U786 ( .A(n1081), .B(n1082), .ZN(G9) );
NOR2_X1 U787 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U788 ( .A1(n1085), .A2(n1086), .ZN(G75) );
NOR2_X1 U789 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND4_X1 U790 ( .A1(n1089), .A2(n1090), .A3(G952), .A4(n1091), .ZN(n1088) );
NAND2_X1 U791 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U792 ( .A(n1094), .B(KEYINPUT9), .Z(n1089) );
NAND2_X1 U793 ( .A1(n1092), .A2(n1095), .ZN(n1094) );
AND3_X1 U794 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1092) );
NAND4_X1 U795 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1087) );
NAND3_X1 U796 ( .A1(n1103), .A2(n1104), .A3(n1098), .ZN(n1100) );
NAND3_X1 U797 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1104) );
NAND2_X1 U798 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U799 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND3_X1 U800 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
XNOR2_X1 U801 ( .A(KEYINPUT7), .B(n1115), .ZN(n1112) );
NAND3_X1 U802 ( .A1(n1096), .A2(n1116), .A3(KEYINPUT49), .ZN(n1110) );
NAND3_X1 U803 ( .A1(n1117), .A2(n1118), .A3(n1096), .ZN(n1106) );
NAND2_X1 U804 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U805 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
INV_X1 U806 ( .A(n1123), .ZN(n1119) );
NAND2_X1 U807 ( .A1(n1097), .A2(n1124), .ZN(n1105) );
NAND2_X1 U808 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
OR2_X1 U809 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND3_X1 U810 ( .A1(n1129), .A2(n1130), .A3(n1096), .ZN(n1099) );
INV_X1 U811 ( .A(KEYINPUT49), .ZN(n1130) );
NAND4_X1 U812 ( .A1(n1098), .A2(n1103), .A3(n1116), .A4(n1108), .ZN(n1129) );
INV_X1 U813 ( .A(n1131), .ZN(n1098) );
NOR3_X1 U814 ( .A1(n1132), .A2(G953), .A3(n1133), .ZN(n1085) );
INV_X1 U815 ( .A(n1101), .ZN(n1133) );
NAND4_X1 U816 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1101) );
NOR3_X1 U817 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1137) );
XOR2_X1 U818 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U819 ( .A1(KEYINPUT63), .A2(n1143), .ZN(n1142) );
NAND3_X1 U820 ( .A1(n1144), .A2(n1127), .A3(n1145), .ZN(n1138) );
NOR3_X1 U821 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1136) );
AND2_X1 U822 ( .A1(n1149), .A2(KEYINPUT60), .ZN(n1148) );
NOR3_X1 U823 ( .A1(KEYINPUT60), .A2(n1150), .A3(n1149), .ZN(n1147) );
XNOR2_X1 U824 ( .A(G475), .B(n1151), .ZN(n1146) );
XOR2_X1 U825 ( .A(n1152), .B(n1153), .Z(n1135) );
XNOR2_X1 U826 ( .A(n1154), .B(n1155), .ZN(n1134) );
XOR2_X1 U827 ( .A(KEYINPUT28), .B(G952), .Z(n1132) );
XOR2_X1 U828 ( .A(n1156), .B(n1157), .Z(G72) );
XOR2_X1 U829 ( .A(n1158), .B(n1159), .Z(n1157) );
AND2_X1 U830 ( .A1(n1102), .A2(n1160), .ZN(n1159) );
NOR2_X1 U831 ( .A1(n1161), .A2(n1162), .ZN(n1158) );
XOR2_X1 U832 ( .A(KEYINPUT39), .B(n1163), .Z(n1162) );
NOR2_X1 U833 ( .A1(G900), .A2(n1102), .ZN(n1163) );
XOR2_X1 U834 ( .A(n1164), .B(n1165), .Z(n1161) );
XNOR2_X1 U835 ( .A(n1166), .B(n1167), .ZN(n1165) );
XNOR2_X1 U836 ( .A(n1168), .B(n1169), .ZN(n1167) );
INV_X1 U837 ( .A(n1170), .ZN(n1166) );
XNOR2_X1 U838 ( .A(n1171), .B(n1172), .ZN(n1164) );
XNOR2_X1 U839 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n1171) );
NOR3_X1 U840 ( .A1(n1102), .A2(KEYINPUT31), .A3(n1173), .ZN(n1156) );
AND2_X1 U841 ( .A1(G227), .A2(G900), .ZN(n1173) );
NAND2_X1 U842 ( .A1(n1174), .A2(n1175), .ZN(G69) );
OR2_X1 U843 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U844 ( .A(n1178), .B(KEYINPUT46), .Z(n1174) );
NAND2_X1 U845 ( .A1(n1177), .A2(n1176), .ZN(n1178) );
NAND2_X1 U846 ( .A1(G953), .A2(n1179), .ZN(n1176) );
XOR2_X1 U847 ( .A(KEYINPUT12), .B(n1180), .Z(n1179) );
AND2_X1 U848 ( .A1(G224), .A2(G898), .ZN(n1180) );
XNOR2_X1 U849 ( .A(n1181), .B(n1182), .ZN(n1177) );
NOR3_X1 U850 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1182) );
NOR2_X1 U851 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NOR2_X1 U852 ( .A1(n1188), .A2(n1189), .ZN(n1184) );
XOR2_X1 U853 ( .A(n1187), .B(KEYINPUT59), .Z(n1189) );
XNOR2_X1 U854 ( .A(n1190), .B(KEYINPUT54), .ZN(n1187) );
NAND2_X1 U855 ( .A1(n1102), .A2(n1191), .ZN(n1181) );
NOR2_X1 U856 ( .A1(n1192), .A2(n1193), .ZN(G66) );
XOR2_X1 U857 ( .A(n1194), .B(n1195), .Z(n1193) );
NOR2_X1 U858 ( .A1(n1149), .A2(n1196), .ZN(n1194) );
NOR2_X1 U859 ( .A1(n1192), .A2(n1197), .ZN(G63) );
XOR2_X1 U860 ( .A(n1198), .B(n1199), .Z(n1197) );
NOR2_X1 U861 ( .A1(n1143), .A2(n1196), .ZN(n1198) );
NOR2_X1 U862 ( .A1(n1192), .A2(n1200), .ZN(G60) );
XOR2_X1 U863 ( .A(n1201), .B(n1202), .Z(n1200) );
XOR2_X1 U864 ( .A(KEYINPUT62), .B(n1203), .Z(n1202) );
AND2_X1 U865 ( .A1(G475), .A2(n1204), .ZN(n1203) );
NAND2_X1 U866 ( .A1(n1205), .A2(n1206), .ZN(G6) );
NAND2_X1 U867 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U868 ( .A(KEYINPUT29), .B(G104), .Z(n1208) );
XOR2_X1 U869 ( .A(n1209), .B(KEYINPUT32), .Z(n1207) );
NAND2_X1 U870 ( .A1(G104), .A2(n1210), .ZN(n1205) );
XNOR2_X1 U871 ( .A(KEYINPUT47), .B(n1209), .ZN(n1210) );
NAND2_X1 U872 ( .A1(n1211), .A2(n1212), .ZN(n1209) );
XOR2_X1 U873 ( .A(KEYINPUT3), .B(n1095), .Z(n1212) );
NOR2_X1 U874 ( .A1(n1192), .A2(n1213), .ZN(G57) );
XNOR2_X1 U875 ( .A(n1214), .B(n1215), .ZN(n1213) );
NOR2_X1 U876 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
XOR2_X1 U877 ( .A(n1218), .B(KEYINPUT25), .Z(n1217) );
NAND4_X1 U878 ( .A1(G902), .A2(G472), .A3(n1219), .A4(n1220), .ZN(n1218) );
XOR2_X1 U879 ( .A(KEYINPUT17), .B(n1090), .Z(n1220) );
NOR2_X1 U880 ( .A1(n1221), .A2(n1219), .ZN(n1216) );
XOR2_X1 U881 ( .A(n1222), .B(n1223), .Z(n1219) );
NOR3_X1 U882 ( .A1(n1155), .A2(n1224), .A3(n1225), .ZN(n1221) );
NOR2_X1 U883 ( .A1(KEYINPUT17), .A2(n1226), .ZN(n1225) );
AND2_X1 U884 ( .A1(G902), .A2(n1090), .ZN(n1226) );
AND2_X1 U885 ( .A1(n1196), .A2(KEYINPUT17), .ZN(n1224) );
INV_X1 U886 ( .A(G472), .ZN(n1155) );
NOR2_X1 U887 ( .A1(n1192), .A2(n1227), .ZN(G54) );
XOR2_X1 U888 ( .A(n1228), .B(n1229), .Z(n1227) );
XOR2_X1 U889 ( .A(n1230), .B(n1231), .Z(n1229) );
AND2_X1 U890 ( .A1(G469), .A2(n1204), .ZN(n1230) );
XNOR2_X1 U891 ( .A(G110), .B(n1232), .ZN(n1228) );
NAND2_X1 U892 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND2_X1 U893 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XOR2_X1 U894 ( .A(n1237), .B(KEYINPUT57), .Z(n1233) );
OR2_X1 U895 ( .A1(n1236), .A2(n1235), .ZN(n1237) );
XOR2_X1 U896 ( .A(n1170), .B(n1238), .Z(n1235) );
XNOR2_X1 U897 ( .A(G128), .B(n1239), .ZN(n1170) );
NOR2_X1 U898 ( .A1(n1192), .A2(n1240), .ZN(G51) );
XOR2_X1 U899 ( .A(n1241), .B(n1242), .Z(n1240) );
XOR2_X1 U900 ( .A(n1243), .B(n1244), .Z(n1242) );
XNOR2_X1 U901 ( .A(G125), .B(KEYINPUT36), .ZN(n1244) );
XNOR2_X1 U902 ( .A(n1245), .B(n1246), .ZN(n1241) );
XOR2_X1 U903 ( .A(n1247), .B(n1248), .Z(n1246) );
NOR2_X1 U904 ( .A1(KEYINPUT18), .A2(n1249), .ZN(n1248) );
NOR2_X1 U905 ( .A1(n1153), .A2(n1196), .ZN(n1247) );
INV_X1 U906 ( .A(n1204), .ZN(n1196) );
NOR2_X1 U907 ( .A1(n1250), .A2(n1090), .ZN(n1204) );
NOR2_X1 U908 ( .A1(n1191), .A2(n1160), .ZN(n1090) );
NAND4_X1 U909 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1160) );
AND4_X1 U910 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1254) );
NAND2_X1 U911 ( .A1(n1259), .A2(n1260), .ZN(n1253) );
NAND2_X1 U912 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
NAND4_X1 U913 ( .A1(n1116), .A2(n1263), .A3(n1264), .A4(n1265), .ZN(n1262) );
NAND2_X1 U914 ( .A1(n1266), .A2(n1267), .ZN(n1261) );
XOR2_X1 U915 ( .A(KEYINPUT2), .B(n1095), .Z(n1267) );
NAND3_X1 U916 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1251) );
OR2_X1 U917 ( .A1(n1271), .A2(KEYINPUT42), .ZN(n1269) );
NAND2_X1 U918 ( .A1(KEYINPUT42), .A2(n1272), .ZN(n1268) );
NAND2_X1 U919 ( .A1(n1259), .A2(n1115), .ZN(n1272) );
NAND4_X1 U920 ( .A1(n1273), .A2(n1274), .A3(n1275), .A4(n1276), .ZN(n1191) );
AND2_X1 U921 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
NAND2_X1 U922 ( .A1(n1211), .A2(n1279), .ZN(n1274) );
OR2_X1 U923 ( .A1(n1095), .A2(n1093), .ZN(n1279) );
INV_X1 U924 ( .A(n1083), .ZN(n1211) );
NAND4_X1 U925 ( .A1(n1263), .A2(n1117), .A3(n1280), .A4(n1281), .ZN(n1083) );
NAND2_X1 U926 ( .A1(n1263), .A2(n1282), .ZN(n1273) );
NAND3_X1 U927 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1282) );
XNOR2_X1 U928 ( .A(n1286), .B(KEYINPUT33), .ZN(n1285) );
NOR2_X1 U929 ( .A1(n1102), .A2(G952), .ZN(n1192) );
XNOR2_X1 U930 ( .A(G146), .B(n1287), .ZN(G48) );
NAND4_X1 U931 ( .A1(n1288), .A2(n1266), .A3(n1095), .A4(n1123), .ZN(n1287) );
XOR2_X1 U932 ( .A(n1289), .B(KEYINPUT35), .Z(n1288) );
XNOR2_X1 U933 ( .A(G143), .B(n1290), .ZN(G45) );
NAND3_X1 U934 ( .A1(n1291), .A2(n1259), .A3(n1292), .ZN(n1290) );
AND3_X1 U935 ( .A1(n1116), .A2(n1265), .A3(n1264), .ZN(n1292) );
XNOR2_X1 U936 ( .A(n1263), .B(KEYINPUT51), .ZN(n1291) );
XNOR2_X1 U937 ( .A(G140), .B(n1293), .ZN(G42) );
NAND2_X1 U938 ( .A1(n1271), .A2(n1270), .ZN(n1293) );
XNOR2_X1 U939 ( .A(n1294), .B(n1252), .ZN(G39) );
NAND4_X1 U940 ( .A1(n1271), .A2(n1103), .A3(n1295), .A4(n1113), .ZN(n1252) );
NAND2_X1 U941 ( .A1(KEYINPUT52), .A2(n1296), .ZN(n1294) );
XNOR2_X1 U942 ( .A(G134), .B(n1258), .ZN(G36) );
NAND3_X1 U943 ( .A1(n1116), .A2(n1093), .A3(n1271), .ZN(n1258) );
XNOR2_X1 U944 ( .A(G131), .B(n1257), .ZN(G33) );
NAND3_X1 U945 ( .A1(n1095), .A2(n1116), .A3(n1271), .ZN(n1257) );
AND2_X1 U946 ( .A1(n1096), .A2(n1259), .ZN(n1271) );
AND2_X1 U947 ( .A1(n1123), .A2(n1289), .ZN(n1259) );
INV_X1 U948 ( .A(n1115), .ZN(n1096) );
NAND2_X1 U949 ( .A1(n1297), .A2(n1127), .ZN(n1115) );
XNOR2_X1 U950 ( .A(G128), .B(n1256), .ZN(G30) );
NAND4_X1 U951 ( .A1(n1266), .A2(n1093), .A3(n1280), .A4(n1289), .ZN(n1256) );
XNOR2_X1 U952 ( .A(G101), .B(n1298), .ZN(G3) );
NAND2_X1 U953 ( .A1(n1263), .A2(n1299), .ZN(n1298) );
XNOR2_X1 U954 ( .A(KEYINPUT6), .B(n1283), .ZN(n1299) );
NAND2_X1 U955 ( .A1(n1300), .A2(n1116), .ZN(n1283) );
XNOR2_X1 U956 ( .A(G125), .B(n1255), .ZN(G27) );
NAND4_X1 U957 ( .A1(n1270), .A2(n1108), .A3(n1263), .A4(n1289), .ZN(n1255) );
NAND2_X1 U958 ( .A1(n1131), .A2(n1301), .ZN(n1289) );
NAND4_X1 U959 ( .A1(G902), .A2(G953), .A3(n1302), .A4(n1303), .ZN(n1301) );
INV_X1 U960 ( .A(G900), .ZN(n1303) );
AND3_X1 U961 ( .A1(n1114), .A2(n1113), .A3(n1095), .ZN(n1270) );
XOR2_X1 U962 ( .A(n1304), .B(n1305), .Z(G24) );
NOR2_X1 U963 ( .A1(G122), .A2(KEYINPUT23), .ZN(n1305) );
NAND2_X1 U964 ( .A1(n1286), .A2(n1263), .ZN(n1304) );
AND4_X1 U965 ( .A1(n1097), .A2(n1264), .A3(n1265), .A4(n1281), .ZN(n1286) );
AND2_X1 U966 ( .A1(n1108), .A2(n1117), .ZN(n1097) );
NOR2_X1 U967 ( .A1(n1113), .A2(n1295), .ZN(n1117) );
XNOR2_X1 U968 ( .A(G119), .B(n1276), .ZN(G21) );
NAND4_X1 U969 ( .A1(n1103), .A2(n1266), .A3(n1108), .A4(n1281), .ZN(n1276) );
AND3_X1 U970 ( .A1(n1295), .A2(n1113), .A3(n1263), .ZN(n1266) );
XNOR2_X1 U971 ( .A(G116), .B(n1278), .ZN(G18) );
NAND2_X1 U972 ( .A1(n1306), .A2(n1093), .ZN(n1278) );
INV_X1 U973 ( .A(n1084), .ZN(n1093) );
NAND2_X1 U974 ( .A1(n1307), .A2(n1265), .ZN(n1084) );
XNOR2_X1 U975 ( .A(n1264), .B(KEYINPUT56), .ZN(n1307) );
XOR2_X1 U976 ( .A(n1277), .B(n1308), .Z(G15) );
XNOR2_X1 U977 ( .A(KEYINPUT44), .B(n1309), .ZN(n1308) );
NAND2_X1 U978 ( .A1(n1095), .A2(n1306), .ZN(n1277) );
AND4_X1 U979 ( .A1(n1116), .A2(n1108), .A3(n1263), .A4(n1281), .ZN(n1306) );
NOR2_X1 U980 ( .A1(n1310), .A2(n1121), .ZN(n1108) );
NOR2_X1 U981 ( .A1(n1113), .A2(n1114), .ZN(n1116) );
NOR2_X1 U982 ( .A1(n1265), .A2(n1311), .ZN(n1095) );
INV_X1 U983 ( .A(n1264), .ZN(n1311) );
NAND2_X1 U984 ( .A1(n1312), .A2(n1313), .ZN(G12) );
NAND3_X1 U985 ( .A1(n1314), .A2(n1315), .A3(n1316), .ZN(n1313) );
INV_X1 U986 ( .A(G110), .ZN(n1315) );
XOR2_X1 U987 ( .A(n1317), .B(KEYINPUT11), .Z(n1312) );
NAND2_X1 U988 ( .A1(G110), .A2(n1318), .ZN(n1317) );
NAND2_X1 U989 ( .A1(n1316), .A2(n1314), .ZN(n1318) );
XNOR2_X1 U990 ( .A(n1263), .B(KEYINPUT5), .ZN(n1314) );
INV_X1 U991 ( .A(n1125), .ZN(n1263) );
NAND2_X1 U992 ( .A1(n1128), .A2(n1127), .ZN(n1125) );
NAND2_X1 U993 ( .A1(G214), .A2(n1319), .ZN(n1127) );
INV_X1 U994 ( .A(n1297), .ZN(n1128) );
XNOR2_X1 U995 ( .A(n1320), .B(n1153), .ZN(n1297) );
NAND2_X1 U996 ( .A1(G210), .A2(n1319), .ZN(n1153) );
NAND2_X1 U997 ( .A1(n1250), .A2(n1321), .ZN(n1319) );
INV_X1 U998 ( .A(G237), .ZN(n1321) );
NAND2_X1 U999 ( .A1(KEYINPUT16), .A2(n1152), .ZN(n1320) );
AND2_X1 U1000 ( .A1(n1322), .A2(n1250), .ZN(n1152) );
XOR2_X1 U1001 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1002 ( .A(n1243), .B(n1249), .Z(n1324) );
NAND2_X1 U1003 ( .A1(G224), .A2(n1102), .ZN(n1249) );
NAND2_X1 U1004 ( .A1(n1325), .A2(n1326), .ZN(n1243) );
NAND2_X1 U1005 ( .A1(n1327), .A2(n1188), .ZN(n1326) );
INV_X1 U1006 ( .A(n1190), .ZN(n1327) );
XOR2_X1 U1007 ( .A(n1328), .B(KEYINPUT38), .Z(n1325) );
NAND2_X1 U1008 ( .A1(n1186), .A2(n1190), .ZN(n1328) );
XOR2_X1 U1009 ( .A(n1223), .B(n1329), .Z(n1190) );
XOR2_X1 U1010 ( .A(n1330), .B(n1331), .Z(n1329) );
NOR2_X1 U1011 ( .A1(G101), .A2(KEYINPUT30), .ZN(n1331) );
NOR2_X1 U1012 ( .A1(n1332), .A2(n1333), .ZN(n1330) );
XOR2_X1 U1013 ( .A(KEYINPUT37), .B(n1334), .Z(n1333) );
NOR2_X1 U1014 ( .A1(G104), .A2(n1335), .ZN(n1334) );
AND2_X1 U1015 ( .A1(n1335), .A2(G104), .ZN(n1332) );
XOR2_X1 U1016 ( .A(G107), .B(KEYINPUT20), .Z(n1335) );
INV_X1 U1017 ( .A(n1188), .ZN(n1186) );
XOR2_X1 U1018 ( .A(G110), .B(G122), .Z(n1188) );
XNOR2_X1 U1019 ( .A(KEYINPUT14), .B(n1336), .ZN(n1323) );
NOR2_X1 U1020 ( .A1(KEYINPUT10), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1021 ( .A(n1338), .B(n1245), .Z(n1337) );
NOR2_X1 U1022 ( .A1(G125), .A2(KEYINPUT0), .ZN(n1338) );
INV_X1 U1023 ( .A(n1284), .ZN(n1316) );
NAND3_X1 U1024 ( .A1(n1114), .A2(n1113), .A3(n1300), .ZN(n1284) );
AND3_X1 U1025 ( .A1(n1280), .A2(n1281), .A3(n1103), .ZN(n1300) );
NOR2_X1 U1026 ( .A1(n1265), .A2(n1264), .ZN(n1103) );
XOR2_X1 U1027 ( .A(n1339), .B(n1151), .Z(n1264) );
NAND2_X1 U1028 ( .A1(n1201), .A2(n1250), .ZN(n1151) );
XNOR2_X1 U1029 ( .A(n1340), .B(n1341), .ZN(n1201) );
NOR2_X1 U1030 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
XOR2_X1 U1031 ( .A(n1344), .B(KEYINPUT4), .Z(n1343) );
NAND2_X1 U1032 ( .A1(G122), .A2(n1309), .ZN(n1344) );
NOR2_X1 U1033 ( .A1(G122), .A2(n1309), .ZN(n1342) );
INV_X1 U1034 ( .A(G113), .ZN(n1309) );
XOR2_X1 U1035 ( .A(n1345), .B(G104), .Z(n1340) );
NAND2_X1 U1036 ( .A1(KEYINPUT34), .A2(n1346), .ZN(n1345) );
XOR2_X1 U1037 ( .A(n1347), .B(n1348), .Z(n1346) );
XNOR2_X1 U1038 ( .A(n1349), .B(G131), .ZN(n1348) );
XOR2_X1 U1039 ( .A(n1350), .B(n1351), .Z(n1347) );
AND2_X1 U1040 ( .A1(n1352), .A2(G214), .ZN(n1351) );
NAND2_X1 U1041 ( .A1(n1353), .A2(n1354), .ZN(n1350) );
NAND2_X1 U1042 ( .A1(G146), .A2(n1355), .ZN(n1354) );
NAND2_X1 U1043 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
XNOR2_X1 U1044 ( .A(n1358), .B(KEYINPUT19), .ZN(n1356) );
NAND2_X1 U1045 ( .A1(n1359), .A2(n1360), .ZN(n1353) );
NAND2_X1 U1046 ( .A1(n1361), .A2(n1362), .ZN(n1359) );
OR2_X1 U1047 ( .A1(n1168), .A2(KEYINPUT19), .ZN(n1362) );
NAND2_X1 U1048 ( .A1(n1358), .A2(KEYINPUT19), .ZN(n1361) );
NAND2_X1 U1049 ( .A1(KEYINPUT61), .A2(G475), .ZN(n1339) );
XNOR2_X1 U1050 ( .A(n1141), .B(n1143), .ZN(n1265) );
INV_X1 U1051 ( .A(G478), .ZN(n1143) );
NOR2_X1 U1052 ( .A1(n1199), .A2(G902), .ZN(n1141) );
XNOR2_X1 U1053 ( .A(n1363), .B(n1364), .ZN(n1199) );
XNOR2_X1 U1054 ( .A(n1365), .B(n1366), .ZN(n1364) );
NAND2_X1 U1055 ( .A1(KEYINPUT50), .A2(n1367), .ZN(n1365) );
INV_X1 U1056 ( .A(G134), .ZN(n1367) );
XOR2_X1 U1057 ( .A(n1368), .B(n1369), .Z(n1363) );
AND2_X1 U1058 ( .A1(n1370), .A2(G217), .ZN(n1369) );
NAND2_X1 U1059 ( .A1(n1371), .A2(KEYINPUT48), .ZN(n1368) );
XOR2_X1 U1060 ( .A(n1372), .B(n1373), .Z(n1371) );
NOR2_X1 U1061 ( .A1(KEYINPUT58), .A2(G107), .ZN(n1373) );
XNOR2_X1 U1062 ( .A(G116), .B(G122), .ZN(n1372) );
NAND2_X1 U1063 ( .A1(n1131), .A2(n1374), .ZN(n1281) );
NAND3_X1 U1064 ( .A1(n1183), .A2(n1302), .A3(G902), .ZN(n1374) );
NOR2_X1 U1065 ( .A1(n1102), .A2(G898), .ZN(n1183) );
NAND3_X1 U1066 ( .A1(n1302), .A2(n1102), .A3(G952), .ZN(n1131) );
NAND2_X1 U1067 ( .A1(G237), .A2(G234), .ZN(n1302) );
XNOR2_X1 U1068 ( .A(n1123), .B(KEYINPUT15), .ZN(n1280) );
NOR2_X1 U1069 ( .A1(n1122), .A2(n1121), .ZN(n1123) );
INV_X1 U1070 ( .A(n1145), .ZN(n1121) );
NAND2_X1 U1071 ( .A1(G221), .A2(n1375), .ZN(n1145) );
INV_X1 U1072 ( .A(n1310), .ZN(n1122) );
XOR2_X1 U1073 ( .A(n1139), .B(KEYINPUT53), .Z(n1310) );
XNOR2_X1 U1074 ( .A(n1376), .B(G469), .ZN(n1139) );
NAND2_X1 U1075 ( .A1(n1377), .A2(n1250), .ZN(n1376) );
XOR2_X1 U1076 ( .A(n1378), .B(n1379), .Z(n1377) );
XNOR2_X1 U1077 ( .A(n1238), .B(n1239), .ZN(n1379) );
NAND2_X1 U1078 ( .A1(n1380), .A2(n1381), .ZN(n1239) );
NAND2_X1 U1079 ( .A1(n1382), .A2(n1383), .ZN(n1381) );
INV_X1 U1080 ( .A(KEYINPUT27), .ZN(n1383) );
XNOR2_X1 U1081 ( .A(G143), .B(G146), .ZN(n1382) );
NAND3_X1 U1082 ( .A1(G143), .A2(n1360), .A3(KEYINPUT27), .ZN(n1380) );
INV_X1 U1083 ( .A(G146), .ZN(n1360) );
XNOR2_X1 U1084 ( .A(n1384), .B(n1385), .ZN(n1238) );
XOR2_X1 U1085 ( .A(G104), .B(G101), .Z(n1385) );
NAND2_X1 U1086 ( .A1(KEYINPUT55), .A2(n1081), .ZN(n1384) );
INV_X1 U1087 ( .A(G107), .ZN(n1081) );
XOR2_X1 U1088 ( .A(n1386), .B(n1387), .Z(n1378) );
XOR2_X1 U1089 ( .A(n1236), .B(n1231), .Z(n1387) );
XNOR2_X1 U1090 ( .A(n1388), .B(n1389), .ZN(n1231) );
XNOR2_X1 U1091 ( .A(KEYINPUT1), .B(n1390), .ZN(n1389) );
INV_X1 U1092 ( .A(G140), .ZN(n1390) );
NAND2_X1 U1093 ( .A1(G227), .A2(n1102), .ZN(n1388) );
NAND3_X1 U1094 ( .A1(n1391), .A2(n1392), .A3(n1144), .ZN(n1113) );
NAND2_X1 U1095 ( .A1(n1150), .A2(n1149), .ZN(n1144) );
NAND2_X1 U1096 ( .A1(n1149), .A2(n1393), .ZN(n1392) );
OR3_X1 U1097 ( .A1(n1149), .A2(n1150), .A3(n1393), .ZN(n1391) );
INV_X1 U1098 ( .A(KEYINPUT8), .ZN(n1393) );
NOR2_X1 U1099 ( .A1(n1195), .A2(G902), .ZN(n1150) );
XNOR2_X1 U1100 ( .A(n1394), .B(n1395), .ZN(n1195) );
XOR2_X1 U1101 ( .A(n1168), .B(n1396), .Z(n1395) );
XNOR2_X1 U1102 ( .A(G119), .B(G146), .ZN(n1396) );
NAND2_X1 U1103 ( .A1(n1357), .A2(n1397), .ZN(n1168) );
INV_X1 U1104 ( .A(n1358), .ZN(n1397) );
NOR2_X1 U1105 ( .A1(n1398), .A2(G140), .ZN(n1358) );
NAND2_X1 U1106 ( .A1(G140), .A2(n1398), .ZN(n1357) );
INV_X1 U1107 ( .A(G125), .ZN(n1398) );
XOR2_X1 U1108 ( .A(n1386), .B(n1399), .Z(n1394) );
NOR2_X1 U1109 ( .A1(KEYINPUT45), .A2(n1400), .ZN(n1399) );
XNOR2_X1 U1110 ( .A(n1401), .B(n1296), .ZN(n1400) );
NAND2_X1 U1111 ( .A1(G221), .A2(n1370), .ZN(n1401) );
AND2_X1 U1112 ( .A1(G234), .A2(n1102), .ZN(n1370) );
INV_X1 U1113 ( .A(G953), .ZN(n1102) );
XNOR2_X1 U1114 ( .A(G110), .B(G128), .ZN(n1386) );
NAND2_X1 U1115 ( .A1(G217), .A2(n1375), .ZN(n1149) );
NAND2_X1 U1116 ( .A1(G234), .A2(n1250), .ZN(n1375) );
INV_X1 U1117 ( .A(n1295), .ZN(n1114) );
XOR2_X1 U1118 ( .A(n1402), .B(n1154), .Z(n1295) );
NAND2_X1 U1119 ( .A1(n1403), .A2(n1250), .ZN(n1154) );
INV_X1 U1120 ( .A(G902), .ZN(n1250) );
XOR2_X1 U1121 ( .A(n1404), .B(n1405), .Z(n1403) );
XNOR2_X1 U1122 ( .A(n1406), .B(n1223), .ZN(n1405) );
XOR2_X1 U1123 ( .A(G113), .B(n1407), .Z(n1223) );
XOR2_X1 U1124 ( .A(G119), .B(G116), .Z(n1407) );
INV_X1 U1125 ( .A(n1214), .ZN(n1406) );
XNOR2_X1 U1126 ( .A(n1408), .B(G101), .ZN(n1214) );
NAND2_X1 U1127 ( .A1(G210), .A2(n1352), .ZN(n1408) );
NOR2_X1 U1128 ( .A1(G953), .A2(G237), .ZN(n1352) );
XNOR2_X1 U1129 ( .A(KEYINPUT13), .B(n1409), .ZN(n1404) );
NOR2_X1 U1130 ( .A1(KEYINPUT26), .A2(n1222), .ZN(n1409) );
XNOR2_X1 U1131 ( .A(n1236), .B(n1245), .ZN(n1222) );
XOR2_X1 U1132 ( .A(G146), .B(n1366), .Z(n1245) );
XNOR2_X1 U1133 ( .A(G128), .B(n1349), .ZN(n1366) );
INV_X1 U1134 ( .A(G143), .ZN(n1349) );
NAND3_X1 U1135 ( .A1(n1410), .A2(n1411), .A3(n1412), .ZN(n1236) );
NAND2_X1 U1136 ( .A1(n1413), .A2(n1172), .ZN(n1412) );
NAND2_X1 U1137 ( .A1(KEYINPUT43), .A2(n1414), .ZN(n1411) );
NAND2_X1 U1138 ( .A1(n1415), .A2(n1169), .ZN(n1414) );
XNOR2_X1 U1139 ( .A(KEYINPUT21), .B(n1172), .ZN(n1415) );
NAND2_X1 U1140 ( .A1(n1416), .A2(n1417), .ZN(n1410) );
INV_X1 U1141 ( .A(KEYINPUT43), .ZN(n1417) );
NAND2_X1 U1142 ( .A1(n1418), .A2(n1419), .ZN(n1416) );
OR3_X1 U1143 ( .A1(n1172), .A2(n1413), .A3(KEYINPUT21), .ZN(n1419) );
INV_X1 U1144 ( .A(n1169), .ZN(n1413) );
XNOR2_X1 U1145 ( .A(G134), .B(n1296), .ZN(n1169) );
INV_X1 U1146 ( .A(G137), .ZN(n1296) );
NAND2_X1 U1147 ( .A1(KEYINPUT21), .A2(n1172), .ZN(n1418) );
INV_X1 U1148 ( .A(G131), .ZN(n1172) );
NAND2_X1 U1149 ( .A1(n1420), .A2(KEYINPUT40), .ZN(n1402) );
XNOR2_X1 U1150 ( .A(G472), .B(KEYINPUT41), .ZN(n1420) );
endmodule


