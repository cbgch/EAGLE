//Key = 0000110000011101111111000001011110011010110010100101111100110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272;

XOR2_X1 U704 ( .A(G107), .B(n969), .Z(G9) );
NOR2_X1 U705 ( .A1(n970), .A2(n971), .ZN(n969) );
XOR2_X1 U706 ( .A(n972), .B(KEYINPUT33), .Z(n970) );
NOR2_X1 U707 ( .A1(n973), .A2(n974), .ZN(G75) );
NOR4_X1 U708 ( .A1(n975), .A2(n976), .A3(n977), .A4(n978), .ZN(n974) );
NAND4_X1 U709 ( .A1(n979), .A2(n980), .A3(n981), .A4(n982), .ZN(n975) );
NAND3_X1 U710 ( .A1(n983), .A2(n984), .A3(n985), .ZN(n980) );
NAND2_X1 U711 ( .A1(n986), .A2(n987), .ZN(n984) );
NAND2_X1 U712 ( .A1(n988), .A2(n989), .ZN(n986) );
NAND2_X1 U713 ( .A1(n990), .A2(n991), .ZN(n989) );
NAND3_X1 U714 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
OR2_X1 U715 ( .A1(n995), .A2(n996), .ZN(n993) );
NAND2_X1 U716 ( .A1(n997), .A2(n998), .ZN(n990) );
NAND2_X1 U717 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND2_X1 U718 ( .A1(n992), .A2(n1001), .ZN(n1000) );
NAND2_X1 U719 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NAND2_X1 U720 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NAND2_X1 U721 ( .A1(n994), .A2(n1006), .ZN(n999) );
NAND2_X1 U722 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND2_X1 U723 ( .A1(n1009), .A2(n1010), .ZN(n983) );
XOR2_X1 U724 ( .A(n1011), .B(KEYINPUT22), .Z(n1010) );
OR2_X1 U725 ( .A1(n1011), .A2(n971), .ZN(n979) );
NAND4_X1 U726 ( .A1(n988), .A2(n994), .A3(n997), .A4(n992), .ZN(n1011) );
INV_X1 U727 ( .A(n1012), .ZN(n988) );
NOR3_X1 U728 ( .A1(n1013), .A2(G953), .A3(G952), .ZN(n973) );
INV_X1 U729 ( .A(n981), .ZN(n1013) );
NAND4_X1 U730 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n981) );
NOR4_X1 U731 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
XNOR2_X1 U732 ( .A(G475), .B(n1022), .ZN(n1021) );
XNOR2_X1 U733 ( .A(n1023), .B(n1024), .ZN(n1020) );
XNOR2_X1 U734 ( .A(n1025), .B(n1026), .ZN(n1019) );
NOR3_X1 U735 ( .A1(n1027), .A2(n1009), .A3(n1004), .ZN(n1016) );
XOR2_X1 U736 ( .A(n1028), .B(n1029), .Z(n1015) );
NAND2_X1 U737 ( .A1(n1030), .A2(KEYINPUT55), .ZN(n1029) );
XNOR2_X1 U738 ( .A(G478), .B(KEYINPUT26), .ZN(n1030) );
XOR2_X1 U739 ( .A(KEYINPUT31), .B(n1031), .Z(n1014) );
XOR2_X1 U740 ( .A(n1032), .B(n1033), .Z(G72) );
XOR2_X1 U741 ( .A(n1034), .B(n1035), .Z(n1033) );
NOR2_X1 U742 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
XOR2_X1 U743 ( .A(n1038), .B(n1039), .Z(n1037) );
XNOR2_X1 U744 ( .A(n1040), .B(n1041), .ZN(n1039) );
XOR2_X1 U745 ( .A(n1042), .B(n1043), .Z(n1038) );
XOR2_X1 U746 ( .A(KEYINPUT45), .B(KEYINPUT27), .Z(n1043) );
NAND2_X1 U747 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
OR2_X1 U748 ( .A1(n1046), .A2(G131), .ZN(n1045) );
XOR2_X1 U749 ( .A(n1047), .B(KEYINPUT24), .Z(n1044) );
NAND2_X1 U750 ( .A1(G131), .A2(n1046), .ZN(n1047) );
NOR2_X1 U751 ( .A1(G900), .A2(n982), .ZN(n1036) );
NAND2_X1 U752 ( .A1(n982), .A2(n1048), .ZN(n1034) );
NAND2_X1 U753 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
INV_X1 U754 ( .A(n976), .ZN(n1049) );
NAND2_X1 U755 ( .A1(G953), .A2(n1051), .ZN(n1032) );
NAND2_X1 U756 ( .A1(G900), .A2(G227), .ZN(n1051) );
XOR2_X1 U757 ( .A(n1052), .B(n1053), .Z(G69) );
NAND2_X1 U758 ( .A1(G953), .A2(n1054), .ZN(n1053) );
NAND2_X1 U759 ( .A1(G898), .A2(G224), .ZN(n1054) );
NAND2_X1 U760 ( .A1(KEYINPUT16), .A2(n1055), .ZN(n1052) );
XOR2_X1 U761 ( .A(n1056), .B(n1057), .Z(n1055) );
NAND2_X1 U762 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U763 ( .A1(n1060), .A2(G953), .ZN(n1059) );
XOR2_X1 U764 ( .A(n1061), .B(n1062), .Z(n1058) );
NAND2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(n1056) );
XNOR2_X1 U766 ( .A(KEYINPUT52), .B(n977), .ZN(n1064) );
XNOR2_X1 U767 ( .A(KEYINPUT59), .B(n982), .ZN(n1063) );
NOR2_X1 U768 ( .A1(n1065), .A2(n1066), .ZN(G66) );
XOR2_X1 U769 ( .A(n1067), .B(n1068), .Z(n1066) );
NOR3_X1 U770 ( .A1(n1069), .A2(KEYINPUT43), .A3(n1070), .ZN(n1068) );
NOR2_X1 U771 ( .A1(n1065), .A2(n1071), .ZN(G63) );
XNOR2_X1 U772 ( .A(n1072), .B(n1073), .ZN(n1071) );
XOR2_X1 U773 ( .A(KEYINPUT57), .B(n1074), .Z(n1073) );
NOR2_X1 U774 ( .A1(n1075), .A2(n1069), .ZN(n1074) );
NOR2_X1 U775 ( .A1(n1065), .A2(n1076), .ZN(G60) );
XOR2_X1 U776 ( .A(n1077), .B(n1078), .Z(n1076) );
XOR2_X1 U777 ( .A(KEYINPUT29), .B(n1079), .Z(n1078) );
NOR2_X1 U778 ( .A1(n1080), .A2(n1069), .ZN(n1079) );
INV_X1 U779 ( .A(G475), .ZN(n1080) );
XNOR2_X1 U780 ( .A(G104), .B(n1081), .ZN(G6) );
NOR2_X1 U781 ( .A1(n1065), .A2(n1082), .ZN(G57) );
NOR3_X1 U782 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
NOR2_X1 U783 ( .A1(G101), .A2(n1086), .ZN(n1085) );
XNOR2_X1 U784 ( .A(n1087), .B(n1088), .ZN(n1086) );
NOR3_X1 U785 ( .A1(n1089), .A2(n1087), .A3(n1088), .ZN(n1084) );
AND2_X1 U786 ( .A1(n1088), .A2(n1090), .ZN(n1083) );
XNOR2_X1 U787 ( .A(n1091), .B(n1092), .ZN(n1088) );
NOR2_X1 U788 ( .A1(n1025), .A2(n1069), .ZN(n1092) );
NOR2_X1 U789 ( .A1(n1065), .A2(n1093), .ZN(G54) );
XOR2_X1 U790 ( .A(n1094), .B(n1095), .Z(n1093) );
XOR2_X1 U791 ( .A(n1096), .B(n1097), .Z(n1095) );
XNOR2_X1 U792 ( .A(n1098), .B(n1099), .ZN(n1097) );
XOR2_X1 U793 ( .A(n1100), .B(n1101), .Z(n1094) );
XNOR2_X1 U794 ( .A(n1102), .B(n1103), .ZN(n1101) );
NOR2_X1 U795 ( .A1(n1104), .A2(n1069), .ZN(n1103) );
INV_X1 U796 ( .A(G469), .ZN(n1104) );
XNOR2_X1 U797 ( .A(KEYINPUT11), .B(n1105), .ZN(n1100) );
NOR2_X1 U798 ( .A1(n1065), .A2(n1106), .ZN(G51) );
XOR2_X1 U799 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U800 ( .A(n1109), .B(n1110), .Z(n1107) );
NOR2_X1 U801 ( .A1(n1111), .A2(n1069), .ZN(n1110) );
NAND2_X1 U802 ( .A1(G902), .A2(n1112), .ZN(n1069) );
OR3_X1 U803 ( .A1(n978), .A2(n977), .A3(n976), .ZN(n1112) );
NAND4_X1 U804 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n976) );
NOR4_X1 U805 ( .A1(n1117), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1116) );
INV_X1 U806 ( .A(n1121), .ZN(n1117) );
NAND2_X1 U807 ( .A1(n1122), .A2(n1123), .ZN(n1115) );
INV_X1 U808 ( .A(n1124), .ZN(n1123) );
XNOR2_X1 U809 ( .A(n1125), .B(KEYINPUT44), .ZN(n1122) );
NAND4_X1 U810 ( .A1(n1081), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n977) );
AND4_X1 U811 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1128) );
NOR3_X1 U812 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1127) );
NOR2_X1 U813 ( .A1(n971), .A2(n972), .ZN(n1135) );
NAND3_X1 U814 ( .A1(n996), .A2(n992), .A3(n1136), .ZN(n972) );
NOR4_X1 U815 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1134) );
NAND2_X1 U816 ( .A1(KEYINPUT23), .A2(n1141), .ZN(n1138) );
NOR2_X1 U817 ( .A1(KEYINPUT23), .A2(n1142), .ZN(n1133) );
INV_X1 U818 ( .A(n1143), .ZN(n1142) );
NAND4_X1 U819 ( .A1(n995), .A2(n1137), .A3(n1136), .A4(n992), .ZN(n1081) );
XNOR2_X1 U820 ( .A(n1050), .B(KEYINPUT34), .ZN(n978) );
INV_X1 U821 ( .A(G210), .ZN(n1111) );
NAND3_X1 U822 ( .A1(KEYINPUT49), .A2(n1144), .A3(n1145), .ZN(n1109) );
XOR2_X1 U823 ( .A(n1146), .B(KEYINPUT48), .Z(n1145) );
NAND2_X1 U824 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U825 ( .A(n1149), .B(n1150), .Z(n1148) );
INV_X1 U826 ( .A(n1151), .ZN(n1147) );
NAND2_X1 U827 ( .A1(n1152), .A2(n1151), .ZN(n1144) );
XNOR2_X1 U828 ( .A(n1150), .B(n1149), .ZN(n1152) );
NAND2_X1 U829 ( .A1(KEYINPUT51), .A2(G125), .ZN(n1149) );
XOR2_X1 U830 ( .A(n1153), .B(KEYINPUT38), .Z(n1150) );
NOR2_X1 U831 ( .A1(n982), .A2(G952), .ZN(n1065) );
XOR2_X1 U832 ( .A(n1113), .B(n1154), .Z(G48) );
NAND2_X1 U833 ( .A1(KEYINPUT15), .A2(G146), .ZN(n1154) );
NAND4_X1 U834 ( .A1(n995), .A2(n1155), .A3(n1125), .A4(n1156), .ZN(n1113) );
XOR2_X1 U835 ( .A(n1157), .B(n1158), .Z(G45) );
NOR2_X1 U836 ( .A1(KEYINPUT9), .A2(n1159), .ZN(n1158) );
NOR2_X1 U837 ( .A1(n1002), .A2(n1124), .ZN(n1159) );
NAND4_X1 U838 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1124) );
NOR2_X1 U839 ( .A1(n971), .A2(n1007), .ZN(n1163) );
INV_X1 U840 ( .A(n1164), .ZN(n1007) );
XNOR2_X1 U841 ( .A(G143), .B(KEYINPUT39), .ZN(n1157) );
XOR2_X1 U842 ( .A(n1114), .B(n1165), .Z(G42) );
NAND2_X1 U843 ( .A1(KEYINPUT46), .A2(G140), .ZN(n1165) );
NAND3_X1 U844 ( .A1(n995), .A2(n1166), .A3(n1141), .ZN(n1114) );
INV_X1 U845 ( .A(n1008), .ZN(n1141) );
XOR2_X1 U846 ( .A(G137), .B(n1120), .Z(G39) );
AND2_X1 U847 ( .A1(n1167), .A2(n1166), .ZN(n1120) );
XNOR2_X1 U848 ( .A(n1168), .B(n1119), .ZN(G36) );
AND3_X1 U849 ( .A1(n1164), .A2(n996), .A3(n1166), .ZN(n1119) );
XNOR2_X1 U850 ( .A(n1118), .B(n1169), .ZN(G33) );
NAND2_X1 U851 ( .A1(KEYINPUT36), .A2(G131), .ZN(n1169) );
AND3_X1 U852 ( .A1(n1166), .A2(n1164), .A3(n995), .ZN(n1118) );
AND4_X1 U853 ( .A1(n1125), .A2(n985), .A3(n987), .A4(n1161), .ZN(n1166) );
XNOR2_X1 U854 ( .A(G128), .B(n1121), .ZN(G30) );
NAND4_X1 U855 ( .A1(n1155), .A2(n996), .A3(n1170), .A4(n1156), .ZN(n1121) );
XNOR2_X1 U856 ( .A(G101), .B(n1126), .ZN(G3) );
NAND4_X1 U857 ( .A1(n997), .A2(n1164), .A3(n1137), .A4(n1136), .ZN(n1126) );
INV_X1 U858 ( .A(n1139), .ZN(n1136) );
XNOR2_X1 U859 ( .A(G125), .B(n1050), .ZN(G27) );
NAND4_X1 U860 ( .A1(n994), .A2(n995), .A3(n1171), .A4(n1155), .ZN(n1050) );
AND3_X1 U861 ( .A1(n1018), .A2(n1161), .A3(n1137), .ZN(n1155) );
NAND2_X1 U862 ( .A1(n1172), .A2(n1012), .ZN(n1161) );
NAND2_X1 U863 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
INV_X1 U864 ( .A(G900), .ZN(n1174) );
XNOR2_X1 U865 ( .A(G122), .B(n1132), .ZN(G24) );
NAND4_X1 U866 ( .A1(n1175), .A2(n992), .A3(n1162), .A4(n1160), .ZN(n1132) );
NOR2_X1 U867 ( .A1(n1018), .A2(n1156), .ZN(n992) );
XNOR2_X1 U868 ( .A(G119), .B(n1131), .ZN(G21) );
NAND2_X1 U869 ( .A1(n1175), .A2(n1167), .ZN(n1131) );
AND3_X1 U870 ( .A1(n1156), .A2(n1018), .A3(n997), .ZN(n1167) );
XNOR2_X1 U871 ( .A(G116), .B(n1130), .ZN(G18) );
NAND3_X1 U872 ( .A1(n1164), .A2(n996), .A3(n1175), .ZN(n1130) );
NOR2_X1 U873 ( .A1(n1176), .A2(n1177), .ZN(n996) );
XNOR2_X1 U874 ( .A(G113), .B(n1129), .ZN(G15) );
NAND3_X1 U875 ( .A1(n995), .A2(n1164), .A3(n1175), .ZN(n1129) );
AND3_X1 U876 ( .A1(n1137), .A2(n1178), .A3(n994), .ZN(n1175) );
AND2_X1 U877 ( .A1(n1005), .A2(n1179), .ZN(n994) );
NOR2_X1 U878 ( .A1(n1018), .A2(n1171), .ZN(n1164) );
AND2_X1 U879 ( .A1(n1176), .A2(n1162), .ZN(n995) );
XNOR2_X1 U880 ( .A(n1177), .B(KEYINPUT54), .ZN(n1162) );
INV_X1 U881 ( .A(n1160), .ZN(n1176) );
NAND2_X1 U882 ( .A1(n1180), .A2(n1181), .ZN(G12) );
NAND2_X1 U883 ( .A1(n1143), .A2(n1105), .ZN(n1181) );
XOR2_X1 U884 ( .A(KEYINPUT40), .B(n1182), .Z(n1180) );
NOR2_X1 U885 ( .A1(n1143), .A2(n1105), .ZN(n1182) );
NOR4_X1 U886 ( .A1(n1008), .A2(n1140), .A3(n971), .A4(n1139), .ZN(n1143) );
NAND2_X1 U887 ( .A1(n1170), .A2(n1178), .ZN(n1139) );
NAND2_X1 U888 ( .A1(n1012), .A2(n1183), .ZN(n1178) );
NAND2_X1 U889 ( .A1(n1060), .A2(n1173), .ZN(n1183) );
AND3_X1 U890 ( .A1(G953), .A2(n1184), .A3(n1185), .ZN(n1173) );
XNOR2_X1 U891 ( .A(G902), .B(KEYINPUT21), .ZN(n1185) );
XNOR2_X1 U892 ( .A(G898), .B(KEYINPUT47), .ZN(n1060) );
NAND3_X1 U893 ( .A1(n1184), .A2(n982), .A3(G952), .ZN(n1012) );
NAND2_X1 U894 ( .A1(G237), .A2(G234), .ZN(n1184) );
XNOR2_X1 U895 ( .A(KEYINPUT62), .B(n1002), .ZN(n1170) );
INV_X1 U896 ( .A(n1125), .ZN(n1002) );
NOR2_X1 U897 ( .A1(n1004), .A2(n1005), .ZN(n1125) );
NOR2_X1 U898 ( .A1(n1031), .A2(n1027), .ZN(n1005) );
AND2_X1 U899 ( .A1(n1186), .A2(G469), .ZN(n1027) );
NOR2_X1 U900 ( .A1(n1186), .A2(G469), .ZN(n1031) );
NAND2_X1 U901 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U902 ( .A(n1098), .B(n1189), .Z(n1187) );
XNOR2_X1 U903 ( .A(n1190), .B(n1191), .ZN(n1189) );
NAND2_X1 U904 ( .A1(KEYINPUT5), .A2(n1099), .ZN(n1191) );
NAND2_X1 U905 ( .A1(KEYINPUT32), .A2(n1192), .ZN(n1190) );
XOR2_X1 U906 ( .A(n1102), .B(n1193), .Z(n1192) );
NAND2_X1 U907 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
OR2_X1 U908 ( .A1(n1196), .A2(n1096), .ZN(n1195) );
XOR2_X1 U909 ( .A(n1197), .B(KEYINPUT56), .Z(n1194) );
NAND2_X1 U910 ( .A1(n1096), .A2(n1196), .ZN(n1197) );
XOR2_X1 U911 ( .A(G110), .B(KEYINPUT1), .Z(n1196) );
XNOR2_X1 U912 ( .A(G140), .B(KEYINPUT63), .ZN(n1096) );
NAND2_X1 U913 ( .A1(G227), .A2(n982), .ZN(n1102) );
XNOR2_X1 U914 ( .A(n1040), .B(n1198), .ZN(n1098) );
XNOR2_X1 U915 ( .A(n1089), .B(n1199), .ZN(n1198) );
NOR2_X1 U916 ( .A1(KEYINPUT42), .A2(n1200), .ZN(n1199) );
XNOR2_X1 U917 ( .A(G104), .B(G107), .ZN(n1200) );
INV_X1 U918 ( .A(n1179), .ZN(n1004) );
NAND2_X1 U919 ( .A1(G221), .A2(n1201), .ZN(n1179) );
NAND2_X1 U920 ( .A1(G234), .A2(n1188), .ZN(n1201) );
INV_X1 U921 ( .A(n1137), .ZN(n971) );
NOR2_X1 U922 ( .A1(n985), .A2(n1009), .ZN(n1137) );
INV_X1 U923 ( .A(n987), .ZN(n1009) );
NAND2_X1 U924 ( .A1(G214), .A2(n1202), .ZN(n987) );
XNOR2_X1 U925 ( .A(n1024), .B(n1203), .ZN(n985) );
NOR2_X1 U926 ( .A1(n1023), .A2(KEYINPUT2), .ZN(n1203) );
AND2_X1 U927 ( .A1(n1204), .A2(n1188), .ZN(n1023) );
XOR2_X1 U928 ( .A(n1205), .B(n1206), .Z(n1204) );
XNOR2_X1 U929 ( .A(n1151), .B(n1207), .ZN(n1206) );
XOR2_X1 U930 ( .A(KEYINPUT61), .B(G125), .Z(n1207) );
NAND2_X1 U931 ( .A1(G224), .A2(n982), .ZN(n1151) );
XOR2_X1 U932 ( .A(n1153), .B(n1108), .Z(n1205) );
XNOR2_X1 U933 ( .A(n1061), .B(n1208), .ZN(n1108) );
NOR2_X1 U934 ( .A1(n1062), .A2(KEYINPUT10), .ZN(n1208) );
AND2_X1 U935 ( .A1(n1209), .A2(n1210), .ZN(n1062) );
NAND2_X1 U936 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XOR2_X1 U937 ( .A(KEYINPUT17), .B(n1213), .Z(n1209) );
NOR2_X1 U938 ( .A1(n1211), .A2(n1212), .ZN(n1213) );
XOR2_X1 U939 ( .A(n1214), .B(n1215), .Z(n1061) );
XNOR2_X1 U940 ( .A(n1089), .B(n1216), .ZN(n1215) );
NOR2_X1 U941 ( .A1(KEYINPUT50), .A2(n1217), .ZN(n1216) );
XNOR2_X1 U942 ( .A(G107), .B(n1218), .ZN(n1214) );
XNOR2_X1 U943 ( .A(G122), .B(n1105), .ZN(n1218) );
NAND2_X1 U944 ( .A1(n1219), .A2(n1202), .ZN(n1024) );
NAND2_X1 U945 ( .A1(n1220), .A2(n1188), .ZN(n1202) );
XNOR2_X1 U946 ( .A(G210), .B(KEYINPUT20), .ZN(n1219) );
INV_X1 U947 ( .A(n997), .ZN(n1140) );
NOR2_X1 U948 ( .A1(n1160), .A2(n1177), .ZN(n997) );
XOR2_X1 U949 ( .A(n1022), .B(n1221), .Z(n1177) );
NOR2_X1 U950 ( .A1(G475), .A2(KEYINPUT25), .ZN(n1221) );
NAND2_X1 U951 ( .A1(n1077), .A2(n1188), .ZN(n1022) );
XOR2_X1 U952 ( .A(n1222), .B(n1223), .Z(n1077) );
XOR2_X1 U953 ( .A(n1224), .B(n1225), .Z(n1223) );
XOR2_X1 U954 ( .A(G143), .B(G131), .Z(n1225) );
XOR2_X1 U955 ( .A(KEYINPUT53), .B(G146), .Z(n1224) );
XOR2_X1 U956 ( .A(n1226), .B(n1227), .Z(n1222) );
XNOR2_X1 U957 ( .A(n1228), .B(n1041), .ZN(n1227) );
AND3_X1 U958 ( .A1(G214), .A2(n982), .A3(n1220), .ZN(n1228) );
XNOR2_X1 U959 ( .A(n1229), .B(n1217), .ZN(n1226) );
INV_X1 U960 ( .A(G104), .ZN(n1217) );
NAND2_X1 U961 ( .A1(n1230), .A2(KEYINPUT18), .ZN(n1229) );
XNOR2_X1 U962 ( .A(G113), .B(n1231), .ZN(n1230) );
NOR2_X1 U963 ( .A1(G122), .A2(KEYINPUT14), .ZN(n1231) );
XOR2_X1 U964 ( .A(n1028), .B(n1075), .Z(n1160) );
INV_X1 U965 ( .A(G478), .ZN(n1075) );
NAND2_X1 U966 ( .A1(n1072), .A2(n1188), .ZN(n1028) );
XNOR2_X1 U967 ( .A(n1232), .B(n1233), .ZN(n1072) );
XNOR2_X1 U968 ( .A(n1168), .B(n1234), .ZN(n1233) );
XOR2_X1 U969 ( .A(KEYINPUT7), .B(G143), .Z(n1234) );
INV_X1 U970 ( .A(G134), .ZN(n1168) );
XOR2_X1 U971 ( .A(n1235), .B(n1236), .Z(n1232) );
AND3_X1 U972 ( .A1(G217), .A2(n982), .A3(G234), .ZN(n1236) );
XNOR2_X1 U973 ( .A(G128), .B(n1237), .ZN(n1235) );
NOR2_X1 U974 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
XOR2_X1 U975 ( .A(n1240), .B(KEYINPUT19), .Z(n1239) );
NAND2_X1 U976 ( .A1(n1241), .A2(G107), .ZN(n1240) );
XNOR2_X1 U977 ( .A(n1242), .B(KEYINPUT13), .ZN(n1241) );
NOR2_X1 U978 ( .A1(G107), .A2(n1242), .ZN(n1238) );
XOR2_X1 U979 ( .A(G116), .B(n1243), .Z(n1242) );
XOR2_X1 U980 ( .A(KEYINPUT37), .B(G122), .Z(n1243) );
NAND2_X1 U981 ( .A1(n1171), .A2(n1018), .ZN(n1008) );
NAND3_X1 U982 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1018) );
NAND2_X1 U983 ( .A1(G217), .A2(G902), .ZN(n1246) );
OR3_X1 U984 ( .A1(n1067), .A2(G902), .A3(n1247), .ZN(n1245) );
NAND2_X1 U985 ( .A1(n1247), .A2(n1067), .ZN(n1244) );
XOR2_X1 U986 ( .A(n1248), .B(n1249), .Z(n1067) );
XNOR2_X1 U987 ( .A(n1250), .B(n1251), .ZN(n1249) );
XOR2_X1 U988 ( .A(n1252), .B(n1253), .Z(n1251) );
NAND2_X1 U989 ( .A1(KEYINPUT4), .A2(n1254), .ZN(n1252) );
INV_X1 U990 ( .A(G119), .ZN(n1254) );
INV_X1 U991 ( .A(n1041), .ZN(n1250) );
XNOR2_X1 U992 ( .A(G140), .B(G125), .ZN(n1041) );
XOR2_X1 U993 ( .A(n1255), .B(n1256), .Z(n1248) );
XOR2_X1 U994 ( .A(KEYINPUT12), .B(G137), .Z(n1256) );
XNOR2_X1 U995 ( .A(n1257), .B(n1105), .ZN(n1255) );
INV_X1 U996 ( .A(G110), .ZN(n1105) );
NAND4_X1 U997 ( .A1(KEYINPUT30), .A2(G221), .A3(G234), .A4(n982), .ZN(n1257) );
NOR2_X1 U998 ( .A1(n1070), .A2(G234), .ZN(n1247) );
INV_X1 U999 ( .A(G217), .ZN(n1070) );
INV_X1 U1000 ( .A(n1156), .ZN(n1171) );
XOR2_X1 U1001 ( .A(n1258), .B(n1025), .Z(n1156) );
INV_X1 U1002 ( .A(G472), .ZN(n1025) );
NAND2_X1 U1003 ( .A1(KEYINPUT41), .A2(n1026), .ZN(n1258) );
AND2_X1 U1004 ( .A1(n1259), .A2(n1188), .ZN(n1026) );
INV_X1 U1005 ( .A(G902), .ZN(n1188) );
XOR2_X1 U1006 ( .A(n1260), .B(n1261), .Z(n1259) );
NOR2_X1 U1007 ( .A1(n1090), .A2(n1262), .ZN(n1261) );
XOR2_X1 U1008 ( .A(KEYINPUT3), .B(n1263), .Z(n1262) );
NOR2_X1 U1009 ( .A1(n1087), .A2(G101), .ZN(n1263) );
INV_X1 U1010 ( .A(n1264), .ZN(n1087) );
NOR2_X1 U1011 ( .A1(n1264), .A2(n1089), .ZN(n1090) );
INV_X1 U1012 ( .A(G101), .ZN(n1089) );
NAND3_X1 U1013 ( .A1(n1265), .A2(n1220), .A3(G210), .ZN(n1264) );
INV_X1 U1014 ( .A(G237), .ZN(n1220) );
XNOR2_X1 U1015 ( .A(KEYINPUT58), .B(n982), .ZN(n1265) );
INV_X1 U1016 ( .A(G953), .ZN(n982) );
NOR2_X1 U1017 ( .A1(KEYINPUT0), .A2(n1091), .ZN(n1260) );
XNOR2_X1 U1018 ( .A(n1266), .B(n1267), .ZN(n1091) );
XOR2_X1 U1019 ( .A(n1268), .B(n1269), .Z(n1267) );
XNOR2_X1 U1020 ( .A(KEYINPUT35), .B(n1212), .ZN(n1269) );
INV_X1 U1021 ( .A(G113), .ZN(n1212) );
NOR2_X1 U1022 ( .A1(KEYINPUT60), .A2(n1270), .ZN(n1268) );
XOR2_X1 U1023 ( .A(n1211), .B(KEYINPUT6), .Z(n1270) );
XNOR2_X1 U1024 ( .A(G116), .B(G119), .ZN(n1211) );
XNOR2_X1 U1025 ( .A(n1153), .B(n1099), .ZN(n1266) );
XOR2_X1 U1026 ( .A(n1271), .B(n1046), .Z(n1099) );
XOR2_X1 U1027 ( .A(G134), .B(G137), .Z(n1046) );
XNOR2_X1 U1028 ( .A(G131), .B(KEYINPUT8), .ZN(n1271) );
XNOR2_X1 U1029 ( .A(n1040), .B(KEYINPUT28), .ZN(n1153) );
XOR2_X1 U1030 ( .A(G143), .B(n1253), .Z(n1040) );
XNOR2_X1 U1031 ( .A(n1272), .B(G146), .ZN(n1253) );
INV_X1 U1032 ( .A(G128), .ZN(n1272) );
endmodule


