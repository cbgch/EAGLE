//Key = 1110001010010000011011000000101001001100101101001101001101000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325;

XOR2_X1 U731 ( .A(n1007), .B(n1008), .Z(G9) );
NAND3_X1 U732 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(G75) );
NAND2_X1 U733 ( .A1(G952), .A2(n1012), .ZN(n1011) );
NAND4_X1 U734 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
NOR3_X1 U735 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1016) );
NAND3_X1 U736 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1015) );
NAND2_X1 U737 ( .A1(n1023), .A2(n1024), .ZN(n1020) );
NAND4_X1 U738 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
NAND2_X1 U739 ( .A1(n1029), .A2(n1030), .ZN(n1023) );
NAND2_X1 U740 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U741 ( .A1(n1033), .A2(n1026), .ZN(n1032) );
NAND2_X1 U742 ( .A1(n1028), .A2(n1034), .ZN(n1031) );
NAND2_X1 U743 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U744 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U745 ( .A1(n1026), .A2(n1039), .ZN(n1013) );
NAND2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U747 ( .A1(n1042), .A2(n1021), .ZN(n1041) );
NAND2_X1 U748 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND3_X1 U749 ( .A1(n1028), .A2(n1045), .A3(n1022), .ZN(n1044) );
NAND2_X1 U750 ( .A1(n1029), .A2(n1046), .ZN(n1043) );
NAND2_X1 U751 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U752 ( .A1(n1049), .A2(n1050), .A3(n1022), .ZN(n1048) );
INV_X1 U753 ( .A(KEYINPUT58), .ZN(n1050) );
NAND2_X1 U754 ( .A1(n1028), .A2(n1051), .ZN(n1047) );
OR2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U756 ( .A1(KEYINPUT58), .A2(n1054), .ZN(n1040) );
NAND4_X1 U757 ( .A1(n1022), .A2(n1049), .A3(n1029), .A4(n1021), .ZN(n1054) );
NAND4_X1 U758 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1009) );
NOR4_X1 U759 ( .A1(n1025), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1058) );
XNOR2_X1 U760 ( .A(n1062), .B(n1063), .ZN(n1060) );
NOR2_X1 U761 ( .A1(G478), .A2(KEYINPUT44), .ZN(n1063) );
NOR2_X1 U762 ( .A1(KEYINPUT48), .A2(n1064), .ZN(n1059) );
NOR2_X1 U763 ( .A1(n1065), .A2(n1066), .ZN(n1057) );
XOR2_X1 U764 ( .A(n1067), .B(n1068), .Z(n1066) );
NAND2_X1 U765 ( .A1(KEYINPUT48), .A2(n1064), .ZN(n1068) );
XOR2_X1 U766 ( .A(n1069), .B(KEYINPUT40), .Z(n1064) );
XOR2_X1 U767 ( .A(n1027), .B(KEYINPUT24), .Z(n1056) );
XNOR2_X1 U768 ( .A(n1070), .B(KEYINPUT31), .ZN(n1055) );
XOR2_X1 U769 ( .A(n1071), .B(n1072), .Z(G72) );
NOR2_X1 U770 ( .A1(n1073), .A2(n1010), .ZN(n1072) );
NOR2_X1 U771 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U772 ( .A1(n1076), .A2(n1077), .ZN(n1071) );
NAND2_X1 U773 ( .A1(n1078), .A2(n1010), .ZN(n1077) );
XNOR2_X1 U774 ( .A(n1019), .B(n1079), .ZN(n1078) );
OR3_X1 U775 ( .A1(n1075), .A2(n1079), .A3(n1010), .ZN(n1076) );
XNOR2_X1 U776 ( .A(n1080), .B(n1081), .ZN(n1079) );
XNOR2_X1 U777 ( .A(n1082), .B(n1083), .ZN(n1081) );
NAND2_X1 U778 ( .A1(KEYINPUT1), .A2(n1084), .ZN(n1082) );
XOR2_X1 U779 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U780 ( .A1(KEYINPUT11), .A2(n1087), .ZN(n1086) );
INV_X1 U781 ( .A(G140), .ZN(n1087) );
NAND2_X1 U782 ( .A1(n1088), .A2(n1089), .ZN(n1080) );
NAND2_X1 U783 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U784 ( .A(n1092), .B(KEYINPUT43), .Z(n1090) );
NAND2_X1 U785 ( .A1(n1093), .A2(G131), .ZN(n1088) );
XOR2_X1 U786 ( .A(n1092), .B(KEYINPUT53), .Z(n1093) );
XOR2_X1 U787 ( .A(n1094), .B(KEYINPUT7), .Z(n1092) );
XOR2_X1 U788 ( .A(n1095), .B(n1096), .Z(G69) );
NOR2_X1 U789 ( .A1(n1097), .A2(n1010), .ZN(n1096) );
AND2_X1 U790 ( .A1(G224), .A2(G898), .ZN(n1097) );
NAND2_X1 U791 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
NAND3_X1 U792 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
NAND2_X1 U793 ( .A1(G953), .A2(n1103), .ZN(n1101) );
OR2_X1 U794 ( .A1(n1102), .A2(n1100), .ZN(n1098) );
NAND2_X1 U795 ( .A1(n1010), .A2(n1104), .ZN(n1102) );
NAND3_X1 U796 ( .A1(n1105), .A2(n1014), .A3(n1106), .ZN(n1104) );
INV_X1 U797 ( .A(n1018), .ZN(n1106) );
XNOR2_X1 U798 ( .A(KEYINPUT47), .B(n1017), .ZN(n1105) );
NOR2_X1 U799 ( .A1(n1107), .A2(n1108), .ZN(G66) );
XNOR2_X1 U800 ( .A(n1109), .B(n1110), .ZN(n1108) );
XOR2_X1 U801 ( .A(KEYINPUT41), .B(n1111), .Z(n1110) );
NOR2_X1 U802 ( .A1(n1069), .A2(n1112), .ZN(n1111) );
NOR2_X1 U803 ( .A1(n1107), .A2(n1113), .ZN(G63) );
NOR3_X1 U804 ( .A1(n1062), .A2(n1114), .A3(n1115), .ZN(n1113) );
AND4_X1 U805 ( .A1(n1116), .A2(KEYINPUT8), .A3(G478), .A4(n1117), .ZN(n1115) );
NOR2_X1 U806 ( .A1(n1118), .A2(n1116), .ZN(n1114) );
AND3_X1 U807 ( .A1(KEYINPUT8), .A2(n1119), .A3(G478), .ZN(n1118) );
NOR2_X1 U808 ( .A1(n1107), .A2(n1120), .ZN(G60) );
NOR2_X1 U809 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U810 ( .A(KEYINPUT46), .B(n1123), .Z(n1122) );
NOR2_X1 U811 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
AND2_X1 U812 ( .A1(n1125), .A2(n1124), .ZN(n1121) );
NAND2_X1 U813 ( .A1(n1117), .A2(G475), .ZN(n1125) );
XNOR2_X1 U814 ( .A(G104), .B(n1126), .ZN(G6) );
NOR2_X1 U815 ( .A1(n1127), .A2(KEYINPUT13), .ZN(n1126) );
INV_X1 U816 ( .A(n1128), .ZN(n1127) );
NOR3_X1 U817 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(G57) );
NOR3_X1 U818 ( .A1(n1132), .A2(G953), .A3(G952), .ZN(n1131) );
AND2_X1 U819 ( .A1(n1132), .A2(n1107), .ZN(n1130) );
INV_X1 U820 ( .A(KEYINPUT38), .ZN(n1132) );
NOR2_X1 U821 ( .A1(n1133), .A2(n1134), .ZN(n1129) );
XOR2_X1 U822 ( .A(n1135), .B(KEYINPUT55), .Z(n1134) );
NAND2_X1 U823 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NOR2_X1 U824 ( .A1(n1136), .A2(n1137), .ZN(n1133) );
XOR2_X1 U825 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U826 ( .A(n1140), .B(n1141), .Z(n1136) );
XOR2_X1 U827 ( .A(n1142), .B(n1143), .Z(n1141) );
AND2_X1 U828 ( .A1(G472), .A2(n1117), .ZN(n1143) );
NOR2_X1 U829 ( .A1(KEYINPUT3), .A2(n1144), .ZN(n1142) );
NAND2_X1 U830 ( .A1(n1145), .A2(n1146), .ZN(n1140) );
XNOR2_X1 U831 ( .A(n1147), .B(KEYINPUT4), .ZN(n1145) );
NOR2_X1 U832 ( .A1(n1107), .A2(n1148), .ZN(G54) );
XOR2_X1 U833 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U834 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U835 ( .A(n1153), .B(n1154), .Z(n1149) );
XNOR2_X1 U836 ( .A(n1155), .B(n1156), .ZN(n1154) );
AND2_X1 U837 ( .A1(G469), .A2(n1117), .ZN(n1153) );
INV_X1 U838 ( .A(n1112), .ZN(n1117) );
NOR2_X1 U839 ( .A1(n1107), .A2(n1157), .ZN(G51) );
XOR2_X1 U840 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U841 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U842 ( .A(n1162), .B(n1163), .Z(n1160) );
XOR2_X1 U843 ( .A(n1164), .B(n1165), .Z(n1158) );
XOR2_X1 U844 ( .A(KEYINPUT29), .B(n1166), .Z(n1165) );
NOR2_X1 U845 ( .A1(n1167), .A2(n1112), .ZN(n1166) );
NAND2_X1 U846 ( .A1(G902), .A2(n1119), .ZN(n1112) );
OR4_X1 U847 ( .A1(n1017), .A2(n1018), .A3(n1168), .A4(n1169), .ZN(n1119) );
INV_X1 U848 ( .A(n1014), .ZN(n1169) );
XOR2_X1 U849 ( .A(KEYINPUT56), .B(n1019), .Z(n1168) );
NAND4_X1 U850 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1019) );
NOR4_X1 U851 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1173) );
INV_X1 U852 ( .A(n1178), .ZN(n1174) );
AND2_X1 U853 ( .A1(n1179), .A2(n1180), .ZN(n1172) );
NAND3_X1 U854 ( .A1(n1181), .A2(n1008), .A3(n1128), .ZN(n1018) );
NAND3_X1 U855 ( .A1(n1182), .A2(n1028), .A3(n1052), .ZN(n1128) );
NAND3_X1 U856 ( .A1(n1053), .A2(n1028), .A3(n1182), .ZN(n1008) );
NAND4_X1 U857 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1017) );
NAND3_X1 U858 ( .A1(n1029), .A2(n1187), .A3(n1188), .ZN(n1183) );
INV_X1 U859 ( .A(n1189), .ZN(n1188) );
XOR2_X1 U860 ( .A(KEYINPUT52), .B(n1190), .Z(n1187) );
NOR2_X1 U861 ( .A1(n1010), .A2(G952), .ZN(n1107) );
XOR2_X1 U862 ( .A(n1191), .B(n1192), .Z(G48) );
XOR2_X1 U863 ( .A(KEYINPUT25), .B(G146), .Z(n1192) );
NAND2_X1 U864 ( .A1(n1193), .A2(n1194), .ZN(n1191) );
NAND3_X1 U865 ( .A1(n1190), .A2(n1195), .A3(n1196), .ZN(n1194) );
NAND2_X1 U866 ( .A1(n1197), .A2(n1052), .ZN(n1195) );
OR2_X1 U867 ( .A1(n1170), .A2(n1196), .ZN(n1193) );
INV_X1 U868 ( .A(KEYINPUT30), .ZN(n1196) );
NAND3_X1 U869 ( .A1(n1052), .A2(n1190), .A3(n1197), .ZN(n1170) );
NAND2_X1 U870 ( .A1(n1198), .A2(n1199), .ZN(G45) );
NAND2_X1 U871 ( .A1(G143), .A2(n1200), .ZN(n1199) );
NAND2_X1 U872 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NAND2_X1 U873 ( .A1(KEYINPUT59), .A2(n1203), .ZN(n1202) );
NAND3_X1 U874 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1198) );
INV_X1 U875 ( .A(KEYINPUT59), .ZN(n1206) );
NAND2_X1 U876 ( .A1(n1171), .A2(n1203), .ZN(n1205) );
NAND2_X1 U877 ( .A1(n1201), .A2(n1207), .ZN(n1204) );
NAND2_X1 U878 ( .A1(n1208), .A2(n1203), .ZN(n1207) );
INV_X1 U879 ( .A(KEYINPUT10), .ZN(n1203) );
INV_X1 U880 ( .A(n1171), .ZN(n1201) );
NAND4_X1 U881 ( .A1(n1209), .A2(n1190), .A3(n1210), .A4(n1070), .ZN(n1171) );
XOR2_X1 U882 ( .A(n1211), .B(G140), .Z(G42) );
NAND2_X1 U883 ( .A1(KEYINPUT18), .A2(n1180), .ZN(n1211) );
NAND3_X1 U884 ( .A1(n1033), .A2(n1052), .A3(n1212), .ZN(n1180) );
AND3_X1 U885 ( .A1(n1026), .A2(n1213), .A3(n1045), .ZN(n1212) );
NAND2_X1 U886 ( .A1(n1214), .A2(n1215), .ZN(G39) );
NAND2_X1 U887 ( .A1(n1176), .A2(n1216), .ZN(n1215) );
XOR2_X1 U888 ( .A(KEYINPUT37), .B(n1217), .Z(n1214) );
NOR2_X1 U889 ( .A1(n1176), .A2(n1216), .ZN(n1217) );
AND3_X1 U890 ( .A1(n1022), .A2(n1026), .A3(n1197), .ZN(n1176) );
XOR2_X1 U891 ( .A(G134), .B(n1218), .Z(G36) );
NOR2_X1 U892 ( .A1(KEYINPUT39), .A2(n1179), .ZN(n1218) );
NAND3_X1 U893 ( .A1(n1026), .A2(n1053), .A3(n1209), .ZN(n1179) );
XOR2_X1 U894 ( .A(G131), .B(n1175), .Z(G33) );
AND3_X1 U895 ( .A1(n1052), .A2(n1026), .A3(n1209), .ZN(n1175) );
AND3_X1 U896 ( .A1(n1045), .A2(n1213), .A3(n1049), .ZN(n1209) );
INV_X1 U897 ( .A(n1065), .ZN(n1026) );
NAND2_X1 U898 ( .A1(n1038), .A2(n1219), .ZN(n1065) );
NAND2_X1 U899 ( .A1(n1220), .A2(n1221), .ZN(G30) );
NAND2_X1 U900 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
XOR2_X1 U901 ( .A(KEYINPUT19), .B(n1177), .Z(n1222) );
INV_X1 U902 ( .A(n1224), .ZN(n1177) );
NAND2_X1 U903 ( .A1(G128), .A2(n1225), .ZN(n1220) );
XOR2_X1 U904 ( .A(n1224), .B(KEYINPUT50), .Z(n1225) );
NAND3_X1 U905 ( .A1(n1053), .A2(n1190), .A3(n1197), .ZN(n1224) );
AND4_X1 U906 ( .A1(n1045), .A2(n1226), .A3(n1061), .A4(n1213), .ZN(n1197) );
XOR2_X1 U907 ( .A(n1227), .B(n1228), .Z(G3) );
XOR2_X1 U908 ( .A(KEYINPUT22), .B(G101), .Z(n1228) );
NAND2_X1 U909 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
OR2_X1 U910 ( .A1(n1014), .A2(KEYINPUT15), .ZN(n1230) );
NAND3_X1 U911 ( .A1(n1049), .A2(n1182), .A3(n1022), .ZN(n1014) );
NAND4_X1 U912 ( .A1(n1182), .A2(n1231), .A3(n1049), .A4(KEYINPUT15), .ZN(n1229) );
INV_X1 U913 ( .A(n1022), .ZN(n1231) );
XOR2_X1 U914 ( .A(n1085), .B(n1178), .Z(G27) );
NAND4_X1 U915 ( .A1(n1033), .A2(n1052), .A3(n1232), .A4(n1029), .ZN(n1178) );
AND2_X1 U916 ( .A1(n1213), .A2(n1190), .ZN(n1232) );
NAND2_X1 U917 ( .A1(n1233), .A2(n1234), .ZN(n1213) );
NAND2_X1 U918 ( .A1(n1235), .A2(n1075), .ZN(n1233) );
INV_X1 U919 ( .A(G900), .ZN(n1075) );
XOR2_X1 U920 ( .A(n1236), .B(n1237), .Z(G24) );
XOR2_X1 U921 ( .A(KEYINPUT61), .B(G122), .Z(n1237) );
NOR3_X1 U922 ( .A1(n1189), .A2(n1238), .A3(n1035), .ZN(n1236) );
INV_X1 U923 ( .A(n1190), .ZN(n1035) );
XNOR2_X1 U924 ( .A(n1029), .B(KEYINPUT62), .ZN(n1238) );
NAND4_X1 U925 ( .A1(n1028), .A2(n1210), .A3(n1070), .A4(n1239), .ZN(n1189) );
AND2_X1 U926 ( .A1(n1240), .A2(n1241), .ZN(n1028) );
XNOR2_X1 U927 ( .A(G119), .B(n1184), .ZN(G21) );
NAND4_X1 U928 ( .A1(n1022), .A2(n1242), .A3(n1226), .A4(n1061), .ZN(n1184) );
XNOR2_X1 U929 ( .A(G116), .B(n1185), .ZN(G18) );
NAND3_X1 U930 ( .A1(n1242), .A2(n1053), .A3(n1049), .ZN(n1185) );
NOR2_X1 U931 ( .A1(n1070), .A2(n1243), .ZN(n1053) );
XOR2_X1 U932 ( .A(n1244), .B(n1245), .Z(G15) );
NAND2_X1 U933 ( .A1(KEYINPUT6), .A2(n1246), .ZN(n1245) );
INV_X1 U934 ( .A(n1186), .ZN(n1246) );
NAND3_X1 U935 ( .A1(n1049), .A2(n1242), .A3(n1052), .ZN(n1186) );
AND2_X1 U936 ( .A1(n1243), .A2(n1070), .ZN(n1052) );
INV_X1 U937 ( .A(n1210), .ZN(n1243) );
AND3_X1 U938 ( .A1(n1190), .A2(n1239), .A3(n1029), .ZN(n1242) );
NOR2_X1 U939 ( .A1(n1247), .A2(n1025), .ZN(n1029) );
INV_X1 U940 ( .A(n1027), .ZN(n1247) );
AND2_X1 U941 ( .A1(n1240), .A2(n1061), .ZN(n1049) );
INV_X1 U942 ( .A(n1241), .ZN(n1061) );
XNOR2_X1 U943 ( .A(G110), .B(n1181), .ZN(G12) );
NAND3_X1 U944 ( .A1(n1022), .A2(n1182), .A3(n1033), .ZN(n1181) );
AND2_X1 U945 ( .A1(n1241), .A2(n1226), .ZN(n1033) );
XNOR2_X1 U946 ( .A(n1240), .B(KEYINPUT16), .ZN(n1226) );
XNOR2_X1 U947 ( .A(n1067), .B(n1069), .ZN(n1240) );
NAND2_X1 U948 ( .A1(G217), .A2(n1248), .ZN(n1069) );
NAND2_X1 U949 ( .A1(n1249), .A2(n1109), .ZN(n1067) );
XNOR2_X1 U950 ( .A(n1250), .B(n1251), .ZN(n1109) );
XOR2_X1 U951 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U952 ( .A(n1216), .B(G140), .Z(n1253) );
NAND2_X1 U953 ( .A1(n1254), .A2(G221), .ZN(n1252) );
XOR2_X1 U954 ( .A(n1162), .B(n1255), .Z(n1250) );
XOR2_X1 U955 ( .A(n1085), .B(n1256), .Z(n1162) );
INV_X1 U956 ( .A(G125), .ZN(n1085) );
XOR2_X1 U957 ( .A(KEYINPUT20), .B(G902), .Z(n1249) );
XOR2_X1 U958 ( .A(n1257), .B(G472), .Z(n1241) );
NAND2_X1 U959 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XOR2_X1 U960 ( .A(n1260), .B(n1261), .Z(n1258) );
XOR2_X1 U961 ( .A(n1262), .B(n1263), .Z(n1261) );
NOR2_X1 U962 ( .A1(KEYINPUT35), .A2(n1144), .ZN(n1263) );
XOR2_X1 U963 ( .A(n1264), .B(G113), .Z(n1144) );
NAND2_X1 U964 ( .A1(n1265), .A2(KEYINPUT21), .ZN(n1264) );
XNOR2_X1 U965 ( .A(G116), .B(n1266), .ZN(n1265) );
XOR2_X1 U966 ( .A(KEYINPUT42), .B(G119), .Z(n1266) );
NAND2_X1 U967 ( .A1(KEYINPUT28), .A2(n1267), .ZN(n1262) );
XNOR2_X1 U968 ( .A(n1138), .B(n1268), .ZN(n1267) );
NOR2_X1 U969 ( .A1(KEYINPUT60), .A2(n1139), .ZN(n1268) );
NAND2_X1 U970 ( .A1(n1269), .A2(G210), .ZN(n1138) );
NAND2_X1 U971 ( .A1(n1270), .A2(n1146), .ZN(n1260) );
NAND2_X1 U972 ( .A1(n1163), .A2(n1156), .ZN(n1146) );
XOR2_X1 U973 ( .A(KEYINPUT49), .B(n1147), .Z(n1270) );
NOR2_X1 U974 ( .A1(n1156), .A2(n1163), .ZN(n1147) );
AND3_X1 U975 ( .A1(n1045), .A2(n1239), .A3(n1190), .ZN(n1182) );
NOR2_X1 U976 ( .A1(n1038), .A2(n1037), .ZN(n1190) );
INV_X1 U977 ( .A(n1219), .ZN(n1037) );
NAND2_X1 U978 ( .A1(G214), .A2(n1271), .ZN(n1219) );
XNOR2_X1 U979 ( .A(n1272), .B(n1167), .ZN(n1038) );
NAND2_X1 U980 ( .A1(G210), .A2(n1271), .ZN(n1167) );
NAND2_X1 U981 ( .A1(n1273), .A2(n1259), .ZN(n1271) );
INV_X1 U982 ( .A(G237), .ZN(n1273) );
NAND3_X1 U983 ( .A1(n1274), .A2(n1259), .A3(n1275), .ZN(n1272) );
XOR2_X1 U984 ( .A(KEYINPUT57), .B(n1276), .Z(n1275) );
NOR2_X1 U985 ( .A1(n1100), .A2(n1277), .ZN(n1276) );
NAND2_X1 U986 ( .A1(n1277), .A2(n1100), .ZN(n1274) );
XNOR2_X1 U987 ( .A(n1161), .B(n1256), .ZN(n1100) );
XOR2_X1 U988 ( .A(G110), .B(G119), .Z(n1256) );
XNOR2_X1 U989 ( .A(n1278), .B(n1279), .ZN(n1161) );
XOR2_X1 U990 ( .A(n1244), .B(n1280), .Z(n1278) );
XOR2_X1 U991 ( .A(n1164), .B(n1281), .Z(n1277) );
NOR2_X1 U992 ( .A1(KEYINPUT32), .A2(n1282), .ZN(n1281) );
XOR2_X1 U993 ( .A(G125), .B(n1163), .Z(n1282) );
XOR2_X1 U994 ( .A(n1083), .B(KEYINPUT12), .Z(n1163) );
NAND2_X1 U995 ( .A1(G224), .A2(n1010), .ZN(n1164) );
NAND2_X1 U996 ( .A1(n1283), .A2(n1234), .ZN(n1239) );
NAND3_X1 U997 ( .A1(n1284), .A2(n1010), .A3(G952), .ZN(n1234) );
XNOR2_X1 U998 ( .A(KEYINPUT36), .B(n1021), .ZN(n1284) );
XOR2_X1 U999 ( .A(n1285), .B(KEYINPUT27), .Z(n1283) );
NAND2_X1 U1000 ( .A1(n1235), .A2(n1103), .ZN(n1285) );
INV_X1 U1001 ( .A(G898), .ZN(n1103) );
AND3_X1 U1002 ( .A1(G953), .A2(n1021), .A3(n1286), .ZN(n1235) );
XOR2_X1 U1003 ( .A(n1259), .B(KEYINPUT51), .Z(n1286) );
NAND2_X1 U1004 ( .A1(G237), .A2(G234), .ZN(n1021) );
NOR2_X1 U1005 ( .A1(n1027), .A2(n1025), .ZN(n1045) );
AND2_X1 U1006 ( .A1(G221), .A2(n1248), .ZN(n1025) );
NAND2_X1 U1007 ( .A1(G234), .A2(n1259), .ZN(n1248) );
XOR2_X1 U1008 ( .A(n1287), .B(G469), .Z(n1027) );
NAND2_X1 U1009 ( .A1(n1288), .A2(n1259), .ZN(n1287) );
XOR2_X1 U1010 ( .A(n1289), .B(n1290), .Z(n1288) );
XNOR2_X1 U1011 ( .A(n1291), .B(n1156), .ZN(n1290) );
NAND2_X1 U1012 ( .A1(n1292), .A2(n1293), .ZN(n1156) );
NAND2_X1 U1013 ( .A1(n1294), .A2(n1091), .ZN(n1293) );
XOR2_X1 U1014 ( .A(KEYINPUT33), .B(n1295), .Z(n1292) );
NOR2_X1 U1015 ( .A1(n1091), .A2(n1294), .ZN(n1295) );
XOR2_X1 U1016 ( .A(KEYINPUT5), .B(n1296), .Z(n1294) );
INV_X1 U1017 ( .A(n1094), .ZN(n1296) );
XOR2_X1 U1018 ( .A(n1216), .B(n1297), .Z(n1094) );
INV_X1 U1019 ( .A(G137), .ZN(n1216) );
INV_X1 U1020 ( .A(G131), .ZN(n1091) );
NOR2_X1 U1021 ( .A1(KEYINPUT14), .A2(n1298), .ZN(n1291) );
XOR2_X1 U1022 ( .A(n1155), .B(n1299), .Z(n1298) );
NOR2_X1 U1023 ( .A1(KEYINPUT63), .A2(n1151), .ZN(n1299) );
XOR2_X1 U1024 ( .A(G110), .B(G140), .Z(n1151) );
NOR2_X1 U1025 ( .A1(n1074), .A2(G953), .ZN(n1155) );
INV_X1 U1026 ( .A(G227), .ZN(n1074) );
NAND2_X1 U1027 ( .A1(KEYINPUT0), .A2(n1152), .ZN(n1289) );
XOR2_X1 U1028 ( .A(n1279), .B(n1083), .Z(n1152) );
XNOR2_X1 U1029 ( .A(n1300), .B(n1255), .ZN(n1083) );
XOR2_X1 U1030 ( .A(G146), .B(G128), .Z(n1255) );
XOR2_X1 U1031 ( .A(n1208), .B(KEYINPUT54), .Z(n1300) );
INV_X1 U1032 ( .A(G143), .ZN(n1208) );
XNOR2_X1 U1033 ( .A(n1301), .B(n1302), .ZN(n1279) );
XOR2_X1 U1034 ( .A(KEYINPUT23), .B(G107), .Z(n1302) );
XOR2_X1 U1035 ( .A(G104), .B(n1139), .Z(n1301) );
INV_X1 U1036 ( .A(G101), .ZN(n1139) );
NOR2_X1 U1037 ( .A1(n1210), .A2(n1070), .ZN(n1022) );
XNOR2_X1 U1038 ( .A(n1303), .B(G475), .ZN(n1070) );
NAND2_X1 U1039 ( .A1(n1124), .A2(n1259), .ZN(n1303) );
INV_X1 U1040 ( .A(G902), .ZN(n1259) );
XNOR2_X1 U1041 ( .A(n1304), .B(n1305), .ZN(n1124) );
XOR2_X1 U1042 ( .A(G104), .B(n1306), .Z(n1305) );
NOR2_X1 U1043 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
XOR2_X1 U1044 ( .A(n1309), .B(KEYINPUT45), .Z(n1308) );
NAND2_X1 U1045 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NOR2_X1 U1046 ( .A1(n1310), .A2(n1311), .ZN(n1307) );
XOR2_X1 U1047 ( .A(G125), .B(n1312), .Z(n1311) );
XOR2_X1 U1048 ( .A(G146), .B(G140), .Z(n1312) );
XOR2_X1 U1049 ( .A(n1313), .B(n1314), .Z(n1310) );
NOR2_X1 U1050 ( .A1(G131), .A2(KEYINPUT9), .ZN(n1314) );
XOR2_X1 U1051 ( .A(n1315), .B(G143), .Z(n1313) );
NAND2_X1 U1052 ( .A1(n1269), .A2(G214), .ZN(n1315) );
NOR2_X1 U1053 ( .A1(G953), .A2(G237), .ZN(n1269) );
XOR2_X1 U1054 ( .A(n1244), .B(n1316), .Z(n1304) );
XOR2_X1 U1055 ( .A(KEYINPUT34), .B(G122), .Z(n1316) );
INV_X1 U1056 ( .A(G113), .ZN(n1244) );
XOR2_X1 U1057 ( .A(n1062), .B(G478), .Z(n1210) );
NOR2_X1 U1058 ( .A1(n1116), .A2(G902), .ZN(n1062) );
XNOR2_X1 U1059 ( .A(n1317), .B(n1318), .ZN(n1116) );
XOR2_X1 U1060 ( .A(n1319), .B(n1320), .Z(n1318) );
XOR2_X1 U1061 ( .A(n1223), .B(G143), .Z(n1320) );
INV_X1 U1062 ( .A(G128), .ZN(n1223) );
NAND2_X1 U1063 ( .A1(G217), .A2(n1254), .ZN(n1319) );
AND2_X1 U1064 ( .A1(G234), .A2(n1010), .ZN(n1254) );
INV_X1 U1065 ( .A(G953), .ZN(n1010) );
XOR2_X1 U1066 ( .A(n1321), .B(n1297), .Z(n1317) );
XOR2_X1 U1067 ( .A(G134), .B(KEYINPUT2), .Z(n1297) );
NAND2_X1 U1068 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
OR2_X1 U1069 ( .A1(n1324), .A2(n1007), .ZN(n1323) );
XOR2_X1 U1070 ( .A(n1325), .B(KEYINPUT26), .Z(n1322) );
NAND2_X1 U1071 ( .A1(n1324), .A2(n1007), .ZN(n1325) );
INV_X1 U1072 ( .A(G107), .ZN(n1007) );
XOR2_X1 U1073 ( .A(n1280), .B(KEYINPUT17), .Z(n1324) );
XOR2_X1 U1074 ( .A(G116), .B(G122), .Z(n1280) );
endmodule


