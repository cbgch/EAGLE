//Key = 0000110111110101001100111001001011010011100111000000000000001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290;

XNOR2_X1 U714 ( .A(G107), .B(n975), .ZN(G9) );
NOR2_X1 U715 ( .A1(n976), .A2(n977), .ZN(G75) );
NOR4_X1 U716 ( .A1(n978), .A2(n979), .A3(KEYINPUT3), .A4(G953), .ZN(n977) );
NAND3_X1 U717 ( .A1(n980), .A2(n981), .A3(n982), .ZN(n978) );
NAND2_X1 U718 ( .A1(n983), .A2(n984), .ZN(n981) );
NAND2_X1 U719 ( .A1(n985), .A2(n986), .ZN(n984) );
NAND3_X1 U720 ( .A1(n987), .A2(n988), .A3(n989), .ZN(n986) );
NAND2_X1 U721 ( .A1(n990), .A2(n991), .ZN(n988) );
NAND2_X1 U722 ( .A1(n992), .A2(n993), .ZN(n991) );
NAND2_X1 U723 ( .A1(n994), .A2(n995), .ZN(n993) );
NAND2_X1 U724 ( .A1(n996), .A2(n997), .ZN(n990) );
NAND2_X1 U725 ( .A1(n998), .A2(n999), .ZN(n997) );
NAND2_X1 U726 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NAND3_X1 U727 ( .A1(n996), .A2(n1002), .A3(n992), .ZN(n985) );
NAND2_X1 U728 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND2_X1 U729 ( .A1(n989), .A2(n1005), .ZN(n1004) );
NAND2_X1 U730 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NAND2_X1 U731 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND2_X1 U732 ( .A1(n987), .A2(n1010), .ZN(n1003) );
NAND2_X1 U733 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND2_X1 U734 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
INV_X1 U735 ( .A(n1015), .ZN(n983) );
NOR3_X1 U736 ( .A1(n979), .A2(G953), .A3(G952), .ZN(n976) );
AND4_X1 U737 ( .A1(n1016), .A2(n1017), .A3(n1018), .A4(n1019), .ZN(n979) );
NOR4_X1 U738 ( .A1(n1020), .A2(n1009), .A3(n1021), .A4(n1022), .ZN(n1019) );
INV_X1 U739 ( .A(n996), .ZN(n1021) );
XOR2_X1 U740 ( .A(n1023), .B(KEYINPUT23), .Z(n1020) );
NAND2_X1 U741 ( .A1(G472), .A2(n1024), .ZN(n1023) );
NOR2_X1 U742 ( .A1(n1000), .A2(n1013), .ZN(n1018) );
INV_X1 U743 ( .A(n1025), .ZN(n1013) );
NAND2_X1 U744 ( .A1(n1026), .A2(n1027), .ZN(n1017) );
XNOR2_X1 U745 ( .A(KEYINPUT17), .B(n1024), .ZN(n1026) );
XNOR2_X1 U746 ( .A(n1028), .B(n1029), .ZN(n1016) );
NOR2_X1 U747 ( .A1(G469), .A2(KEYINPUT51), .ZN(n1029) );
NAND2_X1 U748 ( .A1(n1030), .A2(n1031), .ZN(G72) );
NAND2_X1 U749 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U750 ( .A1(G953), .A2(n1034), .ZN(n1032) );
NAND2_X1 U751 ( .A1(G900), .A2(G227), .ZN(n1034) );
NAND2_X1 U752 ( .A1(n1035), .A2(n1036), .ZN(n1030) );
NAND2_X1 U753 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U754 ( .A1(G953), .A2(n1039), .ZN(n1038) );
INV_X1 U755 ( .A(n1033), .ZN(n1035) );
NAND2_X1 U756 ( .A1(n1040), .A2(n1041), .ZN(n1033) );
NAND2_X1 U757 ( .A1(n1042), .A2(n982), .ZN(n1041) );
XOR2_X1 U758 ( .A(KEYINPUT33), .B(n1043), .Z(n1040) );
NOR3_X1 U759 ( .A1(n1044), .A2(G953), .A3(n982), .ZN(n1043) );
XOR2_X1 U760 ( .A(KEYINPUT20), .B(n1042), .Z(n1044) );
AND2_X1 U761 ( .A1(n1045), .A2(n1037), .ZN(n1042) );
INV_X1 U762 ( .A(n1046), .ZN(n1037) );
XOR2_X1 U763 ( .A(n1047), .B(n1048), .Z(n1045) );
NAND2_X1 U764 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NAND2_X1 U765 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U766 ( .A(KEYINPUT49), .B(n1053), .Z(n1051) );
NAND2_X1 U767 ( .A1(n1054), .A2(n1055), .ZN(n1049) );
XNOR2_X1 U768 ( .A(n1053), .B(KEYINPUT54), .ZN(n1055) );
XOR2_X1 U769 ( .A(n1056), .B(n1057), .Z(G69) );
NOR2_X1 U770 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U771 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U772 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U773 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U774 ( .A1(G953), .A2(n1066), .ZN(n1062) );
AND3_X1 U775 ( .A1(n1061), .A2(n1064), .A3(n1066), .ZN(n1058) );
XNOR2_X1 U776 ( .A(n1067), .B(n1068), .ZN(n1061) );
XOR2_X1 U777 ( .A(KEYINPUT35), .B(n1069), .Z(n1068) );
NOR2_X1 U778 ( .A1(n1070), .A2(n1071), .ZN(n1056) );
NOR2_X1 U779 ( .A1(n1072), .A2(KEYINPUT11), .ZN(n1071) );
NOR2_X1 U780 ( .A1(n1073), .A2(n1064), .ZN(n1072) );
NOR3_X1 U781 ( .A1(n1064), .A2(KEYINPUT25), .A3(n1073), .ZN(n1070) );
AND2_X1 U782 ( .A1(G898), .A2(G224), .ZN(n1073) );
NOR2_X1 U783 ( .A1(n1074), .A2(n1075), .ZN(G66) );
XNOR2_X1 U784 ( .A(n1076), .B(n1077), .ZN(n1075) );
NAND2_X1 U785 ( .A1(n1078), .A2(G217), .ZN(n1076) );
NOR2_X1 U786 ( .A1(n1074), .A2(n1079), .ZN(G63) );
XOR2_X1 U787 ( .A(n1080), .B(n1081), .Z(n1079) );
NAND2_X1 U788 ( .A1(n1078), .A2(G478), .ZN(n1080) );
NOR2_X1 U789 ( .A1(n1074), .A2(n1082), .ZN(G60) );
XOR2_X1 U790 ( .A(n1083), .B(n1084), .Z(n1082) );
XOR2_X1 U791 ( .A(n1085), .B(KEYINPUT2), .Z(n1084) );
NAND2_X1 U792 ( .A1(n1078), .A2(G475), .ZN(n1085) );
XNOR2_X1 U793 ( .A(G104), .B(n1086), .ZN(G6) );
NOR2_X1 U794 ( .A1(n1074), .A2(n1087), .ZN(G57) );
XNOR2_X1 U795 ( .A(n1088), .B(n1089), .ZN(n1087) );
NOR2_X1 U796 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U797 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U798 ( .A(n1094), .B(KEYINPUT58), .Z(n1093) );
AND2_X1 U799 ( .A1(n1094), .A2(n1092), .ZN(n1090) );
NAND2_X1 U800 ( .A1(n1078), .A2(G472), .ZN(n1094) );
NOR2_X1 U801 ( .A1(n1074), .A2(n1095), .ZN(G54) );
XOR2_X1 U802 ( .A(n1096), .B(n1097), .Z(n1095) );
AND2_X1 U803 ( .A1(G469), .A2(n1078), .ZN(n1097) );
INV_X1 U804 ( .A(n1098), .ZN(n1078) );
NOR2_X1 U805 ( .A1(KEYINPUT29), .A2(n1099), .ZN(n1096) );
XOR2_X1 U806 ( .A(n1100), .B(n1101), .Z(n1099) );
XNOR2_X1 U807 ( .A(n1102), .B(n1103), .ZN(n1101) );
XNOR2_X1 U808 ( .A(n1104), .B(n1105), .ZN(n1103) );
NOR2_X1 U809 ( .A1(KEYINPUT47), .A2(n1106), .ZN(n1105) );
XOR2_X1 U810 ( .A(n1107), .B(n1108), .Z(n1100) );
XOR2_X1 U811 ( .A(KEYINPUT57), .B(KEYINPUT30), .Z(n1108) );
NOR2_X1 U812 ( .A1(n1074), .A2(n1109), .ZN(G51) );
NOR2_X1 U813 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U814 ( .A(n1112), .B(KEYINPUT44), .Z(n1111) );
NAND2_X1 U815 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U816 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
XNOR2_X1 U817 ( .A(n1115), .B(n1116), .ZN(n1114) );
NOR2_X1 U818 ( .A1(n1098), .A2(n1117), .ZN(n1113) );
NAND2_X1 U819 ( .A1(G902), .A2(n1118), .ZN(n1098) );
NAND2_X1 U820 ( .A1(n982), .A2(n980), .ZN(n1118) );
INV_X1 U821 ( .A(n1066), .ZN(n980) );
NAND4_X1 U822 ( .A1(n1119), .A2(n1086), .A3(n1120), .A4(n1121), .ZN(n1066) );
AND4_X1 U823 ( .A1(n975), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1121) );
NAND3_X1 U824 ( .A1(n987), .A2(n1125), .A3(n1126), .ZN(n975) );
NAND2_X1 U825 ( .A1(n1127), .A2(n1128), .ZN(n1120) );
NAND2_X1 U826 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND3_X1 U827 ( .A1(n1131), .A2(n1132), .A3(n987), .ZN(n1130) );
NAND2_X1 U828 ( .A1(KEYINPUT38), .A2(n1133), .ZN(n1129) );
NAND3_X1 U829 ( .A1(n987), .A2(n1125), .A3(n1134), .ZN(n1086) );
NAND2_X1 U830 ( .A1(n1135), .A2(n1136), .ZN(n1119) );
NAND2_X1 U831 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U832 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
NAND3_X1 U833 ( .A1(n992), .A2(n1141), .A3(n1133), .ZN(n1140) );
INV_X1 U834 ( .A(KEYINPUT38), .ZN(n1139) );
AND4_X1 U835 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n982) );
AND4_X1 U836 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1145) );
NOR2_X1 U837 ( .A1(n1150), .A2(n1151), .ZN(n1144) );
AND2_X1 U838 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
AND2_X1 U839 ( .A1(n1154), .A2(G953), .ZN(n1074) );
XNOR2_X1 U840 ( .A(G952), .B(KEYINPUT36), .ZN(n1154) );
XOR2_X1 U841 ( .A(G146), .B(n1150), .Z(G48) );
AND4_X1 U842 ( .A1(n1155), .A2(n1134), .A3(n1156), .A4(n1157), .ZN(n1150) );
XNOR2_X1 U843 ( .A(G143), .B(n1142), .ZN(G45) );
NAND4_X1 U844 ( .A1(n1155), .A2(n1135), .A3(n1158), .A4(n1159), .ZN(n1142) );
AND3_X1 U845 ( .A1(n1131), .A2(n1160), .A3(n1132), .ZN(n1159) );
XNOR2_X1 U846 ( .A(G140), .B(n1143), .ZN(G42) );
NAND4_X1 U847 ( .A1(n1152), .A2(n1134), .A3(n1008), .A4(n1009), .ZN(n1143) );
XNOR2_X1 U848 ( .A(G137), .B(n1149), .ZN(G39) );
NAND3_X1 U849 ( .A1(n1152), .A2(n1157), .A3(n1161), .ZN(n1149) );
XNOR2_X1 U850 ( .A(G134), .B(n1162), .ZN(G36) );
NAND4_X1 U851 ( .A1(n1163), .A2(KEYINPUT60), .A3(n1164), .A4(n1153), .ZN(n1162) );
NOR2_X1 U852 ( .A1(n1165), .A2(n998), .ZN(n1164) );
XOR2_X1 U853 ( .A(n1160), .B(KEYINPUT63), .Z(n1163) );
XOR2_X1 U854 ( .A(n1148), .B(n1166), .Z(G33) );
NAND2_X1 U855 ( .A1(KEYINPUT13), .A2(G131), .ZN(n1166) );
NAND2_X1 U856 ( .A1(n1152), .A2(n1133), .ZN(n1148) );
AND3_X1 U857 ( .A1(n1155), .A2(n1160), .A3(n989), .ZN(n1152) );
INV_X1 U858 ( .A(n1165), .ZN(n989) );
NAND2_X1 U859 ( .A1(n1014), .A2(n1025), .ZN(n1165) );
XOR2_X1 U860 ( .A(n1022), .B(KEYINPUT40), .Z(n1014) );
INV_X1 U861 ( .A(n998), .ZN(n1155) );
XOR2_X1 U862 ( .A(n1167), .B(KEYINPUT45), .Z(n998) );
XNOR2_X1 U863 ( .A(G128), .B(n1147), .ZN(G30) );
NAND4_X1 U864 ( .A1(n1156), .A2(n1126), .A3(n1167), .A4(n1157), .ZN(n1147) );
XOR2_X1 U865 ( .A(n1124), .B(n1168), .Z(G3) );
XNOR2_X1 U866 ( .A(G101), .B(KEYINPUT12), .ZN(n1168) );
NAND3_X1 U867 ( .A1(n996), .A2(n1125), .A3(n1158), .ZN(n1124) );
AND2_X1 U868 ( .A1(n1167), .A2(n1169), .ZN(n1125) );
XNOR2_X1 U869 ( .A(G125), .B(n1146), .ZN(G27) );
NAND4_X1 U870 ( .A1(n992), .A2(n1134), .A3(n1008), .A4(n1156), .ZN(n1146) );
AND3_X1 U871 ( .A1(n1160), .A2(n1009), .A3(n1135), .ZN(n1156) );
NAND2_X1 U872 ( .A1(n1015), .A2(n1170), .ZN(n1160) );
NAND3_X1 U873 ( .A1(G902), .A2(n1171), .A3(n1046), .ZN(n1170) );
NOR2_X1 U874 ( .A1(n1064), .A2(G900), .ZN(n1046) );
INV_X1 U875 ( .A(n994), .ZN(n1134) );
XNOR2_X1 U876 ( .A(G122), .B(n1172), .ZN(G24) );
NAND4_X1 U877 ( .A1(n1131), .A2(n1132), .A3(n987), .A4(n1173), .ZN(n1172) );
NOR3_X1 U878 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1173) );
NOR2_X1 U879 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
INV_X1 U880 ( .A(KEYINPUT53), .ZN(n1178) );
NOR2_X1 U881 ( .A1(n1135), .A2(n1179), .ZN(n1177) );
NOR2_X1 U882 ( .A1(KEYINPUT53), .A2(n1169), .ZN(n1175) );
NOR2_X1 U883 ( .A1(n1009), .A2(n1157), .ZN(n987) );
XNOR2_X1 U884 ( .A(n1180), .B(n1181), .ZN(G21) );
NOR2_X1 U885 ( .A1(KEYINPUT1), .A2(n1123), .ZN(n1181) );
NAND3_X1 U886 ( .A1(n1161), .A2(n1157), .A3(n1127), .ZN(n1123) );
XNOR2_X1 U887 ( .A(G116), .B(n1122), .ZN(G18) );
NAND2_X1 U888 ( .A1(n1127), .A2(n1153), .ZN(n1122) );
NOR2_X1 U889 ( .A1(n1006), .A2(n995), .ZN(n1153) );
INV_X1 U890 ( .A(n1126), .ZN(n995) );
NOR2_X1 U891 ( .A1(n1132), .A2(n1182), .ZN(n1126) );
AND2_X1 U892 ( .A1(n992), .A2(n1169), .ZN(n1127) );
NOR2_X1 U893 ( .A1(n1011), .A2(n1179), .ZN(n1169) );
INV_X1 U894 ( .A(n1141), .ZN(n1179) );
XNOR2_X1 U895 ( .A(G113), .B(n1183), .ZN(G15) );
NAND4_X1 U896 ( .A1(n1133), .A2(n992), .A3(n1135), .A4(n1184), .ZN(n1183) );
XNOR2_X1 U897 ( .A(KEYINPUT43), .B(n1141), .ZN(n1184) );
INV_X1 U898 ( .A(n1011), .ZN(n1135) );
INV_X1 U899 ( .A(n1174), .ZN(n992) );
NAND2_X1 U900 ( .A1(n1001), .A2(n1185), .ZN(n1174) );
NOR2_X1 U901 ( .A1(n1006), .A2(n994), .ZN(n1133) );
NAND2_X1 U902 ( .A1(n1182), .A2(n1132), .ZN(n994) );
INV_X1 U903 ( .A(n1131), .ZN(n1182) );
INV_X1 U904 ( .A(n1158), .ZN(n1006) );
NOR2_X1 U905 ( .A1(n1009), .A2(n1008), .ZN(n1158) );
XOR2_X1 U906 ( .A(n1186), .B(n1187), .Z(G12) );
XNOR2_X1 U907 ( .A(KEYINPUT21), .B(n1188), .ZN(n1187) );
NOR2_X1 U908 ( .A1(n1189), .A2(n1011), .ZN(n1186) );
NAND2_X1 U909 ( .A1(n1022), .A2(n1025), .ZN(n1011) );
NAND2_X1 U910 ( .A1(G214), .A2(n1190), .ZN(n1025) );
XNOR2_X1 U911 ( .A(n1191), .B(n1192), .ZN(n1022) );
NOR2_X1 U912 ( .A1(n1117), .A2(n1193), .ZN(n1192) );
XNOR2_X1 U913 ( .A(KEYINPUT46), .B(n1190), .ZN(n1193) );
OR2_X1 U914 ( .A1(G902), .A2(G237), .ZN(n1190) );
INV_X1 U915 ( .A(G210), .ZN(n1117) );
NAND2_X1 U916 ( .A1(n1194), .A2(n1195), .ZN(n1191) );
XOR2_X1 U917 ( .A(n1196), .B(n1116), .Z(n1194) );
XNOR2_X1 U918 ( .A(n1197), .B(n1069), .ZN(n1116) );
XNOR2_X1 U919 ( .A(n1188), .B(G122), .ZN(n1069) );
NAND2_X1 U920 ( .A1(KEYINPUT5), .A2(n1067), .ZN(n1197) );
XNOR2_X1 U921 ( .A(n1198), .B(n1199), .ZN(n1067) );
XOR2_X1 U922 ( .A(n1200), .B(n1201), .Z(n1199) );
XNOR2_X1 U923 ( .A(n1202), .B(n1180), .ZN(n1201) );
NAND2_X1 U924 ( .A1(KEYINPUT18), .A2(n1203), .ZN(n1202) );
XNOR2_X1 U925 ( .A(KEYINPUT50), .B(KEYINPUT15), .ZN(n1200) );
XOR2_X1 U926 ( .A(n1204), .B(n1205), .Z(n1198) );
XNOR2_X1 U927 ( .A(n1206), .B(n1207), .ZN(n1205) );
NAND3_X1 U928 ( .A1(n1208), .A2(n1209), .A3(KEYINPUT4), .ZN(n1196) );
NAND2_X1 U929 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
INV_X1 U930 ( .A(KEYINPUT24), .ZN(n1211) );
XOR2_X1 U931 ( .A(n1212), .B(n1213), .Z(n1210) );
NAND2_X1 U932 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
NAND2_X1 U933 ( .A1(n1115), .A2(KEYINPUT24), .ZN(n1208) );
XNOR2_X1 U934 ( .A(n1216), .B(n1215), .ZN(n1115) );
XOR2_X1 U935 ( .A(G125), .B(KEYINPUT28), .Z(n1215) );
XNOR2_X1 U936 ( .A(n1217), .B(n1213), .ZN(n1216) );
AND2_X1 U937 ( .A1(G224), .A2(n1064), .ZN(n1213) );
XOR2_X1 U938 ( .A(n1138), .B(KEYINPUT52), .Z(n1189) );
NAND4_X1 U939 ( .A1(n1161), .A2(n1167), .A3(n1008), .A4(n1141), .ZN(n1138) );
NAND2_X1 U940 ( .A1(n1218), .A2(n1219), .ZN(n1141) );
NAND4_X1 U941 ( .A1(G953), .A2(G902), .A3(n1171), .A4(n1065), .ZN(n1219) );
INV_X1 U942 ( .A(G898), .ZN(n1065) );
XNOR2_X1 U943 ( .A(KEYINPUT19), .B(n1015), .ZN(n1218) );
NAND3_X1 U944 ( .A1(n1171), .A2(n1064), .A3(G952), .ZN(n1015) );
NAND2_X1 U945 ( .A1(G237), .A2(G234), .ZN(n1171) );
INV_X1 U946 ( .A(n1157), .ZN(n1008) );
XOR2_X1 U947 ( .A(n1024), .B(n1027), .Z(n1157) );
INV_X1 U948 ( .A(G472), .ZN(n1027) );
NAND3_X1 U949 ( .A1(n1220), .A2(n1221), .A3(n1195), .ZN(n1024) );
NAND2_X1 U950 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
INV_X1 U951 ( .A(KEYINPUT0), .ZN(n1223) );
XOR2_X1 U952 ( .A(n1224), .B(n1225), .Z(n1222) );
NAND2_X1 U953 ( .A1(KEYINPUT0), .A2(n1226), .ZN(n1220) );
NAND2_X1 U954 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
OR3_X1 U955 ( .A1(n1229), .A2(KEYINPUT10), .A3(n1225), .ZN(n1228) );
INV_X1 U956 ( .A(n1088), .ZN(n1229) );
NAND2_X1 U957 ( .A1(n1224), .A2(n1225), .ZN(n1227) );
XOR2_X1 U958 ( .A(n1092), .B(KEYINPUT14), .Z(n1225) );
XNOR2_X1 U959 ( .A(n1230), .B(n1102), .ZN(n1092) );
XOR2_X1 U960 ( .A(n1054), .B(n1053), .Z(n1102) );
XOR2_X1 U961 ( .A(n1231), .B(n1214), .Z(n1053) );
XOR2_X1 U962 ( .A(n1232), .B(n1233), .Z(n1230) );
NOR2_X1 U963 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U964 ( .A(n1236), .B(KEYINPUT22), .Z(n1235) );
NAND2_X1 U965 ( .A1(G119), .A2(n1204), .ZN(n1236) );
NOR2_X1 U966 ( .A1(G119), .A2(n1204), .ZN(n1234) );
XNOR2_X1 U967 ( .A(G116), .B(KEYINPUT16), .ZN(n1204) );
NAND2_X1 U968 ( .A1(KEYINPUT39), .A2(n1206), .ZN(n1232) );
XNOR2_X1 U969 ( .A(G113), .B(KEYINPUT48), .ZN(n1206) );
AND2_X1 U970 ( .A1(KEYINPUT10), .A2(n1088), .ZN(n1224) );
XOR2_X1 U971 ( .A(n1237), .B(n1203), .Z(n1088) );
INV_X1 U972 ( .A(G101), .ZN(n1203) );
NAND2_X1 U973 ( .A1(G210), .A2(n1238), .ZN(n1237) );
NOR2_X1 U974 ( .A1(n1001), .A2(n1000), .ZN(n1167) );
INV_X1 U975 ( .A(n1185), .ZN(n1000) );
NAND2_X1 U976 ( .A1(G221), .A2(n1239), .ZN(n1185) );
NAND2_X1 U977 ( .A1(G234), .A2(n1195), .ZN(n1239) );
XNOR2_X1 U978 ( .A(n1028), .B(n1240), .ZN(n1001) );
XOR2_X1 U979 ( .A(KEYINPUT9), .B(G469), .Z(n1240) );
NAND2_X1 U980 ( .A1(n1241), .A2(n1195), .ZN(n1028) );
XOR2_X1 U981 ( .A(n1242), .B(n1243), .Z(n1241) );
XNOR2_X1 U982 ( .A(n1231), .B(n1052), .ZN(n1243) );
INV_X1 U983 ( .A(n1054), .ZN(n1052) );
XOR2_X1 U984 ( .A(G134), .B(KEYINPUT8), .Z(n1054) );
XNOR2_X1 U985 ( .A(G131), .B(G137), .ZN(n1231) );
XNOR2_X1 U986 ( .A(n1244), .B(n1245), .ZN(n1242) );
NOR2_X1 U987 ( .A1(KEYINPUT42), .A2(n1246), .ZN(n1245) );
NOR2_X1 U988 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
XOR2_X1 U989 ( .A(KEYINPUT59), .B(n1249), .Z(n1248) );
AND2_X1 U990 ( .A1(n1106), .A2(n1107), .ZN(n1249) );
NOR2_X1 U991 ( .A1(n1107), .A2(n1106), .ZN(n1247) );
XOR2_X1 U992 ( .A(n1188), .B(G140), .Z(n1106) );
NOR2_X1 U993 ( .A1(n1039), .A2(G953), .ZN(n1107) );
INV_X1 U994 ( .A(G227), .ZN(n1039) );
NOR2_X1 U995 ( .A1(KEYINPUT31), .A2(n1250), .ZN(n1244) );
XOR2_X1 U996 ( .A(n1251), .B(n1252), .Z(n1250) );
XNOR2_X1 U997 ( .A(n1214), .B(n1104), .ZN(n1252) );
XOR2_X1 U998 ( .A(G101), .B(n1207), .Z(n1104) );
XOR2_X1 U999 ( .A(G104), .B(G107), .Z(n1207) );
INV_X1 U1000 ( .A(n1217), .ZN(n1214) );
XOR2_X1 U1001 ( .A(G143), .B(n1253), .Z(n1217) );
XOR2_X1 U1002 ( .A(KEYINPUT6), .B(KEYINPUT41), .Z(n1251) );
AND2_X1 U1003 ( .A1(n996), .A2(n1009), .ZN(n1161) );
NAND3_X1 U1004 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1009) );
NAND2_X1 U1005 ( .A1(n1257), .A2(n1077), .ZN(n1256) );
OR3_X1 U1006 ( .A1(n1077), .A2(n1257), .A3(G902), .ZN(n1255) );
NOR2_X1 U1007 ( .A1(n1258), .A2(G234), .ZN(n1257) );
INV_X1 U1008 ( .A(G217), .ZN(n1258) );
XNOR2_X1 U1009 ( .A(n1259), .B(n1260), .ZN(n1077) );
XOR2_X1 U1010 ( .A(n1261), .B(n1262), .Z(n1260) );
XOR2_X1 U1011 ( .A(n1263), .B(n1264), .Z(n1262) );
AND3_X1 U1012 ( .A1(G221), .A2(n1064), .A3(G234), .ZN(n1264) );
NOR2_X1 U1013 ( .A1(G140), .A2(n1265), .ZN(n1263) );
XNOR2_X1 U1014 ( .A(KEYINPUT55), .B(KEYINPUT32), .ZN(n1265) );
XOR2_X1 U1015 ( .A(KEYINPUT27), .B(G125), .Z(n1261) );
XOR2_X1 U1016 ( .A(n1266), .B(n1267), .Z(n1259) );
XNOR2_X1 U1017 ( .A(n1268), .B(n1269), .ZN(n1267) );
NOR2_X1 U1018 ( .A1(G137), .A2(KEYINPUT26), .ZN(n1269) );
NAND2_X1 U1019 ( .A1(KEYINPUT61), .A2(n1188), .ZN(n1268) );
INV_X1 U1020 ( .A(G110), .ZN(n1188) );
XOR2_X1 U1021 ( .A(n1270), .B(n1253), .Z(n1266) );
XOR2_X1 U1022 ( .A(G128), .B(G146), .Z(n1253) );
NAND2_X1 U1023 ( .A1(KEYINPUT7), .A2(n1180), .ZN(n1270) );
INV_X1 U1024 ( .A(G119), .ZN(n1180) );
NAND2_X1 U1025 ( .A1(G902), .A2(G217), .ZN(n1254) );
NOR2_X1 U1026 ( .A1(n1131), .A2(n1132), .ZN(n996) );
XNOR2_X1 U1027 ( .A(n1271), .B(G475), .ZN(n1132) );
NAND2_X1 U1028 ( .A1(n1083), .A2(n1195), .ZN(n1271) );
XOR2_X1 U1029 ( .A(n1272), .B(n1273), .Z(n1083) );
XOR2_X1 U1030 ( .A(G104), .B(n1274), .Z(n1273) );
NOR2_X1 U1031 ( .A1(KEYINPUT34), .A2(n1275), .ZN(n1274) );
XOR2_X1 U1032 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U1033 ( .A(n1278), .B(n1048), .Z(n1277) );
XOR2_X1 U1034 ( .A(G125), .B(G140), .Z(n1048) );
NAND2_X1 U1035 ( .A1(G214), .A2(n1238), .ZN(n1278) );
NOR2_X1 U1036 ( .A1(G953), .A2(G237), .ZN(n1238) );
XNOR2_X1 U1037 ( .A(G131), .B(n1279), .ZN(n1276) );
XOR2_X1 U1038 ( .A(G146), .B(G143), .Z(n1279) );
XNOR2_X1 U1039 ( .A(G113), .B(G122), .ZN(n1272) );
XNOR2_X1 U1040 ( .A(n1280), .B(G478), .ZN(n1131) );
NAND2_X1 U1041 ( .A1(n1081), .A2(n1195), .ZN(n1280) );
INV_X1 U1042 ( .A(G902), .ZN(n1195) );
XOR2_X1 U1043 ( .A(n1281), .B(n1282), .Z(n1081) );
XOR2_X1 U1044 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U1045 ( .A(G128), .B(G122), .Z(n1284) );
XNOR2_X1 U1046 ( .A(KEYINPUT62), .B(n1285), .ZN(n1283) );
INV_X1 U1047 ( .A(G134), .ZN(n1285) );
XOR2_X1 U1048 ( .A(n1286), .B(n1287), .Z(n1281) );
XOR2_X1 U1049 ( .A(G116), .B(n1288), .Z(n1287) );
AND3_X1 U1050 ( .A1(G234), .A2(n1064), .A3(G217), .ZN(n1288) );
INV_X1 U1051 ( .A(G953), .ZN(n1064) );
XNOR2_X1 U1052 ( .A(n1289), .B(n1290), .ZN(n1286) );
NOR2_X1 U1053 ( .A1(G107), .A2(KEYINPUT56), .ZN(n1290) );
NOR2_X1 U1054 ( .A1(G143), .A2(KEYINPUT37), .ZN(n1289) );
endmodule


