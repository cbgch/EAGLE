//Key = 0110000100001110000010001010111001110001101001101100011100100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395;

XOR2_X1 U775 ( .A(n1059), .B(n1060), .Z(G9) );
NOR2_X1 U776 ( .A1(KEYINPUT4), .A2(n1061), .ZN(n1060) );
NOR4_X1 U777 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1059) );
NOR2_X1 U778 ( .A1(KEYINPUT35), .A2(n1066), .ZN(n1063) );
NOR3_X1 U779 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
NOR2_X1 U780 ( .A1(n1070), .A2(n1071), .ZN(n1062) );
INV_X1 U781 ( .A(KEYINPUT35), .ZN(n1071) );
NOR2_X1 U782 ( .A1(n1072), .A2(n1073), .ZN(G75) );
XOR2_X1 U783 ( .A(n1074), .B(KEYINPUT29), .Z(n1073) );
NAND3_X1 U784 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1074) );
XOR2_X1 U785 ( .A(KEYINPUT14), .B(G952), .Z(n1077) );
NOR4_X1 U786 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1072) );
XOR2_X1 U787 ( .A(KEYINPUT23), .B(n1082), .Z(n1079) );
NOR2_X1 U788 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U789 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NOR3_X1 U790 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NOR2_X1 U791 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U792 ( .A1(n1092), .A2(n1064), .ZN(n1091) );
NOR3_X1 U793 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
NOR3_X1 U794 ( .A1(n1096), .A2(KEYINPUT58), .A3(n1097), .ZN(n1095) );
NOR2_X1 U795 ( .A1(n1098), .A2(n1099), .ZN(n1094) );
NOR2_X1 U796 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
AND2_X1 U797 ( .A1(n1102), .A2(KEYINPUT58), .ZN(n1100) );
NOR2_X1 U798 ( .A1(n1103), .A2(n1104), .ZN(n1093) );
NOR2_X1 U799 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NOR2_X1 U800 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
NOR3_X1 U801 ( .A1(n1104), .A2(n1109), .A3(n1099), .ZN(n1090) );
NOR2_X1 U802 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR4_X1 U803 ( .A1(n1112), .A2(n1064), .A3(n1099), .A4(n1104), .ZN(n1085) );
INV_X1 U804 ( .A(n1113), .ZN(n1064) );
NOR2_X1 U805 ( .A1(n1114), .A2(n1069), .ZN(n1112) );
INV_X1 U806 ( .A(n1115), .ZN(n1069) );
NOR2_X1 U807 ( .A1(n1087), .A2(n1116), .ZN(n1114) );
NAND3_X1 U808 ( .A1(n1075), .A2(n1076), .A3(G952), .ZN(n1078) );
NAND4_X1 U809 ( .A1(n1116), .A2(n1107), .A3(n1117), .A4(n1118), .ZN(n1075) );
NOR4_X1 U810 ( .A1(n1104), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1118) );
XOR2_X1 U811 ( .A(KEYINPUT31), .B(n1122), .Z(n1121) );
XNOR2_X1 U812 ( .A(n1123), .B(n1124), .ZN(n1120) );
INV_X1 U813 ( .A(n1125), .ZN(n1104) );
NOR3_X1 U814 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1117) );
XOR2_X1 U815 ( .A(n1129), .B(n1130), .Z(G72) );
XOR2_X1 U816 ( .A(n1131), .B(n1132), .Z(n1130) );
AND2_X1 U817 ( .A1(n1081), .A2(n1076), .ZN(n1132) );
NOR2_X1 U818 ( .A1(KEYINPUT37), .A2(n1133), .ZN(n1131) );
NOR2_X1 U819 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U820 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND3_X1 U821 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1136) );
NAND2_X1 U822 ( .A1(KEYINPUT59), .A2(n1141), .ZN(n1140) );
OR3_X1 U823 ( .A1(n1141), .A2(KEYINPUT59), .A3(n1142), .ZN(n1139) );
NAND2_X1 U824 ( .A1(n1142), .A2(n1143), .ZN(n1138) );
NAND2_X1 U825 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
INV_X1 U826 ( .A(KEYINPUT59), .ZN(n1145) );
XNOR2_X1 U827 ( .A(n1141), .B(KEYINPUT27), .ZN(n1144) );
XOR2_X1 U828 ( .A(n1146), .B(n1147), .Z(n1141) );
NAND2_X1 U829 ( .A1(n1148), .A2(KEYINPUT42), .ZN(n1146) );
XNOR2_X1 U830 ( .A(n1149), .B(n1150), .ZN(n1148) );
NAND2_X1 U831 ( .A1(KEYINPUT2), .A2(n1151), .ZN(n1149) );
NOR2_X1 U832 ( .A1(G900), .A2(n1076), .ZN(n1134) );
NAND2_X1 U833 ( .A1(G953), .A2(n1152), .ZN(n1129) );
NAND2_X1 U834 ( .A1(G900), .A2(G227), .ZN(n1152) );
XOR2_X1 U835 ( .A(n1153), .B(n1154), .Z(G69) );
NOR2_X1 U836 ( .A1(n1155), .A2(n1076), .ZN(n1154) );
NOR2_X1 U837 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U838 ( .A(n1158), .B(n1159), .Z(n1153) );
NOR2_X1 U839 ( .A1(KEYINPUT17), .A2(n1160), .ZN(n1159) );
NOR2_X1 U840 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XNOR2_X1 U841 ( .A(n1163), .B(n1164), .ZN(n1162) );
XNOR2_X1 U842 ( .A(n1165), .B(n1166), .ZN(n1164) );
NOR2_X1 U843 ( .A1(KEYINPUT61), .A2(n1167), .ZN(n1166) );
NOR2_X1 U844 ( .A1(KEYINPUT25), .A2(n1168), .ZN(n1165) );
NOR2_X1 U845 ( .A1(G898), .A2(n1076), .ZN(n1161) );
NAND2_X1 U846 ( .A1(n1169), .A2(n1080), .ZN(n1158) );
XNOR2_X1 U847 ( .A(KEYINPUT13), .B(n1076), .ZN(n1169) );
NOR2_X1 U848 ( .A1(n1170), .A2(n1171), .ZN(G66) );
XOR2_X1 U849 ( .A(n1172), .B(n1173), .Z(n1171) );
NAND2_X1 U850 ( .A1(n1174), .A2(n1175), .ZN(n1172) );
NOR2_X1 U851 ( .A1(n1170), .A2(n1176), .ZN(G63) );
NOR2_X1 U852 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XOR2_X1 U853 ( .A(KEYINPUT62), .B(n1179), .Z(n1178) );
NOR2_X1 U854 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
AND2_X1 U855 ( .A1(n1181), .A2(n1180), .ZN(n1177) );
NAND2_X1 U856 ( .A1(n1174), .A2(G478), .ZN(n1181) );
NOR2_X1 U857 ( .A1(n1170), .A2(n1182), .ZN(G60) );
XOR2_X1 U858 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND2_X1 U859 ( .A1(n1174), .A2(G475), .ZN(n1183) );
XOR2_X1 U860 ( .A(n1185), .B(n1186), .Z(G6) );
NAND2_X1 U861 ( .A1(KEYINPUT30), .A2(n1187), .ZN(n1185) );
NOR2_X1 U862 ( .A1(n1170), .A2(n1188), .ZN(G57) );
XOR2_X1 U863 ( .A(n1189), .B(n1190), .Z(n1188) );
XNOR2_X1 U864 ( .A(G101), .B(n1191), .ZN(n1190) );
NAND2_X1 U865 ( .A1(n1174), .A2(G472), .ZN(n1191) );
XOR2_X1 U866 ( .A(n1192), .B(n1193), .Z(n1189) );
NOR2_X1 U867 ( .A1(n1170), .A2(n1194), .ZN(G54) );
XOR2_X1 U868 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U869 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U870 ( .A(n1199), .B(n1200), .Z(n1195) );
XNOR2_X1 U871 ( .A(n1201), .B(n1202), .ZN(n1200) );
NAND2_X1 U872 ( .A1(n1174), .A2(G469), .ZN(n1201) );
NOR2_X1 U873 ( .A1(n1170), .A2(n1203), .ZN(G51) );
XOR2_X1 U874 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U875 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U876 ( .A(n1208), .B(n1209), .Z(n1204) );
XNOR2_X1 U877 ( .A(G125), .B(n1210), .ZN(n1209) );
NAND2_X1 U878 ( .A1(n1174), .A2(n1124), .ZN(n1208) );
INV_X1 U879 ( .A(n1211), .ZN(n1124) );
AND2_X1 U880 ( .A1(G902), .A2(n1212), .ZN(n1174) );
OR2_X1 U881 ( .A1(n1081), .A2(n1080), .ZN(n1212) );
NAND4_X1 U882 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1080) );
AND4_X1 U883 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1216) );
NAND2_X1 U884 ( .A1(KEYINPUT40), .A2(n1186), .ZN(n1215) );
AND3_X1 U885 ( .A1(n1102), .A2(n1113), .A3(n1070), .ZN(n1186) );
NAND2_X1 U886 ( .A1(n1113), .A2(n1221), .ZN(n1214) );
NAND2_X1 U887 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NAND3_X1 U888 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1223) );
NAND2_X1 U889 ( .A1(n1070), .A2(n1227), .ZN(n1222) );
NAND2_X1 U890 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
OR2_X1 U891 ( .A1(n1065), .A2(KEYINPUT11), .ZN(n1229) );
OR2_X1 U892 ( .A1(n1102), .A2(KEYINPUT40), .ZN(n1228) );
NAND2_X1 U893 ( .A1(n1101), .A2(n1230), .ZN(n1213) );
NAND2_X1 U894 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND3_X1 U895 ( .A1(n1115), .A2(n1233), .A3(n1234), .ZN(n1232) );
NAND2_X1 U896 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NAND3_X1 U897 ( .A1(n1106), .A2(n1113), .A3(KEYINPUT11), .ZN(n1236) );
NAND3_X1 U898 ( .A1(n1111), .A2(n1237), .A3(n1096), .ZN(n1235) );
OR2_X1 U899 ( .A1(n1237), .A2(n1238), .ZN(n1231) );
INV_X1 U900 ( .A(KEYINPUT34), .ZN(n1237) );
NAND4_X1 U901 ( .A1(n1239), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1081) );
AND4_X1 U902 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1242) );
NOR2_X1 U903 ( .A1(n1247), .A2(n1248), .ZN(n1241) );
NOR2_X1 U904 ( .A1(n1076), .A2(G952), .ZN(n1170) );
XNOR2_X1 U905 ( .A(G146), .B(n1239), .ZN(G48) );
NAND3_X1 U906 ( .A1(n1249), .A2(n1102), .A3(n1250), .ZN(n1239) );
NAND3_X1 U907 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(G45) );
NAND2_X1 U908 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U909 ( .A1(KEYINPUT15), .A2(n1256), .ZN(n1252) );
NAND2_X1 U910 ( .A1(n1257), .A2(G143), .ZN(n1256) );
XNOR2_X1 U911 ( .A(n1254), .B(KEYINPUT16), .ZN(n1257) );
NAND2_X1 U912 ( .A1(n1258), .A2(n1259), .ZN(n1251) );
INV_X1 U913 ( .A(KEYINPUT15), .ZN(n1259) );
NAND2_X1 U914 ( .A1(n1260), .A2(n1261), .ZN(n1258) );
OR3_X1 U915 ( .A1(n1255), .A2(n1254), .A3(KEYINPUT16), .ZN(n1261) );
NAND2_X1 U916 ( .A1(KEYINPUT16), .A2(n1254), .ZN(n1260) );
INV_X1 U917 ( .A(n1240), .ZN(n1254) );
NAND4_X1 U918 ( .A1(n1249), .A2(n1111), .A3(n1224), .A4(n1225), .ZN(n1240) );
XOR2_X1 U919 ( .A(G140), .B(n1248), .Z(G42) );
AND3_X1 U920 ( .A1(n1102), .A2(n1110), .A3(n1262), .ZN(n1248) );
XOR2_X1 U921 ( .A(n1247), .B(n1263), .Z(G39) );
NOR2_X1 U922 ( .A1(KEYINPUT50), .A2(n1150), .ZN(n1263) );
AND3_X1 U923 ( .A1(n1262), .A2(n1250), .A3(n1125), .ZN(n1247) );
XOR2_X1 U924 ( .A(n1246), .B(n1264), .Z(G36) );
NOR2_X1 U925 ( .A1(G134), .A2(KEYINPUT43), .ZN(n1264) );
NAND3_X1 U926 ( .A1(n1101), .A2(n1111), .A3(n1262), .ZN(n1246) );
XNOR2_X1 U927 ( .A(G131), .B(n1245), .ZN(G33) );
NAND3_X1 U928 ( .A1(n1102), .A2(n1111), .A3(n1262), .ZN(n1245) );
NOR3_X1 U929 ( .A1(n1265), .A2(n1088), .A3(n1087), .ZN(n1262) );
INV_X1 U930 ( .A(n1116), .ZN(n1088) );
XNOR2_X1 U931 ( .A(G128), .B(n1244), .ZN(G30) );
NAND3_X1 U932 ( .A1(n1249), .A2(n1101), .A3(n1250), .ZN(n1244) );
INV_X1 U933 ( .A(n1065), .ZN(n1101) );
NOR2_X1 U934 ( .A1(n1265), .A2(n1115), .ZN(n1249) );
NAND2_X1 U935 ( .A1(n1106), .A2(n1266), .ZN(n1265) );
NAND2_X1 U936 ( .A1(n1267), .A2(n1084), .ZN(n1266) );
INV_X1 U937 ( .A(n1067), .ZN(n1106) );
XNOR2_X1 U938 ( .A(G101), .B(n1220), .ZN(G3) );
NAND3_X1 U939 ( .A1(n1125), .A2(n1111), .A3(n1070), .ZN(n1220) );
XNOR2_X1 U940 ( .A(n1268), .B(n1269), .ZN(G27) );
NOR2_X1 U941 ( .A1(KEYINPUT19), .A2(n1243), .ZN(n1269) );
NAND4_X1 U942 ( .A1(n1096), .A2(n1102), .A3(n1270), .A4(n1110), .ZN(n1243) );
NOR2_X1 U943 ( .A1(n1271), .A2(n1115), .ZN(n1270) );
AND2_X1 U944 ( .A1(n1084), .A2(n1267), .ZN(n1271) );
NAND4_X1 U945 ( .A1(n1272), .A2(G953), .A3(G902), .A4(n1273), .ZN(n1267) );
XNOR2_X1 U946 ( .A(G900), .B(KEYINPUT22), .ZN(n1272) );
INV_X1 U947 ( .A(n1099), .ZN(n1096) );
XNOR2_X1 U948 ( .A(G122), .B(n1274), .ZN(G24) );
NAND3_X1 U949 ( .A1(KEYINPUT24), .A2(n1226), .A3(n1275), .ZN(n1274) );
AND3_X1 U950 ( .A1(n1224), .A2(n1225), .A3(n1113), .ZN(n1275) );
NAND2_X1 U951 ( .A1(n1276), .A2(n1277), .ZN(n1113) );
NAND2_X1 U952 ( .A1(n1111), .A2(n1278), .ZN(n1277) );
INV_X1 U953 ( .A(KEYINPUT12), .ZN(n1278) );
NAND3_X1 U954 ( .A1(n1279), .A2(n1280), .A3(KEYINPUT12), .ZN(n1276) );
XNOR2_X1 U955 ( .A(G119), .B(n1219), .ZN(G21) );
NAND3_X1 U956 ( .A1(n1125), .A2(n1250), .A3(n1226), .ZN(n1219) );
NOR2_X1 U957 ( .A1(n1280), .A2(n1279), .ZN(n1250) );
INV_X1 U958 ( .A(n1119), .ZN(n1280) );
XOR2_X1 U959 ( .A(G116), .B(n1281), .Z(G18) );
NOR2_X1 U960 ( .A1(n1065), .A2(n1238), .ZN(n1281) );
NAND2_X1 U961 ( .A1(n1282), .A2(n1224), .ZN(n1065) );
XNOR2_X1 U962 ( .A(n1283), .B(KEYINPUT49), .ZN(n1224) );
XOR2_X1 U963 ( .A(n1284), .B(KEYINPUT3), .Z(n1282) );
XNOR2_X1 U964 ( .A(G113), .B(n1218), .ZN(G15) );
OR2_X1 U965 ( .A1(n1238), .A2(n1097), .ZN(n1218) );
INV_X1 U966 ( .A(n1102), .ZN(n1097) );
NOR2_X1 U967 ( .A1(n1283), .A2(n1284), .ZN(n1102) );
NAND2_X1 U968 ( .A1(n1226), .A2(n1111), .ZN(n1238) );
NOR2_X1 U969 ( .A1(n1119), .A2(n1279), .ZN(n1111) );
NOR3_X1 U970 ( .A1(n1115), .A2(n1068), .A3(n1099), .ZN(n1226) );
NAND2_X1 U971 ( .A1(n1285), .A2(n1286), .ZN(n1099) );
XNOR2_X1 U972 ( .A(G110), .B(n1217), .ZN(G12) );
NAND3_X1 U973 ( .A1(n1125), .A2(n1110), .A3(n1070), .ZN(n1217) );
NOR3_X1 U974 ( .A1(n1067), .A2(n1068), .A3(n1115), .ZN(n1070) );
NAND2_X1 U975 ( .A1(n1087), .A2(n1116), .ZN(n1115) );
NAND2_X1 U976 ( .A1(G214), .A2(n1287), .ZN(n1116) );
NAND3_X1 U977 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n1087) );
NAND2_X1 U978 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
OR3_X1 U979 ( .A1(n1292), .A2(n1291), .A3(n1211), .ZN(n1289) );
INV_X1 U980 ( .A(KEYINPUT63), .ZN(n1292) );
NAND2_X1 U981 ( .A1(n1293), .A2(n1211), .ZN(n1288) );
NAND2_X1 U982 ( .A1(G210), .A2(n1287), .ZN(n1211) );
NAND2_X1 U983 ( .A1(n1294), .A2(n1295), .ZN(n1287) );
INV_X1 U984 ( .A(G237), .ZN(n1294) );
NAND2_X1 U985 ( .A1(n1296), .A2(KEYINPUT63), .ZN(n1293) );
XNOR2_X1 U986 ( .A(n1291), .B(KEYINPUT38), .ZN(n1296) );
XNOR2_X1 U987 ( .A(n1123), .B(KEYINPUT36), .ZN(n1291) );
NAND2_X1 U988 ( .A1(n1297), .A2(n1295), .ZN(n1123) );
XNOR2_X1 U989 ( .A(n1298), .B(n1206), .ZN(n1297) );
XNOR2_X1 U990 ( .A(n1299), .B(n1168), .ZN(n1206) );
XOR2_X1 U991 ( .A(G110), .B(n1300), .Z(n1168) );
NOR2_X1 U992 ( .A1(KEYINPUT51), .A2(n1301), .ZN(n1300) );
NAND2_X1 U993 ( .A1(KEYINPUT55), .A2(n1302), .ZN(n1299) );
XNOR2_X1 U994 ( .A(n1167), .B(n1303), .ZN(n1302) );
INV_X1 U995 ( .A(n1163), .ZN(n1303) );
XNOR2_X1 U996 ( .A(n1304), .B(KEYINPUT10), .ZN(n1163) );
NAND2_X1 U997 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XOR2_X1 U998 ( .A(n1307), .B(G113), .Z(n1167) );
NAND2_X1 U999 ( .A1(n1308), .A2(KEYINPUT53), .ZN(n1298) );
XOR2_X1 U1000 ( .A(n1309), .B(n1310), .Z(n1308) );
XNOR2_X1 U1001 ( .A(n1268), .B(n1210), .ZN(n1310) );
NOR2_X1 U1002 ( .A1(n1156), .A2(G953), .ZN(n1210) );
INV_X1 U1003 ( .A(G224), .ZN(n1156) );
NAND2_X1 U1004 ( .A1(KEYINPUT54), .A2(n1207), .ZN(n1309) );
INV_X1 U1005 ( .A(n1233), .ZN(n1068) );
NAND2_X1 U1006 ( .A1(n1084), .A2(n1311), .ZN(n1233) );
NAND4_X1 U1007 ( .A1(G953), .A2(G902), .A3(n1273), .A4(n1157), .ZN(n1311) );
INV_X1 U1008 ( .A(G898), .ZN(n1157) );
NAND3_X1 U1009 ( .A1(n1273), .A2(n1076), .A3(G952), .ZN(n1084) );
NAND2_X1 U1010 ( .A1(G237), .A2(G234), .ZN(n1273) );
NAND2_X1 U1011 ( .A1(n1285), .A2(n1108), .ZN(n1067) );
INV_X1 U1012 ( .A(n1286), .ZN(n1108) );
NOR2_X1 U1013 ( .A1(n1312), .A2(n1122), .ZN(n1286) );
NOR3_X1 U1014 ( .A1(G469), .A2(G902), .A3(n1313), .ZN(n1122) );
XNOR2_X1 U1015 ( .A(KEYINPUT45), .B(n1126), .ZN(n1312) );
AND2_X1 U1016 ( .A1(G469), .A2(n1314), .ZN(n1126) );
OR2_X1 U1017 ( .A1(n1313), .A2(G902), .ZN(n1314) );
XNOR2_X1 U1018 ( .A(n1315), .B(n1199), .ZN(n1313) );
XOR2_X1 U1019 ( .A(G140), .B(n1316), .Z(n1199) );
AND2_X1 U1020 ( .A1(n1076), .A2(G227), .ZN(n1316) );
XOR2_X1 U1021 ( .A(n1317), .B(G110), .Z(n1315) );
NAND2_X1 U1022 ( .A1(KEYINPUT26), .A2(n1318), .ZN(n1317) );
XOR2_X1 U1023 ( .A(n1319), .B(n1197), .Z(n1318) );
XNOR2_X1 U1024 ( .A(n1320), .B(n1321), .ZN(n1197) );
NAND3_X1 U1025 ( .A1(n1322), .A2(n1323), .A3(n1306), .ZN(n1320) );
NAND2_X1 U1026 ( .A1(n1324), .A2(G104), .ZN(n1306) );
NAND2_X1 U1027 ( .A1(KEYINPUT41), .A2(n1325), .ZN(n1323) );
NAND3_X1 U1028 ( .A1(n1326), .A2(n1327), .A3(n1328), .ZN(n1325) );
INV_X1 U1029 ( .A(n1324), .ZN(n1328) );
NOR2_X1 U1030 ( .A1(n1329), .A2(G107), .ZN(n1324) );
NAND3_X1 U1031 ( .A1(G107), .A2(n1329), .A3(n1187), .ZN(n1327) );
NAND2_X1 U1032 ( .A1(G101), .A2(G104), .ZN(n1326) );
OR2_X1 U1033 ( .A1(n1305), .A2(KEYINPUT41), .ZN(n1322) );
AND2_X1 U1034 ( .A1(n1330), .A2(n1331), .ZN(n1305) );
NAND3_X1 U1035 ( .A1(n1329), .A2(n1187), .A3(n1061), .ZN(n1331) );
INV_X1 U1036 ( .A(G101), .ZN(n1329) );
NAND2_X1 U1037 ( .A1(n1332), .A2(G107), .ZN(n1330) );
XNOR2_X1 U1038 ( .A(n1187), .B(G101), .ZN(n1332) );
NOR2_X1 U1039 ( .A1(KEYINPUT21), .A2(n1333), .ZN(n1319) );
INV_X1 U1040 ( .A(n1142), .ZN(n1333) );
XOR2_X1 U1041 ( .A(G128), .B(n1202), .Z(n1142) );
XOR2_X1 U1042 ( .A(KEYINPUT18), .B(n1107), .Z(n1285) );
NAND2_X1 U1043 ( .A1(G221), .A2(n1334), .ZN(n1107) );
AND2_X1 U1044 ( .A1(n1279), .A2(n1119), .ZN(n1110) );
XNOR2_X1 U1045 ( .A(n1335), .B(n1175), .ZN(n1119) );
AND2_X1 U1046 ( .A1(G217), .A2(n1334), .ZN(n1175) );
NAND2_X1 U1047 ( .A1(G234), .A2(n1295), .ZN(n1334) );
NAND2_X1 U1048 ( .A1(n1173), .A2(n1295), .ZN(n1335) );
XOR2_X1 U1049 ( .A(n1336), .B(n1337), .Z(n1173) );
XOR2_X1 U1050 ( .A(G119), .B(n1338), .Z(n1337) );
XNOR2_X1 U1051 ( .A(KEYINPUT9), .B(n1150), .ZN(n1338) );
XOR2_X1 U1052 ( .A(n1339), .B(n1198), .Z(n1336) );
XNOR2_X1 U1053 ( .A(G110), .B(n1340), .ZN(n1198) );
XOR2_X1 U1054 ( .A(n1341), .B(n1342), .Z(n1339) );
AND3_X1 U1055 ( .A1(G221), .A2(n1076), .A3(G234), .ZN(n1342) );
NAND3_X1 U1056 ( .A1(n1343), .A2(n1344), .A3(n1345), .ZN(n1341) );
NAND2_X1 U1057 ( .A1(KEYINPUT6), .A2(n1137), .ZN(n1345) );
NAND3_X1 U1058 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1344) );
INV_X1 U1059 ( .A(KEYINPUT6), .ZN(n1347) );
OR2_X1 U1060 ( .A1(n1348), .A2(n1346), .ZN(n1343) );
NOR2_X1 U1061 ( .A1(KEYINPUT52), .A2(n1137), .ZN(n1346) );
INV_X1 U1062 ( .A(G146), .ZN(n1348) );
NOR2_X1 U1063 ( .A1(n1349), .A2(n1128), .ZN(n1279) );
NOR2_X1 U1064 ( .A1(n1350), .A2(n1351), .ZN(n1128) );
XOR2_X1 U1065 ( .A(n1127), .B(KEYINPUT5), .Z(n1349) );
AND2_X1 U1066 ( .A1(n1351), .A2(n1350), .ZN(n1127) );
NAND2_X1 U1067 ( .A1(n1352), .A2(n1295), .ZN(n1350) );
XOR2_X1 U1068 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1069 ( .A(KEYINPUT48), .B(n1355), .Z(n1354) );
NOR2_X1 U1070 ( .A1(G101), .A2(KEYINPUT56), .ZN(n1355) );
XOR2_X1 U1071 ( .A(n1192), .B(n1356), .Z(n1353) );
NOR2_X1 U1072 ( .A1(KEYINPUT8), .A2(n1193), .ZN(n1356) );
XOR2_X1 U1073 ( .A(G113), .B(n1357), .Z(n1193) );
NOR2_X1 U1074 ( .A1(KEYINPUT47), .A2(n1307), .ZN(n1357) );
XOR2_X1 U1075 ( .A(G116), .B(n1358), .Z(n1307) );
XOR2_X1 U1076 ( .A(KEYINPUT1), .B(G119), .Z(n1358) );
XOR2_X1 U1077 ( .A(n1359), .B(n1321), .Z(n1192) );
XNOR2_X1 U1078 ( .A(n1147), .B(n1360), .ZN(n1321) );
NOR2_X1 U1079 ( .A1(KEYINPUT44), .A2(n1361), .ZN(n1360) );
XNOR2_X1 U1080 ( .A(n1362), .B(n1150), .ZN(n1361) );
INV_X1 U1081 ( .A(G137), .ZN(n1150) );
NAND2_X1 U1082 ( .A1(KEYINPUT28), .A2(n1151), .ZN(n1362) );
XNOR2_X1 U1083 ( .A(n1207), .B(n1363), .ZN(n1359) );
AND2_X1 U1084 ( .A1(n1364), .A2(G210), .ZN(n1363) );
XNOR2_X1 U1085 ( .A(n1365), .B(n1202), .ZN(n1207) );
XOR2_X1 U1086 ( .A(G146), .B(G143), .Z(n1202) );
NAND2_X1 U1087 ( .A1(KEYINPUT20), .A2(n1340), .ZN(n1365) );
INV_X1 U1088 ( .A(G128), .ZN(n1340) );
XOR2_X1 U1089 ( .A(G472), .B(KEYINPUT60), .Z(n1351) );
NOR2_X1 U1090 ( .A1(n1225), .A2(n1283), .ZN(n1125) );
XNOR2_X1 U1091 ( .A(n1366), .B(G478), .ZN(n1283) );
NAND2_X1 U1092 ( .A1(n1180), .A2(n1295), .ZN(n1366) );
XNOR2_X1 U1093 ( .A(n1367), .B(n1368), .ZN(n1180) );
XOR2_X1 U1094 ( .A(n1369), .B(n1370), .Z(n1368) );
XNOR2_X1 U1095 ( .A(n1151), .B(G128), .ZN(n1370) );
INV_X1 U1096 ( .A(G134), .ZN(n1151) );
XNOR2_X1 U1097 ( .A(KEYINPUT46), .B(n1255), .ZN(n1369) );
XOR2_X1 U1098 ( .A(n1371), .B(n1372), .Z(n1367) );
XNOR2_X1 U1099 ( .A(G116), .B(n1061), .ZN(n1372) );
INV_X1 U1100 ( .A(G107), .ZN(n1061) );
XOR2_X1 U1101 ( .A(n1373), .B(n1374), .Z(n1371) );
AND3_X1 U1102 ( .A1(G234), .A2(n1076), .A3(G217), .ZN(n1374) );
INV_X1 U1103 ( .A(G953), .ZN(n1076) );
NAND2_X1 U1104 ( .A1(KEYINPUT7), .A2(n1375), .ZN(n1373) );
INV_X1 U1105 ( .A(n1284), .ZN(n1225) );
XOR2_X1 U1106 ( .A(n1376), .B(G475), .Z(n1284) );
NAND2_X1 U1107 ( .A1(n1184), .A2(n1295), .ZN(n1376) );
INV_X1 U1108 ( .A(G902), .ZN(n1295) );
XNOR2_X1 U1109 ( .A(n1377), .B(n1378), .ZN(n1184) );
XNOR2_X1 U1110 ( .A(n1187), .B(n1379), .ZN(n1378) );
XOR2_X1 U1111 ( .A(KEYINPUT33), .B(G113), .Z(n1379) );
INV_X1 U1112 ( .A(G104), .ZN(n1187) );
XNOR2_X1 U1113 ( .A(n1380), .B(n1301), .ZN(n1377) );
INV_X1 U1114 ( .A(n1375), .ZN(n1301) );
XOR2_X1 U1115 ( .A(G122), .B(KEYINPUT39), .Z(n1375) );
XOR2_X1 U1116 ( .A(n1381), .B(n1382), .Z(n1380) );
NOR2_X1 U1117 ( .A1(KEYINPUT57), .A2(n1383), .ZN(n1382) );
XNOR2_X1 U1118 ( .A(G146), .B(n1137), .ZN(n1383) );
XOR2_X1 U1119 ( .A(G140), .B(n1268), .Z(n1137) );
INV_X1 U1120 ( .A(G125), .ZN(n1268) );
NAND3_X1 U1121 ( .A1(n1384), .A2(n1385), .A3(n1386), .ZN(n1381) );
NAND2_X1 U1122 ( .A1(n1387), .A2(n1147), .ZN(n1386) );
NAND2_X1 U1123 ( .A1(KEYINPUT0), .A2(n1388), .ZN(n1385) );
NAND2_X1 U1124 ( .A1(n1389), .A2(n1390), .ZN(n1388) );
XNOR2_X1 U1125 ( .A(KEYINPUT32), .B(n1147), .ZN(n1390) );
INV_X1 U1126 ( .A(n1387), .ZN(n1389) );
NAND2_X1 U1127 ( .A1(n1391), .A2(n1392), .ZN(n1384) );
INV_X1 U1128 ( .A(KEYINPUT0), .ZN(n1392) );
NAND2_X1 U1129 ( .A1(n1393), .A2(n1394), .ZN(n1391) );
NAND2_X1 U1130 ( .A1(KEYINPUT32), .A2(n1147), .ZN(n1394) );
OR3_X1 U1131 ( .A1(n1387), .A2(KEYINPUT32), .A3(n1147), .ZN(n1393) );
INV_X1 U1132 ( .A(G131), .ZN(n1147) );
XOR2_X1 U1133 ( .A(n1395), .B(n1255), .Z(n1387) );
INV_X1 U1134 ( .A(G143), .ZN(n1255) );
NAND2_X1 U1135 ( .A1(G214), .A2(n1364), .ZN(n1395) );
NOR2_X1 U1136 ( .A1(G953), .A2(G237), .ZN(n1364) );
endmodule


