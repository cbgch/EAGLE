//Key = 0101001110011001110010011000000000000110111001001110010111011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343;

XOR2_X1 U736 ( .A(n1028), .B(n1029), .Z(G9) );
XNOR2_X1 U737 ( .A(G107), .B(KEYINPUT16), .ZN(n1028) );
NOR2_X1 U738 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U739 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
NOR2_X1 U740 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR3_X1 U741 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1036) );
NOR3_X1 U742 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NOR3_X1 U743 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1039) );
NOR2_X1 U744 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U745 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U746 ( .A1(n1051), .A2(n1052), .ZN(n1047) );
NOR2_X1 U747 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U748 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U749 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
XOR2_X1 U750 ( .A(n1059), .B(KEYINPUT37), .Z(n1038) );
NAND2_X1 U751 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U752 ( .A1(n1062), .A2(n1063), .ZN(n1034) );
XOR2_X1 U753 ( .A(KEYINPUT1), .B(n1064), .Z(n1063) );
NAND3_X1 U754 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1032) );
NAND3_X1 U755 ( .A1(n1068), .A2(n1069), .A3(n1064), .ZN(n1067) );
NOR2_X1 U756 ( .A1(n1041), .A2(n1046), .ZN(n1064) );
INV_X1 U757 ( .A(n1070), .ZN(n1046) );
INV_X1 U758 ( .A(n1060), .ZN(n1041) );
NOR4_X1 U759 ( .A1(n1044), .A2(n1050), .A3(n1052), .A4(n1056), .ZN(n1060) );
NOR3_X1 U760 ( .A1(n1071), .A2(G953), .A3(G952), .ZN(n1030) );
INV_X1 U761 ( .A(n1065), .ZN(n1071) );
NAND4_X1 U762 ( .A1(n1072), .A2(n1070), .A3(n1073), .A4(n1074), .ZN(n1065) );
NOR4_X1 U763 ( .A1(n1069), .A2(n1075), .A3(n1052), .A4(n1076), .ZN(n1074) );
XNOR2_X1 U764 ( .A(n1077), .B(KEYINPUT41), .ZN(n1075) );
XNOR2_X1 U765 ( .A(G475), .B(n1078), .ZN(n1073) );
NOR2_X1 U766 ( .A1(KEYINPUT32), .A2(n1079), .ZN(n1078) );
XOR2_X1 U767 ( .A(n1080), .B(n1081), .Z(n1072) );
XNOR2_X1 U768 ( .A(KEYINPUT10), .B(n1082), .ZN(n1080) );
NOR3_X1 U769 ( .A1(n1083), .A2(KEYINPUT18), .A3(G902), .ZN(n1082) );
XOR2_X1 U770 ( .A(n1084), .B(n1085), .Z(G72) );
NOR2_X1 U771 ( .A1(n1086), .A2(n1066), .ZN(n1085) );
NOR2_X1 U772 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U773 ( .A(KEYINPUT60), .B(G227), .Z(n1088) );
NAND2_X1 U774 ( .A1(n1089), .A2(n1090), .ZN(n1084) );
NAND2_X1 U775 ( .A1(n1091), .A2(n1066), .ZN(n1090) );
XOR2_X1 U776 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND3_X1 U777 ( .A1(G900), .A2(n1092), .A3(G953), .ZN(n1089) );
XOR2_X1 U778 ( .A(n1094), .B(n1095), .Z(n1092) );
NOR2_X1 U779 ( .A1(KEYINPUT35), .A2(n1096), .ZN(n1095) );
XOR2_X1 U780 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U781 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
XOR2_X1 U782 ( .A(KEYINPUT30), .B(n1101), .Z(n1100) );
NOR2_X1 U783 ( .A1(G137), .A2(n1102), .ZN(n1101) );
NOR2_X1 U784 ( .A1(G134), .A2(n1103), .ZN(n1099) );
XOR2_X1 U785 ( .A(n1104), .B(n1105), .Z(G69) );
NOR2_X1 U786 ( .A1(n1106), .A2(n1066), .ZN(n1105) );
AND2_X1 U787 ( .A1(G224), .A2(G898), .ZN(n1106) );
NOR2_X1 U788 ( .A1(KEYINPUT13), .A2(n1107), .ZN(n1104) );
XOR2_X1 U789 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U790 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XNOR2_X1 U791 ( .A(G953), .B(KEYINPUT63), .ZN(n1111) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
XOR2_X1 U793 ( .A(KEYINPUT47), .B(n1114), .Z(n1113) );
NAND2_X1 U794 ( .A1(n1115), .A2(n1116), .ZN(n1108) );
NAND2_X1 U795 ( .A1(G953), .A2(n1117), .ZN(n1116) );
XOR2_X1 U796 ( .A(n1118), .B(n1119), .Z(n1115) );
NAND2_X1 U797 ( .A1(KEYINPUT38), .A2(n1120), .ZN(n1118) );
NOR2_X1 U798 ( .A1(n1121), .A2(n1122), .ZN(G66) );
XOR2_X1 U799 ( .A(KEYINPUT43), .B(n1123), .Z(n1122) );
XNOR2_X1 U800 ( .A(n1124), .B(n1083), .ZN(n1121) );
NAND2_X1 U801 ( .A1(n1125), .A2(n1081), .ZN(n1124) );
NOR2_X1 U802 ( .A1(n1123), .A2(n1126), .ZN(G63) );
XOR2_X1 U803 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR3_X1 U804 ( .A1(n1129), .A2(KEYINPUT44), .A3(n1130), .ZN(n1127) );
NOR2_X1 U805 ( .A1(n1123), .A2(n1131), .ZN(G60) );
XOR2_X1 U806 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U807 ( .A1(n1125), .A2(G475), .ZN(n1132) );
XOR2_X1 U808 ( .A(G104), .B(n1114), .Z(G6) );
NOR3_X1 U809 ( .A1(n1123), .A2(n1134), .A3(n1135), .ZN(G57) );
NOR3_X1 U810 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
NOR2_X1 U811 ( .A1(n1139), .A2(n1140), .ZN(n1134) );
NOR2_X1 U812 ( .A1(n1137), .A2(n1138), .ZN(n1140) );
NOR2_X1 U813 ( .A1(n1141), .A2(n1142), .ZN(n1138) );
AND2_X1 U814 ( .A1(n1143), .A2(n1141), .ZN(n1137) );
XNOR2_X1 U815 ( .A(n1144), .B(n1145), .ZN(n1141) );
NAND2_X1 U816 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
XOR2_X1 U817 ( .A(KEYINPUT5), .B(KEYINPUT23), .Z(n1146) );
XNOR2_X1 U818 ( .A(KEYINPUT45), .B(n1142), .ZN(n1143) );
NAND2_X1 U819 ( .A1(n1125), .A2(G472), .ZN(n1142) );
INV_X1 U820 ( .A(n1136), .ZN(n1139) );
NAND2_X1 U821 ( .A1(n1148), .A2(n1149), .ZN(n1136) );
NOR2_X1 U822 ( .A1(n1123), .A2(n1150), .ZN(G54) );
XOR2_X1 U823 ( .A(n1151), .B(n1152), .Z(n1150) );
XNOR2_X1 U824 ( .A(n1153), .B(n1154), .ZN(n1152) );
NAND2_X1 U825 ( .A1(n1125), .A2(G469), .ZN(n1153) );
XOR2_X1 U826 ( .A(n1155), .B(n1156), .Z(n1151) );
XOR2_X1 U827 ( .A(KEYINPUT53), .B(n1157), .Z(n1156) );
NOR2_X1 U828 ( .A1(KEYINPUT4), .A2(n1158), .ZN(n1155) );
XNOR2_X1 U829 ( .A(G110), .B(G140), .ZN(n1158) );
NOR2_X1 U830 ( .A1(n1123), .A2(n1159), .ZN(G51) );
XOR2_X1 U831 ( .A(n1160), .B(n1161), .Z(n1159) );
XNOR2_X1 U832 ( .A(n1162), .B(n1163), .ZN(n1161) );
XOR2_X1 U833 ( .A(n1164), .B(n1165), .Z(n1160) );
XOR2_X1 U834 ( .A(n1166), .B(n1167), .Z(n1165) );
NAND2_X1 U835 ( .A1(KEYINPUT17), .A2(n1168), .ZN(n1167) );
INV_X1 U836 ( .A(G125), .ZN(n1168) );
NAND2_X1 U837 ( .A1(n1125), .A2(n1169), .ZN(n1164) );
INV_X1 U838 ( .A(n1129), .ZN(n1125) );
NAND2_X1 U839 ( .A1(G902), .A2(n1033), .ZN(n1129) );
OR3_X1 U840 ( .A1(n1112), .A2(n1114), .A3(n1093), .ZN(n1033) );
NAND2_X1 U841 ( .A1(n1170), .A2(n1171), .ZN(n1093) );
AND4_X1 U842 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1171) );
NOR4_X1 U843 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1170) );
NOR2_X1 U844 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NOR2_X1 U845 ( .A1(KEYINPUT51), .A2(n1182), .ZN(n1178) );
NOR2_X1 U846 ( .A1(n1183), .A2(n1037), .ZN(n1177) );
NOR2_X1 U847 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR3_X1 U848 ( .A1(n1186), .A2(n1049), .A3(n1187), .ZN(n1184) );
NAND3_X1 U849 ( .A1(n1061), .A2(n1181), .A3(n1057), .ZN(n1186) );
INV_X1 U850 ( .A(KEYINPUT59), .ZN(n1181) );
NOR2_X1 U851 ( .A1(n1188), .A2(n1189), .ZN(n1176) );
NOR2_X1 U852 ( .A1(n1190), .A2(n1191), .ZN(n1188) );
NOR2_X1 U853 ( .A1(n1037), .A2(n1050), .ZN(n1191) );
AND3_X1 U854 ( .A1(KEYINPUT51), .A2(n1062), .A3(n1058), .ZN(n1190) );
NOR3_X1 U855 ( .A1(n1056), .A2(n1192), .A3(n1193), .ZN(n1114) );
NAND4_X1 U856 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1112) );
NOR3_X1 U857 ( .A1(n1198), .A2(n1029), .A3(n1199), .ZN(n1197) );
AND3_X1 U858 ( .A1(n1200), .A2(n1057), .A3(n1201), .ZN(n1029) );
NAND2_X1 U859 ( .A1(n1054), .A2(n1201), .ZN(n1196) );
INV_X1 U860 ( .A(n1192), .ZN(n1201) );
NAND2_X1 U861 ( .A1(n1202), .A2(n1203), .ZN(n1194) );
NAND2_X1 U862 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
XOR2_X1 U863 ( .A(n1206), .B(KEYINPUT22), .Z(n1204) );
NAND4_X1 U864 ( .A1(n1207), .A2(n1208), .A3(n1058), .A4(n1070), .ZN(n1206) );
XOR2_X1 U865 ( .A(n1209), .B(KEYINPUT19), .Z(n1207) );
NOR2_X1 U866 ( .A1(n1066), .A2(G952), .ZN(n1123) );
XNOR2_X1 U867 ( .A(G146), .B(n1182), .ZN(G48) );
NAND3_X1 U868 ( .A1(n1058), .A2(n1202), .A3(n1210), .ZN(n1182) );
XNOR2_X1 U869 ( .A(G143), .B(n1175), .ZN(G45) );
NAND4_X1 U870 ( .A1(n1211), .A2(n1202), .A3(n1077), .A4(n1212), .ZN(n1175) );
XNOR2_X1 U871 ( .A(n1213), .B(n1214), .ZN(G42) );
NOR2_X1 U872 ( .A1(n1037), .A2(n1215), .ZN(n1214) );
XOR2_X1 U873 ( .A(KEYINPUT11), .B(n1185), .Z(n1215) );
AND2_X1 U874 ( .A1(n1216), .A2(n1217), .ZN(n1185) );
XNOR2_X1 U875 ( .A(G137), .B(n1218), .ZN(G39) );
NAND4_X1 U876 ( .A1(n1054), .A2(n1219), .A3(KEYINPUT6), .A4(n1220), .ZN(n1218) );
NOR3_X1 U877 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1220) );
XOR2_X1 U878 ( .A(n1187), .B(KEYINPUT56), .Z(n1223) );
XNOR2_X1 U879 ( .A(G134), .B(n1180), .ZN(G36) );
NAND3_X1 U880 ( .A1(n1211), .A2(n1057), .A3(n1219), .ZN(n1180) );
XOR2_X1 U881 ( .A(n1174), .B(n1224), .Z(G33) );
XNOR2_X1 U882 ( .A(KEYINPUT55), .B(n1225), .ZN(n1224) );
NAND3_X1 U883 ( .A1(n1211), .A2(n1058), .A3(n1219), .ZN(n1174) );
INV_X1 U884 ( .A(n1037), .ZN(n1219) );
NAND2_X1 U885 ( .A1(n1068), .A2(n1226), .ZN(n1037) );
INV_X1 U886 ( .A(n1076), .ZN(n1068) );
AND2_X1 U887 ( .A1(n1208), .A2(n1216), .ZN(n1211) );
XNOR2_X1 U888 ( .A(n1173), .B(n1227), .ZN(G30) );
NOR2_X1 U889 ( .A1(KEYINPUT25), .A2(n1228), .ZN(n1227) );
INV_X1 U890 ( .A(G128), .ZN(n1228) );
NAND3_X1 U891 ( .A1(n1057), .A2(n1202), .A3(n1210), .ZN(n1173) );
INV_X1 U892 ( .A(n1189), .ZN(n1210) );
NAND3_X1 U893 ( .A1(n1056), .A2(n1052), .A3(n1216), .ZN(n1189) );
AND2_X1 U894 ( .A1(n1061), .A2(n1187), .ZN(n1216) );
XNOR2_X1 U895 ( .A(n1229), .B(n1230), .ZN(G3) );
NOR2_X1 U896 ( .A1(n1231), .A2(n1062), .ZN(n1230) );
XOR2_X1 U897 ( .A(n1205), .B(KEYINPUT52), .Z(n1231) );
NAND4_X1 U898 ( .A1(n1232), .A2(n1208), .A3(n1061), .A4(n1209), .ZN(n1205) );
XNOR2_X1 U899 ( .A(G125), .B(n1172), .ZN(G27) );
NAND4_X1 U900 ( .A1(n1217), .A2(n1070), .A3(n1202), .A4(n1187), .ZN(n1172) );
NAND2_X1 U901 ( .A1(n1044), .A2(n1233), .ZN(n1187) );
NAND4_X1 U902 ( .A1(G953), .A2(G902), .A3(n1234), .A4(n1087), .ZN(n1233) );
INV_X1 U903 ( .A(G900), .ZN(n1087) );
NOR3_X1 U904 ( .A1(n1052), .A2(n1200), .A3(n1193), .ZN(n1217) );
XNOR2_X1 U905 ( .A(G122), .B(n1195), .ZN(G24) );
NAND3_X1 U906 ( .A1(n1200), .A2(n1235), .A3(n1236), .ZN(n1195) );
NOR3_X1 U907 ( .A1(n1052), .A2(n1237), .A3(n1238), .ZN(n1236) );
XOR2_X1 U908 ( .A(G119), .B(n1198), .Z(G21) );
NOR3_X1 U909 ( .A1(n1239), .A2(n1222), .A3(n1240), .ZN(n1198) );
NAND2_X1 U910 ( .A1(n1241), .A2(n1242), .ZN(G18) );
NAND2_X1 U911 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
INV_X1 U912 ( .A(G116), .ZN(n1244) );
NAND2_X1 U913 ( .A1(G116), .A2(n1245), .ZN(n1241) );
NAND2_X1 U914 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
NAND2_X1 U915 ( .A1(KEYINPUT62), .A2(n1199), .ZN(n1247) );
INV_X1 U916 ( .A(n1248), .ZN(n1199) );
OR2_X1 U917 ( .A1(n1243), .A2(KEYINPUT62), .ZN(n1246) );
NOR2_X1 U918 ( .A1(KEYINPUT27), .A2(n1248), .ZN(n1243) );
NAND3_X1 U919 ( .A1(n1208), .A2(n1057), .A3(n1235), .ZN(n1248) );
INV_X1 U920 ( .A(n1239), .ZN(n1235) );
NOR2_X1 U921 ( .A1(n1212), .A2(n1238), .ZN(n1057) );
INV_X1 U922 ( .A(n1077), .ZN(n1238) );
XOR2_X1 U923 ( .A(n1249), .B(n1250), .Z(G15) );
NOR3_X1 U924 ( .A1(n1239), .A2(n1193), .A3(n1049), .ZN(n1250) );
INV_X1 U925 ( .A(n1208), .ZN(n1049) );
NOR2_X1 U926 ( .A1(n1056), .A2(n1222), .ZN(n1208) );
INV_X1 U927 ( .A(n1058), .ZN(n1193) );
NOR2_X1 U928 ( .A1(n1077), .A2(n1237), .ZN(n1058) );
INV_X1 U929 ( .A(n1212), .ZN(n1237) );
NAND3_X1 U930 ( .A1(n1202), .A2(n1209), .A3(n1070), .ZN(n1239) );
NOR2_X1 U931 ( .A1(n1043), .A2(n1251), .ZN(n1070) );
INV_X1 U932 ( .A(n1042), .ZN(n1251) );
XNOR2_X1 U933 ( .A(G113), .B(KEYINPUT7), .ZN(n1249) );
XOR2_X1 U934 ( .A(G110), .B(n1252), .Z(G12) );
NOR3_X1 U935 ( .A1(n1240), .A2(KEYINPUT46), .A3(n1192), .ZN(n1252) );
NAND4_X1 U936 ( .A1(n1061), .A2(n1202), .A3(n1222), .A4(n1209), .ZN(n1192) );
NAND2_X1 U937 ( .A1(n1044), .A2(n1253), .ZN(n1209) );
NAND4_X1 U938 ( .A1(G953), .A2(G902), .A3(n1234), .A4(n1117), .ZN(n1253) );
INV_X1 U939 ( .A(G898), .ZN(n1117) );
NAND3_X1 U940 ( .A1(n1234), .A2(n1066), .A3(G952), .ZN(n1044) );
NAND2_X1 U941 ( .A1(G237), .A2(G234), .ZN(n1234) );
INV_X1 U942 ( .A(n1052), .ZN(n1222) );
XNOR2_X1 U943 ( .A(n1254), .B(n1255), .ZN(n1052) );
XOR2_X1 U944 ( .A(KEYINPUT54), .B(G472), .Z(n1255) );
NAND2_X1 U945 ( .A1(n1256), .A2(n1257), .ZN(n1254) );
XOR2_X1 U946 ( .A(n1258), .B(n1259), .Z(n1256) );
NOR2_X1 U947 ( .A1(KEYINPUT61), .A2(n1260), .ZN(n1259) );
XOR2_X1 U948 ( .A(n1147), .B(n1261), .Z(n1260) );
XOR2_X1 U949 ( .A(KEYINPUT0), .B(n1145), .Z(n1261) );
AND3_X1 U950 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1145) );
NAND2_X1 U951 ( .A1(KEYINPUT28), .A2(n1265), .ZN(n1264) );
OR3_X1 U952 ( .A1(n1265), .A2(KEYINPUT28), .A3(n1266), .ZN(n1263) );
NAND2_X1 U953 ( .A1(n1266), .A2(n1267), .ZN(n1262) );
NAND2_X1 U954 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
INV_X1 U955 ( .A(KEYINPUT28), .ZN(n1269) );
XNOR2_X1 U956 ( .A(KEYINPUT9), .B(n1265), .ZN(n1268) );
XOR2_X1 U957 ( .A(n1270), .B(n1271), .Z(n1266) );
XNOR2_X1 U958 ( .A(G116), .B(KEYINPUT49), .ZN(n1270) );
XOR2_X1 U959 ( .A(KEYINPUT40), .B(n1272), .Z(n1147) );
NOR2_X1 U960 ( .A1(n1273), .A2(n1274), .ZN(n1258) );
XOR2_X1 U961 ( .A(n1148), .B(KEYINPUT57), .Z(n1274) );
NAND2_X1 U962 ( .A1(n1229), .A2(n1275), .ZN(n1148) );
NAND2_X1 U963 ( .A1(n1276), .A2(G210), .ZN(n1275) );
INV_X1 U964 ( .A(G101), .ZN(n1229) );
INV_X1 U965 ( .A(n1149), .ZN(n1273) );
NAND3_X1 U966 ( .A1(G210), .A2(G101), .A3(n1276), .ZN(n1149) );
INV_X1 U967 ( .A(n1062), .ZN(n1202) );
NAND2_X1 U968 ( .A1(n1226), .A2(n1076), .ZN(n1062) );
XNOR2_X1 U969 ( .A(n1277), .B(n1169), .ZN(n1076) );
AND2_X1 U970 ( .A1(G210), .A2(n1278), .ZN(n1169) );
NAND2_X1 U971 ( .A1(n1279), .A2(n1257), .ZN(n1277) );
XOR2_X1 U972 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U973 ( .A(G125), .B(n1282), .ZN(n1281) );
XNOR2_X1 U974 ( .A(KEYINPUT29), .B(KEYINPUT20), .ZN(n1282) );
XOR2_X1 U975 ( .A(n1283), .B(n1162), .Z(n1280) );
XOR2_X1 U976 ( .A(KEYINPUT40), .B(n1284), .Z(n1162) );
XNOR2_X1 U977 ( .A(n1285), .B(n1166), .ZN(n1283) );
NAND2_X1 U978 ( .A1(G224), .A2(n1066), .ZN(n1166) );
NAND2_X1 U979 ( .A1(KEYINPUT42), .A2(n1163), .ZN(n1285) );
XOR2_X1 U980 ( .A(n1120), .B(n1119), .Z(n1163) );
XNOR2_X1 U981 ( .A(n1286), .B(G110), .ZN(n1119) );
NAND2_X1 U982 ( .A1(KEYINPUT24), .A2(n1287), .ZN(n1286) );
XOR2_X1 U983 ( .A(n1288), .B(n1289), .Z(n1120) );
XOR2_X1 U984 ( .A(G104), .B(n1290), .Z(n1289) );
XNOR2_X1 U985 ( .A(KEYINPUT8), .B(n1265), .ZN(n1290) );
INV_X1 U986 ( .A(G113), .ZN(n1265) );
XOR2_X1 U987 ( .A(n1291), .B(n1292), .Z(n1288) );
XNOR2_X1 U988 ( .A(G101), .B(n1271), .ZN(n1291) );
XNOR2_X1 U989 ( .A(n1069), .B(KEYINPUT21), .ZN(n1226) );
AND2_X1 U990 ( .A1(G214), .A2(n1278), .ZN(n1069) );
NAND2_X1 U991 ( .A1(n1257), .A2(n1293), .ZN(n1278) );
INV_X1 U992 ( .A(G237), .ZN(n1293) );
INV_X1 U993 ( .A(n1221), .ZN(n1061) );
NAND2_X1 U994 ( .A1(n1294), .A2(n1043), .ZN(n1221) );
XNOR2_X1 U995 ( .A(n1295), .B(G469), .ZN(n1043) );
NAND3_X1 U996 ( .A1(n1296), .A2(n1297), .A3(n1257), .ZN(n1295) );
NAND2_X1 U997 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
INV_X1 U998 ( .A(KEYINPUT39), .ZN(n1299) );
XNOR2_X1 U999 ( .A(n1300), .B(n1301), .ZN(n1298) );
INV_X1 U1000 ( .A(n1154), .ZN(n1301) );
NAND3_X1 U1001 ( .A1(n1154), .A2(n1300), .A3(KEYINPUT39), .ZN(n1296) );
AND2_X1 U1002 ( .A1(n1302), .A2(n1303), .ZN(n1300) );
NAND2_X1 U1003 ( .A1(G140), .A2(n1304), .ZN(n1303) );
NAND2_X1 U1004 ( .A1(n1305), .A2(n1213), .ZN(n1302) );
INV_X1 U1005 ( .A(G140), .ZN(n1213) );
XNOR2_X1 U1006 ( .A(KEYINPUT58), .B(n1304), .ZN(n1305) );
XNOR2_X1 U1007 ( .A(G110), .B(n1157), .ZN(n1304) );
AND2_X1 U1008 ( .A1(G227), .A2(n1066), .ZN(n1157) );
XNOR2_X1 U1009 ( .A(n1306), .B(n1272), .ZN(n1154) );
XOR2_X1 U1010 ( .A(n1098), .B(n1307), .Z(n1272) );
XNOR2_X1 U1011 ( .A(n1102), .B(n1308), .ZN(n1307) );
NOR2_X1 U1012 ( .A1(G137), .A2(KEYINPUT36), .ZN(n1308) );
INV_X1 U1013 ( .A(G134), .ZN(n1102) );
XOR2_X1 U1014 ( .A(G131), .B(n1284), .Z(n1098) );
XNOR2_X1 U1015 ( .A(n1309), .B(n1310), .ZN(n1284) );
XNOR2_X1 U1016 ( .A(G101), .B(n1311), .ZN(n1306) );
NOR2_X1 U1017 ( .A1(KEYINPUT31), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U1018 ( .A(G107), .B(G104), .ZN(n1312) );
XNOR2_X1 U1019 ( .A(KEYINPUT50), .B(n1042), .ZN(n1294) );
NAND2_X1 U1020 ( .A1(G221), .A2(n1313), .ZN(n1042) );
INV_X1 U1021 ( .A(n1054), .ZN(n1240) );
NOR2_X1 U1022 ( .A1(n1050), .A2(n1200), .ZN(n1054) );
INV_X1 U1023 ( .A(n1056), .ZN(n1200) );
XNOR2_X1 U1024 ( .A(n1314), .B(n1081), .ZN(n1056) );
AND2_X1 U1025 ( .A1(G217), .A2(n1313), .ZN(n1081) );
NAND2_X1 U1026 ( .A1(G234), .A2(n1257), .ZN(n1313) );
NAND2_X1 U1027 ( .A1(n1315), .A2(n1257), .ZN(n1314) );
INV_X1 U1028 ( .A(n1083), .ZN(n1315) );
XNOR2_X1 U1029 ( .A(n1316), .B(n1317), .ZN(n1083) );
XOR2_X1 U1030 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1031 ( .A(n1320), .B(n1321), .Z(n1319) );
NAND2_X1 U1032 ( .A1(KEYINPUT12), .A2(n1103), .ZN(n1321) );
INV_X1 U1033 ( .A(G137), .ZN(n1103) );
NAND2_X1 U1034 ( .A1(n1322), .A2(G221), .ZN(n1320) );
XOR2_X1 U1035 ( .A(G146), .B(G110), .Z(n1318) );
XNOR2_X1 U1036 ( .A(n1310), .B(n1323), .ZN(n1316) );
XOR2_X1 U1037 ( .A(n1271), .B(n1094), .Z(n1323) );
XOR2_X1 U1038 ( .A(G119), .B(KEYINPUT15), .Z(n1271) );
INV_X1 U1039 ( .A(n1232), .ZN(n1050) );
NOR2_X1 U1040 ( .A1(n1077), .A2(n1212), .ZN(n1232) );
XNOR2_X1 U1041 ( .A(n1079), .B(G475), .ZN(n1212) );
NAND2_X1 U1042 ( .A1(n1133), .A2(n1257), .ZN(n1079) );
INV_X1 U1043 ( .A(G902), .ZN(n1257) );
XOR2_X1 U1044 ( .A(n1324), .B(n1325), .Z(n1133) );
XOR2_X1 U1045 ( .A(n1326), .B(n1327), .Z(n1325) );
XOR2_X1 U1046 ( .A(G104), .B(n1328), .Z(n1327) );
NOR4_X1 U1047 ( .A1(n1329), .A2(n1330), .A3(KEYINPUT34), .A4(n1331), .ZN(n1328) );
AND2_X1 U1048 ( .A1(G113), .A2(KEYINPUT2), .ZN(n1331) );
NOR2_X1 U1049 ( .A1(n1332), .A2(n1287), .ZN(n1330) );
INV_X1 U1050 ( .A(G122), .ZN(n1287) );
NOR2_X1 U1051 ( .A1(G113), .A2(KEYINPUT33), .ZN(n1332) );
NOR4_X1 U1052 ( .A1(G122), .A2(G113), .A3(KEYINPUT33), .A4(KEYINPUT2), .ZN(n1329) );
AND2_X1 U1053 ( .A1(G214), .A2(n1276), .ZN(n1326) );
NOR2_X1 U1054 ( .A1(G953), .A2(G237), .ZN(n1276) );
XNOR2_X1 U1055 ( .A(n1333), .B(n1309), .ZN(n1324) );
XNOR2_X1 U1056 ( .A(G143), .B(G146), .ZN(n1309) );
XOR2_X1 U1057 ( .A(n1334), .B(n1094), .Z(n1333) );
XOR2_X1 U1058 ( .A(G125), .B(G140), .Z(n1094) );
NAND2_X1 U1059 ( .A1(KEYINPUT3), .A2(n1225), .ZN(n1334) );
INV_X1 U1060 ( .A(G131), .ZN(n1225) );
XOR2_X1 U1061 ( .A(n1335), .B(n1130), .Z(n1077) );
INV_X1 U1062 ( .A(G478), .ZN(n1130) );
OR2_X1 U1063 ( .A1(n1128), .A2(G902), .ZN(n1335) );
XNOR2_X1 U1064 ( .A(n1336), .B(n1337), .ZN(n1128) );
XNOR2_X1 U1065 ( .A(n1310), .B(n1338), .ZN(n1337) );
XOR2_X1 U1066 ( .A(n1339), .B(n1340), .Z(n1338) );
NOR2_X1 U1067 ( .A1(KEYINPUT14), .A2(n1341), .ZN(n1340) );
XNOR2_X1 U1068 ( .A(G122), .B(n1292), .ZN(n1341) );
XNOR2_X1 U1069 ( .A(n1342), .B(G116), .ZN(n1292) );
INV_X1 U1070 ( .A(G107), .ZN(n1342) );
NAND2_X1 U1071 ( .A1(G217), .A2(n1322), .ZN(n1339) );
AND2_X1 U1072 ( .A1(G234), .A2(n1066), .ZN(n1322) );
INV_X1 U1073 ( .A(G953), .ZN(n1066) );
XOR2_X1 U1074 ( .A(G128), .B(KEYINPUT48), .Z(n1310) );
XNOR2_X1 U1075 ( .A(G134), .B(n1343), .ZN(n1336) );
XOR2_X1 U1076 ( .A(KEYINPUT26), .B(G143), .Z(n1343) );
endmodule


