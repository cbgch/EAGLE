//Key = 0010010000110001000010010100011011111110100100011111000100101101


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229;

OR2_X1 U1253 ( .A1(n2229), .A2(n1683), .ZN(U280) );
OR2_X1 U1254 ( .A1(n1825), .A2(STATO_REG_0__SCAN_IN), .ZN(n1682) );
INV_X2 U1255 ( .A(n1682), .ZN(n1683) );
INV_X2 U1256 ( .A(U280), .ZN(n1684) );
NOR4_X2 U1257 ( .A1(n1824), .A2(n2152), .A3(n2150), .A4(AVERAGE), .ZN(n1932));
INV_X1 U1258 ( .A(n1685), .ZN(U375) );
NAND2_X1 U1259 ( .A1(n1686), .A2(n1687), .ZN(U344) );
NAND2_X1 U1260 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1688), .ZN(n1687) );
NAND2_X1 U1261 ( .A1(n1689), .A2(DATA_IN_7_), .ZN(n1686) );
NAND2_X1 U1262 ( .A1(n1690), .A2(n1691), .ZN(U343) );
NAND2_X1 U1263 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1688), .ZN(n1691) );
NAND2_X1 U1264 ( .A1(n1689), .A2(DATA_IN_6_), .ZN(n1690) );
NAND2_X1 U1265 ( .A1(n1692), .A2(n1693), .ZN(U342) );
NAND2_X1 U1266 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1688), .ZN(n1693) );
NAND2_X1 U1267 ( .A1(n1689), .A2(DATA_IN_5_), .ZN(n1692) );
NAND2_X1 U1268 ( .A1(n1694), .A2(n1695), .ZN(U341) );
NAND2_X1 U1269 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1688), .ZN(n1695) );
NAND2_X1 U1270 ( .A1(n1689), .A2(DATA_IN_4_), .ZN(n1694) );
NAND2_X1 U1271 ( .A1(n1696), .A2(n1697), .ZN(U340) );
NAND2_X1 U1272 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1688), .ZN(n1697) );
NAND2_X1 U1273 ( .A1(n1689), .A2(DATA_IN_3_), .ZN(n1696) );
NAND2_X1 U1274 ( .A1(n1698), .A2(n1699), .ZN(U339) );
NAND2_X1 U1275 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1688), .ZN(n1699) );
NAND2_X1 U1276 ( .A1(n1689), .A2(DATA_IN_2_), .ZN(n1698) );
NAND2_X1 U1277 ( .A1(n1700), .A2(n1701), .ZN(U338) );
NAND2_X1 U1278 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1688), .ZN(n1701) );
NAND2_X1 U1279 ( .A1(n1689), .A2(DATA_IN_1_), .ZN(n1700) );
NAND2_X1 U1280 ( .A1(n1702), .A2(n1703), .ZN(U337) );
NAND2_X1 U1281 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1688), .ZN(n1703) );
NAND2_X1 U1282 ( .A1(n1689), .A2(DATA_IN_0_), .ZN(n1702) );
INV_X1 U1283 ( .A(n1688), .ZN(n1689) );
NAND2_X1 U1284 ( .A1(n1685), .A2(n1704), .ZN(n1688) );
NAND3_X1 U1285 ( .A1(n1705), .A2(n1706), .A3(n1707), .ZN(n1704) );
NAND2_X1 U1286 ( .A1(n1708), .A2(n1709), .ZN(U336) );
NAND2_X1 U1287 ( .A1(n1710), .A2(DATA_IN_7_), .ZN(n1709) );
XOR2_X1 U1288 ( .A(n1711), .B(KEYINPUT23), .Z(n1710) );
NAND2_X1 U1289 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1711), .ZN(n1708) );
NAND2_X1 U1290 ( .A1(n1712), .A2(n1713), .ZN(U335) );
NAND2_X1 U1291 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1711), .ZN(n1713) );
NAND2_X1 U1292 ( .A1(n1714), .A2(DATA_IN_6_), .ZN(n1712) );
NAND2_X1 U1293 ( .A1(n1715), .A2(n1716), .ZN(U334) );
NAND2_X1 U1294 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1711), .ZN(n1716) );
NAND2_X1 U1295 ( .A1(n1714), .A2(DATA_IN_5_), .ZN(n1715) );
NAND2_X1 U1296 ( .A1(n1717), .A2(n1718), .ZN(U333) );
NAND2_X1 U1297 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1711), .ZN(n1718) );
NAND2_X1 U1298 ( .A1(n1714), .A2(DATA_IN_4_), .ZN(n1717) );
NAND2_X1 U1299 ( .A1(n1719), .A2(n1720), .ZN(U332) );
NAND2_X1 U1300 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1711), .ZN(n1720) );
NAND2_X1 U1301 ( .A1(n1714), .A2(DATA_IN_3_), .ZN(n1719) );
NAND2_X1 U1302 ( .A1(n1721), .A2(n1722), .ZN(U331) );
NAND2_X1 U1303 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1711), .ZN(n1722) );
NAND2_X1 U1304 ( .A1(n1714), .A2(DATA_IN_2_), .ZN(n1721) );
NAND2_X1 U1305 ( .A1(n1723), .A2(n1724), .ZN(U330) );
NAND2_X1 U1306 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1711), .ZN(n1724) );
NAND2_X1 U1307 ( .A1(n1714), .A2(DATA_IN_1_), .ZN(n1723) );
NAND2_X1 U1308 ( .A1(n1725), .A2(n1726), .ZN(U329) );
NAND2_X1 U1309 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1711), .ZN(n1726) );
NAND2_X1 U1310 ( .A1(n1714), .A2(n1727), .ZN(n1725) );
XOR2_X1 U1311 ( .A(n1728), .B(KEYINPUT15), .Z(n1727) );
INV_X1 U1312 ( .A(n1711), .ZN(n1714) );
NAND2_X1 U1313 ( .A1(n1685), .A2(n1729), .ZN(n1711) );
NAND2_X1 U1314 ( .A1(n1730), .A2(n1706), .ZN(n1729) );
NAND3_X1 U1315 ( .A1(n1707), .A2(n1705), .A3(n1731), .ZN(n1730) );
NAND2_X1 U1316 ( .A1(n1732), .A2(n1733), .ZN(n1731) );
NAND3_X1 U1317 ( .A1(n1734), .A2(n1735), .A3(n1736), .ZN(n1733) );
NAND2_X1 U1318 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1737), .ZN(n1736) );
NAND3_X1 U1319 ( .A1(n1738), .A2(n1739), .A3(n1740), .ZN(n1735) );
XOR2_X1 U1320 ( .A(n1741), .B(KEYINPUT53), .Z(n1740) );
NAND3_X1 U1321 ( .A1(n1742), .A2(n1743), .A3(n1744), .ZN(n1741) );
XOR2_X1 U1322 ( .A(n1745), .B(KEYINPUT12), .Z(n1744) );
NAND2_X1 U1323 ( .A1(DATA_IN_4_), .A2(n1746), .ZN(n1745) );
NAND3_X1 U1324 ( .A1(n1747), .A2(n1748), .A3(n1749), .ZN(n1743) );
NAND2_X1 U1325 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1750), .ZN(n1749) );
NAND3_X1 U1326 ( .A1(n1751), .A2(n1752), .A3(n1753), .ZN(n1748) );
NAND2_X1 U1327 ( .A1(DATA_IN_3_), .A2(n1754), .ZN(n1753) );
NAND3_X1 U1328 ( .A1(n1755), .A2(n1756), .A3(n1757), .ZN(n1752) );
NAND2_X1 U1329 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1758), .ZN(n1757) );
NAND3_X1 U1330 ( .A1(n1759), .A2(n1728), .A3(n1760), .ZN(n1756) );
XNOR2_X1 U1331 ( .A(RMIN_REG_0__SCAN_IN), .B(KEYINPUT5), .ZN(n1760) );
NAND2_X1 U1332 ( .A1(DATA_IN_1_), .A2(n1761), .ZN(n1759) );
NAND2_X1 U1333 ( .A1(n1762), .A2(RMIN_REG_1__SCAN_IN), .ZN(n1755) );
XOR2_X1 U1334 ( .A(n1763), .B(KEYINPUT41), .Z(n1762) );
NAND2_X1 U1335 ( .A1(DATA_IN_2_), .A2(n1764), .ZN(n1751) );
NAND2_X1 U1336 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1765), .ZN(n1747) );
NAND2_X1 U1337 ( .A1(DATA_IN_5_), .A2(n1766), .ZN(n1742) );
NAND2_X1 U1338 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1767), .ZN(n1739) );
NAND2_X1 U1339 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1768), .ZN(n1738) );
NAND2_X1 U1340 ( .A1(DATA_IN_6_), .A2(n1769), .ZN(n1734) );
NAND2_X1 U1341 ( .A1(n1770), .A2(DATA_IN_7_), .ZN(n1732) );
XOR2_X1 U1342 ( .A(n1771), .B(KEYINPUT7), .Z(n1770) );
NAND3_X1 U1343 ( .A1(n1772), .A2(n1773), .A3(n1774), .ZN(n1705) );
OR2_X1 U1344 ( .A1(n1737), .A2(RMAX_REG_7__SCAN_IN), .ZN(n1774) );
NAND3_X1 U1345 ( .A1(n1775), .A2(n1776), .A3(n1777), .ZN(n1773) );
NAND2_X1 U1346 ( .A1(DATA_IN_6_), .A2(n1778), .ZN(n1777) );
NAND3_X1 U1347 ( .A1(n1779), .A2(n1780), .A3(n1781), .ZN(n1776) );
NAND2_X1 U1348 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1767), .ZN(n1781) );
INV_X1 U1349 ( .A(DATA_IN_5_), .ZN(n1767) );
NAND3_X1 U1350 ( .A1(n1782), .A2(n1783), .A3(n1784), .ZN(n1780) );
NAND2_X1 U1351 ( .A1(DATA_IN_4_), .A2(n1785), .ZN(n1784) );
NAND3_X1 U1352 ( .A1(n1786), .A2(n1787), .A3(n1788), .ZN(n1783) );
NAND2_X1 U1353 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1765), .ZN(n1788) );
NAND3_X1 U1354 ( .A1(n1789), .A2(n1790), .A3(n1791), .ZN(n1787) );
NAND2_X1 U1355 ( .A1(DATA_IN_2_), .A2(n1792), .ZN(n1791) );
NAND3_X1 U1356 ( .A1(n1793), .A2(n1794), .A3(DATA_IN_0_), .ZN(n1790) );
NAND2_X1 U1357 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1763), .ZN(n1794) );
XOR2_X1 U1358 ( .A(RMAX_REG_0__SCAN_IN), .B(KEYINPUT47), .Z(n1793) );
NAND2_X1 U1359 ( .A1(n1795), .A2(n1796), .ZN(n1789) );
XOR2_X1 U1360 ( .A(KEYINPUT17), .B(DATA_IN_1_), .Z(n1795) );
NAND2_X1 U1361 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1758), .ZN(n1786) );
NAND2_X1 U1362 ( .A1(DATA_IN_3_), .A2(n1797), .ZN(n1782) );
NAND2_X1 U1363 ( .A1(n1798), .A2(RMAX_REG_4__SCAN_IN), .ZN(n1779) );
XOR2_X1 U1364 ( .A(n1799), .B(DATA_IN_4_), .Z(n1798) );
XNOR2_X1 U1365 ( .A(KEYINPUT57), .B(KEYINPUT22), .ZN(n1799) );
NAND2_X1 U1366 ( .A1(DATA_IN_5_), .A2(n1800), .ZN(n1775) );
NAND2_X1 U1367 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1768), .ZN(n1772) );
INV_X1 U1368 ( .A(DATA_IN_6_), .ZN(n1768) );
NAND2_X1 U1369 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1737), .ZN(n1707) );
NAND2_X1 U1370 ( .A1(n1801), .A2(n1802), .ZN(U328) );
NAND2_X1 U1371 ( .A1(n1803), .A2(DATA_IN_7_), .ZN(n1802) );
NAND2_X1 U1372 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1804), .ZN(n1801) );
NAND2_X1 U1373 ( .A1(n1805), .A2(n1806), .ZN(U327) );
NAND2_X1 U1374 ( .A1(n1807), .A2(n1804), .ZN(n1806) );
XNOR2_X1 U1375 ( .A(RLAST_REG_6__SCAN_IN), .B(KEYINPUT61), .ZN(n1807) );
NAND2_X1 U1376 ( .A1(n1803), .A2(DATA_IN_6_), .ZN(n1805) );
NAND2_X1 U1377 ( .A1(n1808), .A2(n1809), .ZN(U326) );
NAND2_X1 U1378 ( .A1(n1803), .A2(DATA_IN_5_), .ZN(n1809) );
XOR2_X1 U1379 ( .A(n1810), .B(KEYINPUT39), .Z(n1808) );
NAND2_X1 U1380 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1804), .ZN(n1810) );
NAND2_X1 U1381 ( .A1(n1811), .A2(n1812), .ZN(U325) );
NAND2_X1 U1382 ( .A1(n1803), .A2(DATA_IN_4_), .ZN(n1812) );
NAND2_X1 U1383 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1804), .ZN(n1811) );
NAND2_X1 U1384 ( .A1(n1813), .A2(n1814), .ZN(U324) );
NAND2_X1 U1385 ( .A1(n1803), .A2(DATA_IN_3_), .ZN(n1814) );
NAND2_X1 U1386 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1804), .ZN(n1813) );
NAND2_X1 U1387 ( .A1(n1815), .A2(n1816), .ZN(U323) );
NAND2_X1 U1388 ( .A1(n1817), .A2(n1804), .ZN(n1816) );
XOR2_X1 U1389 ( .A(RLAST_REG_2__SCAN_IN), .B(KEYINPUT59), .Z(n1817) );
NAND2_X1 U1390 ( .A1(n1803), .A2(DATA_IN_2_), .ZN(n1815) );
NAND2_X1 U1391 ( .A1(n1818), .A2(n1819), .ZN(U322) );
NAND2_X1 U1392 ( .A1(n1820), .A2(n1804), .ZN(n1819) );
XNOR2_X1 U1393 ( .A(RLAST_REG_1__SCAN_IN), .B(KEYINPUT35), .ZN(n1820) );
NAND2_X1 U1394 ( .A1(n1803), .A2(DATA_IN_1_), .ZN(n1818) );
NAND2_X1 U1395 ( .A1(n1821), .A2(n1822), .ZN(U321) );
NAND2_X1 U1396 ( .A1(n1803), .A2(DATA_IN_0_), .ZN(n1822) );
AND2_X1 U1397 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1823), .ZN(n1803) );
NAND2_X1 U1398 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1804), .ZN(n1821) );
NAND2_X1 U1399 ( .A1(n1685), .A2(n1823), .ZN(n1804) );
NAND2_X1 U1400 ( .A1(n1706), .A2(n1824), .ZN(n1823) );
NAND2_X1 U1401 ( .A1(n1706), .A2(n1825), .ZN(n1685) );
NAND2_X1 U1402 ( .A1(n1826), .A2(n1827), .ZN(U320) );
NAND2_X1 U1403 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1684), .ZN(n1827) );
NAND2_X1 U1404 ( .A1(n1683), .A2(DATA_IN_7_), .ZN(n1826) );
NAND2_X1 U1405 ( .A1(n1828), .A2(n1829), .ZN(U319) );
NAND2_X1 U1406 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1684), .ZN(n1829) );
NAND2_X1 U1407 ( .A1(n1683), .A2(DATA_IN_6_), .ZN(n1828) );
NAND2_X1 U1408 ( .A1(n1830), .A2(n1831), .ZN(U318) );
NAND2_X1 U1409 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1684), .ZN(n1831) );
NAND2_X1 U1410 ( .A1(n1683), .A2(DATA_IN_5_), .ZN(n1830) );
NAND2_X1 U1411 ( .A1(n1832), .A2(n1833), .ZN(U317) );
NAND2_X1 U1412 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1684), .ZN(n1833) );
NAND2_X1 U1413 ( .A1(n1683), .A2(DATA_IN_4_), .ZN(n1832) );
NAND2_X1 U1414 ( .A1(n1834), .A2(n1835), .ZN(U316) );
NAND2_X1 U1415 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1684), .ZN(n1835) );
NAND2_X1 U1416 ( .A1(n1683), .A2(DATA_IN_3_), .ZN(n1834) );
NAND2_X1 U1417 ( .A1(n1836), .A2(n1837), .ZN(U315) );
NAND2_X1 U1418 ( .A1(n1838), .A2(n1683), .ZN(n1837) );
XOR2_X1 U1419 ( .A(n1758), .B(KEYINPUT25), .Z(n1838) );
NAND2_X1 U1420 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1684), .ZN(n1836) );
NAND2_X1 U1421 ( .A1(n1839), .A2(n1840), .ZN(U314) );
NAND2_X1 U1422 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1684), .ZN(n1840) );
NAND2_X1 U1423 ( .A1(n1683), .A2(DATA_IN_1_), .ZN(n1839) );
NAND2_X1 U1424 ( .A1(n1841), .A2(n1842), .ZN(U313) );
NAND2_X1 U1425 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1684), .ZN(n1842) );
NAND2_X1 U1426 ( .A1(n1683), .A2(DATA_IN_0_), .ZN(n1841) );
NAND2_X1 U1427 ( .A1(n1843), .A2(n1844), .ZN(U312) );
NAND2_X1 U1428 ( .A1(n1683), .A2(n1845), .ZN(n1844) );
XOR2_X1 U1429 ( .A(REG1_REG_7__SCAN_IN), .B(KEYINPUT18), .Z(n1845) );
NAND2_X1 U1430 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1684), .ZN(n1843) );
NAND2_X1 U1431 ( .A1(n1846), .A2(n1847), .ZN(U311) );
NAND2_X1 U1432 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1684), .ZN(n1847) );
NAND2_X1 U1433 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1683), .ZN(n1846) );
NAND2_X1 U1434 ( .A1(n1848), .A2(n1849), .ZN(U310) );
NAND2_X1 U1435 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1684), .ZN(n1849) );
XOR2_X1 U1436 ( .A(KEYINPUT2), .B(n1850), .Z(n1848) );
AND2_X1 U1437 ( .A1(n1683), .A2(REG1_REG_5__SCAN_IN), .ZN(n1850) );
NAND2_X1 U1438 ( .A1(n1851), .A2(n1852), .ZN(U309) );
NAND2_X1 U1439 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1684), .ZN(n1852) );
NAND2_X1 U1440 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1683), .ZN(n1851) );
NAND2_X1 U1441 ( .A1(n1853), .A2(n1854), .ZN(U308) );
NAND2_X1 U1442 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1684), .ZN(n1854) );
NAND2_X1 U1443 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1683), .ZN(n1853) );
NAND2_X1 U1444 ( .A1(n1855), .A2(n1856), .ZN(U307) );
NAND2_X1 U1445 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1684), .ZN(n1856) );
NAND2_X1 U1446 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1683), .ZN(n1855) );
NAND2_X1 U1447 ( .A1(n1857), .A2(n1858), .ZN(U306) );
NAND2_X1 U1448 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1684), .ZN(n1858) );
NAND2_X1 U1449 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1683), .ZN(n1857) );
NAND2_X1 U1450 ( .A1(n1859), .A2(n1860), .ZN(U305) );
NAND2_X1 U1451 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1684), .ZN(n1860) );
NAND2_X1 U1452 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1683), .ZN(n1859) );
NAND2_X1 U1453 ( .A1(n1861), .A2(n1862), .ZN(U304) );
NAND2_X1 U1454 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1684), .ZN(n1862) );
NAND2_X1 U1455 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1683), .ZN(n1861) );
NAND2_X1 U1456 ( .A1(n1863), .A2(n1864), .ZN(U303) );
NAND2_X1 U1457 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1683), .ZN(n1864) );
XOR2_X1 U1458 ( .A(n1865), .B(KEYINPUT46), .Z(n1863) );
NAND2_X1 U1459 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1684), .ZN(n1865) );
NAND2_X1 U1460 ( .A1(n1866), .A2(n1867), .ZN(U302) );
NAND2_X1 U1461 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1684), .ZN(n1867) );
NAND2_X1 U1462 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1683), .ZN(n1866) );
NAND2_X1 U1463 ( .A1(n1868), .A2(n1869), .ZN(U301) );
NAND2_X1 U1464 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1684), .ZN(n1869) );
NAND2_X1 U1465 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1683), .ZN(n1868) );
NAND2_X1 U1466 ( .A1(n1870), .A2(n1871), .ZN(U300) );
NAND2_X1 U1467 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1684), .ZN(n1871) );
NAND2_X1 U1468 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1683), .ZN(n1870) );
NAND2_X1 U1469 ( .A1(n1872), .A2(n1873), .ZN(U299) );
NAND2_X1 U1470 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1874), .ZN(n1873) );
XOR2_X1 U1471 ( .A(KEYINPUT0), .B(n1684), .Z(n1874) );
NAND2_X1 U1472 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1683), .ZN(n1872) );
NAND2_X1 U1473 ( .A1(n1875), .A2(n1876), .ZN(U298) );
NAND2_X1 U1474 ( .A1(n1877), .A2(n1683), .ZN(n1876) );
XNOR2_X1 U1475 ( .A(REG2_REG_1__SCAN_IN), .B(KEYINPUT60), .ZN(n1877) );
XOR2_X1 U1476 ( .A(KEYINPUT36), .B(n1878), .Z(n1875) );
NOR2_X1 U1477 ( .A1(n1879), .A2(n1880), .ZN(n1878) );
INV_X1 U1478 ( .A(REG3_REG_1__SCAN_IN), .ZN(n1880) );
XOR2_X1 U1479 ( .A(U280), .B(KEYINPUT4), .Z(n1879) );
NAND2_X1 U1480 ( .A1(n1881), .A2(n1882), .ZN(U297) );
NAND2_X1 U1481 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1684), .ZN(n1882) );
NAND2_X1 U1482 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1683), .ZN(n1881) );
NAND2_X1 U1483 ( .A1(n1883), .A2(n1884), .ZN(U296) );
NAND2_X1 U1484 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1684), .ZN(n1884) );
NAND2_X1 U1485 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1683), .ZN(n1883) );
NAND2_X1 U1486 ( .A1(n1885), .A2(n1886), .ZN(U295) );
NAND2_X1 U1487 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1684), .ZN(n1886) );
NAND2_X1 U1488 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1683), .ZN(n1885) );
NAND2_X1 U1489 ( .A1(n1887), .A2(n1888), .ZN(U294) );
NAND2_X1 U1490 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1684), .ZN(n1888) );
NAND2_X1 U1491 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1683), .ZN(n1887) );
NAND2_X1 U1492 ( .A1(n1889), .A2(n1890), .ZN(U293) );
NAND2_X1 U1493 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1684), .ZN(n1890) );
NAND2_X1 U1494 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1683), .ZN(n1889) );
NAND2_X1 U1495 ( .A1(n1891), .A2(n1892), .ZN(U292) );
NAND2_X1 U1496 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1684), .ZN(n1892) );
NAND2_X1 U1497 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1683), .ZN(n1891) );
NAND2_X1 U1498 ( .A1(n1893), .A2(n1894), .ZN(U291) );
NAND2_X1 U1499 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1683), .ZN(n1894) );
XOR2_X1 U1500 ( .A(n1895), .B(KEYINPUT19), .Z(n1893) );
NAND2_X1 U1501 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1684), .ZN(n1895) );
NAND2_X1 U1502 ( .A1(n1896), .A2(n1897), .ZN(U290) );
NAND2_X1 U1503 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1684), .ZN(n1897) );
NAND2_X1 U1504 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1683), .ZN(n1896) );
NAND2_X1 U1505 ( .A1(n1898), .A2(n1899), .ZN(U289) );
NAND2_X1 U1506 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1684), .ZN(n1899) );
NAND2_X1 U1507 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1683), .ZN(n1898) );
NAND4_X1 U1508 ( .A1(n1900), .A2(n1901), .A3(n1902), .A4(n1903), .ZN(U288));
NAND2_X1 U1509 ( .A1(n1904), .A2(n1905), .ZN(n1903) );
XNOR2_X1 U1510 ( .A(RLAST_REG_7__SCAN_IN), .B(KEYINPUT40), .ZN(n1904) );
NOR2_X1 U1511 ( .A1(n1906), .A2(n1907), .ZN(n1902) );
NOR3_X1 U1512 ( .A1(n1908), .A2(n1909), .A3(n1910), .ZN(n1907) );
XOR2_X1 U1513 ( .A(n1911), .B(KEYINPUT28), .Z(n1910) );
NAND2_X1 U1514 ( .A1(n1912), .A2(REG4_REG_7__SCAN_IN), .ZN(n1901) );
NAND2_X1 U1515 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1684), .ZN(n1900) );
NAND4_X1 U1516 ( .A1(n1913), .A2(n1914), .A3(n1915), .A4(n1916), .ZN(U287));
NOR3_X1 U1517 ( .A1(n1917), .A2(n1918), .A3(n1919), .ZN(n1916) );
AND2_X1 U1518 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1905), .ZN(n1919) );
NOR2_X1 U1519 ( .A1(n1920), .A2(n1911), .ZN(n1918) );
NOR2_X1 U1520 ( .A1(n1921), .A2(n1922), .ZN(n1920) );
XOR2_X1 U1521 ( .A(n1923), .B(KEYINPUT58), .Z(n1922) );
NAND2_X1 U1522 ( .A1(n1924), .A2(n1909), .ZN(n1923) );
XOR2_X1 U1523 ( .A(n1908), .B(KEYINPUT24), .Z(n1924) );
NOR2_X1 U1524 ( .A1(n1909), .A2(n1908), .ZN(n1921) );
XOR2_X1 U1525 ( .A(KEYINPUT62), .B(n1925), .Z(n1917) );
NOR2_X1 U1526 ( .A1(n1926), .A2(n1927), .ZN(n1925) );
NAND2_X1 U1527 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1928), .ZN(n1915) );
XOR2_X1 U1528 ( .A(KEYINPUT54), .B(n1684), .Z(n1928) );
INV_X1 U1529 ( .A(n1906), .ZN(n1914) );
NOR3_X1 U1530 ( .A1(n1929), .A2(n1930), .A3(n1931), .ZN(n1906) );
NAND3_X1 U1531 ( .A1(n1932), .A2(n1929), .A3(n1930), .ZN(n1913) );
NAND4_X1 U1532 ( .A1(n1933), .A2(n1934), .A3(n1935), .A4(n1936), .ZN(U286));
NOR3_X1 U1533 ( .A1(n1937), .A2(n1938), .A3(n1939), .ZN(n1936) );
NOR3_X1 U1534 ( .A1(n1940), .A2(n1930), .A3(n1931), .ZN(n1939) );
AND2_X1 U1535 ( .A1(n1941), .A2(n1942), .ZN(n1930) );
NAND2_X1 U1536 ( .A1(n1929), .A2(n1943), .ZN(n1942) );
NAND2_X1 U1537 ( .A1(n1944), .A2(n1945), .ZN(n1943) );
NAND2_X1 U1538 ( .A1(n1946), .A2(n1947), .ZN(n1929) );
XOR2_X1 U1539 ( .A(KEYINPUT29), .B(n1945), .Z(n1946) );
XOR2_X1 U1540 ( .A(KEYINPUT13), .B(n1948), .Z(n1940) );
NOR2_X1 U1541 ( .A1(n1941), .A2(n1949), .ZN(n1948) );
XOR2_X1 U1542 ( .A(n1950), .B(n1951), .Z(n1949) );
NAND2_X1 U1543 ( .A1(KEYINPUT29), .A2(n1947), .ZN(n1950) );
INV_X1 U1544 ( .A(n1952), .ZN(n1941) );
NOR3_X1 U1545 ( .A1(n1911), .A2(n1909), .A3(n1953), .ZN(n1938) );
NOR2_X1 U1546 ( .A1(n1954), .A2(n1955), .ZN(n1953) );
AND2_X1 U1547 ( .A1(n1954), .A2(n1955), .ZN(n1909) );
NAND2_X1 U1548 ( .A1(n1908), .A2(n1956), .ZN(n1955) );
NAND2_X1 U1549 ( .A1(n1944), .A2(n1957), .ZN(n1956) );
INV_X1 U1550 ( .A(n1947), .ZN(n1944) );
NAND2_X1 U1551 ( .A1(n1958), .A2(n1947), .ZN(n1908) );
INV_X1 U1552 ( .A(n1959), .ZN(n1954) );
NOR2_X1 U1553 ( .A1(n1947), .A2(n1960), .ZN(n1937) );
NAND2_X1 U1554 ( .A1(n1961), .A2(n1962), .ZN(n1947) );
NAND3_X1 U1555 ( .A1(n1963), .A2(n1964), .A3(n1965), .ZN(n1962) );
XOR2_X1 U1556 ( .A(n1966), .B(n1967), .Z(n1965) );
NAND2_X1 U1557 ( .A1(n1968), .A2(n1969), .ZN(n1963) );
NAND3_X1 U1558 ( .A1(n1970), .A2(n1969), .A3(n1971), .ZN(n1961) );
XOR2_X1 U1559 ( .A(n1972), .B(n1967), .Z(n1971) );
AND2_X1 U1560 ( .A1(n1973), .A2(n1974), .ZN(n1967) );
NAND2_X1 U1561 ( .A1(RESTART), .A2(n1769), .ZN(n1974) );
NAND2_X1 U1562 ( .A1(n1926), .A2(n1975), .ZN(n1973) );
NOR2_X1 U1563 ( .A1(KEYINPUT16), .A2(n1966), .ZN(n1972) );
NAND2_X1 U1564 ( .A1(n1976), .A2(n1977), .ZN(n1966) );
NAND2_X1 U1565 ( .A1(DATA_IN_6_), .A2(n1975), .ZN(n1977) );
NAND2_X1 U1566 ( .A1(RESTART), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1976) );
XOR2_X1 U1567 ( .A(KEYINPUT43), .B(n1978), .Z(n1970) );
NOR2_X1 U1568 ( .A1(n1979), .A2(n1968), .ZN(n1978) );
NAND2_X1 U1569 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1684), .ZN(n1935) );
NAND2_X1 U1570 ( .A1(n1905), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1934) );
NAND2_X1 U1571 ( .A1(n1912), .A2(REG4_REG_5__SCAN_IN), .ZN(n1933) );
NAND3_X1 U1572 ( .A1(n1980), .A2(n1981), .A3(n1982), .ZN(U285) );
XNOR2_X1 U1573 ( .A(n1983), .B(KEYINPUT44), .ZN(n1982) );
NAND4_X1 U1574 ( .A1(n1984), .A2(n1985), .A3(n1986), .A4(n1987), .ZN(n1983));
NAND2_X1 U1575 ( .A1(n1988), .A2(REG4_REG_4__SCAN_IN), .ZN(n1987) );
XOR2_X1 U1576 ( .A(n1927), .B(KEYINPUT11), .Z(n1988) );
NAND2_X1 U1577 ( .A1(n1989), .A2(n1990), .ZN(n1986) );
NAND2_X1 U1578 ( .A1(n1905), .A2(RLAST_REG_4__SCAN_IN), .ZN(n1985) );
NAND2_X1 U1579 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1684), .ZN(n1984) );
NAND3_X1 U1580 ( .A1(n1991), .A2(n1952), .A3(n1932), .ZN(n1981) );
NAND3_X1 U1581 ( .A1(n1992), .A2(n1993), .A3(n1994), .ZN(n1952) );
NAND2_X1 U1582 ( .A1(n1995), .A2(n1945), .ZN(n1992) );
NAND3_X1 U1583 ( .A1(n1996), .A2(n1945), .A3(n1995), .ZN(n1991) );
NAND2_X1 U1584 ( .A1(n1990), .A2(n1997), .ZN(n1995) );
INV_X1 U1585 ( .A(n1951), .ZN(n1945) );
NOR2_X1 U1586 ( .A1(n1997), .A2(n1990), .ZN(n1951) );
NAND2_X1 U1587 ( .A1(n1994), .A2(n1998), .ZN(n1996) );
XNOR2_X1 U1588 ( .A(KEYINPUT34), .B(n1993), .ZN(n1998) );
NAND3_X1 U1589 ( .A1(n1999), .A2(n1959), .A3(n2000), .ZN(n1980) );
NAND2_X1 U1590 ( .A1(n2001), .A2(n2002), .ZN(n1959) );
NAND2_X1 U1591 ( .A1(n2003), .A2(n1957), .ZN(n2002) );
NAND3_X1 U1592 ( .A1(n2004), .A2(n1957), .A3(n2003), .ZN(n1999) );
XOR2_X1 U1593 ( .A(n2005), .B(KEYINPUT3), .Z(n2003) );
NAND2_X1 U1594 ( .A1(n1990), .A2(n2006), .ZN(n2005) );
INV_X1 U1595 ( .A(n1958), .ZN(n1957) );
NOR2_X1 U1596 ( .A1(n2006), .A2(n1990), .ZN(n1958) );
NAND2_X1 U1597 ( .A1(n2007), .A2(n2008), .ZN(n1990) );
NAND2_X1 U1598 ( .A1(n2009), .A2(n2010), .ZN(n2008) );
NAND2_X1 U1599 ( .A1(n1964), .A2(n1969), .ZN(n2009) );
NAND2_X1 U1600 ( .A1(n2011), .A2(n2012), .ZN(n1969) );
INV_X1 U1601 ( .A(n1979), .ZN(n1964) );
NOR2_X1 U1602 ( .A1(n2012), .A2(n2011), .ZN(n1979) );
NAND2_X1 U1603 ( .A1(n2013), .A2(n1968), .ZN(n2007) );
INV_X1 U1604 ( .A(n2010), .ZN(n1968) );
NAND2_X1 U1605 ( .A1(n2014), .A2(n2015), .ZN(n2010) );
NAND2_X1 U1606 ( .A1(n2016), .A2(n2017), .ZN(n2015) );
XOR2_X1 U1607 ( .A(n2018), .B(KEYINPUT42), .Z(n2016) );
XNOR2_X1 U1608 ( .A(KEYINPUT51), .B(n2019), .ZN(n2014) );
XOR2_X1 U1609 ( .A(n2012), .B(n2011), .Z(n2013) );
NAND2_X1 U1610 ( .A1(n2020), .A2(n2021), .ZN(n2011) );
NAND2_X1 U1611 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1975), .ZN(n2021) );
NAND2_X1 U1612 ( .A1(RESTART), .A2(RMIN_REG_5__SCAN_IN), .ZN(n2020) );
NAND2_X1 U1613 ( .A1(n2022), .A2(n2023), .ZN(n2012) );
NAND2_X1 U1614 ( .A1(DATA_IN_5_), .A2(n1975), .ZN(n2023) );
NAND2_X1 U1615 ( .A1(RESTART), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2022) );
XOR2_X1 U1616 ( .A(KEYINPUT50), .B(n2001), .Z(n2004) );
NAND4_X1 U1617 ( .A1(n2024), .A2(n2025), .A3(n2026), .A4(n2027), .ZN(U284));
NOR3_X1 U1618 ( .A1(n2028), .A2(n2029), .A3(n2030), .ZN(n2027) );
NOR3_X1 U1619 ( .A1(n1931), .A2(n2031), .A3(n2032), .ZN(n2030) );
NOR2_X1 U1620 ( .A1(n1993), .A2(n2033), .ZN(n2032) );
XOR2_X1 U1621 ( .A(KEYINPUT8), .B(n1994), .Z(n2033) );
NOR2_X1 U1622 ( .A1(n2034), .A2(n2035), .ZN(n2031) );
XNOR2_X1 U1623 ( .A(KEYINPUT14), .B(n1993), .ZN(n2035) );
NAND2_X1 U1624 ( .A1(n1997), .A2(n2036), .ZN(n1993) );
NAND2_X1 U1625 ( .A1(n2037), .A2(n2038), .ZN(n2036) );
NAND2_X1 U1626 ( .A1(n2039), .A2(n2040), .ZN(n2038) );
XOR2_X1 U1627 ( .A(KEYINPUT9), .B(n2041), .Z(n2039) );
NAND3_X1 U1628 ( .A1(n2041), .A2(n2042), .A3(n2043), .ZN(n1997) );
XNOR2_X1 U1629 ( .A(n2040), .B(KEYINPUT10), .ZN(n2043) );
INV_X1 U1630 ( .A(n1994), .ZN(n2034) );
INV_X1 U1631 ( .A(n1932), .ZN(n1931) );
NOR3_X1 U1632 ( .A1(n1911), .A2(n2001), .A3(n2044), .ZN(n2029) );
NOR2_X1 U1633 ( .A1(n2045), .A2(n2046), .ZN(n2044) );
AND2_X1 U1634 ( .A1(n2045), .A2(n2046), .ZN(n2001) );
NAND2_X1 U1635 ( .A1(n2006), .A2(n2047), .ZN(n2046) );
NAND2_X1 U1636 ( .A1(n2037), .A2(n2048), .ZN(n2047) );
NAND2_X1 U1637 ( .A1(n2041), .A2(n2040), .ZN(n2048) );
NAND3_X1 U1638 ( .A1(n2042), .A2(n2040), .A3(n2041), .ZN(n2006) );
NOR2_X1 U1639 ( .A1(n2042), .A2(n1960), .ZN(n2028) );
INV_X1 U1640 ( .A(n2037), .ZN(n2042) );
XNOR2_X1 U1641 ( .A(n2049), .B(n2018), .ZN(n2037) );
NAND2_X1 U1642 ( .A1(n2050), .A2(n2051), .ZN(n2018) );
NAND2_X1 U1643 ( .A1(n2052), .A2(n2053), .ZN(n2051) );
OR2_X1 U1644 ( .A1(n2054), .A2(n2055), .ZN(n2053) );
NAND2_X1 U1645 ( .A1(n2055), .A2(n2054), .ZN(n2050) );
NAND3_X1 U1646 ( .A1(n2017), .A2(n2019), .A3(KEYINPUT63), .ZN(n2049) );
OR2_X1 U1647 ( .A1(n2056), .A2(n2057), .ZN(n2019) );
NAND2_X1 U1648 ( .A1(n2057), .A2(n2056), .ZN(n2017) );
NAND2_X1 U1649 ( .A1(n2058), .A2(n2059), .ZN(n2056) );
OR2_X1 U1650 ( .A1(REG4_REG_4__SCAN_IN), .A2(RESTART), .ZN(n2059) );
NAND2_X1 U1651 ( .A1(n2060), .A2(RESTART), .ZN(n2058) );
XOR2_X1 U1652 ( .A(RMIN_REG_4__SCAN_IN), .B(KEYINPUT32), .Z(n2060) );
AND2_X1 U1653 ( .A1(n2061), .A2(n2062), .ZN(n2057) );
NAND2_X1 U1654 ( .A1(RESTART), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2062) );
XOR2_X1 U1655 ( .A(n2063), .B(KEYINPUT31), .Z(n2061) );
NAND2_X1 U1656 ( .A1(DATA_IN_4_), .A2(n2064), .ZN(n2063) );
XOR2_X1 U1657 ( .A(RESTART), .B(KEYINPUT33), .Z(n2064) );
XOR2_X1 U1658 ( .A(n2065), .B(KEYINPUT52), .Z(n2026) );
NAND2_X1 U1659 ( .A1(n1905), .A2(RLAST_REG_3__SCAN_IN), .ZN(n2065) );
NAND2_X1 U1660 ( .A1(n1912), .A2(REG4_REG_3__SCAN_IN), .ZN(n2025) );
NAND2_X1 U1661 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1684), .ZN(n2024) );
NAND2_X1 U1662 ( .A1(n2066), .A2(n2067), .ZN(U283) );
NAND3_X1 U1663 ( .A1(n2068), .A2(n2069), .A3(n1932), .ZN(n2067) );
NAND2_X1 U1664 ( .A1(n2070), .A2(n2071), .ZN(n2069) );
NAND2_X1 U1665 ( .A1(n2072), .A2(n2073), .ZN(n2071) );
XOR2_X1 U1666 ( .A(KEYINPUT38), .B(n1994), .Z(n2068) );
NOR3_X1 U1667 ( .A1(n2074), .A2(n2075), .A3(n2070), .ZN(n1994) );
XOR2_X1 U1668 ( .A(n2076), .B(KEYINPUT20), .Z(n2066) );
NAND4_X1 U1669 ( .A1(n2077), .A2(n2078), .A3(n2079), .A4(n2080), .ZN(n2076));
NOR2_X1 U1670 ( .A1(n2081), .A2(n2082), .ZN(n2080) );
NOR2_X1 U1671 ( .A1(n2083), .A2(n1927), .ZN(n2082) );
NOR2_X1 U1672 ( .A1(n2040), .A2(n1960), .ZN(n2081) );
NAND2_X1 U1673 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n2084), .ZN(n2079) );
XOR2_X1 U1674 ( .A(KEYINPUT26), .B(n1905), .Z(n2084) );
NAND3_X1 U1675 ( .A1(n2085), .A2(n2086), .A3(n2000), .ZN(n2078) );
INV_X1 U1676 ( .A(n2045), .ZN(n2086) );
NOR3_X1 U1677 ( .A1(n2075), .A2(n2087), .A3(n2070), .ZN(n2045) );
NAND2_X1 U1678 ( .A1(n2070), .A2(n2088), .ZN(n2085) );
NAND2_X1 U1679 ( .A1(n2073), .A2(n2089), .ZN(n2088) );
XOR2_X1 U1680 ( .A(n2040), .B(n2041), .Z(n2070) );
XOR2_X1 U1681 ( .A(n2090), .B(n2054), .Z(n2040) );
NAND2_X1 U1682 ( .A1(n2091), .A2(n2092), .ZN(n2054) );
NAND2_X1 U1683 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1975), .ZN(n2092) );
NAND2_X1 U1684 ( .A1(RESTART), .A2(RMIN_REG_3__SCAN_IN), .ZN(n2091) );
XNOR2_X1 U1685 ( .A(n2052), .B(n2055), .ZN(n2090) );
AND2_X1 U1686 ( .A1(n2093), .A2(n2094), .ZN(n2055) );
NAND2_X1 U1687 ( .A1(RESTART), .A2(n1797), .ZN(n2094) );
NAND2_X1 U1688 ( .A1(n1765), .A2(n1975), .ZN(n2093) );
INV_X1 U1689 ( .A(DATA_IN_3_), .ZN(n1765) );
AND2_X1 U1690 ( .A1(n2095), .A2(n2096), .ZN(n2052) );
NAND2_X1 U1691 ( .A1(n2097), .A2(n2098), .ZN(n2096) );
NAND2_X1 U1692 ( .A1(n2099), .A2(n2100), .ZN(n2098) );
NAND2_X1 U1693 ( .A1(n2101), .A2(n2102), .ZN(n2095) );
NAND2_X1 U1694 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n2103), .ZN(n2077) );
XOR2_X1 U1695 ( .A(KEYINPUT27), .B(n1684), .Z(n2103) );
NAND4_X1 U1696 ( .A1(n2104), .A2(n2105), .A3(n2106), .A4(n2107), .ZN(U282));
NOR4_X1 U1697 ( .A1(n2108), .A2(n2109), .A3(n2110), .A4(n2111), .ZN(n2107));
AND2_X1 U1698 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1684), .ZN(n2111) );
NOR2_X1 U1699 ( .A1(n2112), .A2(n1927), .ZN(n2110) );
NOR3_X1 U1700 ( .A1(n2073), .A2(n2087), .A3(n1911), .ZN(n2109) );
INV_X1 U1701 ( .A(n2000), .ZN(n1911) );
NOR2_X1 U1702 ( .A1(n2075), .A2(n2113), .ZN(n2108) );
NAND2_X1 U1703 ( .A1(n1905), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2106) );
NAND3_X1 U1704 ( .A1(n2114), .A2(n2115), .A3(n1932), .ZN(n2105) );
NAND2_X1 U1705 ( .A1(n2074), .A2(n2116), .ZN(n2115) );
NAND2_X1 U1706 ( .A1(n2117), .A2(n2072), .ZN(n2114) );
NAND2_X1 U1707 ( .A1(n2075), .A2(n2116), .ZN(n2117) );
INV_X1 U1708 ( .A(KEYINPUT45), .ZN(n2116) );
INV_X1 U1709 ( .A(n2073), .ZN(n2075) );
NAND2_X1 U1710 ( .A1(n2118), .A2(n2119), .ZN(n2073) );
INV_X1 U1711 ( .A(n2041), .ZN(n2119) );
NOR2_X1 U1712 ( .A1(n2120), .A2(n2121), .ZN(n2041) );
NAND2_X1 U1713 ( .A1(n2121), .A2(n2120), .ZN(n2118) );
NAND2_X1 U1714 ( .A1(n1989), .A2(n2121), .ZN(n2104) );
XOR2_X1 U1715 ( .A(n2097), .B(n2122), .Z(n2121) );
NOR2_X1 U1716 ( .A1(n2123), .A2(n2124), .ZN(n2122) );
NOR2_X1 U1717 ( .A1(n2102), .A2(n2125), .ZN(n2124) );
NOR2_X1 U1718 ( .A1(n2126), .A2(n2127), .ZN(n2125) );
AND2_X1 U1719 ( .A1(KEYINPUT56), .A2(n2100), .ZN(n2127) );
NOR2_X1 U1720 ( .A1(KEYINPUT21), .A2(n2100), .ZN(n2126) );
NOR2_X1 U1721 ( .A1(n2099), .A2(n2128), .ZN(n2123) );
NOR2_X1 U1722 ( .A1(n2129), .A2(n2130), .ZN(n2128) );
NOR2_X1 U1723 ( .A1(KEYINPUT56), .A2(n2101), .ZN(n2130) );
NOR2_X1 U1724 ( .A1(KEYINPUT37), .A2(n2100), .ZN(n2129) );
INV_X1 U1725 ( .A(n2101), .ZN(n2100) );
NAND2_X1 U1726 ( .A1(n2131), .A2(n2132), .ZN(n2101) );
NAND2_X1 U1727 ( .A1(RESTART), .A2(n1764), .ZN(n2132) );
NAND2_X1 U1728 ( .A1(n2083), .A2(n1975), .ZN(n2131) );
INV_X1 U1729 ( .A(n2102), .ZN(n2099) );
NAND2_X1 U1730 ( .A1(n2133), .A2(n2134), .ZN(n2102) );
NAND2_X1 U1731 ( .A1(n2135), .A2(n2136), .ZN(n2134) );
OR2_X1 U1732 ( .A1(n2137), .A2(n2138), .ZN(n2136) );
NAND2_X1 U1733 ( .A1(n2138), .A2(n2137), .ZN(n2133) );
NAND2_X1 U1734 ( .A1(n2139), .A2(n2140), .ZN(n2097) );
NAND2_X1 U1735 ( .A1(RESTART), .A2(n1792), .ZN(n2140) );
NAND2_X1 U1736 ( .A1(n1758), .A2(n1975), .ZN(n2139) );
INV_X1 U1737 ( .A(n1960), .ZN(n1989) );
NAND3_X1 U1738 ( .A1(n2113), .A2(n2141), .A3(n2142), .ZN(U281) );
NOR3_X1 U1739 ( .A1(n2143), .A2(n2144), .A3(n2145), .ZN(n2142) );
NOR2_X1 U1740 ( .A1(n2146), .A2(n1960), .ZN(n2145) );
NAND4_X1 U1741 ( .A1(STATO_REG_1__SCAN_IN), .A2(n2147), .A3(n2148), .A4(U280), .ZN(n1960) );
NAND2_X1 U1742 ( .A1(n2149), .A2(n1975), .ZN(n2147) );
NAND3_X1 U1743 ( .A1(n2150), .A2(n2151), .A3(ENABLE), .ZN(n2149) );
AND2_X1 U1744 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1905), .ZN(n2144) );
NOR2_X1 U1745 ( .A1(n2152), .A2(ENABLE), .ZN(n1905) );
NOR2_X1 U1746 ( .A1(n2153), .A2(n1927), .ZN(n2143) );
INV_X1 U1747 ( .A(n1912), .ZN(n1927) );
NOR3_X1 U1748 ( .A1(n1824), .A2(n2152), .A3(n2151), .ZN(n1912) );
INV_X1 U1749 ( .A(AVERAGE), .ZN(n2151) );
NAND2_X1 U1750 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1684), .ZN(n2141) );
AND2_X1 U1751 ( .A1(n2154), .A2(n2155), .ZN(n2113) );
NAND2_X1 U1752 ( .A1(n2087), .A2(n2000), .ZN(n2155) );
NOR3_X1 U1753 ( .A1(n1825), .A2(n1684), .A3(n2148), .ZN(n2000) );
NAND3_X1 U1754 ( .A1(n2156), .A2(n2157), .A3(RESTART), .ZN(n2148) );
NAND2_X1 U1755 ( .A1(n2158), .A2(n1771), .ZN(n2157) );
INV_X1 U1756 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1771) );
NAND2_X1 U1757 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n2159), .ZN(n2158) );
OR2_X1 U1758 ( .A1(n2159), .A2(RMAX_REG_7__SCAN_IN), .ZN(n2156) );
NAND2_X1 U1759 ( .A1(n2160), .A2(n2161), .ZN(n2159) );
NAND2_X1 U1760 ( .A1(n2162), .A2(n1778), .ZN(n2161) );
INV_X1 U1761 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1778) );
NAND2_X1 U1762 ( .A1(n2163), .A2(n2164), .ZN(n2162) );
XOR2_X1 U1763 ( .A(n2165), .B(KEYINPUT1), .Z(n2160) );
NAND2_X1 U1764 ( .A1(n1769), .A2(n2166), .ZN(n2165) );
NAND3_X1 U1765 ( .A1(n2164), .A2(n2163), .A3(RMAX_REG_6__SCAN_IN), .ZN(n2166) );
NAND3_X1 U1766 ( .A1(n2167), .A2(n2168), .A3(n2169), .ZN(n2163) );
NAND2_X1 U1767 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2169) );
NAND3_X1 U1768 ( .A1(n2170), .A2(n2171), .A3(n2172), .ZN(n2168) );
NAND2_X1 U1769 ( .A1(n1785), .A2(n1746), .ZN(n2172) );
INV_X1 U1770 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1746) );
INV_X1 U1771 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1785) );
NAND3_X1 U1772 ( .A1(n2173), .A2(n2174), .A3(n2175), .ZN(n2171) );
NAND2_X1 U1773 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2175) );
NAND3_X1 U1774 ( .A1(n2176), .A2(n2177), .A3(n2178), .ZN(n2174) );
NAND2_X1 U1775 ( .A1(n1792), .A2(n1764), .ZN(n2178) );
INV_X1 U1776 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1764) );
INV_X1 U1777 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1792) );
NAND2_X1 U1778 ( .A1(n2179), .A2(n1761), .ZN(n2177) );
INV_X1 U1779 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1761) );
OR2_X1 U1780 ( .A1(n2180), .A2(n1796), .ZN(n2179) );
NAND2_X1 U1781 ( .A1(n2180), .A2(n1796), .ZN(n2176) );
INV_X1 U1782 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1796) );
NAND2_X1 U1783 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2173) );
NAND2_X1 U1784 ( .A1(n1797), .A2(n1754), .ZN(n2170) );
INV_X1 U1785 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1754) );
INV_X1 U1786 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1797) );
NAND2_X1 U1787 ( .A1(n2181), .A2(RMIN_REG_5__SCAN_IN), .ZN(n2167) );
XOR2_X1 U1788 ( .A(n1800), .B(KEYINPUT30), .Z(n2181) );
NAND2_X1 U1789 ( .A1(n1766), .A2(n1800), .ZN(n2164) );
INV_X1 U1790 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1800) );
INV_X1 U1791 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1766) );
INV_X1 U1792 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1769) );
INV_X1 U1793 ( .A(n2089), .ZN(n2087) );
NAND2_X1 U1794 ( .A1(n2182), .A2(n2183), .ZN(n2089) );
NAND2_X1 U1795 ( .A1(KEYINPUT49), .A2(n2184), .ZN(n2183) );
NAND2_X1 U1796 ( .A1(n2185), .A2(n2186), .ZN(n2182) );
NAND2_X1 U1797 ( .A1(KEYINPUT49), .A2(n2146), .ZN(n2186) );
NAND2_X1 U1798 ( .A1(n2074), .A2(n1932), .ZN(n2154) );
NAND2_X1 U1799 ( .A1(n2187), .A2(n2188), .ZN(n2150) );
NAND2_X1 U1800 ( .A1(n2189), .A2(n2190), .ZN(n2188) );
INV_X1 U1801 ( .A(REG4_REG_7__SCAN_IN), .ZN(n2190) );
OR2_X1 U1802 ( .A1(n2191), .A2(n1737), .ZN(n2189) );
NAND2_X1 U1803 ( .A1(n2191), .A2(n1737), .ZN(n2187) );
INV_X1 U1804 ( .A(DATA_IN_7_), .ZN(n1737) );
NAND2_X1 U1805 ( .A1(n2192), .A2(n2193), .ZN(n2191) );
NAND2_X1 U1806 ( .A1(DATA_IN_6_), .A2(n2194), .ZN(n2193) );
NAND2_X1 U1807 ( .A1(n2195), .A2(n1926), .ZN(n2194) );
INV_X1 U1808 ( .A(REG4_REG_6__SCAN_IN), .ZN(n1926) );
XOR2_X1 U1809 ( .A(KEYINPUT48), .B(n2196), .Z(n2195) );
NAND2_X1 U1810 ( .A1(n2196), .A2(REG4_REG_6__SCAN_IN), .ZN(n2192) );
AND2_X1 U1811 ( .A1(n2197), .A2(n2198), .ZN(n2196) );
NAND2_X1 U1812 ( .A1(n2199), .A2(n2200), .ZN(n2198) );
NAND2_X1 U1813 ( .A1(DATA_IN_5_), .A2(n2201), .ZN(n2200) );
INV_X1 U1814 ( .A(REG4_REG_5__SCAN_IN), .ZN(n2199) );
OR2_X1 U1815 ( .A1(n2201), .A2(DATA_IN_5_), .ZN(n2197) );
NAND2_X1 U1816 ( .A1(n2202), .A2(n2203), .ZN(n2201) );
NAND2_X1 U1817 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2203) );
NAND3_X1 U1818 ( .A1(n2204), .A2(n2205), .A3(n2206), .ZN(n2202) );
OR2_X1 U1819 ( .A1(DATA_IN_3_), .A2(REG4_REG_3__SCAN_IN), .ZN(n2206) );
NAND3_X1 U1820 ( .A1(n2207), .A2(n2208), .A3(n2209), .ZN(n2205) );
NAND2_X1 U1821 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2209) );
NAND3_X1 U1822 ( .A1(n2210), .A2(n2211), .A3(n2212), .ZN(n2208) );
NAND2_X1 U1823 ( .A1(n1758), .A2(n2083), .ZN(n2212) );
INV_X1 U1824 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2083) );
INV_X1 U1825 ( .A(DATA_IN_2_), .ZN(n1758) );
NAND2_X1 U1826 ( .A1(n2213), .A2(n2112), .ZN(n2211) );
INV_X1 U1827 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2112) );
NAND2_X1 U1828 ( .A1(n2214), .A2(n2215), .ZN(n2213) );
XOR2_X1 U1829 ( .A(KEYINPUT6), .B(DATA_IN_1_), .Z(n2215) );
INV_X1 U1830 ( .A(n2216), .ZN(n2214) );
NAND2_X1 U1831 ( .A1(n2216), .A2(n1763), .ZN(n2210) );
INV_X1 U1832 ( .A(DATA_IN_1_), .ZN(n1763) );
NAND2_X1 U1833 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2207) );
NAND2_X1 U1834 ( .A1(n2217), .A2(n1750), .ZN(n2204) );
INV_X1 U1835 ( .A(DATA_IN_4_), .ZN(n1750) );
XOR2_X1 U1836 ( .A(REG4_REG_4__SCAN_IN), .B(KEYINPUT55), .Z(n2217) );
NAND3_X1 U1837 ( .A1(U280), .A2(n1975), .A3(STATO_REG_1__SCAN_IN), .ZN(n2152) );
INV_X1 U1838 ( .A(ENABLE), .ZN(n1824) );
INV_X1 U1839 ( .A(n2072), .ZN(n2074) );
NAND2_X1 U1840 ( .A1(n2120), .A2(n2218), .ZN(n2072) );
NAND2_X1 U1841 ( .A1(n2185), .A2(n2219), .ZN(n2218) );
INV_X1 U1842 ( .A(n2184), .ZN(n2120) );
NOR2_X1 U1843 ( .A1(n2219), .A2(n2185), .ZN(n2184) );
AND3_X1 U1844 ( .A1(n2220), .A2(n2221), .A3(n2137), .ZN(n2185) );
NAND3_X1 U1845 ( .A1(n1728), .A2(n2153), .A3(n1975), .ZN(n2221) );
INV_X1 U1846 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2153) );
INV_X1 U1847 ( .A(DATA_IN_0_), .ZN(n1728) );
OR3_X1 U1848 ( .A1(RMAX_REG_0__SCAN_IN), .A2(RMIN_REG_0__SCAN_IN), .A3(n1975), .ZN(n2220) );
INV_X1 U1849 ( .A(n2146), .ZN(n2219) );
XNOR2_X1 U1850 ( .A(n2135), .B(n2222), .ZN(n2146) );
XNOR2_X1 U1851 ( .A(n2138), .B(n2137), .ZN(n2222) );
NAND2_X1 U1852 ( .A1(n2223), .A2(n2224), .ZN(n2137) );
NAND2_X1 U1853 ( .A1(RESTART), .A2(n2180), .ZN(n2224) );
NAND2_X1 U1854 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2180) );
NAND2_X1 U1855 ( .A1(n2216), .A2(n1975), .ZN(n2223) );
NAND2_X1 U1856 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2216) );
AND2_X1 U1857 ( .A1(n2225), .A2(n2226), .ZN(n2138) );
NAND2_X1 U1858 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1975), .ZN(n2226) );
NAND2_X1 U1859 ( .A1(RESTART), .A2(RMIN_REG_1__SCAN_IN), .ZN(n2225) );
AND2_X1 U1860 ( .A1(n2227), .A2(n2228), .ZN(n2135) );
NAND2_X1 U1861 ( .A1(DATA_IN_1_), .A2(n1975), .ZN(n2228) );
INV_X1 U1862 ( .A(RESTART), .ZN(n1975) );
NAND2_X1 U1863 ( .A1(RESTART), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2227) );
INV_X1 U1864 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1825) );
NOR2_X1 U1865 ( .A1(n1706), .A2(STATO_REG_1__SCAN_IN), .ZN(n2229) );
INV_X1 U1866 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1706) );
endmodule


