//Key = 1010111011110110111010100111011101101101110110101001110110110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317;

XOR2_X1 U729 ( .A(G107), .B(n1005), .Z(G9) );
NOR2_X1 U730 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
XOR2_X1 U731 ( .A(n1008), .B(KEYINPUT24), .Z(n1006) );
NAND3_X1 U732 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(G75) );
NAND2_X1 U733 ( .A1(G952), .A2(n1012), .ZN(n1011) );
NAND4_X1 U734 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
NAND4_X1 U735 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
NAND2_X1 U736 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND3_X1 U737 ( .A1(n1023), .A2(n1024), .A3(KEYINPUT12), .ZN(n1021) );
NAND3_X1 U738 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1019) );
NAND2_X1 U739 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
OR2_X1 U740 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U741 ( .A1(n1023), .A2(n1032), .ZN(n1025) );
NAND2_X1 U742 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
OR2_X1 U743 ( .A1(n1035), .A2(KEYINPUT12), .ZN(n1034) );
NAND2_X1 U744 ( .A1(n1036), .A2(n1037), .ZN(n1033) );
NAND4_X1 U745 ( .A1(n1027), .A2(n1023), .A3(n1028), .A4(n1038), .ZN(n1015) );
NAND2_X1 U746 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U747 ( .A1(n1018), .A2(n1041), .ZN(n1040) );
NAND2_X1 U748 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U749 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U750 ( .A1(n1017), .A2(n1046), .ZN(n1039) );
NAND2_X1 U751 ( .A1(n1007), .A2(n1047), .ZN(n1046) );
NAND2_X1 U752 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
INV_X1 U753 ( .A(n1022), .ZN(n1027) );
XOR2_X1 U754 ( .A(KEYINPUT41), .B(G953), .Z(n1014) );
NAND4_X1 U755 ( .A1(n1036), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1009) );
NOR4_X1 U756 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
XOR2_X1 U757 ( .A(n1057), .B(n1058), .Z(n1056) );
XNOR2_X1 U758 ( .A(G469), .B(n1059), .ZN(n1055) );
XOR2_X1 U759 ( .A(n1060), .B(n1061), .Z(n1054) );
XNOR2_X1 U760 ( .A(n1062), .B(n1063), .ZN(n1053) );
XOR2_X1 U761 ( .A(n1064), .B(KEYINPUT45), .Z(n1063) );
NOR3_X1 U762 ( .A1(n1065), .A2(n1048), .A3(n1044), .ZN(n1051) );
NOR2_X1 U763 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
XOR2_X1 U764 ( .A(KEYINPUT61), .B(n1068), .Z(n1067) );
INV_X1 U765 ( .A(n1069), .ZN(n1066) );
XOR2_X1 U766 ( .A(KEYINPUT43), .B(n1070), .Z(n1050) );
XOR2_X1 U767 ( .A(n1071), .B(n1072), .Z(G72) );
NAND2_X1 U768 ( .A1(G953), .A2(n1073), .ZN(n1072) );
NAND2_X1 U769 ( .A1(G900), .A2(G227), .ZN(n1073) );
NAND2_X1 U770 ( .A1(KEYINPUT2), .A2(n1074), .ZN(n1071) );
XOR2_X1 U771 ( .A(n1075), .B(n1076), .Z(n1074) );
NAND2_X1 U772 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U773 ( .A(KEYINPUT53), .B(G953), .Z(n1077) );
NAND2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1075) );
NAND2_X1 U775 ( .A1(G953), .A2(n1081), .ZN(n1080) );
XOR2_X1 U776 ( .A(n1082), .B(n1083), .Z(n1079) );
NAND2_X1 U777 ( .A1(KEYINPUT5), .A2(n1084), .ZN(n1082) );
XNOR2_X1 U778 ( .A(n1085), .B(n1086), .ZN(n1084) );
NAND2_X1 U779 ( .A1(KEYINPUT48), .A2(n1087), .ZN(n1085) );
XOR2_X1 U780 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U781 ( .A1(KEYINPUT40), .A2(n1090), .ZN(n1088) );
XOR2_X1 U782 ( .A(n1091), .B(n1092), .Z(G69) );
XOR2_X1 U783 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U784 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XOR2_X1 U785 ( .A(n1097), .B(KEYINPUT11), .Z(n1096) );
INV_X1 U786 ( .A(n1098), .ZN(n1095) );
NAND3_X1 U787 ( .A1(n1099), .A2(n1100), .A3(KEYINPUT13), .ZN(n1093) );
NAND2_X1 U788 ( .A1(G953), .A2(n1101), .ZN(n1100) );
NAND2_X1 U789 ( .A1(G953), .A2(n1102), .ZN(n1091) );
NAND2_X1 U790 ( .A1(G898), .A2(G224), .ZN(n1102) );
NOR2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(G66) );
NOR3_X1 U792 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1104) );
NOR3_X1 U793 ( .A1(n1108), .A2(n1060), .A3(n1109), .ZN(n1107) );
NOR2_X1 U794 ( .A1(n1110), .A2(n1111), .ZN(n1106) );
NOR2_X1 U795 ( .A1(n1013), .A2(n1060), .ZN(n1110) );
NOR2_X1 U796 ( .A1(n1103), .A2(n1112), .ZN(G63) );
NOR3_X1 U797 ( .A1(n1062), .A2(n1113), .A3(n1114), .ZN(n1112) );
AND3_X1 U798 ( .A1(n1115), .A2(G478), .A3(n1116), .ZN(n1114) );
NOR2_X1 U799 ( .A1(n1117), .A2(n1115), .ZN(n1113) );
NOR2_X1 U800 ( .A1(n1013), .A2(n1064), .ZN(n1117) );
INV_X1 U801 ( .A(G478), .ZN(n1064) );
NOR2_X1 U802 ( .A1(n1103), .A2(n1118), .ZN(G60) );
XOR2_X1 U803 ( .A(n1119), .B(n1120), .Z(n1118) );
AND2_X1 U804 ( .A1(G475), .A2(n1116), .ZN(n1120) );
NAND2_X1 U805 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
XNOR2_X1 U806 ( .A(KEYINPUT58), .B(KEYINPUT25), .ZN(n1121) );
XOR2_X1 U807 ( .A(n1123), .B(n1124), .Z(G6) );
NOR3_X1 U808 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(G57) );
NOR2_X1 U809 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U810 ( .A(KEYINPUT18), .B(n1130), .Z(n1129) );
NOR2_X1 U811 ( .A1(n1131), .A2(n1132), .ZN(n1126) );
XNOR2_X1 U812 ( .A(n1130), .B(KEYINPUT16), .ZN(n1132) );
XNOR2_X1 U813 ( .A(n1133), .B(n1134), .ZN(n1130) );
AND2_X1 U814 ( .A1(G472), .A2(n1116), .ZN(n1134) );
NAND2_X1 U815 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NAND2_X1 U816 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U817 ( .A(n1139), .B(KEYINPUT23), .Z(n1135) );
OR2_X1 U818 ( .A1(n1138), .A2(n1137), .ZN(n1139) );
INV_X1 U819 ( .A(n1128), .ZN(n1131) );
XOR2_X1 U820 ( .A(n1010), .B(KEYINPUT22), .Z(n1125) );
NOR2_X1 U821 ( .A1(n1103), .A2(n1140), .ZN(G54) );
NOR2_X1 U822 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XOR2_X1 U823 ( .A(n1143), .B(KEYINPUT29), .Z(n1142) );
NAND2_X1 U824 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NOR2_X1 U825 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
XNOR2_X1 U826 ( .A(n1146), .B(n1147), .ZN(n1145) );
XOR2_X1 U827 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U828 ( .A(n1150), .B(n1151), .ZN(n1149) );
XNOR2_X1 U829 ( .A(KEYINPUT31), .B(KEYINPUT26), .ZN(n1148) );
XOR2_X1 U830 ( .A(n1152), .B(n1086), .Z(n1146) );
XOR2_X1 U831 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U832 ( .A1(n1155), .A2(KEYINPUT8), .ZN(n1153) );
XNOR2_X1 U833 ( .A(G140), .B(n1156), .ZN(n1155) );
NOR2_X1 U834 ( .A1(G110), .A2(KEYINPUT50), .ZN(n1156) );
AND2_X1 U835 ( .A1(n1116), .A2(G469), .ZN(n1144) );
NOR3_X1 U836 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(G51) );
NOR3_X1 U837 ( .A1(n1160), .A2(G953), .A3(G952), .ZN(n1159) );
INV_X1 U838 ( .A(KEYINPUT21), .ZN(n1160) );
NOR2_X1 U839 ( .A1(KEYINPUT21), .A2(n1010), .ZN(n1158) );
INV_X1 U840 ( .A(n1103), .ZN(n1010) );
NOR2_X1 U841 ( .A1(n1097), .A2(G952), .ZN(n1103) );
XOR2_X1 U842 ( .A(n1161), .B(n1162), .Z(n1157) );
XOR2_X1 U843 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U844 ( .A1(n1058), .A2(n1109), .ZN(n1164) );
INV_X1 U845 ( .A(n1116), .ZN(n1109) );
NOR2_X1 U846 ( .A1(n1165), .A2(n1013), .ZN(n1116) );
NOR2_X1 U847 ( .A1(n1078), .A2(n1098), .ZN(n1013) );
NAND2_X1 U848 ( .A1(n1166), .A2(n1167), .ZN(n1098) );
NOR4_X1 U849 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
INV_X1 U850 ( .A(n1124), .ZN(n1169) );
NAND4_X1 U851 ( .A1(n1172), .A2(n1030), .A3(n1173), .A4(n1028), .ZN(n1124) );
NOR4_X1 U852 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1166) );
NOR2_X1 U853 ( .A1(n1008), .A2(n1007), .ZN(n1177) );
INV_X1 U854 ( .A(n1178), .ZN(n1007) );
NAND4_X1 U855 ( .A1(n1173), .A2(n1031), .A3(n1028), .A4(n1179), .ZN(n1008) );
NOR4_X1 U856 ( .A1(n1042), .A2(n1035), .A3(n1180), .A4(n1181), .ZN(n1176) );
XOR2_X1 U857 ( .A(KEYINPUT37), .B(n1023), .Z(n1181) );
INV_X1 U858 ( .A(n1173), .ZN(n1042) );
INV_X1 U859 ( .A(n1182), .ZN(n1175) );
INV_X1 U860 ( .A(n1183), .ZN(n1174) );
NAND4_X1 U861 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1078) );
NOR4_X1 U862 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187) );
NOR2_X1 U863 ( .A1(n1192), .A2(n1193), .ZN(n1186) );
INV_X1 U864 ( .A(n1194), .ZN(n1193) );
NOR2_X1 U865 ( .A1(n1195), .A2(n1196), .ZN(n1161) );
NOR2_X1 U866 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NOR2_X1 U867 ( .A1(n1199), .A2(n1200), .ZN(n1195) );
XOR2_X1 U868 ( .A(n1198), .B(KEYINPUT56), .Z(n1200) );
XOR2_X1 U869 ( .A(n1201), .B(G125), .Z(n1198) );
NAND2_X1 U870 ( .A1(KEYINPUT33), .A2(n1202), .ZN(n1201) );
INV_X1 U871 ( .A(n1197), .ZN(n1199) );
XOR2_X1 U872 ( .A(n1192), .B(n1203), .Z(G48) );
XOR2_X1 U873 ( .A(KEYINPUT28), .B(G146), .Z(n1203) );
AND3_X1 U874 ( .A1(n1204), .A2(n1178), .A3(n1030), .ZN(n1192) );
XNOR2_X1 U875 ( .A(G143), .B(n1184), .ZN(G45) );
NAND4_X1 U876 ( .A1(n1205), .A2(n1178), .A3(n1206), .A4(n1207), .ZN(n1184) );
XOR2_X1 U877 ( .A(G140), .B(n1191), .Z(G42) );
AND3_X1 U878 ( .A1(n1018), .A2(n1173), .A3(n1208), .ZN(n1191) );
XOR2_X1 U879 ( .A(G137), .B(n1190), .Z(G39) );
AND3_X1 U880 ( .A1(n1018), .A2(n1204), .A3(n1023), .ZN(n1190) );
XOR2_X1 U881 ( .A(n1090), .B(n1185), .Z(G36) );
NAND3_X1 U882 ( .A1(n1205), .A2(n1031), .A3(n1018), .ZN(n1185) );
INV_X1 U883 ( .A(G134), .ZN(n1090) );
XOR2_X1 U884 ( .A(G131), .B(n1189), .Z(G33) );
AND3_X1 U885 ( .A1(n1018), .A2(n1205), .A3(n1030), .ZN(n1189) );
AND3_X1 U886 ( .A1(n1173), .A2(n1209), .A3(n1024), .ZN(n1205) );
NOR2_X1 U887 ( .A1(n1210), .A2(n1211), .ZN(n1018) );
XOR2_X1 U888 ( .A(G128), .B(n1188), .Z(G30) );
AND3_X1 U889 ( .A1(n1178), .A2(n1031), .A3(n1204), .ZN(n1188) );
AND4_X1 U890 ( .A1(n1173), .A2(n1212), .A3(n1209), .A4(n1037), .ZN(n1204) );
XOR2_X1 U891 ( .A(G101), .B(n1213), .Z(G3) );
NOR2_X1 U892 ( .A1(n1035), .A2(n1214), .ZN(n1213) );
XOR2_X1 U893 ( .A(n1215), .B(n1194), .Z(G27) );
NAND3_X1 U894 ( .A1(n1208), .A2(n1178), .A3(n1017), .ZN(n1194) );
AND4_X1 U895 ( .A1(n1036), .A2(n1030), .A3(n1209), .A4(n1037), .ZN(n1208) );
NAND2_X1 U896 ( .A1(n1022), .A2(n1216), .ZN(n1209) );
NAND4_X1 U897 ( .A1(G953), .A2(G902), .A3(n1217), .A4(n1081), .ZN(n1216) );
INV_X1 U898 ( .A(G900), .ZN(n1081) );
XNOR2_X1 U899 ( .A(n1168), .B(n1218), .ZN(G24) );
NAND2_X1 U900 ( .A1(KEYINPUT34), .A2(G122), .ZN(n1218) );
AND4_X1 U901 ( .A1(n1219), .A2(n1028), .A3(n1206), .A4(n1207), .ZN(n1168) );
NOR2_X1 U902 ( .A1(n1037), .A2(n1212), .ZN(n1028) );
XOR2_X1 U903 ( .A(n1220), .B(n1182), .Z(G21) );
NAND4_X1 U904 ( .A1(n1219), .A2(n1023), .A3(n1212), .A4(n1037), .ZN(n1182) );
NAND2_X1 U905 ( .A1(n1221), .A2(n1222), .ZN(G18) );
NAND2_X1 U906 ( .A1(G116), .A2(n1183), .ZN(n1222) );
XOR2_X1 U907 ( .A(KEYINPUT62), .B(n1223), .Z(n1221) );
NOR2_X1 U908 ( .A1(G116), .A2(n1183), .ZN(n1223) );
NAND3_X1 U909 ( .A1(n1024), .A2(n1031), .A3(n1219), .ZN(n1183) );
AND2_X1 U910 ( .A1(n1224), .A2(n1206), .ZN(n1031) );
XOR2_X1 U911 ( .A(G113), .B(n1171), .Z(G15) );
AND3_X1 U912 ( .A1(n1030), .A2(n1024), .A3(n1219), .ZN(n1171) );
AND2_X1 U913 ( .A1(n1172), .A2(n1017), .ZN(n1219) );
AND2_X1 U914 ( .A1(n1045), .A2(n1225), .ZN(n1017) );
INV_X1 U915 ( .A(n1035), .ZN(n1024) );
NAND2_X1 U916 ( .A1(n1226), .A2(n1212), .ZN(n1035) );
NOR2_X1 U917 ( .A1(n1206), .A2(n1224), .ZN(n1030) );
XOR2_X1 U918 ( .A(G110), .B(n1170), .Z(G12) );
NOR3_X1 U919 ( .A1(n1212), .A2(n1226), .A3(n1214), .ZN(n1170) );
NAND3_X1 U920 ( .A1(n1023), .A2(n1173), .A3(n1172), .ZN(n1214) );
INV_X1 U921 ( .A(n1180), .ZN(n1172) );
NAND2_X1 U922 ( .A1(n1178), .A2(n1179), .ZN(n1180) );
NAND2_X1 U923 ( .A1(n1022), .A2(n1227), .ZN(n1179) );
NAND4_X1 U924 ( .A1(G953), .A2(G902), .A3(n1217), .A4(n1101), .ZN(n1227) );
INV_X1 U925 ( .A(G898), .ZN(n1101) );
NAND3_X1 U926 ( .A1(n1217), .A2(n1097), .A3(G952), .ZN(n1022) );
NAND2_X1 U927 ( .A1(G237), .A2(G234), .ZN(n1217) );
NOR2_X1 U928 ( .A1(n1049), .A2(n1210), .ZN(n1178) );
XNOR2_X1 U929 ( .A(n1048), .B(KEYINPUT51), .ZN(n1210) );
AND2_X1 U930 ( .A1(G214), .A2(n1228), .ZN(n1048) );
INV_X1 U931 ( .A(n1211), .ZN(n1049) );
XOR2_X1 U932 ( .A(n1057), .B(n1229), .Z(n1211) );
NOR2_X1 U933 ( .A1(n1230), .A2(KEYINPUT54), .ZN(n1229) );
INV_X1 U934 ( .A(n1058), .ZN(n1230) );
NAND2_X1 U935 ( .A1(G210), .A2(n1228), .ZN(n1058) );
NAND2_X1 U936 ( .A1(n1165), .A2(n1231), .ZN(n1228) );
INV_X1 U937 ( .A(G237), .ZN(n1231) );
NAND2_X1 U938 ( .A1(n1232), .A2(n1165), .ZN(n1057) );
XOR2_X1 U939 ( .A(n1233), .B(n1234), .Z(n1232) );
XOR2_X1 U940 ( .A(G125), .B(n1163), .Z(n1234) );
AND2_X1 U941 ( .A1(G224), .A2(n1097), .ZN(n1163) );
XOR2_X1 U942 ( .A(n1202), .B(n1197), .Z(n1233) );
XOR2_X1 U943 ( .A(n1099), .B(KEYINPUT3), .Z(n1202) );
XNOR2_X1 U944 ( .A(n1235), .B(n1236), .ZN(n1099) );
XOR2_X1 U945 ( .A(n1237), .B(n1238), .Z(n1236) );
XNOR2_X1 U946 ( .A(n1239), .B(n1240), .ZN(n1238) );
NAND2_X1 U947 ( .A1(KEYINPUT63), .A2(n1220), .ZN(n1240) );
INV_X1 U948 ( .A(G119), .ZN(n1220) );
NAND2_X1 U949 ( .A1(n1241), .A2(KEYINPUT55), .ZN(n1239) );
XOR2_X1 U950 ( .A(n1242), .B(G104), .Z(n1241) );
NAND2_X1 U951 ( .A1(KEYINPUT0), .A2(n1243), .ZN(n1242) );
INV_X1 U952 ( .A(G107), .ZN(n1243) );
XOR2_X1 U953 ( .A(n1244), .B(n1245), .Z(n1235) );
NOR2_X1 U954 ( .A1(KEYINPUT19), .A2(G113), .ZN(n1245) );
XOR2_X1 U955 ( .A(n1246), .B(G110), .Z(n1244) );
NOR2_X1 U956 ( .A1(n1045), .A2(n1044), .ZN(n1173) );
INV_X1 U957 ( .A(n1225), .ZN(n1044) );
NAND2_X1 U958 ( .A1(G221), .A2(n1247), .ZN(n1225) );
XNOR2_X1 U959 ( .A(n1059), .B(n1248), .ZN(n1045) );
NOR2_X1 U960 ( .A1(G469), .A2(KEYINPUT42), .ZN(n1248) );
NAND2_X1 U961 ( .A1(n1249), .A2(n1165), .ZN(n1059) );
XOR2_X1 U962 ( .A(n1250), .B(n1251), .Z(n1249) );
XNOR2_X1 U963 ( .A(n1151), .B(n1252), .ZN(n1251) );
XOR2_X1 U964 ( .A(n1253), .B(n1254), .Z(n1252) );
NOR2_X1 U965 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XOR2_X1 U966 ( .A(n1257), .B(KEYINPUT52), .Z(n1256) );
NAND2_X1 U967 ( .A1(n1150), .A2(n1086), .ZN(n1257) );
NOR2_X1 U968 ( .A1(n1150), .A2(n1086), .ZN(n1255) );
XOR2_X1 U969 ( .A(G128), .B(n1258), .Z(n1086) );
AND2_X1 U970 ( .A1(n1259), .A2(n1260), .ZN(n1150) );
NAND2_X1 U971 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U972 ( .A(n1246), .B(KEYINPUT1), .Z(n1262) );
XOR2_X1 U973 ( .A(n1123), .B(G107), .Z(n1261) );
NAND2_X1 U974 ( .A1(n1263), .A2(n1264), .ZN(n1259) );
XOR2_X1 U975 ( .A(G107), .B(G104), .Z(n1264) );
XOR2_X1 U976 ( .A(n1246), .B(KEYINPUT59), .Z(n1263) );
INV_X1 U977 ( .A(G101), .ZN(n1246) );
NAND2_X1 U978 ( .A1(n1265), .A2(KEYINPUT36), .ZN(n1253) );
XNOR2_X1 U979 ( .A(n1154), .B(KEYINPUT15), .ZN(n1265) );
AND2_X1 U980 ( .A1(G227), .A2(n1097), .ZN(n1151) );
XNOR2_X1 U981 ( .A(G110), .B(n1266), .ZN(n1250) );
XOR2_X1 U982 ( .A(KEYINPUT20), .B(G140), .Z(n1266) );
NOR2_X1 U983 ( .A1(n1207), .A2(n1206), .ZN(n1023) );
XNOR2_X1 U984 ( .A(n1062), .B(n1267), .ZN(n1206) );
NOR2_X1 U985 ( .A1(G478), .A2(KEYINPUT35), .ZN(n1267) );
NOR2_X1 U986 ( .A1(n1115), .A2(G902), .ZN(n1062) );
XNOR2_X1 U987 ( .A(n1268), .B(n1269), .ZN(n1115) );
XOR2_X1 U988 ( .A(G128), .B(n1270), .Z(n1269) );
XOR2_X1 U989 ( .A(G143), .B(G134), .Z(n1270) );
XOR2_X1 U990 ( .A(n1271), .B(n1272), .Z(n1268) );
INV_X1 U991 ( .A(n1237), .ZN(n1272) );
XOR2_X1 U992 ( .A(n1273), .B(n1274), .Z(n1237) );
XOR2_X1 U993 ( .A(n1275), .B(G107), .Z(n1271) );
NAND2_X1 U994 ( .A1(G217), .A2(n1276), .ZN(n1275) );
INV_X1 U995 ( .A(n1224), .ZN(n1207) );
NOR2_X1 U996 ( .A1(n1277), .A2(n1070), .ZN(n1224) );
NOR2_X1 U997 ( .A1(n1069), .A2(n1068), .ZN(n1070) );
AND2_X1 U998 ( .A1(n1068), .A2(n1069), .ZN(n1277) );
NAND2_X1 U999 ( .A1(n1122), .A2(n1165), .ZN(n1069) );
XNOR2_X1 U1000 ( .A(n1278), .B(n1279), .ZN(n1122) );
XOR2_X1 U1001 ( .A(n1083), .B(n1280), .Z(n1279) );
XOR2_X1 U1002 ( .A(n1281), .B(n1258), .Z(n1280) );
NAND2_X1 U1003 ( .A1(n1282), .A2(G214), .ZN(n1281) );
XOR2_X1 U1004 ( .A(n1283), .B(n1284), .Z(n1278) );
NOR2_X1 U1005 ( .A1(KEYINPUT49), .A2(n1285), .ZN(n1284) );
XOR2_X1 U1006 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U1007 ( .A(G113), .B(KEYINPUT47), .ZN(n1287) );
NAND2_X1 U1008 ( .A1(KEYINPUT14), .A2(n1273), .ZN(n1286) );
INV_X1 U1009 ( .A(G122), .ZN(n1273) );
XOR2_X1 U1010 ( .A(G131), .B(n1123), .Z(n1283) );
INV_X1 U1011 ( .A(G104), .ZN(n1123) );
XOR2_X1 U1012 ( .A(G475), .B(KEYINPUT38), .Z(n1068) );
INV_X1 U1013 ( .A(n1037), .ZN(n1226) );
NAND2_X1 U1014 ( .A1(n1288), .A2(n1289), .ZN(n1037) );
NAND2_X1 U1015 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
XOR2_X1 U1016 ( .A(KEYINPUT4), .B(n1292), .Z(n1288) );
NOR2_X1 U1017 ( .A1(n1290), .A2(n1291), .ZN(n1292) );
XOR2_X1 U1018 ( .A(KEYINPUT17), .B(n1105), .Z(n1291) );
INV_X1 U1019 ( .A(n1061), .ZN(n1105) );
NAND2_X1 U1020 ( .A1(n1108), .A2(n1165), .ZN(n1061) );
INV_X1 U1021 ( .A(n1111), .ZN(n1108) );
XOR2_X1 U1022 ( .A(n1293), .B(n1294), .Z(n1111) );
XOR2_X1 U1023 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1024 ( .A(n1297), .B(n1298), .Z(n1296) );
NAND2_X1 U1025 ( .A1(KEYINPUT46), .A2(n1299), .ZN(n1298) );
INV_X1 U1026 ( .A(G146), .ZN(n1299) );
NAND2_X1 U1027 ( .A1(n1276), .A2(G221), .ZN(n1297) );
AND2_X1 U1028 ( .A1(G234), .A2(n1097), .ZN(n1276) );
INV_X1 U1029 ( .A(G953), .ZN(n1097) );
INV_X1 U1030 ( .A(n1083), .ZN(n1295) );
XOR2_X1 U1031 ( .A(n1215), .B(G140), .Z(n1083) );
INV_X1 U1032 ( .A(G125), .ZN(n1215) );
XOR2_X1 U1033 ( .A(n1300), .B(n1301), .Z(n1293) );
XOR2_X1 U1034 ( .A(KEYINPUT44), .B(G137), .Z(n1301) );
NAND2_X1 U1035 ( .A1(n1302), .A2(KEYINPUT30), .ZN(n1300) );
XOR2_X1 U1036 ( .A(n1303), .B(n1304), .Z(n1302) );
NOR2_X1 U1037 ( .A1(KEYINPUT57), .A2(G119), .ZN(n1304) );
XNOR2_X1 U1038 ( .A(G110), .B(G128), .ZN(n1303) );
INV_X1 U1039 ( .A(n1060), .ZN(n1290) );
NAND2_X1 U1040 ( .A1(G217), .A2(n1247), .ZN(n1060) );
NAND2_X1 U1041 ( .A1(G234), .A2(n1165), .ZN(n1247) );
INV_X1 U1042 ( .A(n1036), .ZN(n1212) );
XOR2_X1 U1043 ( .A(n1305), .B(G472), .Z(n1036) );
NAND2_X1 U1044 ( .A1(n1306), .A2(n1165), .ZN(n1305) );
INV_X1 U1045 ( .A(G902), .ZN(n1165) );
XOR2_X1 U1046 ( .A(n1137), .B(n1307), .Z(n1306) );
XNOR2_X1 U1047 ( .A(n1308), .B(n1309), .ZN(n1307) );
NOR2_X1 U1048 ( .A1(KEYINPUT32), .A2(n1128), .ZN(n1309) );
XOR2_X1 U1049 ( .A(n1310), .B(G101), .Z(n1128) );
NAND2_X1 U1050 ( .A1(n1282), .A2(G210), .ZN(n1310) );
NOR2_X1 U1051 ( .A1(G953), .A2(G237), .ZN(n1282) );
NAND2_X1 U1052 ( .A1(KEYINPUT10), .A2(n1138), .ZN(n1308) );
XOR2_X1 U1053 ( .A(G113), .B(n1311), .Z(n1138) );
NOR2_X1 U1054 ( .A1(KEYINPUT60), .A2(n1312), .ZN(n1311) );
XOR2_X1 U1055 ( .A(G119), .B(n1274), .Z(n1312) );
XOR2_X1 U1056 ( .A(G116), .B(KEYINPUT39), .Z(n1274) );
XOR2_X1 U1057 ( .A(n1154), .B(n1197), .Z(n1137) );
XOR2_X1 U1058 ( .A(n1313), .B(n1314), .Z(n1197) );
XOR2_X1 U1059 ( .A(KEYINPUT7), .B(G128), .Z(n1314) );
NAND2_X1 U1060 ( .A1(KEYINPUT9), .A2(n1258), .ZN(n1313) );
XOR2_X1 U1061 ( .A(G143), .B(G146), .Z(n1258) );
XNOR2_X1 U1062 ( .A(n1315), .B(n1316), .ZN(n1154) );
INV_X1 U1063 ( .A(n1089), .ZN(n1316) );
XNOR2_X1 U1064 ( .A(G131), .B(G137), .ZN(n1089) );
XOR2_X1 U1065 ( .A(n1317), .B(KEYINPUT6), .Z(n1315) );
NAND2_X1 U1066 ( .A1(KEYINPUT27), .A2(G134), .ZN(n1317) );
endmodule


