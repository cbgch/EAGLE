//Key = 0111010011000010010001100110111010001000010101000001111101111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356;

XNOR2_X1 U744 ( .A(G107), .B(n1027), .ZN(G9) );
NAND4_X1 U745 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(G75) );
NAND3_X1 U746 ( .A1(n1032), .A2(n1033), .A3(G952), .ZN(n1031) );
NAND2_X1 U747 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NAND4_X1 U748 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
NAND2_X1 U749 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NAND2_X1 U750 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
OR2_X1 U751 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U752 ( .A1(n1046), .A2(n1047), .ZN(n1040) );
OR2_X1 U753 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND3_X1 U754 ( .A1(n1042), .A2(n1050), .A3(n1046), .ZN(n1034) );
NAND2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND3_X1 U756 ( .A1(n1053), .A2(n1054), .A3(n1036), .ZN(n1052) );
OR2_X1 U757 ( .A1(n1039), .A2(n1037), .ZN(n1054) );
NAND3_X1 U758 ( .A1(n1055), .A2(n1056), .A3(n1039), .ZN(n1053) );
OR2_X1 U759 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NAND2_X1 U760 ( .A1(n1037), .A2(n1059), .ZN(n1051) );
NOR2_X1 U761 ( .A1(G953), .A2(n1060), .ZN(n1030) );
NOR4_X1 U762 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1060) );
NOR2_X1 U763 ( .A1(KEYINPUT59), .A2(n1065), .ZN(n1064) );
XOR2_X1 U764 ( .A(n1066), .B(n1067), .Z(n1063) );
NAND2_X1 U765 ( .A1(KEYINPUT51), .A2(n1068), .ZN(n1066) );
NAND3_X1 U766 ( .A1(n1039), .A2(n1058), .A3(n1069), .ZN(n1062) );
XOR2_X1 U767 ( .A(n1070), .B(n1071), .Z(n1069) );
XOR2_X1 U768 ( .A(KEYINPUT5), .B(G472), .Z(n1071) );
NOR2_X1 U769 ( .A1(KEYINPUT42), .A2(n1072), .ZN(n1070) );
NAND4_X1 U770 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1061) );
NOR2_X1 U771 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U772 ( .A(G478), .B(n1079), .Z(n1078) );
XOR2_X1 U773 ( .A(n1080), .B(n1081), .Z(n1075) );
NAND3_X1 U774 ( .A1(KEYINPUT59), .A2(n1065), .A3(G469), .ZN(n1074) );
NAND2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1073) );
INV_X1 U776 ( .A(G469), .ZN(n1083) );
NAND2_X1 U777 ( .A1(KEYINPUT59), .A2(n1084), .ZN(n1082) );
XNOR2_X1 U778 ( .A(KEYINPUT62), .B(n1065), .ZN(n1084) );
XOR2_X1 U779 ( .A(n1085), .B(n1086), .Z(G72) );
NOR2_X1 U780 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U781 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR2_X1 U782 ( .A1(KEYINPUT12), .A2(n1091), .ZN(n1085) );
XOR2_X1 U783 ( .A(n1092), .B(n1093), .Z(n1091) );
NOR3_X1 U784 ( .A1(n1094), .A2(KEYINPUT44), .A3(n1095), .ZN(n1093) );
XOR2_X1 U785 ( .A(n1096), .B(n1097), .Z(n1095) );
XOR2_X1 U786 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U787 ( .A1(KEYINPUT10), .A2(n1100), .ZN(n1098) );
XOR2_X1 U788 ( .A(KEYINPUT34), .B(n1101), .Z(n1094) );
NOR2_X1 U789 ( .A1(G900), .A2(n1088), .ZN(n1101) );
NAND2_X1 U790 ( .A1(n1088), .A2(n1102), .ZN(n1092) );
NAND3_X1 U791 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
XOR2_X1 U792 ( .A(n1106), .B(KEYINPUT48), .Z(n1105) );
XOR2_X1 U793 ( .A(n1107), .B(n1108), .Z(G69) );
XOR2_X1 U794 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U795 ( .A1(n1029), .A2(n1111), .ZN(n1110) );
XOR2_X1 U796 ( .A(KEYINPUT63), .B(G953), .Z(n1111) );
NAND2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(n1109) );
NAND2_X1 U798 ( .A1(G953), .A2(n1114), .ZN(n1113) );
XOR2_X1 U799 ( .A(n1115), .B(n1116), .Z(n1112) );
XNOR2_X1 U800 ( .A(n1117), .B(n1118), .ZN(n1116) );
NAND2_X1 U801 ( .A1(KEYINPUT57), .A2(n1119), .ZN(n1117) );
XOR2_X1 U802 ( .A(G104), .B(n1120), .Z(n1115) );
NOR2_X1 U803 ( .A1(KEYINPUT24), .A2(n1121), .ZN(n1120) );
XOR2_X1 U804 ( .A(G122), .B(G110), .Z(n1121) );
NAND2_X1 U805 ( .A1(G953), .A2(n1122), .ZN(n1107) );
NAND2_X1 U806 ( .A1(G898), .A2(G224), .ZN(n1122) );
NOR2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(G66) );
NOR3_X1 U808 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1124) );
NOR3_X1 U809 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1127) );
AND2_X1 U810 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NAND2_X1 U811 ( .A1(n1081), .A2(n1131), .ZN(n1128) );
XNOR2_X1 U812 ( .A(KEYINPUT21), .B(n1132), .ZN(n1131) );
INV_X1 U813 ( .A(n1080), .ZN(n1125) );
NOR2_X1 U814 ( .A1(n1123), .A2(n1133), .ZN(G63) );
NOR3_X1 U815 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1133) );
NOR2_X1 U816 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U817 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
XNOR2_X1 U818 ( .A(KEYINPUT40), .B(n1141), .ZN(n1140) );
INV_X1 U819 ( .A(KEYINPUT28), .ZN(n1139) );
AND3_X1 U820 ( .A1(n1138), .A2(n1141), .A3(KEYINPUT28), .ZN(n1135) );
NOR2_X1 U821 ( .A1(KEYINPUT28), .A2(n1141), .ZN(n1134) );
NAND2_X1 U822 ( .A1(n1142), .A2(G478), .ZN(n1141) );
NOR2_X1 U823 ( .A1(n1123), .A2(n1143), .ZN(G60) );
XNOR2_X1 U824 ( .A(n1144), .B(n1145), .ZN(n1143) );
AND2_X1 U825 ( .A1(G475), .A2(n1142), .ZN(n1145) );
XNOR2_X1 U826 ( .A(n1146), .B(n1147), .ZN(G6) );
NOR2_X1 U827 ( .A1(KEYINPUT19), .A2(n1148), .ZN(n1147) );
NOR3_X1 U828 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(G57) );
NOR2_X1 U829 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NOR2_X1 U830 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NOR2_X1 U831 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NOR2_X1 U832 ( .A1(n1158), .A2(n1159), .ZN(n1154) );
NOR2_X1 U833 ( .A1(G101), .A2(n1160), .ZN(n1150) );
NOR2_X1 U834 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U835 ( .A1(n1157), .A2(n1159), .ZN(n1162) );
NOR2_X1 U836 ( .A1(n1158), .A2(n1156), .ZN(n1161) );
XOR2_X1 U837 ( .A(n1159), .B(KEYINPUT58), .Z(n1156) );
XOR2_X1 U838 ( .A(n1163), .B(n1164), .Z(n1159) );
XOR2_X1 U839 ( .A(n1165), .B(n1166), .Z(n1163) );
AND2_X1 U840 ( .A1(G472), .A2(n1142), .ZN(n1166) );
NAND2_X1 U841 ( .A1(KEYINPUT60), .A2(n1167), .ZN(n1165) );
INV_X1 U842 ( .A(n1157), .ZN(n1158) );
XOR2_X1 U843 ( .A(KEYINPUT20), .B(n1123), .Z(n1149) );
NOR2_X1 U844 ( .A1(n1123), .A2(n1168), .ZN(G54) );
XOR2_X1 U845 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U846 ( .A1(KEYINPUT38), .A2(n1171), .ZN(n1170) );
XOR2_X1 U847 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U848 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NOR2_X1 U849 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NOR2_X1 U850 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NOR2_X1 U851 ( .A1(n1180), .A2(n1181), .ZN(n1178) );
XOR2_X1 U852 ( .A(KEYINPUT61), .B(n1182), .Z(n1181) );
INV_X1 U853 ( .A(n1183), .ZN(n1176) );
NOR2_X1 U854 ( .A1(n1179), .A2(n1183), .ZN(n1174) );
NAND2_X1 U855 ( .A1(n1180), .A2(n1182), .ZN(n1183) );
XNOR2_X1 U856 ( .A(G110), .B(n1184), .ZN(n1180) );
XOR2_X1 U857 ( .A(KEYINPUT56), .B(G140), .Z(n1184) );
INV_X1 U858 ( .A(KEYINPUT43), .ZN(n1179) );
NAND2_X1 U859 ( .A1(n1142), .A2(G469), .ZN(n1169) );
INV_X1 U860 ( .A(n1185), .ZN(n1142) );
NOR2_X1 U861 ( .A1(n1123), .A2(n1186), .ZN(G51) );
NOR3_X1 U862 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1186) );
NOR3_X1 U863 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1189) );
INV_X1 U864 ( .A(n1193), .ZN(n1192) );
NOR3_X1 U865 ( .A1(n1185), .A2(KEYINPUT4), .A3(n1068), .ZN(n1191) );
NOR2_X1 U866 ( .A1(KEYINPUT30), .A2(n1193), .ZN(n1188) );
NOR3_X1 U867 ( .A1(n1185), .A2(n1194), .A3(n1068), .ZN(n1187) );
NOR2_X1 U868 ( .A1(n1195), .A2(n1190), .ZN(n1194) );
INV_X1 U869 ( .A(KEYINPUT30), .ZN(n1190) );
NOR2_X1 U870 ( .A1(KEYINPUT4), .A2(n1193), .ZN(n1195) );
XNOR2_X1 U871 ( .A(n1196), .B(n1167), .ZN(n1193) );
XOR2_X1 U872 ( .A(n1197), .B(n1198), .Z(n1196) );
NOR2_X1 U873 ( .A1(G125), .A2(KEYINPUT31), .ZN(n1198) );
NAND2_X1 U874 ( .A1(G902), .A2(n1132), .ZN(n1185) );
NAND2_X1 U875 ( .A1(n1199), .A2(n1029), .ZN(n1132) );
AND2_X1 U876 ( .A1(n1200), .A2(n1201), .ZN(n1029) );
AND4_X1 U877 ( .A1(n1202), .A2(n1203), .A3(n1027), .A4(n1204), .ZN(n1201) );
NAND3_X1 U878 ( .A1(n1042), .A2(n1205), .A3(n1045), .ZN(n1027) );
AND4_X1 U879 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1146), .ZN(n1200) );
NAND3_X1 U880 ( .A1(n1042), .A2(n1205), .A3(n1044), .ZN(n1146) );
XNOR2_X1 U881 ( .A(n1028), .B(KEYINPUT2), .ZN(n1199) );
AND3_X1 U882 ( .A1(n1104), .A2(n1106), .A3(n1103), .ZN(n1028) );
AND4_X1 U883 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1103) );
NOR3_X1 U884 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1212) );
NAND3_X1 U885 ( .A1(n1216), .A2(n1059), .A3(n1044), .ZN(n1104) );
NOR2_X1 U886 ( .A1(n1088), .A2(G952), .ZN(n1123) );
XOR2_X1 U887 ( .A(G146), .B(n1217), .Z(G48) );
NOR3_X1 U888 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1217) );
INV_X1 U889 ( .A(n1059), .ZN(n1219) );
XOR2_X1 U890 ( .A(KEYINPUT29), .B(n1044), .Z(n1218) );
XOR2_X1 U891 ( .A(n1221), .B(n1211), .Z(G45) );
NAND4_X1 U892 ( .A1(n1222), .A2(n1059), .A3(n1048), .A4(n1223), .ZN(n1211) );
NOR3_X1 U893 ( .A1(n1056), .A2(n1224), .A3(n1225), .ZN(n1223) );
NAND3_X1 U894 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(G42) );
NAND2_X1 U895 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NAND2_X1 U896 ( .A1(KEYINPUT50), .A2(n1231), .ZN(n1227) );
NAND2_X1 U897 ( .A1(n1232), .A2(n1106), .ZN(n1231) );
XOR2_X1 U898 ( .A(KEYINPUT47), .B(G140), .Z(n1232) );
NAND2_X1 U899 ( .A1(n1233), .A2(n1234), .ZN(n1226) );
INV_X1 U900 ( .A(KEYINPUT50), .ZN(n1234) );
NAND2_X1 U901 ( .A1(n1235), .A2(n1236), .ZN(n1233) );
NAND2_X1 U902 ( .A1(KEYINPUT47), .A2(n1230), .ZN(n1236) );
OR3_X1 U903 ( .A1(n1229), .A2(KEYINPUT47), .A3(n1230), .ZN(n1235) );
INV_X1 U904 ( .A(n1106), .ZN(n1229) );
NAND3_X1 U905 ( .A1(n1044), .A2(n1237), .A3(n1049), .ZN(n1106) );
XNOR2_X1 U906 ( .A(G137), .B(n1209), .ZN(G39) );
NAND4_X1 U907 ( .A1(n1046), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1209) );
XOR2_X1 U908 ( .A(n1210), .B(n1240), .Z(G36) );
NAND2_X1 U909 ( .A1(KEYINPUT9), .A2(G134), .ZN(n1240) );
NAND3_X1 U910 ( .A1(n1237), .A2(n1045), .A3(n1048), .ZN(n1210) );
XOR2_X1 U911 ( .A(n1241), .B(n1215), .Z(G33) );
AND3_X1 U912 ( .A1(n1044), .A2(n1237), .A3(n1048), .ZN(n1215) );
AND3_X1 U913 ( .A1(n1222), .A2(n1059), .A3(n1037), .ZN(n1237) );
NOR2_X1 U914 ( .A1(n1057), .A2(n1242), .ZN(n1037) );
INV_X1 U915 ( .A(n1243), .ZN(n1242) );
NAND2_X1 U916 ( .A1(KEYINPUT17), .A2(n1244), .ZN(n1241) );
XOR2_X1 U917 ( .A(G128), .B(n1214), .Z(G30) );
AND3_X1 U918 ( .A1(n1045), .A2(n1245), .A3(n1216), .ZN(n1214) );
INV_X1 U919 ( .A(n1220), .ZN(n1216) );
NAND4_X1 U920 ( .A1(n1222), .A2(n1246), .A3(n1238), .A4(n1239), .ZN(n1220) );
XOR2_X1 U921 ( .A(n1153), .B(n1208), .Z(G3) );
NAND3_X1 U922 ( .A1(n1048), .A2(n1205), .A3(n1046), .ZN(n1208) );
INV_X1 U923 ( .A(G101), .ZN(n1153) );
XOR2_X1 U924 ( .A(G125), .B(n1213), .Z(G27) );
AND4_X1 U925 ( .A1(n1246), .A2(n1039), .A3(n1222), .A4(n1247), .ZN(n1213) );
AND3_X1 U926 ( .A1(n1049), .A2(n1044), .A3(n1036), .ZN(n1247) );
AND3_X1 U927 ( .A1(n1248), .A2(n1249), .A3(n1033), .ZN(n1222) );
NAND2_X1 U928 ( .A1(G953), .A2(n1250), .ZN(n1248) );
NAND2_X1 U929 ( .A1(G902), .A2(n1090), .ZN(n1250) );
INV_X1 U930 ( .A(G900), .ZN(n1090) );
XOR2_X1 U931 ( .A(n1251), .B(n1207), .Z(G24) );
NAND4_X1 U932 ( .A1(n1252), .A2(n1042), .A3(n1253), .A4(n1077), .ZN(n1207) );
NOR2_X1 U933 ( .A1(n1239), .A2(n1238), .ZN(n1042) );
XOR2_X1 U934 ( .A(n1254), .B(n1255), .Z(G21) );
NAND2_X1 U935 ( .A1(KEYINPUT36), .A2(n1256), .ZN(n1255) );
INV_X1 U936 ( .A(n1203), .ZN(n1256) );
NAND4_X1 U937 ( .A1(n1252), .A2(n1046), .A3(n1238), .A4(n1239), .ZN(n1203) );
XNOR2_X1 U938 ( .A(G116), .B(n1202), .ZN(G18) );
NAND3_X1 U939 ( .A1(n1048), .A2(n1045), .A3(n1252), .ZN(n1202) );
NOR2_X1 U940 ( .A1(n1077), .A2(n1225), .ZN(n1045) );
INV_X1 U941 ( .A(n1253), .ZN(n1225) );
XOR2_X1 U942 ( .A(n1206), .B(n1257), .Z(G15) );
XNOR2_X1 U943 ( .A(G113), .B(KEYINPUT18), .ZN(n1257) );
NAND3_X1 U944 ( .A1(n1048), .A2(n1044), .A3(n1252), .ZN(n1206) );
AND3_X1 U945 ( .A1(n1258), .A2(n1039), .A3(n1036), .ZN(n1252) );
NOR2_X1 U946 ( .A1(n1253), .A2(n1224), .ZN(n1044) );
AND2_X1 U947 ( .A1(n1259), .A2(n1238), .ZN(n1048) );
XNOR2_X1 U948 ( .A(G110), .B(n1204), .ZN(G12) );
NAND3_X1 U949 ( .A1(n1049), .A2(n1205), .A3(n1046), .ZN(n1204) );
NOR2_X1 U950 ( .A1(n1077), .A2(n1253), .ZN(n1046) );
XOR2_X1 U951 ( .A(n1260), .B(n1261), .Z(n1253) );
NOR2_X1 U952 ( .A1(KEYINPUT46), .A2(n1079), .ZN(n1261) );
AND2_X1 U953 ( .A1(n1138), .A2(n1130), .ZN(n1079) );
XOR2_X1 U954 ( .A(n1262), .B(n1263), .Z(n1138) );
XOR2_X1 U955 ( .A(G134), .B(n1264), .Z(n1263) );
NOR2_X1 U956 ( .A1(KEYINPUT0), .A2(n1265), .ZN(n1264) );
XNOR2_X1 U957 ( .A(G107), .B(n1266), .ZN(n1265) );
XOR2_X1 U958 ( .A(G122), .B(G116), .Z(n1266) );
XOR2_X1 U959 ( .A(n1267), .B(n1268), .Z(n1262) );
AND2_X1 U960 ( .A1(n1269), .A2(G217), .ZN(n1268) );
NAND2_X1 U961 ( .A1(n1270), .A2(n1271), .ZN(n1267) );
NAND2_X1 U962 ( .A1(G143), .A2(n1272), .ZN(n1271) );
XOR2_X1 U963 ( .A(KEYINPUT41), .B(n1273), .Z(n1270) );
NOR2_X1 U964 ( .A1(G143), .A2(n1272), .ZN(n1273) );
XNOR2_X1 U965 ( .A(G478), .B(KEYINPUT15), .ZN(n1260) );
INV_X1 U966 ( .A(n1224), .ZN(n1077) );
XOR2_X1 U967 ( .A(n1274), .B(G475), .Z(n1224) );
NAND2_X1 U968 ( .A1(n1144), .A2(n1130), .ZN(n1274) );
XNOR2_X1 U969 ( .A(n1275), .B(n1276), .ZN(n1144) );
XOR2_X1 U970 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U971 ( .A(G113), .B(KEYINPUT25), .ZN(n1278) );
NAND3_X1 U972 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1277) );
OR2_X1 U973 ( .A1(n1282), .A2(KEYINPUT52), .ZN(n1281) );
NAND3_X1 U974 ( .A1(KEYINPUT52), .A2(n1282), .A3(n1221), .ZN(n1280) );
NAND2_X1 U975 ( .A1(G143), .A2(n1283), .ZN(n1279) );
NAND2_X1 U976 ( .A1(n1284), .A2(KEYINPUT52), .ZN(n1283) );
XOR2_X1 U977 ( .A(n1282), .B(KEYINPUT13), .Z(n1284) );
NAND3_X1 U978 ( .A1(n1285), .A2(n1088), .A3(G214), .ZN(n1282) );
XOR2_X1 U979 ( .A(n1096), .B(n1286), .Z(n1275) );
XOR2_X1 U980 ( .A(n1287), .B(n1288), .Z(n1096) );
AND2_X1 U981 ( .A1(n1258), .A2(n1245), .ZN(n1205) );
XOR2_X1 U982 ( .A(n1059), .B(KEYINPUT16), .Z(n1245) );
NOR2_X1 U983 ( .A1(n1036), .A2(n1289), .ZN(n1059) );
INV_X1 U984 ( .A(n1039), .ZN(n1289) );
NAND2_X1 U985 ( .A1(G221), .A2(n1290), .ZN(n1039) );
XOR2_X1 U986 ( .A(n1065), .B(G469), .Z(n1036) );
NAND3_X1 U987 ( .A1(n1291), .A2(n1292), .A3(n1130), .ZN(n1065) );
NAND2_X1 U988 ( .A1(KEYINPUT1), .A2(n1293), .ZN(n1292) );
XOR2_X1 U989 ( .A(n1172), .B(n1294), .Z(n1293) );
OR3_X1 U990 ( .A1(n1172), .A2(n1294), .A3(KEYINPUT1), .ZN(n1291) );
XNOR2_X1 U991 ( .A(n1295), .B(n1182), .ZN(n1294) );
NOR2_X1 U992 ( .A1(n1089), .A2(G953), .ZN(n1182) );
INV_X1 U993 ( .A(G227), .ZN(n1089) );
NAND2_X1 U994 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
OR2_X1 U995 ( .A1(n1230), .A2(G110), .ZN(n1297) );
XOR2_X1 U996 ( .A(n1298), .B(KEYINPUT23), .Z(n1296) );
NAND2_X1 U997 ( .A1(G110), .A2(n1230), .ZN(n1298) );
INV_X1 U998 ( .A(G140), .ZN(n1230) );
XOR2_X1 U999 ( .A(n1299), .B(n1300), .Z(n1172) );
XOR2_X1 U1000 ( .A(n1287), .B(n1301), .Z(n1300) );
XOR2_X1 U1001 ( .A(n1302), .B(n1118), .Z(n1301) );
NAND2_X1 U1002 ( .A1(KEYINPUT54), .A2(n1148), .ZN(n1302) );
XOR2_X1 U1003 ( .A(n1244), .B(n1303), .Z(n1287) );
INV_X1 U1004 ( .A(G131), .ZN(n1244) );
XOR2_X1 U1005 ( .A(n1304), .B(n1099), .Z(n1299) );
XOR2_X1 U1006 ( .A(G128), .B(G143), .Z(n1099) );
AND4_X1 U1007 ( .A1(n1246), .A2(n1033), .A3(n1305), .A4(n1249), .ZN(n1258) );
NAND2_X1 U1008 ( .A1(n1306), .A2(n1088), .ZN(n1249) );
INV_X1 U1009 ( .A(G952), .ZN(n1306) );
NAND2_X1 U1010 ( .A1(G953), .A2(n1307), .ZN(n1305) );
NAND2_X1 U1011 ( .A1(G902), .A2(n1114), .ZN(n1307) );
INV_X1 U1012 ( .A(G898), .ZN(n1114) );
NAND2_X1 U1013 ( .A1(n1308), .A2(G234), .ZN(n1033) );
XOR2_X1 U1014 ( .A(n1285), .B(KEYINPUT26), .Z(n1308) );
INV_X1 U1015 ( .A(n1056), .ZN(n1246) );
NAND2_X1 U1016 ( .A1(n1243), .A2(n1057), .ZN(n1056) );
NAND2_X1 U1017 ( .A1(n1309), .A2(n1310), .ZN(n1057) );
NAND2_X1 U1018 ( .A1(n1067), .A2(n1068), .ZN(n1310) );
XOR2_X1 U1019 ( .A(KEYINPUT22), .B(n1311), .Z(n1309) );
NOR2_X1 U1020 ( .A1(n1067), .A2(n1068), .ZN(n1311) );
NAND2_X1 U1021 ( .A1(G210), .A2(n1312), .ZN(n1068) );
AND2_X1 U1022 ( .A1(n1313), .A2(n1130), .ZN(n1067) );
XOR2_X1 U1023 ( .A(n1314), .B(n1197), .Z(n1313) );
XOR2_X1 U1024 ( .A(n1315), .B(n1316), .Z(n1197) );
XOR2_X1 U1025 ( .A(n1118), .B(n1317), .Z(n1316) );
XOR2_X1 U1026 ( .A(G110), .B(n1318), .Z(n1317) );
AND2_X1 U1027 ( .A1(n1088), .A2(G224), .ZN(n1318) );
XOR2_X1 U1028 ( .A(G107), .B(G101), .Z(n1118) );
XNOR2_X1 U1029 ( .A(n1286), .B(n1119), .ZN(n1315) );
XNOR2_X1 U1030 ( .A(n1319), .B(n1320), .ZN(n1119) );
NOR2_X1 U1031 ( .A1(KEYINPUT11), .A2(n1254), .ZN(n1320) );
INV_X1 U1032 ( .A(G119), .ZN(n1254) );
XOR2_X1 U1033 ( .A(n1148), .B(n1251), .Z(n1286) );
INV_X1 U1034 ( .A(G122), .ZN(n1251) );
INV_X1 U1035 ( .A(G104), .ZN(n1148) );
NAND2_X1 U1036 ( .A1(KEYINPUT53), .A2(n1321), .ZN(n1314) );
XNOR2_X1 U1037 ( .A(G125), .B(n1167), .ZN(n1321) );
XOR2_X1 U1038 ( .A(n1058), .B(KEYINPUT35), .Z(n1243) );
NAND2_X1 U1039 ( .A1(G214), .A2(n1312), .ZN(n1058) );
NAND2_X1 U1040 ( .A1(n1285), .A2(n1130), .ZN(n1312) );
NOR2_X1 U1041 ( .A1(n1238), .A2(n1259), .ZN(n1049) );
INV_X1 U1042 ( .A(n1239), .ZN(n1259) );
NAND3_X1 U1043 ( .A1(n1322), .A2(n1323), .A3(n1324), .ZN(n1239) );
NAND2_X1 U1044 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NAND3_X1 U1045 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1326) );
NAND2_X1 U1046 ( .A1(KEYINPUT32), .A2(KEYINPUT27), .ZN(n1329) );
NAND2_X1 U1047 ( .A1(KEYINPUT37), .A2(n1080), .ZN(n1328) );
NAND2_X1 U1048 ( .A1(n1330), .A2(n1331), .ZN(n1327) );
INV_X1 U1049 ( .A(KEYINPUT37), .ZN(n1331) );
NAND2_X1 U1050 ( .A1(n1080), .A2(n1332), .ZN(n1330) );
NAND2_X1 U1051 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
INV_X1 U1052 ( .A(n1335), .ZN(n1325) );
NAND4_X1 U1053 ( .A1(n1335), .A2(n1080), .A3(KEYINPUT32), .A4(n1333), .ZN(n1323) );
INV_X1 U1054 ( .A(KEYINPUT27), .ZN(n1333) );
NAND2_X1 U1055 ( .A1(KEYINPUT27), .A2(n1336), .ZN(n1322) );
NAND2_X1 U1056 ( .A1(n1080), .A2(n1337), .ZN(n1336) );
NAND2_X1 U1057 ( .A1(n1335), .A2(n1334), .ZN(n1337) );
INV_X1 U1058 ( .A(KEYINPUT32), .ZN(n1334) );
XNOR2_X1 U1059 ( .A(n1081), .B(KEYINPUT45), .ZN(n1335) );
AND2_X1 U1060 ( .A1(G217), .A2(n1290), .ZN(n1081) );
NAND2_X1 U1061 ( .A1(G234), .A2(n1130), .ZN(n1290) );
NAND2_X1 U1062 ( .A1(n1129), .A2(n1130), .ZN(n1080) );
XOR2_X1 U1063 ( .A(n1338), .B(n1288), .Z(n1129) );
XOR2_X1 U1064 ( .A(G125), .B(G140), .Z(n1288) );
XOR2_X1 U1065 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1066 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1067 ( .A(G137), .B(G128), .Z(n1342) );
XOR2_X1 U1068 ( .A(KEYINPUT55), .B(KEYINPUT39), .Z(n1341) );
XOR2_X1 U1069 ( .A(n1343), .B(n1344), .Z(n1339) );
XOR2_X1 U1070 ( .A(n1345), .B(n1303), .Z(n1344) );
NOR2_X1 U1071 ( .A1(G110), .A2(KEYINPUT33), .ZN(n1345) );
XOR2_X1 U1072 ( .A(n1346), .B(G119), .Z(n1343) );
NAND2_X1 U1073 ( .A1(G221), .A2(n1269), .ZN(n1346) );
AND2_X1 U1074 ( .A1(G234), .A2(n1088), .ZN(n1269) );
XNOR2_X1 U1075 ( .A(n1072), .B(G472), .ZN(n1238) );
NAND2_X1 U1076 ( .A1(n1347), .A2(n1130), .ZN(n1072) );
INV_X1 U1077 ( .A(G902), .ZN(n1130) );
XOR2_X1 U1078 ( .A(n1348), .B(n1349), .Z(n1347) );
XOR2_X1 U1079 ( .A(n1164), .B(n1167), .Z(n1349) );
XOR2_X1 U1080 ( .A(n1272), .B(n1350), .Z(n1167) );
NOR2_X1 U1081 ( .A1(KEYINPUT7), .A2(n1351), .ZN(n1350) );
XOR2_X1 U1082 ( .A(n1352), .B(n1303), .Z(n1351) );
XOR2_X1 U1083 ( .A(G146), .B(KEYINPUT14), .Z(n1303) );
XOR2_X1 U1084 ( .A(n1221), .B(KEYINPUT8), .Z(n1352) );
INV_X1 U1085 ( .A(G143), .ZN(n1221) );
INV_X1 U1086 ( .A(G128), .ZN(n1272) );
XNOR2_X1 U1087 ( .A(n1353), .B(n1354), .ZN(n1164) );
XOR2_X1 U1088 ( .A(G131), .B(G119), .Z(n1354) );
XNOR2_X1 U1089 ( .A(n1304), .B(n1319), .ZN(n1353) );
XNOR2_X1 U1090 ( .A(G113), .B(G116), .ZN(n1319) );
XNOR2_X1 U1091 ( .A(n1355), .B(n1100), .ZN(n1304) );
XNOR2_X1 U1092 ( .A(G134), .B(G137), .ZN(n1100) );
XNOR2_X1 U1093 ( .A(KEYINPUT49), .B(KEYINPUT3), .ZN(n1355) );
XOR2_X1 U1094 ( .A(n1157), .B(n1356), .Z(n1348) );
NOR2_X1 U1095 ( .A1(G101), .A2(KEYINPUT6), .ZN(n1356) );
NAND3_X1 U1096 ( .A1(n1285), .A2(n1088), .A3(G210), .ZN(n1157) );
INV_X1 U1097 ( .A(G953), .ZN(n1088) );
INV_X1 U1098 ( .A(G237), .ZN(n1285) );
endmodule


