//Key = 0011101101100110101110010010011011001000000100111100100100011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252;

XOR2_X1 U692 ( .A(G107), .B(n948), .Z(G9) );
NAND4_X1 U693 ( .A1(n949), .A2(n950), .A3(n951), .A4(n952), .ZN(G75) );
NOR3_X1 U694 ( .A1(n953), .A2(G953), .A3(n954), .ZN(n952) );
NOR2_X1 U695 ( .A1(n955), .A2(n956), .ZN(n953) );
NOR2_X1 U696 ( .A1(n957), .A2(n958), .ZN(n955) );
NOR2_X1 U697 ( .A1(n959), .A2(n960), .ZN(n958) );
INV_X1 U698 ( .A(n961), .ZN(n960) );
NOR2_X1 U699 ( .A1(n962), .A2(n963), .ZN(n959) );
NOR2_X1 U700 ( .A1(n964), .A2(n965), .ZN(n963) );
NOR3_X1 U701 ( .A1(n966), .A2(n967), .A3(n968), .ZN(n964) );
NOR3_X1 U702 ( .A1(n969), .A2(KEYINPUT52), .A3(n970), .ZN(n968) );
INV_X1 U703 ( .A(n971), .ZN(n970) );
NOR2_X1 U704 ( .A1(n972), .A2(n973), .ZN(n967) );
NOR2_X1 U705 ( .A1(n974), .A2(n975), .ZN(n972) );
AND2_X1 U706 ( .A1(n971), .A2(KEYINPUT52), .ZN(n974) );
NOR2_X1 U707 ( .A1(n976), .A2(n977), .ZN(n966) );
NOR2_X1 U708 ( .A1(n978), .A2(n979), .ZN(n976) );
INV_X1 U709 ( .A(n980), .ZN(n979) );
NOR2_X1 U710 ( .A1(n981), .A2(n982), .ZN(n978) );
NOR3_X1 U711 ( .A1(n977), .A2(n983), .A3(n973), .ZN(n962) );
NOR2_X1 U712 ( .A1(n984), .A2(n985), .ZN(n983) );
NOR2_X1 U713 ( .A1(n986), .A2(n987), .ZN(n984) );
NOR4_X1 U714 ( .A1(n988), .A2(n973), .A3(n977), .A4(n965), .ZN(n957) );
INV_X1 U715 ( .A(n989), .ZN(n977) );
NOR2_X1 U716 ( .A1(n990), .A2(n991), .ZN(n988) );
NAND4_X1 U717 ( .A1(n992), .A2(n993), .A3(n994), .A4(n995), .ZN(n950) );
NOR4_X1 U718 ( .A1(n996), .A2(n997), .A3(n998), .A4(n999), .ZN(n995) );
XOR2_X1 U719 ( .A(n1000), .B(n1001), .Z(n998) );
NOR2_X1 U720 ( .A1(G472), .A2(KEYINPUT45), .ZN(n1001) );
INV_X1 U721 ( .A(n987), .ZN(n996) );
NOR2_X1 U722 ( .A1(n1002), .A2(n1003), .ZN(n994) );
XNOR2_X1 U723 ( .A(G475), .B(n1004), .ZN(n1003) );
XOR2_X1 U724 ( .A(n1005), .B(n1006), .Z(n1002) );
XOR2_X1 U725 ( .A(n1007), .B(KEYINPUT24), .Z(n993) );
XNOR2_X1 U726 ( .A(n1008), .B(KEYINPUT44), .ZN(n992) );
XOR2_X1 U727 ( .A(n1009), .B(n1010), .Z(G72) );
XOR2_X1 U728 ( .A(n1011), .B(n1012), .Z(n1010) );
NOR2_X1 U729 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
XOR2_X1 U730 ( .A(n1015), .B(n1016), .Z(n1014) );
XOR2_X1 U731 ( .A(n1017), .B(KEYINPUT32), .Z(n1016) );
NAND3_X1 U732 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1017) );
NAND2_X1 U733 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
OR3_X1 U734 ( .A1(n1022), .A2(n1021), .A3(KEYINPUT54), .ZN(n1019) );
NAND2_X1 U735 ( .A1(KEYINPUT20), .A2(n1023), .ZN(n1022) );
NAND2_X1 U736 ( .A1(KEYINPUT54), .A2(n1024), .ZN(n1018) );
INV_X1 U737 ( .A(n1023), .ZN(n1024) );
NOR3_X1 U738 ( .A1(n1025), .A2(KEYINPUT27), .A3(G953), .ZN(n1011) );
NOR2_X1 U739 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
XOR2_X1 U740 ( .A(KEYINPUT21), .B(n954), .Z(n1027) );
NOR2_X1 U741 ( .A1(n1028), .A2(n1029), .ZN(n1009) );
AND2_X1 U742 ( .A1(G227), .A2(G900), .ZN(n1028) );
XOR2_X1 U743 ( .A(n1030), .B(n1031), .Z(G69) );
NOR2_X1 U744 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
XOR2_X1 U745 ( .A(KEYINPUT57), .B(n1034), .Z(n1033) );
NAND3_X1 U746 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1030) );
INV_X1 U747 ( .A(n1032), .ZN(n1037) );
NAND2_X1 U748 ( .A1(G953), .A2(n1038), .ZN(n1036) );
NAND2_X1 U749 ( .A1(n1039), .A2(n1029), .ZN(n1035) );
NAND3_X1 U750 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
XOR2_X1 U751 ( .A(n1043), .B(KEYINPUT51), .Z(n1042) );
XNOR2_X1 U752 ( .A(KEYINPUT23), .B(n1044), .ZN(n1041) );
NOR2_X1 U753 ( .A1(n1045), .A2(n1046), .ZN(G66) );
XOR2_X1 U754 ( .A(n1047), .B(n1048), .Z(n1046) );
NOR2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U756 ( .A1(n1045), .A2(n1051), .ZN(G63) );
XOR2_X1 U757 ( .A(n1052), .B(n1053), .Z(n1051) );
NAND2_X1 U758 ( .A1(KEYINPUT48), .A2(n1054), .ZN(n1053) );
INV_X1 U759 ( .A(n1055), .ZN(n1054) );
NAND2_X1 U760 ( .A1(n1056), .A2(G478), .ZN(n1052) );
NOR2_X1 U761 ( .A1(n1045), .A2(n1057), .ZN(G60) );
XOR2_X1 U762 ( .A(n1058), .B(n1059), .Z(n1057) );
AND2_X1 U763 ( .A1(G475), .A2(n1056), .ZN(n1058) );
XNOR2_X1 U764 ( .A(G104), .B(n1043), .ZN(G6) );
NOR2_X1 U765 ( .A1(n1045), .A2(n1060), .ZN(G57) );
XOR2_X1 U766 ( .A(n1061), .B(n1062), .Z(n1060) );
NAND3_X1 U767 ( .A1(n1056), .A2(G472), .A3(KEYINPUT6), .ZN(n1061) );
INV_X1 U768 ( .A(n1050), .ZN(n1056) );
NOR3_X1 U769 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(G54) );
NOR3_X1 U770 ( .A1(n1066), .A2(G953), .A3(G952), .ZN(n1065) );
AND2_X1 U771 ( .A1(n1066), .A2(n1045), .ZN(n1064) );
INV_X1 U772 ( .A(KEYINPUT1), .ZN(n1066) );
XOR2_X1 U773 ( .A(n1067), .B(n1068), .Z(n1063) );
XOR2_X1 U774 ( .A(n1069), .B(n1070), .Z(n1068) );
XOR2_X1 U775 ( .A(n1071), .B(n1072), .Z(n1070) );
NOR2_X1 U776 ( .A1(n1005), .A2(n1050), .ZN(n1072) );
XOR2_X1 U777 ( .A(n1073), .B(n1074), .Z(n1069) );
XOR2_X1 U778 ( .A(n1075), .B(n1076), .Z(n1067) );
XOR2_X1 U779 ( .A(KEYINPUT38), .B(G140), .Z(n1076) );
XNOR2_X1 U780 ( .A(KEYINPUT43), .B(KEYINPUT50), .ZN(n1075) );
NOR2_X1 U781 ( .A1(n1045), .A2(n1077), .ZN(G51) );
NOR2_X1 U782 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XOR2_X1 U783 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U784 ( .A1(n1082), .A2(n1050), .ZN(n1081) );
NAND2_X1 U785 ( .A1(G902), .A2(n1083), .ZN(n1050) );
NAND3_X1 U786 ( .A1(n1084), .A2(n1085), .A3(n949), .ZN(n1083) );
INV_X1 U787 ( .A(n1026), .ZN(n949) );
NAND4_X1 U788 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1026) );
AND4_X1 U789 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1089) );
OR2_X1 U790 ( .A1(n1094), .A2(n1095), .ZN(n1088) );
NAND2_X1 U791 ( .A1(n1096), .A2(n1097), .ZN(n1086) );
XOR2_X1 U792 ( .A(n1098), .B(KEYINPUT47), .Z(n1096) );
XOR2_X1 U793 ( .A(KEYINPUT22), .B(n951), .Z(n1084) );
AND3_X1 U794 ( .A1(n1043), .A2(n1044), .A3(n1040), .ZN(n951) );
AND4_X1 U795 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1040) );
NOR3_X1 U796 ( .A1(n948), .A2(n1103), .A3(n1104), .ZN(n1102) );
AND3_X1 U797 ( .A1(n961), .A2(n1105), .A3(n971), .ZN(n948) );
NAND3_X1 U798 ( .A1(n961), .A2(n1105), .A3(n975), .ZN(n1043) );
NOR2_X1 U799 ( .A1(KEYINPUT12), .A2(n1106), .ZN(n1080) );
AND2_X1 U800 ( .A1(n1106), .A2(KEYINPUT12), .ZN(n1078) );
XNOR2_X1 U801 ( .A(n1107), .B(KEYINPUT2), .ZN(n1106) );
NOR2_X1 U802 ( .A1(n1029), .A2(G952), .ZN(n1045) );
XNOR2_X1 U803 ( .A(G146), .B(n1087), .ZN(G48) );
NAND3_X1 U804 ( .A1(n975), .A2(n1108), .A3(n1109), .ZN(n1087) );
XOR2_X1 U805 ( .A(n1093), .B(n1110), .Z(G45) );
NAND2_X1 U806 ( .A1(KEYINPUT7), .A2(G143), .ZN(n1110) );
NAND4_X1 U807 ( .A1(n1109), .A2(n990), .A3(n999), .A4(n1111), .ZN(n1093) );
XOR2_X1 U808 ( .A(n1112), .B(n1092), .Z(G42) );
NAND3_X1 U809 ( .A1(n991), .A2(n975), .A3(n1113), .ZN(n1092) );
XNOR2_X1 U810 ( .A(n1091), .B(n1114), .ZN(G39) );
NOR2_X1 U811 ( .A1(KEYINPUT42), .A2(n1115), .ZN(n1114) );
NAND3_X1 U812 ( .A1(n989), .A2(n1108), .A3(n1113), .ZN(n1091) );
NAND2_X1 U813 ( .A1(n1116), .A2(n1117), .ZN(G36) );
NAND2_X1 U814 ( .A1(G134), .A2(n1090), .ZN(n1117) );
XOR2_X1 U815 ( .A(KEYINPUT18), .B(n1118), .Z(n1116) );
NOR2_X1 U816 ( .A1(G134), .A2(n1090), .ZN(n1118) );
NAND2_X1 U817 ( .A1(n1097), .A2(n971), .ZN(n1090) );
INV_X1 U818 ( .A(n1119), .ZN(n1097) );
XOR2_X1 U819 ( .A(G131), .B(n1120), .Z(G33) );
NOR2_X1 U820 ( .A1(n1098), .A2(n1119), .ZN(n1120) );
NAND2_X1 U821 ( .A1(n1113), .A2(n990), .ZN(n1119) );
NOR3_X1 U822 ( .A1(n980), .A2(n1121), .A3(n965), .ZN(n1113) );
NAND2_X1 U823 ( .A1(n1007), .A2(n987), .ZN(n965) );
INV_X1 U824 ( .A(n1122), .ZN(n1121) );
XOR2_X1 U825 ( .A(G128), .B(n954), .Z(G30) );
INV_X1 U826 ( .A(n1085), .ZN(n954) );
NAND3_X1 U827 ( .A1(n1108), .A2(n971), .A3(n1109), .ZN(n1085) );
AND2_X1 U828 ( .A1(n1123), .A2(n1122), .ZN(n1109) );
XOR2_X1 U829 ( .A(n1124), .B(n1101), .Z(G3) );
NAND3_X1 U830 ( .A1(n989), .A2(n1105), .A3(n990), .ZN(n1101) );
XOR2_X1 U831 ( .A(G125), .B(n1125), .Z(G27) );
NOR2_X1 U832 ( .A1(n1126), .A2(n1095), .ZN(n1125) );
XOR2_X1 U833 ( .A(n1094), .B(KEYINPUT34), .Z(n1126) );
NAND4_X1 U834 ( .A1(n991), .A2(n975), .A3(n969), .A4(n1122), .ZN(n1094) );
NAND2_X1 U835 ( .A1(n956), .A2(n1127), .ZN(n1122) );
NAND3_X1 U836 ( .A1(G902), .A2(n1128), .A3(n1013), .ZN(n1127) );
NOR2_X1 U837 ( .A1(n1029), .A2(G900), .ZN(n1013) );
XOR2_X1 U838 ( .A(n1099), .B(n1129), .Z(G24) );
NAND2_X1 U839 ( .A1(KEYINPUT30), .A2(G122), .ZN(n1129) );
NAND4_X1 U840 ( .A1(n1130), .A2(n961), .A3(n999), .A4(n1111), .ZN(n1099) );
NOR2_X1 U841 ( .A1(n1008), .A2(n1131), .ZN(n961) );
XNOR2_X1 U842 ( .A(G119), .B(n1044), .ZN(G21) );
NAND3_X1 U843 ( .A1(n1130), .A2(n1108), .A3(n989), .ZN(n1044) );
AND2_X1 U844 ( .A1(n1132), .A2(n1008), .ZN(n1108) );
XOR2_X1 U845 ( .A(n1133), .B(KEYINPUT14), .Z(n1132) );
XNOR2_X1 U846 ( .A(G116), .B(n1134), .ZN(G18) );
NOR2_X1 U847 ( .A1(n1104), .A2(KEYINPUT15), .ZN(n1134) );
AND3_X1 U848 ( .A1(n1130), .A2(n971), .A3(n990), .ZN(n1104) );
NOR2_X1 U849 ( .A1(n1111), .A2(n1135), .ZN(n971) );
NAND2_X1 U850 ( .A1(n1136), .A2(n1137), .ZN(G15) );
NAND2_X1 U851 ( .A1(n1103), .A2(n1138), .ZN(n1137) );
XOR2_X1 U852 ( .A(KEYINPUT4), .B(n1139), .Z(n1136) );
NOR2_X1 U853 ( .A1(n1103), .A2(n1138), .ZN(n1139) );
AND3_X1 U854 ( .A1(n975), .A2(n1130), .A3(n990), .ZN(n1103) );
NOR2_X1 U855 ( .A1(n1008), .A2(n1133), .ZN(n990) );
NOR3_X1 U856 ( .A1(n1095), .A2(n1140), .A3(n973), .ZN(n1130) );
INV_X1 U857 ( .A(n969), .ZN(n973) );
NOR2_X1 U858 ( .A1(n981), .A2(n997), .ZN(n969) );
INV_X1 U859 ( .A(n982), .ZN(n997) );
INV_X1 U860 ( .A(n1098), .ZN(n975) );
NAND2_X1 U861 ( .A1(n1141), .A2(n1111), .ZN(n1098) );
XOR2_X1 U862 ( .A(n1135), .B(KEYINPUT11), .Z(n1141) );
XOR2_X1 U863 ( .A(n1142), .B(n1143), .Z(G12) );
NOR2_X1 U864 ( .A1(KEYINPUT62), .A2(n1144), .ZN(n1143) );
NAND2_X1 U865 ( .A1(n1145), .A2(n1146), .ZN(n1142) );
OR2_X1 U866 ( .A1(n1100), .A2(KEYINPUT58), .ZN(n1146) );
NAND3_X1 U867 ( .A1(n989), .A2(n1105), .A3(n991), .ZN(n1100) );
AND2_X1 U868 ( .A1(n1123), .A2(n1147), .ZN(n1105) );
NOR2_X1 U869 ( .A1(n1095), .A2(n980), .ZN(n1123) );
NAND4_X1 U870 ( .A1(n991), .A2(n989), .A3(n1148), .A4(KEYINPUT58), .ZN(n1145) );
NOR3_X1 U871 ( .A1(n980), .A2(n1140), .A3(n985), .ZN(n1148) );
INV_X1 U872 ( .A(n1095), .ZN(n985) );
NAND2_X1 U873 ( .A1(n986), .A2(n987), .ZN(n1095) );
NAND2_X1 U874 ( .A1(G214), .A2(n1149), .ZN(n987) );
INV_X1 U875 ( .A(n1007), .ZN(n986) );
XNOR2_X1 U876 ( .A(n1150), .B(n1082), .ZN(n1007) );
NAND2_X1 U877 ( .A1(G210), .A2(n1149), .ZN(n1082) );
NAND2_X1 U878 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
XOR2_X1 U879 ( .A(n1153), .B(KEYINPUT40), .Z(n1151) );
NAND2_X1 U880 ( .A1(n1154), .A2(n1152), .ZN(n1150) );
XOR2_X1 U881 ( .A(KEYINPUT17), .B(n1155), .Z(n1154) );
INV_X1 U882 ( .A(n1107), .ZN(n1155) );
XOR2_X1 U883 ( .A(n1156), .B(n1157), .Z(n1107) );
XOR2_X1 U884 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U885 ( .A(KEYINPUT25), .B(G125), .Z(n1159) );
NOR2_X1 U886 ( .A1(n1160), .A2(n1038), .ZN(n1158) );
INV_X1 U887 ( .A(G224), .ZN(n1038) );
XNOR2_X1 U888 ( .A(n1034), .B(n1023), .ZN(n1156) );
XNOR2_X1 U889 ( .A(n1161), .B(n1162), .ZN(n1034) );
XOR2_X1 U890 ( .A(G113), .B(n1163), .Z(n1162) );
XOR2_X1 U891 ( .A(KEYINPUT16), .B(G119), .Z(n1163) );
XOR2_X1 U892 ( .A(n1073), .B(n1164), .Z(n1161) );
XNOR2_X1 U893 ( .A(n1165), .B(n1166), .ZN(n1164) );
NAND2_X1 U894 ( .A1(KEYINPUT36), .A2(n1124), .ZN(n1165) );
INV_X1 U895 ( .A(G101), .ZN(n1124) );
XOR2_X1 U896 ( .A(n1144), .B(n1167), .Z(n1073) );
INV_X1 U897 ( .A(n1147), .ZN(n1140) );
NAND2_X1 U898 ( .A1(n956), .A2(n1168), .ZN(n1147) );
NAND3_X1 U899 ( .A1(G902), .A2(n1128), .A3(n1032), .ZN(n1168) );
NOR2_X1 U900 ( .A1(G898), .A2(n1029), .ZN(n1032) );
NAND3_X1 U901 ( .A1(n1128), .A2(n1029), .A3(G952), .ZN(n956) );
NAND2_X1 U902 ( .A1(G234), .A2(G237), .ZN(n1128) );
NAND2_X1 U903 ( .A1(n981), .A2(n982), .ZN(n980) );
NAND2_X1 U904 ( .A1(G221), .A2(n1169), .ZN(n982) );
NAND3_X1 U905 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n981) );
NAND2_X1 U906 ( .A1(G469), .A2(n1006), .ZN(n1172) );
NAND2_X1 U907 ( .A1(KEYINPUT35), .A2(n1173), .ZN(n1171) );
NAND2_X1 U908 ( .A1(n1174), .A2(n1005), .ZN(n1173) );
INV_X1 U909 ( .A(G469), .ZN(n1005) );
XOR2_X1 U910 ( .A(n1006), .B(KEYINPUT61), .Z(n1174) );
NAND2_X1 U911 ( .A1(n1175), .A2(n1176), .ZN(n1170) );
INV_X1 U912 ( .A(KEYINPUT35), .ZN(n1176) );
NAND2_X1 U913 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
NAND2_X1 U914 ( .A1(n1006), .A2(n1179), .ZN(n1178) );
OR3_X1 U915 ( .A1(n1006), .A2(G469), .A3(n1179), .ZN(n1177) );
INV_X1 U916 ( .A(KEYINPUT61), .ZN(n1179) );
NAND2_X1 U917 ( .A1(n1180), .A2(n1152), .ZN(n1006) );
XOR2_X1 U918 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U919 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U920 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NOR2_X1 U921 ( .A1(KEYINPUT49), .A2(n1187), .ZN(n1186) );
AND2_X1 U922 ( .A1(KEYINPUT26), .A2(n1187), .ZN(n1185) );
XNOR2_X1 U923 ( .A(n1188), .B(n1189), .ZN(n1187) );
XNOR2_X1 U924 ( .A(KEYINPUT43), .B(n1167), .ZN(n1188) );
XNOR2_X1 U925 ( .A(G104), .B(n1190), .ZN(n1167) );
XOR2_X1 U926 ( .A(n1191), .B(n1192), .Z(n1183) );
NOR2_X1 U927 ( .A1(KEYINPUT0), .A2(n1193), .ZN(n1192) );
XOR2_X1 U928 ( .A(n1112), .B(KEYINPUT56), .Z(n1193) );
INV_X1 U929 ( .A(G140), .ZN(n1112) );
XOR2_X1 U930 ( .A(n1194), .B(n1071), .Z(n1181) );
AND2_X1 U931 ( .A1(G227), .A2(n1195), .ZN(n1071) );
XOR2_X1 U932 ( .A(n1144), .B(KEYINPUT31), .Z(n1194) );
INV_X1 U933 ( .A(G110), .ZN(n1144) );
NOR2_X1 U934 ( .A1(n999), .A2(n1111), .ZN(n989) );
NAND2_X1 U935 ( .A1(n1196), .A2(n1197), .ZN(n1111) );
NAND2_X1 U936 ( .A1(G475), .A2(n1004), .ZN(n1197) );
XOR2_X1 U937 ( .A(KEYINPUT3), .B(n1198), .Z(n1196) );
NOR2_X1 U938 ( .A1(n1199), .A2(n1004), .ZN(n1198) );
OR2_X1 U939 ( .A1(n1059), .A2(G902), .ZN(n1004) );
XNOR2_X1 U940 ( .A(n1200), .B(n1201), .ZN(n1059) );
XOR2_X1 U941 ( .A(G104), .B(n1202), .Z(n1201) );
NOR2_X1 U942 ( .A1(KEYINPUT37), .A2(G113), .ZN(n1202) );
XOR2_X1 U943 ( .A(n1203), .B(n1204), .Z(n1200) );
NOR3_X1 U944 ( .A1(n1205), .A2(n1206), .A3(n1160), .ZN(n1204) );
INV_X1 U945 ( .A(n1195), .ZN(n1160) );
XOR2_X1 U946 ( .A(n1153), .B(KEYINPUT33), .Z(n1206) );
INV_X1 U947 ( .A(G214), .ZN(n1205) );
XOR2_X1 U948 ( .A(n1207), .B(n1208), .Z(n1203) );
XOR2_X1 U949 ( .A(n1209), .B(n1210), .Z(n1208) );
XNOR2_X1 U950 ( .A(G122), .B(n1211), .ZN(n1210) );
NOR2_X1 U951 ( .A1(G140), .A2(KEYINPUT53), .ZN(n1211) );
XOR2_X1 U952 ( .A(n1212), .B(n1213), .Z(n1207) );
XOR2_X1 U953 ( .A(KEYINPUT46), .B(G131), .Z(n1213) );
XNOR2_X1 U954 ( .A(G475), .B(KEYINPUT10), .ZN(n1199) );
INV_X1 U955 ( .A(n1135), .ZN(n999) );
XOR2_X1 U956 ( .A(n1214), .B(G478), .Z(n1135) );
NAND2_X1 U957 ( .A1(n1215), .A2(n1055), .ZN(n1214) );
XOR2_X1 U958 ( .A(n1216), .B(n1217), .Z(n1055) );
AND3_X1 U959 ( .A1(G234), .A2(G217), .A3(n1195), .ZN(n1217) );
NAND2_X1 U960 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
NAND2_X1 U961 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
INV_X1 U962 ( .A(n1222), .ZN(n1221) );
XOR2_X1 U963 ( .A(n1190), .B(n1166), .Z(n1220) );
INV_X1 U964 ( .A(G107), .ZN(n1190) );
XOR2_X1 U965 ( .A(n1223), .B(KEYINPUT8), .Z(n1218) );
NAND2_X1 U966 ( .A1(n1222), .A2(n1224), .ZN(n1223) );
XOR2_X1 U967 ( .A(G107), .B(n1166), .Z(n1224) );
XOR2_X1 U968 ( .A(G116), .B(G122), .Z(n1166) );
XOR2_X1 U969 ( .A(n1225), .B(n1226), .Z(n1222) );
XOR2_X1 U970 ( .A(G134), .B(n1227), .Z(n1226) );
NOR2_X1 U971 ( .A1(G128), .A2(KEYINPUT39), .ZN(n1227) );
XNOR2_X1 U972 ( .A(G143), .B(KEYINPUT55), .ZN(n1225) );
XOR2_X1 U973 ( .A(n1152), .B(KEYINPUT63), .Z(n1215) );
AND2_X1 U974 ( .A1(n1228), .A2(n1008), .ZN(n991) );
XOR2_X1 U975 ( .A(n1229), .B(n1049), .Z(n1008) );
NAND2_X1 U976 ( .A1(G217), .A2(n1169), .ZN(n1049) );
NAND2_X1 U977 ( .A1(G234), .A2(n1152), .ZN(n1169) );
OR2_X1 U978 ( .A1(n1048), .A2(G902), .ZN(n1229) );
XNOR2_X1 U979 ( .A(n1230), .B(n1231), .ZN(n1048) );
XOR2_X1 U980 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U981 ( .A(G146), .B(G110), .Z(n1233) );
NOR2_X1 U982 ( .A1(KEYINPUT28), .A2(n1234), .ZN(n1232) );
XOR2_X1 U983 ( .A(n1115), .B(n1235), .Z(n1234) );
AND3_X1 U984 ( .A1(G221), .A2(G234), .A3(n1195), .ZN(n1235) );
INV_X1 U985 ( .A(G137), .ZN(n1115) );
XNOR2_X1 U986 ( .A(n1236), .B(n1237), .ZN(n1230) );
NAND2_X1 U987 ( .A1(KEYINPUT29), .A2(n1015), .ZN(n1237) );
XOR2_X1 U988 ( .A(n1212), .B(G140), .Z(n1015) );
INV_X1 U989 ( .A(G125), .ZN(n1212) );
NAND2_X1 U990 ( .A1(KEYINPUT59), .A2(n1238), .ZN(n1236) );
XOR2_X1 U991 ( .A(G128), .B(G119), .Z(n1238) );
XOR2_X1 U992 ( .A(KEYINPUT19), .B(n1131), .Z(n1228) );
INV_X1 U993 ( .A(n1133), .ZN(n1131) );
XOR2_X1 U994 ( .A(n1000), .B(G472), .Z(n1133) );
NAND2_X1 U995 ( .A1(n1239), .A2(n1152), .ZN(n1000) );
INV_X1 U996 ( .A(G902), .ZN(n1152) );
XOR2_X1 U997 ( .A(KEYINPUT9), .B(n1240), .Z(n1239) );
INV_X1 U998 ( .A(n1062), .ZN(n1240) );
XOR2_X1 U999 ( .A(n1241), .B(n1242), .Z(n1062) );
XOR2_X1 U1000 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U1001 ( .A(KEYINPUT60), .B(KEYINPUT25), .Z(n1244) );
NOR2_X1 U1002 ( .A1(n1245), .A2(n1246), .ZN(n1243) );
XOR2_X1 U1003 ( .A(n1247), .B(KEYINPUT13), .Z(n1246) );
NAND2_X1 U1004 ( .A1(n1248), .A2(n1138), .ZN(n1247) );
NOR2_X1 U1005 ( .A1(n1248), .A2(n1138), .ZN(n1245) );
INV_X1 U1006 ( .A(G113), .ZN(n1138) );
XNOR2_X1 U1007 ( .A(G116), .B(n1249), .ZN(n1248) );
XOR2_X1 U1008 ( .A(KEYINPUT5), .B(G119), .Z(n1249) );
XOR2_X1 U1009 ( .A(n1250), .B(n1074), .Z(n1241) );
XOR2_X1 U1010 ( .A(n1021), .B(n1189), .Z(n1074) );
XOR2_X1 U1011 ( .A(G101), .B(n1023), .Z(n1189) );
XOR2_X1 U1012 ( .A(n1251), .B(n1209), .Z(n1023) );
XNOR2_X1 U1013 ( .A(G143), .B(G146), .ZN(n1209) );
INV_X1 U1014 ( .A(G128), .ZN(n1251) );
INV_X1 U1015 ( .A(n1191), .ZN(n1021) );
XNOR2_X1 U1016 ( .A(G131), .B(n1252), .ZN(n1191) );
XOR2_X1 U1017 ( .A(G137), .B(G134), .Z(n1252) );
NAND3_X1 U1018 ( .A1(n1195), .A2(n1153), .A3(G210), .ZN(n1250) );
INV_X1 U1019 ( .A(G237), .ZN(n1153) );
XOR2_X1 U1020 ( .A(n1029), .B(KEYINPUT41), .Z(n1195) );
INV_X1 U1021 ( .A(G953), .ZN(n1029) );
endmodule


