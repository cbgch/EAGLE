//Key = 1111110101110101011001011100101111101111010011101101011001110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284;

XNOR2_X1 U716 ( .A(G107), .B(n978), .ZN(G9) );
NOR2_X1 U717 ( .A1(n979), .A2(n980), .ZN(G75) );
NOR4_X1 U718 ( .A1(G953), .A2(n981), .A3(n982), .A4(n983), .ZN(n980) );
NOR2_X1 U719 ( .A1(n984), .A2(n985), .ZN(n982) );
NOR2_X1 U720 ( .A1(n986), .A2(n987), .ZN(n985) );
NOR3_X1 U721 ( .A1(n988), .A2(n989), .A3(n990), .ZN(n987) );
NOR2_X1 U722 ( .A1(n991), .A2(n992), .ZN(n989) );
AND2_X1 U723 ( .A1(n993), .A2(n994), .ZN(n992) );
NOR3_X1 U724 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n991) );
NOR2_X1 U725 ( .A1(n998), .A2(n999), .ZN(n997) );
XNOR2_X1 U726 ( .A(n994), .B(KEYINPUT18), .ZN(n999) );
NOR3_X1 U727 ( .A1(n1000), .A2(n1001), .A3(n1002), .ZN(n996) );
NOR2_X1 U728 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NOR4_X1 U729 ( .A1(n1005), .A2(n1000), .A3(n1006), .A4(n995), .ZN(n986) );
NOR3_X1 U730 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1005) );
AND3_X1 U731 ( .A1(n988), .A2(n1010), .A3(KEYINPUT60), .ZN(n1009) );
NOR2_X1 U732 ( .A1(n1011), .A2(n988), .ZN(n1008) );
INV_X1 U733 ( .A(n1012), .ZN(n988) );
NOR2_X1 U734 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
NOR2_X1 U735 ( .A1(KEYINPUT60), .A2(n1015), .ZN(n1013) );
NOR2_X1 U736 ( .A1(n1016), .A2(n990), .ZN(n1007) );
NOR2_X1 U737 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
INV_X1 U738 ( .A(n1019), .ZN(n984) );
NOR3_X1 U739 ( .A1(n981), .A2(G953), .A3(G952), .ZN(n979) );
AND4_X1 U740 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n981) );
NOR3_X1 U741 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
NAND3_X1 U742 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1024) );
XNOR2_X1 U743 ( .A(n1030), .B(n1031), .ZN(n1029) );
OR2_X1 U744 ( .A1(G478), .A2(KEYINPUT25), .ZN(n1028) );
NAND2_X1 U745 ( .A1(KEYINPUT25), .A2(n1032), .ZN(n1027) );
AND3_X1 U746 ( .A1(n998), .A2(n1033), .A3(n1003), .ZN(n1022) );
XOR2_X1 U747 ( .A(n1034), .B(n1035), .Z(n1021) );
NAND2_X1 U748 ( .A1(KEYINPUT13), .A2(n1036), .ZN(n1035) );
XOR2_X1 U749 ( .A(n1037), .B(n1038), .Z(n1020) );
XNOR2_X1 U750 ( .A(n1039), .B(KEYINPUT24), .ZN(n1038) );
XOR2_X1 U751 ( .A(n1040), .B(n1041), .Z(G72) );
NOR2_X1 U752 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NAND2_X1 U754 ( .A1(n1046), .A2(n1047), .ZN(n1040) );
NAND2_X1 U755 ( .A1(n1048), .A2(n1043), .ZN(n1047) );
XNOR2_X1 U756 ( .A(n1049), .B(n1050), .ZN(n1048) );
NAND3_X1 U757 ( .A1(G900), .A2(n1050), .A3(G953), .ZN(n1046) );
XOR2_X1 U758 ( .A(n1051), .B(n1052), .Z(n1050) );
XOR2_X1 U759 ( .A(n1053), .B(n1054), .Z(n1052) );
XNOR2_X1 U760 ( .A(G131), .B(G134), .ZN(n1054) );
NAND2_X1 U761 ( .A1(KEYINPUT39), .A2(n1055), .ZN(n1053) );
XOR2_X1 U762 ( .A(n1056), .B(n1057), .Z(n1051) );
NAND3_X1 U763 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1056) );
NAND2_X1 U764 ( .A1(G125), .A2(n1061), .ZN(n1060) );
OR3_X1 U765 ( .A1(n1061), .A2(n1062), .A3(G140), .ZN(n1059) );
INV_X1 U766 ( .A(KEYINPUT45), .ZN(n1061) );
NAND2_X1 U767 ( .A1(G140), .A2(n1062), .ZN(n1058) );
NAND2_X1 U768 ( .A1(KEYINPUT9), .A2(n1063), .ZN(n1062) );
XOR2_X1 U769 ( .A(n1064), .B(n1065), .Z(G69) );
XOR2_X1 U770 ( .A(n1066), .B(n1067), .Z(n1065) );
NOR2_X1 U771 ( .A1(n1068), .A2(n1043), .ZN(n1067) );
NOR2_X1 U772 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U773 ( .A1(n1071), .A2(n1072), .ZN(n1066) );
NAND2_X1 U774 ( .A1(n1073), .A2(n1070), .ZN(n1072) );
XNOR2_X1 U775 ( .A(KEYINPUT27), .B(n1043), .ZN(n1073) );
XOR2_X1 U776 ( .A(n1074), .B(n1075), .Z(n1071) );
XNOR2_X1 U777 ( .A(n1076), .B(KEYINPUT23), .ZN(n1075) );
NAND2_X1 U778 ( .A1(n1077), .A2(KEYINPUT11), .ZN(n1076) );
XOR2_X1 U779 ( .A(n1078), .B(n1079), .Z(n1077) );
XOR2_X1 U780 ( .A(n1080), .B(n1081), .Z(n1078) );
NAND2_X1 U781 ( .A1(n1043), .A2(n1082), .ZN(n1064) );
NAND2_X1 U782 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XNOR2_X1 U783 ( .A(KEYINPUT51), .B(n978), .ZN(n1084) );
NOR2_X1 U784 ( .A1(n1085), .A2(n1086), .ZN(G66) );
NOR3_X1 U785 ( .A1(n1039), .A2(n1087), .A3(n1088), .ZN(n1086) );
NOR4_X1 U786 ( .A1(n1089), .A2(n1090), .A3(n1037), .A4(n1091), .ZN(n1088) );
INV_X1 U787 ( .A(n1092), .ZN(n1089) );
NOR2_X1 U788 ( .A1(n1093), .A2(n1092), .ZN(n1087) );
NOR3_X1 U789 ( .A1(n1090), .A2(n1094), .A3(n1037), .ZN(n1093) );
INV_X1 U790 ( .A(KEYINPUT36), .ZN(n1090) );
NOR2_X1 U791 ( .A1(n1085), .A2(n1095), .ZN(G63) );
XNOR2_X1 U792 ( .A(n1096), .B(n1097), .ZN(n1095) );
XOR2_X1 U793 ( .A(KEYINPUT61), .B(n1098), .Z(n1097) );
NOR2_X1 U794 ( .A1(n1099), .A2(n1091), .ZN(n1098) );
NOR2_X1 U795 ( .A1(n1085), .A2(n1100), .ZN(G60) );
XOR2_X1 U796 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U797 ( .A1(n1103), .A2(n1091), .ZN(n1101) );
XNOR2_X1 U798 ( .A(G104), .B(n1104), .ZN(G6) );
NOR2_X1 U799 ( .A1(n1105), .A2(n1106), .ZN(G57) );
XOR2_X1 U800 ( .A(n1107), .B(n1108), .Z(n1106) );
XNOR2_X1 U801 ( .A(KEYINPUT41), .B(n1109), .ZN(n1108) );
NOR4_X1 U802 ( .A1(KEYINPUT50), .A2(n1094), .A3(n1031), .A4(n1110), .ZN(n1109) );
XNOR2_X1 U803 ( .A(KEYINPUT59), .B(n1111), .ZN(n1110) );
INV_X1 U804 ( .A(G472), .ZN(n1031) );
NOR2_X1 U805 ( .A1(n1043), .A2(n1112), .ZN(n1105) );
XNOR2_X1 U806 ( .A(KEYINPUT55), .B(n1113), .ZN(n1112) );
NOR2_X1 U807 ( .A1(n1085), .A2(n1114), .ZN(G54) );
XOR2_X1 U808 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U809 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U810 ( .A(n1119), .B(n1120), .Z(n1118) );
NOR3_X1 U811 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1120) );
NOR2_X1 U812 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
AND3_X1 U813 ( .A1(n1125), .A2(n1126), .A3(n1124), .ZN(n1122) );
AND2_X1 U814 ( .A1(KEYINPUT34), .A2(n1127), .ZN(n1124) );
NOR2_X1 U815 ( .A1(n1127), .A2(n1126), .ZN(n1121) );
INV_X1 U816 ( .A(KEYINPUT63), .ZN(n1126) );
XOR2_X1 U817 ( .A(n1128), .B(KEYINPUT21), .Z(n1127) );
NOR2_X1 U818 ( .A1(G110), .A2(KEYINPUT52), .ZN(n1119) );
NOR2_X1 U819 ( .A1(n1129), .A2(n1091), .ZN(n1117) );
NAND2_X1 U820 ( .A1(G902), .A2(n983), .ZN(n1091) );
XOR2_X1 U821 ( .A(n1130), .B(n1131), .Z(n1115) );
XOR2_X1 U822 ( .A(KEYINPUT38), .B(G140), .Z(n1131) );
NOR2_X1 U823 ( .A1(n1085), .A2(n1132), .ZN(G51) );
XOR2_X1 U824 ( .A(n1133), .B(n1134), .Z(n1132) );
XNOR2_X1 U825 ( .A(n1135), .B(n1136), .ZN(n1134) );
NOR3_X1 U826 ( .A1(KEYINPUT35), .A2(n1137), .A3(n1138), .ZN(n1136) );
AND3_X1 U827 ( .A1(KEYINPUT19), .A2(n1063), .A3(n1139), .ZN(n1138) );
NOR2_X1 U828 ( .A1(KEYINPUT19), .A2(n1140), .ZN(n1137) );
NAND4_X1 U829 ( .A1(n1141), .A2(KEYINPUT15), .A3(G902), .A4(n1142), .ZN(n1135) );
INV_X1 U830 ( .A(n1036), .ZN(n1142) );
XNOR2_X1 U831 ( .A(n1094), .B(KEYINPUT26), .ZN(n1141) );
INV_X1 U832 ( .A(n983), .ZN(n1094) );
NAND3_X1 U833 ( .A1(n1083), .A2(n978), .A3(n1049), .ZN(n983) );
AND4_X1 U834 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1049) );
NOR4_X1 U835 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1146) );
NOR2_X1 U836 ( .A1(n1151), .A2(n1152), .ZN(n1145) );
NOR2_X1 U837 ( .A1(n1006), .A2(n1153), .ZN(n1152) );
XOR2_X1 U838 ( .A(KEYINPUT46), .B(n1154), .Z(n1153) );
INV_X1 U839 ( .A(n994), .ZN(n1006) );
INV_X1 U840 ( .A(n1155), .ZN(n1151) );
NAND3_X1 U841 ( .A1(n1156), .A2(n1157), .A3(n1017), .ZN(n978) );
AND4_X1 U842 ( .A1(n1104), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1083) );
AND4_X1 U843 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1160) );
NAND3_X1 U844 ( .A1(n1018), .A2(n1014), .A3(n1165), .ZN(n1159) );
NAND3_X1 U845 ( .A1(n1156), .A2(n1157), .A3(n1018), .ZN(n1104) );
NOR2_X1 U846 ( .A1(n1043), .A2(G952), .ZN(n1085) );
XOR2_X1 U847 ( .A(G146), .B(n1150), .Z(G48) );
AND3_X1 U848 ( .A1(n1166), .A2(n1001), .A3(n1018), .ZN(n1150) );
XNOR2_X1 U849 ( .A(n1167), .B(n1168), .ZN(G45) );
NAND2_X1 U850 ( .A1(KEYINPUT4), .A2(n1155), .ZN(n1167) );
NAND4_X1 U851 ( .A1(n1169), .A2(n993), .A3(n1014), .A4(n1170), .ZN(n1155) );
AND3_X1 U852 ( .A1(n1001), .A2(n1171), .A3(n1026), .ZN(n1170) );
XNOR2_X1 U853 ( .A(G140), .B(n1143), .ZN(G42) );
NAND3_X1 U854 ( .A1(n994), .A2(n993), .A3(n1172), .ZN(n1143) );
XNOR2_X1 U855 ( .A(G137), .B(n1173), .ZN(G39) );
NAND2_X1 U856 ( .A1(n1154), .A2(n994), .ZN(n1173) );
AND2_X1 U857 ( .A1(n1012), .A2(n1166), .ZN(n1154) );
XOR2_X1 U858 ( .A(G134), .B(n1149), .Z(G36) );
AND2_X1 U859 ( .A1(n1174), .A2(n1017), .ZN(n1149) );
XNOR2_X1 U860 ( .A(n1175), .B(n1148), .ZN(G33) );
AND2_X1 U861 ( .A1(n1174), .A2(n1018), .ZN(n1148) );
AND4_X1 U862 ( .A1(n1014), .A2(n994), .A3(n1169), .A4(n993), .ZN(n1174) );
NOR2_X1 U863 ( .A1(n1004), .A2(n1176), .ZN(n994) );
XOR2_X1 U864 ( .A(G128), .B(n1147), .Z(G30) );
AND3_X1 U865 ( .A1(n1017), .A2(n1001), .A3(n1166), .ZN(n1147) );
AND4_X1 U866 ( .A1(n1177), .A2(n1169), .A3(n993), .A4(n1178), .ZN(n1166) );
XNOR2_X1 U867 ( .A(G101), .B(n1158), .ZN(G3) );
NAND3_X1 U868 ( .A1(n1014), .A2(n1157), .A3(n1012), .ZN(n1158) );
XNOR2_X1 U869 ( .A(G125), .B(n1144), .ZN(G27) );
NAND4_X1 U870 ( .A1(n1179), .A2(n1172), .A3(n1001), .A4(n998), .ZN(n1144) );
AND3_X1 U871 ( .A1(n1018), .A2(n1169), .A3(n1010), .ZN(n1172) );
AND3_X1 U872 ( .A1(n1180), .A2(n1181), .A3(n1019), .ZN(n1169) );
NAND2_X1 U873 ( .A1(G953), .A2(n1182), .ZN(n1180) );
NAND2_X1 U874 ( .A1(G902), .A2(n1045), .ZN(n1182) );
INV_X1 U875 ( .A(G900), .ZN(n1045) );
XNOR2_X1 U876 ( .A(G122), .B(n1163), .ZN(G24) );
NAND4_X1 U877 ( .A1(n1165), .A2(n1156), .A3(n1026), .A4(n1171), .ZN(n1163) );
INV_X1 U878 ( .A(n990), .ZN(n1156) );
NAND2_X1 U879 ( .A1(n1183), .A2(n1184), .ZN(n990) );
XNOR2_X1 U880 ( .A(G119), .B(n1164), .ZN(G21) );
NAND4_X1 U881 ( .A1(n1165), .A2(n1012), .A3(n1177), .A4(n1178), .ZN(n1164) );
XNOR2_X1 U882 ( .A(G116), .B(n1162), .ZN(G18) );
NAND3_X1 U883 ( .A1(n1014), .A2(n1017), .A3(n1165), .ZN(n1162) );
AND2_X1 U884 ( .A1(n1185), .A2(n1171), .ZN(n1017) );
XNOR2_X1 U885 ( .A(G113), .B(n1186), .ZN(G15) );
NAND3_X1 U886 ( .A1(n1165), .A2(n1018), .A3(n1187), .ZN(n1186) );
XNOR2_X1 U887 ( .A(n1014), .B(KEYINPUT7), .ZN(n1187) );
AND2_X1 U888 ( .A1(n1184), .A2(n1178), .ZN(n1014) );
NOR2_X1 U889 ( .A1(n1171), .A2(n1185), .ZN(n1018) );
INV_X1 U890 ( .A(n1026), .ZN(n1185) );
AND3_X1 U891 ( .A1(n1188), .A2(n998), .A3(n1179), .ZN(n1165) );
XNOR2_X1 U892 ( .A(G110), .B(n1161), .ZN(G12) );
NAND3_X1 U893 ( .A1(n1010), .A2(n1157), .A3(n1012), .ZN(n1161) );
NOR2_X1 U894 ( .A1(n1171), .A2(n1026), .ZN(n1012) );
XOR2_X1 U895 ( .A(n1189), .B(n1103), .Z(n1026) );
INV_X1 U896 ( .A(G475), .ZN(n1103) );
OR2_X1 U897 ( .A1(n1102), .A2(G902), .ZN(n1189) );
XNOR2_X1 U898 ( .A(n1190), .B(n1191), .ZN(n1102) );
XOR2_X1 U899 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U900 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U901 ( .A(n1196), .B(n1197), .Z(n1195) );
NAND2_X1 U902 ( .A1(KEYINPUT1), .A2(n1063), .ZN(n1197) );
NAND2_X1 U903 ( .A1(G214), .A2(n1198), .ZN(n1196) );
XNOR2_X1 U904 ( .A(n1199), .B(n1200), .ZN(n1194) );
NOR2_X1 U905 ( .A1(G146), .A2(KEYINPUT42), .ZN(n1200) );
XOR2_X1 U906 ( .A(n1201), .B(n1202), .Z(n1192) );
XOR2_X1 U907 ( .A(KEYINPUT20), .B(G140), .Z(n1202) );
XNOR2_X1 U908 ( .A(G104), .B(G122), .ZN(n1201) );
XNOR2_X1 U909 ( .A(G143), .B(KEYINPUT30), .ZN(n1190) );
NAND3_X1 U910 ( .A1(n1203), .A2(n1204), .A3(n1033), .ZN(n1171) );
NAND3_X1 U911 ( .A1(n1099), .A2(n1111), .A3(n1096), .ZN(n1033) );
INV_X1 U912 ( .A(G478), .ZN(n1099) );
OR2_X1 U913 ( .A1(G478), .A2(KEYINPUT57), .ZN(n1204) );
NAND2_X1 U914 ( .A1(n1032), .A2(KEYINPUT57), .ZN(n1203) );
AND2_X1 U915 ( .A1(G478), .A2(n1205), .ZN(n1032) );
NAND2_X1 U916 ( .A1(n1096), .A2(n1111), .ZN(n1205) );
XOR2_X1 U917 ( .A(n1206), .B(n1207), .Z(n1096) );
XOR2_X1 U918 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U919 ( .A(G128), .B(n1210), .Z(n1209) );
NOR2_X1 U920 ( .A1(KEYINPUT16), .A2(n1211), .ZN(n1210) );
XNOR2_X1 U921 ( .A(n1212), .B(n1213), .ZN(n1211) );
XOR2_X1 U922 ( .A(G122), .B(G116), .Z(n1213) );
AND2_X1 U923 ( .A1(n1214), .A2(G217), .ZN(n1208) );
XNOR2_X1 U924 ( .A(G134), .B(n1215), .ZN(n1206) );
XNOR2_X1 U925 ( .A(KEYINPUT22), .B(n1168), .ZN(n1215) );
AND2_X1 U926 ( .A1(n1188), .A2(n993), .ZN(n1157) );
NOR2_X1 U927 ( .A1(n1179), .A2(n1000), .ZN(n993) );
INV_X1 U928 ( .A(n998), .ZN(n1000) );
NAND2_X1 U929 ( .A1(G221), .A2(n1216), .ZN(n998) );
INV_X1 U930 ( .A(n995), .ZN(n1179) );
XOR2_X1 U931 ( .A(n1025), .B(KEYINPUT14), .Z(n995) );
XOR2_X1 U932 ( .A(n1217), .B(n1129), .Z(n1025) );
INV_X1 U933 ( .A(G469), .ZN(n1129) );
NAND2_X1 U934 ( .A1(n1218), .A2(n1111), .ZN(n1217) );
XOR2_X1 U935 ( .A(n1219), .B(n1220), .Z(n1218) );
XOR2_X1 U936 ( .A(n1221), .B(n1222), .Z(n1220) );
XOR2_X1 U937 ( .A(G140), .B(n1130), .Z(n1222) );
NOR2_X1 U938 ( .A1(n1044), .A2(G953), .ZN(n1130) );
INV_X1 U939 ( .A(G227), .ZN(n1044) );
NOR2_X1 U940 ( .A1(G110), .A2(KEYINPUT29), .ZN(n1221) );
XNOR2_X1 U941 ( .A(n1125), .B(n1128), .ZN(n1219) );
XOR2_X1 U942 ( .A(n1223), .B(n1175), .Z(n1128) );
INV_X1 U943 ( .A(G131), .ZN(n1175) );
XNOR2_X1 U944 ( .A(n1224), .B(n1225), .ZN(n1125) );
XOR2_X1 U945 ( .A(n1226), .B(n1057), .Z(n1225) );
XNOR2_X1 U946 ( .A(n1227), .B(n1228), .ZN(n1057) );
XOR2_X1 U947 ( .A(n1229), .B(KEYINPUT48), .Z(n1227) );
NAND2_X1 U948 ( .A1(KEYINPUT53), .A2(G128), .ZN(n1229) );
NOR2_X1 U949 ( .A1(KEYINPUT40), .A2(n1230), .ZN(n1226) );
XNOR2_X1 U950 ( .A(n1231), .B(n1232), .ZN(n1224) );
INV_X1 U951 ( .A(G104), .ZN(n1232) );
NAND2_X1 U952 ( .A1(KEYINPUT33), .A2(G107), .ZN(n1231) );
AND4_X1 U953 ( .A1(n1001), .A2(n1019), .A3(n1233), .A4(n1181), .ZN(n1188) );
NAND2_X1 U954 ( .A1(n1113), .A2(n1043), .ZN(n1181) );
INV_X1 U955 ( .A(G952), .ZN(n1113) );
NAND2_X1 U956 ( .A1(G953), .A2(n1234), .ZN(n1233) );
NAND2_X1 U957 ( .A1(G902), .A2(n1070), .ZN(n1234) );
INV_X1 U958 ( .A(G898), .ZN(n1070) );
NAND2_X1 U959 ( .A1(n1235), .A2(G234), .ZN(n1019) );
XNOR2_X1 U960 ( .A(G237), .B(KEYINPUT10), .ZN(n1235) );
NOR2_X1 U961 ( .A1(n1176), .A2(n1236), .ZN(n1001) );
INV_X1 U962 ( .A(n1004), .ZN(n1236) );
XOR2_X1 U963 ( .A(n1034), .B(n1036), .Z(n1004) );
NAND2_X1 U964 ( .A1(G210), .A2(n1237), .ZN(n1036) );
NAND2_X1 U965 ( .A1(n1238), .A2(n1111), .ZN(n1034) );
XNOR2_X1 U966 ( .A(n1133), .B(n1140), .ZN(n1238) );
XNOR2_X1 U967 ( .A(n1139), .B(n1063), .ZN(n1140) );
INV_X1 U968 ( .A(G125), .ZN(n1063) );
XOR2_X1 U969 ( .A(n1239), .B(n1240), .Z(n1133) );
XOR2_X1 U970 ( .A(n1241), .B(n1074), .Z(n1240) );
XNOR2_X1 U971 ( .A(n1242), .B(n1243), .ZN(n1074) );
XOR2_X1 U972 ( .A(KEYINPUT5), .B(G122), .Z(n1243) );
INV_X1 U973 ( .A(G110), .ZN(n1242) );
NOR2_X1 U974 ( .A1(G953), .A2(n1069), .ZN(n1241) );
INV_X1 U975 ( .A(G224), .ZN(n1069) );
XNOR2_X1 U976 ( .A(KEYINPUT12), .B(n1244), .ZN(n1239) );
NOR2_X1 U977 ( .A1(KEYINPUT8), .A2(n1245), .ZN(n1244) );
XOR2_X1 U978 ( .A(n1080), .B(n1246), .Z(n1245) );
XNOR2_X1 U979 ( .A(n1247), .B(n1230), .ZN(n1246) );
NAND2_X1 U980 ( .A1(KEYINPUT44), .A2(n1248), .ZN(n1247) );
XOR2_X1 U981 ( .A(G116), .B(n1081), .Z(n1248) );
XNOR2_X1 U982 ( .A(n1249), .B(G119), .ZN(n1081) );
INV_X1 U983 ( .A(G113), .ZN(n1249) );
NAND3_X1 U984 ( .A1(n1250), .A2(n1251), .A3(KEYINPUT54), .ZN(n1080) );
NAND2_X1 U985 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
INV_X1 U986 ( .A(KEYINPUT6), .ZN(n1253) );
XNOR2_X1 U987 ( .A(G104), .B(G107), .ZN(n1252) );
NAND3_X1 U988 ( .A1(G104), .A2(n1212), .A3(KEYINPUT6), .ZN(n1250) );
INV_X1 U989 ( .A(G107), .ZN(n1212) );
XNOR2_X1 U990 ( .A(n1003), .B(KEYINPUT47), .ZN(n1176) );
NAND2_X1 U991 ( .A1(G214), .A2(n1237), .ZN(n1003) );
NAND2_X1 U992 ( .A1(n1254), .A2(n1111), .ZN(n1237) );
INV_X1 U993 ( .A(G237), .ZN(n1254) );
INV_X1 U994 ( .A(n1015), .ZN(n1010) );
NAND2_X1 U995 ( .A1(n1177), .A2(n1183), .ZN(n1015) );
XOR2_X1 U996 ( .A(n1178), .B(KEYINPUT17), .Z(n1183) );
NAND3_X1 U997 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1178) );
NAND2_X1 U998 ( .A1(G472), .A2(n1258), .ZN(n1257) );
OR3_X1 U999 ( .A1(n1258), .A2(G472), .A3(KEYINPUT56), .ZN(n1256) );
AND2_X1 U1000 ( .A1(KEYINPUT28), .A2(n1030), .ZN(n1258) );
NAND2_X1 U1001 ( .A1(KEYINPUT56), .A2(n1259), .ZN(n1255) );
OR2_X1 U1002 ( .A1(n1030), .A2(G472), .ZN(n1259) );
NAND2_X1 U1003 ( .A1(n1260), .A2(n1111), .ZN(n1030) );
XOR2_X1 U1004 ( .A(n1107), .B(KEYINPUT49), .Z(n1260) );
XOR2_X1 U1005 ( .A(n1261), .B(n1262), .Z(n1107) );
XOR2_X1 U1006 ( .A(n1199), .B(n1263), .Z(n1262) );
XNOR2_X1 U1007 ( .A(n1264), .B(n1079), .ZN(n1263) );
XNOR2_X1 U1008 ( .A(n1230), .B(G116), .ZN(n1079) );
INV_X1 U1009 ( .A(G101), .ZN(n1230) );
INV_X1 U1010 ( .A(n1139), .ZN(n1264) );
XOR2_X1 U1011 ( .A(G128), .B(n1228), .Z(n1139) );
XNOR2_X1 U1012 ( .A(n1168), .B(G146), .ZN(n1228) );
INV_X1 U1013 ( .A(G143), .ZN(n1168) );
XOR2_X1 U1014 ( .A(G113), .B(G131), .Z(n1199) );
XOR2_X1 U1015 ( .A(n1265), .B(n1266), .Z(n1261) );
XNOR2_X1 U1016 ( .A(n1267), .B(KEYINPUT0), .ZN(n1266) );
NAND2_X1 U1017 ( .A1(KEYINPUT58), .A2(G119), .ZN(n1267) );
XOR2_X1 U1018 ( .A(n1223), .B(n1268), .Z(n1265) );
AND2_X1 U1019 ( .A1(n1198), .A2(G210), .ZN(n1268) );
NOR2_X1 U1020 ( .A1(G953), .A2(G237), .ZN(n1198) );
XNOR2_X1 U1021 ( .A(n1269), .B(n1055), .ZN(n1223) );
NAND2_X1 U1022 ( .A1(n1270), .A2(KEYINPUT31), .ZN(n1269) );
XNOR2_X1 U1023 ( .A(G134), .B(KEYINPUT43), .ZN(n1270) );
INV_X1 U1024 ( .A(n1184), .ZN(n1177) );
XOR2_X1 U1025 ( .A(n1271), .B(n1272), .Z(n1184) );
INV_X1 U1026 ( .A(n1039), .ZN(n1272) );
NOR2_X1 U1027 ( .A1(n1092), .A2(G902), .ZN(n1039) );
XNOR2_X1 U1028 ( .A(n1273), .B(n1274), .ZN(n1092) );
XOR2_X1 U1029 ( .A(n1275), .B(n1276), .Z(n1274) );
XNOR2_X1 U1030 ( .A(G140), .B(n1055), .ZN(n1276) );
INV_X1 U1031 ( .A(G137), .ZN(n1055) );
XOR2_X1 U1032 ( .A(KEYINPUT3), .B(G146), .Z(n1275) );
XOR2_X1 U1033 ( .A(n1277), .B(n1278), .Z(n1273) );
XOR2_X1 U1034 ( .A(n1279), .B(n1280), .Z(n1278) );
NAND2_X1 U1035 ( .A1(G221), .A2(n1214), .ZN(n1280) );
AND2_X1 U1036 ( .A1(G234), .A2(n1043), .ZN(n1214) );
INV_X1 U1037 ( .A(G953), .ZN(n1043) );
NAND2_X1 U1038 ( .A1(n1281), .A2(KEYINPUT2), .ZN(n1279) );
XOR2_X1 U1039 ( .A(n1282), .B(G128), .Z(n1281) );
NAND2_X1 U1040 ( .A1(KEYINPUT37), .A2(n1283), .ZN(n1282) );
INV_X1 U1041 ( .A(G119), .ZN(n1283) );
XNOR2_X1 U1042 ( .A(G110), .B(G125), .ZN(n1277) );
NAND2_X1 U1043 ( .A1(KEYINPUT62), .A2(n1037), .ZN(n1271) );
NAND2_X1 U1044 ( .A1(G217), .A2(n1216), .ZN(n1037) );
NAND2_X1 U1045 ( .A1(n1284), .A2(n1111), .ZN(n1216) );
INV_X1 U1046 ( .A(G902), .ZN(n1111) );
XNOR2_X1 U1047 ( .A(G234), .B(KEYINPUT32), .ZN(n1284) );
endmodule


