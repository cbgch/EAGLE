//Key = 0000101110100010001011000000111011100110101000001110011110011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341;

XOR2_X1 U727 ( .A(n1021), .B(n1022), .Z(G9) );
XNOR2_X1 U728 ( .A(KEYINPUT60), .B(n1023), .ZN(n1022) );
NAND4_X1 U729 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1021) );
XNOR2_X1 U730 ( .A(KEYINPUT45), .B(n1028), .ZN(n1027) );
NOR2_X1 U731 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U732 ( .A1(G953), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1030) );
NOR3_X1 U733 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1032) );
NOR2_X1 U734 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR3_X1 U735 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NOR2_X1 U736 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U737 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U738 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U739 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U740 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
XNOR2_X1 U741 ( .A(KEYINPUT17), .B(n1052), .ZN(n1051) );
NOR2_X1 U742 ( .A1(n1053), .A2(n1054), .ZN(n1050) );
NOR2_X1 U743 ( .A1(n1055), .A2(n1056), .ZN(n1046) );
NOR2_X1 U744 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U745 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR3_X1 U746 ( .A1(n1049), .A2(n1061), .A3(n1056), .ZN(n1042) );
NOR4_X1 U747 ( .A1(n1062), .A2(n1045), .A3(n1056), .A4(n1049), .ZN(n1037) );
INV_X1 U748 ( .A(n1063), .ZN(n1045) );
NOR2_X1 U749 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U750 ( .A1(n1066), .A2(n1039), .ZN(n1064) );
INV_X1 U751 ( .A(n1067), .ZN(n1035) );
NOR3_X1 U752 ( .A1(n1031), .A2(G953), .A3(G952), .ZN(n1029) );
AND4_X1 U753 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1031) );
NOR4_X1 U754 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1071) );
XNOR2_X1 U755 ( .A(KEYINPUT36), .B(n1076), .ZN(n1075) );
XNOR2_X1 U756 ( .A(G478), .B(n1077), .ZN(n1073) );
NOR2_X1 U757 ( .A1(KEYINPUT24), .A2(n1078), .ZN(n1077) );
XOR2_X1 U758 ( .A(n1079), .B(KEYINPUT59), .Z(n1078) );
XNOR2_X1 U759 ( .A(n1080), .B(KEYINPUT14), .ZN(n1072) );
AND3_X1 U760 ( .A1(n1081), .A2(n1060), .A3(n1066), .ZN(n1070) );
OR2_X1 U761 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XNOR2_X1 U762 ( .A(G469), .B(KEYINPUT33), .ZN(n1083) );
XOR2_X1 U763 ( .A(n1084), .B(KEYINPUT26), .Z(n1082) );
XOR2_X1 U764 ( .A(n1085), .B(n1086), .Z(n1069) );
NOR2_X1 U765 ( .A1(n1087), .A2(KEYINPUT58), .ZN(n1086) );
XOR2_X1 U766 ( .A(KEYINPUT4), .B(n1088), .Z(n1068) );
NOR2_X1 U767 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XNOR2_X1 U768 ( .A(KEYINPUT26), .B(n1084), .ZN(n1090) );
XOR2_X1 U769 ( .A(n1091), .B(n1092), .Z(G72) );
XOR2_X1 U770 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U771 ( .A1(G953), .A2(n1095), .ZN(n1094) );
NAND2_X1 U772 ( .A1(n1096), .A2(n1097), .ZN(n1093) );
NAND2_X1 U773 ( .A1(G953), .A2(n1098), .ZN(n1097) );
XOR2_X1 U774 ( .A(n1099), .B(n1100), .Z(n1096) );
XNOR2_X1 U775 ( .A(n1101), .B(n1102), .ZN(n1100) );
NAND2_X1 U776 ( .A1(n1103), .A2(KEYINPUT49), .ZN(n1101) );
XNOR2_X1 U777 ( .A(G125), .B(G140), .ZN(n1103) );
XOR2_X1 U778 ( .A(n1104), .B(n1105), .Z(n1099) );
NOR2_X1 U779 ( .A1(KEYINPUT57), .A2(G137), .ZN(n1105) );
XNOR2_X1 U780 ( .A(G131), .B(G134), .ZN(n1104) );
NAND2_X1 U781 ( .A1(G953), .A2(n1106), .ZN(n1091) );
NAND2_X1 U782 ( .A1(G900), .A2(G227), .ZN(n1106) );
XOR2_X1 U783 ( .A(n1107), .B(n1108), .Z(G69) );
NOR2_X1 U784 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U785 ( .A1(n1111), .A2(n1112), .ZN(n1109) );
NAND2_X1 U786 ( .A1(n1113), .A2(n1114), .ZN(n1107) );
NAND3_X1 U787 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
XNOR2_X1 U788 ( .A(n1118), .B(n1119), .ZN(n1116) );
NAND2_X1 U789 ( .A1(G953), .A2(n1112), .ZN(n1115) );
XOR2_X1 U790 ( .A(n1120), .B(KEYINPUT61), .Z(n1113) );
NAND3_X1 U791 ( .A1(n1121), .A2(n1110), .A3(n1122), .ZN(n1120) );
XNOR2_X1 U792 ( .A(n1119), .B(n1123), .ZN(n1122) );
NOR2_X1 U793 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XOR2_X1 U794 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U795 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NOR2_X1 U796 ( .A1(n1124), .A2(n1130), .ZN(G63) );
XNOR2_X1 U797 ( .A(n1131), .B(n1132), .ZN(n1130) );
XOR2_X1 U798 ( .A(KEYINPUT62), .B(n1133), .Z(n1132) );
NOR2_X1 U799 ( .A1(n1134), .A2(n1129), .ZN(n1133) );
NOR2_X1 U800 ( .A1(n1124), .A2(n1135), .ZN(G60) );
XNOR2_X1 U801 ( .A(n1136), .B(n1137), .ZN(n1135) );
AND2_X1 U802 ( .A1(G475), .A2(n1138), .ZN(n1137) );
XNOR2_X1 U803 ( .A(n1139), .B(n1140), .ZN(G6) );
NOR3_X1 U804 ( .A1(n1141), .A2(n1028), .A3(n1056), .ZN(n1140) );
NAND3_X1 U805 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1141) );
OR2_X1 U806 ( .A1(n1026), .A2(KEYINPUT52), .ZN(n1143) );
NAND2_X1 U807 ( .A1(KEYINPUT52), .A2(n1145), .ZN(n1142) );
NOR2_X1 U808 ( .A1(n1124), .A2(n1146), .ZN(G57) );
XOR2_X1 U809 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U810 ( .A(n1149), .B(n1150), .Z(n1148) );
NAND3_X1 U811 ( .A1(n1151), .A2(n1152), .A3(G472), .ZN(n1149) );
NAND2_X1 U812 ( .A1(KEYINPUT8), .A2(n1129), .ZN(n1152) );
NAND2_X1 U813 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
INV_X1 U814 ( .A(KEYINPUT8), .ZN(n1154) );
NAND2_X1 U815 ( .A1(n1155), .A2(n1033), .ZN(n1153) );
XOR2_X1 U816 ( .A(n1156), .B(n1157), .Z(n1147) );
NAND2_X1 U817 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
INV_X1 U818 ( .A(n1160), .ZN(n1159) );
NAND2_X1 U819 ( .A1(n1161), .A2(n1162), .ZN(n1158) );
XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n1163), .ZN(n1161) );
NAND4_X1 U821 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1156) );
NAND2_X1 U822 ( .A1(KEYINPUT13), .A2(n1102), .ZN(n1167) );
NAND3_X1 U823 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1166) );
INV_X1 U824 ( .A(KEYINPUT13), .ZN(n1169) );
XNOR2_X1 U825 ( .A(n1171), .B(KEYINPUT1), .ZN(n1168) );
NAND3_X1 U826 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1165) );
INV_X1 U827 ( .A(KEYINPUT32), .ZN(n1174) );
NAND2_X1 U828 ( .A1(KEYINPUT1), .A2(n1170), .ZN(n1173) );
NAND3_X1 U829 ( .A1(n1171), .A2(n1175), .A3(KEYINPUT32), .ZN(n1164) );
OR2_X1 U830 ( .A1(n1102), .A2(KEYINPUT1), .ZN(n1175) );
NOR2_X1 U831 ( .A1(n1124), .A2(n1176), .ZN(G54) );
NOR2_X1 U832 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XOR2_X1 U833 ( .A(n1179), .B(n1180), .Z(n1178) );
AND2_X1 U834 ( .A1(n1181), .A2(KEYINPUT28), .ZN(n1180) );
NOR2_X1 U835 ( .A1(n1089), .A2(n1129), .ZN(n1179) );
NOR2_X1 U836 ( .A1(KEYINPUT28), .A2(n1181), .ZN(n1177) );
XNOR2_X1 U837 ( .A(n1182), .B(n1183), .ZN(n1181) );
XNOR2_X1 U838 ( .A(n1184), .B(n1172), .ZN(n1183) );
INV_X1 U839 ( .A(n1171), .ZN(n1172) );
XOR2_X1 U840 ( .A(n1185), .B(n1186), .Z(n1182) );
NOR2_X1 U841 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U842 ( .A(KEYINPUT19), .B(n1189), .Z(n1188) );
AND2_X1 U843 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U844 ( .A1(n1191), .A2(n1190), .ZN(n1187) );
NAND2_X1 U845 ( .A1(KEYINPUT21), .A2(n1192), .ZN(n1185) );
XOR2_X1 U846 ( .A(KEYINPUT53), .B(n1193), .Z(n1192) );
NOR2_X1 U847 ( .A1(n1124), .A2(n1194), .ZN(G51) );
XOR2_X1 U848 ( .A(n1195), .B(n1196), .Z(n1194) );
NOR2_X1 U849 ( .A1(KEYINPUT51), .A2(n1197), .ZN(n1196) );
NAND2_X1 U850 ( .A1(n1138), .A2(n1198), .ZN(n1195) );
XOR2_X1 U851 ( .A(KEYINPUT9), .B(n1085), .Z(n1198) );
INV_X1 U852 ( .A(n1129), .ZN(n1138) );
NAND2_X1 U853 ( .A1(G902), .A2(n1033), .ZN(n1129) );
NAND2_X1 U854 ( .A1(n1117), .A2(n1095), .ZN(n1033) );
AND2_X1 U855 ( .A1(n1199), .A2(n1200), .ZN(n1095) );
NOR4_X1 U856 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
NOR4_X1 U857 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1199) );
NOR3_X1 U858 ( .A1(n1209), .A2(n1028), .A3(n1210), .ZN(n1208) );
INV_X1 U859 ( .A(n1211), .ZN(n1205) );
INV_X1 U860 ( .A(n1121), .ZN(n1117) );
NAND4_X1 U861 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1121) );
AND3_X1 U862 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
NAND2_X1 U863 ( .A1(n1058), .A2(n1219), .ZN(n1214) );
NAND2_X1 U864 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NAND4_X1 U865 ( .A1(n1222), .A2(n1063), .A3(n1223), .A4(n1224), .ZN(n1221) );
OR2_X1 U866 ( .A1(n1026), .A2(KEYINPUT63), .ZN(n1224) );
NAND2_X1 U867 ( .A1(KEYINPUT63), .A2(n1145), .ZN(n1223) );
NAND2_X1 U868 ( .A1(n1225), .A2(n1226), .ZN(n1145) );
OR3_X1 U869 ( .A1(n1227), .A2(n1061), .A3(n1056), .ZN(n1220) );
INV_X1 U870 ( .A(n1025), .ZN(n1056) );
NOR2_X1 U871 ( .A1(n1024), .A2(n1144), .ZN(n1061) );
NOR2_X1 U872 ( .A1(n1110), .A2(G952), .ZN(n1124) );
XNOR2_X1 U873 ( .A(G146), .B(n1228), .ZN(G48) );
NAND3_X1 U874 ( .A1(n1229), .A2(n1144), .A3(n1230), .ZN(n1228) );
XNOR2_X1 U875 ( .A(n1058), .B(KEYINPUT6), .ZN(n1230) );
NAND2_X1 U876 ( .A1(n1231), .A2(n1232), .ZN(G45) );
NAND2_X1 U877 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
XOR2_X1 U878 ( .A(KEYINPUT46), .B(n1206), .Z(n1233) );
NAND2_X1 U879 ( .A1(n1235), .A2(G143), .ZN(n1231) );
XOR2_X1 U880 ( .A(KEYINPUT56), .B(n1206), .Z(n1235) );
NOR4_X1 U881 ( .A1(n1052), .A2(n1028), .A3(n1236), .A4(n1237), .ZN(n1206) );
NAND3_X1 U882 ( .A1(n1065), .A2(n1074), .A3(n1238), .ZN(n1237) );
XOR2_X1 U883 ( .A(G140), .B(n1207), .Z(G42) );
AND4_X1 U884 ( .A1(n1239), .A2(n1144), .A3(n1076), .A4(n1080), .ZN(n1207) );
XNOR2_X1 U885 ( .A(G137), .B(n1211), .ZN(G39) );
NAND4_X1 U886 ( .A1(n1239), .A2(n1063), .A3(n1080), .A4(n1054), .ZN(n1211) );
XOR2_X1 U887 ( .A(G134), .B(n1204), .Z(G36) );
AND3_X1 U888 ( .A1(n1222), .A2(n1024), .A3(n1239), .ZN(n1204) );
XOR2_X1 U889 ( .A(G131), .B(n1203), .Z(G33) );
AND3_X1 U890 ( .A1(n1222), .A2(n1144), .A3(n1239), .ZN(n1203) );
NOR4_X1 U891 ( .A1(n1039), .A2(n1236), .A3(n1041), .A4(n1028), .ZN(n1239) );
XOR2_X1 U892 ( .A(G128), .B(n1202), .Z(G30) );
NOR3_X1 U893 ( .A1(n1240), .A2(n1028), .A3(n1209), .ZN(n1202) );
INV_X1 U894 ( .A(n1229), .ZN(n1209) );
NOR2_X1 U895 ( .A1(n1241), .A2(n1076), .ZN(n1229) );
XNOR2_X1 U896 ( .A(n1163), .B(n1242), .ZN(G3) );
NOR2_X1 U897 ( .A1(n1243), .A2(n1052), .ZN(n1242) );
INV_X1 U898 ( .A(n1222), .ZN(n1052) );
XOR2_X1 U899 ( .A(G125), .B(n1201), .Z(G27) );
NOR4_X1 U900 ( .A1(n1241), .A2(n1210), .A3(n1054), .A4(n1049), .ZN(n1201) );
OR3_X1 U901 ( .A1(n1226), .A2(n1053), .A3(n1236), .ZN(n1241) );
NAND2_X1 U902 ( .A1(n1067), .A2(n1244), .ZN(n1236) );
NAND2_X1 U903 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND3_X1 U904 ( .A1(G902), .A2(n1098), .A3(G953), .ZN(n1245) );
INV_X1 U905 ( .A(G900), .ZN(n1098) );
XNOR2_X1 U906 ( .A(G122), .B(n1212), .ZN(G24) );
NAND4_X1 U907 ( .A1(n1247), .A2(n1025), .A3(n1238), .A4(n1074), .ZN(n1212) );
NOR2_X1 U908 ( .A1(n1054), .A2(n1080), .ZN(n1025) );
XNOR2_X1 U909 ( .A(G119), .B(n1213), .ZN(G21) );
NAND4_X1 U910 ( .A1(n1247), .A2(n1063), .A3(n1080), .A4(n1054), .ZN(n1213) );
XNOR2_X1 U911 ( .A(G116), .B(n1216), .ZN(G18) );
NAND3_X1 U912 ( .A1(n1247), .A2(n1024), .A3(n1222), .ZN(n1216) );
XNOR2_X1 U913 ( .A(G113), .B(n1218), .ZN(G15) );
NAND3_X1 U914 ( .A1(n1144), .A2(n1247), .A3(n1222), .ZN(n1218) );
NOR2_X1 U915 ( .A1(n1080), .A2(n1076), .ZN(n1222) );
INV_X1 U916 ( .A(n1054), .ZN(n1076) );
NOR2_X1 U917 ( .A1(n1049), .A2(n1227), .ZN(n1247) );
NAND2_X1 U918 ( .A1(n1248), .A2(n1060), .ZN(n1049) );
INV_X1 U919 ( .A(n1059), .ZN(n1248) );
INV_X1 U920 ( .A(n1210), .ZN(n1144) );
NAND2_X1 U921 ( .A1(n1249), .A2(n1074), .ZN(n1210) );
XNOR2_X1 U922 ( .A(KEYINPUT48), .B(n1250), .ZN(n1249) );
XNOR2_X1 U923 ( .A(G110), .B(n1217), .ZN(G12) );
OR3_X1 U924 ( .A1(n1054), .A2(n1053), .A3(n1243), .ZN(n1217) );
NAND3_X1 U925 ( .A1(n1058), .A2(n1063), .A3(n1026), .ZN(n1243) );
INV_X1 U926 ( .A(n1227), .ZN(n1026) );
NAND2_X1 U927 ( .A1(n1225), .A2(n1065), .ZN(n1227) );
INV_X1 U928 ( .A(n1226), .ZN(n1065) );
NAND2_X1 U929 ( .A1(n1251), .A2(n1039), .ZN(n1226) );
XOR2_X1 U930 ( .A(n1087), .B(n1252), .Z(n1039) );
XOR2_X1 U931 ( .A(KEYINPUT39), .B(n1085), .Z(n1252) );
AND2_X1 U932 ( .A1(G210), .A2(n1253), .ZN(n1085) );
NOR2_X1 U933 ( .A1(n1197), .A2(G902), .ZN(n1087) );
XOR2_X1 U934 ( .A(n1254), .B(n1255), .Z(n1197) );
XOR2_X1 U935 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U936 ( .A(G125), .B(n1258), .Z(n1257) );
NOR2_X1 U937 ( .A1(KEYINPUT31), .A2(n1123), .ZN(n1258) );
INV_X1 U938 ( .A(n1118), .ZN(n1123) );
XNOR2_X1 U939 ( .A(n1259), .B(n1260), .ZN(n1118) );
NAND2_X1 U940 ( .A1(KEYINPUT29), .A2(n1023), .ZN(n1259) );
NOR2_X1 U941 ( .A1(G953), .A2(n1111), .ZN(n1256) );
INV_X1 U942 ( .A(G224), .ZN(n1111) );
XNOR2_X1 U943 ( .A(n1119), .B(n1102), .ZN(n1254) );
XOR2_X1 U944 ( .A(n1261), .B(n1262), .Z(n1119) );
XOR2_X1 U945 ( .A(n1263), .B(G113), .Z(n1261) );
NAND2_X1 U946 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NAND2_X1 U947 ( .A1(G122), .A2(n1266), .ZN(n1265) );
XOR2_X1 U948 ( .A(KEYINPUT55), .B(n1267), .Z(n1264) );
NOR2_X1 U949 ( .A1(G122), .A2(n1266), .ZN(n1267) );
INV_X1 U950 ( .A(G110), .ZN(n1266) );
INV_X1 U951 ( .A(n1041), .ZN(n1251) );
XNOR2_X1 U952 ( .A(n1066), .B(KEYINPUT16), .ZN(n1041) );
NAND2_X1 U953 ( .A1(G214), .A2(n1253), .ZN(n1066) );
NAND2_X1 U954 ( .A1(n1268), .A2(n1269), .ZN(n1253) );
AND2_X1 U955 ( .A1(n1270), .A2(n1067), .ZN(n1225) );
NAND2_X1 U956 ( .A1(G237), .A2(G234), .ZN(n1067) );
NAND2_X1 U957 ( .A1(n1246), .A2(n1271), .ZN(n1270) );
NAND3_X1 U958 ( .A1(G902), .A2(n1112), .A3(G953), .ZN(n1271) );
INV_X1 U959 ( .A(G898), .ZN(n1112) );
NAND2_X1 U960 ( .A1(n1272), .A2(n1110), .ZN(n1246) );
XNOR2_X1 U961 ( .A(KEYINPUT23), .B(n1034), .ZN(n1272) );
XNOR2_X1 U962 ( .A(G952), .B(KEYINPUT41), .ZN(n1034) );
NAND2_X1 U963 ( .A1(n1273), .A2(n1274), .ZN(n1063) );
OR2_X1 U964 ( .A1(n1240), .A2(KEYINPUT48), .ZN(n1274) );
INV_X1 U965 ( .A(n1024), .ZN(n1240) );
NOR2_X1 U966 ( .A1(n1074), .A2(n1250), .ZN(n1024) );
NAND3_X1 U967 ( .A1(n1275), .A2(n1250), .A3(KEYINPUT48), .ZN(n1273) );
INV_X1 U968 ( .A(n1238), .ZN(n1250) );
XOR2_X1 U969 ( .A(n1079), .B(n1134), .Z(n1238) );
INV_X1 U970 ( .A(G478), .ZN(n1134) );
NAND2_X1 U971 ( .A1(n1131), .A2(n1155), .ZN(n1079) );
XNOR2_X1 U972 ( .A(n1276), .B(n1277), .ZN(n1131) );
XOR2_X1 U973 ( .A(n1278), .B(n1279), .Z(n1277) );
XNOR2_X1 U974 ( .A(G107), .B(G122), .ZN(n1279) );
NAND2_X1 U975 ( .A1(G217), .A2(n1280), .ZN(n1278) );
XNOR2_X1 U976 ( .A(n1281), .B(n1282), .ZN(n1276) );
XOR2_X1 U977 ( .A(n1283), .B(n1284), .Z(n1282) );
NOR2_X1 U978 ( .A1(G134), .A2(KEYINPUT44), .ZN(n1283) );
INV_X1 U979 ( .A(n1074), .ZN(n1275) );
XNOR2_X1 U980 ( .A(n1285), .B(G475), .ZN(n1074) );
NAND2_X1 U981 ( .A1(n1136), .A2(n1155), .ZN(n1285) );
XNOR2_X1 U982 ( .A(n1286), .B(n1287), .ZN(n1136) );
XOR2_X1 U983 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U984 ( .A(n1290), .B(n1291), .Z(n1289) );
NAND2_X1 U985 ( .A1(KEYINPUT38), .A2(n1292), .ZN(n1291) );
NAND2_X1 U986 ( .A1(n1293), .A2(n1294), .ZN(n1290) );
NAND2_X1 U987 ( .A1(n1295), .A2(n1139), .ZN(n1294) );
XOR2_X1 U988 ( .A(KEYINPUT18), .B(n1296), .Z(n1293) );
NOR2_X1 U989 ( .A1(n1295), .A2(n1139), .ZN(n1296) );
INV_X1 U990 ( .A(G104), .ZN(n1139) );
XOR2_X1 U991 ( .A(G122), .B(n1297), .Z(n1295) );
NOR2_X1 U992 ( .A1(G113), .A2(KEYINPUT25), .ZN(n1297) );
NOR2_X1 U993 ( .A1(G140), .A2(KEYINPUT11), .ZN(n1288) );
XOR2_X1 U994 ( .A(n1298), .B(n1299), .Z(n1286) );
XOR2_X1 U995 ( .A(G125), .B(n1300), .Z(n1299) );
AND3_X1 U996 ( .A1(G214), .A2(n1110), .A3(n1269), .ZN(n1300) );
XNOR2_X1 U997 ( .A(G131), .B(G143), .ZN(n1298) );
INV_X1 U998 ( .A(n1028), .ZN(n1058) );
NAND2_X1 U999 ( .A1(n1059), .A2(n1060), .ZN(n1028) );
NAND2_X1 U1000 ( .A1(G221), .A2(n1301), .ZN(n1060) );
XNOR2_X1 U1001 ( .A(n1084), .B(n1302), .ZN(n1059) );
XNOR2_X1 U1002 ( .A(KEYINPUT27), .B(n1089), .ZN(n1302) );
INV_X1 U1003 ( .A(G469), .ZN(n1089) );
NAND2_X1 U1004 ( .A1(n1303), .A2(n1155), .ZN(n1084) );
XOR2_X1 U1005 ( .A(n1304), .B(n1305), .Z(n1303) );
XNOR2_X1 U1006 ( .A(n1306), .B(n1191), .ZN(n1305) );
NAND2_X1 U1007 ( .A1(KEYINPUT40), .A2(n1307), .ZN(n1306) );
XOR2_X1 U1008 ( .A(n1193), .B(n1308), .Z(n1307) );
XOR2_X1 U1009 ( .A(n1309), .B(n1184), .Z(n1308) );
XNOR2_X1 U1010 ( .A(n1102), .B(KEYINPUT15), .ZN(n1184) );
INV_X1 U1011 ( .A(n1170), .ZN(n1102) );
NOR2_X1 U1012 ( .A1(KEYINPUT35), .A2(n1171), .ZN(n1309) );
XNOR2_X1 U1013 ( .A(n1310), .B(n1260), .ZN(n1193) );
XNOR2_X1 U1014 ( .A(n1163), .B(G104), .ZN(n1260) );
NAND2_X1 U1015 ( .A1(KEYINPUT10), .A2(n1311), .ZN(n1310) );
XNOR2_X1 U1016 ( .A(KEYINPUT3), .B(n1023), .ZN(n1311) );
INV_X1 U1017 ( .A(G107), .ZN(n1023) );
XNOR2_X1 U1018 ( .A(KEYINPUT54), .B(n1190), .ZN(n1304) );
NAND2_X1 U1019 ( .A1(G227), .A2(n1110), .ZN(n1190) );
INV_X1 U1020 ( .A(n1080), .ZN(n1053) );
XOR2_X1 U1021 ( .A(n1312), .B(n1128), .Z(n1080) );
NAND2_X1 U1022 ( .A1(G217), .A2(n1301), .ZN(n1128) );
NAND2_X1 U1023 ( .A1(n1268), .A2(n1313), .ZN(n1301) );
XOR2_X1 U1024 ( .A(KEYINPUT2), .B(G234), .Z(n1313) );
XNOR2_X1 U1025 ( .A(G902), .B(KEYINPUT0), .ZN(n1268) );
OR2_X1 U1026 ( .A1(n1127), .A2(G902), .ZN(n1312) );
XNOR2_X1 U1027 ( .A(n1314), .B(n1315), .ZN(n1127) );
XOR2_X1 U1028 ( .A(n1316), .B(n1317), .Z(n1315) );
XOR2_X1 U1029 ( .A(G128), .B(G125), .Z(n1317) );
XNOR2_X1 U1030 ( .A(KEYINPUT5), .B(n1318), .ZN(n1316) );
INV_X1 U1031 ( .A(G137), .ZN(n1318) );
XOR2_X1 U1032 ( .A(n1319), .B(n1320), .Z(n1314) );
XNOR2_X1 U1033 ( .A(G119), .B(n1321), .ZN(n1320) );
NAND2_X1 U1034 ( .A1(KEYINPUT37), .A2(n1292), .ZN(n1321) );
INV_X1 U1035 ( .A(G146), .ZN(n1292) );
XOR2_X1 U1036 ( .A(n1322), .B(n1191), .Z(n1319) );
XOR2_X1 U1037 ( .A(G110), .B(G140), .Z(n1191) );
NAND2_X1 U1038 ( .A1(G221), .A2(n1280), .ZN(n1322) );
AND2_X1 U1039 ( .A1(G234), .A2(n1110), .ZN(n1280) );
XNOR2_X1 U1040 ( .A(n1323), .B(G472), .ZN(n1054) );
NAND2_X1 U1041 ( .A1(n1324), .A2(n1155), .ZN(n1323) );
INV_X1 U1042 ( .A(G902), .ZN(n1155) );
XOR2_X1 U1043 ( .A(n1325), .B(n1326), .Z(n1324) );
NOR2_X1 U1044 ( .A1(n1160), .A2(n1327), .ZN(n1326) );
NOR2_X1 U1045 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
XNOR2_X1 U1046 ( .A(G101), .B(KEYINPUT42), .ZN(n1329) );
INV_X1 U1047 ( .A(n1162), .ZN(n1328) );
NOR2_X1 U1048 ( .A1(n1163), .A2(n1162), .ZN(n1160) );
NAND3_X1 U1049 ( .A1(n1269), .A2(n1110), .A3(G210), .ZN(n1162) );
INV_X1 U1050 ( .A(G953), .ZN(n1110) );
INV_X1 U1051 ( .A(G237), .ZN(n1269) );
INV_X1 U1052 ( .A(G101), .ZN(n1163) );
NOR2_X1 U1053 ( .A1(KEYINPUT22), .A2(n1330), .ZN(n1325) );
NOR3_X1 U1054 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(n1330) );
AND2_X1 U1055 ( .A1(n1334), .A2(n1150), .ZN(n1333) );
NOR3_X1 U1056 ( .A1(n1150), .A2(KEYINPUT43), .A3(n1334), .ZN(n1332) );
NAND2_X1 U1057 ( .A1(KEYINPUT34), .A2(n1335), .ZN(n1334) );
XNOR2_X1 U1058 ( .A(n1262), .B(n1336), .ZN(n1150) );
NOR2_X1 U1059 ( .A1(G113), .A2(KEYINPUT47), .ZN(n1336) );
XOR2_X1 U1060 ( .A(G119), .B(n1281), .Z(n1262) );
XOR2_X1 U1061 ( .A(G116), .B(KEYINPUT7), .Z(n1281) );
NOR2_X1 U1062 ( .A1(n1335), .A2(n1337), .ZN(n1331) );
INV_X1 U1063 ( .A(KEYINPUT43), .ZN(n1337) );
XNOR2_X1 U1064 ( .A(n1171), .B(n1170), .ZN(n1335) );
XNOR2_X1 U1065 ( .A(n1338), .B(n1284), .ZN(n1170) );
XNOR2_X1 U1066 ( .A(G128), .B(n1234), .ZN(n1284) );
INV_X1 U1067 ( .A(G143), .ZN(n1234) );
XNOR2_X1 U1068 ( .A(G146), .B(KEYINPUT20), .ZN(n1338) );
XNOR2_X1 U1069 ( .A(n1339), .B(n1340), .ZN(n1171) );
NOR2_X1 U1070 ( .A1(KEYINPUT12), .A2(n1341), .ZN(n1340) );
XNOR2_X1 U1071 ( .A(G131), .B(KEYINPUT50), .ZN(n1341) );
XNOR2_X1 U1072 ( .A(G134), .B(G137), .ZN(n1339) );
endmodule


