//Key = 1110111110000010011000100101000111101100101100100111011111000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399;

XNOR2_X1 U759 ( .A(n1064), .B(n1065), .ZN(G9) );
AND2_X1 U760 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(G75) );
NOR4_X1 U762 ( .A1(n1070), .A2(n1071), .A3(G953), .A4(n1072), .ZN(n1069) );
NOR3_X1 U763 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1071) );
NOR2_X1 U764 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U765 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U766 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR2_X1 U767 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR3_X1 U768 ( .A1(n1084), .A2(n1066), .A3(n1085), .ZN(n1082) );
NOR2_X1 U769 ( .A1(KEYINPUT17), .A2(n1086), .ZN(n1085) );
NOR2_X1 U770 ( .A1(n1087), .A2(n1088), .ZN(n1084) );
NOR2_X1 U771 ( .A1(n1089), .A2(n1090), .ZN(n1080) );
XNOR2_X1 U772 ( .A(KEYINPUT55), .B(n1086), .ZN(n1090) );
NOR3_X1 U773 ( .A1(n1086), .A2(n1091), .A3(n1083), .ZN(n1076) );
NAND3_X1 U774 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1070) );
NAND2_X1 U775 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NAND2_X1 U776 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U777 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U778 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND3_X1 U779 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
NAND2_X1 U780 ( .A1(n1106), .A2(n1107), .ZN(n1101) );
NAND2_X1 U781 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND3_X1 U782 ( .A1(n1103), .A2(n1110), .A3(n1111), .ZN(n1109) );
INV_X1 U783 ( .A(KEYINPUT19), .ZN(n1110) );
NAND2_X1 U784 ( .A1(n1104), .A2(n1112), .ZN(n1108) );
NAND2_X1 U785 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND3_X1 U786 ( .A1(n1115), .A2(n1116), .A3(KEYINPUT17), .ZN(n1114) );
NAND2_X1 U787 ( .A1(KEYINPUT19), .A2(n1117), .ZN(n1097) );
NAND4_X1 U788 ( .A1(n1099), .A2(n1106), .A3(n1111), .A4(n1103), .ZN(n1117) );
INV_X1 U789 ( .A(n1073), .ZN(n1099) );
NOR3_X1 U790 ( .A1(n1072), .A2(G953), .A3(G952), .ZN(n1068) );
AND4_X1 U791 ( .A1(n1118), .A2(n1095), .A3(n1119), .A4(n1120), .ZN(n1072) );
NOR4_X1 U792 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1120) );
XNOR2_X1 U793 ( .A(n1125), .B(KEYINPUT63), .ZN(n1122) );
XNOR2_X1 U794 ( .A(n1126), .B(n1127), .ZN(n1121) );
NAND2_X1 U795 ( .A1(KEYINPUT18), .A2(n1128), .ZN(n1126) );
XNOR2_X1 U796 ( .A(KEYINPUT14), .B(n1129), .ZN(n1128) );
XNOR2_X1 U797 ( .A(n1116), .B(KEYINPUT35), .ZN(n1119) );
XOR2_X1 U798 ( .A(n1130), .B(n1131), .Z(G72) );
NOR2_X1 U799 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NOR2_X1 U800 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
NAND3_X1 U801 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1130) );
NAND3_X1 U802 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1138) );
NAND2_X1 U803 ( .A1(G953), .A2(n1135), .ZN(n1139) );
OR4_X1 U804 ( .A1(n1092), .A2(G953), .A3(n1141), .A4(KEYINPUT62), .ZN(n1137) );
XOR2_X1 U805 ( .A(n1142), .B(n1143), .Z(n1141) );
XNOR2_X1 U806 ( .A(n1144), .B(n1145), .ZN(n1143) );
XOR2_X1 U807 ( .A(n1146), .B(n1147), .Z(n1142) );
NOR2_X1 U808 ( .A1(KEYINPUT38), .A2(G134), .ZN(n1147) );
XNOR2_X1 U809 ( .A(G125), .B(G140), .ZN(n1146) );
NAND2_X1 U810 ( .A1(KEYINPUT62), .A2(n1140), .ZN(n1136) );
NAND2_X1 U811 ( .A1(n1148), .A2(n1133), .ZN(n1140) );
NAND2_X1 U812 ( .A1(n1149), .A2(n1150), .ZN(G69) );
NAND2_X1 U813 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U814 ( .A(KEYINPUT22), .B(n1153), .Z(n1149) );
NOR2_X1 U815 ( .A1(n1151), .A2(n1152), .ZN(n1153) );
NAND2_X1 U816 ( .A1(G953), .A2(n1154), .ZN(n1152) );
NAND2_X1 U817 ( .A1(G898), .A2(G224), .ZN(n1154) );
XNOR2_X1 U818 ( .A(n1155), .B(n1156), .ZN(n1151) );
NOR2_X1 U819 ( .A1(n1094), .A2(G953), .ZN(n1156) );
NAND2_X1 U820 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
NAND2_X1 U821 ( .A1(G953), .A2(n1159), .ZN(n1158) );
XOR2_X1 U822 ( .A(n1160), .B(KEYINPUT10), .Z(n1157) );
NOR2_X1 U823 ( .A1(n1161), .A2(n1162), .ZN(G66) );
XOR2_X1 U824 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U825 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
NOR2_X1 U826 ( .A1(n1161), .A2(n1167), .ZN(G63) );
XOR2_X1 U827 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U828 ( .A1(n1170), .A2(n1166), .ZN(n1168) );
NOR2_X1 U829 ( .A1(n1161), .A2(n1171), .ZN(G60) );
XNOR2_X1 U830 ( .A(n1172), .B(n1173), .ZN(n1171) );
NOR2_X1 U831 ( .A1(n1174), .A2(n1166), .ZN(n1173) );
XNOR2_X1 U832 ( .A(G104), .B(n1175), .ZN(G6) );
NOR2_X1 U833 ( .A1(n1176), .A2(n1177), .ZN(G57) );
XOR2_X1 U834 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U835 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U836 ( .A1(n1129), .A2(n1166), .ZN(n1180) );
XOR2_X1 U837 ( .A(n1182), .B(n1183), .Z(n1178) );
NAND2_X1 U838 ( .A1(KEYINPUT46), .A2(n1184), .ZN(n1182) );
NOR2_X1 U839 ( .A1(G952), .A2(n1185), .ZN(n1176) );
XOR2_X1 U840 ( .A(KEYINPUT51), .B(n1186), .Z(n1185) );
NOR4_X1 U841 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(G54) );
AND2_X1 U842 ( .A1(KEYINPUT54), .A2(n1161), .ZN(n1190) );
NOR3_X1 U843 ( .A1(KEYINPUT54), .A2(G952), .A3(n1186), .ZN(n1189) );
INV_X1 U844 ( .A(n1191), .ZN(n1186) );
NOR2_X1 U845 ( .A1(n1192), .A2(n1193), .ZN(n1188) );
XNOR2_X1 U846 ( .A(n1194), .B(KEYINPUT9), .ZN(n1193) );
INV_X1 U847 ( .A(n1195), .ZN(n1192) );
NOR2_X1 U848 ( .A1(n1194), .A2(n1195), .ZN(n1187) );
XOR2_X1 U849 ( .A(n1196), .B(n1197), .Z(n1195) );
XOR2_X1 U850 ( .A(n1198), .B(n1199), .Z(n1197) );
XOR2_X1 U851 ( .A(n1200), .B(n1201), .Z(n1196) );
NOR2_X1 U852 ( .A1(n1166), .A2(n1202), .ZN(n1194) );
INV_X1 U853 ( .A(G469), .ZN(n1202) );
NOR2_X1 U854 ( .A1(n1161), .A2(n1203), .ZN(G51) );
XOR2_X1 U855 ( .A(n1204), .B(n1205), .Z(n1203) );
NOR2_X1 U856 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
XOR2_X1 U857 ( .A(KEYINPUT21), .B(n1208), .Z(n1207) );
NOR2_X1 U858 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
AND2_X1 U859 ( .A1(n1209), .A2(n1210), .ZN(n1206) );
XOR2_X1 U860 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U861 ( .A(KEYINPUT48), .B(n1213), .Z(n1212) );
NOR2_X1 U862 ( .A1(n1214), .A2(n1166), .ZN(n1204) );
NAND2_X1 U863 ( .A1(G902), .A2(n1215), .ZN(n1166) );
NAND2_X1 U864 ( .A1(n1094), .A2(n1092), .ZN(n1215) );
INV_X1 U865 ( .A(n1148), .ZN(n1092) );
NAND4_X1 U866 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1148) );
AND4_X1 U867 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1219) );
NAND2_X1 U868 ( .A1(n1066), .A2(n1224), .ZN(n1218) );
XNOR2_X1 U869 ( .A(KEYINPUT45), .B(n1225), .ZN(n1224) );
NAND3_X1 U870 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1217) );
NAND2_X1 U871 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
NAND2_X1 U872 ( .A1(n1111), .A2(n1231), .ZN(n1230) );
XNOR2_X1 U873 ( .A(KEYINPUT61), .B(n1086), .ZN(n1231) );
NAND2_X1 U874 ( .A1(n1232), .A2(n1066), .ZN(n1229) );
NAND2_X1 U875 ( .A1(n1233), .A2(n1095), .ZN(n1216) );
XOR2_X1 U876 ( .A(n1234), .B(KEYINPUT56), .Z(n1233) );
AND4_X1 U877 ( .A1(n1175), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1094) );
AND4_X1 U878 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1237) );
OR2_X1 U879 ( .A1(n1242), .A2(n1243), .ZN(n1238) );
XOR2_X1 U880 ( .A(KEYINPUT34), .B(n1067), .Z(n1243) );
NOR4_X1 U881 ( .A1(n1113), .A2(n1083), .A3(n1091), .A4(n1244), .ZN(n1067) );
INV_X1 U882 ( .A(n1104), .ZN(n1083) );
NOR3_X1 U883 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1236) );
AND3_X1 U884 ( .A1(n1106), .A2(n1248), .A3(n1232), .ZN(n1247) );
AND4_X1 U885 ( .A1(n1079), .A2(KEYINPUT26), .A3(n1249), .A4(n1250), .ZN(n1246) );
INV_X1 U886 ( .A(n1106), .ZN(n1079) );
NOR2_X1 U887 ( .A1(KEYINPUT26), .A2(n1251), .ZN(n1245) );
NAND3_X1 U888 ( .A1(n1105), .A2(n1104), .A3(n1249), .ZN(n1175) );
NOR2_X1 U889 ( .A1(n1191), .A2(G952), .ZN(n1161) );
XOR2_X1 U890 ( .A(n1133), .B(KEYINPUT11), .Z(n1191) );
XNOR2_X1 U891 ( .A(n1252), .B(n1253), .ZN(G48) );
NOR2_X1 U892 ( .A1(n1242), .A2(n1225), .ZN(n1253) );
NAND2_X1 U893 ( .A1(n1254), .A2(n1232), .ZN(n1225) );
XNOR2_X1 U894 ( .A(G143), .B(n1223), .ZN(G45) );
NAND3_X1 U895 ( .A1(n1228), .A2(n1111), .A3(n1255), .ZN(n1223) );
NOR3_X1 U896 ( .A1(n1242), .A2(n1118), .A3(n1256), .ZN(n1255) );
INV_X1 U897 ( .A(n1257), .ZN(n1118) );
XNOR2_X1 U898 ( .A(G140), .B(n1222), .ZN(G42) );
NAND3_X1 U899 ( .A1(n1250), .A2(n1095), .A3(n1254), .ZN(n1222) );
XNOR2_X1 U900 ( .A(G137), .B(n1258), .ZN(G39) );
NAND2_X1 U901 ( .A1(KEYINPUT4), .A2(n1259), .ZN(n1258) );
INV_X1 U902 ( .A(n1220), .ZN(n1259) );
NAND4_X1 U903 ( .A1(n1228), .A2(n1232), .A3(n1106), .A4(n1095), .ZN(n1220) );
NAND2_X1 U904 ( .A1(n1260), .A2(n1261), .ZN(G36) );
NAND3_X1 U905 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1261) );
NAND2_X1 U906 ( .A1(KEYINPUT30), .A2(n1265), .ZN(n1263) );
NAND2_X1 U907 ( .A1(KEYINPUT31), .A2(G134), .ZN(n1262) );
NAND3_X1 U908 ( .A1(G134), .A2(n1266), .A3(KEYINPUT31), .ZN(n1260) );
NAND2_X1 U909 ( .A1(n1264), .A2(n1267), .ZN(n1266) );
INV_X1 U910 ( .A(KEYINPUT30), .ZN(n1267) );
AND4_X1 U911 ( .A1(n1228), .A2(n1111), .A3(n1095), .A4(n1226), .ZN(n1264) );
XOR2_X1 U912 ( .A(G131), .B(n1268), .Z(G33) );
NOR2_X1 U913 ( .A1(n1086), .A2(n1234), .ZN(n1268) );
NAND2_X1 U914 ( .A1(n1254), .A2(n1111), .ZN(n1234) );
AND2_X1 U915 ( .A1(n1228), .A2(n1105), .ZN(n1254) );
NOR2_X1 U916 ( .A1(n1113), .A2(n1269), .ZN(n1228) );
INV_X1 U917 ( .A(n1095), .ZN(n1086) );
NOR2_X1 U918 ( .A1(n1087), .A2(n1270), .ZN(n1095) );
INV_X1 U919 ( .A(n1088), .ZN(n1270) );
XNOR2_X1 U920 ( .A(G128), .B(n1271), .ZN(G30) );
NAND4_X1 U921 ( .A1(n1226), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1271) );
NOR2_X1 U922 ( .A1(n1242), .A2(n1275), .ZN(n1274) );
XOR2_X1 U923 ( .A(KEYINPUT25), .B(n1269), .Z(n1272) );
XNOR2_X1 U924 ( .A(G101), .B(n1235), .ZN(G3) );
NAND3_X1 U925 ( .A1(n1249), .A2(n1111), .A3(n1106), .ZN(n1235) );
XNOR2_X1 U926 ( .A(G125), .B(n1221), .ZN(G27) );
NAND4_X1 U927 ( .A1(n1250), .A2(n1105), .A3(n1276), .A4(n1103), .ZN(n1221) );
NOR2_X1 U928 ( .A1(n1269), .A2(n1242), .ZN(n1276) );
AND2_X1 U929 ( .A1(n1073), .A2(n1277), .ZN(n1269) );
NAND4_X1 U930 ( .A1(G953), .A2(G902), .A3(n1278), .A4(n1135), .ZN(n1277) );
INV_X1 U931 ( .A(G900), .ZN(n1135) );
XNOR2_X1 U932 ( .A(G122), .B(n1241), .ZN(G24) );
NAND4_X1 U933 ( .A1(n1248), .A2(n1104), .A3(n1279), .A4(n1257), .ZN(n1241) );
NOR2_X1 U934 ( .A1(n1123), .A2(n1280), .ZN(n1104) );
XNOR2_X1 U935 ( .A(G119), .B(n1281), .ZN(G21) );
NAND4_X1 U936 ( .A1(n1232), .A2(n1106), .A3(n1282), .A4(n1103), .ZN(n1281) );
NOR2_X1 U937 ( .A1(n1244), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U938 ( .A(n1066), .B(KEYINPUT15), .ZN(n1283) );
INV_X1 U939 ( .A(n1242), .ZN(n1066) );
INV_X1 U940 ( .A(n1275), .ZN(n1232) );
NAND2_X1 U941 ( .A1(n1280), .A2(n1123), .ZN(n1275) );
XNOR2_X1 U942 ( .A(G116), .B(n1240), .ZN(G18) );
NAND3_X1 U943 ( .A1(n1248), .A2(n1226), .A3(n1111), .ZN(n1240) );
INV_X1 U944 ( .A(n1091), .ZN(n1226) );
NAND2_X1 U945 ( .A1(n1284), .A2(n1257), .ZN(n1091) );
XNOR2_X1 U946 ( .A(KEYINPUT29), .B(n1279), .ZN(n1284) );
NAND2_X1 U947 ( .A1(n1285), .A2(n1286), .ZN(G15) );
OR2_X1 U948 ( .A1(n1239), .A2(G113), .ZN(n1286) );
XOR2_X1 U949 ( .A(n1287), .B(KEYINPUT44), .Z(n1285) );
NAND2_X1 U950 ( .A1(G113), .A2(n1239), .ZN(n1287) );
NAND3_X1 U951 ( .A1(n1105), .A2(n1248), .A3(n1111), .ZN(n1239) );
NOR2_X1 U952 ( .A1(n1123), .A2(n1288), .ZN(n1111) );
NOR3_X1 U953 ( .A1(n1242), .A2(n1244), .A3(n1075), .ZN(n1248) );
INV_X1 U954 ( .A(n1103), .ZN(n1075) );
NOR2_X1 U955 ( .A1(n1125), .A2(n1116), .ZN(n1103) );
INV_X1 U956 ( .A(n1115), .ZN(n1125) );
NOR2_X1 U957 ( .A1(n1257), .A2(n1256), .ZN(n1105) );
XNOR2_X1 U958 ( .A(G110), .B(n1251), .ZN(G12) );
NAND3_X1 U959 ( .A1(n1106), .A2(n1249), .A3(n1250), .ZN(n1251) );
INV_X1 U960 ( .A(n1089), .ZN(n1250) );
NAND2_X1 U961 ( .A1(n1288), .A2(n1123), .ZN(n1089) );
NAND3_X1 U962 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1123) );
NAND2_X1 U963 ( .A1(n1292), .A2(n1164), .ZN(n1291) );
OR3_X1 U964 ( .A1(n1164), .A2(n1292), .A3(G902), .ZN(n1290) );
NOR2_X1 U965 ( .A1(n1165), .A2(G234), .ZN(n1292) );
INV_X1 U966 ( .A(G217), .ZN(n1165) );
XNOR2_X1 U967 ( .A(n1293), .B(n1294), .ZN(n1164) );
XNOR2_X1 U968 ( .A(KEYINPUT23), .B(n1295), .ZN(n1294) );
INV_X1 U969 ( .A(G119), .ZN(n1295) );
XOR2_X1 U970 ( .A(n1296), .B(n1297), .Z(n1293) );
XOR2_X1 U971 ( .A(n1298), .B(n1299), .Z(n1297) );
XOR2_X1 U972 ( .A(n1300), .B(n1201), .Z(n1299) );
NOR2_X1 U973 ( .A1(G140), .A2(KEYINPUT24), .ZN(n1300) );
XOR2_X1 U974 ( .A(n1301), .B(n1302), .Z(n1298) );
NAND2_X1 U975 ( .A1(KEYINPUT6), .A2(n1252), .ZN(n1302) );
NAND2_X1 U976 ( .A1(n1303), .A2(G221), .ZN(n1301) );
XOR2_X1 U977 ( .A(n1304), .B(n1305), .Z(n1296) );
XNOR2_X1 U978 ( .A(KEYINPUT2), .B(n1306), .ZN(n1305) );
INV_X1 U979 ( .A(G137), .ZN(n1306) );
XNOR2_X1 U980 ( .A(G128), .B(G125), .ZN(n1304) );
NAND2_X1 U981 ( .A1(G217), .A2(G902), .ZN(n1289) );
INV_X1 U982 ( .A(n1280), .ZN(n1288) );
XNOR2_X1 U983 ( .A(n1127), .B(n1307), .ZN(n1280) );
XNOR2_X1 U984 ( .A(KEYINPUT59), .B(n1129), .ZN(n1307) );
INV_X1 U985 ( .A(G472), .ZN(n1129) );
NAND2_X1 U986 ( .A1(n1308), .A2(n1309), .ZN(n1127) );
XOR2_X1 U987 ( .A(n1310), .B(n1311), .Z(n1308) );
XNOR2_X1 U988 ( .A(G101), .B(n1312), .ZN(n1311) );
XNOR2_X1 U989 ( .A(KEYINPUT52), .B(KEYINPUT13), .ZN(n1312) );
XNOR2_X1 U990 ( .A(n1181), .B(n1183), .ZN(n1310) );
NOR2_X1 U991 ( .A1(n1214), .A2(n1313), .ZN(n1183) );
INV_X1 U992 ( .A(G210), .ZN(n1214) );
XNOR2_X1 U993 ( .A(n1314), .B(n1315), .ZN(n1181) );
XOR2_X1 U994 ( .A(n1316), .B(n1317), .Z(n1315) );
NAND2_X1 U995 ( .A1(KEYINPUT57), .A2(n1318), .ZN(n1316) );
XNOR2_X1 U996 ( .A(n1200), .B(n1144), .ZN(n1314) );
INV_X1 U997 ( .A(n1211), .ZN(n1144) );
NOR3_X1 U998 ( .A1(n1113), .A2(n1244), .A3(n1242), .ZN(n1249) );
NAND2_X1 U999 ( .A1(n1087), .A2(n1088), .ZN(n1242) );
NAND2_X1 U1000 ( .A1(G214), .A2(n1319), .ZN(n1088) );
NAND2_X1 U1001 ( .A1(n1320), .A2(n1309), .ZN(n1319) );
NAND2_X1 U1002 ( .A1(n1321), .A2(n1322), .ZN(n1087) );
NAND2_X1 U1003 ( .A1(G210), .A2(n1323), .ZN(n1322) );
NAND2_X1 U1004 ( .A1(n1309), .A2(n1324), .ZN(n1323) );
OR2_X1 U1005 ( .A1(n1320), .A2(n1325), .ZN(n1324) );
NAND3_X1 U1006 ( .A1(n1326), .A2(n1309), .A3(n1325), .ZN(n1321) );
XOR2_X1 U1007 ( .A(n1327), .B(n1209), .Z(n1325) );
NAND2_X1 U1008 ( .A1(n1328), .A2(n1329), .ZN(n1209) );
OR2_X1 U1009 ( .A1(n1160), .A2(KEYINPUT3), .ZN(n1329) );
NAND3_X1 U1010 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n1160) );
NAND2_X1 U1011 ( .A1(n1333), .A2(n1334), .ZN(n1331) );
INV_X1 U1012 ( .A(n1335), .ZN(n1334) );
XOR2_X1 U1013 ( .A(n1336), .B(n1337), .Z(n1333) );
NAND3_X1 U1014 ( .A1(n1336), .A2(n1337), .A3(n1335), .ZN(n1330) );
NAND2_X1 U1015 ( .A1(KEYINPUT3), .A2(n1338), .ZN(n1328) );
NAND2_X1 U1016 ( .A1(n1332), .A2(n1339), .ZN(n1338) );
OR2_X1 U1017 ( .A1(n1335), .A2(n1340), .ZN(n1339) );
NAND2_X1 U1018 ( .A1(n1340), .A2(n1335), .ZN(n1332) );
XNOR2_X1 U1019 ( .A(n1341), .B(G122), .ZN(n1335) );
NAND2_X1 U1020 ( .A1(KEYINPUT0), .A2(n1342), .ZN(n1341) );
XOR2_X1 U1021 ( .A(KEYINPUT49), .B(n1201), .Z(n1342) );
NOR2_X1 U1022 ( .A1(n1337), .A2(n1336), .ZN(n1340) );
XOR2_X1 U1023 ( .A(n1317), .B(n1318), .Z(n1336) );
XNOR2_X1 U1024 ( .A(G119), .B(G113), .ZN(n1317) );
XNOR2_X1 U1025 ( .A(n1343), .B(KEYINPUT36), .ZN(n1337) );
NAND2_X1 U1026 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
NAND2_X1 U1027 ( .A1(n1346), .A2(n1184), .ZN(n1345) );
XOR2_X1 U1028 ( .A(KEYINPUT8), .B(n1347), .Z(n1344) );
NOR2_X1 U1029 ( .A1(n1346), .A2(n1184), .ZN(n1347) );
INV_X1 U1030 ( .A(G101), .ZN(n1184) );
XOR2_X1 U1031 ( .A(n1348), .B(n1213), .Z(n1327) );
XOR2_X1 U1032 ( .A(G125), .B(n1349), .Z(n1213) );
AND2_X1 U1033 ( .A1(n1133), .A2(G224), .ZN(n1349) );
NAND2_X1 U1034 ( .A1(KEYINPUT27), .A2(n1211), .ZN(n1348) );
NAND2_X1 U1035 ( .A1(G210), .A2(G237), .ZN(n1326) );
AND2_X1 U1036 ( .A1(n1350), .A2(n1073), .ZN(n1244) );
NAND3_X1 U1037 ( .A1(n1278), .A2(n1133), .A3(G952), .ZN(n1073) );
NAND4_X1 U1038 ( .A1(G953), .A2(G902), .A3(n1351), .A4(n1159), .ZN(n1350) );
INV_X1 U1039 ( .A(G898), .ZN(n1159) );
XNOR2_X1 U1040 ( .A(KEYINPUT43), .B(n1278), .ZN(n1351) );
NAND2_X1 U1041 ( .A1(G237), .A2(G234), .ZN(n1278) );
INV_X1 U1042 ( .A(n1273), .ZN(n1113) );
NOR2_X1 U1043 ( .A1(n1115), .A2(n1116), .ZN(n1273) );
AND2_X1 U1044 ( .A1(G221), .A2(n1352), .ZN(n1116) );
NAND2_X1 U1045 ( .A1(G234), .A2(n1309), .ZN(n1352) );
XOR2_X1 U1046 ( .A(n1353), .B(G469), .Z(n1115) );
NAND2_X1 U1047 ( .A1(n1354), .A2(n1309), .ZN(n1353) );
XOR2_X1 U1048 ( .A(n1355), .B(n1356), .Z(n1354) );
XOR2_X1 U1049 ( .A(n1357), .B(n1199), .Z(n1356) );
XOR2_X1 U1050 ( .A(G140), .B(n1358), .Z(n1199) );
NOR2_X1 U1051 ( .A1(G953), .A2(n1134), .ZN(n1358) );
INV_X1 U1052 ( .A(G227), .ZN(n1134) );
XOR2_X1 U1053 ( .A(n1359), .B(n1198), .Z(n1357) );
XNOR2_X1 U1054 ( .A(n1360), .B(n1211), .ZN(n1198) );
XNOR2_X1 U1055 ( .A(n1361), .B(n1362), .ZN(n1211) );
XNOR2_X1 U1056 ( .A(G146), .B(KEYINPUT33), .ZN(n1361) );
NAND2_X1 U1057 ( .A1(n1363), .A2(n1364), .ZN(n1360) );
NAND2_X1 U1058 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
XNOR2_X1 U1059 ( .A(G101), .B(KEYINPUT41), .ZN(n1365) );
XOR2_X1 U1060 ( .A(KEYINPUT50), .B(n1367), .Z(n1363) );
NOR2_X1 U1061 ( .A1(n1366), .A2(n1368), .ZN(n1367) );
XNOR2_X1 U1062 ( .A(G101), .B(KEYINPUT16), .ZN(n1368) );
XOR2_X1 U1063 ( .A(n1346), .B(KEYINPUT47), .Z(n1366) );
XNOR2_X1 U1064 ( .A(G104), .B(G107), .ZN(n1346) );
NAND2_X1 U1065 ( .A1(KEYINPUT42), .A2(n1201), .ZN(n1359) );
XOR2_X1 U1066 ( .A(G110), .B(KEYINPUT20), .Z(n1201) );
XOR2_X1 U1067 ( .A(n1369), .B(n1370), .Z(n1355) );
XOR2_X1 U1068 ( .A(KEYINPUT60), .B(KEYINPUT28), .Z(n1370) );
NAND2_X1 U1069 ( .A1(KEYINPUT7), .A2(n1200), .ZN(n1369) );
XNOR2_X1 U1070 ( .A(G134), .B(n1145), .ZN(n1200) );
XOR2_X1 U1071 ( .A(G131), .B(G137), .Z(n1145) );
NOR2_X1 U1072 ( .A1(n1257), .A2(n1279), .ZN(n1106) );
INV_X1 U1073 ( .A(n1256), .ZN(n1279) );
XOR2_X1 U1074 ( .A(n1124), .B(KEYINPUT37), .Z(n1256) );
XOR2_X1 U1075 ( .A(n1371), .B(n1174), .Z(n1124) );
INV_X1 U1076 ( .A(G475), .ZN(n1174) );
NAND2_X1 U1077 ( .A1(n1172), .A2(n1309), .ZN(n1371) );
INV_X1 U1078 ( .A(G902), .ZN(n1309) );
XNOR2_X1 U1079 ( .A(n1372), .B(n1373), .ZN(n1172) );
XOR2_X1 U1080 ( .A(n1374), .B(n1375), .Z(n1373) );
XOR2_X1 U1081 ( .A(G122), .B(G113), .Z(n1375) );
XOR2_X1 U1082 ( .A(G143), .B(G131), .Z(n1374) );
XOR2_X1 U1083 ( .A(n1376), .B(n1377), .Z(n1372) );
NOR2_X1 U1084 ( .A1(n1313), .A2(n1378), .ZN(n1377) );
INV_X1 U1085 ( .A(G214), .ZN(n1378) );
NAND2_X1 U1086 ( .A1(n1133), .A2(n1320), .ZN(n1313) );
INV_X1 U1087 ( .A(G237), .ZN(n1320) );
XNOR2_X1 U1088 ( .A(G104), .B(n1379), .ZN(n1376) );
NOR2_X1 U1089 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
XOR2_X1 U1090 ( .A(n1382), .B(KEYINPUT32), .Z(n1381) );
NAND2_X1 U1091 ( .A1(n1383), .A2(n1252), .ZN(n1382) );
NOR2_X1 U1092 ( .A1(n1252), .A2(n1383), .ZN(n1380) );
XNOR2_X1 U1093 ( .A(G140), .B(n1384), .ZN(n1383) );
NAND2_X1 U1094 ( .A1(n1385), .A2(KEYINPUT1), .ZN(n1384) );
XNOR2_X1 U1095 ( .A(G125), .B(KEYINPUT58), .ZN(n1385) );
INV_X1 U1096 ( .A(G146), .ZN(n1252) );
XOR2_X1 U1097 ( .A(n1386), .B(n1170), .Z(n1257) );
INV_X1 U1098 ( .A(G478), .ZN(n1170) );
OR2_X1 U1099 ( .A1(n1169), .A2(G902), .ZN(n1386) );
XNOR2_X1 U1100 ( .A(n1387), .B(n1388), .ZN(n1169) );
NOR2_X1 U1101 ( .A1(n1389), .A2(n1390), .ZN(n1388) );
XOR2_X1 U1102 ( .A(n1391), .B(KEYINPUT53), .Z(n1390) );
NAND2_X1 U1103 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
NOR2_X1 U1104 ( .A1(n1393), .A2(n1392), .ZN(n1389) );
XNOR2_X1 U1105 ( .A(n1265), .B(n1362), .ZN(n1392) );
XOR2_X1 U1106 ( .A(G128), .B(G143), .Z(n1362) );
INV_X1 U1107 ( .A(G134), .ZN(n1265) );
NAND2_X1 U1108 ( .A1(n1394), .A2(n1395), .ZN(n1393) );
NAND2_X1 U1109 ( .A1(n1396), .A2(n1064), .ZN(n1395) );
XOR2_X1 U1110 ( .A(n1397), .B(KEYINPUT39), .Z(n1394) );
OR2_X1 U1111 ( .A1(n1396), .A2(n1064), .ZN(n1397) );
INV_X1 U1112 ( .A(G107), .ZN(n1064) );
XOR2_X1 U1113 ( .A(n1398), .B(n1318), .Z(n1396) );
XNOR2_X1 U1114 ( .A(G116), .B(KEYINPUT5), .ZN(n1318) );
XNOR2_X1 U1115 ( .A(KEYINPUT40), .B(n1399), .ZN(n1398) );
NOR2_X1 U1116 ( .A1(G122), .A2(KEYINPUT12), .ZN(n1399) );
NAND2_X1 U1117 ( .A1(n1303), .A2(G217), .ZN(n1387) );
AND2_X1 U1118 ( .A1(G234), .A2(n1133), .ZN(n1303) );
INV_X1 U1119 ( .A(G953), .ZN(n1133) );
endmodule


