//Key = 0111111101101010110010000101101110010100011011011110010011000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370;

NAND3_X1 U748 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(G9) );
OR2_X1 U749 ( .A1(n1047), .A2(KEYINPUT35), .ZN(n1046) );
NAND3_X1 U750 ( .A1(KEYINPUT35), .A2(n1047), .A3(n1048), .ZN(n1045) );
NAND2_X1 U751 ( .A1(G107), .A2(n1049), .ZN(n1044) );
NAND2_X1 U752 ( .A1(n1050), .A2(KEYINPUT35), .ZN(n1049) );
XNOR2_X1 U753 ( .A(n1047), .B(KEYINPUT49), .ZN(n1050) );
INV_X1 U754 ( .A(n1051), .ZN(n1047) );
NOR2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(G75) );
NOR4_X1 U756 ( .A1(n1054), .A2(n1055), .A3(G953), .A4(n1056), .ZN(n1053) );
NOR3_X1 U757 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1055) );
NOR2_X1 U758 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U761 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
AND2_X1 U762 ( .A1(n1068), .A2(n1069), .ZN(n1064) );
NOR3_X1 U763 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1060) );
XNOR2_X1 U764 ( .A(n1073), .B(KEYINPUT59), .ZN(n1071) );
NAND3_X1 U765 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1054) );
NAND2_X1 U766 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
XOR2_X1 U767 ( .A(KEYINPUT24), .B(n1079), .Z(n1074) );
NOR2_X1 U768 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR2_X1 U769 ( .A1(n1082), .A2(n1063), .ZN(n1081) );
NOR2_X1 U770 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U771 ( .A1(n1085), .A2(n1057), .ZN(n1084) );
NOR2_X1 U772 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U773 ( .A1(n1088), .A2(n1067), .ZN(n1087) );
NOR2_X1 U774 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR3_X1 U775 ( .A1(n1091), .A2(n1059), .A3(n1092), .ZN(n1090) );
NOR3_X1 U776 ( .A1(n1093), .A2(KEYINPUT21), .A3(n1072), .ZN(n1089) );
NOR4_X1 U777 ( .A1(n1094), .A2(n1059), .A3(n1072), .A4(n1095), .ZN(n1086) );
INV_X1 U778 ( .A(n1096), .ZN(n1059) );
AND3_X1 U779 ( .A1(KEYINPUT21), .A2(n1093), .A3(n1077), .ZN(n1083) );
INV_X1 U780 ( .A(n1097), .ZN(n1093) );
AND3_X1 U781 ( .A1(n1077), .A2(n1096), .A3(n1098), .ZN(n1080) );
NOR3_X1 U782 ( .A1(n1067), .A2(n1072), .A3(n1057), .ZN(n1077) );
NOR3_X1 U783 ( .A1(n1056), .A2(G953), .A3(G952), .ZN(n1052) );
AND4_X1 U784 ( .A1(n1099), .A2(n1069), .A3(n1100), .A4(n1101), .ZN(n1056) );
NOR4_X1 U785 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1101) );
XNOR2_X1 U786 ( .A(n1106), .B(n1107), .ZN(n1104) );
NAND2_X1 U787 ( .A1(KEYINPUT12), .A2(n1108), .ZN(n1106) );
NOR3_X1 U788 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1103) );
NOR2_X1 U789 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
AND3_X1 U790 ( .A1(n1113), .A2(n1112), .A3(KEYINPUT20), .ZN(n1110) );
NOR2_X1 U791 ( .A1(n1114), .A2(KEYINPUT60), .ZN(n1112) );
INV_X1 U792 ( .A(n1115), .ZN(n1114) );
NOR2_X1 U793 ( .A1(KEYINPUT20), .A2(n1115), .ZN(n1109) );
XOR2_X1 U794 ( .A(n1116), .B(G472), .Z(n1100) );
XNOR2_X1 U795 ( .A(n1117), .B(KEYINPUT34), .ZN(n1099) );
XOR2_X1 U796 ( .A(n1118), .B(n1119), .Z(G72) );
NOR2_X1 U797 ( .A1(KEYINPUT58), .A2(n1120), .ZN(n1119) );
XOR2_X1 U798 ( .A(n1121), .B(n1122), .Z(n1120) );
NAND2_X1 U799 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U800 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U801 ( .A1(n1127), .A2(n1128), .ZN(n1121) );
OR2_X1 U802 ( .A1(n1123), .A2(G900), .ZN(n1128) );
XNOR2_X1 U803 ( .A(n1129), .B(n1130), .ZN(n1127) );
XOR2_X1 U804 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U805 ( .A1(KEYINPUT19), .A2(n1133), .ZN(n1132) );
XNOR2_X1 U806 ( .A(n1134), .B(G125), .ZN(n1133) );
NAND4_X1 U807 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1131) );
NAND3_X1 U808 ( .A1(G134), .A2(n1139), .A3(n1140), .ZN(n1138) );
NAND3_X1 U809 ( .A1(n1141), .A2(n1142), .A3(G131), .ZN(n1137) );
NAND2_X1 U810 ( .A1(KEYINPUT47), .A2(n1143), .ZN(n1141) );
OR2_X1 U811 ( .A1(n1144), .A2(n1139), .ZN(n1135) );
INV_X1 U812 ( .A(KEYINPUT47), .ZN(n1139) );
NAND2_X1 U813 ( .A1(G953), .A2(n1145), .ZN(n1118) );
NAND2_X1 U814 ( .A1(G900), .A2(G227), .ZN(n1145) );
XOR2_X1 U815 ( .A(n1146), .B(n1147), .Z(G69) );
NOR2_X1 U816 ( .A1(n1148), .A2(n1123), .ZN(n1147) );
AND2_X1 U817 ( .A1(G898), .A2(G224), .ZN(n1148) );
NAND2_X1 U818 ( .A1(n1149), .A2(n1150), .ZN(n1146) );
NAND2_X1 U819 ( .A1(n1151), .A2(n1123), .ZN(n1150) );
XNOR2_X1 U820 ( .A(n1152), .B(n1153), .ZN(n1151) );
NAND3_X1 U821 ( .A1(G898), .A2(n1153), .A3(G953), .ZN(n1149) );
NOR2_X1 U822 ( .A1(n1154), .A2(n1155), .ZN(G66) );
XOR2_X1 U823 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U824 ( .A1(n1158), .A2(G217), .ZN(n1156) );
NOR3_X1 U825 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(G63) );
AND2_X1 U826 ( .A1(KEYINPUT10), .A2(n1154), .ZN(n1161) );
NOR3_X1 U827 ( .A1(KEYINPUT10), .A2(G953), .A3(G952), .ZN(n1160) );
NOR3_X1 U828 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1159) );
NOR4_X1 U829 ( .A1(n1165), .A2(n1166), .A3(n1107), .A4(n1167), .ZN(n1164) );
NOR2_X1 U830 ( .A1(n1168), .A2(n1169), .ZN(n1163) );
NOR3_X1 U831 ( .A1(n1166), .A2(n1076), .A3(n1107), .ZN(n1168) );
INV_X1 U832 ( .A(KEYINPUT16), .ZN(n1166) );
NOR2_X1 U833 ( .A1(n1154), .A2(n1170), .ZN(G60) );
XOR2_X1 U834 ( .A(n1171), .B(n1172), .Z(n1170) );
NAND2_X1 U835 ( .A1(n1158), .A2(G475), .ZN(n1171) );
XOR2_X1 U836 ( .A(G104), .B(n1173), .Z(G6) );
NOR2_X1 U837 ( .A1(n1066), .A2(n1174), .ZN(n1173) );
NOR2_X1 U838 ( .A1(n1154), .A2(n1175), .ZN(G57) );
XOR2_X1 U839 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U840 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U841 ( .A(n1180), .B(n1181), .Z(n1176) );
XNOR2_X1 U842 ( .A(n1182), .B(n1183), .ZN(n1181) );
NAND2_X1 U843 ( .A1(n1158), .A2(G472), .ZN(n1183) );
NAND2_X1 U844 ( .A1(KEYINPUT41), .A2(n1184), .ZN(n1180) );
NOR2_X1 U845 ( .A1(n1154), .A2(n1185), .ZN(G54) );
XOR2_X1 U846 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U847 ( .A(n1188), .B(n1189), .Z(n1187) );
NOR3_X1 U848 ( .A1(n1167), .A2(KEYINPUT18), .A3(n1113), .ZN(n1189) );
INV_X1 U849 ( .A(n1158), .ZN(n1167) );
XOR2_X1 U850 ( .A(n1190), .B(n1191), .Z(n1186) );
NOR2_X1 U851 ( .A1(KEYINPUT13), .A2(n1192), .ZN(n1191) );
XNOR2_X1 U852 ( .A(n1182), .B(n1193), .ZN(n1192) );
NOR2_X1 U853 ( .A1(KEYINPUT39), .A2(n1194), .ZN(n1193) );
XNOR2_X1 U854 ( .A(n1195), .B(n1196), .ZN(n1194) );
XNOR2_X1 U855 ( .A(n1129), .B(G101), .ZN(n1196) );
NOR3_X1 U856 ( .A1(KEYINPUT26), .A2(n1197), .A3(n1198), .ZN(n1190) );
AND3_X1 U857 ( .A1(KEYINPUT38), .A2(n1134), .A3(G110), .ZN(n1198) );
NOR2_X1 U858 ( .A1(KEYINPUT38), .A2(n1199), .ZN(n1197) );
XNOR2_X1 U859 ( .A(n1134), .B(G110), .ZN(n1199) );
NOR2_X1 U860 ( .A1(n1154), .A2(n1200), .ZN(G51) );
XOR2_X1 U861 ( .A(n1201), .B(n1202), .Z(n1200) );
XOR2_X1 U862 ( .A(n1203), .B(n1204), .Z(n1202) );
NOR2_X1 U863 ( .A1(KEYINPUT46), .A2(n1205), .ZN(n1204) );
NAND2_X1 U864 ( .A1(KEYINPUT25), .A2(n1153), .ZN(n1203) );
XOR2_X1 U865 ( .A(n1206), .B(n1207), .Z(n1201) );
NAND2_X1 U866 ( .A1(n1158), .A2(n1208), .ZN(n1206) );
NOR2_X1 U867 ( .A1(n1209), .A2(n1076), .ZN(n1158) );
AND3_X1 U868 ( .A1(n1152), .A2(n1125), .A3(n1210), .ZN(n1076) );
XOR2_X1 U869 ( .A(n1126), .B(KEYINPUT15), .Z(n1210) );
AND4_X1 U870 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1125) );
NOR4_X1 U871 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
NAND3_X1 U872 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1213) );
XNOR2_X1 U873 ( .A(KEYINPUT55), .B(n1067), .ZN(n1220) );
INV_X1 U874 ( .A(n1073), .ZN(n1067) );
AND4_X1 U875 ( .A1(n1222), .A2(n1051), .A3(n1223), .A4(n1224), .ZN(n1152) );
NOR4_X1 U876 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1224) );
NOR3_X1 U877 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1223) );
AND2_X1 U878 ( .A1(KEYINPUT6), .A2(n1232), .ZN(n1231) );
NOR2_X1 U879 ( .A1(KEYINPUT6), .A2(n1233), .ZN(n1230) );
NAND4_X1 U880 ( .A1(n1078), .A2(n1068), .A3(n1066), .A4(n1234), .ZN(n1233) );
NOR3_X1 U881 ( .A1(n1105), .A2(n1235), .A3(n1063), .ZN(n1078) );
INV_X1 U882 ( .A(n1236), .ZN(n1063) );
NOR2_X1 U883 ( .A1(n1237), .A2(n1066), .ZN(n1229) );
XOR2_X1 U884 ( .A(n1174), .B(KEYINPUT40), .Z(n1237) );
NAND4_X1 U885 ( .A1(n1238), .A2(n1096), .A3(n1068), .A4(n1234), .ZN(n1174) );
NAND4_X1 U886 ( .A1(n1098), .A2(n1096), .A3(n1239), .A4(n1068), .ZN(n1051) );
NOR2_X1 U887 ( .A1(n1123), .A2(G952), .ZN(n1154) );
XNOR2_X1 U888 ( .A(G146), .B(n1211), .ZN(G48) );
NAND2_X1 U889 ( .A1(n1221), .A2(n1240), .ZN(n1211) );
XNOR2_X1 U890 ( .A(G143), .B(n1126), .ZN(G45) );
NAND4_X1 U891 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1117), .ZN(n1126) );
XNOR2_X1 U892 ( .A(G140), .B(n1212), .ZN(G42) );
NAND4_X1 U893 ( .A1(n1219), .A2(n1238), .A3(n1069), .A4(n1068), .ZN(n1212) );
XNOR2_X1 U894 ( .A(n1143), .B(n1218), .ZN(G39) );
AND3_X1 U895 ( .A1(n1236), .A2(n1069), .A3(n1240), .ZN(n1218) );
XNOR2_X1 U896 ( .A(n1217), .B(n1244), .ZN(G36) );
NOR2_X1 U897 ( .A1(G134), .A2(KEYINPUT29), .ZN(n1244) );
AND3_X1 U898 ( .A1(n1069), .A2(n1098), .A3(n1241), .ZN(n1217) );
XNOR2_X1 U899 ( .A(n1140), .B(n1216), .ZN(G33) );
AND3_X1 U900 ( .A1(n1238), .A2(n1069), .A3(n1241), .ZN(n1216) );
AND4_X1 U901 ( .A1(n1245), .A2(n1068), .A3(n1246), .A4(n1247), .ZN(n1241) );
INV_X1 U902 ( .A(n1072), .ZN(n1069) );
NAND2_X1 U903 ( .A1(n1248), .A2(n1091), .ZN(n1072) );
INV_X1 U904 ( .A(n1092), .ZN(n1248) );
XOR2_X1 U905 ( .A(G128), .B(n1215), .Z(G30) );
AND3_X1 U906 ( .A1(n1098), .A2(n1242), .A3(n1240), .ZN(n1215) );
AND4_X1 U907 ( .A1(n1245), .A2(n1068), .A3(n1105), .A4(n1247), .ZN(n1240) );
XNOR2_X1 U908 ( .A(n1249), .B(n1232), .ZN(G3) );
AND3_X1 U909 ( .A1(n1246), .A2(n1245), .A3(n1250), .ZN(n1232) );
XNOR2_X1 U910 ( .A(G125), .B(n1251), .ZN(G27) );
NAND3_X1 U911 ( .A1(n1219), .A2(n1073), .A3(n1221), .ZN(n1251) );
NOR2_X1 U912 ( .A1(n1070), .A2(n1066), .ZN(n1221) );
INV_X1 U913 ( .A(n1238), .ZN(n1070) );
AND2_X1 U914 ( .A1(n1097), .A2(n1247), .ZN(n1219) );
NAND2_X1 U915 ( .A1(n1057), .A2(n1252), .ZN(n1247) );
NAND2_X1 U916 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
XOR2_X1 U917 ( .A(KEYINPUT45), .B(G900), .Z(n1254) );
XOR2_X1 U918 ( .A(n1255), .B(n1228), .Z(G24) );
AND4_X1 U919 ( .A1(n1073), .A2(n1096), .A3(n1256), .A4(n1239), .ZN(n1228) );
NOR2_X1 U920 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NOR2_X1 U921 ( .A1(n1105), .A2(n1245), .ZN(n1096) );
NAND2_X1 U922 ( .A1(KEYINPUT7), .A2(n1259), .ZN(n1255) );
XOR2_X1 U923 ( .A(G119), .B(n1227), .Z(G21) );
AND3_X1 U924 ( .A1(n1260), .A2(n1105), .A3(n1236), .ZN(n1227) );
XOR2_X1 U925 ( .A(n1261), .B(n1226), .Z(G18) );
AND3_X1 U926 ( .A1(n1246), .A2(n1098), .A3(n1260), .ZN(n1226) );
NOR2_X1 U927 ( .A1(n1258), .A2(n1117), .ZN(n1098) );
NAND2_X1 U928 ( .A1(KEYINPUT37), .A2(n1262), .ZN(n1261) );
XNOR2_X1 U929 ( .A(KEYINPUT28), .B(n1263), .ZN(n1262) );
XOR2_X1 U930 ( .A(G113), .B(n1225), .Z(G15) );
AND3_X1 U931 ( .A1(n1246), .A2(n1260), .A3(n1238), .ZN(n1225) );
NOR2_X1 U932 ( .A1(n1257), .A2(n1243), .ZN(n1238) );
INV_X1 U933 ( .A(n1117), .ZN(n1257) );
AND3_X1 U934 ( .A1(n1245), .A2(n1239), .A3(n1073), .ZN(n1260) );
NOR2_X1 U935 ( .A1(n1094), .A2(n1102), .ZN(n1073) );
INV_X1 U936 ( .A(n1095), .ZN(n1102) );
NAND2_X1 U937 ( .A1(n1264), .A2(n1265), .ZN(G12) );
NAND2_X1 U938 ( .A1(G110), .A2(n1222), .ZN(n1265) );
XOR2_X1 U939 ( .A(n1266), .B(KEYINPUT52), .Z(n1264) );
OR2_X1 U940 ( .A1(n1222), .A2(G110), .ZN(n1266) );
NAND2_X1 U941 ( .A1(n1097), .A2(n1250), .ZN(n1222) );
AND3_X1 U942 ( .A1(n1239), .A2(n1068), .A3(n1236), .ZN(n1250) );
NOR2_X1 U943 ( .A1(n1117), .A2(n1243), .ZN(n1236) );
INV_X1 U944 ( .A(n1258), .ZN(n1243) );
NAND2_X1 U945 ( .A1(n1267), .A2(n1268), .ZN(n1258) );
NAND2_X1 U946 ( .A1(n1162), .A2(n1269), .ZN(n1268) );
NAND2_X1 U947 ( .A1(KEYINPUT4), .A2(n1270), .ZN(n1269) );
NAND2_X1 U948 ( .A1(G478), .A2(n1271), .ZN(n1270) );
NAND2_X1 U949 ( .A1(n1272), .A2(n1107), .ZN(n1267) );
INV_X1 U950 ( .A(G478), .ZN(n1107) );
NAND2_X1 U951 ( .A1(n1271), .A2(n1273), .ZN(n1272) );
NAND2_X1 U952 ( .A1(KEYINPUT4), .A2(n1108), .ZN(n1273) );
INV_X1 U953 ( .A(n1162), .ZN(n1108) );
NOR2_X1 U954 ( .A1(n1169), .A2(G902), .ZN(n1162) );
INV_X1 U955 ( .A(n1165), .ZN(n1169) );
XNOR2_X1 U956 ( .A(n1274), .B(n1275), .ZN(n1165) );
XOR2_X1 U957 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U958 ( .A(n1259), .B(G116), .ZN(n1277) );
NOR2_X1 U959 ( .A1(KEYINPUT0), .A2(n1278), .ZN(n1276) );
XNOR2_X1 U960 ( .A(G134), .B(KEYINPUT31), .ZN(n1278) );
XNOR2_X1 U961 ( .A(n1279), .B(n1280), .ZN(n1274) );
XOR2_X1 U962 ( .A(n1281), .B(n1282), .Z(n1280) );
NAND2_X1 U963 ( .A1(G217), .A2(n1283), .ZN(n1282) );
NAND2_X1 U964 ( .A1(KEYINPUT48), .A2(n1048), .ZN(n1281) );
INV_X1 U965 ( .A(G107), .ZN(n1048) );
INV_X1 U966 ( .A(KEYINPUT43), .ZN(n1271) );
XNOR2_X1 U967 ( .A(n1284), .B(G475), .ZN(n1117) );
NAND2_X1 U968 ( .A1(n1172), .A2(n1209), .ZN(n1284) );
XNOR2_X1 U969 ( .A(n1285), .B(n1286), .ZN(n1172) );
XOR2_X1 U970 ( .A(n1287), .B(n1288), .Z(n1286) );
NAND2_X1 U971 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
XNOR2_X1 U972 ( .A(G125), .B(n1291), .ZN(n1290) );
XNOR2_X1 U973 ( .A(KEYINPUT62), .B(KEYINPUT3), .ZN(n1289) );
XOR2_X1 U974 ( .A(n1292), .B(n1293), .Z(n1285) );
XOR2_X1 U975 ( .A(KEYINPUT42), .B(n1294), .Z(n1293) );
NOR2_X1 U976 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
XOR2_X1 U977 ( .A(n1297), .B(KEYINPUT61), .Z(n1296) );
NAND2_X1 U978 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NAND2_X1 U979 ( .A1(G214), .A2(n1300), .ZN(n1299) );
AND3_X1 U980 ( .A1(G214), .A2(G143), .A3(n1300), .ZN(n1295) );
NAND2_X1 U981 ( .A1(KEYINPUT32), .A2(G131), .ZN(n1292) );
AND2_X1 U982 ( .A1(n1094), .A2(n1095), .ZN(n1068) );
NAND2_X1 U983 ( .A1(G221), .A2(n1301), .ZN(n1095) );
XNOR2_X1 U984 ( .A(n1302), .B(n1113), .ZN(n1094) );
INV_X1 U985 ( .A(G469), .ZN(n1113) );
NAND2_X1 U986 ( .A1(KEYINPUT2), .A2(n1115), .ZN(n1302) );
NAND2_X1 U987 ( .A1(n1303), .A2(n1209), .ZN(n1115) );
XOR2_X1 U988 ( .A(n1304), .B(n1305), .Z(n1303) );
XOR2_X1 U989 ( .A(n1306), .B(n1307), .Z(n1305) );
XNOR2_X1 U990 ( .A(n1182), .B(G140), .ZN(n1307) );
XNOR2_X1 U991 ( .A(KEYINPUT50), .B(KEYINPUT22), .ZN(n1306) );
XOR2_X1 U992 ( .A(n1308), .B(n1309), .Z(n1304) );
XNOR2_X1 U993 ( .A(n1310), .B(n1311), .ZN(n1309) );
INV_X1 U994 ( .A(n1195), .ZN(n1310) );
XNOR2_X1 U995 ( .A(n1312), .B(G104), .ZN(n1195) );
NAND2_X1 U996 ( .A1(KEYINPUT14), .A2(G107), .ZN(n1312) );
XOR2_X1 U997 ( .A(n1313), .B(n1188), .Z(n1308) );
AND2_X1 U998 ( .A1(G227), .A2(n1123), .ZN(n1188) );
NAND2_X1 U999 ( .A1(KEYINPUT5), .A2(n1129), .ZN(n1313) );
XOR2_X1 U1000 ( .A(G146), .B(n1279), .Z(n1129) );
AND2_X1 U1001 ( .A1(n1242), .A2(n1234), .ZN(n1239) );
NAND2_X1 U1002 ( .A1(n1057), .A2(n1314), .ZN(n1234) );
NAND2_X1 U1003 ( .A1(n1315), .A2(n1253), .ZN(n1314) );
AND3_X1 U1004 ( .A1(G902), .A2(n1316), .A3(G953), .ZN(n1253) );
XNOR2_X1 U1005 ( .A(G898), .B(KEYINPUT8), .ZN(n1315) );
NAND3_X1 U1006 ( .A1(n1316), .A2(n1123), .A3(G952), .ZN(n1057) );
NAND2_X1 U1007 ( .A1(G237), .A2(n1317), .ZN(n1316) );
INV_X1 U1008 ( .A(n1066), .ZN(n1242) );
NAND2_X1 U1009 ( .A1(n1092), .A2(n1091), .ZN(n1066) );
NAND2_X1 U1010 ( .A1(G214), .A2(n1318), .ZN(n1091) );
XNOR2_X1 U1011 ( .A(n1319), .B(n1208), .ZN(n1092) );
AND2_X1 U1012 ( .A1(G210), .A2(n1318), .ZN(n1208) );
NAND2_X1 U1013 ( .A1(n1320), .A2(n1209), .ZN(n1318) );
INV_X1 U1014 ( .A(G237), .ZN(n1320) );
NAND2_X1 U1015 ( .A1(n1321), .A2(n1209), .ZN(n1319) );
XOR2_X1 U1016 ( .A(n1153), .B(n1322), .Z(n1321) );
XNOR2_X1 U1017 ( .A(KEYINPUT57), .B(n1323), .ZN(n1322) );
NOR2_X1 U1018 ( .A1(KEYINPUT54), .A2(n1324), .ZN(n1323) );
XNOR2_X1 U1019 ( .A(n1207), .B(n1205), .ZN(n1324) );
XNOR2_X1 U1020 ( .A(n1179), .B(n1325), .ZN(n1205) );
INV_X1 U1021 ( .A(G125), .ZN(n1325) );
AND2_X1 U1022 ( .A1(G224), .A2(n1123), .ZN(n1207) );
XOR2_X1 U1023 ( .A(n1326), .B(n1327), .Z(n1153) );
XOR2_X1 U1024 ( .A(n1328), .B(n1329), .Z(n1327) );
XNOR2_X1 U1025 ( .A(G107), .B(KEYINPUT44), .ZN(n1329) );
NAND2_X1 U1026 ( .A1(n1330), .A2(KEYINPUT9), .ZN(n1328) );
XNOR2_X1 U1027 ( .A(G116), .B(G119), .ZN(n1330) );
XOR2_X1 U1028 ( .A(n1288), .B(n1311), .Z(n1326) );
XNOR2_X1 U1029 ( .A(n1249), .B(G110), .ZN(n1311) );
INV_X1 U1030 ( .A(G101), .ZN(n1249) );
XNOR2_X1 U1031 ( .A(G104), .B(n1331), .ZN(n1288) );
XNOR2_X1 U1032 ( .A(n1259), .B(G113), .ZN(n1331) );
INV_X1 U1033 ( .A(G122), .ZN(n1259) );
NOR2_X1 U1034 ( .A1(n1245), .A2(n1246), .ZN(n1097) );
INV_X1 U1035 ( .A(n1105), .ZN(n1246) );
XNOR2_X1 U1036 ( .A(n1332), .B(n1333), .ZN(n1105) );
AND2_X1 U1037 ( .A1(n1301), .A2(G217), .ZN(n1333) );
NAND2_X1 U1038 ( .A1(n1317), .A2(n1209), .ZN(n1301) );
XNOR2_X1 U1039 ( .A(G234), .B(KEYINPUT30), .ZN(n1317) );
NAND2_X1 U1040 ( .A1(n1334), .A2(n1157), .ZN(n1332) );
XOR2_X1 U1041 ( .A(n1335), .B(n1336), .Z(n1157) );
AND2_X1 U1042 ( .A1(n1283), .A2(G221), .ZN(n1336) );
AND2_X1 U1043 ( .A1(G234), .A2(n1123), .ZN(n1283) );
INV_X1 U1044 ( .A(G953), .ZN(n1123) );
XNOR2_X1 U1045 ( .A(n1337), .B(n1143), .ZN(n1335) );
NAND3_X1 U1046 ( .A1(n1338), .A2(n1339), .A3(n1340), .ZN(n1337) );
OR2_X1 U1047 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
NAND2_X1 U1048 ( .A1(n1343), .A2(n1344), .ZN(n1339) );
INV_X1 U1049 ( .A(KEYINPUT17), .ZN(n1344) );
NAND2_X1 U1050 ( .A1(n1345), .A2(n1342), .ZN(n1343) );
XNOR2_X1 U1051 ( .A(KEYINPUT1), .B(n1341), .ZN(n1345) );
NAND2_X1 U1052 ( .A1(KEYINPUT17), .A2(n1346), .ZN(n1338) );
NAND2_X1 U1053 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
OR2_X1 U1054 ( .A1(n1341), .A2(KEYINPUT1), .ZN(n1348) );
NAND3_X1 U1055 ( .A1(n1342), .A2(n1341), .A3(KEYINPUT1), .ZN(n1347) );
XOR2_X1 U1056 ( .A(n1291), .B(n1349), .Z(n1341) );
NOR2_X1 U1057 ( .A1(G125), .A2(KEYINPUT33), .ZN(n1349) );
XNOR2_X1 U1058 ( .A(G146), .B(n1134), .ZN(n1291) );
INV_X1 U1059 ( .A(G140), .ZN(n1134) );
XNOR2_X1 U1060 ( .A(n1350), .B(G110), .ZN(n1342) );
NAND2_X1 U1061 ( .A1(KEYINPUT63), .A2(n1351), .ZN(n1350) );
XOR2_X1 U1062 ( .A(G128), .B(G119), .Z(n1351) );
XNOR2_X1 U1063 ( .A(G902), .B(KEYINPUT36), .ZN(n1334) );
INV_X1 U1064 ( .A(n1235), .ZN(n1245) );
XNOR2_X1 U1065 ( .A(n1352), .B(G472), .ZN(n1235) );
NAND2_X1 U1066 ( .A1(KEYINPUT27), .A2(n1116), .ZN(n1352) );
NAND2_X1 U1067 ( .A1(n1353), .A2(n1209), .ZN(n1116) );
INV_X1 U1068 ( .A(G902), .ZN(n1209) );
XNOR2_X1 U1069 ( .A(n1354), .B(n1184), .ZN(n1353) );
XOR2_X1 U1070 ( .A(n1355), .B(G101), .Z(n1184) );
NAND2_X1 U1071 ( .A1(G210), .A2(n1300), .ZN(n1355) );
NOR2_X1 U1072 ( .A1(G953), .A2(G237), .ZN(n1300) );
NOR2_X1 U1073 ( .A1(n1356), .A2(n1357), .ZN(n1354) );
XOR2_X1 U1074 ( .A(n1358), .B(KEYINPUT53), .Z(n1357) );
NAND2_X1 U1075 ( .A1(n1178), .A2(n1359), .ZN(n1358) );
NOR2_X1 U1076 ( .A1(n1178), .A2(n1359), .ZN(n1356) );
XOR2_X1 U1077 ( .A(n1179), .B(n1360), .Z(n1359) );
NOR2_X1 U1078 ( .A1(n1182), .A2(KEYINPUT23), .ZN(n1360) );
AND3_X1 U1079 ( .A1(n1136), .A2(n1144), .A3(n1361), .ZN(n1182) );
NAND3_X1 U1080 ( .A1(G131), .A2(n1142), .A3(G137), .ZN(n1361) );
INV_X1 U1081 ( .A(G134), .ZN(n1142) );
NAND2_X1 U1082 ( .A1(n1362), .A2(n1143), .ZN(n1144) );
INV_X1 U1083 ( .A(G137), .ZN(n1143) );
XNOR2_X1 U1084 ( .A(G131), .B(G134), .ZN(n1362) );
NAND3_X1 U1085 ( .A1(G134), .A2(n1140), .A3(G137), .ZN(n1136) );
INV_X1 U1086 ( .A(G131), .ZN(n1140) );
NAND2_X1 U1087 ( .A1(n1363), .A2(n1364), .ZN(n1179) );
NAND2_X1 U1088 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
INV_X1 U1089 ( .A(G146), .ZN(n1366) );
XOR2_X1 U1090 ( .A(KEYINPUT56), .B(n1279), .Z(n1365) );
NAND2_X1 U1091 ( .A1(n1279), .A2(G146), .ZN(n1363) );
XNOR2_X1 U1092 ( .A(G128), .B(n1298), .ZN(n1279) );
INV_X1 U1093 ( .A(G143), .ZN(n1298) );
XOR2_X1 U1094 ( .A(n1367), .B(n1368), .Z(n1178) );
NOR2_X1 U1095 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
AND2_X1 U1096 ( .A1(KEYINPUT11), .A2(n1263), .ZN(n1370) );
NOR2_X1 U1097 ( .A1(KEYINPUT51), .A2(n1263), .ZN(n1369) );
INV_X1 U1098 ( .A(G116), .ZN(n1263) );
XNOR2_X1 U1099 ( .A(G113), .B(G119), .ZN(n1367) );
endmodule


