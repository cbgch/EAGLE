//Key = 0100101111001101111000011000101000000010010000010011111001001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242;

XNOR2_X1 U689 ( .A(n945), .B(n946), .ZN(G9) );
NOR2_X1 U690 ( .A1(KEYINPUT21), .A2(n947), .ZN(n946) );
NAND3_X1 U691 ( .A1(n948), .A2(n949), .A3(n950), .ZN(G75) );
NAND2_X1 U692 ( .A1(G952), .A2(n951), .ZN(n950) );
NAND4_X1 U693 ( .A1(n952), .A2(n953), .A3(n954), .A4(n955), .ZN(n951) );
NAND3_X1 U694 ( .A1(n956), .A2(n957), .A3(KEYINPUT25), .ZN(n955) );
NAND4_X1 U695 ( .A1(n958), .A2(n959), .A3(n960), .A4(n961), .ZN(n957) );
NAND2_X1 U696 ( .A1(n962), .A2(n961), .ZN(n954) );
NAND2_X1 U697 ( .A1(n963), .A2(n964), .ZN(n962) );
NAND3_X1 U698 ( .A1(n965), .A2(n966), .A3(n960), .ZN(n964) );
NAND2_X1 U699 ( .A1(n967), .A2(n968), .ZN(n966) );
NAND2_X1 U700 ( .A1(n956), .A2(n969), .ZN(n968) );
NAND2_X1 U701 ( .A1(n970), .A2(n971), .ZN(n969) );
NAND3_X1 U702 ( .A1(n972), .A2(n973), .A3(n974), .ZN(n971) );
NAND2_X1 U703 ( .A1(n959), .A2(n975), .ZN(n967) );
NAND3_X1 U704 ( .A1(n976), .A2(n977), .A3(n978), .ZN(n975) );
NAND2_X1 U705 ( .A1(n956), .A2(n979), .ZN(n978) );
NAND2_X1 U706 ( .A1(n973), .A2(n980), .ZN(n979) );
INV_X1 U707 ( .A(KEYINPUT39), .ZN(n973) );
INV_X1 U708 ( .A(n981), .ZN(n977) );
NAND4_X1 U709 ( .A1(n982), .A2(G214), .A3(n983), .A4(n980), .ZN(n976) );
INV_X1 U710 ( .A(KEYINPUT36), .ZN(n980) );
NAND3_X1 U711 ( .A1(n956), .A2(n984), .A3(n959), .ZN(n963) );
NAND3_X1 U712 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n984) );
NAND2_X1 U713 ( .A1(n960), .A2(n988), .ZN(n987) );
NAND2_X1 U714 ( .A1(n989), .A2(n990), .ZN(n988) );
NAND2_X1 U715 ( .A1(n958), .A2(n991), .ZN(n990) );
INV_X1 U716 ( .A(KEYINPUT25), .ZN(n991) );
NAND2_X1 U717 ( .A1(n965), .A2(n992), .ZN(n986) );
NAND2_X1 U718 ( .A1(n993), .A2(n994), .ZN(n992) );
NAND2_X1 U719 ( .A1(n995), .A2(n996), .ZN(n994) );
OR3_X1 U720 ( .A1(n996), .A2(n997), .A3(n965), .ZN(n985) );
INV_X1 U721 ( .A(KEYINPUT55), .ZN(n996) );
NAND4_X1 U722 ( .A1(n998), .A2(n999), .A3(n1000), .A4(n1001), .ZN(n948) );
NOR4_X1 U723 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n1001) );
NOR2_X1 U724 ( .A1(n1006), .A2(n1007), .ZN(n1003) );
INV_X1 U725 ( .A(KEYINPUT19), .ZN(n1007) );
NOR2_X1 U726 ( .A1(n972), .A2(n974), .ZN(n1006) );
INV_X1 U727 ( .A(n1008), .ZN(n974) );
NOR2_X1 U728 ( .A1(KEYINPUT19), .A2(n959), .ZN(n1002) );
XOR2_X1 U729 ( .A(n1009), .B(n1010), .Z(G72) );
NOR2_X1 U730 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NOR3_X1 U731 ( .A1(n949), .A2(n1013), .A3(n1014), .ZN(n1012) );
NOR2_X1 U732 ( .A1(G953), .A2(n1015), .ZN(n1011) );
XNOR2_X1 U733 ( .A(n952), .B(n1014), .ZN(n1015) );
XOR2_X1 U734 ( .A(n1016), .B(n1017), .Z(n1014) );
XNOR2_X1 U735 ( .A(n1018), .B(G125), .ZN(n1017) );
XNOR2_X1 U736 ( .A(n1019), .B(n1020), .ZN(n1016) );
NAND3_X1 U737 ( .A1(G953), .A2(n1021), .A3(KEYINPUT18), .ZN(n1009) );
NAND2_X1 U738 ( .A1(G900), .A2(G227), .ZN(n1021) );
XOR2_X1 U739 ( .A(n1022), .B(n1023), .Z(G69) );
NOR2_X1 U740 ( .A1(n1024), .A2(n949), .ZN(n1023) );
AND2_X1 U741 ( .A1(G224), .A2(G898), .ZN(n1024) );
NAND2_X1 U742 ( .A1(n1025), .A2(n1026), .ZN(n1022) );
NAND2_X1 U743 ( .A1(n1027), .A2(n949), .ZN(n1026) );
XNOR2_X1 U744 ( .A(n1028), .B(n953), .ZN(n1027) );
NAND3_X1 U745 ( .A1(n1028), .A2(n1029), .A3(G953), .ZN(n1025) );
NOR2_X1 U746 ( .A1(KEYINPUT22), .A2(n1030), .ZN(n1028) );
XOR2_X1 U747 ( .A(n1031), .B(n1032), .Z(n1030) );
NOR2_X1 U748 ( .A1(n1033), .A2(n1034), .ZN(G66) );
XNOR2_X1 U749 ( .A(n1035), .B(n1036), .ZN(n1034) );
XOR2_X1 U750 ( .A(KEYINPUT5), .B(n1037), .Z(n1036) );
NOR2_X1 U751 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR2_X1 U752 ( .A1(n1033), .A2(n1040), .ZN(G63) );
XNOR2_X1 U753 ( .A(n1041), .B(n1042), .ZN(n1040) );
NOR2_X1 U754 ( .A1(n1043), .A2(n1039), .ZN(n1042) );
NOR2_X1 U755 ( .A1(n1033), .A2(n1044), .ZN(G60) );
XNOR2_X1 U756 ( .A(n1045), .B(n1046), .ZN(n1044) );
NOR2_X1 U757 ( .A1(n1047), .A2(n1039), .ZN(n1046) );
XNOR2_X1 U758 ( .A(G475), .B(KEYINPUT46), .ZN(n1047) );
XNOR2_X1 U759 ( .A(G104), .B(n1048), .ZN(G6) );
NOR2_X1 U760 ( .A1(n1033), .A2(n1049), .ZN(G57) );
XOR2_X1 U761 ( .A(n1050), .B(n1051), .Z(n1049) );
XOR2_X1 U762 ( .A(n1052), .B(n1053), .Z(n1051) );
NOR2_X1 U763 ( .A1(KEYINPUT3), .A2(n1054), .ZN(n1053) );
XOR2_X1 U764 ( .A(n1055), .B(n1056), .Z(n1054) );
NOR2_X1 U765 ( .A1(n1057), .A2(n1039), .ZN(n1056) );
NOR2_X1 U766 ( .A1(KEYINPUT61), .A2(n1058), .ZN(n1055) );
XOR2_X1 U767 ( .A(n1059), .B(n1060), .Z(n1058) );
XNOR2_X1 U768 ( .A(KEYINPUT2), .B(n1061), .ZN(n1050) );
INV_X1 U769 ( .A(G101), .ZN(n1061) );
NOR2_X1 U770 ( .A1(n1033), .A2(n1062), .ZN(G54) );
XOR2_X1 U771 ( .A(n1063), .B(n1064), .Z(n1062) );
NOR2_X1 U772 ( .A1(n1065), .A2(n1039), .ZN(n1064) );
NOR2_X1 U773 ( .A1(n1066), .A2(n1067), .ZN(n1063) );
XOR2_X1 U774 ( .A(KEYINPUT11), .B(n1068), .Z(n1067) );
NOR2_X1 U775 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
INV_X1 U776 ( .A(n1071), .ZN(n1069) );
NOR2_X1 U777 ( .A1(n1072), .A2(n1071), .ZN(n1066) );
XNOR2_X1 U778 ( .A(n1019), .B(n1073), .ZN(n1071) );
XOR2_X1 U779 ( .A(n1074), .B(n1075), .Z(n1019) );
XOR2_X1 U780 ( .A(n1070), .B(KEYINPUT15), .Z(n1072) );
XNOR2_X1 U781 ( .A(n1076), .B(n1077), .ZN(n1070) );
NAND2_X1 U782 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NAND2_X1 U783 ( .A1(G110), .A2(n1018), .ZN(n1079) );
XOR2_X1 U784 ( .A(KEYINPUT62), .B(n1080), .Z(n1078) );
NOR2_X1 U785 ( .A1(G110), .A2(n1018), .ZN(n1080) );
NOR2_X1 U786 ( .A1(n1033), .A2(n1081), .ZN(G51) );
XOR2_X1 U787 ( .A(n1082), .B(n1083), .Z(n1081) );
XOR2_X1 U788 ( .A(n1084), .B(n1085), .Z(n1083) );
NOR2_X1 U789 ( .A1(n1086), .A2(n1039), .ZN(n1085) );
NAND2_X1 U790 ( .A1(G902), .A2(n1087), .ZN(n1039) );
NAND2_X1 U791 ( .A1(n952), .A2(n953), .ZN(n1087) );
AND4_X1 U792 ( .A1(n1048), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n953) );
AND4_X1 U793 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n945), .ZN(n1090) );
NAND3_X1 U794 ( .A1(n1094), .A2(n1095), .A3(n960), .ZN(n945) );
NAND2_X1 U795 ( .A1(n1096), .A2(n1097), .ZN(n1089) );
NAND2_X1 U796 ( .A1(n1098), .A2(n997), .ZN(n1097) );
XNOR2_X1 U797 ( .A(KEYINPUT8), .B(n993), .ZN(n1098) );
NAND3_X1 U798 ( .A1(n960), .A2(n1094), .A3(n958), .ZN(n1048) );
AND4_X1 U799 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n952) );
NOR4_X1 U800 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1102) );
AND2_X1 U801 ( .A1(n1107), .A2(n1108), .ZN(n1101) );
NAND2_X1 U802 ( .A1(n1109), .A2(n956), .ZN(n1100) );
XOR2_X1 U803 ( .A(n1110), .B(KEYINPUT53), .Z(n1109) );
NAND2_X1 U804 ( .A1(n1111), .A2(n1112), .ZN(n1099) );
XNOR2_X1 U805 ( .A(KEYINPUT20), .B(n1004), .ZN(n1112) );
NOR2_X1 U806 ( .A1(n1113), .A2(n1114), .ZN(n1084) );
XOR2_X1 U807 ( .A(n1115), .B(KEYINPUT16), .Z(n1114) );
NAND2_X1 U808 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NOR2_X1 U809 ( .A1(n1117), .A2(n1116), .ZN(n1113) );
XNOR2_X1 U810 ( .A(n1118), .B(n1119), .ZN(n1116) );
NAND2_X1 U811 ( .A1(KEYINPUT47), .A2(n1120), .ZN(n1118) );
AND2_X1 U812 ( .A1(n1121), .A2(G953), .ZN(n1033) );
XNOR2_X1 U813 ( .A(G952), .B(KEYINPUT29), .ZN(n1121) );
XOR2_X1 U814 ( .A(n1107), .B(n1122), .Z(G48) );
NAND2_X1 U815 ( .A1(KEYINPUT28), .A2(G146), .ZN(n1122) );
NAND3_X1 U816 ( .A1(n958), .A2(n981), .A3(n1123), .ZN(n1107) );
XNOR2_X1 U817 ( .A(n1124), .B(n1125), .ZN(G45) );
NAND2_X1 U818 ( .A1(KEYINPUT51), .A2(n1108), .ZN(n1124) );
NAND4_X1 U819 ( .A1(n1126), .A2(n1127), .A3(n981), .A4(n1005), .ZN(n1108) );
XNOR2_X1 U820 ( .A(n1018), .B(n1128), .ZN(G42) );
NOR2_X1 U821 ( .A1(n1004), .A2(n1110), .ZN(n1128) );
NAND4_X1 U822 ( .A1(n958), .A2(n995), .A3(n1129), .A4(n1130), .ZN(n1110) );
INV_X1 U823 ( .A(G140), .ZN(n1018) );
XNOR2_X1 U824 ( .A(n1131), .B(n1106), .ZN(G39) );
AND3_X1 U825 ( .A1(n956), .A2(n965), .A3(n1123), .ZN(n1106) );
XNOR2_X1 U826 ( .A(G134), .B(n1132), .ZN(G36) );
NAND2_X1 U827 ( .A1(n1111), .A2(n956), .ZN(n1132) );
AND2_X1 U828 ( .A1(n1127), .A2(n1095), .ZN(n1111) );
XOR2_X1 U829 ( .A(G131), .B(n1105), .Z(G33) );
AND3_X1 U830 ( .A1(n958), .A2(n956), .A3(n1127), .ZN(n1105) );
AND3_X1 U831 ( .A1(n1129), .A2(n1130), .A3(n1133), .ZN(n1127) );
INV_X1 U832 ( .A(n1004), .ZN(n956) );
NAND2_X1 U833 ( .A1(n982), .A2(n1134), .ZN(n1004) );
NAND2_X1 U834 ( .A1(G214), .A2(n983), .ZN(n1134) );
XOR2_X1 U835 ( .A(G128), .B(n1104), .Z(G30) );
AND3_X1 U836 ( .A1(n1095), .A2(n981), .A3(n1123), .ZN(n1104) );
AND4_X1 U837 ( .A1(n1135), .A2(n1129), .A3(n1136), .A4(n1130), .ZN(n1123) );
XNOR2_X1 U838 ( .A(G101), .B(n1137), .ZN(G3) );
NAND2_X1 U839 ( .A1(n1096), .A2(n1133), .ZN(n1137) );
NAND2_X1 U840 ( .A1(n1138), .A2(n1139), .ZN(G27) );
NAND2_X1 U841 ( .A1(n1103), .A2(n1120), .ZN(n1139) );
XOR2_X1 U842 ( .A(KEYINPUT24), .B(n1140), .Z(n1138) );
NOR2_X1 U843 ( .A1(n1103), .A2(n1120), .ZN(n1140) );
AND4_X1 U844 ( .A1(n981), .A2(n1130), .A3(n995), .A4(n1141), .ZN(n1103) );
AND2_X1 U845 ( .A1(n959), .A2(n958), .ZN(n1141) );
NAND2_X1 U846 ( .A1(n1142), .A2(n1143), .ZN(n1130) );
NAND4_X1 U847 ( .A1(G953), .A2(G902), .A3(n1013), .A4(n961), .ZN(n1143) );
XOR2_X1 U848 ( .A(G900), .B(KEYINPUT60), .Z(n1013) );
XNOR2_X1 U849 ( .A(G122), .B(n1093), .ZN(G24) );
NAND4_X1 U850 ( .A1(n1144), .A2(n960), .A3(n1126), .A4(n1005), .ZN(n1093) );
AND2_X1 U851 ( .A1(n1145), .A2(n1000), .ZN(n960) );
XOR2_X1 U852 ( .A(n998), .B(KEYINPUT59), .Z(n1145) );
XNOR2_X1 U853 ( .A(G119), .B(n1088), .ZN(G21) );
NAND4_X1 U854 ( .A1(n1135), .A2(n1144), .A3(n965), .A4(n1136), .ZN(n1088) );
XNOR2_X1 U855 ( .A(G116), .B(n1092), .ZN(G18) );
NAND3_X1 U856 ( .A1(n1133), .A2(n1095), .A3(n1144), .ZN(n1092) );
INV_X1 U857 ( .A(n989), .ZN(n1095) );
NAND2_X1 U858 ( .A1(n1146), .A2(n1005), .ZN(n989) );
XNOR2_X1 U859 ( .A(KEYINPUT12), .B(n999), .ZN(n1146) );
XNOR2_X1 U860 ( .A(G113), .B(n1091), .ZN(G15) );
NAND3_X1 U861 ( .A1(n1133), .A2(n958), .A3(n1144), .ZN(n1091) );
AND3_X1 U862 ( .A1(n981), .A2(n1147), .A3(n959), .ZN(n1144) );
NOR2_X1 U863 ( .A1(n1008), .A2(n972), .ZN(n959) );
INV_X1 U864 ( .A(n993), .ZN(n1133) );
NAND2_X1 U865 ( .A1(n998), .A2(n1136), .ZN(n993) );
XNOR2_X1 U866 ( .A(G110), .B(n1148), .ZN(G12) );
NAND2_X1 U867 ( .A1(n1096), .A2(n995), .ZN(n1148) );
INV_X1 U868 ( .A(n997), .ZN(n995) );
NAND2_X1 U869 ( .A1(n1135), .A2(n1000), .ZN(n997) );
INV_X1 U870 ( .A(n1136), .ZN(n1000) );
XOR2_X1 U871 ( .A(n1149), .B(n1057), .Z(n1136) );
INV_X1 U872 ( .A(G472), .ZN(n1057) );
NAND2_X1 U873 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XOR2_X1 U874 ( .A(n1152), .B(n1153), .Z(n1150) );
XOR2_X1 U875 ( .A(n1059), .B(n1154), .Z(n1153) );
XOR2_X1 U876 ( .A(n1155), .B(n1156), .Z(n1059) );
XOR2_X1 U877 ( .A(KEYINPUT52), .B(n1157), .Z(n1156) );
XNOR2_X1 U878 ( .A(n1075), .B(n1158), .ZN(n1155) );
XOR2_X1 U879 ( .A(G137), .B(n1159), .Z(n1075) );
XNOR2_X1 U880 ( .A(n1052), .B(KEYINPUT37), .ZN(n1152) );
NOR3_X1 U881 ( .A1(G237), .A2(G953), .A3(n1086), .ZN(n1052) );
XOR2_X1 U882 ( .A(n998), .B(KEYINPUT63), .Z(n1135) );
XNOR2_X1 U883 ( .A(n1160), .B(n1038), .ZN(n998) );
NAND2_X1 U884 ( .A1(G217), .A2(n1161), .ZN(n1038) );
NAND2_X1 U885 ( .A1(n1035), .A2(n1151), .ZN(n1160) );
XNOR2_X1 U886 ( .A(n1162), .B(n1163), .ZN(n1035) );
XOR2_X1 U887 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U888 ( .A1(n1166), .A2(n1167), .ZN(n1164) );
OR2_X1 U889 ( .A1(n1168), .A2(G110), .ZN(n1167) );
XOR2_X1 U890 ( .A(n1169), .B(KEYINPUT49), .Z(n1166) );
NAND2_X1 U891 ( .A1(G110), .A2(n1168), .ZN(n1169) );
XOR2_X1 U892 ( .A(G119), .B(n1170), .Z(n1168) );
XOR2_X1 U893 ( .A(n1171), .B(n1172), .Z(n1162) );
XNOR2_X1 U894 ( .A(n1131), .B(G125), .ZN(n1172) );
NAND2_X1 U895 ( .A1(G221), .A2(n1173), .ZN(n1171) );
AND2_X1 U896 ( .A1(n1094), .A2(n965), .ZN(n1096) );
NAND2_X1 U897 ( .A1(n1174), .A2(n1175), .ZN(n965) );
NAND2_X1 U898 ( .A1(n958), .A2(n1176), .ZN(n1175) );
NOR2_X1 U899 ( .A1(n1005), .A2(n999), .ZN(n958) );
OR3_X1 U900 ( .A1(n1126), .A2(n1005), .A3(n1176), .ZN(n1174) );
INV_X1 U901 ( .A(KEYINPUT12), .ZN(n1176) );
XOR2_X1 U902 ( .A(n1177), .B(n1043), .Z(n1005) );
INV_X1 U903 ( .A(G478), .ZN(n1043) );
NAND2_X1 U904 ( .A1(n1041), .A2(n1151), .ZN(n1177) );
XNOR2_X1 U905 ( .A(n1178), .B(n1179), .ZN(n1041) );
XOR2_X1 U906 ( .A(n1159), .B(n1180), .Z(n1179) );
XNOR2_X1 U907 ( .A(n1181), .B(n1182), .ZN(n1180) );
NOR2_X1 U908 ( .A1(G107), .A2(KEYINPUT43), .ZN(n1182) );
NAND2_X1 U909 ( .A1(KEYINPUT4), .A2(n1183), .ZN(n1181) );
XOR2_X1 U910 ( .A(G134), .B(n1170), .Z(n1159) );
XOR2_X1 U911 ( .A(n1184), .B(n1185), .Z(n1178) );
AND2_X1 U912 ( .A1(G217), .A2(n1173), .ZN(n1185) );
AND2_X1 U913 ( .A1(G234), .A2(n949), .ZN(n1173) );
XNOR2_X1 U914 ( .A(G122), .B(n1186), .ZN(n1184) );
NOR2_X1 U915 ( .A1(KEYINPUT0), .A2(n1125), .ZN(n1186) );
INV_X1 U916 ( .A(n999), .ZN(n1126) );
XNOR2_X1 U917 ( .A(n1187), .B(n1188), .ZN(n999) );
XOR2_X1 U918 ( .A(KEYINPUT50), .B(G475), .Z(n1188) );
NAND2_X1 U919 ( .A1(n1045), .A2(n1151), .ZN(n1187) );
XNOR2_X1 U920 ( .A(n1189), .B(n1190), .ZN(n1045) );
XOR2_X1 U921 ( .A(G104), .B(n1191), .Z(n1190) );
XOR2_X1 U922 ( .A(G122), .B(G113), .Z(n1191) );
XOR2_X1 U923 ( .A(n1165), .B(n1192), .Z(n1189) );
XNOR2_X1 U924 ( .A(n1193), .B(n1194), .ZN(n1192) );
NOR2_X1 U925 ( .A1(KEYINPUT34), .A2(n1195), .ZN(n1194) );
XNOR2_X1 U926 ( .A(n1196), .B(n1020), .ZN(n1195) );
NAND2_X1 U927 ( .A1(KEYINPUT57), .A2(n1197), .ZN(n1196) );
XNOR2_X1 U928 ( .A(G143), .B(n1198), .ZN(n1197) );
NAND4_X1 U929 ( .A1(n1199), .A2(G214), .A3(n1200), .A4(n949), .ZN(n1198) );
INV_X1 U930 ( .A(G237), .ZN(n1200) );
XNOR2_X1 U931 ( .A(KEYINPUT42), .B(KEYINPUT27), .ZN(n1199) );
NAND2_X1 U932 ( .A1(KEYINPUT1), .A2(G125), .ZN(n1193) );
XNOR2_X1 U933 ( .A(G146), .B(G140), .ZN(n1165) );
AND3_X1 U934 ( .A1(n1129), .A2(n1147), .A3(n981), .ZN(n1094) );
NOR2_X1 U935 ( .A1(n982), .A2(n1201), .ZN(n981) );
AND2_X1 U936 ( .A1(G214), .A2(n983), .ZN(n1201) );
XOR2_X1 U937 ( .A(n1202), .B(n1203), .Z(n982) );
NOR2_X1 U938 ( .A1(n1086), .A2(n1204), .ZN(n1203) );
XNOR2_X1 U939 ( .A(KEYINPUT56), .B(n983), .ZN(n1204) );
NAND2_X1 U940 ( .A1(n1205), .A2(n1151), .ZN(n983) );
XNOR2_X1 U941 ( .A(G237), .B(KEYINPUT48), .ZN(n1205) );
INV_X1 U942 ( .A(G210), .ZN(n1086) );
NAND2_X1 U943 ( .A1(n1206), .A2(n1151), .ZN(n1202) );
XOR2_X1 U944 ( .A(n1207), .B(n1208), .Z(n1206) );
XNOR2_X1 U945 ( .A(n1117), .B(n1209), .ZN(n1208) );
XNOR2_X1 U946 ( .A(KEYINPUT32), .B(n1120), .ZN(n1209) );
INV_X1 U947 ( .A(G125), .ZN(n1120) );
NAND2_X1 U948 ( .A1(G224), .A2(n949), .ZN(n1117) );
XNOR2_X1 U949 ( .A(n1082), .B(n1119), .ZN(n1207) );
XOR2_X1 U950 ( .A(n1158), .B(n1170), .Z(n1119) );
XNOR2_X1 U951 ( .A(n1210), .B(G146), .ZN(n1158) );
NAND2_X1 U952 ( .A1(KEYINPUT13), .A2(n1125), .ZN(n1210) );
XNOR2_X1 U953 ( .A(n1031), .B(n1211), .ZN(n1082) );
NOR2_X1 U954 ( .A1(KEYINPUT35), .A2(n1032), .ZN(n1211) );
XNOR2_X1 U955 ( .A(n1212), .B(n1213), .ZN(n1032) );
XOR2_X1 U956 ( .A(KEYINPUT38), .B(G122), .Z(n1213) );
NAND2_X1 U957 ( .A1(KEYINPUT30), .A2(n1214), .ZN(n1212) );
XOR2_X1 U958 ( .A(n1215), .B(n1216), .Z(n1031) );
XNOR2_X1 U959 ( .A(n947), .B(G104), .ZN(n1216) );
XNOR2_X1 U960 ( .A(n1157), .B(n1217), .ZN(n1215) );
NOR2_X1 U961 ( .A1(G101), .A2(KEYINPUT45), .ZN(n1217) );
XOR2_X1 U962 ( .A(G113), .B(n1218), .Z(n1157) );
XNOR2_X1 U963 ( .A(G119), .B(n1183), .ZN(n1218) );
INV_X1 U964 ( .A(G116), .ZN(n1183) );
NAND2_X1 U965 ( .A1(n1219), .A2(n1142), .ZN(n1147) );
NAND3_X1 U966 ( .A1(G952), .A2(n949), .A3(n1220), .ZN(n1142) );
XOR2_X1 U967 ( .A(n961), .B(KEYINPUT10), .Z(n1220) );
XOR2_X1 U968 ( .A(n1221), .B(KEYINPUT40), .Z(n1219) );
NAND4_X1 U969 ( .A1(G953), .A2(G902), .A3(n1222), .A4(n961), .ZN(n1221) );
NAND2_X1 U970 ( .A1(G237), .A2(G234), .ZN(n961) );
INV_X1 U971 ( .A(n1029), .ZN(n1222) );
XOR2_X1 U972 ( .A(G898), .B(KEYINPUT58), .Z(n1029) );
INV_X1 U973 ( .A(n970), .ZN(n1129) );
NAND2_X1 U974 ( .A1(n1223), .A2(n1008), .ZN(n970) );
XOR2_X1 U975 ( .A(n1224), .B(n1065), .Z(n1008) );
INV_X1 U976 ( .A(G469), .ZN(n1065) );
NAND2_X1 U977 ( .A1(n1225), .A2(n1151), .ZN(n1224) );
XOR2_X1 U978 ( .A(n1226), .B(n1227), .Z(n1225) );
XOR2_X1 U979 ( .A(n1228), .B(n1229), .Z(n1227) );
XNOR2_X1 U980 ( .A(n1131), .B(G134), .ZN(n1229) );
INV_X1 U981 ( .A(G137), .ZN(n1131) );
NOR2_X1 U982 ( .A1(KEYINPUT31), .A2(n1230), .ZN(n1228) );
XNOR2_X1 U983 ( .A(n1231), .B(n1214), .ZN(n1230) );
INV_X1 U984 ( .A(G110), .ZN(n1214) );
NAND2_X1 U985 ( .A1(KEYINPUT9), .A2(G140), .ZN(n1231) );
XNOR2_X1 U986 ( .A(n1073), .B(n1232), .ZN(n1226) );
XOR2_X1 U987 ( .A(n1077), .B(n1233), .Z(n1232) );
NAND2_X1 U988 ( .A1(n1234), .A2(KEYINPUT6), .ZN(n1233) );
XOR2_X1 U989 ( .A(n1074), .B(n1170), .Z(n1234) );
XOR2_X1 U990 ( .A(G128), .B(KEYINPUT44), .Z(n1170) );
NAND2_X1 U991 ( .A1(n1235), .A2(n1236), .ZN(n1074) );
NAND2_X1 U992 ( .A1(G146), .A2(n1125), .ZN(n1236) );
XOR2_X1 U993 ( .A(KEYINPUT54), .B(n1237), .Z(n1235) );
NOR2_X1 U994 ( .A1(G146), .A2(n1125), .ZN(n1237) );
INV_X1 U995 ( .A(G143), .ZN(n1125) );
NAND2_X1 U996 ( .A1(G227), .A2(n949), .ZN(n1077) );
INV_X1 U997 ( .A(G953), .ZN(n949) );
XNOR2_X1 U998 ( .A(n1238), .B(n1239), .ZN(n1073) );
XNOR2_X1 U999 ( .A(KEYINPUT33), .B(n947), .ZN(n1239) );
INV_X1 U1000 ( .A(G107), .ZN(n947) );
XNOR2_X1 U1001 ( .A(n1154), .B(n1240), .ZN(n1238) );
NOR2_X1 U1002 ( .A1(G104), .A2(KEYINPUT26), .ZN(n1240) );
XOR2_X1 U1003 ( .A(G101), .B(n1060), .Z(n1154) );
XNOR2_X1 U1004 ( .A(n1241), .B(KEYINPUT23), .ZN(n1060) );
NAND2_X1 U1005 ( .A1(KEYINPUT7), .A2(n1020), .ZN(n1241) );
XNOR2_X1 U1006 ( .A(G131), .B(KEYINPUT14), .ZN(n1020) );
XOR2_X1 U1007 ( .A(KEYINPUT41), .B(n972), .Z(n1223) );
AND2_X1 U1008 ( .A1(G221), .A2(n1161), .ZN(n972) );
NAND2_X1 U1009 ( .A1(n1242), .A2(n1151), .ZN(n1161) );
INV_X1 U1010 ( .A(G902), .ZN(n1151) );
XNOR2_X1 U1011 ( .A(G234), .B(KEYINPUT17), .ZN(n1242) );
endmodule


