//Key = 0001001100101001110000101110011011001010001101010010100010110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389;

NAND2_X1 U762 ( .A1(n1060), .A2(n1061), .ZN(G9) );
NAND2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND2_X1 U765 ( .A1(KEYINPUT31), .A2(n1066), .ZN(n1065) );
OR2_X1 U766 ( .A1(n1067), .A2(KEYINPUT31), .ZN(n1064) );
NAND2_X1 U767 ( .A1(G107), .A2(n1067), .ZN(n1060) );
NOR2_X1 U768 ( .A1(n1068), .A2(KEYINPUT2), .ZN(n1067) );
INV_X1 U769 ( .A(n1066), .ZN(n1068) );
NOR2_X1 U770 ( .A1(n1069), .A2(n1070), .ZN(G75) );
NOR3_X1 U771 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1070) );
NOR2_X1 U772 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR2_X1 U776 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR3_X1 U777 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1082) );
NOR2_X1 U778 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR2_X1 U780 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR2_X1 U781 ( .A1(KEYINPUT39), .A2(n1093), .ZN(n1089) );
NOR2_X1 U782 ( .A1(n1094), .A2(n1095), .ZN(n1085) );
XOR2_X1 U783 ( .A(KEYINPUT33), .B(n1096), .Z(n1095) );
AND2_X1 U784 ( .A1(n1097), .A2(n1096), .ZN(n1084) );
NOR3_X1 U785 ( .A1(n1098), .A2(n1088), .A3(n1099), .ZN(n1080) );
INV_X1 U786 ( .A(n1100), .ZN(n1088) );
INV_X1 U787 ( .A(n1096), .ZN(n1098) );
NOR3_X1 U788 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1076) );
NAND3_X1 U789 ( .A1(n1104), .A2(n1100), .A3(n1105), .ZN(n1101) );
XOR2_X1 U790 ( .A(KEYINPUT14), .B(n1106), .Z(n1105) );
XOR2_X1 U791 ( .A(KEYINPUT61), .B(n1096), .Z(n1104) );
NAND3_X1 U792 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1071) );
NAND4_X1 U793 ( .A1(n1106), .A2(n1110), .A3(n1100), .A4(n1111), .ZN(n1109) );
NAND2_X1 U794 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND3_X1 U795 ( .A1(n1114), .A2(n1075), .A3(KEYINPUT39), .ZN(n1113) );
INV_X1 U796 ( .A(n1115), .ZN(n1075) );
NAND2_X1 U797 ( .A1(n1096), .A2(n1116), .ZN(n1112) );
NAND2_X1 U798 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
INV_X1 U800 ( .A(n1079), .ZN(n1106) );
NOR3_X1 U801 ( .A1(n1121), .A2(G953), .A3(G952), .ZN(n1069) );
INV_X1 U802 ( .A(n1107), .ZN(n1121) );
NAND4_X1 U803 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1107) );
NOR4_X1 U804 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n1125) );
XOR2_X1 U805 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U806 ( .A(n1132), .B(n1133), .Z(n1128) );
NOR3_X1 U807 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1124) );
INV_X1 U808 ( .A(n1102), .ZN(n1135) );
NOR3_X1 U809 ( .A1(n1137), .A2(G902), .A3(n1138), .ZN(n1134) );
XNOR2_X1 U810 ( .A(n1139), .B(n1140), .ZN(n1122) );
NOR2_X1 U811 ( .A1(G469), .A2(KEYINPUT37), .ZN(n1140) );
XOR2_X1 U812 ( .A(n1141), .B(n1142), .Z(G72) );
NOR2_X1 U813 ( .A1(n1143), .A2(n1108), .ZN(n1142) );
NOR2_X1 U814 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U815 ( .A(KEYINPUT32), .B(G227), .Z(n1145) );
NAND2_X1 U816 ( .A1(n1146), .A2(n1147), .ZN(n1141) );
NAND2_X1 U817 ( .A1(n1148), .A2(n1108), .ZN(n1147) );
XOR2_X1 U818 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U819 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
OR3_X1 U820 ( .A1(n1144), .A2(n1150), .A3(n1108), .ZN(n1146) );
XNOR2_X1 U821 ( .A(n1153), .B(n1154), .ZN(n1150) );
XOR2_X1 U822 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U823 ( .A(G140), .B(G125), .Z(n1156) );
XOR2_X1 U824 ( .A(n1157), .B(n1158), .Z(n1153) );
XOR2_X1 U825 ( .A(n1159), .B(n1160), .Z(G69) );
XOR2_X1 U826 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U827 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U828 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U829 ( .A1(KEYINPUT46), .A2(n1167), .ZN(n1166) );
XOR2_X1 U830 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U831 ( .A1(n1170), .A2(KEYINPUT48), .ZN(n1168) );
NOR2_X1 U832 ( .A1(G898), .A2(n1108), .ZN(n1163) );
NOR2_X1 U833 ( .A1(n1171), .A2(n1172), .ZN(n1161) );
XOR2_X1 U834 ( .A(KEYINPUT27), .B(G953), .Z(n1172) );
NOR2_X1 U835 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
XOR2_X1 U836 ( .A(KEYINPUT34), .B(n1175), .Z(n1174) );
NOR2_X1 U837 ( .A1(n1176), .A2(n1108), .ZN(n1159) );
AND2_X1 U838 ( .A1(G224), .A2(G898), .ZN(n1176) );
NOR2_X1 U839 ( .A1(n1177), .A2(n1178), .ZN(G66) );
XOR2_X1 U840 ( .A(n1179), .B(n1180), .Z(n1178) );
NAND2_X1 U841 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
NOR2_X1 U842 ( .A1(n1177), .A2(n1183), .ZN(G63) );
XOR2_X1 U843 ( .A(n1184), .B(n1185), .Z(n1183) );
NAND2_X1 U844 ( .A1(n1181), .A2(G478), .ZN(n1184) );
NOR3_X1 U845 ( .A1(n1177), .A2(n1186), .A3(n1187), .ZN(G60) );
NOR4_X1 U846 ( .A1(n1188), .A2(n1189), .A3(KEYINPUT18), .A4(n1130), .ZN(n1187) );
NOR2_X1 U847 ( .A1(n1190), .A2(n1191), .ZN(n1186) );
NOR3_X1 U848 ( .A1(n1189), .A2(n1192), .A3(n1130), .ZN(n1191) );
INV_X1 U849 ( .A(G475), .ZN(n1130) );
NOR2_X1 U850 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
INV_X1 U851 ( .A(KEYINPUT18), .ZN(n1194) );
INV_X1 U852 ( .A(n1188), .ZN(n1190) );
NAND2_X1 U853 ( .A1(KEYINPUT16), .A2(n1193), .ZN(n1188) );
XOR2_X1 U854 ( .A(G104), .B(n1195), .Z(G6) );
NOR2_X1 U855 ( .A1(n1093), .A2(n1196), .ZN(n1195) );
NOR2_X1 U856 ( .A1(n1177), .A2(n1197), .ZN(G57) );
NOR2_X1 U857 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U858 ( .A(KEYINPUT51), .B(n1200), .Z(n1199) );
AND2_X1 U859 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NOR2_X1 U860 ( .A1(n1201), .A2(n1202), .ZN(n1198) );
XNOR2_X1 U861 ( .A(n1203), .B(n1204), .ZN(n1202) );
XOR2_X1 U862 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U863 ( .A(n1207), .B(KEYINPUT8), .Z(n1206) );
NAND2_X1 U864 ( .A1(KEYINPUT25), .A2(n1208), .ZN(n1207) );
NAND2_X1 U865 ( .A1(n1181), .A2(G472), .ZN(n1205) );
XNOR2_X1 U866 ( .A(n1209), .B(n1210), .ZN(n1203) );
NOR2_X1 U867 ( .A1(n1177), .A2(n1211), .ZN(G54) );
XOR2_X1 U868 ( .A(n1212), .B(n1213), .Z(n1211) );
XNOR2_X1 U869 ( .A(n1214), .B(n1215), .ZN(n1213) );
NAND2_X1 U870 ( .A1(n1181), .A2(G469), .ZN(n1214) );
XOR2_X1 U871 ( .A(n1216), .B(KEYINPUT30), .Z(n1212) );
NAND2_X1 U872 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NAND2_X1 U873 ( .A1(G140), .A2(n1219), .ZN(n1218) );
XOR2_X1 U874 ( .A(n1220), .B(KEYINPUT5), .Z(n1217) );
NAND2_X1 U875 ( .A1(G110), .A2(n1221), .ZN(n1220) );
NOR2_X1 U876 ( .A1(n1177), .A2(n1222), .ZN(G51) );
XOR2_X1 U877 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U878 ( .A(n1225), .B(n1226), .Z(n1224) );
NAND2_X1 U879 ( .A1(KEYINPUT42), .A2(n1227), .ZN(n1226) );
NAND2_X1 U880 ( .A1(n1181), .A2(G210), .ZN(n1225) );
INV_X1 U881 ( .A(n1189), .ZN(n1181) );
NAND2_X1 U882 ( .A1(G902), .A2(n1073), .ZN(n1189) );
OR4_X1 U883 ( .A1(n1228), .A2(n1173), .A3(n1152), .A4(n1175), .ZN(n1073) );
INV_X1 U884 ( .A(n1229), .ZN(n1175) );
NAND4_X1 U885 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1152) );
NAND3_X1 U886 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1231) );
XOR2_X1 U887 ( .A(n1117), .B(KEYINPUT29), .Z(n1236) );
NAND4_X1 U888 ( .A1(n1237), .A2(n1097), .A3(n1238), .A4(n1239), .ZN(n1230) );
OR2_X1 U889 ( .A1(n1234), .A2(KEYINPUT4), .ZN(n1239) );
NAND2_X1 U890 ( .A1(KEYINPUT4), .A2(n1240), .ZN(n1238) );
NAND3_X1 U891 ( .A1(n1241), .A2(n1099), .A3(n1096), .ZN(n1240) );
NAND4_X1 U892 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1173) );
AND4_X1 U893 ( .A1(n1246), .A2(n1247), .A3(n1066), .A4(n1248), .ZN(n1245) );
NAND4_X1 U894 ( .A1(n1115), .A2(n1235), .A3(n1249), .A4(n1250), .ZN(n1066) );
NAND2_X1 U895 ( .A1(n1251), .A2(n1114), .ZN(n1244) );
XOR2_X1 U896 ( .A(n1196), .B(KEYINPUT3), .Z(n1251) );
NAND4_X1 U897 ( .A1(n1097), .A2(n1115), .A3(n1252), .A4(n1250), .ZN(n1196) );
XNOR2_X1 U898 ( .A(n1151), .B(KEYINPUT10), .ZN(n1228) );
NAND4_X1 U899 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1151) );
XOR2_X1 U900 ( .A(n1257), .B(n1258), .Z(n1223) );
NOR2_X1 U901 ( .A1(n1108), .A2(G952), .ZN(n1177) );
XNOR2_X1 U902 ( .A(G146), .B(n1253), .ZN(G48) );
NAND2_X1 U903 ( .A1(n1259), .A2(n1097), .ZN(n1253) );
XNOR2_X1 U904 ( .A(n1254), .B(n1260), .ZN(G45) );
NOR2_X1 U905 ( .A1(KEYINPUT23), .A2(n1261), .ZN(n1260) );
NAND3_X1 U906 ( .A1(n1237), .A2(n1249), .A3(n1262), .ZN(n1254) );
AND3_X1 U907 ( .A1(n1263), .A2(n1241), .A3(n1126), .ZN(n1262) );
XNOR2_X1 U908 ( .A(n1255), .B(n1264), .ZN(G42) );
NOR2_X1 U909 ( .A1(KEYINPUT35), .A2(n1221), .ZN(n1264) );
INV_X1 U910 ( .A(G140), .ZN(n1221) );
NAND2_X1 U911 ( .A1(n1234), .A2(n1265), .ZN(n1255) );
XNOR2_X1 U912 ( .A(G137), .B(n1256), .ZN(G39) );
NAND3_X1 U913 ( .A1(n1266), .A2(n1100), .A3(n1234), .ZN(n1256) );
INV_X1 U914 ( .A(n1267), .ZN(n1234) );
XNOR2_X1 U915 ( .A(G134), .B(n1268), .ZN(G36) );
NAND2_X1 U916 ( .A1(n1269), .A2(n1235), .ZN(n1268) );
XOR2_X1 U917 ( .A(n1270), .B(n1271), .Z(G33) );
XNOR2_X1 U918 ( .A(G131), .B(KEYINPUT44), .ZN(n1271) );
NAND2_X1 U919 ( .A1(n1269), .A2(n1097), .ZN(n1270) );
NOR2_X1 U920 ( .A1(n1267), .A2(n1117), .ZN(n1269) );
INV_X1 U921 ( .A(n1237), .ZN(n1117) );
NAND3_X1 U922 ( .A1(n1252), .A2(n1241), .A3(n1096), .ZN(n1267) );
NOR2_X1 U923 ( .A1(n1092), .A2(n1136), .ZN(n1096) );
INV_X1 U924 ( .A(n1099), .ZN(n1252) );
XOR2_X1 U925 ( .A(n1272), .B(n1232), .Z(G30) );
NAND2_X1 U926 ( .A1(n1259), .A2(n1235), .ZN(n1232) );
AND3_X1 U927 ( .A1(n1249), .A2(n1241), .A3(n1266), .ZN(n1259) );
XOR2_X1 U928 ( .A(G101), .B(n1273), .Z(G3) );
NOR2_X1 U929 ( .A1(KEYINPUT41), .A2(n1229), .ZN(n1273) );
NAND2_X1 U930 ( .A1(n1237), .A2(n1274), .ZN(n1229) );
XOR2_X1 U931 ( .A(n1275), .B(n1233), .Z(G27) );
NAND4_X1 U932 ( .A1(n1265), .A2(n1110), .A3(n1114), .A4(n1241), .ZN(n1233) );
NAND2_X1 U933 ( .A1(n1079), .A2(n1276), .ZN(n1241) );
NAND4_X1 U934 ( .A1(n1277), .A2(G953), .A3(G902), .A4(n1278), .ZN(n1276) );
XOR2_X1 U935 ( .A(n1144), .B(KEYINPUT57), .Z(n1277) );
INV_X1 U936 ( .A(G900), .ZN(n1144) );
AND3_X1 U937 ( .A1(n1119), .A2(n1120), .A3(n1097), .ZN(n1265) );
XNOR2_X1 U938 ( .A(G122), .B(n1242), .ZN(G24) );
NAND4_X1 U939 ( .A1(n1279), .A2(n1115), .A3(n1263), .A4(n1126), .ZN(n1242) );
NOR2_X1 U940 ( .A1(n1127), .A2(n1120), .ZN(n1115) );
XOR2_X1 U941 ( .A(n1280), .B(n1243), .Z(G21) );
NAND3_X1 U942 ( .A1(n1279), .A2(n1100), .A3(n1266), .ZN(n1243) );
AND2_X1 U943 ( .A1(n1120), .A2(n1127), .ZN(n1266) );
INV_X1 U944 ( .A(n1119), .ZN(n1127) );
XOR2_X1 U945 ( .A(n1281), .B(n1247), .Z(G18) );
NAND3_X1 U946 ( .A1(n1237), .A2(n1235), .A3(n1279), .ZN(n1247) );
INV_X1 U947 ( .A(n1094), .ZN(n1235) );
NAND2_X1 U948 ( .A1(n1282), .A2(n1126), .ZN(n1094) );
XOR2_X1 U949 ( .A(KEYINPUT21), .B(n1283), .Z(n1282) );
XOR2_X1 U950 ( .A(n1284), .B(n1246), .Z(G15) );
NAND3_X1 U951 ( .A1(n1237), .A2(n1097), .A3(n1279), .ZN(n1246) );
AND3_X1 U952 ( .A1(n1114), .A2(n1250), .A3(n1110), .ZN(n1279) );
INV_X1 U953 ( .A(n1083), .ZN(n1110) );
NAND2_X1 U954 ( .A1(n1285), .A2(n1102), .ZN(n1083) );
INV_X1 U955 ( .A(n1093), .ZN(n1114) );
NOR2_X1 U956 ( .A1(n1120), .A2(n1119), .ZN(n1237) );
NAND3_X1 U957 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(G12) );
OR2_X1 U958 ( .A1(n1248), .A2(KEYINPUT45), .ZN(n1288) );
NAND3_X1 U959 ( .A1(KEYINPUT45), .A2(n1248), .A3(G110), .ZN(n1287) );
NAND2_X1 U960 ( .A1(n1289), .A2(n1219), .ZN(n1286) );
NAND2_X1 U961 ( .A1(n1290), .A2(KEYINPUT45), .ZN(n1289) );
XOR2_X1 U962 ( .A(n1248), .B(KEYINPUT63), .Z(n1290) );
NAND3_X1 U963 ( .A1(n1119), .A2(n1120), .A3(n1274), .ZN(n1248) );
AND3_X1 U964 ( .A1(n1100), .A2(n1250), .A3(n1249), .ZN(n1274) );
NOR2_X1 U965 ( .A1(n1099), .A2(n1093), .ZN(n1249) );
NAND2_X1 U966 ( .A1(n1291), .A2(n1092), .ZN(n1093) );
NAND3_X1 U967 ( .A1(n1292), .A2(n1293), .A3(n1123), .ZN(n1092) );
NAND2_X1 U968 ( .A1(G210), .A2(n1294), .ZN(n1123) );
NAND2_X1 U969 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
NAND2_X1 U970 ( .A1(n1137), .A2(n1297), .ZN(n1296) );
NAND2_X1 U971 ( .A1(KEYINPUT49), .A2(n1298), .ZN(n1293) );
OR3_X1 U972 ( .A1(n1138), .A2(KEYINPUT49), .A3(n1298), .ZN(n1292) );
OR2_X1 U973 ( .A1(n1137), .A2(G902), .ZN(n1298) );
XNOR2_X1 U974 ( .A(n1299), .B(n1300), .ZN(n1137) );
NOR2_X1 U975 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NOR3_X1 U976 ( .A1(KEYINPUT22), .A2(n1209), .A3(n1303), .ZN(n1302) );
NOR2_X1 U977 ( .A1(n1258), .A2(n1304), .ZN(n1301) );
INV_X1 U978 ( .A(KEYINPUT22), .ZN(n1304) );
XNOR2_X1 U979 ( .A(n1303), .B(n1209), .ZN(n1258) );
XOR2_X1 U980 ( .A(n1275), .B(KEYINPUT11), .Z(n1303) );
XNOR2_X1 U981 ( .A(n1257), .B(n1227), .ZN(n1299) );
NAND2_X1 U982 ( .A1(G224), .A2(n1108), .ZN(n1227) );
XOR2_X1 U983 ( .A(n1305), .B(n1306), .Z(n1257) );
XNOR2_X1 U984 ( .A(n1170), .B(n1165), .ZN(n1306) );
XOR2_X1 U985 ( .A(n1307), .B(n1308), .Z(n1165) );
XOR2_X1 U986 ( .A(KEYINPUT12), .B(G122), .Z(n1308) );
NAND2_X1 U987 ( .A1(KEYINPUT7), .A2(n1219), .ZN(n1307) );
AND2_X1 U988 ( .A1(n1309), .A2(n1310), .ZN(n1170) );
NAND2_X1 U989 ( .A1(n1311), .A2(n1284), .ZN(n1310) );
XOR2_X1 U990 ( .A(n1280), .B(n1312), .Z(n1311) );
NAND2_X1 U991 ( .A1(n1313), .A2(n1314), .ZN(n1309) );
XOR2_X1 U992 ( .A(KEYINPUT54), .B(G113), .Z(n1314) );
XOR2_X1 U993 ( .A(n1312), .B(G119), .Z(n1313) );
NAND2_X1 U994 ( .A1(KEYINPUT59), .A2(n1281), .ZN(n1312) );
AND2_X1 U995 ( .A1(G210), .A2(n1297), .ZN(n1138) );
XOR2_X1 U996 ( .A(KEYINPUT52), .B(n1136), .Z(n1291) );
INV_X1 U997 ( .A(n1091), .ZN(n1136) );
NAND2_X1 U998 ( .A1(G214), .A2(n1315), .ZN(n1091) );
OR2_X1 U999 ( .A1(n1297), .A2(G902), .ZN(n1315) );
XOR2_X1 U1000 ( .A(G237), .B(KEYINPUT62), .Z(n1297) );
NAND2_X1 U1001 ( .A1(n1103), .A2(n1102), .ZN(n1099) );
NAND2_X1 U1002 ( .A1(G221), .A2(n1316), .ZN(n1102) );
INV_X1 U1003 ( .A(n1285), .ZN(n1103) );
XOR2_X1 U1004 ( .A(n1139), .B(G469), .Z(n1285) );
NAND2_X1 U1005 ( .A1(n1317), .A2(n1295), .ZN(n1139) );
XOR2_X1 U1006 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1007 ( .A(KEYINPUT24), .B(G140), .Z(n1319) );
XOR2_X1 U1008 ( .A(n1219), .B(n1215), .Z(n1318) );
XNOR2_X1 U1009 ( .A(n1320), .B(n1321), .ZN(n1215) );
XNOR2_X1 U1010 ( .A(n1155), .B(n1208), .ZN(n1321) );
XOR2_X1 U1011 ( .A(G128), .B(n1322), .Z(n1155) );
NOR2_X1 U1012 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1013 ( .A(n1325), .B(KEYINPUT50), .Z(n1324) );
NAND2_X1 U1014 ( .A1(n1326), .A2(n1261), .ZN(n1325) );
XOR2_X1 U1015 ( .A(KEYINPUT53), .B(G146), .Z(n1326) );
NOR2_X1 U1016 ( .A1(G146), .A2(n1261), .ZN(n1323) );
XOR2_X1 U1017 ( .A(n1327), .B(n1169), .Z(n1320) );
INV_X1 U1018 ( .A(n1305), .ZN(n1169) );
XOR2_X1 U1019 ( .A(n1328), .B(n1329), .Z(n1305) );
XOR2_X1 U1020 ( .A(n1330), .B(G107), .Z(n1328) );
XOR2_X1 U1021 ( .A(n1331), .B(KEYINPUT38), .Z(n1327) );
NAND2_X1 U1022 ( .A1(G227), .A2(n1108), .ZN(n1331) );
INV_X1 U1023 ( .A(G110), .ZN(n1219) );
NAND2_X1 U1024 ( .A1(n1079), .A2(n1332), .ZN(n1250) );
NAND4_X1 U1025 ( .A1(G953), .A2(G902), .A3(n1278), .A4(n1333), .ZN(n1332) );
INV_X1 U1026 ( .A(G898), .ZN(n1333) );
NAND3_X1 U1027 ( .A1(n1278), .A2(n1108), .A3(G952), .ZN(n1079) );
NAND2_X1 U1028 ( .A1(G234), .A2(G237), .ZN(n1278) );
NAND2_X1 U1029 ( .A1(n1334), .A2(n1335), .ZN(n1100) );
OR3_X1 U1030 ( .A1(n1263), .A2(n1126), .A3(KEYINPUT21), .ZN(n1335) );
NAND2_X1 U1031 ( .A1(KEYINPUT21), .A2(n1097), .ZN(n1334) );
NOR2_X1 U1032 ( .A1(n1126), .A2(n1283), .ZN(n1097) );
INV_X1 U1033 ( .A(n1263), .ZN(n1283) );
XOR2_X1 U1034 ( .A(n1131), .B(n1336), .Z(n1263) );
NOR2_X1 U1035 ( .A1(G475), .A2(KEYINPUT0), .ZN(n1336) );
NAND2_X1 U1036 ( .A1(n1193), .A2(n1295), .ZN(n1131) );
XNOR2_X1 U1037 ( .A(n1337), .B(n1338), .ZN(n1193) );
XOR2_X1 U1038 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1039 ( .A(n1341), .B(n1342), .Z(n1340) );
NOR2_X1 U1040 ( .A1(KEYINPUT40), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1041 ( .A(n1344), .B(n1345), .Z(n1343) );
XOR2_X1 U1042 ( .A(n1346), .B(G125), .Z(n1344) );
NAND2_X1 U1043 ( .A1(KEYINPUT26), .A2(G140), .ZN(n1346) );
NAND3_X1 U1044 ( .A1(n1347), .A2(n1108), .A3(G214), .ZN(n1341) );
NAND2_X1 U1045 ( .A1(KEYINPUT36), .A2(n1330), .ZN(n1339) );
INV_X1 U1046 ( .A(G104), .ZN(n1330) );
XOR2_X1 U1047 ( .A(n1348), .B(n1349), .Z(n1337) );
XOR2_X1 U1048 ( .A(G122), .B(G113), .Z(n1349) );
XOR2_X1 U1049 ( .A(G131), .B(n1261), .Z(n1348) );
INV_X1 U1050 ( .A(G143), .ZN(n1261) );
XNOR2_X1 U1051 ( .A(n1350), .B(G478), .ZN(n1126) );
NAND2_X1 U1052 ( .A1(n1185), .A2(n1295), .ZN(n1350) );
XOR2_X1 U1053 ( .A(n1351), .B(n1352), .Z(n1185) );
XOR2_X1 U1054 ( .A(n1063), .B(n1353), .Z(n1352) );
NAND2_X1 U1055 ( .A1(n1354), .A2(KEYINPUT6), .ZN(n1353) );
XOR2_X1 U1056 ( .A(n1281), .B(G122), .Z(n1354) );
INV_X1 U1057 ( .A(G107), .ZN(n1063) );
XOR2_X1 U1058 ( .A(n1355), .B(n1356), .Z(n1351) );
NOR2_X1 U1059 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
XOR2_X1 U1060 ( .A(KEYINPUT1), .B(n1359), .Z(n1358) );
NOR2_X1 U1061 ( .A1(G134), .A2(n1360), .ZN(n1359) );
AND2_X1 U1062 ( .A1(n1360), .A2(G134), .ZN(n1357) );
NAND2_X1 U1063 ( .A1(n1361), .A2(G217), .ZN(n1355) );
XNOR2_X1 U1064 ( .A(n1362), .B(n1182), .ZN(n1120) );
INV_X1 U1065 ( .A(n1132), .ZN(n1182) );
NAND2_X1 U1066 ( .A1(G217), .A2(n1316), .ZN(n1132) );
NAND2_X1 U1067 ( .A1(G234), .A2(n1295), .ZN(n1316) );
NAND2_X1 U1068 ( .A1(KEYINPUT15), .A2(n1363), .ZN(n1362) );
INV_X1 U1069 ( .A(n1133), .ZN(n1363) );
NAND2_X1 U1070 ( .A1(n1180), .A2(n1295), .ZN(n1133) );
XNOR2_X1 U1071 ( .A(n1364), .B(n1365), .ZN(n1180) );
XNOR2_X1 U1072 ( .A(n1345), .B(n1366), .ZN(n1365) );
XOR2_X1 U1073 ( .A(n1367), .B(n1368), .Z(n1366) );
NOR2_X1 U1074 ( .A1(KEYINPUT13), .A2(n1275), .ZN(n1368) );
INV_X1 U1075 ( .A(G125), .ZN(n1275) );
NAND2_X1 U1076 ( .A1(G221), .A2(n1361), .ZN(n1367) );
AND2_X1 U1077 ( .A1(G234), .A2(n1108), .ZN(n1361) );
XOR2_X1 U1078 ( .A(G146), .B(KEYINPUT17), .Z(n1345) );
XOR2_X1 U1079 ( .A(n1369), .B(n1370), .Z(n1364) );
XOR2_X1 U1080 ( .A(G140), .B(n1371), .Z(n1370) );
NOR2_X1 U1081 ( .A1(KEYINPUT20), .A2(G137), .ZN(n1371) );
NAND2_X1 U1082 ( .A1(n1372), .A2(n1373), .ZN(n1369) );
OR2_X1 U1083 ( .A1(n1374), .A2(G110), .ZN(n1373) );
XOR2_X1 U1084 ( .A(n1375), .B(KEYINPUT60), .Z(n1372) );
NAND2_X1 U1085 ( .A1(G110), .A2(n1374), .ZN(n1375) );
XOR2_X1 U1086 ( .A(n1280), .B(n1272), .Z(n1374) );
XOR2_X1 U1087 ( .A(n1376), .B(G472), .Z(n1119) );
NAND2_X1 U1088 ( .A1(n1377), .A2(n1295), .ZN(n1376) );
INV_X1 U1089 ( .A(G902), .ZN(n1295) );
XNOR2_X1 U1090 ( .A(n1378), .B(n1201), .ZN(n1377) );
XNOR2_X1 U1091 ( .A(n1379), .B(n1329), .ZN(n1201) );
XOR2_X1 U1092 ( .A(G101), .B(KEYINPUT43), .Z(n1329) );
NAND3_X1 U1093 ( .A1(n1347), .A2(n1108), .A3(G210), .ZN(n1379) );
INV_X1 U1094 ( .A(G953), .ZN(n1108) );
XNOR2_X1 U1095 ( .A(G237), .B(KEYINPUT28), .ZN(n1347) );
NAND3_X1 U1096 ( .A1(n1380), .A2(n1381), .A3(n1382), .ZN(n1378) );
OR2_X1 U1097 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
NAND3_X1 U1098 ( .A1(n1385), .A2(n1383), .A3(n1210), .ZN(n1381) );
INV_X1 U1099 ( .A(KEYINPUT9), .ZN(n1383) );
OR2_X1 U1100 ( .A1(n1210), .A2(n1385), .ZN(n1380) );
AND2_X1 U1101 ( .A1(KEYINPUT56), .A2(n1384), .ZN(n1385) );
XNOR2_X1 U1102 ( .A(n1209), .B(n1208), .ZN(n1384) );
XNOR2_X1 U1103 ( .A(n1386), .B(n1157), .ZN(n1208) );
XNOR2_X1 U1104 ( .A(G131), .B(G137), .ZN(n1157) );
NAND2_X1 U1105 ( .A1(KEYINPUT58), .A2(n1158), .ZN(n1386) );
XOR2_X1 U1106 ( .A(G134), .B(KEYINPUT47), .Z(n1158) );
XOR2_X1 U1107 ( .A(G146), .B(n1360), .Z(n1209) );
XNOR2_X1 U1108 ( .A(n1272), .B(G143), .ZN(n1360) );
INV_X1 U1109 ( .A(G128), .ZN(n1272) );
XNOR2_X1 U1110 ( .A(n1284), .B(n1387), .ZN(n1210) );
NOR2_X1 U1111 ( .A1(KEYINPUT55), .A2(n1388), .ZN(n1387) );
XOR2_X1 U1112 ( .A(n1281), .B(n1389), .Z(n1388) );
NOR2_X1 U1113 ( .A1(KEYINPUT19), .A2(n1280), .ZN(n1389) );
INV_X1 U1114 ( .A(G119), .ZN(n1280) );
INV_X1 U1115 ( .A(G116), .ZN(n1281) );
INV_X1 U1116 ( .A(G113), .ZN(n1284) );
endmodule


