//Key = 0100101101111100101101111101111100001011110101000011100010011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450;

XOR2_X1 U797 ( .A(G107), .B(n1101), .Z(G9) );
NOR3_X1 U798 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
XNOR2_X1 U799 ( .A(n1105), .B(KEYINPUT15), .ZN(n1103) );
NOR2_X1 U800 ( .A1(n1106), .A2(n1107), .ZN(G75) );
NOR3_X1 U801 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1107) );
NAND3_X1 U802 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1108) );
NAND2_X1 U803 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
NAND2_X1 U804 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND3_X1 U805 ( .A1(n1118), .A2(n1119), .A3(n1105), .ZN(n1117) );
NAND2_X1 U806 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U807 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U808 ( .A1(n1124), .A2(n1104), .ZN(n1123) );
NAND2_X1 U809 ( .A1(n1125), .A2(n1126), .ZN(n1120) );
NAND2_X1 U810 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U811 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
INV_X1 U812 ( .A(n1131), .ZN(n1127) );
NAND3_X1 U813 ( .A1(n1122), .A2(n1132), .A3(n1125), .ZN(n1116) );
NAND2_X1 U814 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U815 ( .A1(n1118), .A2(n1135), .ZN(n1134) );
OR2_X1 U816 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U817 ( .A1(n1105), .A2(n1138), .ZN(n1133) );
NAND2_X1 U818 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NAND2_X1 U819 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
INV_X1 U820 ( .A(n1143), .ZN(n1114) );
AND3_X1 U821 ( .A1(n1113), .A2(n1112), .A3(n1144), .ZN(n1106) );
XNOR2_X1 U822 ( .A(n1109), .B(KEYINPUT1), .ZN(n1144) );
INV_X1 U823 ( .A(G952), .ZN(n1109) );
NAND4_X1 U824 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1112) );
NOR4_X1 U825 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1148) );
XNOR2_X1 U826 ( .A(G469), .B(n1153), .ZN(n1152) );
XOR2_X1 U827 ( .A(G478), .B(n1154), .Z(n1151) );
XNOR2_X1 U828 ( .A(n1155), .B(n1156), .ZN(n1149) );
NAND2_X1 U829 ( .A1(KEYINPUT16), .A2(n1157), .ZN(n1155) );
NOR2_X1 U830 ( .A1(n1129), .A2(n1141), .ZN(n1147) );
XNOR2_X1 U831 ( .A(n1158), .B(n1159), .ZN(n1146) );
NAND2_X1 U832 ( .A1(KEYINPUT43), .A2(n1160), .ZN(n1159) );
XOR2_X1 U833 ( .A(n1161), .B(n1162), .Z(n1145) );
NAND2_X1 U834 ( .A1(KEYINPUT51), .A2(n1163), .ZN(n1162) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(G72) );
NOR2_X1 U836 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
AND2_X1 U837 ( .A1(G227), .A2(G900), .ZN(n1166) );
NAND2_X1 U838 ( .A1(n1168), .A2(n1169), .ZN(n1164) );
NAND2_X1 U839 ( .A1(n1170), .A2(n1167), .ZN(n1169) );
XNOR2_X1 U840 ( .A(n1171), .B(n1172), .ZN(n1170) );
NOR2_X1 U841 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XNOR2_X1 U842 ( .A(n1175), .B(KEYINPUT30), .ZN(n1173) );
NAND3_X1 U843 ( .A1(G900), .A2(n1171), .A3(G953), .ZN(n1168) );
XNOR2_X1 U844 ( .A(n1176), .B(n1177), .ZN(n1171) );
XOR2_X1 U845 ( .A(n1178), .B(n1179), .Z(n1176) );
NAND2_X1 U846 ( .A1(n1180), .A2(KEYINPUT25), .ZN(n1178) );
XNOR2_X1 U847 ( .A(n1181), .B(n1182), .ZN(n1180) );
XNOR2_X1 U848 ( .A(n1183), .B(n1184), .ZN(n1182) );
NOR2_X1 U849 ( .A1(G137), .A2(KEYINPUT49), .ZN(n1184) );
XOR2_X1 U850 ( .A(n1185), .B(n1186), .Z(G69) );
NOR3_X1 U851 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1186) );
NOR3_X1 U852 ( .A1(n1167), .A2(KEYINPUT26), .A3(n1190), .ZN(n1189) );
NOR3_X1 U853 ( .A1(G953), .A2(KEYINPUT48), .A3(n1191), .ZN(n1188) );
NOR2_X1 U854 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U855 ( .A(n1194), .B(KEYINPUT55), .Z(n1192) );
AND3_X1 U856 ( .A1(KEYINPUT26), .A2(G953), .A3(n1190), .ZN(n1187) );
AND2_X1 U857 ( .A1(G898), .A2(G224), .ZN(n1190) );
NAND3_X1 U858 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1185) );
NAND2_X1 U859 ( .A1(G953), .A2(n1198), .ZN(n1197) );
NAND2_X1 U860 ( .A1(n1199), .A2(n1200), .ZN(n1196) );
NAND2_X1 U861 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
XNOR2_X1 U862 ( .A(KEYINPUT38), .B(n1203), .ZN(n1199) );
NAND3_X1 U863 ( .A1(n1204), .A2(n1202), .A3(n1201), .ZN(n1195) );
XOR2_X1 U864 ( .A(n1205), .B(KEYINPUT53), .Z(n1201) );
NOR2_X1 U865 ( .A1(n1206), .A2(n1207), .ZN(G66) );
XNOR2_X1 U866 ( .A(n1208), .B(n1209), .ZN(n1207) );
NOR2_X1 U867 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NOR2_X1 U868 ( .A1(n1206), .A2(n1212), .ZN(G63) );
NOR3_X1 U869 ( .A1(n1154), .A2(n1213), .A3(n1214), .ZN(n1212) );
AND4_X1 U870 ( .A1(n1215), .A2(KEYINPUT59), .A3(G478), .A4(n1216), .ZN(n1214) );
NOR2_X1 U871 ( .A1(n1217), .A2(n1215), .ZN(n1213) );
AND3_X1 U872 ( .A1(KEYINPUT59), .A2(n1110), .A3(G478), .ZN(n1217) );
INV_X1 U873 ( .A(n1218), .ZN(n1110) );
NOR2_X1 U874 ( .A1(n1206), .A2(n1219), .ZN(G60) );
NOR3_X1 U875 ( .A1(n1158), .A2(n1220), .A3(n1221), .ZN(n1219) );
AND3_X1 U876 ( .A1(n1222), .A2(G475), .A3(n1216), .ZN(n1221) );
NOR2_X1 U877 ( .A1(n1223), .A2(n1222), .ZN(n1220) );
NOR2_X1 U878 ( .A1(n1218), .A2(n1160), .ZN(n1223) );
XNOR2_X1 U879 ( .A(G104), .B(n1224), .ZN(G6) );
NAND3_X1 U880 ( .A1(n1225), .A2(n1105), .A3(n1226), .ZN(n1224) );
NOR3_X1 U881 ( .A1(n1206), .A2(n1227), .A3(n1228), .ZN(G57) );
NOR3_X1 U882 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1228) );
NOR2_X1 U883 ( .A1(n1232), .A2(n1233), .ZN(n1227) );
INV_X1 U884 ( .A(n1229), .ZN(n1233) );
XNOR2_X1 U885 ( .A(n1234), .B(n1235), .ZN(n1229) );
NOR2_X1 U886 ( .A1(G101), .A2(KEYINPUT5), .ZN(n1235) );
NOR2_X1 U887 ( .A1(n1230), .A2(n1231), .ZN(n1232) );
XNOR2_X1 U888 ( .A(n1236), .B(KEYINPUT42), .ZN(n1231) );
NAND2_X1 U889 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NOR2_X1 U890 ( .A1(n1238), .A2(n1237), .ZN(n1230) );
NAND2_X1 U891 ( .A1(n1216), .A2(G472), .ZN(n1238) );
NOR2_X1 U892 ( .A1(n1206), .A2(n1239), .ZN(G54) );
XOR2_X1 U893 ( .A(n1240), .B(n1241), .Z(n1239) );
XNOR2_X1 U894 ( .A(n1242), .B(n1243), .ZN(n1241) );
NAND3_X1 U895 ( .A1(n1216), .A2(G469), .A3(KEYINPUT41), .ZN(n1242) );
XNOR2_X1 U896 ( .A(n1244), .B(KEYINPUT8), .ZN(n1240) );
NAND2_X1 U897 ( .A1(KEYINPUT40), .A2(n1245), .ZN(n1244) );
XNOR2_X1 U898 ( .A(n1246), .B(n1247), .ZN(n1245) );
NOR2_X1 U899 ( .A1(n1206), .A2(n1248), .ZN(G51) );
XNOR2_X1 U900 ( .A(n1249), .B(n1250), .ZN(n1248) );
XOR2_X1 U901 ( .A(n1251), .B(n1252), .Z(n1250) );
NOR2_X1 U902 ( .A1(n1161), .A2(n1211), .ZN(n1252) );
INV_X1 U903 ( .A(n1216), .ZN(n1211) );
NOR2_X1 U904 ( .A1(n1253), .A2(n1218), .ZN(n1216) );
NOR4_X1 U905 ( .A1(n1194), .A2(n1174), .A3(n1193), .A4(n1175), .ZN(n1218) );
INV_X1 U906 ( .A(n1254), .ZN(n1175) );
OR4_X1 U907 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1193) );
INV_X1 U908 ( .A(n1259), .ZN(n1258) );
AND4_X1 U909 ( .A1(n1260), .A2(n1261), .A3(n1122), .A4(n1262), .ZN(n1255) );
XNOR2_X1 U910 ( .A(KEYINPUT9), .B(n1263), .ZN(n1262) );
XNOR2_X1 U911 ( .A(n1264), .B(KEYINPUT6), .ZN(n1260) );
NAND4_X1 U912 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1174) );
NAND3_X1 U913 ( .A1(n1269), .A2(n1270), .A3(n1131), .ZN(n1268) );
NAND2_X1 U914 ( .A1(n1271), .A2(n1272), .ZN(n1269) );
OR3_X1 U915 ( .A1(n1118), .A2(KEYINPUT29), .A3(n1273), .ZN(n1272) );
NAND2_X1 U916 ( .A1(n1264), .A2(n1274), .ZN(n1271) );
NAND2_X1 U917 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NAND3_X1 U918 ( .A1(n1150), .A2(n1277), .A3(n1278), .ZN(n1276) );
NAND3_X1 U919 ( .A1(n1279), .A2(n1280), .A3(n1137), .ZN(n1275) );
AND2_X1 U920 ( .A1(n1281), .A2(n1282), .ZN(n1267) );
NAND2_X1 U921 ( .A1(n1283), .A2(n1284), .ZN(n1266) );
NAND2_X1 U922 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND2_X1 U923 ( .A1(KEYINPUT29), .A2(n1261), .ZN(n1286) );
INV_X1 U924 ( .A(n1273), .ZN(n1261) );
NAND2_X1 U925 ( .A1(n1137), .A2(n1226), .ZN(n1285) );
OR2_X1 U926 ( .A1(n1287), .A2(n1139), .ZN(n1265) );
NAND4_X1 U927 ( .A1(n1288), .A2(n1289), .A3(n1290), .A4(n1291), .ZN(n1194) );
NAND4_X1 U928 ( .A1(n1131), .A2(n1292), .A3(n1263), .A4(n1139), .ZN(n1290) );
NAND2_X1 U929 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
NAND3_X1 U930 ( .A1(n1125), .A2(n1136), .A3(KEYINPUT47), .ZN(n1294) );
NAND2_X1 U931 ( .A1(n1105), .A2(n1295), .ZN(n1293) );
NAND2_X1 U932 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
NAND2_X1 U933 ( .A1(KEYINPUT17), .A2(n1278), .ZN(n1297) );
OR2_X1 U934 ( .A1(n1124), .A2(KEYINPUT31), .ZN(n1296) );
NAND3_X1 U935 ( .A1(n1105), .A2(n1298), .A3(n1225), .ZN(n1289) );
NAND2_X1 U936 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
OR2_X1 U937 ( .A1(n1104), .A2(KEYINPUT17), .ZN(n1300) );
NAND2_X1 U938 ( .A1(KEYINPUT31), .A2(n1226), .ZN(n1299) );
OR2_X1 U939 ( .A1(n1301), .A2(KEYINPUT47), .ZN(n1288) );
NAND2_X1 U940 ( .A1(n1302), .A2(KEYINPUT56), .ZN(n1251) );
XNOR2_X1 U941 ( .A(n1303), .B(KEYINPUT0), .ZN(n1302) );
NOR2_X1 U942 ( .A1(n1167), .A2(G952), .ZN(n1206) );
NAND2_X1 U943 ( .A1(n1304), .A2(n1305), .ZN(G48) );
NAND2_X1 U944 ( .A1(G146), .A2(n1306), .ZN(n1305) );
XOR2_X1 U945 ( .A(KEYINPUT24), .B(n1307), .Z(n1304) );
NOR2_X1 U946 ( .A1(G146), .A2(n1306), .ZN(n1307) );
NAND2_X1 U947 ( .A1(n1308), .A2(n1264), .ZN(n1306) );
XOR2_X1 U948 ( .A(n1287), .B(KEYINPUT22), .Z(n1308) );
NAND2_X1 U949 ( .A1(n1309), .A2(n1226), .ZN(n1287) );
XNOR2_X1 U950 ( .A(G143), .B(n1310), .ZN(G45) );
NAND4_X1 U951 ( .A1(n1279), .A2(n1137), .A3(n1311), .A4(n1312), .ZN(n1310) );
NOR3_X1 U952 ( .A1(n1139), .A2(n1313), .A3(n1314), .ZN(n1312) );
XNOR2_X1 U953 ( .A(n1131), .B(KEYINPUT10), .ZN(n1311) );
XNOR2_X1 U954 ( .A(G140), .B(n1282), .ZN(G42) );
NAND3_X1 U955 ( .A1(n1136), .A2(n1226), .A3(n1283), .ZN(n1282) );
INV_X1 U956 ( .A(n1315), .ZN(n1283) );
XNOR2_X1 U957 ( .A(n1316), .B(n1317), .ZN(G39) );
NOR2_X1 U958 ( .A1(n1315), .A2(n1273), .ZN(n1317) );
NAND3_X1 U959 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(G36) );
NAND2_X1 U960 ( .A1(G134), .A2(n1281), .ZN(n1320) );
INV_X1 U961 ( .A(n1321), .ZN(n1281) );
NAND2_X1 U962 ( .A1(n1322), .A2(n1323), .ZN(n1319) );
INV_X1 U963 ( .A(KEYINPUT39), .ZN(n1323) );
NAND2_X1 U964 ( .A1(n1321), .A2(n1324), .ZN(n1322) );
XNOR2_X1 U965 ( .A(KEYINPUT4), .B(n1183), .ZN(n1324) );
NAND2_X1 U966 ( .A1(KEYINPUT39), .A2(n1325), .ZN(n1318) );
NAND2_X1 U967 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
NAND3_X1 U968 ( .A1(KEYINPUT4), .A2(n1321), .A3(n1183), .ZN(n1327) );
NOR3_X1 U969 ( .A1(n1328), .A2(n1104), .A3(n1315), .ZN(n1321) );
OR2_X1 U970 ( .A1(n1183), .A2(KEYINPUT4), .ZN(n1326) );
XOR2_X1 U971 ( .A(G131), .B(n1329), .Z(G33) );
NOR4_X1 U972 ( .A1(KEYINPUT44), .A2(n1124), .A3(n1328), .A4(n1315), .ZN(n1329) );
NAND3_X1 U973 ( .A1(n1118), .A2(n1270), .A3(n1131), .ZN(n1315) );
NAND2_X1 U974 ( .A1(n1330), .A2(n1331), .ZN(n1118) );
OR2_X1 U975 ( .A1(n1139), .A2(KEYINPUT60), .ZN(n1331) );
NAND3_X1 U976 ( .A1(n1142), .A2(n1332), .A3(KEYINPUT60), .ZN(n1330) );
XNOR2_X1 U977 ( .A(G128), .B(n1333), .ZN(G30) );
NAND4_X1 U978 ( .A1(KEYINPUT52), .A2(n1309), .A3(n1278), .A4(n1264), .ZN(n1333) );
INV_X1 U979 ( .A(n1104), .ZN(n1278) );
AND4_X1 U980 ( .A1(n1131), .A2(n1150), .A3(n1277), .A4(n1270), .ZN(n1309) );
XNOR2_X1 U981 ( .A(G101), .B(n1291), .ZN(G3) );
NAND3_X1 U982 ( .A1(n1137), .A2(n1225), .A3(n1125), .ZN(n1291) );
INV_X1 U983 ( .A(n1328), .ZN(n1137) );
XNOR2_X1 U984 ( .A(G125), .B(n1254), .ZN(G27) );
NAND4_X1 U985 ( .A1(n1136), .A2(n1226), .A3(n1334), .A4(n1122), .ZN(n1254) );
NOR2_X1 U986 ( .A1(n1313), .A2(n1139), .ZN(n1334) );
INV_X1 U987 ( .A(n1264), .ZN(n1139) );
INV_X1 U988 ( .A(n1270), .ZN(n1313) );
NAND2_X1 U989 ( .A1(n1143), .A2(n1335), .ZN(n1270) );
NAND4_X1 U990 ( .A1(G953), .A2(G902), .A3(n1336), .A4(n1337), .ZN(n1335) );
INV_X1 U991 ( .A(G900), .ZN(n1337) );
XNOR2_X1 U992 ( .A(n1338), .B(n1339), .ZN(G24) );
NOR2_X1 U993 ( .A1(KEYINPUT35), .A2(n1259), .ZN(n1339) );
NAND4_X1 U994 ( .A1(n1340), .A2(n1105), .A3(n1279), .A4(n1280), .ZN(n1259) );
NOR2_X1 U995 ( .A1(n1277), .A2(n1150), .ZN(n1105) );
INV_X1 U996 ( .A(n1341), .ZN(n1340) );
XOR2_X1 U997 ( .A(G119), .B(n1342), .Z(G21) );
NOR2_X1 U998 ( .A1(n1273), .A2(n1341), .ZN(n1342) );
NAND3_X1 U999 ( .A1(n1150), .A2(n1277), .A3(n1125), .ZN(n1273) );
XNOR2_X1 U1000 ( .A(n1343), .B(n1256), .ZN(G18) );
NOR3_X1 U1001 ( .A1(n1328), .A2(n1104), .A3(n1341), .ZN(n1256) );
NAND2_X1 U1002 ( .A1(n1279), .A2(n1314), .ZN(n1104) );
XOR2_X1 U1003 ( .A(G113), .B(n1257), .Z(G15) );
NOR3_X1 U1004 ( .A1(n1328), .A2(n1124), .A3(n1341), .ZN(n1257) );
NAND3_X1 U1005 ( .A1(n1264), .A2(n1263), .A3(n1122), .ZN(n1341) );
NOR2_X1 U1006 ( .A1(n1344), .A2(n1129), .ZN(n1122) );
INV_X1 U1007 ( .A(n1226), .ZN(n1124) );
NOR2_X1 U1008 ( .A1(n1314), .A2(n1279), .ZN(n1226) );
NAND2_X1 U1009 ( .A1(n1345), .A2(n1277), .ZN(n1328) );
XOR2_X1 U1010 ( .A(n1301), .B(n1346), .Z(G12) );
XOR2_X1 U1011 ( .A(KEYINPUT12), .B(G110), .Z(n1346) );
NAND3_X1 U1012 ( .A1(n1136), .A2(n1225), .A3(n1125), .ZN(n1301) );
NOR2_X1 U1013 ( .A1(n1280), .A2(n1279), .ZN(n1125) );
XNOR2_X1 U1014 ( .A(n1154), .B(n1347), .ZN(n1279) );
NOR2_X1 U1015 ( .A1(G478), .A2(KEYINPUT3), .ZN(n1347) );
NOR2_X1 U1016 ( .A1(n1215), .A2(G902), .ZN(n1154) );
XNOR2_X1 U1017 ( .A(n1348), .B(n1349), .ZN(n1215) );
XOR2_X1 U1018 ( .A(n1350), .B(n1351), .Z(n1349) );
XNOR2_X1 U1019 ( .A(G116), .B(n1352), .ZN(n1351) );
NOR2_X1 U1020 ( .A1(G107), .A2(KEYINPUT34), .ZN(n1352) );
NAND2_X1 U1021 ( .A1(G217), .A2(n1353), .ZN(n1350) );
XOR2_X1 U1022 ( .A(n1354), .B(n1355), .Z(n1348) );
XNOR2_X1 U1023 ( .A(n1356), .B(G134), .ZN(n1355) );
XNOR2_X1 U1024 ( .A(G122), .B(G128), .ZN(n1354) );
INV_X1 U1025 ( .A(n1314), .ZN(n1280) );
XOR2_X1 U1026 ( .A(n1158), .B(n1160), .Z(n1314) );
INV_X1 U1027 ( .A(G475), .ZN(n1160) );
NOR2_X1 U1028 ( .A1(n1222), .A2(G902), .ZN(n1158) );
XOR2_X1 U1029 ( .A(n1357), .B(n1358), .Z(n1222) );
XOR2_X1 U1030 ( .A(G113), .B(n1359), .Z(n1358) );
XNOR2_X1 U1031 ( .A(G131), .B(n1338), .ZN(n1359) );
XOR2_X1 U1032 ( .A(n1360), .B(n1361), .Z(n1357) );
XNOR2_X1 U1033 ( .A(n1362), .B(n1363), .ZN(n1361) );
NOR2_X1 U1034 ( .A1(KEYINPUT37), .A2(n1364), .ZN(n1363) );
XNOR2_X1 U1035 ( .A(n1356), .B(n1365), .ZN(n1364) );
AND3_X1 U1036 ( .A1(G214), .A2(n1167), .A3(n1366), .ZN(n1365) );
NAND2_X1 U1037 ( .A1(n1367), .A2(KEYINPUT61), .ZN(n1360) );
XNOR2_X1 U1038 ( .A(n1368), .B(n1369), .ZN(n1367) );
NAND3_X1 U1039 ( .A1(n1370), .A2(n1371), .A3(KEYINPUT50), .ZN(n1368) );
OR2_X1 U1040 ( .A1(n1179), .A2(KEYINPUT63), .ZN(n1371) );
NAND3_X1 U1041 ( .A1(G125), .A2(n1372), .A3(KEYINPUT63), .ZN(n1370) );
INV_X1 U1042 ( .A(n1102), .ZN(n1225) );
NAND3_X1 U1043 ( .A1(n1264), .A2(n1263), .A3(n1131), .ZN(n1102) );
NOR2_X1 U1044 ( .A1(n1130), .A2(n1129), .ZN(n1131) );
AND2_X1 U1045 ( .A1(G221), .A2(n1373), .ZN(n1129) );
INV_X1 U1046 ( .A(n1344), .ZN(n1130) );
NAND3_X1 U1047 ( .A1(n1374), .A2(n1375), .A3(n1376), .ZN(n1344) );
NAND2_X1 U1048 ( .A1(G469), .A2(n1377), .ZN(n1376) );
NAND2_X1 U1049 ( .A1(n1378), .A2(n1379), .ZN(n1375) );
INV_X1 U1050 ( .A(KEYINPUT23), .ZN(n1379) );
NAND2_X1 U1051 ( .A1(n1380), .A2(n1381), .ZN(n1378) );
INV_X1 U1052 ( .A(G469), .ZN(n1381) );
XNOR2_X1 U1053 ( .A(KEYINPUT57), .B(n1377), .ZN(n1380) );
NAND2_X1 U1054 ( .A1(KEYINPUT23), .A2(n1382), .ZN(n1374) );
NAND2_X1 U1055 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
OR3_X1 U1056 ( .A1(n1377), .A2(G469), .A3(KEYINPUT57), .ZN(n1384) );
NAND2_X1 U1057 ( .A1(KEYINPUT57), .A2(n1377), .ZN(n1383) );
XOR2_X1 U1058 ( .A(n1153), .B(KEYINPUT62), .Z(n1377) );
NAND3_X1 U1059 ( .A1(n1385), .A2(n1386), .A3(n1387), .ZN(n1153) );
XNOR2_X1 U1060 ( .A(KEYINPUT36), .B(n1253), .ZN(n1387) );
NAND2_X1 U1061 ( .A1(n1388), .A2(n1389), .ZN(n1386) );
NAND2_X1 U1062 ( .A1(KEYINPUT27), .A2(n1247), .ZN(n1389) );
XNOR2_X1 U1063 ( .A(n1390), .B(n1391), .ZN(n1388) );
NOR2_X1 U1064 ( .A1(n1246), .A2(n1392), .ZN(n1390) );
NAND3_X1 U1065 ( .A1(n1247), .A2(n1393), .A3(KEYINPUT27), .ZN(n1385) );
XNOR2_X1 U1066 ( .A(n1394), .B(n1391), .ZN(n1393) );
INV_X1 U1067 ( .A(n1243), .ZN(n1391) );
XNOR2_X1 U1068 ( .A(n1395), .B(n1396), .ZN(n1243) );
XNOR2_X1 U1069 ( .A(n1372), .B(G110), .ZN(n1396) );
NAND2_X1 U1070 ( .A1(G227), .A2(n1167), .ZN(n1395) );
NOR2_X1 U1071 ( .A1(n1397), .A2(n1392), .ZN(n1394) );
INV_X1 U1072 ( .A(KEYINPUT28), .ZN(n1392) );
INV_X1 U1073 ( .A(n1246), .ZN(n1397) );
XOR2_X1 U1074 ( .A(n1398), .B(n1177), .Z(n1247) );
XNOR2_X1 U1075 ( .A(n1399), .B(G128), .ZN(n1177) );
NAND2_X1 U1076 ( .A1(n1400), .A2(KEYINPUT13), .ZN(n1399) );
XNOR2_X1 U1077 ( .A(n1401), .B(n1356), .ZN(n1400) );
INV_X1 U1078 ( .A(G143), .ZN(n1356) );
NAND2_X1 U1079 ( .A1(KEYINPUT18), .A2(n1369), .ZN(n1401) );
NAND2_X1 U1080 ( .A1(n1402), .A2(n1403), .ZN(n1398) );
NAND2_X1 U1081 ( .A1(n1404), .A2(n1405), .ZN(n1403) );
XOR2_X1 U1082 ( .A(KEYINPUT11), .B(n1406), .Z(n1402) );
NOR2_X1 U1083 ( .A1(n1405), .A2(n1404), .ZN(n1406) );
XNOR2_X1 U1084 ( .A(G107), .B(n1362), .ZN(n1404) );
NAND2_X1 U1085 ( .A1(n1143), .A2(n1407), .ZN(n1263) );
NAND4_X1 U1086 ( .A1(G953), .A2(G902), .A3(n1336), .A4(n1198), .ZN(n1407) );
INV_X1 U1087 ( .A(G898), .ZN(n1198) );
NAND3_X1 U1088 ( .A1(n1113), .A2(n1336), .A3(G952), .ZN(n1143) );
NAND2_X1 U1089 ( .A1(G237), .A2(G234), .ZN(n1336) );
XNOR2_X1 U1090 ( .A(G953), .B(KEYINPUT33), .ZN(n1113) );
NOR2_X1 U1091 ( .A1(n1142), .A2(n1141), .ZN(n1264) );
INV_X1 U1092 ( .A(n1332), .ZN(n1141) );
NAND2_X1 U1093 ( .A1(G214), .A2(n1408), .ZN(n1332) );
XNOR2_X1 U1094 ( .A(n1163), .B(n1161), .ZN(n1142) );
NAND2_X1 U1095 ( .A1(G210), .A2(n1408), .ZN(n1161) );
NAND2_X1 U1096 ( .A1(n1366), .A2(n1253), .ZN(n1408) );
NAND2_X1 U1097 ( .A1(n1409), .A2(n1253), .ZN(n1163) );
XNOR2_X1 U1098 ( .A(n1410), .B(n1303), .ZN(n1409) );
XOR2_X1 U1099 ( .A(G125), .B(n1411), .Z(n1303) );
INV_X1 U1100 ( .A(n1249), .ZN(n1410) );
XNOR2_X1 U1101 ( .A(n1412), .B(n1413), .ZN(n1249) );
XNOR2_X1 U1102 ( .A(n1204), .B(n1414), .ZN(n1413) );
NAND2_X1 U1103 ( .A1(G224), .A2(n1167), .ZN(n1414) );
INV_X1 U1104 ( .A(n1203), .ZN(n1204) );
NAND2_X1 U1105 ( .A1(n1415), .A2(n1416), .ZN(n1203) );
OR2_X1 U1106 ( .A1(n1338), .A2(G110), .ZN(n1416) );
XOR2_X1 U1107 ( .A(n1417), .B(KEYINPUT14), .Z(n1415) );
NAND2_X1 U1108 ( .A1(G110), .A2(n1338), .ZN(n1417) );
INV_X1 U1109 ( .A(G122), .ZN(n1338) );
NAND2_X1 U1110 ( .A1(n1202), .A2(n1205), .ZN(n1412) );
NAND2_X1 U1111 ( .A1(n1418), .A2(n1419), .ZN(n1205) );
XNOR2_X1 U1112 ( .A(n1420), .B(n1405), .ZN(n1419) );
NAND2_X1 U1113 ( .A1(n1421), .A2(n1422), .ZN(n1202) );
XNOR2_X1 U1114 ( .A(n1420), .B(n1423), .ZN(n1421) );
INV_X1 U1115 ( .A(n1405), .ZN(n1423) );
XOR2_X1 U1116 ( .A(G101), .B(KEYINPUT20), .Z(n1405) );
XOR2_X1 U1117 ( .A(n1424), .B(G107), .Z(n1420) );
NAND2_X1 U1118 ( .A1(KEYINPUT19), .A2(n1362), .ZN(n1424) );
INV_X1 U1119 ( .A(G104), .ZN(n1362) );
NOR2_X1 U1120 ( .A1(n1277), .A2(n1345), .ZN(n1136) );
INV_X1 U1121 ( .A(n1150), .ZN(n1345) );
XOR2_X1 U1122 ( .A(n1425), .B(n1210), .Z(n1150) );
NAND2_X1 U1123 ( .A1(G217), .A2(n1373), .ZN(n1210) );
NAND2_X1 U1124 ( .A1(G234), .A2(n1253), .ZN(n1373) );
NAND2_X1 U1125 ( .A1(n1208), .A2(n1253), .ZN(n1425) );
XNOR2_X1 U1126 ( .A(n1426), .B(n1427), .ZN(n1208) );
XOR2_X1 U1127 ( .A(n1428), .B(n1429), .Z(n1427) );
XOR2_X1 U1128 ( .A(G119), .B(G110), .Z(n1429) );
XNOR2_X1 U1129 ( .A(n1369), .B(G137), .ZN(n1428) );
INV_X1 U1130 ( .A(G146), .ZN(n1369) );
XNOR2_X1 U1131 ( .A(n1179), .B(n1430), .ZN(n1426) );
XNOR2_X1 U1132 ( .A(n1431), .B(n1432), .ZN(n1430) );
NOR2_X1 U1133 ( .A1(KEYINPUT2), .A2(n1433), .ZN(n1432) );
NAND3_X1 U1134 ( .A1(n1353), .A2(G221), .A3(KEYINPUT45), .ZN(n1431) );
AND2_X1 U1135 ( .A1(G234), .A2(n1167), .ZN(n1353) );
XNOR2_X1 U1136 ( .A(G125), .B(n1372), .ZN(n1179) );
INV_X1 U1137 ( .A(G140), .ZN(n1372) );
XNOR2_X1 U1138 ( .A(n1156), .B(n1434), .ZN(n1277) );
XNOR2_X1 U1139 ( .A(KEYINPUT46), .B(n1157), .ZN(n1434) );
INV_X1 U1140 ( .A(G472), .ZN(n1157) );
NAND2_X1 U1141 ( .A1(n1435), .A2(n1253), .ZN(n1156) );
INV_X1 U1142 ( .A(G902), .ZN(n1253) );
XNOR2_X1 U1143 ( .A(n1237), .B(n1436), .ZN(n1435) );
XNOR2_X1 U1144 ( .A(G101), .B(n1234), .ZN(n1436) );
NAND3_X1 U1145 ( .A1(n1366), .A2(n1167), .A3(G210), .ZN(n1234) );
INV_X1 U1146 ( .A(G953), .ZN(n1167) );
INV_X1 U1147 ( .A(G237), .ZN(n1366) );
XNOR2_X1 U1148 ( .A(n1411), .B(n1437), .ZN(n1237) );
XNOR2_X1 U1149 ( .A(n1246), .B(n1418), .ZN(n1437) );
INV_X1 U1150 ( .A(n1422), .ZN(n1418) );
XOR2_X1 U1151 ( .A(G113), .B(n1438), .Z(n1422) );
XNOR2_X1 U1152 ( .A(G119), .B(n1343), .ZN(n1438) );
INV_X1 U1153 ( .A(G116), .ZN(n1343) );
XOR2_X1 U1154 ( .A(n1439), .B(n1440), .Z(n1246) );
INV_X1 U1155 ( .A(n1181), .ZN(n1440) );
XOR2_X1 U1156 ( .A(G131), .B(KEYINPUT7), .Z(n1181) );
NAND2_X1 U1157 ( .A1(n1441), .A2(n1442), .ZN(n1439) );
NAND2_X1 U1158 ( .A1(n1443), .A2(n1183), .ZN(n1442) );
INV_X1 U1159 ( .A(G134), .ZN(n1183) );
NAND2_X1 U1160 ( .A1(n1444), .A2(n1445), .ZN(n1443) );
NAND2_X1 U1161 ( .A1(KEYINPUT21), .A2(n1316), .ZN(n1445) );
INV_X1 U1162 ( .A(G137), .ZN(n1316) );
NAND2_X1 U1163 ( .A1(G137), .A2(n1446), .ZN(n1441) );
NAND2_X1 U1164 ( .A1(KEYINPUT21), .A2(n1447), .ZN(n1446) );
NAND2_X1 U1165 ( .A1(G134), .A2(n1444), .ZN(n1447) );
INV_X1 U1166 ( .A(KEYINPUT58), .ZN(n1444) );
XNOR2_X1 U1167 ( .A(n1448), .B(n1449), .ZN(n1411) );
XNOR2_X1 U1168 ( .A(n1433), .B(n1450), .ZN(n1449) );
NOR2_X1 U1169 ( .A1(G146), .A2(KEYINPUT54), .ZN(n1450) );
INV_X1 U1170 ( .A(G128), .ZN(n1433) );
XNOR2_X1 U1171 ( .A(G143), .B(KEYINPUT32), .ZN(n1448) );
endmodule


