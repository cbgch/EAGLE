//Key = 0111000000011111111101110110010100001111011100000100101001111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305;

XOR2_X1 U724 ( .A(n995), .B(n996), .Z(G9) );
NAND2_X1 U725 ( .A1(n997), .A2(n998), .ZN(n996) );
NOR2_X1 U726 ( .A1(n999), .A2(n1000), .ZN(G75) );
NOR4_X1 U727 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n1000) );
NOR3_X1 U728 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n1003) );
NOR2_X1 U729 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
NOR2_X1 U730 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NOR2_X1 U731 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NOR2_X1 U732 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NOR2_X1 U733 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR2_X1 U734 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NOR2_X1 U735 ( .A1(n1020), .A2(n1021), .ZN(n1012) );
NOR2_X1 U736 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U737 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR3_X1 U738 ( .A1(n1015), .A2(n1026), .A3(n1021), .ZN(n1008) );
INV_X1 U739 ( .A(n1027), .ZN(n1021) );
NOR2_X1 U740 ( .A1(n997), .A2(n1028), .ZN(n1026) );
NAND3_X1 U741 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1001) );
NAND4_X1 U742 ( .A1(n1027), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1031) );
NOR2_X1 U743 ( .A1(n1015), .A2(n1005), .ZN(n1034) );
NAND2_X1 U744 ( .A1(n1035), .A2(n1036), .ZN(n1032) );
XOR2_X1 U745 ( .A(n1037), .B(KEYINPUT24), .Z(n1035) );
AND3_X1 U746 ( .A1(n1029), .A2(n1030), .A3(n1038), .ZN(n999) );
NAND4_X1 U747 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1029) );
NOR4_X1 U748 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
XOR2_X1 U749 ( .A(KEYINPUT40), .B(n1047), .Z(n1046) );
XNOR2_X1 U750 ( .A(G469), .B(n1048), .ZN(n1045) );
XOR2_X1 U751 ( .A(n1049), .B(n1050), .Z(n1044) );
XOR2_X1 U752 ( .A(n1051), .B(KEYINPUT32), .Z(n1050) );
NOR2_X1 U753 ( .A1(n1052), .A2(n1053), .ZN(n1041) );
XNOR2_X1 U754 ( .A(n1054), .B(n1055), .ZN(n1040) );
NAND2_X1 U755 ( .A1(KEYINPUT22), .A2(n1056), .ZN(n1055) );
XOR2_X1 U756 ( .A(KEYINPUT13), .B(n1057), .Z(n1039) );
XOR2_X1 U757 ( .A(n1058), .B(n1059), .Z(G72) );
XOR2_X1 U758 ( .A(n1060), .B(n1061), .Z(n1059) );
NAND2_X1 U759 ( .A1(n1030), .A2(n1004), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NAND2_X1 U761 ( .A1(G953), .A2(n1064), .ZN(n1063) );
XOR2_X1 U762 ( .A(n1065), .B(n1066), .Z(n1062) );
NAND2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NAND2_X1 U764 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XOR2_X1 U765 ( .A(n1071), .B(KEYINPUT49), .Z(n1069) );
NAND2_X1 U766 ( .A1(n1072), .A2(n1073), .ZN(n1067) );
XOR2_X1 U767 ( .A(KEYINPUT57), .B(n1074), .Z(n1072) );
INV_X1 U768 ( .A(n1071), .ZN(n1074) );
NOR2_X1 U769 ( .A1(n1075), .A2(n1030), .ZN(n1058) );
NOR2_X1 U770 ( .A1(n1076), .A2(n1064), .ZN(n1075) );
XOR2_X1 U771 ( .A(n1077), .B(n1078), .Z(G69) );
XOR2_X1 U772 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND2_X1 U773 ( .A1(G953), .A2(n1081), .ZN(n1080) );
NAND2_X1 U774 ( .A1(G898), .A2(G224), .ZN(n1081) );
NAND2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1079) );
NAND2_X1 U776 ( .A1(G953), .A2(n1084), .ZN(n1083) );
XOR2_X1 U777 ( .A(n1085), .B(n1086), .Z(n1082) );
NAND2_X1 U778 ( .A1(KEYINPUT3), .A2(n1087), .ZN(n1085) );
AND2_X1 U779 ( .A1(n1002), .A2(n1030), .ZN(n1077) );
NOR2_X1 U780 ( .A1(n1088), .A2(n1089), .ZN(G66) );
NOR3_X1 U781 ( .A1(n1054), .A2(n1090), .A3(n1091), .ZN(n1089) );
NOR3_X1 U782 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
INV_X1 U783 ( .A(n1095), .ZN(n1092) );
NOR2_X1 U784 ( .A1(n1096), .A2(n1095), .ZN(n1090) );
NOR2_X1 U785 ( .A1(n1097), .A2(n1093), .ZN(n1096) );
XOR2_X1 U786 ( .A(G217), .B(KEYINPUT39), .Z(n1093) );
NOR2_X1 U787 ( .A1(n1004), .A2(n1002), .ZN(n1097) );
NOR2_X1 U788 ( .A1(n1088), .A2(n1098), .ZN(G63) );
XOR2_X1 U789 ( .A(n1099), .B(n1100), .Z(n1098) );
NAND2_X1 U790 ( .A1(n1101), .A2(G478), .ZN(n1099) );
NOR3_X1 U791 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(G60) );
NOR3_X1 U792 ( .A1(n1105), .A2(n1030), .A3(n1038), .ZN(n1104) );
INV_X1 U793 ( .A(G952), .ZN(n1038) );
AND2_X1 U794 ( .A1(n1105), .A2(n1088), .ZN(n1103) );
INV_X1 U795 ( .A(KEYINPUT34), .ZN(n1105) );
XOR2_X1 U796 ( .A(n1106), .B(n1107), .Z(n1102) );
NAND2_X1 U797 ( .A1(n1101), .A2(G475), .ZN(n1106) );
XNOR2_X1 U798 ( .A(n1108), .B(n1109), .ZN(G6) );
NOR2_X1 U799 ( .A1(KEYINPUT10), .A2(n1110), .ZN(n1109) );
NOR2_X1 U800 ( .A1(n1088), .A2(n1111), .ZN(G57) );
XOR2_X1 U801 ( .A(n1112), .B(n1113), .Z(n1111) );
XNOR2_X1 U802 ( .A(n1114), .B(n1115), .ZN(n1113) );
NOR2_X1 U803 ( .A1(KEYINPUT45), .A2(n1116), .ZN(n1115) );
XOR2_X1 U804 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U805 ( .A(n1119), .B(KEYINPUT51), .Z(n1118) );
INV_X1 U806 ( .A(G101), .ZN(n1119) );
NAND2_X1 U807 ( .A1(n1120), .A2(KEYINPUT23), .ZN(n1114) );
XOR2_X1 U808 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U809 ( .A(KEYINPUT43), .B(G119), .Z(n1122) );
NAND2_X1 U810 ( .A1(n1101), .A2(G472), .ZN(n1112) );
NOR2_X1 U811 ( .A1(n1088), .A2(n1123), .ZN(G54) );
XOR2_X1 U812 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U813 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U814 ( .A1(n1101), .A2(G469), .ZN(n1126) );
INV_X1 U815 ( .A(n1094), .ZN(n1101) );
XOR2_X1 U816 ( .A(n1128), .B(n1129), .Z(n1124) );
XNOR2_X1 U817 ( .A(G140), .B(n1130), .ZN(n1129) );
NAND2_X1 U818 ( .A1(n1131), .A2(KEYINPUT29), .ZN(n1130) );
XOR2_X1 U819 ( .A(n1132), .B(n1073), .Z(n1131) );
INV_X1 U820 ( .A(n1070), .ZN(n1073) );
NAND2_X1 U821 ( .A1(n1133), .A2(KEYINPUT63), .ZN(n1128) );
XOR2_X1 U822 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U823 ( .A1(n1088), .A2(n1136), .ZN(G51) );
NOR2_X1 U824 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U825 ( .A(n1139), .B(KEYINPUT11), .Z(n1138) );
NAND2_X1 U826 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR2_X1 U827 ( .A1(n1140), .A2(n1141), .ZN(n1137) );
XNOR2_X1 U828 ( .A(n1142), .B(n1143), .ZN(n1141) );
NOR2_X1 U829 ( .A1(KEYINPUT53), .A2(n1144), .ZN(n1143) );
XOR2_X1 U830 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR2_X1 U831 ( .A1(n1094), .A2(n1049), .ZN(n1140) );
NAND2_X1 U832 ( .A1(G902), .A2(n1147), .ZN(n1094) );
OR2_X1 U833 ( .A1(n1002), .A2(n1004), .ZN(n1147) );
NAND4_X1 U834 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1004) );
AND3_X1 U835 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
OR2_X1 U836 ( .A1(n1155), .A2(KEYINPUT28), .ZN(n1150) );
NAND4_X1 U837 ( .A1(n1156), .A2(n1157), .A3(n997), .A4(n1027), .ZN(n1149) );
NAND2_X1 U838 ( .A1(n1017), .A2(n1158), .ZN(n1148) );
NAND3_X1 U839 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1158) );
XNOR2_X1 U840 ( .A(KEYINPUT36), .B(n1162), .ZN(n1161) );
NAND2_X1 U841 ( .A1(n1028), .A2(n1163), .ZN(n1160) );
NAND2_X1 U842 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND4_X1 U843 ( .A1(KEYINPUT28), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1165) );
NAND2_X1 U844 ( .A1(n1169), .A2(n1156), .ZN(n1164) );
XNOR2_X1 U845 ( .A(n1170), .B(KEYINPUT42), .ZN(n1169) );
XNOR2_X1 U846 ( .A(KEYINPUT38), .B(n1171), .ZN(n1159) );
NAND4_X1 U847 ( .A1(n1108), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1002) );
AND4_X1 U848 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1174) );
INV_X1 U849 ( .A(n1179), .ZN(n1175) );
NOR2_X1 U850 ( .A1(n1180), .A2(n1181), .ZN(n1173) );
NOR3_X1 U851 ( .A1(n1037), .A2(n1182), .A3(n1011), .ZN(n1181) );
NOR4_X1 U852 ( .A1(n1183), .A2(n1184), .A3(n1007), .A4(n1185), .ZN(n1180) );
NOR2_X1 U853 ( .A1(KEYINPUT54), .A2(n1186), .ZN(n1184) );
NOR3_X1 U854 ( .A1(n1187), .A2(n1188), .A3(n1017), .ZN(n1186) );
AND2_X1 U855 ( .A1(n1182), .A2(KEYINPUT54), .ZN(n1183) );
NAND2_X1 U856 ( .A1(n1028), .A2(n998), .ZN(n1108) );
NOR2_X1 U857 ( .A1(n1007), .A2(n1182), .ZN(n998) );
INV_X1 U858 ( .A(n1189), .ZN(n1007) );
NOR2_X1 U859 ( .A1(n1030), .A2(G952), .ZN(n1088) );
XNOR2_X1 U860 ( .A(G146), .B(n1190), .ZN(G48) );
NAND3_X1 U861 ( .A1(n1170), .A2(n1017), .A3(n1191), .ZN(n1190) );
XOR2_X1 U862 ( .A(G143), .B(n1192), .Z(G45) );
NOR2_X1 U863 ( .A1(n1193), .A2(n1162), .ZN(n1192) );
NAND4_X1 U864 ( .A1(n1156), .A2(n1157), .A3(n1043), .A4(n1047), .ZN(n1162) );
XNOR2_X1 U865 ( .A(G140), .B(n1152), .ZN(G42) );
NAND3_X1 U866 ( .A1(n1168), .A2(n1027), .A3(n1191), .ZN(n1152) );
XNOR2_X1 U867 ( .A(G137), .B(n1154), .ZN(G39) );
NAND4_X1 U868 ( .A1(n1156), .A2(n1170), .A3(n1033), .A4(n1027), .ZN(n1154) );
XNOR2_X1 U869 ( .A(G134), .B(n1194), .ZN(G36) );
NAND4_X1 U870 ( .A1(n1027), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1194) );
NOR2_X1 U871 ( .A1(n1185), .A2(n1037), .ZN(n1197) );
XOR2_X1 U872 ( .A(KEYINPUT20), .B(n1023), .Z(n1196) );
INV_X1 U873 ( .A(n1187), .ZN(n1023) );
XNOR2_X1 U874 ( .A(G131), .B(n1153), .ZN(G33) );
NAND3_X1 U875 ( .A1(n1157), .A2(n1027), .A3(n1191), .ZN(n1153) );
AND2_X1 U876 ( .A1(n1156), .A2(n1028), .ZN(n1191) );
NAND2_X1 U877 ( .A1(n1198), .A2(n1199), .ZN(n1027) );
OR3_X1 U878 ( .A1(n1018), .A2(n1053), .A3(KEYINPUT56), .ZN(n1199) );
INV_X1 U879 ( .A(n1019), .ZN(n1053) );
NAND2_X1 U880 ( .A1(KEYINPUT56), .A2(n1017), .ZN(n1198) );
INV_X1 U881 ( .A(n1193), .ZN(n1017) );
XOR2_X1 U882 ( .A(G128), .B(n1200), .Z(G30) );
NOR2_X1 U883 ( .A1(n1193), .A2(n1171), .ZN(n1200) );
NAND3_X1 U884 ( .A1(n1170), .A2(n997), .A3(n1156), .ZN(n1171) );
NOR2_X1 U885 ( .A1(n1187), .A2(n1166), .ZN(n1156) );
XOR2_X1 U886 ( .A(G101), .B(n1201), .Z(G3) );
NOR4_X1 U887 ( .A1(KEYINPUT35), .A2(n1182), .A3(n1011), .A4(n1037), .ZN(n1201) );
INV_X1 U888 ( .A(n1157), .ZN(n1037) );
XOR2_X1 U889 ( .A(n1155), .B(n1202), .Z(G27) );
NAND2_X1 U890 ( .A1(KEYINPUT61), .A2(G125), .ZN(n1202) );
NAND4_X1 U891 ( .A1(n1028), .A2(n1167), .A3(n1203), .A4(n1168), .ZN(n1155) );
INV_X1 U892 ( .A(n1036), .ZN(n1168) );
NOR2_X1 U893 ( .A1(n1166), .A2(n1193), .ZN(n1203) );
INV_X1 U894 ( .A(n1195), .ZN(n1166) );
NAND2_X1 U895 ( .A1(n1204), .A2(n1005), .ZN(n1195) );
NAND4_X1 U896 ( .A1(G902), .A2(n1205), .A3(n1206), .A4(n1064), .ZN(n1204) );
INV_X1 U897 ( .A(G900), .ZN(n1064) );
XOR2_X1 U898 ( .A(KEYINPUT46), .B(G953), .Z(n1205) );
XOR2_X1 U899 ( .A(n1207), .B(n1172), .Z(G24) );
NAND4_X1 U900 ( .A1(n1208), .A2(n1189), .A3(n1043), .A4(n1047), .ZN(n1172) );
NOR2_X1 U901 ( .A1(n1209), .A2(n1057), .ZN(n1189) );
XNOR2_X1 U902 ( .A(G119), .B(n1178), .ZN(G21) );
NAND3_X1 U903 ( .A1(n1208), .A2(n1033), .A3(n1170), .ZN(n1178) );
AND2_X1 U904 ( .A1(n1057), .A2(n1209), .ZN(n1170) );
INV_X1 U905 ( .A(n1210), .ZN(n1057) );
INV_X1 U906 ( .A(n1011), .ZN(n1033) );
XNOR2_X1 U907 ( .A(G116), .B(n1177), .ZN(G18) );
NAND3_X1 U908 ( .A1(n1208), .A2(n997), .A3(n1157), .ZN(n1177) );
INV_X1 U909 ( .A(n1185), .ZN(n997) );
NAND2_X1 U910 ( .A1(n1211), .A2(n1047), .ZN(n1185) );
INV_X1 U911 ( .A(n1212), .ZN(n1047) );
XOR2_X1 U912 ( .A(KEYINPUT5), .B(n1213), .Z(n1211) );
INV_X1 U913 ( .A(n1214), .ZN(n1213) );
XOR2_X1 U914 ( .A(n1176), .B(n1215), .Z(G15) );
NAND2_X1 U915 ( .A1(KEYINPUT25), .A2(G113), .ZN(n1215) );
NAND3_X1 U916 ( .A1(n1208), .A2(n1028), .A3(n1157), .ZN(n1176) );
NOR2_X1 U917 ( .A1(n1209), .A2(n1210), .ZN(n1157) );
AND2_X1 U918 ( .A1(n1212), .A2(n1043), .ZN(n1028) );
NOR3_X1 U919 ( .A1(n1193), .A2(n1188), .A3(n1015), .ZN(n1208) );
INV_X1 U920 ( .A(n1167), .ZN(n1015) );
NOR2_X1 U921 ( .A1(n1024), .A2(n1052), .ZN(n1167) );
INV_X1 U922 ( .A(n1025), .ZN(n1052) );
XOR2_X1 U923 ( .A(G110), .B(n1179), .Z(G12) );
NOR3_X1 U924 ( .A1(n1036), .A2(n1182), .A3(n1011), .ZN(n1179) );
NAND2_X1 U925 ( .A1(n1216), .A2(n1212), .ZN(n1011) );
XOR2_X1 U926 ( .A(n1217), .B(G478), .Z(n1212) );
NAND2_X1 U927 ( .A1(n1100), .A2(n1218), .ZN(n1217) );
XOR2_X1 U928 ( .A(n1219), .B(n1220), .Z(n1100) );
XOR2_X1 U929 ( .A(n1221), .B(n1222), .Z(n1220) );
XOR2_X1 U930 ( .A(n1223), .B(G116), .Z(n1222) );
NAND2_X1 U931 ( .A1(KEYINPUT15), .A2(n1224), .ZN(n1223) );
NAND3_X1 U932 ( .A1(G217), .A2(n1030), .A3(G234), .ZN(n1224) );
NAND2_X1 U933 ( .A1(KEYINPUT12), .A2(n1207), .ZN(n1221) );
XOR2_X1 U934 ( .A(n1225), .B(n1226), .Z(n1219) );
NOR2_X1 U935 ( .A1(G107), .A2(KEYINPUT0), .ZN(n1226) );
NAND2_X1 U936 ( .A1(n1227), .A2(n1228), .ZN(n1225) );
OR2_X1 U937 ( .A1(n1135), .A2(n1070), .ZN(n1228) );
XOR2_X1 U938 ( .A(n1229), .B(KEYINPUT7), .Z(n1227) );
NAND2_X1 U939 ( .A1(n1070), .A2(n1135), .ZN(n1229) );
XOR2_X1 U940 ( .A(n1214), .B(KEYINPUT37), .Z(n1216) );
XNOR2_X1 U941 ( .A(n1043), .B(KEYINPUT31), .ZN(n1214) );
XNOR2_X1 U942 ( .A(n1230), .B(G475), .ZN(n1043) );
NAND2_X1 U943 ( .A1(n1231), .A2(n1218), .ZN(n1230) );
XOR2_X1 U944 ( .A(KEYINPUT21), .B(n1232), .Z(n1231) );
INV_X1 U945 ( .A(n1107), .ZN(n1232) );
XOR2_X1 U946 ( .A(n1233), .B(n1234), .Z(n1107) );
XNOR2_X1 U947 ( .A(n1235), .B(n1236), .ZN(n1234) );
XOR2_X1 U948 ( .A(n1237), .B(n1238), .Z(n1236) );
NOR2_X1 U949 ( .A1(G125), .A2(KEYINPUT62), .ZN(n1238) );
NAND2_X1 U950 ( .A1(G214), .A2(n1239), .ZN(n1237) );
XOR2_X1 U951 ( .A(n1240), .B(n1241), .Z(n1233) );
XOR2_X1 U952 ( .A(G143), .B(G131), .Z(n1241) );
NAND2_X1 U953 ( .A1(KEYINPUT16), .A2(n1242), .ZN(n1240) );
XOR2_X1 U954 ( .A(n1110), .B(n1243), .Z(n1242) );
NAND2_X1 U955 ( .A1(KEYINPUT26), .A2(n1244), .ZN(n1243) );
XOR2_X1 U956 ( .A(G122), .B(G113), .Z(n1244) );
INV_X1 U957 ( .A(G104), .ZN(n1110) );
OR3_X1 U958 ( .A1(n1193), .A2(n1188), .A3(n1187), .ZN(n1182) );
NAND2_X1 U959 ( .A1(n1024), .A2(n1025), .ZN(n1187) );
NAND2_X1 U960 ( .A1(G221), .A2(n1245), .ZN(n1025) );
XOR2_X1 U961 ( .A(n1246), .B(G469), .Z(n1024) );
NAND2_X1 U962 ( .A1(KEYINPUT59), .A2(n1048), .ZN(n1246) );
NAND2_X1 U963 ( .A1(n1247), .A2(n1218), .ZN(n1048) );
XOR2_X1 U964 ( .A(n1248), .B(n1249), .Z(n1247) );
XOR2_X1 U965 ( .A(n1250), .B(n1251), .Z(n1249) );
XOR2_X1 U966 ( .A(KEYINPUT27), .B(n1252), .Z(n1251) );
NOR2_X1 U967 ( .A1(G140), .A2(KEYINPUT8), .ZN(n1252) );
XOR2_X1 U968 ( .A(n1127), .B(n1253), .Z(n1248) );
INV_X1 U969 ( .A(n1134), .ZN(n1253) );
XNOR2_X1 U970 ( .A(G146), .B(KEYINPUT52), .ZN(n1134) );
XOR2_X1 U971 ( .A(n1254), .B(n1255), .Z(n1127) );
XOR2_X1 U972 ( .A(G104), .B(n1256), .Z(n1255) );
XOR2_X1 U973 ( .A(KEYINPUT60), .B(G110), .Z(n1256) );
XOR2_X1 U974 ( .A(n1257), .B(n1258), .Z(n1254) );
XOR2_X1 U975 ( .A(G101), .B(n1259), .Z(n1258) );
NOR2_X1 U976 ( .A1(G953), .A2(n1076), .ZN(n1259) );
INV_X1 U977 ( .A(G227), .ZN(n1076) );
NAND2_X1 U978 ( .A1(KEYINPUT2), .A2(n995), .ZN(n1257) );
INV_X1 U979 ( .A(G107), .ZN(n995) );
AND2_X1 U980 ( .A1(n1005), .A2(n1260), .ZN(n1188) );
NAND4_X1 U981 ( .A1(G953), .A2(G902), .A3(n1206), .A4(n1084), .ZN(n1260) );
INV_X1 U982 ( .A(G898), .ZN(n1084) );
NAND3_X1 U983 ( .A1(n1206), .A2(n1030), .A3(G952), .ZN(n1005) );
NAND2_X1 U984 ( .A1(G237), .A2(n1261), .ZN(n1206) );
XOR2_X1 U985 ( .A(KEYINPUT47), .B(G234), .Z(n1261) );
NAND2_X1 U986 ( .A1(n1018), .A2(n1019), .ZN(n1193) );
NAND2_X1 U987 ( .A1(G214), .A2(n1262), .ZN(n1019) );
XNOR2_X1 U988 ( .A(n1263), .B(n1051), .ZN(n1018) );
NAND2_X1 U989 ( .A1(n1264), .A2(n1218), .ZN(n1051) );
XOR2_X1 U990 ( .A(n1265), .B(n1146), .Z(n1264) );
XOR2_X1 U991 ( .A(G125), .B(n1266), .Z(n1146) );
AND2_X1 U992 ( .A1(G224), .A2(n1030), .ZN(n1266) );
XNOR2_X1 U993 ( .A(n1267), .B(n1268), .ZN(n1265) );
NAND2_X1 U994 ( .A1(KEYINPUT58), .A2(n1142), .ZN(n1268) );
XNOR2_X1 U995 ( .A(n1269), .B(n1086), .ZN(n1142) );
XNOR2_X1 U996 ( .A(n1270), .B(n1271), .ZN(n1086) );
XOR2_X1 U997 ( .A(n1272), .B(n1273), .Z(n1271) );
NOR2_X1 U998 ( .A1(G116), .A2(KEYINPUT30), .ZN(n1272) );
XOR2_X1 U999 ( .A(n1274), .B(n1275), .Z(n1270) );
NOR2_X1 U1000 ( .A1(KEYINPUT4), .A2(n1276), .ZN(n1275) );
NAND2_X1 U1001 ( .A1(KEYINPUT14), .A2(n1277), .ZN(n1274) );
XOR2_X1 U1002 ( .A(G107), .B(G104), .Z(n1277) );
XNOR2_X1 U1003 ( .A(n1087), .B(KEYINPUT50), .ZN(n1269) );
AND2_X1 U1004 ( .A1(n1278), .A2(n1279), .ZN(n1087) );
NAND2_X1 U1005 ( .A1(n1280), .A2(G110), .ZN(n1279) );
XOR2_X1 U1006 ( .A(KEYINPUT33), .B(n1207), .Z(n1280) );
INV_X1 U1007 ( .A(G122), .ZN(n1207) );
XOR2_X1 U1008 ( .A(n1281), .B(KEYINPUT44), .Z(n1278) );
NAND2_X1 U1009 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
INV_X1 U1010 ( .A(G110), .ZN(n1283) );
XOR2_X1 U1011 ( .A(KEYINPUT33), .B(G122), .Z(n1282) );
NAND2_X1 U1012 ( .A1(KEYINPUT18), .A2(n1145), .ZN(n1267) );
XOR2_X1 U1013 ( .A(n1284), .B(n1135), .Z(n1145) );
NAND2_X1 U1014 ( .A1(KEYINPUT41), .A2(n1049), .ZN(n1263) );
NAND2_X1 U1015 ( .A1(G210), .A2(n1262), .ZN(n1049) );
NAND2_X1 U1016 ( .A1(n1285), .A2(n1218), .ZN(n1262) );
INV_X1 U1017 ( .A(G237), .ZN(n1285) );
NAND2_X1 U1018 ( .A1(n1210), .A2(n1209), .ZN(n1036) );
XNOR2_X1 U1019 ( .A(n1054), .B(n1056), .ZN(n1209) );
NAND2_X1 U1020 ( .A1(G217), .A2(n1245), .ZN(n1056) );
NAND2_X1 U1021 ( .A1(G234), .A2(n1218), .ZN(n1245) );
NOR2_X1 U1022 ( .A1(n1095), .A2(G902), .ZN(n1054) );
XOR2_X1 U1023 ( .A(n1286), .B(n1287), .Z(n1095) );
XOR2_X1 U1024 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U1025 ( .A(G137), .B(G110), .Z(n1289) );
NOR2_X1 U1026 ( .A1(KEYINPUT6), .A2(n1290), .ZN(n1288) );
NOR2_X1 U1027 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XOR2_X1 U1028 ( .A(n1293), .B(KEYINPUT17), .Z(n1292) );
NAND2_X1 U1029 ( .A1(G119), .A2(n1294), .ZN(n1293) );
NOR2_X1 U1030 ( .A1(G119), .A2(n1294), .ZN(n1291) );
XNOR2_X1 U1031 ( .A(n1066), .B(n1295), .ZN(n1286) );
AND3_X1 U1032 ( .A1(G221), .A2(n1030), .A3(G234), .ZN(n1295) );
INV_X1 U1033 ( .A(G953), .ZN(n1030) );
XOR2_X1 U1034 ( .A(G125), .B(n1235), .Z(n1066) );
XOR2_X1 U1035 ( .A(G140), .B(G146), .Z(n1235) );
XOR2_X1 U1036 ( .A(n1296), .B(G472), .Z(n1210) );
NAND2_X1 U1037 ( .A1(n1297), .A2(n1218), .ZN(n1296) );
INV_X1 U1038 ( .A(G902), .ZN(n1218) );
XOR2_X1 U1039 ( .A(n1298), .B(n1299), .Z(n1297) );
XNOR2_X1 U1040 ( .A(KEYINPUT55), .B(n1117), .ZN(n1299) );
NAND2_X1 U1041 ( .A1(G210), .A2(n1239), .ZN(n1117) );
NOR2_X1 U1042 ( .A1(G953), .A2(G237), .ZN(n1239) );
XOR2_X1 U1043 ( .A(n1121), .B(n1273), .Z(n1298) );
XOR2_X1 U1044 ( .A(G101), .B(G119), .Z(n1273) );
XOR2_X1 U1045 ( .A(n1300), .B(n1301), .Z(n1121) );
XOR2_X1 U1046 ( .A(n1284), .B(n1302), .Z(n1301) );
NAND2_X1 U1047 ( .A1(KEYINPUT1), .A2(n1276), .ZN(n1302) );
INV_X1 U1048 ( .A(G113), .ZN(n1276) );
NAND2_X1 U1049 ( .A1(n1303), .A2(G146), .ZN(n1284) );
INV_X1 U1050 ( .A(KEYINPUT9), .ZN(n1303) );
XNOR2_X1 U1051 ( .A(n1250), .B(n1304), .ZN(n1300) );
NOR2_X1 U1052 ( .A1(G116), .A2(KEYINPUT48), .ZN(n1304) );
XOR2_X1 U1053 ( .A(n1070), .B(n1071), .Z(n1250) );
XOR2_X1 U1054 ( .A(n1132), .B(n1135), .Z(n1071) );
XOR2_X1 U1055 ( .A(n1305), .B(n1294), .Z(n1135) );
INV_X1 U1056 ( .A(G128), .ZN(n1294) );
INV_X1 U1057 ( .A(G143), .ZN(n1305) );
XNOR2_X1 U1058 ( .A(G131), .B(G137), .ZN(n1132) );
XNOR2_X1 U1059 ( .A(G134), .B(KEYINPUT19), .ZN(n1070) );
endmodule


