//Key = 1010111010011011011100011000111111010011100110100110011111110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292;

XOR2_X1 U706 ( .A(G107), .B(n982), .Z(G9) );
NOR2_X1 U707 ( .A1(n983), .A2(n984), .ZN(G75) );
NOR4_X1 U708 ( .A1(n985), .A2(n986), .A3(G953), .A4(n987), .ZN(n984) );
NOR2_X1 U709 ( .A1(n988), .A2(n989), .ZN(n986) );
NOR2_X1 U710 ( .A1(n990), .A2(n991), .ZN(n988) );
NOR3_X1 U711 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
NOR4_X1 U712 ( .A1(n995), .A2(n996), .A3(n997), .A4(n998), .ZN(n993) );
NOR3_X1 U713 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n998) );
NOR3_X1 U714 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(n997) );
NOR3_X1 U715 ( .A1(n1002), .A2(n1005), .A3(n1000), .ZN(n990) );
NOR2_X1 U716 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
AND2_X1 U717 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NOR2_X1 U718 ( .A1(n1010), .A2(n994), .ZN(n1006) );
NAND3_X1 U719 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n985) );
XOR2_X1 U720 ( .A(KEYINPUT46), .B(n1014), .Z(n1012) );
NOR4_X1 U721 ( .A1(n1015), .A2(n992), .A3(n1016), .A4(n1017), .ZN(n1014) );
NAND3_X1 U722 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1015) );
XOR2_X1 U723 ( .A(n1000), .B(KEYINPUT57), .Z(n1020) );
INV_X1 U724 ( .A(n989), .ZN(n1018) );
NOR3_X1 U725 ( .A1(n987), .A2(G953), .A3(G952), .ZN(n983) );
AND4_X1 U726 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n987) );
NOR4_X1 U727 ( .A1(n1025), .A2(n1026), .A3(n994), .A4(n1027), .ZN(n1024) );
XOR2_X1 U728 ( .A(n1028), .B(n1029), .Z(n1027) );
NAND2_X1 U729 ( .A1(KEYINPUT14), .A2(G469), .ZN(n1029) );
INV_X1 U730 ( .A(n999), .ZN(n1026) );
XOR2_X1 U731 ( .A(n1030), .B(G475), .Z(n1023) );
XOR2_X1 U732 ( .A(n1031), .B(KEYINPUT63), .Z(n1022) );
XOR2_X1 U733 ( .A(n1032), .B(KEYINPUT22), .Z(n1021) );
XOR2_X1 U734 ( .A(n1033), .B(n1034), .Z(G72) );
NOR2_X1 U735 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U736 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NAND2_X1 U737 ( .A1(n1039), .A2(n1040), .ZN(n1033) );
NAND3_X1 U738 ( .A1(n1041), .A2(n1036), .A3(n1042), .ZN(n1040) );
XOR2_X1 U739 ( .A(KEYINPUT53), .B(n1043), .Z(n1039) );
NOR2_X1 U740 ( .A1(n1041), .A2(n1042), .ZN(n1043) );
NAND2_X1 U741 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NAND2_X1 U742 ( .A1(n1046), .A2(n1038), .ZN(n1045) );
XOR2_X1 U743 ( .A(n1047), .B(n1048), .Z(n1044) );
XOR2_X1 U744 ( .A(n1049), .B(n1050), .Z(G69) );
NOR2_X1 U745 ( .A1(n1051), .A2(n1036), .ZN(n1050) );
NOR2_X1 U746 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U747 ( .A1(n1054), .A2(n1055), .ZN(n1049) );
NAND2_X1 U748 ( .A1(KEYINPUT26), .A2(n1056), .ZN(n1055) );
XOR2_X1 U749 ( .A(n1057), .B(n1058), .Z(n1054) );
NOR2_X1 U750 ( .A1(n1013), .A2(G953), .ZN(n1058) );
OR2_X1 U751 ( .A1(n1056), .A2(KEYINPUT26), .ZN(n1057) );
NAND2_X1 U752 ( .A1(n1059), .A2(n1060), .ZN(n1056) );
NAND2_X1 U753 ( .A1(n1061), .A2(n1046), .ZN(n1060) );
XOR2_X1 U754 ( .A(KEYINPUT12), .B(G898), .Z(n1061) );
XOR2_X1 U755 ( .A(n1062), .B(n1063), .Z(n1059) );
NOR2_X1 U756 ( .A1(n1064), .A2(n1065), .ZN(G66) );
XOR2_X1 U757 ( .A(n1066), .B(n1067), .Z(n1065) );
NOR2_X1 U758 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U759 ( .A1(n1064), .A2(n1070), .ZN(G63) );
XOR2_X1 U760 ( .A(n1071), .B(n1072), .Z(n1070) );
NOR2_X1 U761 ( .A1(n1073), .A2(n1069), .ZN(n1072) );
INV_X1 U762 ( .A(G478), .ZN(n1073) );
NAND2_X1 U763 ( .A1(KEYINPUT19), .A2(n1074), .ZN(n1071) );
NOR3_X1 U764 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(G60) );
AND2_X1 U765 ( .A1(KEYINPUT62), .A2(n1064), .ZN(n1077) );
NOR3_X1 U766 ( .A1(KEYINPUT62), .A2(n1036), .A3(n1078), .ZN(n1076) );
XOR2_X1 U767 ( .A(n1079), .B(n1080), .Z(n1075) );
NOR2_X1 U768 ( .A1(n1081), .A2(n1069), .ZN(n1079) );
NAND2_X1 U769 ( .A1(n1082), .A2(n1083), .ZN(G6) );
NAND2_X1 U770 ( .A1(G104), .A2(n1084), .ZN(n1083) );
XOR2_X1 U771 ( .A(KEYINPUT50), .B(n1085), .Z(n1082) );
NOR2_X1 U772 ( .A1(G104), .A2(n1084), .ZN(n1085) );
NOR3_X1 U773 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(G57) );
NOR3_X1 U774 ( .A1(n1089), .A2(n1036), .A3(n1078), .ZN(n1088) );
INV_X1 U775 ( .A(G952), .ZN(n1078) );
AND2_X1 U776 ( .A1(n1089), .A2(n1064), .ZN(n1087) );
INV_X1 U777 ( .A(KEYINPUT47), .ZN(n1089) );
XOR2_X1 U778 ( .A(n1090), .B(n1091), .Z(n1086) );
XOR2_X1 U779 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND2_X1 U780 ( .A1(KEYINPUT32), .A2(n1094), .ZN(n1093) );
NAND2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1090) );
NAND2_X1 U782 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U783 ( .A(KEYINPUT44), .B(n1099), .Z(n1097) );
NOR2_X1 U784 ( .A1(n1100), .A2(n1069), .ZN(n1099) );
OR3_X1 U785 ( .A1(n1069), .A2(n1100), .A3(n1098), .ZN(n1095) );
XOR2_X1 U786 ( .A(n1101), .B(n1102), .Z(n1098) );
NAND2_X1 U787 ( .A1(KEYINPUT59), .A2(n1103), .ZN(n1101) );
INV_X1 U788 ( .A(G472), .ZN(n1100) );
NOR2_X1 U789 ( .A1(n1064), .A2(n1104), .ZN(G54) );
XOR2_X1 U790 ( .A(n1105), .B(n1106), .Z(n1104) );
XOR2_X1 U791 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND2_X1 U792 ( .A1(KEYINPUT15), .A2(n1109), .ZN(n1108) );
NAND3_X1 U793 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1107) );
NAND2_X1 U794 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
INV_X1 U795 ( .A(KEYINPUT55), .ZN(n1114) );
NAND2_X1 U796 ( .A1(n1115), .A2(G110), .ZN(n1113) );
XOR2_X1 U797 ( .A(KEYINPUT16), .B(n1116), .Z(n1115) );
NAND2_X1 U798 ( .A1(KEYINPUT55), .A2(n1117), .ZN(n1110) );
NAND2_X1 U799 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
OR3_X1 U800 ( .A1(n1120), .A2(G140), .A3(KEYINPUT16), .ZN(n1119) );
NAND2_X1 U801 ( .A1(KEYINPUT16), .A2(G140), .ZN(n1118) );
XOR2_X1 U802 ( .A(n1121), .B(n1122), .Z(n1105) );
NOR2_X1 U803 ( .A1(n1123), .A2(n1069), .ZN(n1122) );
INV_X1 U804 ( .A(G469), .ZN(n1123) );
NOR2_X1 U805 ( .A1(n1064), .A2(n1124), .ZN(G51) );
XNOR2_X1 U806 ( .A(n1125), .B(n1126), .ZN(n1124) );
XOR2_X1 U807 ( .A(KEYINPUT45), .B(n1127), .Z(n1126) );
NOR2_X1 U808 ( .A1(n1128), .A2(n1069), .ZN(n1127) );
NAND2_X1 U809 ( .A1(G902), .A2(n1129), .ZN(n1069) );
NAND2_X1 U810 ( .A1(n1013), .A2(n1011), .ZN(n1129) );
INV_X1 U811 ( .A(n1041), .ZN(n1011) );
NAND4_X1 U812 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1041) );
NOR4_X1 U813 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1133) );
OR3_X1 U814 ( .A1(n1002), .A2(n1010), .A3(n1138), .ZN(n1132) );
NOR2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(n1010) );
NAND4_X1 U816 ( .A1(n1141), .A2(n1140), .A3(n1142), .A4(n1143), .ZN(n1130) );
AND4_X1 U817 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1013) );
NOR4_X1 U818 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1147) );
NOR2_X1 U819 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U820 ( .A(n1154), .B(KEYINPUT25), .Z(n1152) );
INV_X1 U821 ( .A(n1084), .ZN(n1150) );
NAND3_X1 U822 ( .A1(n1155), .A2(n1156), .A3(n1139), .ZN(n1084) );
INV_X1 U823 ( .A(n1157), .ZN(n1148) );
NOR2_X1 U824 ( .A1(n1158), .A2(n982), .ZN(n1146) );
AND3_X1 U825 ( .A1(n1140), .A2(n1156), .A3(n1155), .ZN(n982) );
NOR2_X1 U826 ( .A1(n1036), .A2(G952), .ZN(n1064) );
XNOR2_X1 U827 ( .A(G146), .B(n1131), .ZN(G48) );
NAND4_X1 U828 ( .A1(n1141), .A2(n1139), .A3(n1143), .A4(n1159), .ZN(n1131) );
XOR2_X1 U829 ( .A(G143), .B(n1137), .Z(G45) );
NOR4_X1 U830 ( .A1(n1138), .A2(n1153), .A3(n1160), .A4(n1161), .ZN(n1137) );
XOR2_X1 U831 ( .A(G140), .B(n1136), .Z(G42) );
AND2_X1 U832 ( .A1(n996), .A2(n1162), .ZN(n1136) );
XOR2_X1 U833 ( .A(G137), .B(n1135), .Z(G39) );
AND3_X1 U834 ( .A1(n996), .A2(n1008), .A3(n1141), .ZN(n1135) );
AND2_X1 U835 ( .A1(n1019), .A2(n1159), .ZN(n996) );
XOR2_X1 U836 ( .A(G134), .B(n1163), .Z(G36) );
NOR3_X1 U837 ( .A1(n1164), .A2(n1002), .A3(n1138), .ZN(n1163) );
XOR2_X1 U838 ( .A(KEYINPUT56), .B(n1140), .Z(n1164) );
XNOR2_X1 U839 ( .A(G131), .B(n1165), .ZN(G33) );
NAND2_X1 U840 ( .A1(n1019), .A2(n1166), .ZN(n1165) );
XOR2_X1 U841 ( .A(KEYINPUT7), .B(n1167), .Z(n1166) );
NOR2_X1 U842 ( .A1(n1168), .A2(n1138), .ZN(n1167) );
NAND3_X1 U843 ( .A1(n1159), .A2(n1169), .A3(n1009), .ZN(n1138) );
INV_X1 U844 ( .A(n1002), .ZN(n1019) );
NAND2_X1 U845 ( .A1(n1032), .A2(n999), .ZN(n1002) );
XOR2_X1 U846 ( .A(n1170), .B(n1171), .Z(G30) );
NAND4_X1 U847 ( .A1(n1172), .A2(n1173), .A3(n1142), .A4(n1141), .ZN(n1171) );
AND3_X1 U848 ( .A1(n1174), .A2(n1169), .A3(n1017), .ZN(n1141) );
INV_X1 U849 ( .A(n1175), .ZN(n1017) );
XOR2_X1 U850 ( .A(n1176), .B(KEYINPUT49), .Z(n1173) );
XOR2_X1 U851 ( .A(n1153), .B(KEYINPUT4), .Z(n1172) );
XOR2_X1 U852 ( .A(n1149), .B(n1177), .Z(G3) );
XOR2_X1 U853 ( .A(KEYINPUT42), .B(G101), .Z(n1177) );
AND3_X1 U854 ( .A1(n1008), .A2(n1155), .A3(n1009), .ZN(n1149) );
XOR2_X1 U855 ( .A(n1178), .B(n1134), .Z(G27) );
AND2_X1 U856 ( .A1(n1162), .A2(n995), .ZN(n1134) );
AND4_X1 U857 ( .A1(n1175), .A2(n1139), .A3(n1174), .A4(n1169), .ZN(n1162) );
NAND2_X1 U858 ( .A1(n989), .A2(n1179), .ZN(n1169) );
NAND4_X1 U859 ( .A1(G902), .A2(n1046), .A3(n1180), .A4(n1038), .ZN(n1179) );
INV_X1 U860 ( .A(G900), .ZN(n1038) );
XNOR2_X1 U861 ( .A(G125), .B(KEYINPUT28), .ZN(n1178) );
XOR2_X1 U862 ( .A(G122), .B(n1181), .Z(G24) );
NOR2_X1 U863 ( .A1(n1153), .A2(n1154), .ZN(n1181) );
NAND3_X1 U864 ( .A1(n1182), .A2(n1156), .A3(n1183), .ZN(n1154) );
NOR3_X1 U865 ( .A1(n1160), .A2(n1184), .A3(n1161), .ZN(n1183) );
INV_X1 U866 ( .A(n994), .ZN(n1156) );
NAND2_X1 U867 ( .A1(n1016), .A2(n1175), .ZN(n994) );
XOR2_X1 U868 ( .A(n1185), .B(n1158), .Z(G21) );
AND3_X1 U869 ( .A1(n995), .A2(n1008), .A3(n1186), .ZN(n1158) );
NOR3_X1 U870 ( .A1(n1175), .A2(n1184), .A3(n1016), .ZN(n1186) );
INV_X1 U871 ( .A(n1187), .ZN(n1184) );
NAND2_X1 U872 ( .A1(KEYINPUT6), .A2(n1188), .ZN(n1185) );
INV_X1 U873 ( .A(G119), .ZN(n1188) );
NAND2_X1 U874 ( .A1(n1189), .A2(n1190), .ZN(G18) );
NAND2_X1 U875 ( .A1(G116), .A2(n1157), .ZN(n1190) );
XOR2_X1 U876 ( .A(n1191), .B(KEYINPUT21), .Z(n1189) );
OR2_X1 U877 ( .A1(n1157), .A2(G116), .ZN(n1191) );
NAND4_X1 U878 ( .A1(n1009), .A2(n995), .A3(n1140), .A4(n1187), .ZN(n1157) );
INV_X1 U879 ( .A(n1176), .ZN(n1140) );
NAND2_X1 U880 ( .A1(n1161), .A2(n1192), .ZN(n1176) );
XNOR2_X1 U881 ( .A(G113), .B(n1144), .ZN(G15) );
NAND4_X1 U882 ( .A1(n1009), .A2(n995), .A3(n1139), .A4(n1187), .ZN(n1144) );
INV_X1 U883 ( .A(n1168), .ZN(n1139) );
NAND2_X1 U884 ( .A1(n1193), .A2(n1194), .ZN(n1168) );
INV_X1 U885 ( .A(n1161), .ZN(n1194) );
XOR2_X1 U886 ( .A(KEYINPUT33), .B(n1192), .Z(n1193) );
INV_X1 U887 ( .A(n1160), .ZN(n1192) );
NOR2_X1 U888 ( .A1(n1000), .A2(n1153), .ZN(n995) );
INV_X1 U889 ( .A(n1182), .ZN(n1000) );
NOR2_X1 U890 ( .A1(n1004), .A2(n1195), .ZN(n1182) );
INV_X1 U891 ( .A(n1196), .ZN(n1004) );
NOR2_X1 U892 ( .A1(n1174), .A2(n1175), .ZN(n1009) );
XOR2_X1 U893 ( .A(n1145), .B(n1197), .Z(G12) );
NAND2_X1 U894 ( .A1(n1198), .A2(KEYINPUT2), .ZN(n1197) );
XOR2_X1 U895 ( .A(n1120), .B(KEYINPUT23), .Z(n1198) );
NAND4_X1 U896 ( .A1(n1008), .A2(n1155), .A3(n1175), .A4(n1174), .ZN(n1145) );
INV_X1 U897 ( .A(n1016), .ZN(n1174) );
XNOR2_X1 U898 ( .A(n1199), .B(n1068), .ZN(n1016) );
NAND2_X1 U899 ( .A1(G217), .A2(n1200), .ZN(n1068) );
OR2_X1 U900 ( .A1(n1067), .A2(G902), .ZN(n1199) );
XNOR2_X1 U901 ( .A(n1201), .B(n1202), .ZN(n1067) );
XOR2_X1 U902 ( .A(G110), .B(n1203), .Z(n1202) );
XOR2_X1 U903 ( .A(KEYINPUT9), .B(G119), .Z(n1203) );
XOR2_X1 U904 ( .A(n1204), .B(n1048), .Z(n1201) );
XOR2_X1 U905 ( .A(G140), .B(n1205), .Z(n1048) );
XOR2_X1 U906 ( .A(n1206), .B(n1207), .Z(n1204) );
NAND4_X1 U907 ( .A1(KEYINPUT40), .A2(G221), .A3(G234), .A4(n1036), .ZN(n1206) );
XOR2_X1 U908 ( .A(n1208), .B(G472), .Z(n1175) );
NAND2_X1 U909 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XOR2_X1 U910 ( .A(n1211), .B(n1212), .Z(n1209) );
XOR2_X1 U911 ( .A(n1103), .B(n1102), .Z(n1212) );
XNOR2_X1 U912 ( .A(n1213), .B(KEYINPUT35), .ZN(n1102) );
XOR2_X1 U913 ( .A(n1214), .B(n1215), .Z(n1103) );
XNOR2_X1 U914 ( .A(n1094), .B(n1216), .ZN(n1211) );
XOR2_X1 U915 ( .A(n1092), .B(KEYINPUT60), .Z(n1216) );
INV_X1 U916 ( .A(G101), .ZN(n1092) );
AND3_X1 U917 ( .A1(n1217), .A2(n1036), .A3(G210), .ZN(n1094) );
AND3_X1 U918 ( .A1(n1142), .A2(n1187), .A3(n1143), .ZN(n1155) );
INV_X1 U919 ( .A(n1153), .ZN(n1143) );
NAND2_X1 U920 ( .A1(n1001), .A2(n999), .ZN(n1153) );
NAND2_X1 U921 ( .A1(G214), .A2(n1218), .ZN(n999) );
INV_X1 U922 ( .A(n1032), .ZN(n1001) );
XNOR2_X1 U923 ( .A(n1219), .B(n1128), .ZN(n1032) );
NAND2_X1 U924 ( .A1(G210), .A2(n1218), .ZN(n1128) );
NAND2_X1 U925 ( .A1(n1217), .A2(n1210), .ZN(n1218) );
NAND2_X1 U926 ( .A1(n1125), .A2(n1210), .ZN(n1219) );
XNOR2_X1 U927 ( .A(n1220), .B(n1221), .ZN(n1125) );
XOR2_X1 U928 ( .A(n1215), .B(n1222), .Z(n1221) );
XOR2_X1 U929 ( .A(n1223), .B(n1224), .Z(n1222) );
NOR2_X1 U930 ( .A1(G953), .A2(n1052), .ZN(n1223) );
INV_X1 U931 ( .A(G224), .ZN(n1052) );
XOR2_X1 U932 ( .A(G143), .B(KEYINPUT48), .Z(n1215) );
XOR2_X1 U933 ( .A(n1225), .B(n1205), .Z(n1220) );
NAND2_X1 U934 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
OR2_X1 U935 ( .A1(n1062), .A2(n1063), .ZN(n1227) );
NAND2_X1 U936 ( .A1(n1063), .A2(n1228), .ZN(n1226) );
XOR2_X1 U937 ( .A(n1062), .B(KEYINPUT52), .Z(n1228) );
XOR2_X1 U938 ( .A(n1229), .B(n1230), .Z(n1062) );
XOR2_X1 U939 ( .A(n1231), .B(n1232), .Z(n1230) );
XNOR2_X1 U940 ( .A(KEYINPUT43), .B(KEYINPUT24), .ZN(n1232) );
XOR2_X1 U941 ( .A(n1213), .B(G110), .Z(n1229) );
XNOR2_X1 U942 ( .A(G113), .B(n1233), .ZN(n1213) );
XOR2_X1 U943 ( .A(G119), .B(G116), .Z(n1233) );
XNOR2_X1 U944 ( .A(n1234), .B(n1235), .ZN(n1063) );
NAND2_X1 U945 ( .A1(n1236), .A2(n1237), .ZN(n1234) );
XOR2_X1 U946 ( .A(G107), .B(G104), .Z(n1237) );
XNOR2_X1 U947 ( .A(KEYINPUT61), .B(KEYINPUT58), .ZN(n1236) );
NAND2_X1 U948 ( .A1(n989), .A2(n1238), .ZN(n1187) );
NAND4_X1 U949 ( .A1(G902), .A2(n1046), .A3(n1180), .A4(n1053), .ZN(n1238) );
INV_X1 U950 ( .A(G898), .ZN(n1053) );
XOR2_X1 U951 ( .A(G953), .B(KEYINPUT41), .Z(n1046) );
NAND3_X1 U952 ( .A1(n1180), .A2(n1036), .A3(G952), .ZN(n989) );
NAND2_X1 U953 ( .A1(G237), .A2(G234), .ZN(n1180) );
XNOR2_X1 U954 ( .A(n1159), .B(KEYINPUT38), .ZN(n1142) );
NOR2_X1 U955 ( .A1(n1195), .A2(n1196), .ZN(n1159) );
XOR2_X1 U956 ( .A(n1028), .B(n1239), .Z(n1196) );
XOR2_X1 U957 ( .A(KEYINPUT20), .B(G469), .Z(n1239) );
NAND2_X1 U958 ( .A1(n1240), .A2(n1210), .ZN(n1028) );
XOR2_X1 U959 ( .A(n1241), .B(n1242), .Z(n1240) );
INV_X1 U960 ( .A(n1121), .ZN(n1242) );
XOR2_X1 U961 ( .A(n1243), .B(n1244), .Z(n1121) );
XOR2_X1 U962 ( .A(G107), .B(n1245), .Z(n1244) );
NOR2_X1 U963 ( .A1(G104), .A2(KEYINPUT10), .ZN(n1245) );
XOR2_X1 U964 ( .A(n1047), .B(n1246), .Z(n1243) );
NOR2_X1 U965 ( .A1(KEYINPUT1), .A2(n1235), .ZN(n1246) );
XOR2_X1 U966 ( .A(G101), .B(KEYINPUT27), .Z(n1235) );
XOR2_X1 U967 ( .A(n1247), .B(n1214), .Z(n1047) );
XNOR2_X1 U968 ( .A(n1248), .B(n1249), .ZN(n1214) );
XOR2_X1 U969 ( .A(KEYINPUT18), .B(G131), .Z(n1249) );
XOR2_X1 U970 ( .A(n1207), .B(n1250), .Z(n1248) );
XOR2_X1 U971 ( .A(G137), .B(n1224), .Z(n1207) );
XOR2_X1 U972 ( .A(G128), .B(G146), .Z(n1224) );
NAND2_X1 U973 ( .A1(KEYINPUT30), .A2(G143), .ZN(n1247) );
NAND2_X1 U974 ( .A1(n1251), .A2(KEYINPUT39), .ZN(n1241) );
XOR2_X1 U975 ( .A(n1252), .B(n1109), .Z(n1251) );
NOR2_X1 U976 ( .A1(n1037), .A2(G953), .ZN(n1109) );
INV_X1 U977 ( .A(G227), .ZN(n1037) );
NAND3_X1 U978 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1252) );
XOR2_X1 U979 ( .A(KEYINPUT29), .B(n1256), .Z(n1255) );
NOR2_X1 U980 ( .A1(G140), .A2(n1257), .ZN(n1256) );
XOR2_X1 U981 ( .A(KEYINPUT8), .B(G110), .Z(n1257) );
OR3_X1 U982 ( .A1(n1116), .A2(n1120), .A3(KEYINPUT8), .ZN(n1254) );
INV_X1 U983 ( .A(G140), .ZN(n1116) );
NAND2_X1 U984 ( .A1(n1258), .A2(KEYINPUT8), .ZN(n1253) );
INV_X1 U985 ( .A(n1112), .ZN(n1258) );
NAND2_X1 U986 ( .A1(G140), .A2(n1120), .ZN(n1112) );
INV_X1 U987 ( .A(G110), .ZN(n1120) );
XNOR2_X1 U988 ( .A(n1025), .B(KEYINPUT31), .ZN(n1195) );
INV_X1 U989 ( .A(n1003), .ZN(n1025) );
NAND2_X1 U990 ( .A1(G221), .A2(n1200), .ZN(n1003) );
NAND2_X1 U991 ( .A1(G234), .A2(n1210), .ZN(n1200) );
INV_X1 U992 ( .A(n992), .ZN(n1008) );
NAND2_X1 U993 ( .A1(n1160), .A2(n1161), .ZN(n992) );
XOR2_X1 U994 ( .A(n1081), .B(n1259), .Z(n1161) );
NOR2_X1 U995 ( .A1(KEYINPUT37), .A2(n1030), .ZN(n1259) );
NAND2_X1 U996 ( .A1(n1260), .A2(n1210), .ZN(n1030) );
XOR2_X1 U997 ( .A(KEYINPUT54), .B(n1080), .Z(n1260) );
XNOR2_X1 U998 ( .A(n1261), .B(n1262), .ZN(n1080) );
XOR2_X1 U999 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U1000 ( .A(n1265), .B(n1266), .ZN(n1264) );
NOR2_X1 U1001 ( .A1(KEYINPUT34), .A2(n1267), .ZN(n1266) );
INV_X1 U1002 ( .A(G104), .ZN(n1267) );
NOR2_X1 U1003 ( .A1(KEYINPUT3), .A2(n1268), .ZN(n1265) );
XNOR2_X1 U1004 ( .A(n1205), .B(n1269), .ZN(n1268) );
XNOR2_X1 U1005 ( .A(G146), .B(n1270), .ZN(n1269) );
NOR2_X1 U1006 ( .A1(G140), .A2(KEYINPUT36), .ZN(n1270) );
XOR2_X1 U1007 ( .A(G125), .B(KEYINPUT0), .Z(n1205) );
NAND3_X1 U1008 ( .A1(n1217), .A2(n1036), .A3(G214), .ZN(n1263) );
INV_X1 U1009 ( .A(G237), .ZN(n1217) );
XOR2_X1 U1010 ( .A(n1271), .B(n1272), .Z(n1261) );
XOR2_X1 U1011 ( .A(G143), .B(G131), .Z(n1272) );
XOR2_X1 U1012 ( .A(G113), .B(n1231), .Z(n1271) );
INV_X1 U1013 ( .A(G122), .ZN(n1231) );
INV_X1 U1014 ( .A(G475), .ZN(n1081) );
XOR2_X1 U1015 ( .A(n1031), .B(KEYINPUT51), .Z(n1160) );
XOR2_X1 U1016 ( .A(n1273), .B(G478), .Z(n1031) );
NAND2_X1 U1017 ( .A1(n1210), .A2(n1074), .ZN(n1273) );
NAND2_X1 U1018 ( .A1(n1274), .A2(n1275), .ZN(n1074) );
NAND4_X1 U1019 ( .A1(n1276), .A2(n1036), .A3(n1277), .A4(n1278), .ZN(n1275) );
AND2_X1 U1020 ( .A1(G234), .A2(G217), .ZN(n1278) );
NAND2_X1 U1021 ( .A1(n1279), .A2(n1280), .ZN(n1274) );
NAND3_X1 U1022 ( .A1(G234), .A2(n1036), .A3(G217), .ZN(n1280) );
INV_X1 U1023 ( .A(G953), .ZN(n1036) );
NAND2_X1 U1024 ( .A1(n1277), .A2(n1276), .ZN(n1279) );
NAND2_X1 U1025 ( .A1(n1281), .A2(n1282), .ZN(n1276) );
XOR2_X1 U1026 ( .A(n1283), .B(n1284), .Z(n1281) );
NAND2_X1 U1027 ( .A1(n1285), .A2(n1286), .ZN(n1277) );
XNOR2_X1 U1028 ( .A(n1283), .B(n1284), .ZN(n1286) );
XOR2_X1 U1029 ( .A(n1170), .B(n1287), .Z(n1284) );
INV_X1 U1030 ( .A(G143), .ZN(n1287) );
INV_X1 U1031 ( .A(G128), .ZN(n1170) );
NAND2_X1 U1032 ( .A1(KEYINPUT5), .A2(n1250), .ZN(n1283) );
XNOR2_X1 U1033 ( .A(G134), .B(KEYINPUT13), .ZN(n1250) );
INV_X1 U1034 ( .A(n1282), .ZN(n1285) );
NAND2_X1 U1035 ( .A1(n1288), .A2(n1289), .ZN(n1282) );
NAND2_X1 U1036 ( .A1(G107), .A2(n1290), .ZN(n1289) );
XOR2_X1 U1037 ( .A(KEYINPUT11), .B(n1291), .Z(n1288) );
NOR2_X1 U1038 ( .A1(G107), .A2(n1292), .ZN(n1291) );
XNOR2_X1 U1039 ( .A(n1290), .B(KEYINPUT17), .ZN(n1292) );
XOR2_X1 U1040 ( .A(G116), .B(G122), .Z(n1290) );
INV_X1 U1041 ( .A(G902), .ZN(n1210) );
endmodule


