//Key = 0101011111010100111111110100011100001010111001100101011101011011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269;

XOR2_X1 U705 ( .A(G107), .B(n971), .Z(G9) );
NOR2_X1 U706 ( .A1(n972), .A2(n973), .ZN(G75) );
NOR4_X1 U707 ( .A1(n974), .A2(n975), .A3(n976), .A4(n977), .ZN(n973) );
NOR2_X1 U708 ( .A1(n978), .A2(n979), .ZN(n975) );
NOR2_X1 U709 ( .A1(n980), .A2(n981), .ZN(n978) );
NOR2_X1 U710 ( .A1(n982), .A2(n983), .ZN(n981) );
NOR2_X1 U711 ( .A1(n984), .A2(n985), .ZN(n982) );
NOR2_X1 U712 ( .A1(n986), .A2(n987), .ZN(n985) );
NOR2_X1 U713 ( .A1(n988), .A2(n989), .ZN(n986) );
NOR2_X1 U714 ( .A1(n990), .A2(n991), .ZN(n989) );
NOR2_X1 U715 ( .A1(n992), .A2(n993), .ZN(n990) );
AND2_X1 U716 ( .A1(n994), .A2(n995), .ZN(n992) );
NOR2_X1 U717 ( .A1(n996), .A2(n997), .ZN(n988) );
NOR2_X1 U718 ( .A1(n998), .A2(n999), .ZN(n996) );
NOR2_X1 U719 ( .A1(n1000), .A2(n1001), .ZN(n998) );
NOR3_X1 U720 ( .A1(n997), .A2(n1002), .A3(n991), .ZN(n984) );
NOR2_X1 U721 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
AND2_X1 U722 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
NOR4_X1 U723 ( .A1(n1007), .A2(n991), .A3(n987), .A4(n997), .ZN(n980) );
NOR2_X1 U724 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NOR3_X1 U725 ( .A1(n976), .A2(G952), .A3(n974), .ZN(n972) );
AND4_X1 U726 ( .A1(n1010), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n974) );
NOR3_X1 U727 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
XOR2_X1 U728 ( .A(KEYINPUT15), .B(n1017), .Z(n1016) );
NOR2_X1 U729 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
XOR2_X1 U730 ( .A(n1020), .B(n1021), .Z(n1015) );
NAND3_X1 U731 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1014) );
XOR2_X1 U732 ( .A(KEYINPUT49), .B(n1025), .Z(n1024) );
NOR2_X1 U733 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
XOR2_X1 U734 ( .A(n1028), .B(KEYINPUT17), .Z(n1027) );
XOR2_X1 U735 ( .A(n1029), .B(n1030), .Z(n1023) );
NAND2_X1 U736 ( .A1(KEYINPUT11), .A2(n1031), .ZN(n1030) );
XOR2_X1 U737 ( .A(KEYINPUT36), .B(n1032), .Z(n1022) );
NOR3_X1 U738 ( .A1(n1033), .A2(n1006), .A3(n995), .ZN(n1012) );
NOR3_X1 U739 ( .A1(n1034), .A2(G902), .A3(n1028), .ZN(n1033) );
XNOR2_X1 U740 ( .A(G469), .B(KEYINPUT41), .ZN(n1028) );
NAND2_X1 U741 ( .A1(n1018), .A2(n1019), .ZN(n1011) );
XNOR2_X1 U742 ( .A(KEYINPUT42), .B(G472), .ZN(n1018) );
XOR2_X1 U743 ( .A(KEYINPUT14), .B(n1035), .Z(n1010) );
NOR3_X1 U744 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NOR3_X1 U745 ( .A1(n1039), .A2(KEYINPUT10), .A3(n1040), .ZN(n1038) );
AND2_X1 U746 ( .A1(n1039), .A2(KEYINPUT10), .ZN(n1037) );
XOR2_X1 U747 ( .A(n1041), .B(n1042), .Z(G72) );
NOR2_X1 U748 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U749 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U750 ( .A1(G227), .A2(n1047), .ZN(n1045) );
NOR2_X1 U751 ( .A1(n1048), .A2(n1047), .ZN(n1043) );
NOR2_X1 U752 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U753 ( .A1(G227), .A2(n1051), .ZN(n1049) );
INV_X1 U754 ( .A(n1046), .ZN(n1051) );
XOR2_X1 U755 ( .A(n1052), .B(n1053), .Z(n1046) );
XOR2_X1 U756 ( .A(G140), .B(G125), .Z(n1053) );
XOR2_X1 U757 ( .A(n1054), .B(n1055), .Z(n1052) );
NOR2_X1 U758 ( .A1(KEYINPUT48), .A2(n1056), .ZN(n1055) );
NAND2_X1 U759 ( .A1(n1047), .A2(n1057), .ZN(n1041) );
NAND2_X1 U760 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U761 ( .A1(n1060), .A2(n1061), .ZN(G69) );
NAND3_X1 U762 ( .A1(n1062), .A2(n1063), .A3(G953), .ZN(n1061) );
XOR2_X1 U763 ( .A(n1064), .B(KEYINPUT24), .Z(n1060) );
NAND3_X1 U764 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NAND2_X1 U765 ( .A1(n1068), .A2(n1063), .ZN(n1067) );
OR3_X1 U766 ( .A1(n1063), .A2(n1068), .A3(G953), .ZN(n1066) );
NAND2_X1 U767 ( .A1(G953), .A2(n1069), .ZN(n1065) );
OR2_X1 U768 ( .A1(n1063), .A2(n1062), .ZN(n1069) );
NAND2_X1 U769 ( .A1(G898), .A2(G224), .ZN(n1062) );
NAND2_X1 U770 ( .A1(n1070), .A2(n1071), .ZN(n1063) );
NAND2_X1 U771 ( .A1(n1072), .A2(G953), .ZN(n1071) );
XNOR2_X1 U772 ( .A(G898), .B(KEYINPUT37), .ZN(n1072) );
XOR2_X1 U773 ( .A(n1073), .B(n1074), .Z(n1070) );
NAND2_X1 U774 ( .A1(KEYINPUT5), .A2(n1075), .ZN(n1074) );
NAND2_X1 U775 ( .A1(n1076), .A2(n1077), .ZN(n1073) );
XOR2_X1 U776 ( .A(n1078), .B(KEYINPUT52), .Z(n1076) );
NOR2_X1 U777 ( .A1(n1079), .A2(n1080), .ZN(G66) );
NOR2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XOR2_X1 U779 ( .A(n1083), .B(KEYINPUT38), .Z(n1082) );
NAND2_X1 U780 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U781 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
NAND2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XNOR2_X1 U783 ( .A(G217), .B(KEYINPUT51), .ZN(n1086) );
NOR2_X1 U784 ( .A1(n1079), .A2(n1088), .ZN(G63) );
XOR2_X1 U785 ( .A(n1089), .B(n1090), .Z(n1088) );
NAND3_X1 U786 ( .A1(n1087), .A2(G478), .A3(KEYINPUT29), .ZN(n1089) );
NOR2_X1 U787 ( .A1(n1079), .A2(n1091), .ZN(G60) );
XNOR2_X1 U788 ( .A(n1092), .B(n1093), .ZN(n1091) );
NOR4_X1 U789 ( .A1(n1094), .A2(n1095), .A3(KEYINPUT61), .A4(n1020), .ZN(n1093) );
INV_X1 U790 ( .A(G475), .ZN(n1020) );
NOR2_X1 U791 ( .A1(KEYINPUT55), .A2(n1096), .ZN(n1095) );
AND2_X1 U792 ( .A1(n1097), .A2(n977), .ZN(n1096) );
AND2_X1 U793 ( .A1(n1098), .A2(KEYINPUT55), .ZN(n1094) );
XOR2_X1 U794 ( .A(G104), .B(n1099), .Z(G6) );
NOR2_X1 U795 ( .A1(n1079), .A2(n1100), .ZN(G57) );
XOR2_X1 U796 ( .A(n1101), .B(n1102), .Z(n1100) );
XOR2_X1 U797 ( .A(n1103), .B(n1104), .Z(n1102) );
AND2_X1 U798 ( .A1(G472), .A2(n1087), .ZN(n1103) );
XOR2_X1 U799 ( .A(n1105), .B(n1106), .Z(n1101) );
NOR2_X1 U800 ( .A1(n1079), .A2(n1107), .ZN(G54) );
XOR2_X1 U801 ( .A(n1108), .B(n1034), .Z(n1107) );
AND2_X1 U802 ( .A1(G469), .A2(n1087), .ZN(n1108) );
INV_X1 U803 ( .A(n1098), .ZN(n1087) );
NOR2_X1 U804 ( .A1(n1079), .A2(n1109), .ZN(G51) );
XNOR2_X1 U805 ( .A(n1110), .B(n1111), .ZN(n1109) );
XOR2_X1 U806 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U807 ( .A1(n1029), .A2(n1098), .ZN(n1113) );
NAND2_X1 U808 ( .A1(G902), .A2(n977), .ZN(n1098) );
NAND3_X1 U809 ( .A1(n1058), .A2(n1114), .A3(n1068), .ZN(n977) );
AND2_X1 U810 ( .A1(n1115), .A2(n1116), .ZN(n1068) );
NOR4_X1 U811 ( .A1(n971), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1116) );
AND3_X1 U812 ( .A1(n1120), .A2(n1121), .A3(n1008), .ZN(n971) );
NOR4_X1 U813 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1099), .ZN(n1115) );
AND3_X1 U814 ( .A1(n1120), .A2(n1121), .A3(n1009), .ZN(n1099) );
INV_X1 U815 ( .A(n1125), .ZN(n1121) );
NOR3_X1 U816 ( .A1(n1126), .A2(n1125), .A3(n1127), .ZN(n1124) );
XOR2_X1 U817 ( .A(KEYINPUT30), .B(n1128), .Z(n1126) );
INV_X1 U818 ( .A(n1129), .ZN(n1123) );
XNOR2_X1 U819 ( .A(KEYINPUT20), .B(n1059), .ZN(n1114) );
AND4_X1 U820 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1058) );
AND4_X1 U821 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1133) );
NAND3_X1 U822 ( .A1(n1138), .A2(n993), .A3(n1139), .ZN(n1132) );
NAND2_X1 U823 ( .A1(KEYINPUT18), .A2(n1140), .ZN(n1112) );
NOR2_X1 U824 ( .A1(n1047), .A2(G952), .ZN(n1079) );
XNOR2_X1 U825 ( .A(G146), .B(n1130), .ZN(G48) );
NAND3_X1 U826 ( .A1(n1009), .A2(n993), .A3(n1141), .ZN(n1130) );
XOR2_X1 U827 ( .A(n1142), .B(n1131), .Z(G45) );
NAND4_X1 U828 ( .A1(n1143), .A2(n993), .A3(n1032), .A4(n1144), .ZN(n1131) );
XOR2_X1 U829 ( .A(n1145), .B(n1137), .Z(G42) );
NAND3_X1 U830 ( .A1(n1146), .A2(n1004), .A3(n1139), .ZN(n1137) );
XOR2_X1 U831 ( .A(n1059), .B(n1147), .Z(G39) );
XOR2_X1 U832 ( .A(n1148), .B(KEYINPUT39), .Z(n1147) );
NAND3_X1 U833 ( .A1(n1141), .A2(n1128), .A3(n1146), .ZN(n1059) );
XOR2_X1 U834 ( .A(n1136), .B(n1149), .Z(G36) );
NAND2_X1 U835 ( .A1(KEYINPUT3), .A2(G134), .ZN(n1149) );
NAND3_X1 U836 ( .A1(n1143), .A2(n1008), .A3(n1146), .ZN(n1136) );
XNOR2_X1 U837 ( .A(G131), .B(n1135), .ZN(G33) );
NAND3_X1 U838 ( .A1(n1143), .A2(n1009), .A3(n1146), .ZN(n1135) );
INV_X1 U839 ( .A(n997), .ZN(n1146) );
NAND2_X1 U840 ( .A1(n994), .A2(n1150), .ZN(n997) );
AND3_X1 U841 ( .A1(n1004), .A2(n1151), .A3(n999), .ZN(n1143) );
XOR2_X1 U842 ( .A(n1152), .B(n1134), .Z(G30) );
NAND3_X1 U843 ( .A1(n1008), .A2(n993), .A3(n1141), .ZN(n1134) );
AND4_X1 U844 ( .A1(n1004), .A2(n1151), .A3(n1153), .A4(n1001), .ZN(n1141) );
XOR2_X1 U845 ( .A(n1105), .B(n1154), .Z(G3) );
NAND2_X1 U846 ( .A1(n999), .A2(n1155), .ZN(n1154) );
XNOR2_X1 U847 ( .A(G125), .B(n1156), .ZN(G27) );
NAND3_X1 U848 ( .A1(n993), .A2(n1157), .A3(n1139), .ZN(n1156) );
AND4_X1 U849 ( .A1(n1009), .A2(n1158), .A3(n1151), .A4(n1153), .ZN(n1139) );
NAND2_X1 U850 ( .A1(n979), .A2(n1159), .ZN(n1151) );
NAND4_X1 U851 ( .A1(G953), .A2(G902), .A3(n1160), .A4(n1050), .ZN(n1159) );
INV_X1 U852 ( .A(G900), .ZN(n1050) );
XOR2_X1 U853 ( .A(KEYINPUT12), .B(n1138), .Z(n1157) );
XOR2_X1 U854 ( .A(n1161), .B(n1129), .Z(G24) );
NAND4_X1 U855 ( .A1(n1162), .A2(n1120), .A3(n1032), .A4(n1144), .ZN(n1129) );
INV_X1 U856 ( .A(n991), .ZN(n1120) );
NAND2_X1 U857 ( .A1(n1158), .A2(n1000), .ZN(n991) );
XOR2_X1 U858 ( .A(G119), .B(n1122), .Z(G21) );
AND4_X1 U859 ( .A1(n1162), .A2(n1128), .A3(n1153), .A4(n1001), .ZN(n1122) );
INV_X1 U860 ( .A(n983), .ZN(n1128) );
XOR2_X1 U861 ( .A(G116), .B(n1119), .Z(G18) );
AND3_X1 U862 ( .A1(n1162), .A2(n1008), .A3(n999), .ZN(n1119) );
NOR2_X1 U863 ( .A1(n1144), .A2(n1163), .ZN(n1008) );
INV_X1 U864 ( .A(n1164), .ZN(n1144) );
XOR2_X1 U865 ( .A(G113), .B(n1118), .Z(G15) );
AND3_X1 U866 ( .A1(n1009), .A2(n1162), .A3(n999), .ZN(n1118) );
INV_X1 U867 ( .A(n1127), .ZN(n999) );
NAND2_X1 U868 ( .A1(n1000), .A2(n1001), .ZN(n1127) );
AND3_X1 U869 ( .A1(n993), .A2(n1165), .A3(n1138), .ZN(n1162) );
INV_X1 U870 ( .A(n987), .ZN(n1138) );
NAND2_X1 U871 ( .A1(n1005), .A2(n1166), .ZN(n987) );
NOR2_X1 U872 ( .A1(n1032), .A2(n1164), .ZN(n1009) );
INV_X1 U873 ( .A(n1163), .ZN(n1032) );
XOR2_X1 U874 ( .A(G110), .B(n1117), .Z(G12) );
AND3_X1 U875 ( .A1(n1158), .A2(n1153), .A3(n1155), .ZN(n1117) );
NOR2_X1 U876 ( .A1(n983), .A2(n1125), .ZN(n1155) );
NAND3_X1 U877 ( .A1(n993), .A2(n1165), .A3(n1004), .ZN(n1125) );
NOR2_X1 U878 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
INV_X1 U879 ( .A(n1166), .ZN(n1006) );
NAND2_X1 U880 ( .A1(G221), .A2(n1167), .ZN(n1166) );
XOR2_X1 U881 ( .A(n1168), .B(n1169), .Z(n1005) );
NOR2_X1 U882 ( .A1(KEYINPUT0), .A2(n1026), .ZN(n1169) );
NOR2_X1 U883 ( .A1(G902), .A2(n1034), .ZN(n1026) );
XNOR2_X1 U884 ( .A(n1170), .B(n1171), .ZN(n1034) );
XNOR2_X1 U885 ( .A(G107), .B(n1172), .ZN(n1171) );
NAND2_X1 U886 ( .A1(KEYINPUT1), .A2(n1105), .ZN(n1172) );
XOR2_X1 U887 ( .A(n1173), .B(n1174), .Z(n1170) );
XOR2_X1 U888 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U889 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U890 ( .A(G140), .B(G110), .Z(n1178) );
XOR2_X1 U891 ( .A(n1179), .B(n1180), .Z(n1177) );
NAND2_X1 U892 ( .A1(G227), .A2(n1047), .ZN(n1179) );
XOR2_X1 U893 ( .A(n1181), .B(n1182), .Z(n1175) );
XOR2_X1 U894 ( .A(KEYINPUT63), .B(KEYINPUT58), .Z(n1182) );
XNOR2_X1 U895 ( .A(KEYINPUT57), .B(KEYINPUT19), .ZN(n1181) );
XNOR2_X1 U896 ( .A(G469), .B(KEYINPUT8), .ZN(n1168) );
NAND2_X1 U897 ( .A1(n979), .A2(n1183), .ZN(n1165) );
NAND4_X1 U898 ( .A1(n1184), .A2(G953), .A3(G902), .A4(n1160), .ZN(n1183) );
XNOR2_X1 U899 ( .A(G898), .B(KEYINPUT43), .ZN(n1184) );
NAND3_X1 U900 ( .A1(n1185), .A2(n1160), .A3(G952), .ZN(n979) );
NAND2_X1 U901 ( .A1(G237), .A2(G234), .ZN(n1160) );
INV_X1 U902 ( .A(n976), .ZN(n1185) );
XOR2_X1 U903 ( .A(n1047), .B(KEYINPUT40), .Z(n976) );
NOR2_X1 U904 ( .A1(n994), .A2(n995), .ZN(n993) );
INV_X1 U905 ( .A(n1150), .ZN(n995) );
NAND2_X1 U906 ( .A1(G214), .A2(n1186), .ZN(n1150) );
XNOR2_X1 U907 ( .A(n1031), .B(n1029), .ZN(n994) );
NAND2_X1 U908 ( .A1(G210), .A2(n1186), .ZN(n1029) );
NAND2_X1 U909 ( .A1(n1187), .A2(n1097), .ZN(n1186) );
NAND2_X1 U910 ( .A1(n1188), .A2(n1097), .ZN(n1031) );
XNOR2_X1 U911 ( .A(n1140), .B(n1110), .ZN(n1188) );
XOR2_X1 U912 ( .A(n1075), .B(n1189), .Z(n1110) );
XOR2_X1 U913 ( .A(n1190), .B(n1191), .Z(n1189) );
AND2_X1 U914 ( .A1(n1047), .A2(G224), .ZN(n1191) );
NOR2_X1 U915 ( .A1(KEYINPUT26), .A2(n1192), .ZN(n1190) );
NOR2_X1 U916 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XOR2_X1 U917 ( .A(n1078), .B(KEYINPUT7), .Z(n1194) );
NAND2_X1 U918 ( .A1(n1195), .A2(n1196), .ZN(n1078) );
XOR2_X1 U919 ( .A(n1197), .B(n1198), .Z(n1196) );
INV_X1 U920 ( .A(G113), .ZN(n1197) );
XOR2_X1 U921 ( .A(n1199), .B(n1200), .Z(n1195) );
INV_X1 U922 ( .A(n1077), .ZN(n1193) );
NAND2_X1 U923 ( .A1(n1201), .A2(n1202), .ZN(n1077) );
XOR2_X1 U924 ( .A(G113), .B(n1198), .Z(n1202) );
NOR2_X1 U925 ( .A1(KEYINPUT44), .A2(n1203), .ZN(n1198) );
XNOR2_X1 U926 ( .A(n1200), .B(n1199), .ZN(n1201) );
NAND2_X1 U927 ( .A1(n1204), .A2(n1205), .ZN(n1199) );
NAND2_X1 U928 ( .A1(G107), .A2(n1180), .ZN(n1205) );
XOR2_X1 U929 ( .A(n1206), .B(KEYINPUT4), .Z(n1204) );
OR2_X1 U930 ( .A1(n1180), .A2(G107), .ZN(n1206) );
XOR2_X1 U931 ( .A(G104), .B(KEYINPUT53), .Z(n1180) );
NOR2_X1 U932 ( .A1(KEYINPUT35), .A2(n1105), .ZN(n1200) );
XOR2_X1 U933 ( .A(G110), .B(n1207), .Z(n1075) );
XOR2_X1 U934 ( .A(KEYINPUT45), .B(G122), .Z(n1207) );
XOR2_X1 U935 ( .A(n1054), .B(G125), .Z(n1140) );
NAND2_X1 U936 ( .A1(n1163), .A2(n1164), .ZN(n983) );
XOR2_X1 U937 ( .A(n1021), .B(n1208), .Z(n1164) );
XOR2_X1 U938 ( .A(KEYINPUT25), .B(n1209), .Z(n1208) );
NOR2_X1 U939 ( .A1(KEYINPUT27), .A2(G475), .ZN(n1209) );
NAND2_X1 U940 ( .A1(n1092), .A2(n1097), .ZN(n1021) );
XNOR2_X1 U941 ( .A(n1210), .B(n1211), .ZN(n1092) );
XOR2_X1 U942 ( .A(n1212), .B(n1213), .Z(n1211) );
XOR2_X1 U943 ( .A(n1214), .B(n1215), .Z(n1213) );
NOR2_X1 U944 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
XOR2_X1 U945 ( .A(n1218), .B(KEYINPUT31), .Z(n1217) );
NAND2_X1 U946 ( .A1(n1219), .A2(n1161), .ZN(n1218) );
XOR2_X1 U947 ( .A(KEYINPUT50), .B(G113), .Z(n1219) );
NOR2_X1 U948 ( .A1(G113), .A2(n1161), .ZN(n1216) );
INV_X1 U949 ( .A(G122), .ZN(n1161) );
NAND2_X1 U950 ( .A1(KEYINPUT13), .A2(n1220), .ZN(n1214) );
XOR2_X1 U951 ( .A(n1221), .B(n1222), .Z(n1220) );
XNOR2_X1 U952 ( .A(G146), .B(G125), .ZN(n1222) );
NAND2_X1 U953 ( .A1(KEYINPUT22), .A2(n1145), .ZN(n1221) );
INV_X1 U954 ( .A(G140), .ZN(n1145) );
NAND3_X1 U955 ( .A1(n1187), .A2(n1047), .A3(G214), .ZN(n1212) );
XNOR2_X1 U956 ( .A(G104), .B(n1223), .ZN(n1210) );
XOR2_X1 U957 ( .A(G143), .B(G131), .Z(n1223) );
XOR2_X1 U958 ( .A(n1224), .B(G478), .Z(n1163) );
NAND2_X1 U959 ( .A1(n1090), .A2(n1097), .ZN(n1224) );
XOR2_X1 U960 ( .A(n1225), .B(n1226), .Z(n1090) );
XOR2_X1 U961 ( .A(n1227), .B(n1228), .Z(n1226) );
NAND3_X1 U962 ( .A1(G217), .A2(n1047), .A3(G234), .ZN(n1228) );
NAND2_X1 U963 ( .A1(n1229), .A2(KEYINPUT60), .ZN(n1227) );
XOR2_X1 U964 ( .A(n1230), .B(n1231), .Z(n1229) );
XOR2_X1 U965 ( .A(KEYINPUT33), .B(G122), .Z(n1231) );
INV_X1 U966 ( .A(G116), .ZN(n1230) );
XOR2_X1 U967 ( .A(n1232), .B(n1233), .Z(n1225) );
XOR2_X1 U968 ( .A(G134), .B(G107), .Z(n1233) );
NAND2_X1 U969 ( .A1(n1234), .A2(KEYINPUT62), .ZN(n1232) );
XNOR2_X1 U970 ( .A(n1235), .B(KEYINPUT46), .ZN(n1234) );
INV_X1 U971 ( .A(n1000), .ZN(n1153) );
NOR2_X1 U972 ( .A1(n1036), .A2(n1236), .ZN(n1000) );
NOR2_X1 U973 ( .A1(n1039), .A2(n1040), .ZN(n1236) );
AND2_X1 U974 ( .A1(n1040), .A2(n1039), .ZN(n1036) );
NAND2_X1 U975 ( .A1(G217), .A2(n1167), .ZN(n1039) );
NAND2_X1 U976 ( .A1(G234), .A2(n1097), .ZN(n1167) );
AND2_X1 U977 ( .A1(n1084), .A2(n1097), .ZN(n1040) );
XNOR2_X1 U978 ( .A(n1237), .B(n1238), .ZN(n1084) );
XOR2_X1 U979 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U980 ( .A(n1241), .B(G110), .Z(n1240) );
NAND2_X1 U981 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND2_X1 U982 ( .A1(n1244), .A2(G146), .ZN(n1243) );
XOR2_X1 U983 ( .A(KEYINPUT6), .B(n1245), .Z(n1242) );
NOR2_X1 U984 ( .A1(G146), .A2(n1244), .ZN(n1245) );
XNOR2_X1 U985 ( .A(G125), .B(n1246), .ZN(n1244) );
NOR2_X1 U986 ( .A1(G140), .A2(KEYINPUT47), .ZN(n1246) );
NAND2_X1 U987 ( .A1(n1247), .A2(n1248), .ZN(n1239) );
NAND2_X1 U988 ( .A1(n1249), .A2(n1148), .ZN(n1248) );
XOR2_X1 U989 ( .A(n1250), .B(KEYINPUT2), .Z(n1247) );
OR2_X1 U990 ( .A1(n1249), .A2(n1148), .ZN(n1250) );
INV_X1 U991 ( .A(G137), .ZN(n1148) );
NAND3_X1 U992 ( .A1(n1251), .A2(n1047), .A3(G234), .ZN(n1249) );
XOR2_X1 U993 ( .A(KEYINPUT34), .B(G221), .Z(n1251) );
XNOR2_X1 U994 ( .A(G119), .B(n1252), .ZN(n1237) );
XOR2_X1 U995 ( .A(KEYINPUT28), .B(G128), .Z(n1252) );
INV_X1 U996 ( .A(n1001), .ZN(n1158) );
NAND2_X1 U997 ( .A1(n1253), .A2(n1254), .ZN(n1001) );
OR2_X1 U998 ( .A1(n1019), .A2(G472), .ZN(n1254) );
XOR2_X1 U999 ( .A(n1255), .B(KEYINPUT32), .Z(n1253) );
NAND2_X1 U1000 ( .A1(G472), .A2(n1019), .ZN(n1255) );
NAND2_X1 U1001 ( .A1(n1256), .A2(n1097), .ZN(n1019) );
INV_X1 U1002 ( .A(G902), .ZN(n1097) );
XNOR2_X1 U1003 ( .A(n1104), .B(n1257), .ZN(n1256) );
NOR2_X1 U1004 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XOR2_X1 U1005 ( .A(n1260), .B(KEYINPUT16), .Z(n1259) );
OR2_X1 U1006 ( .A1(n1105), .A2(n1106), .ZN(n1260) );
INV_X1 U1007 ( .A(G101), .ZN(n1105) );
NOR2_X1 U1008 ( .A1(n1261), .A2(n1262), .ZN(n1258) );
XOR2_X1 U1009 ( .A(KEYINPUT56), .B(G101), .Z(n1262) );
XOR2_X1 U1010 ( .A(n1106), .B(KEYINPUT54), .Z(n1261) );
NAND3_X1 U1011 ( .A1(n1187), .A2(n1047), .A3(G210), .ZN(n1106) );
INV_X1 U1012 ( .A(G953), .ZN(n1047) );
INV_X1 U1013 ( .A(G237), .ZN(n1187) );
XNOR2_X1 U1014 ( .A(n1263), .B(n1264), .ZN(n1104) );
XOR2_X1 U1015 ( .A(KEYINPUT9), .B(G113), .Z(n1264) );
XOR2_X1 U1016 ( .A(n1265), .B(n1266), .Z(n1263) );
INV_X1 U1017 ( .A(n1173), .ZN(n1266) );
XOR2_X1 U1018 ( .A(n1267), .B(n1268), .Z(n1173) );
XOR2_X1 U1019 ( .A(KEYINPUT59), .B(KEYINPUT23), .Z(n1268) );
XOR2_X1 U1020 ( .A(n1054), .B(n1056), .Z(n1267) );
XOR2_X1 U1021 ( .A(G131), .B(n1269), .Z(n1056) );
XOR2_X1 U1022 ( .A(G137), .B(G134), .Z(n1269) );
XNOR2_X1 U1023 ( .A(G146), .B(n1235), .ZN(n1054) );
XOR2_X1 U1024 ( .A(n1152), .B(n1142), .Z(n1235) );
INV_X1 U1025 ( .A(G143), .ZN(n1142) );
INV_X1 U1026 ( .A(G128), .ZN(n1152) );
NAND2_X1 U1027 ( .A1(KEYINPUT21), .A2(n1203), .ZN(n1265) );
XOR2_X1 U1028 ( .A(G116), .B(G119), .Z(n1203) );
endmodule


