//Key = 1000100101010011001010100100010100000111100111111110010011011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416;

XOR2_X1 U764 ( .A(G107), .B(n1063), .Z(G9) );
NOR2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
AND2_X1 U766 ( .A1(KEYINPUT38), .A2(n1066), .ZN(n1065) );
NOR2_X1 U767 ( .A1(KEYINPUT37), .A2(n1066), .ZN(n1064) );
NAND4_X1 U768 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(G75) );
NAND4_X1 U769 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1069) );
NOR3_X1 U770 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1074) );
XOR2_X1 U771 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U772 ( .A1(n1080), .A2(KEYINPUT27), .ZN(n1079) );
NOR2_X1 U773 ( .A1(n1081), .A2(n1082), .ZN(n1076) );
AND2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NAND3_X1 U775 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1075) );
NOR3_X1 U776 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1073) );
NOR3_X1 U777 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
INV_X1 U778 ( .A(KEYINPUT49), .ZN(n1091) );
NOR2_X1 U779 ( .A1(KEYINPUT49), .A2(G472), .ZN(n1089) );
XNOR2_X1 U780 ( .A(KEYINPUT54), .B(n1094), .ZN(n1088) );
XOR2_X1 U781 ( .A(n1095), .B(n1096), .Z(n1071) );
NOR2_X1 U782 ( .A1(KEYINPUT8), .A2(n1097), .ZN(n1096) );
NAND2_X1 U783 ( .A1(n1098), .A2(n1099), .ZN(n1068) );
NAND2_X1 U784 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND3_X1 U785 ( .A1(n1102), .A2(n1103), .A3(n1072), .ZN(n1101) );
NAND2_X1 U786 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U787 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U788 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U789 ( .A1(n1110), .A2(n1111), .ZN(n1104) );
NAND2_X1 U790 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
OR2_X1 U791 ( .A1(n1086), .A2(n1114), .ZN(n1113) );
NAND3_X1 U792 ( .A1(n1110), .A2(n1115), .A3(n1106), .ZN(n1100) );
NAND3_X1 U793 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
NAND2_X1 U794 ( .A1(n1102), .A2(n1119), .ZN(n1118) );
NAND2_X1 U795 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U796 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U797 ( .A1(n1072), .A2(n1124), .ZN(n1117) );
NAND2_X1 U798 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U799 ( .A1(KEYINPUT57), .A2(n1127), .ZN(n1126) );
NAND3_X1 U800 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1116) );
INV_X1 U801 ( .A(KEYINPUT57), .ZN(n1128) );
INV_X1 U802 ( .A(n1130), .ZN(n1098) );
NAND2_X1 U803 ( .A1(n1131), .A2(n1132), .ZN(G72) );
NAND2_X1 U804 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U805 ( .A(KEYINPUT53), .B(n1135), .Z(n1131) );
NOR2_X1 U806 ( .A1(n1133), .A2(n1134), .ZN(n1135) );
NAND2_X1 U807 ( .A1(G953), .A2(n1136), .ZN(n1134) );
NAND2_X1 U808 ( .A1(G900), .A2(G227), .ZN(n1136) );
NAND2_X1 U809 ( .A1(n1137), .A2(n1138), .ZN(n1133) );
NAND2_X1 U810 ( .A1(n1139), .A2(n1070), .ZN(n1138) );
XOR2_X1 U811 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND3_X1 U812 ( .A1(G900), .A2(n1141), .A3(G953), .ZN(n1137) );
XNOR2_X1 U813 ( .A(n1142), .B(n1143), .ZN(n1141) );
XOR2_X1 U814 ( .A(n1144), .B(n1145), .Z(n1142) );
NOR2_X1 U815 ( .A1(KEYINPUT52), .A2(n1146), .ZN(n1145) );
NAND2_X1 U816 ( .A1(n1147), .A2(n1148), .ZN(n1144) );
NAND2_X1 U817 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NAND2_X1 U818 ( .A1(KEYINPUT61), .A2(n1151), .ZN(n1150) );
NAND2_X1 U819 ( .A1(KEYINPUT45), .A2(n1152), .ZN(n1151) );
INV_X1 U820 ( .A(n1153), .ZN(n1149) );
NAND2_X1 U821 ( .A1(G131), .A2(n1154), .ZN(n1147) );
NAND2_X1 U822 ( .A1(KEYINPUT45), .A2(n1155), .ZN(n1154) );
NAND2_X1 U823 ( .A1(KEYINPUT61), .A2(n1153), .ZN(n1155) );
XOR2_X1 U824 ( .A(n1156), .B(n1157), .Z(G69) );
NOR2_X1 U825 ( .A1(n1158), .A2(n1070), .ZN(n1157) );
NOR2_X1 U826 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NAND2_X1 U827 ( .A1(n1161), .A2(n1162), .ZN(n1156) );
NAND2_X1 U828 ( .A1(n1163), .A2(n1070), .ZN(n1162) );
XOR2_X1 U829 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND3_X1 U830 ( .A1(n1164), .A2(G898), .A3(G953), .ZN(n1161) );
XNOR2_X1 U831 ( .A(n1166), .B(n1167), .ZN(n1164) );
XOR2_X1 U832 ( .A(n1168), .B(KEYINPUT28), .Z(n1166) );
NOR2_X1 U833 ( .A1(n1169), .A2(n1170), .ZN(G66) );
XOR2_X1 U834 ( .A(n1171), .B(n1172), .Z(n1170) );
NAND2_X1 U835 ( .A1(n1173), .A2(n1080), .ZN(n1172) );
NOR2_X1 U836 ( .A1(n1169), .A2(n1174), .ZN(G63) );
XOR2_X1 U837 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U838 ( .A1(n1173), .A2(G478), .ZN(n1175) );
NOR2_X1 U839 ( .A1(n1169), .A2(n1177), .ZN(G60) );
XOR2_X1 U840 ( .A(n1178), .B(n1084), .Z(n1177) );
NAND2_X1 U841 ( .A1(n1173), .A2(G475), .ZN(n1178) );
XOR2_X1 U842 ( .A(n1179), .B(n1180), .Z(G6) );
NOR2_X1 U843 ( .A1(n1169), .A2(n1181), .ZN(G57) );
XOR2_X1 U844 ( .A(n1182), .B(n1183), .Z(n1181) );
NAND2_X1 U845 ( .A1(KEYINPUT11), .A2(n1184), .ZN(n1182) );
NAND2_X1 U846 ( .A1(n1173), .A2(G472), .ZN(n1184) );
NOR2_X1 U847 ( .A1(n1169), .A2(n1185), .ZN(G54) );
XOR2_X1 U848 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U849 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U850 ( .A(n1190), .B(n1191), .Z(n1189) );
XOR2_X1 U851 ( .A(n1192), .B(n1193), .Z(n1186) );
XNOR2_X1 U852 ( .A(n1194), .B(KEYINPUT46), .ZN(n1193) );
NAND2_X1 U853 ( .A1(KEYINPUT0), .A2(n1195), .ZN(n1194) );
NAND2_X1 U854 ( .A1(n1173), .A2(G469), .ZN(n1195) );
NAND2_X1 U855 ( .A1(KEYINPUT15), .A2(n1196), .ZN(n1192) );
INV_X1 U856 ( .A(n1197), .ZN(n1196) );
NOR2_X1 U857 ( .A1(n1169), .A2(n1198), .ZN(G51) );
XOR2_X1 U858 ( .A(n1199), .B(n1200), .Z(n1198) );
XNOR2_X1 U859 ( .A(n1201), .B(n1202), .ZN(n1200) );
NAND2_X1 U860 ( .A1(n1203), .A2(n1204), .ZN(n1201) );
NAND2_X1 U861 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XOR2_X1 U862 ( .A(n1207), .B(KEYINPUT26), .Z(n1205) );
NAND2_X1 U863 ( .A1(n1208), .A2(G125), .ZN(n1203) );
XOR2_X1 U864 ( .A(KEYINPUT21), .B(n1209), .Z(n1208) );
INV_X1 U865 ( .A(n1207), .ZN(n1209) );
XOR2_X1 U866 ( .A(n1210), .B(n1211), .Z(n1207) );
NAND2_X1 U867 ( .A1(n1173), .A2(n1212), .ZN(n1210) );
NOR2_X1 U868 ( .A1(n1083), .A2(n1067), .ZN(n1173) );
NOR2_X1 U869 ( .A1(n1165), .A2(n1140), .ZN(n1067) );
NAND4_X1 U870 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1140) );
AND4_X1 U871 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1216) );
NAND2_X1 U872 ( .A1(n1221), .A2(n1222), .ZN(n1215) );
INV_X1 U873 ( .A(KEYINPUT58), .ZN(n1222) );
NAND2_X1 U874 ( .A1(n1106), .A2(n1223), .ZN(n1213) );
NAND2_X1 U875 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NAND4_X1 U876 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1225) );
NAND2_X1 U877 ( .A1(n1230), .A2(n1120), .ZN(n1229) );
NAND2_X1 U878 ( .A1(KEYINPUT10), .A2(n1231), .ZN(n1230) );
NAND3_X1 U879 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1228) );
OR2_X1 U880 ( .A1(n1109), .A2(KEYINPUT10), .ZN(n1233) );
NAND2_X1 U881 ( .A1(KEYINPUT58), .A2(n1108), .ZN(n1232) );
NAND2_X1 U882 ( .A1(n1235), .A2(n1236), .ZN(n1165) );
NOR4_X1 U883 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1236) );
INV_X1 U884 ( .A(n1241), .ZN(n1240) );
INV_X1 U885 ( .A(n1066), .ZN(n1239) );
NAND3_X1 U886 ( .A1(n1102), .A2(n1242), .A3(n1243), .ZN(n1066) );
NOR4_X1 U887 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1247), .ZN(n1235) );
AND2_X1 U888 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
AND3_X1 U889 ( .A1(n1127), .A2(n1110), .A3(n1242), .ZN(n1246) );
INV_X1 U890 ( .A(n1180), .ZN(n1245) );
NAND3_X1 U891 ( .A1(n1102), .A2(n1242), .A3(n1231), .ZN(n1180) );
INV_X1 U892 ( .A(n1250), .ZN(n1244) );
XNOR2_X1 U893 ( .A(n1251), .B(KEYINPUT19), .ZN(n1199) );
NOR2_X1 U894 ( .A1(n1070), .A2(G952), .ZN(n1169) );
XOR2_X1 U895 ( .A(n1252), .B(n1214), .Z(G48) );
NAND3_X1 U896 ( .A1(n1231), .A2(n1248), .A3(n1253), .ZN(n1214) );
XOR2_X1 U897 ( .A(n1219), .B(n1254), .Z(G45) );
XOR2_X1 U898 ( .A(n1255), .B(KEYINPUT63), .Z(n1254) );
NAND4_X1 U899 ( .A1(n1234), .A2(n1248), .A3(n1226), .A4(n1256), .ZN(n1219) );
NOR3_X1 U900 ( .A1(n1094), .A2(n1257), .A3(n1258), .ZN(n1256) );
XOR2_X1 U901 ( .A(G140), .B(n1259), .Z(G42) );
NOR2_X1 U902 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XOR2_X1 U903 ( .A(n1224), .B(KEYINPUT34), .Z(n1260) );
NAND4_X1 U904 ( .A1(n1127), .A2(n1231), .A3(n1234), .A4(n1227), .ZN(n1224) );
INV_X1 U905 ( .A(n1109), .ZN(n1231) );
XNOR2_X1 U906 ( .A(G137), .B(n1218), .ZN(G39) );
NAND3_X1 U907 ( .A1(n1106), .A2(n1110), .A3(n1253), .ZN(n1218) );
XNOR2_X1 U908 ( .A(n1221), .B(n1262), .ZN(G36) );
XOR2_X1 U909 ( .A(n1263), .B(KEYINPUT1), .Z(n1262) );
NOR3_X1 U910 ( .A1(n1108), .A2(n1258), .A3(n1264), .ZN(n1221) );
XOR2_X1 U911 ( .A(G131), .B(n1265), .Z(G33) );
NOR3_X1 U912 ( .A1(n1264), .A2(n1266), .A3(n1109), .ZN(n1265) );
XOR2_X1 U913 ( .A(n1227), .B(KEYINPUT31), .Z(n1266) );
NAND3_X1 U914 ( .A1(n1226), .A2(n1234), .A3(n1106), .ZN(n1264) );
INV_X1 U915 ( .A(n1261), .ZN(n1106) );
NAND2_X1 U916 ( .A1(n1267), .A2(n1086), .ZN(n1261) );
INV_X1 U917 ( .A(n1114), .ZN(n1267) );
XOR2_X1 U918 ( .A(G128), .B(n1268), .Z(G30) );
NOR2_X1 U919 ( .A1(KEYINPUT24), .A2(n1220), .ZN(n1268) );
NAND3_X1 U920 ( .A1(n1243), .A2(n1248), .A3(n1253), .ZN(n1220) );
NOR4_X1 U921 ( .A1(n1120), .A2(n1269), .A3(n1258), .A4(n1270), .ZN(n1253) );
INV_X1 U922 ( .A(n1227), .ZN(n1258) );
XOR2_X1 U923 ( .A(n1238), .B(n1271), .Z(G3) );
NOR2_X1 U924 ( .A1(KEYINPUT51), .A2(n1272), .ZN(n1271) );
AND3_X1 U925 ( .A1(n1242), .A2(n1110), .A3(n1226), .ZN(n1238) );
NOR3_X1 U926 ( .A1(n1112), .A2(n1273), .A3(n1120), .ZN(n1242) );
INV_X1 U927 ( .A(n1234), .ZN(n1120) );
XOR2_X1 U928 ( .A(n1206), .B(n1217), .Z(G27) );
NAND3_X1 U929 ( .A1(n1274), .A2(n1227), .A3(n1127), .ZN(n1217) );
NOR2_X1 U930 ( .A1(n1275), .A2(n1269), .ZN(n1127) );
NAND2_X1 U931 ( .A1(n1130), .A2(n1276), .ZN(n1227) );
NAND4_X1 U932 ( .A1(G953), .A2(G902), .A3(n1277), .A4(n1278), .ZN(n1276) );
INV_X1 U933 ( .A(G900), .ZN(n1278) );
INV_X1 U934 ( .A(G125), .ZN(n1206) );
XOR2_X1 U935 ( .A(n1279), .B(n1250), .Z(G24) );
NAND4_X1 U936 ( .A1(n1102), .A2(n1248), .A3(n1072), .A4(n1280), .ZN(n1250) );
NOR3_X1 U937 ( .A1(n1094), .A2(n1257), .A3(n1273), .ZN(n1280) );
NOR2_X1 U938 ( .A1(n1275), .A2(n1281), .ZN(n1102) );
XOR2_X1 U939 ( .A(n1282), .B(n1241), .Z(G21) );
NAND4_X1 U940 ( .A1(n1283), .A2(n1072), .A3(n1248), .A4(n1275), .ZN(n1241) );
INV_X1 U941 ( .A(n1129), .ZN(n1072) );
NAND2_X1 U942 ( .A1(n1284), .A2(n1285), .ZN(G18) );
OR2_X1 U943 ( .A1(n1286), .A2(G116), .ZN(n1285) );
XOR2_X1 U944 ( .A(n1287), .B(KEYINPUT6), .Z(n1284) );
NAND2_X1 U945 ( .A1(G116), .A2(n1286), .ZN(n1287) );
NAND2_X1 U946 ( .A1(n1248), .A2(n1288), .ZN(n1286) );
XOR2_X1 U947 ( .A(KEYINPUT17), .B(n1249), .Z(n1288) );
NOR4_X1 U948 ( .A1(n1125), .A2(n1129), .A3(n1108), .A4(n1273), .ZN(n1249) );
INV_X1 U949 ( .A(n1289), .ZN(n1273) );
INV_X1 U950 ( .A(n1112), .ZN(n1248) );
XOR2_X1 U951 ( .A(n1290), .B(n1237), .Z(G15) );
AND3_X1 U952 ( .A1(n1274), .A2(n1289), .A3(n1226), .ZN(n1237) );
INV_X1 U953 ( .A(n1125), .ZN(n1226) );
NAND2_X1 U954 ( .A1(n1269), .A2(n1275), .ZN(n1125) );
NOR3_X1 U955 ( .A1(n1129), .A2(n1112), .A3(n1109), .ZN(n1274) );
NAND2_X1 U956 ( .A1(n1291), .A2(n1292), .ZN(n1109) );
XNOR2_X1 U957 ( .A(KEYINPUT22), .B(n1094), .ZN(n1291) );
NAND2_X1 U958 ( .A1(n1123), .A2(n1293), .ZN(n1129) );
NAND2_X1 U959 ( .A1(KEYINPUT62), .A2(n1294), .ZN(n1290) );
XOR2_X1 U960 ( .A(n1295), .B(n1296), .Z(G12) );
NAND4_X1 U961 ( .A1(n1297), .A2(n1283), .A3(n1270), .A4(n1298), .ZN(n1296) );
XOR2_X1 U962 ( .A(KEYINPUT42), .B(n1234), .Z(n1298) );
NOR2_X1 U963 ( .A1(n1123), .A2(n1122), .ZN(n1234) );
INV_X1 U964 ( .A(n1293), .ZN(n1122) );
NAND2_X1 U965 ( .A1(G221), .A2(n1299), .ZN(n1293) );
XOR2_X1 U966 ( .A(n1300), .B(G469), .Z(n1123) );
NAND2_X1 U967 ( .A1(n1301), .A2(n1083), .ZN(n1300) );
XOR2_X1 U968 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U969 ( .A(n1304), .B(KEYINPUT13), .ZN(n1303) );
NAND2_X1 U970 ( .A1(KEYINPUT7), .A2(n1190), .ZN(n1304) );
XOR2_X1 U971 ( .A(n1305), .B(KEYINPUT16), .Z(n1190) );
INV_X1 U972 ( .A(G140), .ZN(n1305) );
XOR2_X1 U973 ( .A(n1306), .B(n1191), .Z(n1302) );
XOR2_X1 U974 ( .A(G110), .B(n1307), .Z(n1191) );
AND2_X1 U975 ( .A1(n1070), .A2(G227), .ZN(n1307) );
NAND2_X1 U976 ( .A1(n1308), .A2(n1309), .ZN(n1306) );
NAND2_X1 U977 ( .A1(n1197), .A2(n1188), .ZN(n1309) );
XOR2_X1 U978 ( .A(KEYINPUT29), .B(n1310), .Z(n1308) );
NOR2_X1 U979 ( .A1(n1197), .A2(n1188), .ZN(n1310) );
XOR2_X1 U980 ( .A(n1311), .B(n1312), .Z(n1188) );
XOR2_X1 U981 ( .A(G107), .B(G104), .Z(n1312) );
XOR2_X1 U982 ( .A(n1143), .B(G101), .Z(n1311) );
NAND2_X1 U983 ( .A1(n1313), .A2(n1314), .ZN(n1143) );
NAND2_X1 U984 ( .A1(n1315), .A2(n1252), .ZN(n1314) );
XOR2_X1 U985 ( .A(KEYINPUT56), .B(n1316), .Z(n1315) );
NAND2_X1 U986 ( .A1(n1316), .A2(G146), .ZN(n1313) );
XOR2_X1 U987 ( .A(n1317), .B(KEYINPUT33), .Z(n1197) );
INV_X1 U988 ( .A(n1275), .ZN(n1270) );
NAND2_X1 U989 ( .A1(n1087), .A2(n1318), .ZN(n1275) );
OR2_X1 U990 ( .A1(n1093), .A2(n1092), .ZN(n1318) );
NAND2_X1 U991 ( .A1(n1092), .A2(n1093), .ZN(n1087) );
INV_X1 U992 ( .A(G472), .ZN(n1093) );
NOR2_X1 U993 ( .A1(n1183), .A2(G902), .ZN(n1092) );
XOR2_X1 U994 ( .A(n1319), .B(n1320), .Z(n1183) );
XOR2_X1 U995 ( .A(n1211), .B(n1321), .Z(n1320) );
XOR2_X1 U996 ( .A(G101), .B(n1322), .Z(n1321) );
NOR3_X1 U997 ( .A1(n1323), .A2(G953), .A3(G237), .ZN(n1322) );
INV_X1 U998 ( .A(G210), .ZN(n1323) );
INV_X1 U999 ( .A(n1324), .ZN(n1211) );
XOR2_X1 U1000 ( .A(n1325), .B(n1326), .Z(n1319) );
INV_X1 U1001 ( .A(n1317), .ZN(n1326) );
XOR2_X1 U1002 ( .A(n1152), .B(n1327), .Z(n1317) );
NOR2_X1 U1003 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NOR3_X1 U1004 ( .A1(KEYINPUT39), .A2(G137), .A3(n1263), .ZN(n1329) );
AND2_X1 U1005 ( .A1(n1153), .A2(KEYINPUT39), .ZN(n1328) );
XOR2_X1 U1006 ( .A(n1263), .B(G137), .Z(n1153) );
INV_X1 U1007 ( .A(G131), .ZN(n1152) );
NAND2_X1 U1008 ( .A1(n1330), .A2(n1331), .ZN(n1325) );
OR2_X1 U1009 ( .A1(n1332), .A2(G116), .ZN(n1331) );
NAND2_X1 U1010 ( .A1(n1333), .A2(G116), .ZN(n1330) );
XOR2_X1 U1011 ( .A(KEYINPUT41), .B(n1332), .Z(n1333) );
AND3_X1 U1012 ( .A1(n1281), .A2(n1289), .A3(n1110), .ZN(n1283) );
NAND2_X1 U1013 ( .A1(n1334), .A2(n1335), .ZN(n1110) );
OR2_X1 U1014 ( .A1(n1108), .A2(KEYINPUT22), .ZN(n1335) );
INV_X1 U1015 ( .A(n1243), .ZN(n1108) );
NOR2_X1 U1016 ( .A1(n1292), .A2(n1094), .ZN(n1243) );
NAND3_X1 U1017 ( .A1(n1257), .A2(n1094), .A3(KEYINPUT22), .ZN(n1334) );
XOR2_X1 U1018 ( .A(n1336), .B(G478), .Z(n1094) );
NAND2_X1 U1019 ( .A1(n1176), .A2(n1083), .ZN(n1336) );
XNOR2_X1 U1020 ( .A(n1337), .B(n1338), .ZN(n1176) );
AND2_X1 U1021 ( .A1(n1339), .A2(G217), .ZN(n1338) );
XOR2_X1 U1022 ( .A(n1340), .B(n1341), .Z(n1337) );
NOR2_X1 U1023 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NOR2_X1 U1024 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
XOR2_X1 U1025 ( .A(n1346), .B(G107), .Z(n1345) );
OR2_X1 U1026 ( .A1(n1279), .A2(KEYINPUT30), .ZN(n1346) );
NOR2_X1 U1027 ( .A1(G116), .A2(n1347), .ZN(n1344) );
NOR3_X1 U1028 ( .A1(n1347), .A2(G116), .A3(n1348), .ZN(n1342) );
XOR2_X1 U1029 ( .A(n1349), .B(n1350), .Z(n1348) );
NOR2_X1 U1030 ( .A1(G122), .A2(KEYINPUT30), .ZN(n1350) );
INV_X1 U1031 ( .A(KEYINPUT44), .ZN(n1347) );
NAND2_X1 U1032 ( .A1(n1351), .A2(n1352), .ZN(n1340) );
NAND2_X1 U1033 ( .A1(n1353), .A2(n1263), .ZN(n1352) );
XOR2_X1 U1034 ( .A(KEYINPUT47), .B(n1354), .Z(n1351) );
NOR2_X1 U1035 ( .A1(n1353), .A2(n1263), .ZN(n1354) );
INV_X1 U1036 ( .A(G134), .ZN(n1263) );
XNOR2_X1 U1037 ( .A(KEYINPUT35), .B(n1316), .ZN(n1353) );
INV_X1 U1038 ( .A(n1292), .ZN(n1257) );
NAND2_X1 U1039 ( .A1(n1355), .A2(n1085), .ZN(n1292) );
NAND3_X1 U1040 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1085) );
NAND2_X1 U1041 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
NAND2_X1 U1042 ( .A1(n1084), .A2(n1083), .ZN(n1357) );
XNOR2_X1 U1043 ( .A(n1358), .B(n1359), .ZN(n1084) );
XOR2_X1 U1044 ( .A(n1360), .B(n1361), .Z(n1359) );
XOR2_X1 U1045 ( .A(G131), .B(n1362), .Z(n1361) );
NOR2_X1 U1046 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
XOR2_X1 U1047 ( .A(n1365), .B(KEYINPUT25), .Z(n1364) );
NAND2_X1 U1048 ( .A1(n1366), .A2(n1367), .ZN(n1365) );
XOR2_X1 U1049 ( .A(KEYINPUT48), .B(n1368), .Z(n1367) );
XOR2_X1 U1050 ( .A(KEYINPUT50), .B(G104), .Z(n1366) );
AND2_X1 U1051 ( .A1(n1368), .A2(G104), .ZN(n1363) );
XOR2_X1 U1052 ( .A(n1294), .B(n1279), .Z(n1368) );
NOR2_X1 U1053 ( .A1(KEYINPUT23), .A2(n1255), .ZN(n1360) );
INV_X1 U1054 ( .A(G143), .ZN(n1255) );
XOR2_X1 U1055 ( .A(n1369), .B(n1370), .Z(n1358) );
NOR3_X1 U1056 ( .A1(n1371), .A2(G953), .A3(G237), .ZN(n1370) );
INV_X1 U1057 ( .A(G214), .ZN(n1371) );
NAND2_X1 U1058 ( .A1(KEYINPUT59), .A2(n1372), .ZN(n1369) );
XOR2_X1 U1059 ( .A(n1082), .B(KEYINPUT9), .Z(n1356) );
INV_X1 U1060 ( .A(G475), .ZN(n1082) );
NAND2_X1 U1061 ( .A1(n1130), .A2(n1373), .ZN(n1289) );
NAND4_X1 U1062 ( .A1(G953), .A2(G902), .A3(n1277), .A4(n1160), .ZN(n1373) );
INV_X1 U1063 ( .A(G898), .ZN(n1160) );
NAND3_X1 U1064 ( .A1(n1277), .A2(n1070), .A3(G952), .ZN(n1130) );
NAND2_X1 U1065 ( .A1(G237), .A2(G234), .ZN(n1277) );
INV_X1 U1066 ( .A(n1269), .ZN(n1281) );
XOR2_X1 U1067 ( .A(n1078), .B(n1080), .Z(n1269) );
AND2_X1 U1068 ( .A1(G217), .A2(n1299), .ZN(n1080) );
NAND2_X1 U1069 ( .A1(G234), .A2(n1083), .ZN(n1299) );
NAND2_X1 U1070 ( .A1(n1374), .A2(n1171), .ZN(n1078) );
NAND3_X1 U1071 ( .A1(n1375), .A2(n1376), .A3(n1377), .ZN(n1171) );
NAND2_X1 U1072 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
NAND2_X1 U1073 ( .A1(n1380), .A2(n1381), .ZN(n1376) );
INV_X1 U1074 ( .A(KEYINPUT40), .ZN(n1381) );
NAND2_X1 U1075 ( .A1(n1382), .A2(n1383), .ZN(n1380) );
INV_X1 U1076 ( .A(n1378), .ZN(n1383) );
XNOR2_X1 U1077 ( .A(KEYINPUT36), .B(n1379), .ZN(n1382) );
NAND2_X1 U1078 ( .A1(KEYINPUT40), .A2(n1384), .ZN(n1375) );
NAND2_X1 U1079 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
OR3_X1 U1080 ( .A1(n1378), .A2(n1379), .A3(KEYINPUT36), .ZN(n1386) );
XOR2_X1 U1081 ( .A(n1387), .B(G137), .Z(n1378) );
NAND2_X1 U1082 ( .A1(G221), .A2(n1339), .ZN(n1387) );
AND2_X1 U1083 ( .A1(G234), .A2(n1070), .ZN(n1339) );
INV_X1 U1084 ( .A(G953), .ZN(n1070) );
NAND2_X1 U1085 ( .A1(KEYINPUT36), .A2(n1379), .ZN(n1385) );
XNOR2_X1 U1086 ( .A(n1372), .B(n1388), .ZN(n1379) );
XOR2_X1 U1087 ( .A(n1295), .B(n1389), .Z(n1388) );
NAND2_X1 U1088 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
NAND2_X1 U1089 ( .A1(n1392), .A2(n1282), .ZN(n1391) );
XOR2_X1 U1090 ( .A(n1393), .B(KEYINPUT55), .Z(n1390) );
OR2_X1 U1091 ( .A1(n1392), .A2(n1282), .ZN(n1393) );
INV_X1 U1092 ( .A(G119), .ZN(n1282) );
XNOR2_X1 U1093 ( .A(n1394), .B(KEYINPUT3), .ZN(n1392) );
INV_X1 U1094 ( .A(G128), .ZN(n1394) );
XOR2_X1 U1095 ( .A(n1395), .B(n1146), .Z(n1372) );
XOR2_X1 U1096 ( .A(G140), .B(G125), .Z(n1146) );
XOR2_X1 U1097 ( .A(n1252), .B(KEYINPUT4), .Z(n1395) );
XOR2_X1 U1098 ( .A(n1083), .B(KEYINPUT2), .Z(n1374) );
XOR2_X1 U1099 ( .A(n1112), .B(KEYINPUT18), .Z(n1297) );
NAND2_X1 U1100 ( .A1(n1114), .A2(n1086), .ZN(n1112) );
NAND2_X1 U1101 ( .A1(G214), .A2(n1396), .ZN(n1086) );
XNOR2_X1 U1102 ( .A(n1097), .B(n1212), .ZN(n1114) );
INV_X1 U1103 ( .A(n1095), .ZN(n1212) );
NAND2_X1 U1104 ( .A1(G210), .A2(n1396), .ZN(n1095) );
NAND2_X1 U1105 ( .A1(n1397), .A2(n1083), .ZN(n1396) );
XOR2_X1 U1106 ( .A(KEYINPUT43), .B(G237), .Z(n1397) );
NAND2_X1 U1107 ( .A1(n1398), .A2(n1083), .ZN(n1097) );
INV_X1 U1108 ( .A(G902), .ZN(n1083) );
XOR2_X1 U1109 ( .A(n1399), .B(n1400), .Z(n1398) );
XOR2_X1 U1110 ( .A(n1401), .B(n1324), .Z(n1400) );
XOR2_X1 U1111 ( .A(n1252), .B(n1316), .Z(n1324) );
XOR2_X1 U1112 ( .A(G128), .B(G143), .Z(n1316) );
INV_X1 U1113 ( .A(G146), .ZN(n1252) );
NAND2_X1 U1114 ( .A1(KEYINPUT20), .A2(n1202), .ZN(n1401) );
NAND3_X1 U1115 ( .A1(n1402), .A2(n1403), .A3(n1404), .ZN(n1202) );
NAND2_X1 U1116 ( .A1(n1405), .A2(n1406), .ZN(n1404) );
NAND2_X1 U1117 ( .A1(KEYINPUT60), .A2(n1407), .ZN(n1406) );
XOR2_X1 U1118 ( .A(KEYINPUT5), .B(n1408), .Z(n1407) );
NAND3_X1 U1119 ( .A1(KEYINPUT60), .A2(n1167), .A3(n1408), .ZN(n1403) );
INV_X1 U1120 ( .A(n1405), .ZN(n1167) );
XOR2_X1 U1121 ( .A(n1409), .B(n1410), .Z(n1405) );
XNOR2_X1 U1122 ( .A(n1332), .B(n1411), .ZN(n1410) );
NAND2_X1 U1123 ( .A1(n1412), .A2(n1413), .ZN(n1411) );
NAND2_X1 U1124 ( .A1(n1414), .A2(n1349), .ZN(n1413) );
INV_X1 U1125 ( .A(G107), .ZN(n1349) );
XOR2_X1 U1126 ( .A(n1179), .B(KEYINPUT12), .Z(n1414) );
INV_X1 U1127 ( .A(G104), .ZN(n1179) );
NAND2_X1 U1128 ( .A1(n1415), .A2(G107), .ZN(n1412) );
XOR2_X1 U1129 ( .A(KEYINPUT32), .B(G104), .Z(n1415) );
XNOR2_X1 U1130 ( .A(n1294), .B(G119), .ZN(n1332) );
INV_X1 U1131 ( .A(G113), .ZN(n1294) );
XOR2_X1 U1132 ( .A(n1272), .B(G116), .Z(n1409) );
INV_X1 U1133 ( .A(G101), .ZN(n1272) );
OR2_X1 U1134 ( .A1(n1408), .A2(KEYINPUT60), .ZN(n1402) );
INV_X1 U1135 ( .A(n1168), .ZN(n1408) );
XOR2_X1 U1136 ( .A(n1416), .B(G110), .Z(n1168) );
NAND2_X1 U1137 ( .A1(KEYINPUT14), .A2(n1279), .ZN(n1416) );
INV_X1 U1138 ( .A(G122), .ZN(n1279) );
XOR2_X1 U1139 ( .A(G125), .B(n1251), .Z(n1399) );
NOR2_X1 U1140 ( .A1(n1159), .A2(G953), .ZN(n1251) );
INV_X1 U1141 ( .A(G224), .ZN(n1159) );
INV_X1 U1142 ( .A(G110), .ZN(n1295) );
endmodule


