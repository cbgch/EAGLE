//Key = 1011000111000000110101100011010111011001011101111000011011000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352;

XNOR2_X1 U742 ( .A(G107), .B(n1026), .ZN(G9) );
NAND3_X1 U743 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
XNOR2_X1 U744 ( .A(KEYINPUT14), .B(n1030), .ZN(n1028) );
NOR2_X1 U745 ( .A1(n1031), .A2(n1032), .ZN(G75) );
NOR3_X1 U746 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1032) );
NAND3_X1 U747 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1033) );
NAND2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND3_X1 U750 ( .A1(n1027), .A2(n1043), .A3(n1044), .ZN(n1042) );
NAND2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NAND2_X1 U752 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U753 ( .A1(n1049), .A2(n1030), .ZN(n1048) );
NAND2_X1 U754 ( .A1(n1050), .A2(n1051), .ZN(n1045) );
NAND2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U756 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND3_X1 U757 ( .A1(n1047), .A2(n1056), .A3(n1050), .ZN(n1041) );
NAND2_X1 U758 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U759 ( .A1(n1044), .A2(n1059), .ZN(n1058) );
NAND2_X1 U760 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U761 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U762 ( .A1(n1027), .A2(n1064), .ZN(n1057) );
NAND2_X1 U763 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U764 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
INV_X1 U765 ( .A(n1069), .ZN(n1039) );
NOR3_X1 U766 ( .A1(n1070), .A2(G953), .A3(G952), .ZN(n1031) );
INV_X1 U767 ( .A(n1036), .ZN(n1070) );
NAND4_X1 U768 ( .A1(n1071), .A2(n1072), .A3(n1047), .A4(n1073), .ZN(n1036) );
NOR4_X1 U769 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1073) );
XOR2_X1 U770 ( .A(KEYINPUT34), .B(n1078), .Z(n1077) );
XNOR2_X1 U771 ( .A(n1079), .B(n1080), .ZN(n1076) );
XNOR2_X1 U772 ( .A(n1081), .B(KEYINPUT29), .ZN(n1080) );
NOR2_X1 U773 ( .A1(KEYINPUT22), .A2(n1082), .ZN(n1075) );
NOR2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U775 ( .A1(n1027), .A2(n1085), .ZN(n1074) );
INV_X1 U776 ( .A(KEYINPUT22), .ZN(n1085) );
NAND2_X1 U777 ( .A1(n1086), .A2(n1087), .ZN(G72) );
NAND2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U779 ( .A1(G953), .A2(n1090), .ZN(n1088) );
NAND2_X1 U780 ( .A1(G900), .A2(G227), .ZN(n1090) );
NAND2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1086) );
NAND2_X1 U782 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
OR2_X1 U783 ( .A1(n1037), .A2(G227), .ZN(n1094) );
INV_X1 U784 ( .A(n1089), .ZN(n1091) );
NAND2_X1 U785 ( .A1(n1095), .A2(n1096), .ZN(n1089) );
NAND2_X1 U786 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U787 ( .A(KEYINPUT0), .B(n1099), .Z(n1095) );
NOR3_X1 U788 ( .A1(n1100), .A2(G953), .A3(n1098), .ZN(n1099) );
XOR2_X1 U789 ( .A(KEYINPUT6), .B(n1097), .Z(n1100) );
AND2_X1 U790 ( .A1(n1101), .A2(n1093), .ZN(n1097) );
INV_X1 U791 ( .A(n1102), .ZN(n1093) );
XOR2_X1 U792 ( .A(n1103), .B(n1104), .Z(n1101) );
XOR2_X1 U793 ( .A(KEYINPUT30), .B(n1105), .Z(n1104) );
XNOR2_X1 U794 ( .A(n1106), .B(n1107), .ZN(n1103) );
XOR2_X1 U795 ( .A(n1108), .B(n1109), .Z(G69) );
XOR2_X1 U796 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR3_X1 U797 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
NOR3_X1 U798 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
INV_X1 U799 ( .A(n1118), .ZN(n1115) );
NOR2_X1 U800 ( .A1(n1119), .A2(n1118), .ZN(n1113) );
XNOR2_X1 U801 ( .A(n1120), .B(KEYINPUT53), .ZN(n1118) );
NOR2_X1 U802 ( .A1(n1116), .A2(n1117), .ZN(n1119) );
NAND2_X1 U803 ( .A1(n1121), .A2(n1122), .ZN(n1117) );
OR2_X1 U804 ( .A1(n1123), .A2(KEYINPUT19), .ZN(n1122) );
NAND3_X1 U805 ( .A1(n1124), .A2(n1123), .A3(KEYINPUT19), .ZN(n1121) );
NOR2_X1 U806 ( .A1(G898), .A2(n1125), .ZN(n1112) );
XNOR2_X1 U807 ( .A(G953), .B(KEYINPUT55), .ZN(n1125) );
NAND2_X1 U808 ( .A1(n1037), .A2(n1035), .ZN(n1110) );
NAND2_X1 U809 ( .A1(G953), .A2(n1126), .ZN(n1108) );
NAND2_X1 U810 ( .A1(G898), .A2(G224), .ZN(n1126) );
NOR2_X1 U811 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XNOR2_X1 U812 ( .A(n1129), .B(n1130), .ZN(n1128) );
NAND2_X1 U813 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
NOR2_X1 U814 ( .A1(n1127), .A2(n1133), .ZN(G63) );
XOR2_X1 U815 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U816 ( .A1(n1131), .A2(G478), .ZN(n1134) );
NOR2_X1 U817 ( .A1(n1127), .A2(n1136), .ZN(G60) );
NOR3_X1 U818 ( .A1(n1081), .A2(n1137), .A3(n1138), .ZN(n1136) );
AND3_X1 U819 ( .A1(n1139), .A2(G475), .A3(n1131), .ZN(n1138) );
NOR2_X1 U820 ( .A1(n1140), .A2(n1139), .ZN(n1137) );
AND2_X1 U821 ( .A1(n1141), .A2(G475), .ZN(n1140) );
XNOR2_X1 U822 ( .A(G104), .B(n1142), .ZN(G6) );
NAND2_X1 U823 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U824 ( .A(n1145), .B(KEYINPUT36), .Z(n1143) );
NOR2_X1 U825 ( .A1(n1127), .A2(n1146), .ZN(G57) );
XOR2_X1 U826 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U827 ( .A(n1149), .B(n1150), .ZN(n1148) );
XOR2_X1 U828 ( .A(n1151), .B(n1152), .Z(n1147) );
NAND3_X1 U829 ( .A1(n1153), .A2(n1141), .A3(G472), .ZN(n1151) );
XNOR2_X1 U830 ( .A(KEYINPUT28), .B(n1154), .ZN(n1153) );
NOR2_X1 U831 ( .A1(n1155), .A2(n1156), .ZN(G54) );
XOR2_X1 U832 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U833 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U834 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U835 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U836 ( .A(n1165), .B(KEYINPUT27), .Z(n1164) );
NOR2_X1 U837 ( .A1(n1166), .A2(n1165), .ZN(n1161) );
NAND3_X1 U838 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1165) );
NAND2_X1 U839 ( .A1(G140), .A2(n1170), .ZN(n1169) );
NAND3_X1 U840 ( .A1(n1171), .A2(n1172), .A3(KEYINPUT26), .ZN(n1168) );
INV_X1 U841 ( .A(n1170), .ZN(n1171) );
NAND2_X1 U842 ( .A1(KEYINPUT43), .A2(n1173), .ZN(n1170) );
OR2_X1 U843 ( .A1(n1173), .A2(KEYINPUT26), .ZN(n1167) );
INV_X1 U844 ( .A(n1163), .ZN(n1166) );
XOR2_X1 U845 ( .A(n1174), .B(n1175), .Z(n1157) );
NAND3_X1 U846 ( .A1(G469), .A2(n1141), .A3(n1176), .ZN(n1174) );
XNOR2_X1 U847 ( .A(G902), .B(KEYINPUT17), .ZN(n1176) );
INV_X1 U848 ( .A(n1177), .ZN(n1141) );
XNOR2_X1 U849 ( .A(n1127), .B(KEYINPUT56), .ZN(n1155) );
NOR2_X1 U850 ( .A1(n1127), .A2(n1178), .ZN(G51) );
XOR2_X1 U851 ( .A(n1179), .B(n1180), .Z(n1178) );
XNOR2_X1 U852 ( .A(n1181), .B(n1182), .ZN(n1180) );
NOR2_X1 U853 ( .A1(KEYINPUT40), .A2(n1183), .ZN(n1181) );
XNOR2_X1 U854 ( .A(n1184), .B(n1185), .ZN(n1183) );
NOR2_X1 U855 ( .A1(KEYINPUT23), .A2(n1186), .ZN(n1185) );
XNOR2_X1 U856 ( .A(KEYINPUT33), .B(n1187), .ZN(n1186) );
NAND2_X1 U857 ( .A1(n1131), .A2(n1188), .ZN(n1179) );
NOR2_X1 U858 ( .A1(n1154), .A2(n1177), .ZN(n1131) );
NOR2_X1 U859 ( .A1(n1035), .A2(n1189), .ZN(n1177) );
XNOR2_X1 U860 ( .A(KEYINPUT24), .B(n1098), .ZN(n1189) );
INV_X1 U861 ( .A(n1034), .ZN(n1098) );
NAND4_X1 U862 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1034) );
NOR4_X1 U863 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
NOR2_X1 U864 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XNOR2_X1 U865 ( .A(n1200), .B(KEYINPUT4), .ZN(n1198) );
NOR3_X1 U866 ( .A1(n1201), .A2(n1065), .A3(n1202), .ZN(n1196) );
INV_X1 U867 ( .A(n1203), .ZN(n1195) );
NOR2_X1 U868 ( .A1(n1204), .A2(n1205), .ZN(n1192) );
NAND4_X1 U869 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1035) );
AND4_X1 U870 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1209) );
NAND2_X1 U871 ( .A1(n1144), .A2(n1214), .ZN(n1208) );
NAND2_X1 U872 ( .A1(n1215), .A2(n1145), .ZN(n1214) );
NAND4_X1 U873 ( .A1(n1200), .A2(n1027), .A3(n1216), .A4(n1217), .ZN(n1145) );
XOR2_X1 U874 ( .A(n1218), .B(KEYINPUT15), .Z(n1215) );
NAND3_X1 U875 ( .A1(n1027), .A2(n1219), .A3(n1029), .ZN(n1206) );
NOR2_X1 U876 ( .A1(n1037), .A2(G952), .ZN(n1127) );
XOR2_X1 U877 ( .A(G146), .B(n1194), .Z(G48) );
AND3_X1 U878 ( .A1(n1200), .A2(n1144), .A3(n1220), .ZN(n1194) );
NAND2_X1 U879 ( .A1(n1221), .A2(n1222), .ZN(G45) );
NAND2_X1 U880 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XOR2_X1 U881 ( .A(n1225), .B(KEYINPUT38), .Z(n1221) );
OR2_X1 U882 ( .A1(n1224), .A2(n1223), .ZN(n1225) );
NOR3_X1 U883 ( .A1(n1202), .A2(n1226), .A3(n1201), .ZN(n1223) );
NAND4_X1 U884 ( .A1(n1227), .A2(n1216), .A3(n1228), .A4(n1229), .ZN(n1201) );
XNOR2_X1 U885 ( .A(KEYINPUT18), .B(n1144), .ZN(n1226) );
INV_X1 U886 ( .A(G143), .ZN(n1224) );
XNOR2_X1 U887 ( .A(G140), .B(n1191), .ZN(G42) );
NAND4_X1 U888 ( .A1(n1044), .A2(n1230), .A3(n1063), .A4(n1200), .ZN(n1191) );
XOR2_X1 U889 ( .A(G137), .B(n1205), .Z(G39) );
AND3_X1 U890 ( .A1(n1044), .A2(n1050), .A3(n1220), .ZN(n1205) );
XNOR2_X1 U891 ( .A(n1204), .B(n1231), .ZN(G36) );
NAND2_X1 U892 ( .A1(KEYINPUT48), .A2(G134), .ZN(n1231) );
NOR2_X1 U893 ( .A1(n1199), .A2(n1030), .ZN(n1204) );
INV_X1 U894 ( .A(n1219), .ZN(n1030) );
XOR2_X1 U895 ( .A(G131), .B(n1232), .Z(G33) );
NOR2_X1 U896 ( .A1(n1049), .A2(n1199), .ZN(n1232) );
NAND4_X1 U897 ( .A1(n1044), .A2(n1227), .A3(n1216), .A4(n1229), .ZN(n1199) );
NOR2_X1 U898 ( .A1(n1233), .A2(n1067), .ZN(n1044) );
NAND2_X1 U899 ( .A1(n1234), .A2(n1235), .ZN(G30) );
NAND2_X1 U900 ( .A1(n1236), .A2(n1203), .ZN(n1235) );
XOR2_X1 U901 ( .A(KEYINPUT2), .B(n1237), .Z(n1234) );
NOR2_X1 U902 ( .A1(n1236), .A2(n1203), .ZN(n1237) );
NAND3_X1 U903 ( .A1(n1219), .A2(n1144), .A3(n1220), .ZN(n1203) );
AND2_X1 U904 ( .A1(n1230), .A2(n1084), .ZN(n1220) );
AND3_X1 U905 ( .A1(n1216), .A2(n1229), .A3(n1062), .ZN(n1230) );
XNOR2_X1 U906 ( .A(n1238), .B(KEYINPUT59), .ZN(n1236) );
XNOR2_X1 U907 ( .A(G101), .B(n1211), .ZN(G3) );
NAND3_X1 U908 ( .A1(n1050), .A2(n1029), .A3(n1227), .ZN(n1211) );
XNOR2_X1 U909 ( .A(G125), .B(n1190), .ZN(G27) );
NAND4_X1 U910 ( .A1(n1144), .A2(n1229), .A3(n1063), .A4(n1239), .ZN(n1190) );
AND3_X1 U911 ( .A1(n1200), .A2(n1047), .A3(n1062), .ZN(n1239) );
INV_X1 U912 ( .A(n1240), .ZN(n1047) );
NAND2_X1 U913 ( .A1(n1069), .A2(n1241), .ZN(n1229) );
NAND3_X1 U914 ( .A1(G902), .A2(n1242), .A3(n1102), .ZN(n1241) );
NOR2_X1 U915 ( .A1(n1037), .A2(G900), .ZN(n1102) );
XOR2_X1 U916 ( .A(n1207), .B(n1243), .Z(G24) );
NOR2_X1 U917 ( .A1(G122), .A2(KEYINPUT25), .ZN(n1243) );
NAND4_X1 U918 ( .A1(n1244), .A2(n1245), .A3(n1027), .A4(n1228), .ZN(n1207) );
AND2_X1 U919 ( .A1(n1063), .A2(n1083), .ZN(n1027) );
XOR2_X1 U920 ( .A(n1246), .B(n1247), .Z(G21) );
NOR2_X1 U921 ( .A1(n1248), .A2(n1218), .ZN(n1247) );
NAND3_X1 U922 ( .A1(n1062), .A2(n1050), .A3(n1249), .ZN(n1218) );
NOR3_X1 U923 ( .A1(n1240), .A2(n1250), .A3(n1063), .ZN(n1249) );
XNOR2_X1 U924 ( .A(n1144), .B(KEYINPUT1), .ZN(n1248) );
NAND2_X1 U925 ( .A1(KEYINPUT57), .A2(n1251), .ZN(n1246) );
XNOR2_X1 U926 ( .A(G116), .B(n1213), .ZN(G18) );
NAND3_X1 U927 ( .A1(n1227), .A2(n1219), .A3(n1245), .ZN(n1213) );
NOR2_X1 U928 ( .A1(n1071), .A2(n1244), .ZN(n1219) );
XNOR2_X1 U929 ( .A(G113), .B(n1212), .ZN(G15) );
NAND3_X1 U930 ( .A1(n1245), .A2(n1227), .A3(n1200), .ZN(n1212) );
INV_X1 U931 ( .A(n1049), .ZN(n1200) );
NAND2_X1 U932 ( .A1(n1244), .A2(n1252), .ZN(n1049) );
INV_X1 U933 ( .A(n1202), .ZN(n1244) );
INV_X1 U934 ( .A(n1060), .ZN(n1227) );
NAND2_X1 U935 ( .A1(n1083), .A2(n1084), .ZN(n1060) );
NOR3_X1 U936 ( .A1(n1065), .A2(n1250), .A3(n1240), .ZN(n1245) );
NAND2_X1 U937 ( .A1(n1055), .A2(n1253), .ZN(n1240) );
XNOR2_X1 U938 ( .A(G110), .B(n1210), .ZN(G12) );
NAND4_X1 U939 ( .A1(n1062), .A2(n1050), .A3(n1063), .A4(n1029), .ZN(n1210) );
NOR3_X1 U940 ( .A1(n1052), .A2(n1250), .A3(n1065), .ZN(n1029) );
INV_X1 U941 ( .A(n1144), .ZN(n1065) );
NOR2_X1 U942 ( .A1(n1068), .A2(n1067), .ZN(n1144) );
INV_X1 U943 ( .A(n1072), .ZN(n1067) );
NAND2_X1 U944 ( .A1(G214), .A2(n1254), .ZN(n1072) );
INV_X1 U945 ( .A(n1233), .ZN(n1068) );
XOR2_X1 U946 ( .A(n1078), .B(KEYINPUT20), .Z(n1233) );
XNOR2_X1 U947 ( .A(n1255), .B(n1188), .ZN(n1078) );
AND2_X1 U948 ( .A1(G210), .A2(n1254), .ZN(n1188) );
NAND2_X1 U949 ( .A1(n1154), .A2(n1256), .ZN(n1254) );
NAND3_X1 U950 ( .A1(n1257), .A2(n1154), .A3(n1258), .ZN(n1255) );
XOR2_X1 U951 ( .A(n1259), .B(KEYINPUT51), .Z(n1258) );
NAND2_X1 U952 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XOR2_X1 U953 ( .A(n1262), .B(KEYINPUT37), .Z(n1261) );
XNOR2_X1 U954 ( .A(n1263), .B(KEYINPUT13), .ZN(n1260) );
INV_X1 U955 ( .A(n1182), .ZN(n1263) );
NAND2_X1 U956 ( .A1(n1264), .A2(n1265), .ZN(n1257) );
XNOR2_X1 U957 ( .A(KEYINPUT37), .B(n1262), .ZN(n1265) );
NAND3_X1 U958 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(n1262) );
OR2_X1 U959 ( .A1(n1184), .A2(n1269), .ZN(n1268) );
NAND3_X1 U960 ( .A1(n1269), .A2(n1184), .A3(KEYINPUT32), .ZN(n1267) );
XNOR2_X1 U961 ( .A(n1270), .B(n1238), .ZN(n1184) );
NOR2_X1 U962 ( .A1(KEYINPUT44), .A2(n1187), .ZN(n1269) );
NAND2_X1 U963 ( .A1(n1187), .A2(n1271), .ZN(n1266) );
INV_X1 U964 ( .A(KEYINPUT32), .ZN(n1271) );
NAND2_X1 U965 ( .A1(G224), .A2(n1037), .ZN(n1187) );
XNOR2_X1 U966 ( .A(KEYINPUT13), .B(n1182), .ZN(n1264) );
NAND3_X1 U967 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n1182) );
NAND2_X1 U968 ( .A1(n1275), .A2(n1124), .ZN(n1274) );
XNOR2_X1 U969 ( .A(n1120), .B(n1123), .ZN(n1275) );
OR3_X1 U970 ( .A1(n1276), .A2(n1124), .A3(n1120), .ZN(n1273) );
NAND2_X1 U971 ( .A1(n1116), .A2(n1120), .ZN(n1272) );
XOR2_X1 U972 ( .A(n1277), .B(n1278), .Z(n1120) );
XOR2_X1 U973 ( .A(KEYINPUT8), .B(G122), .Z(n1278) );
NAND2_X1 U974 ( .A1(KEYINPUT16), .A2(n1173), .ZN(n1277) );
INV_X1 U975 ( .A(G110), .ZN(n1173) );
NOR2_X1 U976 ( .A1(n1123), .A2(n1124), .ZN(n1116) );
XOR2_X1 U977 ( .A(n1279), .B(n1280), .Z(n1124) );
NOR2_X1 U978 ( .A1(KEYINPUT52), .A2(n1281), .ZN(n1280) );
INV_X1 U979 ( .A(n1276), .ZN(n1123) );
XOR2_X1 U980 ( .A(G113), .B(n1282), .Z(n1276) );
INV_X1 U981 ( .A(n1217), .ZN(n1250) );
NAND2_X1 U982 ( .A1(n1069), .A2(n1283), .ZN(n1217) );
NAND4_X1 U983 ( .A1(G953), .A2(G902), .A3(n1242), .A4(n1284), .ZN(n1283) );
INV_X1 U984 ( .A(G898), .ZN(n1284) );
NAND3_X1 U985 ( .A1(n1242), .A2(n1037), .A3(G952), .ZN(n1069) );
NAND2_X1 U986 ( .A1(G237), .A2(G234), .ZN(n1242) );
INV_X1 U987 ( .A(n1216), .ZN(n1052) );
NOR2_X1 U988 ( .A1(n1055), .A2(n1054), .ZN(n1216) );
INV_X1 U989 ( .A(n1253), .ZN(n1054) );
NAND2_X1 U990 ( .A1(G221), .A2(n1285), .ZN(n1253) );
XOR2_X1 U991 ( .A(n1286), .B(G469), .Z(n1055) );
NAND2_X1 U992 ( .A1(n1287), .A2(n1154), .ZN(n1286) );
XOR2_X1 U993 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U994 ( .A(n1290), .B(n1106), .Z(n1289) );
XNOR2_X1 U995 ( .A(n1291), .B(n1172), .ZN(n1106) );
NAND2_X1 U996 ( .A1(KEYINPUT63), .A2(n1292), .ZN(n1290) );
XNOR2_X1 U997 ( .A(n1293), .B(n1159), .ZN(n1292) );
XOR2_X1 U998 ( .A(n1294), .B(n1295), .Z(n1159) );
INV_X1 U999 ( .A(n1279), .ZN(n1295) );
XOR2_X1 U1000 ( .A(G101), .B(KEYINPUT54), .Z(n1279) );
XNOR2_X1 U1001 ( .A(n1105), .B(n1281), .ZN(n1294) );
XNOR2_X1 U1002 ( .A(G104), .B(n1296), .ZN(n1281) );
NOR2_X1 U1003 ( .A1(KEYINPUT58), .A2(n1238), .ZN(n1105) );
XOR2_X1 U1004 ( .A(n1297), .B(n1298), .Z(n1288) );
NOR2_X1 U1005 ( .A1(KEYINPUT5), .A2(n1163), .ZN(n1298) );
NAND2_X1 U1006 ( .A1(G227), .A2(n1037), .ZN(n1163) );
XNOR2_X1 U1007 ( .A(G110), .B(KEYINPUT49), .ZN(n1297) );
INV_X1 U1008 ( .A(n1084), .ZN(n1063) );
XNOR2_X1 U1009 ( .A(n1299), .B(G472), .ZN(n1084) );
NAND2_X1 U1010 ( .A1(n1300), .A2(n1154), .ZN(n1299) );
XNOR2_X1 U1011 ( .A(n1152), .B(n1301), .ZN(n1300) );
NOR3_X1 U1012 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1301) );
NOR2_X1 U1013 ( .A1(KEYINPUT35), .A2(n1150), .ZN(n1304) );
INV_X1 U1014 ( .A(n1305), .ZN(n1150) );
AND3_X1 U1015 ( .A1(KEYINPUT35), .A2(n1149), .A3(n1306), .ZN(n1303) );
NOR2_X1 U1016 ( .A1(n1306), .A2(n1149), .ZN(n1302) );
INV_X1 U1017 ( .A(G101), .ZN(n1149) );
NOR2_X1 U1018 ( .A1(KEYINPUT12), .A2(n1305), .ZN(n1306) );
NAND3_X1 U1019 ( .A1(n1256), .A2(n1037), .A3(G210), .ZN(n1305) );
XNOR2_X1 U1020 ( .A(n1307), .B(n1308), .ZN(n1152) );
XNOR2_X1 U1021 ( .A(n1238), .B(G113), .ZN(n1308) );
XNOR2_X1 U1022 ( .A(n1175), .B(n1309), .ZN(n1307) );
NOR2_X1 U1023 ( .A1(KEYINPUT11), .A2(n1282), .ZN(n1309) );
XOR2_X1 U1024 ( .A(n1251), .B(G116), .Z(n1282) );
INV_X1 U1025 ( .A(G119), .ZN(n1251) );
XOR2_X1 U1026 ( .A(n1291), .B(n1293), .Z(n1175) );
XNOR2_X1 U1027 ( .A(G131), .B(n1310), .ZN(n1291) );
XOR2_X1 U1028 ( .A(G137), .B(G134), .Z(n1310) );
AND2_X1 U1029 ( .A1(n1252), .A2(n1202), .ZN(n1050) );
XNOR2_X1 U1030 ( .A(n1311), .B(n1081), .ZN(n1202) );
NOR2_X1 U1031 ( .A1(n1139), .A2(G902), .ZN(n1081) );
XOR2_X1 U1032 ( .A(n1312), .B(n1313), .Z(n1139) );
XNOR2_X1 U1033 ( .A(n1107), .B(n1314), .ZN(n1313) );
XNOR2_X1 U1034 ( .A(n1315), .B(n1316), .ZN(n1314) );
NOR2_X1 U1035 ( .A1(G104), .A2(KEYINPUT10), .ZN(n1316) );
NAND4_X1 U1036 ( .A1(KEYINPUT46), .A2(G214), .A3(n1256), .A4(n1037), .ZN(n1315) );
INV_X1 U1037 ( .A(G237), .ZN(n1256) );
INV_X1 U1038 ( .A(n1270), .ZN(n1107) );
XNOR2_X1 U1039 ( .A(G125), .B(n1293), .ZN(n1270) );
XNOR2_X1 U1040 ( .A(G146), .B(G143), .ZN(n1293) );
XOR2_X1 U1041 ( .A(n1317), .B(n1318), .Z(n1312) );
XNOR2_X1 U1042 ( .A(KEYINPUT61), .B(n1172), .ZN(n1318) );
INV_X1 U1043 ( .A(G140), .ZN(n1172) );
XOR2_X1 U1044 ( .A(n1319), .B(G131), .Z(n1317) );
NAND2_X1 U1045 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NAND2_X1 U1046 ( .A1(G122), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1047 ( .A(KEYINPUT39), .B(n1323), .Z(n1320) );
NOR2_X1 U1048 ( .A1(G122), .A2(n1322), .ZN(n1323) );
INV_X1 U1049 ( .A(G113), .ZN(n1322) );
NAND2_X1 U1050 ( .A1(KEYINPUT47), .A2(n1079), .ZN(n1311) );
XOR2_X1 U1051 ( .A(G475), .B(KEYINPUT9), .Z(n1079) );
XNOR2_X1 U1052 ( .A(n1071), .B(KEYINPUT31), .ZN(n1252) );
INV_X1 U1053 ( .A(n1228), .ZN(n1071) );
XNOR2_X1 U1054 ( .A(n1324), .B(G478), .ZN(n1228) );
NAND2_X1 U1055 ( .A1(n1135), .A2(n1154), .ZN(n1324) );
XNOR2_X1 U1056 ( .A(n1325), .B(n1326), .ZN(n1135) );
AND3_X1 U1057 ( .A1(G217), .A2(n1037), .A3(G234), .ZN(n1326) );
XOR2_X1 U1058 ( .A(n1327), .B(n1328), .Z(n1325) );
NOR2_X1 U1059 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XOR2_X1 U1060 ( .A(KEYINPUT50), .B(n1331), .Z(n1330) );
NOR2_X1 U1061 ( .A1(G134), .A2(n1332), .ZN(n1331) );
AND2_X1 U1062 ( .A1(n1332), .A2(G134), .ZN(n1329) );
XNOR2_X1 U1063 ( .A(G143), .B(n1238), .ZN(n1332) );
NAND2_X1 U1064 ( .A1(n1333), .A2(n1334), .ZN(n1327) );
NAND2_X1 U1065 ( .A1(n1335), .A2(n1296), .ZN(n1334) );
XOR2_X1 U1066 ( .A(KEYINPUT3), .B(n1336), .Z(n1333) );
NOR2_X1 U1067 ( .A1(n1335), .A2(n1296), .ZN(n1336) );
INV_X1 U1068 ( .A(G107), .ZN(n1296) );
XNOR2_X1 U1069 ( .A(G116), .B(G122), .ZN(n1335) );
XOR2_X1 U1070 ( .A(n1083), .B(KEYINPUT41), .Z(n1062) );
XNOR2_X1 U1071 ( .A(n1132), .B(n1337), .ZN(n1083) );
NOR2_X1 U1072 ( .A1(G902), .A2(n1130), .ZN(n1337) );
XNOR2_X1 U1073 ( .A(n1338), .B(n1339), .ZN(n1130) );
NOR2_X1 U1074 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
XOR2_X1 U1075 ( .A(n1342), .B(KEYINPUT42), .Z(n1341) );
NAND2_X1 U1076 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
NOR2_X1 U1077 ( .A1(n1343), .A2(n1344), .ZN(n1340) );
XNOR2_X1 U1078 ( .A(n1345), .B(n1346), .ZN(n1344) );
NOR2_X1 U1079 ( .A1(KEYINPUT62), .A2(n1347), .ZN(n1346) );
XOR2_X1 U1080 ( .A(KEYINPUT45), .B(G146), .Z(n1347) );
XNOR2_X1 U1081 ( .A(G125), .B(G140), .ZN(n1345) );
XOR2_X1 U1082 ( .A(n1348), .B(n1349), .Z(n1343) );
XNOR2_X1 U1083 ( .A(KEYINPUT60), .B(n1238), .ZN(n1349) );
INV_X1 U1084 ( .A(G128), .ZN(n1238) );
XNOR2_X1 U1085 ( .A(G119), .B(G110), .ZN(n1348) );
NAND2_X1 U1086 ( .A1(n1350), .A2(KEYINPUT21), .ZN(n1338) );
XOR2_X1 U1087 ( .A(n1351), .B(G137), .Z(n1350) );
NAND2_X1 U1088 ( .A1(KEYINPUT7), .A2(n1352), .ZN(n1351) );
NAND3_X1 U1089 ( .A1(G234), .A2(n1037), .A3(G221), .ZN(n1352) );
INV_X1 U1090 ( .A(G953), .ZN(n1037) );
AND2_X1 U1091 ( .A1(G217), .A2(n1285), .ZN(n1132) );
NAND2_X1 U1092 ( .A1(G234), .A2(n1154), .ZN(n1285) );
INV_X1 U1093 ( .A(G902), .ZN(n1154) );
endmodule


