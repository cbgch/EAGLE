//Key = 1100001110010111010001001111010110100010010001001000111101010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361;

XNOR2_X1 U748 ( .A(G107), .B(n1035), .ZN(G9) );
NAND4_X1 U749 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
XOR2_X1 U750 ( .A(KEYINPUT3), .B(n1040), .Z(n1039) );
NOR2_X1 U751 ( .A1(n1041), .A2(n1042), .ZN(n1038) );
NOR2_X1 U752 ( .A1(n1043), .A2(n1044), .ZN(G75) );
NOR4_X1 U753 ( .A1(G953), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1044) );
NOR2_X1 U754 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U755 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR2_X1 U756 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U757 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U758 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U759 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U760 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U761 ( .A1(n1062), .A2(n1040), .ZN(n1060) );
NOR2_X1 U762 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U763 ( .A1(n1065), .A2(n1066), .ZN(n1058) );
NOR2_X1 U764 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR3_X1 U765 ( .A1(n1066), .A2(n1069), .A3(n1061), .ZN(n1054) );
NOR2_X1 U766 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR4_X1 U768 ( .A1(n1074), .A2(n1061), .A3(n1066), .A4(n1057), .ZN(n1050) );
NOR2_X1 U769 ( .A1(n1037), .A2(n1075), .ZN(n1074) );
NOR3_X1 U770 ( .A1(n1045), .A2(G953), .A3(G952), .ZN(n1043) );
AND4_X1 U771 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1045) );
NOR4_X1 U772 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1079) );
XOR2_X1 U773 ( .A(n1084), .B(KEYINPUT32), .Z(n1082) );
XOR2_X1 U774 ( .A(n1085), .B(n1086), .Z(n1081) );
NAND2_X1 U775 ( .A1(KEYINPUT1), .A2(n1087), .ZN(n1085) );
XOR2_X1 U776 ( .A(n1088), .B(KEYINPUT51), .Z(n1078) );
XOR2_X1 U777 ( .A(n1089), .B(n1090), .Z(G72) );
XOR2_X1 U778 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U779 ( .A1(G953), .A2(n1093), .ZN(n1092) );
NAND2_X1 U780 ( .A1(G900), .A2(G227), .ZN(n1093) );
NAND2_X1 U781 ( .A1(n1094), .A2(n1095), .ZN(n1091) );
NAND2_X1 U782 ( .A1(G953), .A2(n1096), .ZN(n1095) );
XOR2_X1 U783 ( .A(n1097), .B(n1098), .Z(n1094) );
XNOR2_X1 U784 ( .A(n1099), .B(n1100), .ZN(n1098) );
XNOR2_X1 U785 ( .A(G131), .B(n1101), .ZN(n1100) );
NOR2_X1 U786 ( .A1(KEYINPUT35), .A2(n1102), .ZN(n1101) );
XOR2_X1 U787 ( .A(G137), .B(n1103), .Z(n1097) );
XOR2_X1 U788 ( .A(KEYINPUT14), .B(G140), .Z(n1103) );
NOR2_X1 U789 ( .A1(n1104), .A2(G953), .ZN(n1089) );
XOR2_X1 U790 ( .A(n1105), .B(n1106), .Z(G69) );
NOR2_X1 U791 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XOR2_X1 U792 ( .A(n1109), .B(KEYINPUT56), .Z(n1108) );
AND2_X1 U793 ( .A1(G224), .A2(G898), .ZN(n1107) );
NOR2_X1 U794 ( .A1(KEYINPUT43), .A2(n1110), .ZN(n1105) );
XOR2_X1 U795 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U796 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U797 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U798 ( .A1(KEYINPUT10), .A2(n1117), .ZN(n1115) );
XNOR2_X1 U799 ( .A(n1118), .B(KEYINPUT55), .ZN(n1117) );
XNOR2_X1 U800 ( .A(n1119), .B(KEYINPUT48), .ZN(n1113) );
NAND2_X1 U801 ( .A1(n1120), .A2(n1121), .ZN(n1111) );
NAND2_X1 U802 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XOR2_X1 U803 ( .A(n1124), .B(KEYINPUT60), .Z(n1122) );
XOR2_X1 U804 ( .A(n1109), .B(KEYINPUT42), .Z(n1120) );
NOR2_X1 U805 ( .A1(n1125), .A2(n1126), .ZN(G66) );
XNOR2_X1 U806 ( .A(n1127), .B(n1128), .ZN(n1126) );
NOR2_X1 U807 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U808 ( .A1(n1125), .A2(n1131), .ZN(G63) );
NOR3_X1 U809 ( .A1(n1086), .A2(n1132), .A3(n1133), .ZN(n1131) );
AND3_X1 U810 ( .A1(n1134), .A2(G478), .A3(n1135), .ZN(n1133) );
NOR2_X1 U811 ( .A1(n1136), .A2(n1134), .ZN(n1132) );
AND2_X1 U812 ( .A1(n1047), .A2(G478), .ZN(n1136) );
NOR2_X1 U813 ( .A1(n1125), .A2(n1137), .ZN(G60) );
XOR2_X1 U814 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U815 ( .A1(n1140), .A2(KEYINPUT20), .ZN(n1139) );
INV_X1 U816 ( .A(n1141), .ZN(n1140) );
NAND2_X1 U817 ( .A1(n1135), .A2(G475), .ZN(n1138) );
XNOR2_X1 U818 ( .A(G104), .B(n1142), .ZN(G6) );
NOR2_X1 U819 ( .A1(n1125), .A2(n1143), .ZN(G57) );
XOR2_X1 U820 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U821 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U822 ( .A(n1148), .B(n1149), .Z(n1144) );
XNOR2_X1 U823 ( .A(n1150), .B(n1151), .ZN(n1149) );
NAND2_X1 U824 ( .A1(KEYINPUT63), .A2(n1152), .ZN(n1151) );
NAND3_X1 U825 ( .A1(n1135), .A2(G472), .A3(KEYINPUT29), .ZN(n1150) );
NOR3_X1 U826 ( .A1(n1125), .A2(n1153), .A3(n1154), .ZN(G54) );
NOR3_X1 U827 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1154) );
NOR2_X1 U828 ( .A1(KEYINPUT38), .A2(n1158), .ZN(n1157) );
NOR2_X1 U829 ( .A1(n1159), .A2(n1160), .ZN(n1153) );
NOR2_X1 U830 ( .A1(n1158), .A2(n1161), .ZN(n1160) );
INV_X1 U831 ( .A(KEYINPUT38), .ZN(n1161) );
XOR2_X1 U832 ( .A(n1156), .B(KEYINPUT2), .Z(n1158) );
AND2_X1 U833 ( .A1(n1162), .A2(n1163), .ZN(n1156) );
NAND2_X1 U834 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XOR2_X1 U835 ( .A(KEYINPUT59), .B(n1166), .Z(n1162) );
NOR2_X1 U836 ( .A1(n1164), .A2(n1165), .ZN(n1166) );
XOR2_X1 U837 ( .A(n1167), .B(n1168), .Z(n1165) );
NAND2_X1 U838 ( .A1(KEYINPUT31), .A2(n1169), .ZN(n1167) );
XOR2_X1 U839 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U840 ( .A(n1172), .B(n1173), .Z(n1164) );
NAND2_X1 U841 ( .A1(KEYINPUT27), .A2(n1174), .ZN(n1172) );
INV_X1 U842 ( .A(n1155), .ZN(n1159) );
NAND2_X1 U843 ( .A1(n1175), .A2(n1135), .ZN(n1155) );
INV_X1 U844 ( .A(n1130), .ZN(n1135) );
XNOR2_X1 U845 ( .A(G469), .B(KEYINPUT26), .ZN(n1175) );
NOR2_X1 U846 ( .A1(n1109), .A2(G952), .ZN(n1125) );
NOR2_X1 U847 ( .A1(n1176), .A2(n1177), .ZN(G51) );
XOR2_X1 U848 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U849 ( .A(KEYINPUT44), .B(n1180), .Z(n1179) );
NOR2_X1 U850 ( .A1(n1181), .A2(n1130), .ZN(n1180) );
NAND2_X1 U851 ( .A1(G902), .A2(n1047), .ZN(n1130) );
NAND3_X1 U852 ( .A1(n1123), .A2(n1124), .A3(n1104), .ZN(n1047) );
AND4_X1 U853 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1104) );
NOR4_X1 U854 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1185) );
INV_X1 U855 ( .A(n1190), .ZN(n1189) );
NOR4_X1 U856 ( .A1(n1042), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1188) );
XOR2_X1 U857 ( .A(KEYINPUT7), .B(n1040), .Z(n1193) );
NOR2_X1 U858 ( .A1(n1194), .A2(n1195), .ZN(n1184) );
NOR3_X1 U859 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1195) );
XOR2_X1 U860 ( .A(KEYINPUT52), .B(n1037), .Z(n1198) );
XOR2_X1 U861 ( .A(KEYINPUT45), .B(n1077), .Z(n1196) );
INV_X1 U862 ( .A(n1199), .ZN(n1194) );
AND4_X1 U863 ( .A1(n1200), .A2(n1201), .A3(n1142), .A4(n1202), .ZN(n1123) );
NOR3_X1 U864 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1202) );
NOR3_X1 U865 ( .A1(n1206), .A2(n1207), .A3(n1191), .ZN(n1205) );
NOR2_X1 U866 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
AND2_X1 U867 ( .A1(n1067), .A2(n1210), .ZN(n1209) );
NOR2_X1 U868 ( .A1(n1042), .A2(n1061), .ZN(n1208) );
INV_X1 U869 ( .A(n1211), .ZN(n1204) );
NOR3_X1 U870 ( .A1(n1212), .A2(n1042), .A3(n1053), .ZN(n1203) );
NAND3_X1 U871 ( .A1(n1213), .A2(n1214), .A3(n1068), .ZN(n1212) );
NAND2_X1 U872 ( .A1(KEYINPUT24), .A2(n1206), .ZN(n1214) );
NAND2_X1 U873 ( .A1(n1215), .A2(n1216), .ZN(n1213) );
INV_X1 U874 ( .A(KEYINPUT24), .ZN(n1216) );
NAND2_X1 U875 ( .A1(n1041), .A2(n1040), .ZN(n1215) );
INV_X1 U876 ( .A(n1217), .ZN(n1041) );
NAND4_X1 U877 ( .A1(n1218), .A2(n1075), .A3(n1036), .A4(n1219), .ZN(n1142) );
XOR2_X1 U878 ( .A(n1220), .B(n1221), .Z(n1178) );
NAND2_X1 U879 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
NOR2_X1 U880 ( .A1(n1109), .A2(n1224), .ZN(n1176) );
XOR2_X1 U881 ( .A(KEYINPUT37), .B(G952), .Z(n1224) );
XOR2_X1 U882 ( .A(n1225), .B(n1199), .Z(G48) );
NAND4_X1 U883 ( .A1(n1226), .A2(n1075), .A3(n1040), .A4(n1071), .ZN(n1199) );
XNOR2_X1 U884 ( .A(G143), .B(n1182), .ZN(G45) );
NAND4_X1 U885 ( .A1(n1227), .A2(n1040), .A3(n1228), .A4(n1083), .ZN(n1182) );
XNOR2_X1 U886 ( .A(G140), .B(n1183), .ZN(G42) );
NAND3_X1 U887 ( .A1(n1077), .A2(n1071), .A3(n1229), .ZN(n1183) );
XNOR2_X1 U888 ( .A(n1187), .B(n1230), .ZN(G39) );
XOR2_X1 U889 ( .A(KEYINPUT21), .B(G137), .Z(n1230) );
AND4_X1 U890 ( .A1(n1231), .A2(n1226), .A3(n1077), .A4(n1071), .ZN(n1187) );
XOR2_X1 U891 ( .A(n1232), .B(n1233), .Z(G36) );
NOR3_X1 U892 ( .A1(n1197), .A2(n1191), .A3(n1066), .ZN(n1233) );
INV_X1 U893 ( .A(n1077), .ZN(n1066) );
XOR2_X1 U894 ( .A(n1102), .B(KEYINPUT41), .Z(n1232) );
INV_X1 U895 ( .A(G134), .ZN(n1102) );
XOR2_X1 U896 ( .A(G131), .B(n1186), .Z(G33) );
AND3_X1 U897 ( .A1(n1227), .A2(n1077), .A3(n1075), .ZN(n1186) );
NOR2_X1 U898 ( .A1(n1064), .A2(n1234), .ZN(n1077) );
INV_X1 U899 ( .A(n1197), .ZN(n1227) );
NAND3_X1 U900 ( .A1(n1071), .A2(n1235), .A3(n1067), .ZN(n1197) );
XNOR2_X1 U901 ( .A(G128), .B(n1236), .ZN(G30) );
NAND4_X1 U902 ( .A1(n1226), .A2(n1037), .A3(n1040), .A4(n1219), .ZN(n1236) );
INV_X1 U903 ( .A(n1192), .ZN(n1226) );
NAND3_X1 U904 ( .A1(n1237), .A2(n1235), .A3(n1238), .ZN(n1192) );
XNOR2_X1 U905 ( .A(G101), .B(n1200), .ZN(G3) );
NAND4_X1 U906 ( .A1(n1218), .A2(n1231), .A3(n1067), .A4(n1219), .ZN(n1200) );
XOR2_X1 U907 ( .A(n1239), .B(G125), .Z(G27) );
NAND2_X1 U908 ( .A1(KEYINPUT57), .A2(n1190), .ZN(n1239) );
NAND3_X1 U909 ( .A1(n1229), .A2(n1040), .A3(n1210), .ZN(n1190) );
AND3_X1 U910 ( .A1(n1075), .A2(n1235), .A3(n1068), .ZN(n1229) );
NAND2_X1 U911 ( .A1(n1240), .A2(n1049), .ZN(n1235) );
XOR2_X1 U912 ( .A(n1241), .B(KEYINPUT5), .Z(n1240) );
NAND4_X1 U913 ( .A1(G902), .A2(G953), .A3(n1242), .A4(n1096), .ZN(n1241) );
INV_X1 U914 ( .A(G900), .ZN(n1096) );
NAND3_X1 U915 ( .A1(n1243), .A2(n1244), .A3(n1245), .ZN(G24) );
NAND2_X1 U916 ( .A1(G122), .A2(n1201), .ZN(n1245) );
NAND2_X1 U917 ( .A1(n1246), .A2(n1247), .ZN(n1244) );
INV_X1 U918 ( .A(KEYINPUT61), .ZN(n1247) );
NAND2_X1 U919 ( .A1(n1248), .A2(n1249), .ZN(n1246) );
XNOR2_X1 U920 ( .A(KEYINPUT49), .B(n1201), .ZN(n1248) );
NAND2_X1 U921 ( .A1(KEYINPUT61), .A2(n1250), .ZN(n1243) );
NAND2_X1 U922 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U923 ( .A1(KEYINPUT49), .A2(n1201), .ZN(n1252) );
OR3_X1 U924 ( .A1(G122), .A2(KEYINPUT49), .A3(n1201), .ZN(n1251) );
NAND4_X1 U925 ( .A1(n1218), .A2(n1210), .A3(n1253), .A4(n1036), .ZN(n1201) );
INV_X1 U926 ( .A(n1061), .ZN(n1036) );
NAND2_X1 U927 ( .A1(n1254), .A2(n1088), .ZN(n1061) );
AND2_X1 U928 ( .A1(n1083), .A2(n1228), .ZN(n1253) );
XOR2_X1 U929 ( .A(n1255), .B(n1124), .Z(G21) );
NAND3_X1 U930 ( .A1(n1218), .A2(n1210), .A3(n1256), .ZN(n1124) );
NOR3_X1 U931 ( .A1(n1053), .A2(n1254), .A3(n1088), .ZN(n1256) );
XNOR2_X1 U932 ( .A(G116), .B(n1257), .ZN(G18) );
NAND4_X1 U933 ( .A1(n1258), .A2(n1218), .A3(n1067), .A4(n1037), .ZN(n1257) );
INV_X1 U934 ( .A(n1191), .ZN(n1037) );
NAND2_X1 U935 ( .A1(n1228), .A2(n1259), .ZN(n1191) );
XOR2_X1 U936 ( .A(n1260), .B(KEYINPUT0), .Z(n1228) );
XOR2_X1 U937 ( .A(n1057), .B(KEYINPUT13), .Z(n1258) );
INV_X1 U938 ( .A(n1210), .ZN(n1057) );
XOR2_X1 U939 ( .A(n1261), .B(n1211), .Z(G15) );
NAND4_X1 U940 ( .A1(n1218), .A2(n1210), .A3(n1075), .A4(n1067), .ZN(n1211) );
NOR2_X1 U941 ( .A1(n1238), .A2(n1254), .ZN(n1067) );
INV_X1 U942 ( .A(n1088), .ZN(n1238) );
AND2_X1 U943 ( .A1(n1260), .A2(n1083), .ZN(n1075) );
INV_X1 U944 ( .A(n1259), .ZN(n1083) );
NOR2_X1 U945 ( .A1(n1072), .A2(n1080), .ZN(n1210) );
XOR2_X1 U946 ( .A(n1076), .B(KEYINPUT15), .Z(n1072) );
XOR2_X1 U947 ( .A(n1174), .B(n1262), .Z(G12) );
NAND4_X1 U948 ( .A1(n1218), .A2(n1231), .A3(n1263), .A4(n1219), .ZN(n1262) );
INV_X1 U949 ( .A(n1042), .ZN(n1219) );
XNOR2_X1 U950 ( .A(n1071), .B(KEYINPUT30), .ZN(n1042) );
NOR2_X1 U951 ( .A1(n1264), .A2(n1076), .ZN(n1071) );
XOR2_X1 U952 ( .A(n1265), .B(G469), .Z(n1076) );
NAND2_X1 U953 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XOR2_X1 U954 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U955 ( .A(G110), .B(n1173), .Z(n1269) );
XOR2_X1 U956 ( .A(G140), .B(n1270), .Z(n1173) );
AND2_X1 U957 ( .A1(n1109), .A2(G227), .ZN(n1270) );
XNOR2_X1 U958 ( .A(n1170), .B(n1271), .ZN(n1268) );
XNOR2_X1 U959 ( .A(n1272), .B(n1273), .ZN(n1170) );
NAND2_X1 U960 ( .A1(KEYINPUT17), .A2(n1274), .ZN(n1272) );
XOR2_X1 U961 ( .A(n1275), .B(KEYINPUT9), .Z(n1266) );
XOR2_X1 U962 ( .A(n1080), .B(KEYINPUT40), .Z(n1264) );
INV_X1 U963 ( .A(n1073), .ZN(n1080) );
NAND2_X1 U964 ( .A1(G221), .A2(n1276), .ZN(n1073) );
XOR2_X1 U965 ( .A(KEYINPUT4), .B(n1068), .Z(n1263) );
NOR2_X1 U966 ( .A1(n1237), .A2(n1088), .ZN(n1068) );
XNOR2_X1 U967 ( .A(n1277), .B(n1129), .ZN(n1088) );
NAND2_X1 U968 ( .A1(G217), .A2(n1276), .ZN(n1129) );
NAND2_X1 U969 ( .A1(G234), .A2(n1275), .ZN(n1276) );
NAND2_X1 U970 ( .A1(n1127), .A2(n1275), .ZN(n1277) );
XNOR2_X1 U971 ( .A(n1278), .B(n1279), .ZN(n1127) );
XOR2_X1 U972 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U973 ( .A(G110), .B(n1282), .Z(n1281) );
NOR2_X1 U974 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NOR3_X1 U975 ( .A1(n1285), .A2(G953), .A3(n1286), .ZN(n1280) );
XNOR2_X1 U976 ( .A(G234), .B(KEYINPUT22), .ZN(n1286) );
INV_X1 U977 ( .A(G221), .ZN(n1285) );
XOR2_X1 U978 ( .A(n1255), .B(n1287), .Z(n1278) );
XOR2_X1 U979 ( .A(G137), .B(G128), .Z(n1287) );
INV_X1 U980 ( .A(n1254), .ZN(n1237) );
XOR2_X1 U981 ( .A(n1084), .B(KEYINPUT19), .Z(n1254) );
XOR2_X1 U982 ( .A(n1288), .B(G472), .Z(n1084) );
NAND2_X1 U983 ( .A1(n1289), .A2(n1275), .ZN(n1288) );
XOR2_X1 U984 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U985 ( .A(n1273), .B(n1147), .Z(n1291) );
XNOR2_X1 U986 ( .A(n1261), .B(n1292), .ZN(n1147) );
NOR2_X1 U987 ( .A1(KEYINPUT23), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U988 ( .A(G116), .B(n1294), .ZN(n1293) );
NAND2_X1 U989 ( .A1(KEYINPUT34), .A2(n1255), .ZN(n1294) );
INV_X1 U990 ( .A(n1148), .ZN(n1273) );
XOR2_X1 U991 ( .A(n1295), .B(n1152), .Z(n1290) );
AND3_X1 U992 ( .A1(n1296), .A2(n1109), .A3(G210), .ZN(n1152) );
NAND2_X1 U993 ( .A1(KEYINPUT8), .A2(n1146), .ZN(n1295) );
XOR2_X1 U994 ( .A(n1271), .B(KEYINPUT6), .Z(n1146) );
XOR2_X1 U995 ( .A(n1171), .B(n1297), .Z(n1271) );
INV_X1 U996 ( .A(n1168), .ZN(n1297) );
XOR2_X1 U997 ( .A(n1298), .B(n1299), .Z(n1168) );
XOR2_X1 U998 ( .A(KEYINPUT53), .B(G134), .Z(n1299) );
XNOR2_X1 U999 ( .A(n1300), .B(n1301), .ZN(n1298) );
NOR2_X1 U1000 ( .A1(G131), .A2(KEYINPUT50), .ZN(n1301) );
NOR2_X1 U1001 ( .A1(KEYINPUT12), .A2(n1302), .ZN(n1300) );
INV_X1 U1002 ( .A(G137), .ZN(n1302) );
INV_X1 U1003 ( .A(n1053), .ZN(n1231) );
NAND2_X1 U1004 ( .A1(n1259), .A2(n1260), .ZN(n1053) );
XOR2_X1 U1005 ( .A(n1086), .B(n1087), .Z(n1260) );
INV_X1 U1006 ( .A(G478), .ZN(n1087) );
NOR2_X1 U1007 ( .A1(n1134), .A2(G902), .ZN(n1086) );
XOR2_X1 U1008 ( .A(n1303), .B(n1304), .Z(n1134) );
XOR2_X1 U1009 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U1010 ( .A(G107), .B(n1307), .Z(n1306) );
AND3_X1 U1011 ( .A1(G217), .A2(n1109), .A3(G234), .ZN(n1307) );
XNOR2_X1 U1012 ( .A(G116), .B(n1308), .ZN(n1303) );
XOR2_X1 U1013 ( .A(G134), .B(G122), .Z(n1308) );
XOR2_X1 U1014 ( .A(n1309), .B(G475), .Z(n1259) );
NAND2_X1 U1015 ( .A1(n1275), .A2(n1141), .ZN(n1309) );
NAND3_X1 U1016 ( .A1(n1310), .A2(n1311), .A3(n1312), .ZN(n1141) );
NAND2_X1 U1017 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
NAND2_X1 U1018 ( .A1(KEYINPUT62), .A2(n1315), .ZN(n1311) );
NAND2_X1 U1019 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XNOR2_X1 U1020 ( .A(n1313), .B(KEYINPUT16), .ZN(n1317) );
NAND2_X1 U1021 ( .A1(n1318), .A2(n1319), .ZN(n1310) );
INV_X1 U1022 ( .A(KEYINPUT62), .ZN(n1319) );
NAND2_X1 U1023 ( .A1(n1320), .A2(n1321), .ZN(n1318) );
OR3_X1 U1024 ( .A1(n1313), .A2(n1314), .A3(KEYINPUT16), .ZN(n1321) );
INV_X1 U1025 ( .A(n1316), .ZN(n1314) );
XOR2_X1 U1026 ( .A(n1322), .B(n1323), .Z(n1316) );
XOR2_X1 U1027 ( .A(G143), .B(G131), .Z(n1323) );
XOR2_X1 U1028 ( .A(n1324), .B(n1325), .Z(n1322) );
NOR3_X1 U1029 ( .A1(n1326), .A2(G953), .A3(n1327), .ZN(n1325) );
XOR2_X1 U1030 ( .A(n1296), .B(KEYINPUT54), .Z(n1327) );
INV_X1 U1031 ( .A(G237), .ZN(n1296) );
INV_X1 U1032 ( .A(G214), .ZN(n1326) );
NAND3_X1 U1033 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1324) );
INV_X1 U1034 ( .A(n1283), .ZN(n1330) );
NOR3_X1 U1035 ( .A1(n1331), .A2(n1225), .A3(n1332), .ZN(n1283) );
NAND2_X1 U1036 ( .A1(n1284), .A2(n1333), .ZN(n1329) );
INV_X1 U1037 ( .A(KEYINPUT28), .ZN(n1333) );
NAND2_X1 U1038 ( .A1(n1334), .A2(n1335), .ZN(n1284) );
NAND2_X1 U1039 ( .A1(n1336), .A2(n1225), .ZN(n1335) );
XOR2_X1 U1040 ( .A(n1332), .B(n1331), .Z(n1336) );
NAND3_X1 U1041 ( .A1(n1331), .A2(n1332), .A3(G146), .ZN(n1334) );
NAND2_X1 U1042 ( .A1(n1337), .A2(KEYINPUT28), .ZN(n1328) );
XOR2_X1 U1043 ( .A(n1225), .B(n1338), .Z(n1337) );
NAND2_X1 U1044 ( .A1(n1331), .A2(n1332), .ZN(n1338) );
INV_X1 U1045 ( .A(G125), .ZN(n1332) );
XOR2_X1 U1046 ( .A(G140), .B(KEYINPUT47), .Z(n1331) );
NAND2_X1 U1047 ( .A1(KEYINPUT16), .A2(n1313), .ZN(n1320) );
AND2_X1 U1048 ( .A1(n1339), .A2(n1340), .ZN(n1313) );
NAND2_X1 U1049 ( .A1(n1341), .A2(G122), .ZN(n1340) );
NAND2_X1 U1050 ( .A1(n1342), .A2(n1249), .ZN(n1339) );
XNOR2_X1 U1051 ( .A(KEYINPUT46), .B(n1341), .ZN(n1342) );
XOR2_X1 U1052 ( .A(G104), .B(n1261), .Z(n1341) );
INV_X1 U1053 ( .A(n1206), .ZN(n1218) );
NAND2_X1 U1054 ( .A1(n1040), .A2(n1217), .ZN(n1206) );
NAND2_X1 U1055 ( .A1(n1049), .A2(n1343), .ZN(n1217) );
NAND3_X1 U1056 ( .A1(n1119), .A2(n1242), .A3(G902), .ZN(n1343) );
NOR2_X1 U1057 ( .A1(n1109), .A2(G898), .ZN(n1119) );
NAND3_X1 U1058 ( .A1(n1242), .A2(n1109), .A3(G952), .ZN(n1049) );
NAND2_X1 U1059 ( .A1(G237), .A2(G234), .ZN(n1242) );
AND2_X1 U1060 ( .A1(n1344), .A2(n1064), .ZN(n1040) );
XOR2_X1 U1061 ( .A(n1345), .B(n1181), .Z(n1064) );
NAND2_X1 U1062 ( .A1(G210), .A2(n1346), .ZN(n1181) );
NAND2_X1 U1063 ( .A1(n1347), .A2(n1275), .ZN(n1345) );
XOR2_X1 U1064 ( .A(n1348), .B(n1221), .Z(n1347) );
XOR2_X1 U1065 ( .A(n1116), .B(n1118), .Z(n1221) );
XNOR2_X1 U1066 ( .A(n1349), .B(n1350), .ZN(n1118) );
XOR2_X1 U1067 ( .A(n1148), .B(n1274), .Z(n1350) );
XNOR2_X1 U1068 ( .A(G104), .B(G107), .ZN(n1274) );
XNOR2_X1 U1069 ( .A(G101), .B(KEYINPUT18), .ZN(n1148) );
XOR2_X1 U1070 ( .A(n1351), .B(KEYINPUT11), .Z(n1349) );
NAND2_X1 U1071 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
OR2_X1 U1072 ( .A1(n1354), .A2(n1261), .ZN(n1353) );
XOR2_X1 U1073 ( .A(n1355), .B(KEYINPUT39), .Z(n1352) );
NAND2_X1 U1074 ( .A1(n1354), .A2(n1261), .ZN(n1355) );
INV_X1 U1075 ( .A(G113), .ZN(n1261) );
XNOR2_X1 U1076 ( .A(n1255), .B(n1356), .ZN(n1354) );
NOR2_X1 U1077 ( .A1(G116), .A2(KEYINPUT58), .ZN(n1356) );
INV_X1 U1078 ( .A(G119), .ZN(n1255) );
XOR2_X1 U1079 ( .A(n1174), .B(n1249), .Z(n1116) );
INV_X1 U1080 ( .A(G122), .ZN(n1249) );
NOR2_X1 U1081 ( .A1(n1357), .A2(n1358), .ZN(n1348) );
XNOR2_X1 U1082 ( .A(KEYINPUT33), .B(n1223), .ZN(n1358) );
NAND2_X1 U1083 ( .A1(n1099), .A2(n1359), .ZN(n1223) );
NAND2_X1 U1084 ( .A1(G224), .A2(n1109), .ZN(n1359) );
INV_X1 U1085 ( .A(n1222), .ZN(n1357) );
NAND3_X1 U1086 ( .A1(n1360), .A2(n1109), .A3(G224), .ZN(n1222) );
INV_X1 U1087 ( .A(G953), .ZN(n1109) );
INV_X1 U1088 ( .A(n1099), .ZN(n1360) );
XOR2_X1 U1089 ( .A(n1171), .B(G125), .Z(n1099) );
XNOR2_X1 U1090 ( .A(n1225), .B(n1305), .ZN(n1171) );
XOR2_X1 U1091 ( .A(G128), .B(G143), .Z(n1305) );
INV_X1 U1092 ( .A(G146), .ZN(n1225) );
XNOR2_X1 U1093 ( .A(n1234), .B(KEYINPUT36), .ZN(n1344) );
INV_X1 U1094 ( .A(n1063), .ZN(n1234) );
NAND2_X1 U1095 ( .A1(G214), .A2(n1346), .ZN(n1063) );
NAND2_X1 U1096 ( .A1(n1361), .A2(n1275), .ZN(n1346) );
INV_X1 U1097 ( .A(G902), .ZN(n1275) );
XOR2_X1 U1098 ( .A(KEYINPUT25), .B(G237), .Z(n1361) );
INV_X1 U1099 ( .A(G110), .ZN(n1174) );
endmodule


