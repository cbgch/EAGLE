//Key = 1010001101111110010101110101010011010010111011011101110001010110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341;

XNOR2_X1 U733 ( .A(G107), .B(n1015), .ZN(G9) );
NOR2_X1 U734 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
NOR2_X1 U736 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U737 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U738 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR3_X1 U739 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1024) );
INV_X1 U740 ( .A(n1031), .ZN(n1030) );
NAND3_X1 U741 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1028) );
NAND2_X1 U742 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NAND2_X1 U743 ( .A1(n1037), .A2(n1038), .ZN(n1032) );
NAND2_X1 U744 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
XOR2_X1 U745 ( .A(KEYINPUT42), .B(n1041), .Z(n1019) );
NOR2_X1 U746 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR4_X1 U747 ( .A1(n1044), .A2(n1023), .A3(n1029), .A4(n1045), .ZN(n1043) );
INV_X1 U748 ( .A(n1046), .ZN(n1023) );
NOR2_X1 U749 ( .A1(n1047), .A2(n1048), .ZN(n1044) );
NOR2_X1 U750 ( .A1(n1049), .A2(n1027), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U752 ( .A1(n1052), .A2(n1029), .ZN(n1051) );
AND2_X1 U753 ( .A1(n1046), .A2(n1053), .ZN(n1050) );
NAND3_X1 U754 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1018) );
NAND3_X1 U755 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
XOR2_X1 U756 ( .A(n1029), .B(KEYINPUT10), .Z(n1059) );
INV_X1 U757 ( .A(n1027), .ZN(n1057) );
NAND4_X1 U758 ( .A1(n1034), .A2(n1060), .A3(n1031), .A4(n1038), .ZN(n1027) );
INV_X1 U759 ( .A(n1045), .ZN(n1034) );
NOR3_X1 U760 ( .A1(n1061), .A2(G953), .A3(G952), .ZN(n1016) );
INV_X1 U761 ( .A(n1054), .ZN(n1061) );
NAND4_X1 U762 ( .A1(n1062), .A2(n1063), .A3(n1060), .A4(n1038), .ZN(n1054) );
XOR2_X1 U763 ( .A(n1064), .B(KEYINPUT32), .Z(n1063) );
NAND4_X1 U764 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1064) );
NOR4_X1 U765 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1068) );
XOR2_X1 U766 ( .A(KEYINPUT31), .B(n1073), .Z(n1072) );
NOR3_X1 U767 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1070) );
INV_X1 U768 ( .A(KEYINPUT29), .ZN(n1074) );
NOR2_X1 U769 ( .A1(KEYINPUT29), .A2(G475), .ZN(n1069) );
NAND2_X1 U770 ( .A1(G478), .A2(n1077), .ZN(n1065) );
XOR2_X1 U771 ( .A(n1031), .B(KEYINPUT30), .Z(n1062) );
XOR2_X1 U772 ( .A(n1078), .B(n1079), .Z(G72) );
NAND2_X1 U773 ( .A1(n1055), .A2(n1080), .ZN(n1079) );
NAND2_X1 U774 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(n1078) );
NAND3_X1 U776 ( .A1(n1085), .A2(n1086), .A3(G900), .ZN(n1084) );
NAND2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U778 ( .A1(G953), .A2(n1089), .ZN(n1087) );
NAND2_X1 U779 ( .A1(G227), .A2(n1089), .ZN(n1085) );
OR2_X1 U780 ( .A1(n1089), .A2(G953), .ZN(n1083) );
XNOR2_X1 U781 ( .A(n1090), .B(n1091), .ZN(n1089) );
NOR2_X1 U782 ( .A1(KEYINPUT36), .A2(n1092), .ZN(n1091) );
XOR2_X1 U783 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U784 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND2_X1 U785 ( .A1(KEYINPUT51), .A2(n1097), .ZN(n1095) );
NAND2_X1 U786 ( .A1(n1098), .A2(n1099), .ZN(n1090) );
NAND2_X1 U787 ( .A1(G125), .A2(n1100), .ZN(n1099) );
XOR2_X1 U788 ( .A(KEYINPUT14), .B(n1101), .Z(n1098) );
NOR2_X1 U789 ( .A1(G125), .A2(n1100), .ZN(n1101) );
NAND2_X1 U790 ( .A1(n1102), .A2(n1103), .ZN(G69) );
NAND2_X1 U791 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XNOR2_X1 U792 ( .A(KEYINPUT49), .B(n1106), .ZN(n1105) );
XNOR2_X1 U793 ( .A(n1107), .B(KEYINPUT40), .ZN(n1104) );
XOR2_X1 U794 ( .A(KEYINPUT27), .B(n1108), .Z(n1102) );
NOR2_X1 U795 ( .A1(n1106), .A2(n1107), .ZN(n1108) );
XNOR2_X1 U796 ( .A(n1109), .B(n1110), .ZN(n1107) );
NOR2_X1 U797 ( .A1(G953), .A2(n1111), .ZN(n1110) );
NAND3_X1 U798 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1109) );
XOR2_X1 U799 ( .A(KEYINPUT12), .B(n1115), .Z(n1114) );
NOR2_X1 U800 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1113) );
NAND2_X1 U802 ( .A1(G953), .A2(n1118), .ZN(n1112) );
NAND2_X1 U803 ( .A1(n1119), .A2(G953), .ZN(n1106) );
XOR2_X1 U804 ( .A(n1120), .B(KEYINPUT46), .Z(n1119) );
NAND2_X1 U805 ( .A1(G898), .A2(G224), .ZN(n1120) );
NOR2_X1 U806 ( .A1(n1121), .A2(n1122), .ZN(G66) );
NOR2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U808 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U809 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U810 ( .A1(KEYINPUT39), .A2(n1129), .ZN(n1125) );
AND2_X1 U811 ( .A1(n1129), .A2(KEYINPUT39), .ZN(n1123) );
NOR3_X1 U812 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(G63) );
AND3_X1 U813 ( .A1(KEYINPUT20), .A2(n1055), .A3(n1133), .ZN(n1132) );
NOR2_X1 U814 ( .A1(KEYINPUT20), .A2(n1134), .ZN(n1131) );
NOR2_X1 U815 ( .A1(n1135), .A2(n1136), .ZN(n1130) );
XOR2_X1 U816 ( .A(n1137), .B(n1138), .Z(n1136) );
AND2_X1 U817 ( .A1(G478), .A2(n1139), .ZN(n1138) );
NOR2_X1 U818 ( .A1(n1140), .A2(n1141), .ZN(n1137) );
AND2_X1 U819 ( .A1(n1141), .A2(n1140), .ZN(n1135) );
INV_X1 U820 ( .A(KEYINPUT47), .ZN(n1141) );
NOR2_X1 U821 ( .A1(n1121), .A2(n1142), .ZN(G60) );
XOR2_X1 U822 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U823 ( .A1(n1076), .A2(n1128), .ZN(n1144) );
XNOR2_X1 U824 ( .A(n1145), .B(n1146), .ZN(G6) );
NAND2_X1 U825 ( .A1(n1147), .A2(KEYINPUT48), .ZN(n1146) );
XNOR2_X1 U826 ( .A(G104), .B(KEYINPUT61), .ZN(n1147) );
NOR3_X1 U827 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(G57) );
AND3_X1 U828 ( .A1(KEYINPUT55), .A2(n1055), .A3(n1133), .ZN(n1150) );
NOR2_X1 U829 ( .A1(KEYINPUT55), .A2(n1134), .ZN(n1149) );
XOR2_X1 U830 ( .A(n1151), .B(n1152), .Z(n1148) );
XOR2_X1 U831 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U832 ( .A1(KEYINPUT35), .A2(n1155), .ZN(n1153) );
XOR2_X1 U833 ( .A(KEYINPUT63), .B(n1156), .Z(n1151) );
AND2_X1 U834 ( .A1(G472), .A2(n1139), .ZN(n1156) );
NOR2_X1 U835 ( .A1(n1121), .A2(n1157), .ZN(G54) );
XOR2_X1 U836 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U837 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U838 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U839 ( .A1(KEYINPUT15), .A2(n1164), .ZN(n1163) );
NAND2_X1 U840 ( .A1(n1165), .A2(n1166), .ZN(n1160) );
NAND2_X1 U841 ( .A1(KEYINPUT26), .A2(n1167), .ZN(n1166) );
NAND2_X1 U842 ( .A1(KEYINPUT13), .A2(n1168), .ZN(n1165) );
INV_X1 U843 ( .A(n1167), .ZN(n1168) );
NAND2_X1 U844 ( .A1(n1139), .A2(G469), .ZN(n1167) );
INV_X1 U845 ( .A(n1128), .ZN(n1139) );
XOR2_X1 U846 ( .A(n1169), .B(n1170), .Z(n1158) );
NOR2_X1 U847 ( .A1(KEYINPUT28), .A2(n1171), .ZN(n1170) );
XNOR2_X1 U848 ( .A(KEYINPUT6), .B(n1172), .ZN(n1169) );
NOR2_X1 U849 ( .A1(KEYINPUT5), .A2(n1173), .ZN(n1172) );
XOR2_X1 U850 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND2_X1 U851 ( .A1(KEYINPUT45), .A2(n1176), .ZN(n1174) );
XOR2_X1 U852 ( .A(n1177), .B(n1178), .Z(n1176) );
NOR2_X1 U853 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NOR2_X1 U854 ( .A1(KEYINPUT0), .A2(n1181), .ZN(n1180) );
AND2_X1 U855 ( .A1(KEYINPUT59), .A2(n1181), .ZN(n1179) );
NOR2_X1 U856 ( .A1(n1121), .A2(n1182), .ZN(G51) );
XOR2_X1 U857 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U858 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U859 ( .A1(n1187), .A2(n1128), .ZN(n1186) );
NAND2_X1 U860 ( .A1(G902), .A2(n1021), .ZN(n1128) );
NAND3_X1 U861 ( .A1(n1081), .A2(n1111), .A3(n1188), .ZN(n1021) );
XOR2_X1 U862 ( .A(n1082), .B(KEYINPUT56), .Z(n1188) );
AND4_X1 U863 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1111) );
AND4_X1 U864 ( .A1(n1015), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1192) );
NAND3_X1 U865 ( .A1(n1196), .A2(n1046), .A3(n1197), .ZN(n1015) );
NOR2_X1 U866 ( .A1(n1145), .A2(n1198), .ZN(n1191) );
NOR3_X1 U867 ( .A1(n1029), .A2(n1199), .A3(n1052), .ZN(n1198) );
AND3_X1 U868 ( .A1(n1197), .A2(n1046), .A3(n1053), .ZN(n1145) );
AND4_X1 U869 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1081) );
NOR4_X1 U870 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203) );
NOR3_X1 U871 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1207) );
XNOR2_X1 U872 ( .A(KEYINPUT54), .B(n1211), .ZN(n1210) );
NAND3_X1 U873 ( .A1(n1212), .A2(n1213), .A3(n1196), .ZN(n1208) );
OR2_X1 U874 ( .A1(n1214), .A2(n1052), .ZN(n1202) );
NAND2_X1 U875 ( .A1(KEYINPUT11), .A2(n1215), .ZN(n1185) );
INV_X1 U876 ( .A(n1134), .ZN(n1121) );
NAND2_X1 U877 ( .A1(G953), .A2(n1133), .ZN(n1134) );
XOR2_X1 U878 ( .A(G952), .B(KEYINPUT21), .Z(n1133) );
NAND2_X1 U879 ( .A1(n1216), .A2(n1217), .ZN(G48) );
NAND2_X1 U880 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XOR2_X1 U881 ( .A(KEYINPUT41), .B(n1220), .Z(n1216) );
NOR2_X1 U882 ( .A1(n1218), .A2(n1219), .ZN(n1220) );
INV_X1 U883 ( .A(G146), .ZN(n1219) );
INV_X1 U884 ( .A(n1082), .ZN(n1218) );
NAND3_X1 U885 ( .A1(n1053), .A2(n1213), .A3(n1221), .ZN(n1082) );
INV_X1 U886 ( .A(n1222), .ZN(n1221) );
XOR2_X1 U887 ( .A(G143), .B(n1223), .Z(G45) );
NOR2_X1 U888 ( .A1(n1224), .A2(n1214), .ZN(n1223) );
NAND3_X1 U889 ( .A1(n1211), .A2(n1212), .A3(n1225), .ZN(n1214) );
AND3_X1 U890 ( .A1(n1213), .A2(n1226), .A3(n1227), .ZN(n1225) );
XOR2_X1 U891 ( .A(n1052), .B(KEYINPUT18), .Z(n1224) );
XOR2_X1 U892 ( .A(n1100), .B(n1200), .Z(G42) );
NAND3_X1 U893 ( .A1(n1053), .A2(n1058), .A3(n1228), .ZN(n1200) );
XNOR2_X1 U894 ( .A(n1201), .B(n1229), .ZN(G39) );
NOR2_X1 U895 ( .A1(KEYINPUT34), .A2(n1230), .ZN(n1229) );
NAND3_X1 U896 ( .A1(n1231), .A2(n1228), .A3(n1232), .ZN(n1201) );
XOR2_X1 U897 ( .A(G134), .B(n1206), .Z(G36) );
AND3_X1 U898 ( .A1(n1228), .A2(n1196), .A3(n1233), .ZN(n1206) );
NAND2_X1 U899 ( .A1(n1234), .A2(n1235), .ZN(G33) );
NAND2_X1 U900 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U901 ( .A1(G131), .A2(n1238), .ZN(n1234) );
NAND2_X1 U902 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
NAND2_X1 U903 ( .A1(KEYINPUT37), .A2(n1205), .ZN(n1240) );
OR2_X1 U904 ( .A1(n1236), .A2(KEYINPUT37), .ZN(n1239) );
AND2_X1 U905 ( .A1(KEYINPUT22), .A2(n1205), .ZN(n1236) );
AND3_X1 U906 ( .A1(n1228), .A2(n1053), .A3(n1233), .ZN(n1205) );
AND2_X1 U907 ( .A1(n1048), .A2(n1213), .ZN(n1228) );
AND3_X1 U908 ( .A1(n1212), .A2(n1038), .A3(n1031), .ZN(n1048) );
XOR2_X1 U909 ( .A(G128), .B(n1241), .Z(G30) );
NOR3_X1 U910 ( .A1(n1222), .A2(n1242), .A3(n1026), .ZN(n1241) );
INV_X1 U911 ( .A(n1196), .ZN(n1026) );
XOR2_X1 U912 ( .A(n1213), .B(KEYINPUT62), .Z(n1242) );
NAND3_X1 U913 ( .A1(n1211), .A2(n1212), .A3(n1231), .ZN(n1222) );
XNOR2_X1 U914 ( .A(G101), .B(n1243), .ZN(G3) );
NAND4_X1 U915 ( .A1(n1212), .A2(n1244), .A3(n1233), .A4(n1245), .ZN(n1243) );
NOR2_X1 U916 ( .A1(n1029), .A2(n1246), .ZN(n1245) );
XNOR2_X1 U917 ( .A(KEYINPUT50), .B(n1247), .ZN(n1246) );
INV_X1 U918 ( .A(n1232), .ZN(n1029) );
XNOR2_X1 U919 ( .A(n1204), .B(n1248), .ZN(G27) );
NAND2_X1 U920 ( .A1(KEYINPUT7), .A2(G125), .ZN(n1248) );
AND4_X1 U921 ( .A1(n1053), .A2(n1047), .A3(n1058), .A4(n1213), .ZN(n1204) );
NAND2_X1 U922 ( .A1(n1045), .A2(n1249), .ZN(n1213) );
NAND4_X1 U923 ( .A1(G953), .A2(G902), .A3(n1250), .A4(n1251), .ZN(n1249) );
INV_X1 U924 ( .A(G900), .ZN(n1251) );
XNOR2_X1 U925 ( .A(G122), .B(n1189), .ZN(G24) );
NAND4_X1 U926 ( .A1(n1252), .A2(n1046), .A3(n1227), .A4(n1226), .ZN(n1189) );
NOR2_X1 U927 ( .A1(n1071), .A2(n1253), .ZN(n1046) );
XOR2_X1 U928 ( .A(KEYINPUT44), .B(n1067), .Z(n1253) );
XNOR2_X1 U929 ( .A(G119), .B(n1190), .ZN(G21) );
NAND3_X1 U930 ( .A1(n1232), .A2(n1231), .A3(n1252), .ZN(n1190) );
INV_X1 U931 ( .A(n1209), .ZN(n1231) );
NAND2_X1 U932 ( .A1(n1254), .A2(n1071), .ZN(n1209) );
INV_X1 U933 ( .A(n1067), .ZN(n1254) );
XOR2_X1 U934 ( .A(n1255), .B(n1195), .Z(G18) );
NAND3_X1 U935 ( .A1(n1233), .A2(n1196), .A3(n1252), .ZN(n1195) );
AND2_X1 U936 ( .A1(n1047), .A2(n1247), .ZN(n1252) );
AND2_X1 U937 ( .A1(n1211), .A2(n1060), .ZN(n1047) );
XNOR2_X1 U938 ( .A(n1244), .B(KEYINPUT17), .ZN(n1211) );
NOR2_X1 U939 ( .A1(n1226), .A2(n1256), .ZN(n1196) );
XNOR2_X1 U940 ( .A(G113), .B(n1194), .ZN(G15) );
NAND4_X1 U941 ( .A1(n1233), .A2(n1053), .A3(n1257), .A4(n1060), .ZN(n1194) );
INV_X1 U942 ( .A(n1036), .ZN(n1060) );
NAND2_X1 U943 ( .A1(n1040), .A2(n1258), .ZN(n1036) );
AND2_X1 U944 ( .A1(n1247), .A2(n1244), .ZN(n1257) );
AND2_X1 U945 ( .A1(n1256), .A2(n1226), .ZN(n1053) );
INV_X1 U946 ( .A(n1052), .ZN(n1233) );
NAND2_X1 U947 ( .A1(n1067), .A2(n1071), .ZN(n1052) );
XOR2_X1 U948 ( .A(n1177), .B(n1193), .Z(G12) );
NAND3_X1 U949 ( .A1(n1058), .A2(n1197), .A3(n1232), .ZN(n1193) );
NOR2_X1 U950 ( .A1(n1227), .A2(n1226), .ZN(n1232) );
NAND2_X1 U951 ( .A1(n1259), .A2(n1066), .ZN(n1226) );
NAND2_X1 U952 ( .A1(n1075), .A2(n1076), .ZN(n1066) );
OR2_X1 U953 ( .A1(n1076), .A2(n1075), .ZN(n1259) );
NOR2_X1 U954 ( .A1(n1143), .A2(G902), .ZN(n1075) );
XOR2_X1 U955 ( .A(n1260), .B(n1261), .Z(n1143) );
XOR2_X1 U956 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U957 ( .A(G131), .B(G122), .Z(n1263) );
XOR2_X1 U958 ( .A(KEYINPUT38), .B(KEYINPUT2), .Z(n1262) );
XOR2_X1 U959 ( .A(n1264), .B(n1265), .Z(n1260) );
XOR2_X1 U960 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U961 ( .A(n1268), .B(n1269), .Z(n1264) );
NAND2_X1 U962 ( .A1(n1270), .A2(G214), .ZN(n1268) );
INV_X1 U963 ( .A(G475), .ZN(n1076) );
INV_X1 U964 ( .A(n1256), .ZN(n1227) );
NOR2_X1 U965 ( .A1(n1073), .A2(n1271), .ZN(n1256) );
AND2_X1 U966 ( .A1(G478), .A2(n1077), .ZN(n1271) );
NOR2_X1 U967 ( .A1(n1077), .A2(G478), .ZN(n1073) );
OR2_X1 U968 ( .A1(n1140), .A2(G902), .ZN(n1077) );
XNOR2_X1 U969 ( .A(n1272), .B(n1273), .ZN(n1140) );
XOR2_X1 U970 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U971 ( .A(n1276), .B(n1277), .Z(n1275) );
NOR2_X1 U972 ( .A1(n1278), .A2(n1279), .ZN(n1276) );
INV_X1 U973 ( .A(G217), .ZN(n1279) );
XOR2_X1 U974 ( .A(G116), .B(G107), .Z(n1274) );
XOR2_X1 U975 ( .A(n1280), .B(n1281), .Z(n1272) );
XOR2_X1 U976 ( .A(G128), .B(G122), .Z(n1281) );
XNOR2_X1 U977 ( .A(G143), .B(KEYINPUT33), .ZN(n1280) );
INV_X1 U978 ( .A(n1199), .ZN(n1197) );
NAND3_X1 U979 ( .A1(n1244), .A2(n1247), .A3(n1212), .ZN(n1199) );
NOR2_X1 U980 ( .A1(n1040), .A2(n1039), .ZN(n1212) );
INV_X1 U981 ( .A(n1258), .ZN(n1039) );
NAND2_X1 U982 ( .A1(G221), .A2(n1282), .ZN(n1258) );
XOR2_X1 U983 ( .A(n1283), .B(G469), .Z(n1040) );
NAND4_X1 U984 ( .A1(n1284), .A2(n1285), .A3(n1286), .A4(n1287), .ZN(n1283) );
OR3_X1 U985 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n1287) );
INV_X1 U986 ( .A(KEYINPUT53), .ZN(n1288) );
NAND2_X1 U987 ( .A1(n1290), .A2(n1289), .ZN(n1286) );
NAND2_X1 U988 ( .A1(KEYINPUT52), .A2(n1291), .ZN(n1289) );
XOR2_X1 U989 ( .A(n1181), .B(n1292), .Z(n1290) );
XOR2_X1 U990 ( .A(G110), .B(n1175), .Z(n1292) );
NOR2_X1 U991 ( .A1(n1088), .A2(G953), .ZN(n1175) );
INV_X1 U992 ( .A(G227), .ZN(n1088) );
XNOR2_X1 U993 ( .A(n1100), .B(KEYINPUT9), .ZN(n1181) );
INV_X1 U994 ( .A(G140), .ZN(n1100) );
OR2_X1 U995 ( .A1(n1291), .A2(KEYINPUT53), .ZN(n1284) );
XNOR2_X1 U996 ( .A(n1162), .B(n1293), .ZN(n1291) );
XOR2_X1 U997 ( .A(n1294), .B(n1171), .Z(n1293) );
XNOR2_X1 U998 ( .A(G104), .B(n1295), .ZN(n1171) );
INV_X1 U999 ( .A(n1093), .ZN(n1162) );
XOR2_X1 U1000 ( .A(n1296), .B(n1297), .Z(n1093) );
NAND2_X1 U1001 ( .A1(n1045), .A2(n1298), .ZN(n1247) );
NAND4_X1 U1002 ( .A1(G953), .A2(G902), .A3(n1250), .A4(n1118), .ZN(n1298) );
INV_X1 U1003 ( .A(G898), .ZN(n1118) );
NAND3_X1 U1004 ( .A1(n1250), .A2(n1055), .A3(G952), .ZN(n1045) );
NAND2_X1 U1005 ( .A1(G237), .A2(G234), .ZN(n1250) );
NOR2_X1 U1006 ( .A1(n1031), .A2(n1035), .ZN(n1244) );
INV_X1 U1007 ( .A(n1038), .ZN(n1035) );
NAND2_X1 U1008 ( .A1(G214), .A2(n1299), .ZN(n1038) );
XNOR2_X1 U1009 ( .A(n1300), .B(n1187), .ZN(n1031) );
NAND2_X1 U1010 ( .A1(G210), .A2(n1299), .ZN(n1187) );
NAND2_X1 U1011 ( .A1(n1301), .A2(n1285), .ZN(n1299) );
INV_X1 U1012 ( .A(G237), .ZN(n1301) );
NAND2_X1 U1013 ( .A1(n1302), .A2(n1285), .ZN(n1300) );
XOR2_X1 U1014 ( .A(n1215), .B(n1183), .Z(n1302) );
XOR2_X1 U1015 ( .A(n1303), .B(n1304), .Z(n1183) );
XNOR2_X1 U1016 ( .A(G125), .B(n1305), .ZN(n1303) );
AND2_X1 U1017 ( .A1(n1055), .A2(G224), .ZN(n1305) );
NAND3_X1 U1018 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1215) );
NAND2_X1 U1019 ( .A1(KEYINPUT43), .A2(n1309), .ZN(n1308) );
NAND3_X1 U1020 ( .A1(n1116), .A2(n1310), .A3(n1117), .ZN(n1307) );
INV_X1 U1021 ( .A(n1311), .ZN(n1117) );
NAND2_X1 U1022 ( .A1(n1311), .A2(n1312), .ZN(n1306) );
NAND2_X1 U1023 ( .A1(n1313), .A2(n1310), .ZN(n1312) );
INV_X1 U1024 ( .A(KEYINPUT43), .ZN(n1310) );
XOR2_X1 U1025 ( .A(KEYINPUT8), .B(n1116), .Z(n1313) );
INV_X1 U1026 ( .A(n1309), .ZN(n1116) );
XOR2_X1 U1027 ( .A(n1314), .B(n1315), .Z(n1309) );
XOR2_X1 U1028 ( .A(n1295), .B(n1316), .Z(n1315) );
NOR2_X1 U1029 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NOR2_X1 U1030 ( .A1(KEYINPUT57), .A2(G116), .ZN(n1318) );
NOR2_X1 U1031 ( .A1(KEYINPUT16), .A2(n1255), .ZN(n1317) );
XOR2_X1 U1032 ( .A(G101), .B(G107), .Z(n1295) );
XNOR2_X1 U1033 ( .A(G119), .B(n1267), .ZN(n1314) );
XOR2_X1 U1034 ( .A(G104), .B(G113), .Z(n1267) );
XOR2_X1 U1035 ( .A(n1177), .B(G122), .Z(n1311) );
NOR2_X1 U1036 ( .A1(n1071), .A2(n1067), .ZN(n1058) );
XNOR2_X1 U1037 ( .A(n1319), .B(n1127), .ZN(n1067) );
NAND2_X1 U1038 ( .A1(G217), .A2(n1282), .ZN(n1127) );
NAND2_X1 U1039 ( .A1(G234), .A2(n1285), .ZN(n1282) );
OR2_X1 U1040 ( .A1(n1129), .A2(G902), .ZN(n1319) );
XOR2_X1 U1041 ( .A(n1320), .B(n1321), .Z(n1129) );
XOR2_X1 U1042 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U1043 ( .A(G110), .B(n1324), .Z(n1323) );
NOR2_X1 U1044 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1045 ( .A(n1327), .B(KEYINPUT19), .Z(n1326) );
NAND2_X1 U1046 ( .A1(G146), .A2(n1269), .ZN(n1327) );
NOR2_X1 U1047 ( .A1(G146), .A2(n1269), .ZN(n1325) );
XOR2_X1 U1048 ( .A(G125), .B(G140), .Z(n1269) );
NOR2_X1 U1049 ( .A1(n1328), .A2(n1278), .ZN(n1322) );
NAND2_X1 U1050 ( .A1(n1329), .A2(n1055), .ZN(n1278) );
INV_X1 U1051 ( .A(G953), .ZN(n1055) );
XOR2_X1 U1052 ( .A(KEYINPUT24), .B(G234), .Z(n1329) );
INV_X1 U1053 ( .A(G221), .ZN(n1328) );
XNOR2_X1 U1054 ( .A(G119), .B(n1330), .ZN(n1320) );
XOR2_X1 U1055 ( .A(G137), .B(G128), .Z(n1330) );
XNOR2_X1 U1056 ( .A(n1331), .B(G472), .ZN(n1071) );
NAND2_X1 U1057 ( .A1(n1332), .A2(n1285), .ZN(n1331) );
INV_X1 U1058 ( .A(G902), .ZN(n1285) );
XNOR2_X1 U1059 ( .A(n1155), .B(n1333), .ZN(n1332) );
XOR2_X1 U1060 ( .A(KEYINPUT60), .B(n1334), .Z(n1333) );
INV_X1 U1061 ( .A(n1154), .ZN(n1334) );
XOR2_X1 U1062 ( .A(n1335), .B(G101), .Z(n1154) );
NAND2_X1 U1063 ( .A1(n1270), .A2(G210), .ZN(n1335) );
NOR2_X1 U1064 ( .A1(G953), .A2(G237), .ZN(n1270) );
XNOR2_X1 U1065 ( .A(n1336), .B(n1337), .ZN(n1155) );
XOR2_X1 U1066 ( .A(n1304), .B(n1164), .Z(n1337) );
INV_X1 U1067 ( .A(n1294), .ZN(n1164) );
XOR2_X1 U1068 ( .A(n1096), .B(n1338), .Z(n1294) );
NOR2_X1 U1069 ( .A1(KEYINPUT58), .A2(n1097), .ZN(n1338) );
XOR2_X1 U1070 ( .A(n1230), .B(n1277), .Z(n1097) );
XOR2_X1 U1071 ( .A(G134), .B(KEYINPUT3), .Z(n1277) );
INV_X1 U1072 ( .A(G137), .ZN(n1230) );
XOR2_X1 U1073 ( .A(n1237), .B(KEYINPUT25), .Z(n1096) );
INV_X1 U1074 ( .A(G131), .ZN(n1237) );
XNOR2_X1 U1075 ( .A(n1296), .B(n1339), .ZN(n1304) );
NOR2_X1 U1076 ( .A1(KEYINPUT1), .A2(n1297), .ZN(n1339) );
XNOR2_X1 U1077 ( .A(n1266), .B(KEYINPUT23), .ZN(n1297) );
XOR2_X1 U1078 ( .A(G143), .B(G146), .Z(n1266) );
INV_X1 U1079 ( .A(G128), .ZN(n1296) );
XOR2_X1 U1080 ( .A(n1340), .B(n1341), .Z(n1336) );
NOR2_X1 U1081 ( .A1(G119), .A2(KEYINPUT4), .ZN(n1341) );
XOR2_X1 U1082 ( .A(G113), .B(n1255), .Z(n1340) );
INV_X1 U1083 ( .A(G116), .ZN(n1255) );
INV_X1 U1084 ( .A(G110), .ZN(n1177) );
endmodule


