//Key = 0010110100100011010001000011011101011111101101011000001010111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385;

XNOR2_X1 U765 ( .A(G107), .B(n1052), .ZN(G9) );
NAND3_X1 U766 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
AND3_X1 U767 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
XNOR2_X1 U768 ( .A(n1059), .B(KEYINPUT7), .ZN(n1053) );
NOR2_X1 U769 ( .A1(n1060), .A2(n1061), .ZN(G75) );
NOR3_X1 U770 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
NOR3_X1 U771 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1063) );
NOR4_X1 U772 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1067) );
NOR2_X1 U773 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U774 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
AND2_X1 U775 ( .A1(n1058), .A2(n1054), .ZN(n1075) );
NOR3_X1 U776 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1074) );
NOR3_X1 U777 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NOR2_X1 U778 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U779 ( .A1(n1058), .A2(n1084), .ZN(n1077) );
NOR3_X1 U780 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1070) );
NOR2_X1 U781 ( .A1(KEYINPUT63), .A2(n1088), .ZN(n1069) );
INV_X1 U782 ( .A(n1089), .ZN(n1088) );
NOR2_X1 U783 ( .A1(n1090), .A2(n1091), .ZN(n1066) );
AND2_X1 U784 ( .A1(n1089), .A2(KEYINPUT63), .ZN(n1091) );
NAND3_X1 U785 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1062) );
NAND4_X1 U786 ( .A1(n1090), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1094) );
NAND2_X1 U787 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
INV_X1 U788 ( .A(n1086), .ZN(n1095) );
INV_X1 U789 ( .A(n1068), .ZN(n1090) );
NOR3_X1 U790 ( .A1(n1100), .A2(G953), .A3(G952), .ZN(n1060) );
INV_X1 U791 ( .A(n1092), .ZN(n1100) );
NAND4_X1 U792 ( .A1(n1101), .A2(n1096), .A3(n1102), .A4(n1103), .ZN(n1092) );
NOR3_X1 U793 ( .A1(n1083), .A2(n1079), .A3(n1104), .ZN(n1103) );
XOR2_X1 U794 ( .A(n1082), .B(KEYINPUT38), .Z(n1104) );
XNOR2_X1 U795 ( .A(n1105), .B(n1106), .ZN(n1102) );
NAND2_X1 U796 ( .A1(KEYINPUT47), .A2(n1107), .ZN(n1105) );
XOR2_X1 U797 ( .A(n1108), .B(n1109), .Z(G72) );
XOR2_X1 U798 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U799 ( .A1(G953), .A2(n1112), .ZN(n1111) );
NAND2_X1 U800 ( .A1(G900), .A2(G227), .ZN(n1112) );
NAND3_X1 U801 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1110) );
OR2_X1 U802 ( .A1(n1093), .A2(G900), .ZN(n1115) );
NAND2_X1 U803 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NAND2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
OR2_X1 U805 ( .A1(n1120), .A2(KEYINPUT5), .ZN(n1119) );
NAND3_X1 U806 ( .A1(n1121), .A2(n1122), .A3(KEYINPUT5), .ZN(n1113) );
NAND2_X1 U807 ( .A1(KEYINPUT15), .A2(n1123), .ZN(n1122) );
NAND2_X1 U808 ( .A1(n1124), .A2(n1118), .ZN(n1123) );
INV_X1 U809 ( .A(n1116), .ZN(n1124) );
XNOR2_X1 U810 ( .A(n1125), .B(n1126), .ZN(n1116) );
XOR2_X1 U811 ( .A(n1127), .B(n1128), .Z(n1126) );
XNOR2_X1 U812 ( .A(G131), .B(KEYINPUT35), .ZN(n1128) );
NAND2_X1 U813 ( .A1(KEYINPUT43), .A2(n1129), .ZN(n1127) );
XNOR2_X1 U814 ( .A(n1130), .B(n1131), .ZN(n1125) );
NAND2_X1 U815 ( .A1(n1118), .A2(n1120), .ZN(n1121) );
INV_X1 U816 ( .A(KEYINPUT15), .ZN(n1120) );
XNOR2_X1 U817 ( .A(n1132), .B(n1133), .ZN(n1118) );
XNOR2_X1 U818 ( .A(KEYINPUT58), .B(n1134), .ZN(n1133) );
NOR2_X1 U819 ( .A1(n1135), .A2(G953), .ZN(n1108) );
XOR2_X1 U820 ( .A(n1136), .B(n1137), .Z(G69) );
NOR3_X1 U821 ( .A1(n1093), .A2(KEYINPUT41), .A3(n1138), .ZN(n1137) );
NOR2_X1 U822 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NAND2_X1 U823 ( .A1(n1141), .A2(n1142), .ZN(n1136) );
NAND2_X1 U824 ( .A1(KEYINPUT13), .A2(n1143), .ZN(n1142) );
XOR2_X1 U825 ( .A(n1144), .B(n1145), .Z(n1141) );
NOR2_X1 U826 ( .A1(KEYINPUT13), .A2(n1143), .ZN(n1145) );
NAND2_X1 U827 ( .A1(n1146), .A2(n1147), .ZN(n1143) );
NAND2_X1 U828 ( .A1(G953), .A2(n1140), .ZN(n1147) );
XOR2_X1 U829 ( .A(n1148), .B(KEYINPUT28), .Z(n1146) );
NAND2_X1 U830 ( .A1(n1093), .A2(n1149), .ZN(n1144) );
NOR2_X1 U831 ( .A1(n1150), .A2(n1151), .ZN(G66) );
XOR2_X1 U832 ( .A(KEYINPUT24), .B(n1152), .Z(n1151) );
XOR2_X1 U833 ( .A(n1153), .B(n1154), .Z(n1150) );
NOR2_X1 U834 ( .A1(n1155), .A2(n1156), .ZN(n1153) );
NOR2_X1 U835 ( .A1(n1152), .A2(n1157), .ZN(G63) );
XOR2_X1 U836 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U837 ( .A1(n1160), .A2(n1156), .ZN(n1158) );
NOR2_X1 U838 ( .A1(n1152), .A2(n1161), .ZN(G60) );
XOR2_X1 U839 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND3_X1 U840 ( .A1(n1164), .A2(n1064), .A3(G475), .ZN(n1162) );
XNOR2_X1 U841 ( .A(KEYINPUT25), .B(n1165), .ZN(n1164) );
XOR2_X1 U842 ( .A(G104), .B(n1166), .Z(G6) );
NOR2_X1 U843 ( .A1(n1152), .A2(n1167), .ZN(G57) );
XOR2_X1 U844 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U845 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U846 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
NAND2_X1 U847 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
INV_X1 U848 ( .A(KEYINPUT1), .ZN(n1175) );
NAND3_X1 U849 ( .A1(n1176), .A2(n1177), .A3(KEYINPUT1), .ZN(n1172) );
XOR2_X1 U850 ( .A(n1178), .B(n1179), .Z(n1168) );
NOR2_X1 U851 ( .A1(n1180), .A2(n1156), .ZN(n1179) );
NOR2_X1 U852 ( .A1(n1152), .A2(n1181), .ZN(G54) );
XOR2_X1 U853 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U854 ( .A(n1184), .B(n1185), .Z(n1182) );
NOR2_X1 U855 ( .A1(n1186), .A2(n1156), .ZN(n1185) );
NAND2_X1 U856 ( .A1(KEYINPUT21), .A2(n1187), .ZN(n1184) );
NOR2_X1 U857 ( .A1(n1152), .A2(n1188), .ZN(G51) );
XOR2_X1 U858 ( .A(n1148), .B(n1189), .Z(n1188) );
XOR2_X1 U859 ( .A(n1190), .B(n1191), .Z(n1189) );
NOR2_X1 U860 ( .A1(n1192), .A2(n1156), .ZN(n1191) );
NAND2_X1 U861 ( .A1(G902), .A2(n1064), .ZN(n1156) );
NAND2_X1 U862 ( .A1(n1193), .A2(n1135), .ZN(n1064) );
AND4_X1 U863 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1135) );
NOR4_X1 U864 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
NOR2_X1 U865 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NOR2_X1 U866 ( .A1(n1204), .A2(n1205), .ZN(n1202) );
NOR2_X1 U867 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NOR2_X1 U868 ( .A1(n1208), .A2(n1209), .ZN(n1206) );
NOR2_X1 U869 ( .A1(n1210), .A2(n1098), .ZN(n1209) );
XNOR2_X1 U870 ( .A(n1096), .B(KEYINPUT55), .ZN(n1210) );
NOR2_X1 U871 ( .A1(n1099), .A2(n1211), .ZN(n1208) );
XNOR2_X1 U872 ( .A(KEYINPUT30), .B(n1073), .ZN(n1211) );
NOR3_X1 U873 ( .A1(n1212), .A2(n1073), .A3(n1065), .ZN(n1204) );
INV_X1 U874 ( .A(n1101), .ZN(n1065) );
INV_X1 U875 ( .A(n1213), .ZN(n1200) );
NOR2_X1 U876 ( .A1(n1214), .A2(n1215), .ZN(n1199) );
INV_X1 U877 ( .A(KEYINPUT59), .ZN(n1214) );
NOR2_X1 U878 ( .A1(KEYINPUT59), .A2(n1216), .ZN(n1198) );
NAND4_X1 U879 ( .A1(n1217), .A2(n1054), .A3(n1218), .A4(n1068), .ZN(n1216) );
INV_X1 U880 ( .A(n1149), .ZN(n1193) );
NAND4_X1 U881 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1149) );
NOR4_X1 U882 ( .A1(n1223), .A2(n1166), .A3(n1224), .A4(n1225), .ZN(n1222) );
AND3_X1 U883 ( .A1(n1226), .A2(n1058), .A3(n1227), .ZN(n1166) );
NAND2_X1 U884 ( .A1(n1227), .A2(n1228), .ZN(n1221) );
NAND2_X1 U885 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NAND2_X1 U886 ( .A1(n1231), .A2(n1080), .ZN(n1230) );
XNOR2_X1 U887 ( .A(n1101), .B(KEYINPUT56), .ZN(n1231) );
NAND2_X1 U888 ( .A1(n1056), .A2(n1058), .ZN(n1229) );
NAND3_X1 U889 ( .A1(n1232), .A2(n1057), .A3(n1089), .ZN(n1219) );
NAND2_X1 U890 ( .A1(n1233), .A2(n1234), .ZN(n1190) );
NAND2_X1 U891 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NAND2_X1 U892 ( .A1(G224), .A2(n1093), .ZN(n1236) );
INV_X1 U893 ( .A(n1237), .ZN(n1233) );
NOR2_X1 U894 ( .A1(n1093), .A2(G952), .ZN(n1152) );
XNOR2_X1 U895 ( .A(n1215), .B(n1238), .ZN(G48) );
NOR2_X1 U896 ( .A1(KEYINPUT12), .A2(n1239), .ZN(n1238) );
INV_X1 U897 ( .A(G146), .ZN(n1239) );
NAND2_X1 U898 ( .A1(n1217), .A2(n1240), .ZN(n1215) );
NOR3_X1 U899 ( .A1(n1098), .A2(n1241), .A3(n1212), .ZN(n1217) );
XNOR2_X1 U900 ( .A(G143), .B(n1213), .ZN(G45) );
NAND4_X1 U901 ( .A1(n1240), .A2(n1232), .A3(n1080), .A4(n1059), .ZN(n1213) );
XNOR2_X1 U902 ( .A(G140), .B(n1196), .ZN(G42) );
NAND3_X1 U903 ( .A1(n1242), .A2(n1096), .A3(n1240), .ZN(n1196) );
NAND2_X1 U904 ( .A1(n1243), .A2(n1244), .ZN(G39) );
NAND4_X1 U905 ( .A1(n1245), .A2(n1096), .A3(n1246), .A4(n1247), .ZN(n1244) );
NAND2_X1 U906 ( .A1(KEYINPUT44), .A2(n1129), .ZN(n1247) );
NAND2_X1 U907 ( .A1(KEYINPUT4), .A2(G137), .ZN(n1246) );
NAND3_X1 U908 ( .A1(G137), .A2(n1248), .A3(KEYINPUT4), .ZN(n1243) );
NAND3_X1 U909 ( .A1(n1096), .A2(n1249), .A3(n1245), .ZN(n1248) );
XOR2_X1 U910 ( .A(n1250), .B(KEYINPUT14), .Z(n1245) );
NAND3_X1 U911 ( .A1(n1101), .A2(n1251), .A3(n1240), .ZN(n1250) );
XNOR2_X1 U912 ( .A(KEYINPUT11), .B(n1212), .ZN(n1251) );
INV_X1 U913 ( .A(n1252), .ZN(n1212) );
INV_X1 U914 ( .A(KEYINPUT44), .ZN(n1249) );
XOR2_X1 U915 ( .A(G134), .B(n1253), .Z(G36) );
NOR2_X1 U916 ( .A1(n1099), .A2(n1254), .ZN(n1253) );
INV_X1 U917 ( .A(n1056), .ZN(n1099) );
XNOR2_X1 U918 ( .A(n1255), .B(n1256), .ZN(G33) );
NOR2_X1 U919 ( .A1(n1098), .A2(n1254), .ZN(n1256) );
NAND3_X1 U920 ( .A1(n1080), .A2(n1096), .A3(n1240), .ZN(n1254) );
INV_X1 U921 ( .A(n1073), .ZN(n1096) );
NAND2_X1 U922 ( .A1(n1257), .A2(n1085), .ZN(n1073) );
INV_X1 U923 ( .A(n1087), .ZN(n1257) );
XNOR2_X1 U924 ( .A(G128), .B(n1194), .ZN(G30) );
NAND4_X1 U925 ( .A1(n1240), .A2(n1252), .A3(n1056), .A4(n1059), .ZN(n1194) );
INV_X1 U926 ( .A(n1203), .ZN(n1240) );
NAND2_X1 U927 ( .A1(n1054), .A2(n1258), .ZN(n1203) );
NAND2_X1 U928 ( .A1(n1218), .A2(n1068), .ZN(n1258) );
XOR2_X1 U929 ( .A(n1259), .B(n1260), .Z(G3) );
NOR2_X1 U930 ( .A1(n1207), .A2(n1261), .ZN(n1260) );
NOR2_X1 U931 ( .A1(KEYINPUT34), .A2(n1262), .ZN(n1259) );
XNOR2_X1 U932 ( .A(G101), .B(KEYINPUT50), .ZN(n1262) );
XNOR2_X1 U933 ( .A(n1132), .B(n1263), .ZN(G27) );
NOR2_X1 U934 ( .A1(KEYINPUT22), .A2(n1195), .ZN(n1263) );
NAND3_X1 U935 ( .A1(n1242), .A2(n1059), .A3(n1264), .ZN(n1195) );
NOR3_X1 U936 ( .A1(n1076), .A2(n1079), .A3(n1265), .ZN(n1264) );
AND2_X1 U937 ( .A1(n1068), .A2(n1218), .ZN(n1265) );
XOR2_X1 U938 ( .A(n1266), .B(KEYINPUT0), .Z(n1218) );
NAND2_X1 U939 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
XOR2_X1 U940 ( .A(KEYINPUT54), .B(G900), .Z(n1268) );
NOR3_X1 U941 ( .A1(n1083), .A2(n1082), .A3(n1098), .ZN(n1242) );
XNOR2_X1 U942 ( .A(G122), .B(n1269), .ZN(G24) );
NAND3_X1 U943 ( .A1(n1270), .A2(n1057), .A3(n1089), .ZN(n1269) );
NOR2_X1 U944 ( .A1(n1086), .A2(n1241), .ZN(n1089) );
NAND3_X1 U945 ( .A1(n1271), .A2(n1084), .A3(n1058), .ZN(n1086) );
AND2_X1 U946 ( .A1(n1082), .A2(n1272), .ZN(n1058) );
XOR2_X1 U947 ( .A(KEYINPUT6), .B(n1232), .Z(n1270) );
AND2_X1 U948 ( .A1(n1273), .A2(n1274), .ZN(n1232) );
XNOR2_X1 U949 ( .A(G119), .B(n1220), .ZN(G21) );
NAND3_X1 U950 ( .A1(n1275), .A2(n1101), .A3(n1252), .ZN(n1220) );
NOR2_X1 U951 ( .A1(n1272), .A2(n1082), .ZN(n1252) );
INV_X1 U952 ( .A(n1083), .ZN(n1272) );
XOR2_X1 U953 ( .A(G116), .B(n1223), .Z(G18) );
AND3_X1 U954 ( .A1(n1275), .A2(n1056), .A3(n1080), .ZN(n1223) );
NOR2_X1 U955 ( .A1(n1274), .A2(n1276), .ZN(n1056) );
XOR2_X1 U956 ( .A(n1225), .B(n1277), .Z(G15) );
XOR2_X1 U957 ( .A(KEYINPUT32), .B(G113), .Z(n1277) );
AND3_X1 U958 ( .A1(n1080), .A2(n1275), .A3(n1226), .ZN(n1225) );
INV_X1 U959 ( .A(n1098), .ZN(n1226) );
NAND2_X1 U960 ( .A1(n1276), .A2(n1274), .ZN(n1098) );
INV_X1 U961 ( .A(n1273), .ZN(n1276) );
AND4_X1 U962 ( .A1(n1059), .A2(n1271), .A3(n1084), .A4(n1057), .ZN(n1275) );
INV_X1 U963 ( .A(n1207), .ZN(n1080) );
NAND2_X1 U964 ( .A1(n1082), .A2(n1083), .ZN(n1207) );
XNOR2_X1 U965 ( .A(n1224), .B(n1278), .ZN(G12) );
NAND2_X1 U966 ( .A1(KEYINPUT29), .A2(G110), .ZN(n1278) );
NOR3_X1 U967 ( .A1(n1083), .A2(n1082), .A3(n1261), .ZN(n1224) );
NAND2_X1 U968 ( .A1(n1227), .A2(n1101), .ZN(n1261) );
NOR2_X1 U969 ( .A1(n1273), .A2(n1274), .ZN(n1101) );
XNOR2_X1 U970 ( .A(n1279), .B(G475), .ZN(n1274) );
NAND2_X1 U971 ( .A1(n1163), .A2(n1165), .ZN(n1279) );
XNOR2_X1 U972 ( .A(n1280), .B(n1281), .ZN(n1163) );
XOR2_X1 U973 ( .A(n1282), .B(n1283), .Z(n1281) );
XOR2_X1 U974 ( .A(n1284), .B(n1285), .Z(n1283) );
NOR3_X1 U975 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1285) );
NOR2_X1 U976 ( .A1(KEYINPUT8), .A2(n1289), .ZN(n1288) );
NOR2_X1 U977 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NOR2_X1 U978 ( .A1(KEYINPUT48), .A2(n1132), .ZN(n1291) );
AND3_X1 U979 ( .A1(n1132), .A2(G140), .A3(KEYINPUT48), .ZN(n1290) );
NOR2_X1 U980 ( .A1(n1292), .A2(n1293), .ZN(n1287) );
INV_X1 U981 ( .A(KEYINPUT8), .ZN(n1293) );
NOR2_X1 U982 ( .A1(n1294), .A2(n1134), .ZN(n1292) );
XNOR2_X1 U983 ( .A(KEYINPUT48), .B(G125), .ZN(n1294) );
NOR2_X1 U984 ( .A1(G140), .A2(n1132), .ZN(n1286) );
NOR2_X1 U985 ( .A1(KEYINPUT3), .A2(n1295), .ZN(n1284) );
XOR2_X1 U986 ( .A(n1296), .B(n1297), .Z(n1295) );
NOR2_X1 U987 ( .A1(KEYINPUT49), .A2(n1298), .ZN(n1297) );
XNOR2_X1 U988 ( .A(n1299), .B(n1255), .ZN(n1296) );
NAND2_X1 U989 ( .A1(G214), .A2(n1300), .ZN(n1299) );
NOR2_X1 U990 ( .A1(G146), .A2(KEYINPUT53), .ZN(n1282) );
XNOR2_X1 U991 ( .A(G104), .B(n1301), .ZN(n1280) );
XOR2_X1 U992 ( .A(G122), .B(G113), .Z(n1301) );
XOR2_X1 U993 ( .A(n1302), .B(n1160), .Z(n1273) );
INV_X1 U994 ( .A(G478), .ZN(n1160) );
OR2_X1 U995 ( .A1(n1159), .A2(G902), .ZN(n1302) );
XNOR2_X1 U996 ( .A(n1303), .B(n1304), .ZN(n1159) );
XOR2_X1 U997 ( .A(G116), .B(n1305), .Z(n1304) );
XOR2_X1 U998 ( .A(G134), .B(G122), .Z(n1305) );
XOR2_X1 U999 ( .A(n1306), .B(n1307), .Z(n1303) );
XOR2_X1 U1000 ( .A(n1308), .B(n1309), .Z(n1307) );
AND3_X1 U1001 ( .A1(G217), .A2(n1093), .A3(G234), .ZN(n1309) );
NOR2_X1 U1002 ( .A1(KEYINPUT18), .A2(n1310), .ZN(n1308) );
XNOR2_X1 U1003 ( .A(G128), .B(G143), .ZN(n1310) );
NAND2_X1 U1004 ( .A1(KEYINPUT31), .A2(n1311), .ZN(n1306) );
INV_X1 U1005 ( .A(G107), .ZN(n1311) );
AND3_X1 U1006 ( .A1(n1059), .A2(n1057), .A3(n1054), .ZN(n1227) );
NOR2_X1 U1007 ( .A1(n1271), .A2(n1079), .ZN(n1054) );
INV_X1 U1008 ( .A(n1084), .ZN(n1079) );
NAND2_X1 U1009 ( .A1(G221), .A2(n1312), .ZN(n1084) );
INV_X1 U1010 ( .A(n1076), .ZN(n1271) );
XNOR2_X1 U1011 ( .A(n1106), .B(n1107), .ZN(n1076) );
XOR2_X1 U1012 ( .A(n1186), .B(KEYINPUT37), .Z(n1107) );
INV_X1 U1013 ( .A(G469), .ZN(n1186) );
NAND2_X1 U1014 ( .A1(n1313), .A2(n1165), .ZN(n1106) );
XOR2_X1 U1015 ( .A(n1183), .B(n1187), .Z(n1313) );
XOR2_X1 U1016 ( .A(n1314), .B(n1315), .Z(n1187) );
XOR2_X1 U1017 ( .A(n1316), .B(n1131), .Z(n1315) );
XNOR2_X1 U1018 ( .A(n1317), .B(G128), .ZN(n1131) );
NAND2_X1 U1019 ( .A1(n1318), .A2(KEYINPUT62), .ZN(n1317) );
XNOR2_X1 U1020 ( .A(G146), .B(n1319), .ZN(n1318) );
NOR2_X1 U1021 ( .A1(G101), .A2(KEYINPUT46), .ZN(n1316) );
XNOR2_X1 U1022 ( .A(G104), .B(G107), .ZN(n1314) );
XNOR2_X1 U1023 ( .A(n1320), .B(n1321), .ZN(n1183) );
XOR2_X1 U1024 ( .A(n1322), .B(n1176), .Z(n1321) );
AND2_X1 U1025 ( .A1(n1093), .A2(G227), .ZN(n1322) );
XNOR2_X1 U1026 ( .A(G110), .B(G140), .ZN(n1320) );
NAND2_X1 U1027 ( .A1(n1323), .A2(n1068), .ZN(n1057) );
NAND3_X1 U1028 ( .A1(n1324), .A2(n1093), .A3(G952), .ZN(n1068) );
NAND2_X1 U1029 ( .A1(n1267), .A2(n1140), .ZN(n1323) );
INV_X1 U1030 ( .A(G898), .ZN(n1140) );
AND3_X1 U1031 ( .A1(G902), .A2(n1324), .A3(G953), .ZN(n1267) );
NAND2_X1 U1032 ( .A1(G237), .A2(G234), .ZN(n1324) );
INV_X1 U1033 ( .A(n1241), .ZN(n1059) );
NAND2_X1 U1034 ( .A1(n1087), .A2(n1085), .ZN(n1241) );
NAND2_X1 U1035 ( .A1(n1325), .A2(G214), .ZN(n1085) );
XOR2_X1 U1036 ( .A(n1326), .B(KEYINPUT23), .Z(n1325) );
XOR2_X1 U1037 ( .A(n1327), .B(n1192), .Z(n1087) );
NAND2_X1 U1038 ( .A1(G210), .A2(n1326), .ZN(n1192) );
OR2_X1 U1039 ( .A1(G902), .A2(G237), .ZN(n1326) );
NAND2_X1 U1040 ( .A1(n1328), .A2(n1165), .ZN(n1327) );
XOR2_X1 U1041 ( .A(n1148), .B(n1329), .Z(n1328) );
NOR2_X1 U1042 ( .A1(n1237), .A2(n1330), .ZN(n1329) );
NOR2_X1 U1043 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XNOR2_X1 U1044 ( .A(n1235), .B(KEYINPUT51), .ZN(n1332) );
NOR2_X1 U1045 ( .A1(G953), .A2(n1139), .ZN(n1331) );
NOR3_X1 U1046 ( .A1(n1235), .A2(G953), .A3(n1139), .ZN(n1237) );
INV_X1 U1047 ( .A(G224), .ZN(n1139) );
XNOR2_X1 U1048 ( .A(n1177), .B(n1132), .ZN(n1235) );
XOR2_X1 U1049 ( .A(n1333), .B(n1334), .Z(n1148) );
XOR2_X1 U1050 ( .A(n1335), .B(n1336), .Z(n1334) );
XNOR2_X1 U1051 ( .A(G122), .B(n1337), .ZN(n1336) );
XOR2_X1 U1052 ( .A(KEYINPUT40), .B(KEYINPUT16), .Z(n1335) );
XNOR2_X1 U1053 ( .A(n1338), .B(n1339), .ZN(n1333) );
XNOR2_X1 U1054 ( .A(n1340), .B(n1341), .ZN(n1338) );
NAND2_X1 U1055 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
NAND2_X1 U1056 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
NAND2_X1 U1057 ( .A1(KEYINPUT36), .A2(n1346), .ZN(n1345) );
OR2_X1 U1058 ( .A1(G101), .A2(KEYINPUT57), .ZN(n1346) );
INV_X1 U1059 ( .A(n1347), .ZN(n1344) );
NAND2_X1 U1060 ( .A1(G101), .A2(n1348), .ZN(n1342) );
NAND2_X1 U1061 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1062 ( .A1(KEYINPUT36), .A2(n1347), .ZN(n1350) );
XNOR2_X1 U1063 ( .A(n1351), .B(n1352), .ZN(n1347) );
NOR2_X1 U1064 ( .A1(KEYINPUT19), .A2(G104), .ZN(n1352) );
XNOR2_X1 U1065 ( .A(G107), .B(KEYINPUT61), .ZN(n1351) );
INV_X1 U1066 ( .A(KEYINPUT57), .ZN(n1349) );
XNOR2_X1 U1067 ( .A(n1353), .B(n1155), .ZN(n1082) );
NAND2_X1 U1068 ( .A1(G217), .A2(n1312), .ZN(n1155) );
NAND2_X1 U1069 ( .A1(G234), .A2(n1165), .ZN(n1312) );
OR2_X1 U1070 ( .A1(n1154), .A2(G902), .ZN(n1353) );
XNOR2_X1 U1071 ( .A(n1354), .B(n1355), .ZN(n1154) );
XOR2_X1 U1072 ( .A(n1356), .B(n1357), .Z(n1355) );
NAND2_X1 U1073 ( .A1(KEYINPUT60), .A2(n1337), .ZN(n1356) );
INV_X1 U1074 ( .A(G119), .ZN(n1337) );
XOR2_X1 U1075 ( .A(n1358), .B(n1359), .Z(n1354) );
NOR2_X1 U1076 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NOR2_X1 U1077 ( .A1(G140), .A2(n1362), .ZN(n1361) );
NOR2_X1 U1078 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
NOR2_X1 U1079 ( .A1(G125), .A2(n1365), .ZN(n1363) );
NOR2_X1 U1080 ( .A1(n1366), .A2(n1132), .ZN(n1360) );
INV_X1 U1081 ( .A(G125), .ZN(n1132) );
NOR2_X1 U1082 ( .A1(n1367), .A2(n1365), .ZN(n1366) );
INV_X1 U1083 ( .A(KEYINPUT39), .ZN(n1365) );
NOR2_X1 U1084 ( .A1(n1134), .A2(n1364), .ZN(n1367) );
INV_X1 U1085 ( .A(KEYINPUT45), .ZN(n1364) );
INV_X1 U1086 ( .A(G140), .ZN(n1134) );
XNOR2_X1 U1087 ( .A(n1368), .B(n1341), .ZN(n1358) );
INV_X1 U1088 ( .A(G110), .ZN(n1341) );
NAND2_X1 U1089 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
NAND2_X1 U1090 ( .A1(n1371), .A2(n1129), .ZN(n1370) );
XOR2_X1 U1091 ( .A(KEYINPUT42), .B(n1372), .Z(n1369) );
NOR2_X1 U1092 ( .A1(n1129), .A2(n1371), .ZN(n1372) );
NAND3_X1 U1093 ( .A1(G234), .A2(n1093), .A3(G221), .ZN(n1371) );
INV_X1 U1094 ( .A(G953), .ZN(n1093) );
INV_X1 U1095 ( .A(G137), .ZN(n1129) );
XOR2_X1 U1096 ( .A(n1373), .B(n1180), .Z(n1083) );
INV_X1 U1097 ( .A(G472), .ZN(n1180) );
NAND2_X1 U1098 ( .A1(n1374), .A2(n1165), .ZN(n1373) );
INV_X1 U1099 ( .A(G902), .ZN(n1165) );
XOR2_X1 U1100 ( .A(n1174), .B(n1375), .Z(n1374) );
XOR2_X1 U1101 ( .A(n1376), .B(n1171), .Z(n1375) );
XNOR2_X1 U1102 ( .A(n1339), .B(n1377), .ZN(n1171) );
XNOR2_X1 U1103 ( .A(G101), .B(n1378), .ZN(n1377) );
NAND2_X1 U1104 ( .A1(KEYINPUT33), .A2(G119), .ZN(n1378) );
XNOR2_X1 U1105 ( .A(G113), .B(n1379), .ZN(n1339) );
XOR2_X1 U1106 ( .A(KEYINPUT20), .B(G116), .Z(n1379) );
NOR2_X1 U1107 ( .A1(KEYINPUT9), .A2(n1380), .ZN(n1376) );
XNOR2_X1 U1108 ( .A(KEYINPUT17), .B(n1178), .ZN(n1380) );
NAND2_X1 U1109 ( .A1(G210), .A2(n1300), .ZN(n1178) );
NOR2_X1 U1110 ( .A1(G953), .A2(G237), .ZN(n1300) );
XOR2_X1 U1111 ( .A(n1177), .B(n1176), .Z(n1174) );
XNOR2_X1 U1112 ( .A(n1255), .B(n1381), .ZN(n1176) );
NOR2_X1 U1113 ( .A1(KEYINPUT52), .A2(n1382), .ZN(n1381) );
XNOR2_X1 U1114 ( .A(n1383), .B(n1384), .ZN(n1382) );
INV_X1 U1115 ( .A(n1130), .ZN(n1384) );
XOR2_X1 U1116 ( .A(G134), .B(KEYINPUT2), .Z(n1130) );
XNOR2_X1 U1117 ( .A(G137), .B(KEYINPUT27), .ZN(n1383) );
INV_X1 U1118 ( .A(G131), .ZN(n1255) );
XNOR2_X1 U1119 ( .A(n1357), .B(n1385), .ZN(n1177) );
XOR2_X1 U1120 ( .A(KEYINPUT26), .B(n1319), .Z(n1385) );
XNOR2_X1 U1121 ( .A(n1298), .B(KEYINPUT10), .ZN(n1319) );
INV_X1 U1122 ( .A(G143), .ZN(n1298) );
XNOR2_X1 U1123 ( .A(G128), .B(G146), .ZN(n1357) );
endmodule


