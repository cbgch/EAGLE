//Key = 0011110110110010101000111011111111010000101101101010101111000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298;

XNOR2_X1 U730 ( .A(G107), .B(n994), .ZN(G9) );
NOR2_X1 U731 ( .A1(n995), .A2(n996), .ZN(G75) );
NOR4_X1 U732 ( .A1(n997), .A2(n998), .A3(n999), .A4(n1000), .ZN(n996) );
NAND3_X1 U733 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n997) );
NAND2_X1 U734 ( .A1(n1004), .A2(n1005), .ZN(n1001) );
NAND2_X1 U735 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NAND2_X1 U736 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND2_X1 U737 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND4_X1 U738 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1011) );
XNOR2_X1 U739 ( .A(n1016), .B(KEYINPUT2), .ZN(n1012) );
NAND3_X1 U740 ( .A1(n1017), .A2(n1018), .A3(n1016), .ZN(n1010) );
OR2_X1 U741 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND2_X1 U742 ( .A1(n1015), .A2(n1021), .ZN(n1006) );
NAND3_X1 U743 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1021) );
NAND3_X1 U744 ( .A1(n1025), .A2(n1026), .A3(n1016), .ZN(n1024) );
XOR2_X1 U745 ( .A(KEYINPUT1), .B(n1008), .Z(n1026) );
NAND2_X1 U746 ( .A1(n1017), .A2(n1027), .ZN(n1023) );
NAND2_X1 U747 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U748 ( .A1(n1016), .A2(n1030), .ZN(n1029) );
NAND2_X1 U749 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U750 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U751 ( .A1(n1008), .A2(n1035), .ZN(n1028) );
NAND2_X1 U752 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U753 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
INV_X1 U754 ( .A(KEYINPUT36), .ZN(n1039) );
NAND2_X1 U755 ( .A1(n1040), .A2(n1041), .ZN(n1036) );
NAND4_X1 U756 ( .A1(n1008), .A2(n1038), .A3(KEYINPUT36), .A4(n1042), .ZN(n1022) );
INV_X1 U757 ( .A(n1043), .ZN(n1004) );
AND3_X1 U758 ( .A1(n1003), .A2(n1044), .A3(n1002), .ZN(n995) );
NAND2_X1 U759 ( .A1(n1045), .A2(n1046), .ZN(n1002) );
NOR4_X1 U760 ( .A1(n1041), .A2(n1014), .A3(n1047), .A4(n1048), .ZN(n1046) );
XOR2_X1 U761 ( .A(n1049), .B(n1050), .Z(n1048) );
NAND2_X1 U762 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
XOR2_X1 U763 ( .A(KEYINPUT7), .B(KEYINPUT53), .Z(n1051) );
XNOR2_X1 U764 ( .A(n1053), .B(n1054), .ZN(n1047) );
NAND2_X1 U765 ( .A1(KEYINPUT56), .A2(n1055), .ZN(n1053) );
NOR4_X1 U766 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1045) );
XNOR2_X1 U767 ( .A(n1060), .B(KEYINPUT16), .ZN(n1058) );
XNOR2_X1 U768 ( .A(n1034), .B(KEYINPUT62), .ZN(n1057) );
XOR2_X1 U769 ( .A(n1061), .B(n1062), .Z(n1056) );
NOR2_X1 U770 ( .A1(G902), .A2(n1063), .ZN(n1062) );
XNOR2_X1 U771 ( .A(G475), .B(KEYINPUT40), .ZN(n1061) );
XOR2_X1 U772 ( .A(n1064), .B(n1065), .Z(G72) );
XOR2_X1 U773 ( .A(n1066), .B(n1067), .Z(n1065) );
NOR2_X1 U774 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
AND2_X1 U775 ( .A1(G227), .A2(G900), .ZN(n1068) );
NAND2_X1 U776 ( .A1(n1070), .A2(n1071), .ZN(n1066) );
NAND2_X1 U777 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XNOR2_X1 U778 ( .A(G953), .B(KEYINPUT50), .ZN(n1072) );
XOR2_X1 U779 ( .A(n1074), .B(n1075), .Z(n1070) );
NOR3_X1 U780 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NOR2_X1 U781 ( .A1(KEYINPUT33), .A2(n1079), .ZN(n1078) );
NOR3_X1 U782 ( .A1(n1080), .A2(G125), .A3(n1081), .ZN(n1077) );
INV_X1 U783 ( .A(KEYINPUT33), .ZN(n1080) );
AND2_X1 U784 ( .A1(n1081), .A2(G125), .ZN(n1076) );
NAND2_X1 U785 ( .A1(KEYINPUT42), .A2(n1079), .ZN(n1081) );
NAND3_X1 U786 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1074) );
NAND2_X1 U787 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U788 ( .A1(KEYINPUT63), .A2(n1087), .ZN(n1083) );
NAND2_X1 U789 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XNOR2_X1 U790 ( .A(KEYINPUT48), .B(n1090), .ZN(n1089) );
NAND2_X1 U791 ( .A1(n1091), .A2(n1092), .ZN(n1082) );
INV_X1 U792 ( .A(KEYINPUT63), .ZN(n1092) );
NAND2_X1 U793 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NAND3_X1 U794 ( .A1(KEYINPUT48), .A2(n1088), .A3(n1090), .ZN(n1094) );
OR2_X1 U795 ( .A1(n1090), .A2(KEYINPUT48), .ZN(n1093) );
INV_X1 U796 ( .A(n1085), .ZN(n1090) );
NAND2_X1 U797 ( .A1(n1069), .A2(n1095), .ZN(n1064) );
NAND2_X1 U798 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
INV_X1 U799 ( .A(n999), .ZN(n1096) );
XOR2_X1 U800 ( .A(n1098), .B(n1099), .Z(G69) );
NAND2_X1 U801 ( .A1(KEYINPUT28), .A2(n1100), .ZN(n1099) );
NAND2_X1 U802 ( .A1(G953), .A2(n1101), .ZN(n1100) );
NAND2_X1 U803 ( .A1(G898), .A2(n1102), .ZN(n1101) );
XOR2_X1 U804 ( .A(KEYINPUT37), .B(G224), .Z(n1102) );
NAND2_X1 U805 ( .A1(n1103), .A2(n1104), .ZN(n1098) );
NAND2_X1 U806 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U807 ( .A1(n1107), .A2(n998), .ZN(n1106) );
XOR2_X1 U808 ( .A(n1108), .B(KEYINPUT10), .Z(n1105) );
XOR2_X1 U809 ( .A(n1109), .B(KEYINPUT25), .Z(n1103) );
NAND3_X1 U810 ( .A1(n1108), .A2(n998), .A3(n1107), .ZN(n1109) );
XNOR2_X1 U811 ( .A(KEYINPUT60), .B(G953), .ZN(n1107) );
NAND2_X1 U812 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NAND2_X1 U813 ( .A1(G953), .A2(n1112), .ZN(n1111) );
XOR2_X1 U814 ( .A(n1113), .B(KEYINPUT35), .Z(n1110) );
NAND2_X1 U815 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XNOR2_X1 U816 ( .A(KEYINPUT55), .B(n1116), .ZN(n1114) );
NOR3_X1 U817 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(G66) );
AND2_X1 U818 ( .A1(KEYINPUT18), .A2(n1120), .ZN(n1119) );
NOR3_X1 U819 ( .A1(KEYINPUT18), .A2(n1069), .A3(n1044), .ZN(n1118) );
XNOR2_X1 U820 ( .A(n1121), .B(n1122), .ZN(n1117) );
NOR2_X1 U821 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U822 ( .A1(n1120), .A2(n1125), .ZN(G63) );
XOR2_X1 U823 ( .A(n1126), .B(n1127), .Z(n1125) );
AND2_X1 U824 ( .A1(G478), .A2(n1128), .ZN(n1126) );
NOR2_X1 U825 ( .A1(n1120), .A2(n1129), .ZN(G60) );
XOR2_X1 U826 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U827 ( .A1(KEYINPUT58), .A2(n1063), .ZN(n1131) );
NAND2_X1 U828 ( .A1(n1128), .A2(G475), .ZN(n1130) );
XOR2_X1 U829 ( .A(n1132), .B(G104), .Z(G6) );
NAND2_X1 U830 ( .A1(KEYINPUT23), .A2(n1133), .ZN(n1132) );
NOR3_X1 U831 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(G57) );
NOR3_X1 U832 ( .A1(n1137), .A2(n1069), .A3(n1044), .ZN(n1136) );
INV_X1 U833 ( .A(G952), .ZN(n1044) );
AND2_X1 U834 ( .A1(n1137), .A2(n1120), .ZN(n1135) );
INV_X1 U835 ( .A(KEYINPUT21), .ZN(n1137) );
XOR2_X1 U836 ( .A(n1138), .B(n1139), .Z(n1134) );
XOR2_X1 U837 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U838 ( .A(n1142), .B(n1143), .Z(n1138) );
AND2_X1 U839 ( .A1(G472), .A2(n1128), .ZN(n1143) );
NAND2_X1 U840 ( .A1(KEYINPUT43), .A2(n1144), .ZN(n1142) );
XNOR2_X1 U841 ( .A(G101), .B(n1145), .ZN(n1144) );
NOR2_X1 U842 ( .A1(n1120), .A2(n1146), .ZN(G54) );
XOR2_X1 U843 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U844 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U845 ( .A1(n1054), .A2(n1124), .ZN(n1150) );
INV_X1 U846 ( .A(G469), .ZN(n1054) );
NOR2_X1 U847 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
XOR2_X1 U848 ( .A(n1153), .B(n1154), .Z(n1152) );
XNOR2_X1 U849 ( .A(n1155), .B(KEYINPUT0), .ZN(n1154) );
XNOR2_X1 U850 ( .A(KEYINPUT17), .B(KEYINPUT14), .ZN(n1151) );
NOR2_X1 U851 ( .A1(n1120), .A2(n1156), .ZN(G51) );
XOR2_X1 U852 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U853 ( .A1(KEYINPUT47), .A2(n1159), .ZN(n1158) );
XOR2_X1 U854 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U855 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
AND3_X1 U856 ( .A1(KEYINPUT51), .A2(n1164), .A3(G125), .ZN(n1163) );
NOR2_X1 U857 ( .A1(KEYINPUT51), .A2(n1165), .ZN(n1162) );
XNOR2_X1 U858 ( .A(G125), .B(n1164), .ZN(n1165) );
XOR2_X1 U859 ( .A(n1166), .B(n1167), .Z(n1160) );
NOR2_X1 U860 ( .A1(n1168), .A2(KEYINPUT39), .ZN(n1167) );
NAND2_X1 U861 ( .A1(n1128), .A2(n1050), .ZN(n1157) );
INV_X1 U862 ( .A(n1124), .ZN(n1128) );
NAND2_X1 U863 ( .A1(G902), .A2(n1169), .ZN(n1124) );
OR3_X1 U864 ( .A1(n1000), .A2(n999), .A3(n998), .ZN(n1169) );
NAND4_X1 U865 ( .A1(n1170), .A2(n1171), .A3(n994), .A4(n1172), .ZN(n998) );
NOR3_X1 U866 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1172) );
INV_X1 U867 ( .A(n1133), .ZN(n1175) );
NAND3_X1 U868 ( .A1(n1176), .A2(n1008), .A3(n1019), .ZN(n1133) );
NOR2_X1 U869 ( .A1(n1177), .A2(n1178), .ZN(n1173) );
NOR3_X1 U870 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1177) );
NOR2_X1 U871 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
INV_X1 U872 ( .A(n1184), .ZN(n1180) );
NOR2_X1 U873 ( .A1(n1185), .A2(n1031), .ZN(n1179) );
NAND3_X1 U874 ( .A1(n1020), .A2(n1008), .A3(n1176), .ZN(n994) );
NAND4_X1 U875 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n999) );
NOR4_X1 U876 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
XNOR2_X1 U877 ( .A(n1097), .B(KEYINPUT34), .ZN(n1000) );
NOR2_X1 U878 ( .A1(n1069), .A2(G952), .ZN(n1120) );
XNOR2_X1 U879 ( .A(G146), .B(n1188), .ZN(G48) );
NAND3_X1 U880 ( .A1(n1194), .A2(n1019), .A3(n1195), .ZN(n1188) );
XNOR2_X1 U881 ( .A(G143), .B(n1186), .ZN(G45) );
NAND4_X1 U882 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1059), .ZN(n1186) );
XNOR2_X1 U883 ( .A(G140), .B(n1097), .ZN(G42) );
NAND2_X1 U884 ( .A1(n1198), .A2(n1199), .ZN(n1097) );
XNOR2_X1 U885 ( .A(G137), .B(n1187), .ZN(G39) );
NAND3_X1 U886 ( .A1(n1194), .A2(n1015), .A3(n1198), .ZN(n1187) );
XOR2_X1 U887 ( .A(G134), .B(n1193), .Z(G36) );
AND3_X1 U888 ( .A1(n1196), .A2(n1020), .A3(n1198), .ZN(n1193) );
NAND2_X1 U889 ( .A1(n1200), .A2(n1201), .ZN(G33) );
NAND2_X1 U890 ( .A1(n1192), .A2(n1202), .ZN(n1201) );
XOR2_X1 U891 ( .A(KEYINPUT52), .B(n1203), .Z(n1200) );
NOR2_X1 U892 ( .A1(n1192), .A2(n1202), .ZN(n1203) );
AND3_X1 U893 ( .A1(n1196), .A2(n1019), .A3(n1198), .ZN(n1192) );
AND3_X1 U894 ( .A1(n1025), .A2(n1204), .A3(n1016), .ZN(n1198) );
AND2_X1 U895 ( .A1(n1205), .A2(n1040), .ZN(n1016) );
XNOR2_X1 U896 ( .A(KEYINPUT49), .B(n1041), .ZN(n1205) );
XOR2_X1 U897 ( .A(G128), .B(n1191), .Z(G30) );
AND3_X1 U898 ( .A1(n1194), .A2(n1020), .A3(n1195), .ZN(n1191) );
AND3_X1 U899 ( .A1(n1038), .A2(n1204), .A3(n1025), .ZN(n1195) );
XOR2_X1 U900 ( .A(n1206), .B(n1174), .Z(G3) );
AND3_X1 U901 ( .A1(n1015), .A2(n1176), .A3(n1196), .ZN(n1174) );
XNOR2_X1 U902 ( .A(G101), .B(KEYINPUT22), .ZN(n1206) );
XOR2_X1 U903 ( .A(G125), .B(n1190), .Z(G27) );
AND4_X1 U904 ( .A1(n1199), .A2(n1017), .A3(n1038), .A4(n1204), .ZN(n1190) );
NAND2_X1 U905 ( .A1(n1043), .A2(n1207), .ZN(n1204) );
NAND4_X1 U906 ( .A1(G953), .A2(G902), .A3(n1208), .A4(n1073), .ZN(n1207) );
INV_X1 U907 ( .A(G900), .ZN(n1073) );
AND3_X1 U908 ( .A1(n1033), .A2(n1034), .A3(n1019), .ZN(n1199) );
XOR2_X1 U909 ( .A(n1209), .B(n1210), .Z(G24) );
NOR2_X1 U910 ( .A1(KEYINPUT38), .A2(n1211), .ZN(n1210) );
NOR3_X1 U911 ( .A1(n1184), .A2(n1212), .A3(n1213), .ZN(n1209) );
NOR2_X1 U912 ( .A1(KEYINPUT5), .A2(n1214), .ZN(n1213) );
NOR3_X1 U913 ( .A1(n1042), .A2(n1038), .A3(n1215), .ZN(n1214) );
INV_X1 U914 ( .A(n1216), .ZN(n1215) );
AND2_X1 U915 ( .A1(n1178), .A2(KEYINPUT5), .ZN(n1212) );
NAND3_X1 U916 ( .A1(n1008), .A2(n1059), .A3(n1197), .ZN(n1184) );
NOR2_X1 U917 ( .A1(n1034), .A2(n1060), .ZN(n1008) );
XOR2_X1 U918 ( .A(G119), .B(n1217), .Z(G21) );
NOR3_X1 U919 ( .A1(n1178), .A2(n1218), .A3(n1182), .ZN(n1217) );
INV_X1 U920 ( .A(n1015), .ZN(n1182) );
XNOR2_X1 U921 ( .A(n1194), .B(KEYINPUT41), .ZN(n1218) );
INV_X1 U922 ( .A(n1183), .ZN(n1194) );
NAND2_X1 U923 ( .A1(n1060), .A2(n1034), .ZN(n1183) );
XOR2_X1 U924 ( .A(G116), .B(n1219), .Z(G18) );
NOR4_X1 U925 ( .A1(n1185), .A2(n1178), .A3(n1031), .A4(n1220), .ZN(n1219) );
XOR2_X1 U926 ( .A(KEYINPUT61), .B(KEYINPUT32), .Z(n1220) );
INV_X1 U927 ( .A(n1196), .ZN(n1031) );
INV_X1 U928 ( .A(n1020), .ZN(n1185) );
NOR2_X1 U929 ( .A1(n1197), .A2(n1221), .ZN(n1020) );
INV_X1 U930 ( .A(n1059), .ZN(n1221) );
XNOR2_X1 U931 ( .A(G113), .B(n1170), .ZN(G15) );
NAND3_X1 U932 ( .A1(n1019), .A2(n1222), .A3(n1196), .ZN(n1170) );
NOR2_X1 U933 ( .A1(n1034), .A2(n1033), .ZN(n1196) );
INV_X1 U934 ( .A(n1178), .ZN(n1222) );
NAND3_X1 U935 ( .A1(n1038), .A2(n1216), .A3(n1017), .ZN(n1178) );
INV_X1 U936 ( .A(n1042), .ZN(n1017) );
NAND2_X1 U937 ( .A1(n1013), .A2(n1223), .ZN(n1042) );
XOR2_X1 U938 ( .A(KEYINPUT11), .B(n1014), .Z(n1223) );
NOR2_X1 U939 ( .A1(n1224), .A2(n1059), .ZN(n1019) );
XNOR2_X1 U940 ( .A(G110), .B(n1225), .ZN(G12) );
NAND2_X1 U941 ( .A1(KEYINPUT4), .A2(n1226), .ZN(n1225) );
INV_X1 U942 ( .A(n1171), .ZN(n1226) );
NAND4_X1 U943 ( .A1(n1015), .A2(n1176), .A3(n1033), .A4(n1034), .ZN(n1171) );
XOR2_X1 U944 ( .A(n1227), .B(n1123), .Z(n1034) );
NAND2_X1 U945 ( .A1(G217), .A2(n1228), .ZN(n1123) );
NAND2_X1 U946 ( .A1(n1121), .A2(n1229), .ZN(n1227) );
XNOR2_X1 U947 ( .A(n1230), .B(n1231), .ZN(n1121) );
XOR2_X1 U948 ( .A(n1232), .B(n1233), .Z(n1231) );
XNOR2_X1 U949 ( .A(n1234), .B(n1235), .ZN(n1233) );
NAND2_X1 U950 ( .A1(n1236), .A2(G221), .ZN(n1234) );
XOR2_X1 U951 ( .A(n1237), .B(n1238), .Z(n1230) );
XOR2_X1 U952 ( .A(KEYINPUT24), .B(G125), .Z(n1238) );
XOR2_X1 U953 ( .A(n1239), .B(G119), .Z(n1237) );
NAND2_X1 U954 ( .A1(KEYINPUT46), .A2(n1240), .ZN(n1239) );
XOR2_X1 U955 ( .A(KEYINPUT3), .B(G137), .Z(n1240) );
INV_X1 U956 ( .A(n1060), .ZN(n1033) );
XNOR2_X1 U957 ( .A(n1241), .B(G472), .ZN(n1060) );
NAND2_X1 U958 ( .A1(n1242), .A2(n1229), .ZN(n1241) );
XNOR2_X1 U959 ( .A(n1243), .B(n1244), .ZN(n1242) );
INV_X1 U960 ( .A(n1245), .ZN(n1244) );
XNOR2_X1 U961 ( .A(n1140), .B(n1145), .ZN(n1243) );
NAND2_X1 U962 ( .A1(n1246), .A2(G210), .ZN(n1145) );
XOR2_X1 U963 ( .A(n1247), .B(n1155), .Z(n1140) );
XOR2_X1 U964 ( .A(n1085), .B(n1248), .Z(n1155) );
XOR2_X1 U965 ( .A(n1249), .B(KEYINPUT9), .Z(n1247) );
NAND2_X1 U966 ( .A1(KEYINPUT31), .A2(n1250), .ZN(n1249) );
INV_X1 U967 ( .A(G113), .ZN(n1250) );
AND3_X1 U968 ( .A1(n1038), .A2(n1216), .A3(n1025), .ZN(n1176) );
NOR2_X1 U969 ( .A1(n1013), .A2(n1014), .ZN(n1025) );
AND2_X1 U970 ( .A1(G221), .A2(n1228), .ZN(n1014) );
NAND2_X1 U971 ( .A1(G234), .A2(n1229), .ZN(n1228) );
XOR2_X1 U972 ( .A(n1055), .B(G469), .Z(n1013) );
NAND2_X1 U973 ( .A1(n1251), .A2(n1229), .ZN(n1055) );
XOR2_X1 U974 ( .A(n1252), .B(n1253), .Z(n1251) );
XNOR2_X1 U975 ( .A(n1153), .B(n1147), .ZN(n1253) );
XNOR2_X1 U976 ( .A(n1254), .B(n1232), .ZN(n1147) );
XNOR2_X1 U977 ( .A(G110), .B(n1079), .ZN(n1232) );
NAND2_X1 U978 ( .A1(n1255), .A2(n1069), .ZN(n1254) );
XNOR2_X1 U979 ( .A(G227), .B(KEYINPUT30), .ZN(n1255) );
XOR2_X1 U980 ( .A(n1256), .B(n1257), .Z(n1153) );
NOR2_X1 U981 ( .A1(KEYINPUT19), .A2(n1258), .ZN(n1257) );
XNOR2_X1 U982 ( .A(G101), .B(KEYINPUT59), .ZN(n1256) );
XNOR2_X1 U983 ( .A(n1259), .B(n1085), .ZN(n1252) );
XOR2_X1 U984 ( .A(G131), .B(n1260), .Z(n1085) );
XOR2_X1 U985 ( .A(G137), .B(G134), .Z(n1260) );
NAND2_X1 U986 ( .A1(KEYINPUT8), .A2(n1086), .ZN(n1259) );
INV_X1 U987 ( .A(n1088), .ZN(n1086) );
XOR2_X1 U988 ( .A(KEYINPUT0), .B(n1164), .Z(n1088) );
INV_X1 U989 ( .A(n1248), .ZN(n1164) );
NAND2_X1 U990 ( .A1(n1043), .A2(n1261), .ZN(n1216) );
NAND4_X1 U991 ( .A1(G953), .A2(G902), .A3(n1208), .A4(n1112), .ZN(n1261) );
INV_X1 U992 ( .A(G898), .ZN(n1112) );
NAND3_X1 U993 ( .A1(n1003), .A2(n1208), .A3(G952), .ZN(n1043) );
NAND2_X1 U994 ( .A1(G237), .A2(G234), .ZN(n1208) );
XOR2_X1 U995 ( .A(n1069), .B(KEYINPUT13), .Z(n1003) );
NOR2_X1 U996 ( .A1(n1262), .A2(n1040), .ZN(n1038) );
XOR2_X1 U997 ( .A(n1052), .B(n1050), .Z(n1040) );
AND2_X1 U998 ( .A1(G210), .A2(n1263), .ZN(n1050) );
NAND2_X1 U999 ( .A1(n1264), .A2(n1229), .ZN(n1052) );
XOR2_X1 U1000 ( .A(n1168), .B(n1265), .Z(n1264) );
XOR2_X1 U1001 ( .A(n1266), .B(n1166), .Z(n1265) );
NAND2_X1 U1002 ( .A1(n1116), .A2(n1115), .ZN(n1166) );
NAND2_X1 U1003 ( .A1(n1267), .A2(n1268), .ZN(n1115) );
OR2_X1 U1004 ( .A1(n1267), .A2(n1268), .ZN(n1116) );
XNOR2_X1 U1005 ( .A(n1269), .B(n1258), .ZN(n1268) );
XOR2_X1 U1006 ( .A(G104), .B(n1270), .Z(n1258) );
XOR2_X1 U1007 ( .A(KEYINPUT26), .B(G107), .Z(n1270) );
XNOR2_X1 U1008 ( .A(n1245), .B(G113), .ZN(n1269) );
XOR2_X1 U1009 ( .A(G101), .B(n1141), .Z(n1245) );
XOR2_X1 U1010 ( .A(G116), .B(G119), .Z(n1141) );
XOR2_X1 U1011 ( .A(G110), .B(n1271), .Z(n1267) );
NOR2_X1 U1012 ( .A1(KEYINPUT20), .A2(n1211), .ZN(n1271) );
NAND2_X1 U1013 ( .A1(n1272), .A2(KEYINPUT57), .ZN(n1266) );
XNOR2_X1 U1014 ( .A(n1248), .B(G125), .ZN(n1272) );
XOR2_X1 U1015 ( .A(G143), .B(n1235), .Z(n1248) );
XOR2_X1 U1016 ( .A(G128), .B(G146), .Z(n1235) );
AND2_X1 U1017 ( .A1(G224), .A2(n1069), .ZN(n1168) );
XOR2_X1 U1018 ( .A(KEYINPUT49), .B(n1041), .Z(n1262) );
AND2_X1 U1019 ( .A1(G214), .A2(n1263), .ZN(n1041) );
NAND2_X1 U1020 ( .A1(n1229), .A2(n1273), .ZN(n1263) );
INV_X1 U1021 ( .A(G237), .ZN(n1273) );
INV_X1 U1022 ( .A(G902), .ZN(n1229) );
NOR2_X1 U1023 ( .A1(n1059), .A2(n1197), .ZN(n1015) );
INV_X1 U1024 ( .A(n1224), .ZN(n1197) );
XNOR2_X1 U1025 ( .A(n1274), .B(G475), .ZN(n1224) );
NAND2_X1 U1026 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
OR2_X1 U1027 ( .A1(n1063), .A2(G902), .ZN(n1276) );
XOR2_X1 U1028 ( .A(n1277), .B(n1278), .Z(n1063) );
XOR2_X1 U1029 ( .A(G104), .B(n1279), .Z(n1278) );
NOR2_X1 U1030 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
XOR2_X1 U1031 ( .A(n1282), .B(KEYINPUT54), .Z(n1281) );
NAND2_X1 U1032 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NOR2_X1 U1033 ( .A1(n1283), .A2(n1284), .ZN(n1280) );
XOR2_X1 U1034 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U1035 ( .A(G143), .B(n1202), .ZN(n1286) );
INV_X1 U1036 ( .A(G131), .ZN(n1202) );
NAND2_X1 U1037 ( .A1(n1246), .A2(G214), .ZN(n1285) );
NOR2_X1 U1038 ( .A1(G953), .A2(G237), .ZN(n1246) );
XOR2_X1 U1039 ( .A(n1287), .B(n1288), .Z(n1283) );
XOR2_X1 U1040 ( .A(KEYINPUT15), .B(G146), .Z(n1288) );
XOR2_X1 U1041 ( .A(G125), .B(n1079), .Z(n1287) );
XNOR2_X1 U1042 ( .A(G140), .B(KEYINPUT12), .ZN(n1079) );
XNOR2_X1 U1043 ( .A(G113), .B(G122), .ZN(n1277) );
XOR2_X1 U1044 ( .A(KEYINPUT6), .B(KEYINPUT45), .Z(n1275) );
XNOR2_X1 U1045 ( .A(n1289), .B(G478), .ZN(n1059) );
OR2_X1 U1046 ( .A1(n1127), .A2(G902), .ZN(n1289) );
XNOR2_X1 U1047 ( .A(n1290), .B(n1291), .ZN(n1127) );
XOR2_X1 U1048 ( .A(G107), .B(n1292), .Z(n1291) );
XNOR2_X1 U1049 ( .A(n1211), .B(G116), .ZN(n1292) );
INV_X1 U1050 ( .A(G122), .ZN(n1211) );
XOR2_X1 U1051 ( .A(n1293), .B(n1294), .Z(n1290) );
NOR2_X1 U1052 ( .A1(KEYINPUT44), .A2(n1295), .ZN(n1294) );
XOR2_X1 U1053 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U1054 ( .A(KEYINPUT27), .B(G134), .Z(n1297) );
NAND2_X1 U1055 ( .A1(KEYINPUT29), .A2(n1298), .ZN(n1296) );
XOR2_X1 U1056 ( .A(G143), .B(G128), .Z(n1298) );
NAND2_X1 U1057 ( .A1(G217), .A2(n1236), .ZN(n1293) );
AND2_X1 U1058 ( .A1(G234), .A2(n1069), .ZN(n1236) );
INV_X1 U1059 ( .A(G953), .ZN(n1069) );
endmodule


