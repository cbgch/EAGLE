//Key = 1001100111000100101011001000100100010111011101010101010110111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376;

XNOR2_X1 U750 ( .A(G107), .B(n1045), .ZN(G9) );
NAND2_X1 U751 ( .A1(KEYINPUT35), .A2(n1046), .ZN(n1045) );
INV_X1 U752 ( .A(n1047), .ZN(n1046) );
NOR2_X1 U753 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR4_X1 U754 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1049) );
NAND3_X1 U755 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1050) );
NAND2_X1 U756 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND4_X1 U758 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1060) );
NAND2_X1 U759 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U760 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND3_X1 U761 ( .A1(n1069), .A2(n1070), .A3(n1068), .ZN(n1059) );
NAND2_X1 U762 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NAND3_X1 U763 ( .A1(n1063), .A2(n1073), .A3(n1062), .ZN(n1072) );
NAND2_X1 U764 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U765 ( .A1(n1061), .A2(n1076), .ZN(n1071) );
NAND2_X1 U766 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U767 ( .A1(n1063), .A2(n1079), .ZN(n1078) );
NAND2_X1 U768 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U769 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U770 ( .A1(n1062), .A2(n1084), .ZN(n1077) );
NAND2_X1 U771 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
INV_X1 U772 ( .A(n1087), .ZN(n1057) );
NOR3_X1 U773 ( .A1(n1088), .A2(G953), .A3(n1089), .ZN(n1048) );
INV_X1 U774 ( .A(n1054), .ZN(n1089) );
NAND4_X1 U775 ( .A1(n1063), .A2(n1070), .A3(n1062), .A4(n1090), .ZN(n1054) );
NOR4_X1 U776 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1090) );
XNOR2_X1 U777 ( .A(n1095), .B(n1096), .ZN(n1094) );
NOR2_X1 U778 ( .A1(KEYINPUT17), .A2(n1097), .ZN(n1095) );
XOR2_X1 U779 ( .A(KEYINPUT53), .B(n1098), .Z(n1097) );
XOR2_X1 U780 ( .A(KEYINPUT58), .B(n1099), .Z(n1093) );
NOR2_X1 U781 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U782 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XNOR2_X1 U783 ( .A(KEYINPUT42), .B(n1104), .ZN(n1103) );
XNOR2_X1 U784 ( .A(G475), .B(KEYINPUT45), .ZN(n1102) );
NOR2_X1 U785 ( .A1(n1105), .A2(n1106), .ZN(n1100) );
XNOR2_X1 U786 ( .A(G475), .B(KEYINPUT14), .ZN(n1106) );
XOR2_X1 U787 ( .A(n1104), .B(KEYINPUT42), .Z(n1105) );
AND2_X1 U788 ( .A1(n1107), .A2(KEYINPUT9), .ZN(n1092) );
NOR2_X1 U789 ( .A1(KEYINPUT9), .A2(n1108), .ZN(n1091) );
NOR2_X1 U790 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
INV_X1 U791 ( .A(G478), .ZN(n1110) );
AND2_X1 U792 ( .A1(n1111), .A2(n1112), .ZN(n1109) );
XOR2_X1 U793 ( .A(n1052), .B(KEYINPUT59), .Z(n1088) );
INV_X1 U794 ( .A(G952), .ZN(n1052) );
XOR2_X1 U795 ( .A(n1113), .B(n1114), .Z(G72) );
XOR2_X1 U796 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U797 ( .A1(n1117), .A2(n1055), .ZN(n1116) );
AND2_X1 U798 ( .A1(G227), .A2(G900), .ZN(n1117) );
NAND2_X1 U799 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
NAND2_X1 U800 ( .A1(G953), .A2(n1120), .ZN(n1119) );
XOR2_X1 U801 ( .A(n1121), .B(n1122), .Z(n1118) );
XOR2_X1 U802 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U803 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND2_X1 U804 ( .A1(KEYINPUT3), .A2(n1127), .ZN(n1126) );
XOR2_X1 U805 ( .A(G134), .B(n1128), .Z(n1121) );
XOR2_X1 U806 ( .A(KEYINPUT51), .B(G137), .Z(n1128) );
NAND2_X1 U807 ( .A1(n1055), .A2(n1053), .ZN(n1113) );
XOR2_X1 U808 ( .A(n1129), .B(n1130), .Z(G69) );
XOR2_X1 U809 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U810 ( .A1(n1133), .A2(n1055), .ZN(n1132) );
NOR2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND2_X1 U812 ( .A1(n1136), .A2(n1137), .ZN(n1131) );
NAND2_X1 U813 ( .A1(G953), .A2(n1135), .ZN(n1137) );
XNOR2_X1 U814 ( .A(n1138), .B(n1139), .ZN(n1136) );
NOR2_X1 U815 ( .A1(KEYINPUT29), .A2(n1140), .ZN(n1139) );
NAND2_X1 U816 ( .A1(n1055), .A2(n1051), .ZN(n1129) );
NOR2_X1 U817 ( .A1(n1141), .A2(n1142), .ZN(G66) );
XOR2_X1 U818 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U819 ( .A1(n1145), .A2(n1146), .ZN(n1143) );
NOR2_X1 U820 ( .A1(n1141), .A2(n1147), .ZN(G63) );
XOR2_X1 U821 ( .A(n1148), .B(n1112), .Z(n1147) );
NAND2_X1 U822 ( .A1(n1145), .A2(G478), .ZN(n1148) );
NOR2_X1 U823 ( .A1(n1141), .A2(n1149), .ZN(G60) );
XOR2_X1 U824 ( .A(n1150), .B(n1151), .Z(n1149) );
XNOR2_X1 U825 ( .A(n1152), .B(n1153), .ZN(n1151) );
NAND2_X1 U826 ( .A1(n1145), .A2(G475), .ZN(n1152) );
XNOR2_X1 U827 ( .A(KEYINPUT30), .B(KEYINPUT23), .ZN(n1150) );
XOR2_X1 U828 ( .A(G104), .B(n1154), .Z(G6) );
NOR3_X1 U829 ( .A1(n1074), .A2(n1155), .A3(n1156), .ZN(n1154) );
XNOR2_X1 U830 ( .A(n1063), .B(KEYINPUT6), .ZN(n1155) );
NOR2_X1 U831 ( .A1(n1141), .A2(n1157), .ZN(G57) );
NOR2_X1 U832 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U833 ( .A(KEYINPUT44), .B(n1160), .Z(n1159) );
NOR2_X1 U834 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
AND2_X1 U835 ( .A1(n1162), .A2(n1161), .ZN(n1158) );
AND3_X1 U836 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1161) );
NAND3_X1 U837 ( .A1(KEYINPUT49), .A2(n1166), .A3(n1167), .ZN(n1164) );
OR2_X1 U838 ( .A1(n1167), .A2(KEYINPUT49), .ZN(n1163) );
XNOR2_X1 U839 ( .A(n1168), .B(n1169), .ZN(n1162) );
XOR2_X1 U840 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U841 ( .A1(n1172), .A2(KEYINPUT4), .ZN(n1170) );
XOR2_X1 U842 ( .A(n1173), .B(KEYINPUT24), .Z(n1172) );
XOR2_X1 U843 ( .A(n1174), .B(n1175), .Z(n1168) );
NAND2_X1 U844 ( .A1(n1145), .A2(G472), .ZN(n1174) );
NOR3_X1 U845 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(G54) );
NOR3_X1 U846 ( .A1(n1179), .A2(G953), .A3(G952), .ZN(n1178) );
AND2_X1 U847 ( .A1(n1179), .A2(n1141), .ZN(n1177) );
INV_X1 U848 ( .A(KEYINPUT1), .ZN(n1179) );
XOR2_X1 U849 ( .A(n1180), .B(n1181), .Z(n1176) );
XOR2_X1 U850 ( .A(n1182), .B(n1183), .Z(n1181) );
NAND3_X1 U851 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1182) );
NAND2_X1 U852 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
INV_X1 U853 ( .A(KEYINPUT61), .ZN(n1188) );
NAND3_X1 U854 ( .A1(KEYINPUT61), .A2(n1189), .A3(n1173), .ZN(n1185) );
OR2_X1 U855 ( .A1(n1173), .A2(n1189), .ZN(n1184) );
NOR2_X1 U856 ( .A1(KEYINPUT15), .A2(n1187), .ZN(n1189) );
XOR2_X1 U857 ( .A(n1190), .B(n1191), .Z(n1180) );
XOR2_X1 U858 ( .A(n1192), .B(n1175), .Z(n1191) );
NAND2_X1 U859 ( .A1(n1145), .A2(G469), .ZN(n1190) );
NOR2_X1 U860 ( .A1(n1141), .A2(n1193), .ZN(G51) );
XOR2_X1 U861 ( .A(n1194), .B(n1123), .Z(n1193) );
XOR2_X1 U862 ( .A(G125), .B(n1195), .Z(n1123) );
INV_X1 U863 ( .A(n1173), .ZN(n1195) );
XOR2_X1 U864 ( .A(n1196), .B(n1197), .Z(n1194) );
NAND2_X1 U865 ( .A1(n1145), .A2(n1098), .ZN(n1196) );
AND2_X1 U866 ( .A1(G902), .A2(n1198), .ZN(n1145) );
OR2_X1 U867 ( .A1(n1051), .A2(n1053), .ZN(n1198) );
NAND4_X1 U868 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1053) );
NOR4_X1 U869 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
INV_X1 U870 ( .A(n1207), .ZN(n1206) );
NOR2_X1 U871 ( .A1(n1208), .A2(n1209), .ZN(n1201) );
NOR3_X1 U872 ( .A1(n1210), .A2(n1075), .A3(n1211), .ZN(n1209) );
NAND4_X1 U873 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1051) );
AND4_X1 U874 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1047), .ZN(n1215) );
NAND3_X1 U875 ( .A1(n1219), .A2(n1063), .A3(n1220), .ZN(n1047) );
NAND2_X1 U876 ( .A1(n1221), .A2(n1222), .ZN(n1214) );
NAND3_X1 U877 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1222) );
NAND3_X1 U878 ( .A1(n1061), .A2(n1220), .A3(KEYINPUT13), .ZN(n1225) );
NAND3_X1 U879 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1224) );
NAND2_X1 U880 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
OR3_X1 U881 ( .A1(n1080), .A2(KEYINPUT13), .A3(n1231), .ZN(n1230) );
NAND3_X1 U882 ( .A1(n1232), .A2(n1062), .A3(KEYINPUT57), .ZN(n1229) );
NAND3_X1 U883 ( .A1(n1233), .A2(n1234), .A3(n1232), .ZN(n1223) );
INV_X1 U884 ( .A(KEYINPUT57), .ZN(n1234) );
NAND3_X1 U885 ( .A1(n1220), .A2(n1063), .A3(n1232), .ZN(n1212) );
NOR2_X1 U886 ( .A1(n1055), .A2(G952), .ZN(n1141) );
XOR2_X1 U887 ( .A(G146), .B(n1208), .Z(G48) );
NOR3_X1 U888 ( .A1(n1074), .A2(n1211), .A3(n1210), .ZN(n1208) );
XNOR2_X1 U889 ( .A(G143), .B(n1199), .ZN(G45) );
NAND4_X1 U890 ( .A1(n1235), .A2(n1221), .A3(n1236), .A4(n1107), .ZN(n1199) );
XOR2_X1 U891 ( .A(n1205), .B(n1237), .Z(G42) );
NOR2_X1 U892 ( .A1(KEYINPUT48), .A2(n1127), .ZN(n1237) );
AND3_X1 U893 ( .A1(n1232), .A2(n1238), .A3(n1239), .ZN(n1205) );
XOR2_X1 U894 ( .A(G137), .B(n1204), .Z(G39) );
AND3_X1 U895 ( .A1(n1240), .A2(n1061), .A3(n1239), .ZN(n1204) );
NAND3_X1 U896 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(G36) );
NAND2_X1 U897 ( .A1(KEYINPUT2), .A2(G134), .ZN(n1243) );
OR3_X1 U898 ( .A1(G134), .A2(KEYINPUT2), .A3(n1200), .ZN(n1242) );
NAND2_X1 U899 ( .A1(n1244), .A2(n1200), .ZN(n1241) );
NAND3_X1 U900 ( .A1(n1219), .A2(n1221), .A3(n1239), .ZN(n1200) );
NAND2_X1 U901 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
INV_X1 U902 ( .A(KEYINPUT2), .ZN(n1246) );
XOR2_X1 U903 ( .A(n1247), .B(KEYINPUT34), .Z(n1245) );
XOR2_X1 U904 ( .A(G131), .B(n1203), .Z(G33) );
AND3_X1 U905 ( .A1(n1232), .A2(n1221), .A3(n1239), .ZN(n1203) );
NOR4_X1 U906 ( .A1(n1248), .A2(n1080), .A3(n1249), .A4(n1067), .ZN(n1239) );
INV_X1 U907 ( .A(n1070), .ZN(n1067) );
XOR2_X1 U908 ( .A(G128), .B(n1250), .Z(G30) );
NOR3_X1 U909 ( .A1(n1210), .A2(n1251), .A3(n1075), .ZN(n1250) );
INV_X1 U910 ( .A(n1219), .ZN(n1075) );
XOR2_X1 U911 ( .A(n1211), .B(KEYINPUT5), .Z(n1251) );
INV_X1 U912 ( .A(n1235), .ZN(n1210) );
NOR3_X1 U913 ( .A1(n1080), .A2(n1249), .A3(n1065), .ZN(n1235) );
XOR2_X1 U914 ( .A(G101), .B(n1252), .Z(G3) );
NOR3_X1 U915 ( .A1(n1231), .A2(n1085), .A3(n1156), .ZN(n1252) );
INV_X1 U916 ( .A(n1220), .ZN(n1156) );
INV_X1 U917 ( .A(n1221), .ZN(n1085) );
INV_X1 U918 ( .A(n1061), .ZN(n1231) );
XOR2_X1 U919 ( .A(n1253), .B(G125), .Z(G27) );
NAND2_X1 U920 ( .A1(KEYINPUT39), .A2(n1207), .ZN(n1253) );
NAND4_X1 U921 ( .A1(n1232), .A2(n1238), .A3(n1254), .A4(n1062), .ZN(n1207) );
NOR2_X1 U922 ( .A1(n1249), .A2(n1065), .ZN(n1254) );
AND2_X1 U923 ( .A1(n1087), .A2(n1255), .ZN(n1249) );
NAND4_X1 U924 ( .A1(G953), .A2(G902), .A3(n1256), .A4(n1120), .ZN(n1255) );
INV_X1 U925 ( .A(G900), .ZN(n1120) );
XNOR2_X1 U926 ( .A(G122), .B(n1213), .ZN(G24) );
NAND4_X1 U927 ( .A1(n1233), .A2(n1063), .A3(n1236), .A4(n1107), .ZN(n1213) );
XNOR2_X1 U928 ( .A(G119), .B(n1218), .ZN(G21) );
NAND3_X1 U929 ( .A1(n1233), .A2(n1061), .A3(n1240), .ZN(n1218) );
INV_X1 U930 ( .A(n1211), .ZN(n1240) );
NAND2_X1 U931 ( .A1(n1257), .A2(n1258), .ZN(n1211) );
XNOR2_X1 U932 ( .A(G116), .B(n1217), .ZN(G18) );
NAND3_X1 U933 ( .A1(n1219), .A2(n1221), .A3(n1233), .ZN(n1217) );
NOR2_X1 U934 ( .A1(n1236), .A2(n1259), .ZN(n1219) );
XOR2_X1 U935 ( .A(n1260), .B(n1261), .Z(G15) );
NAND3_X1 U936 ( .A1(n1233), .A2(n1221), .A3(n1232), .ZN(n1261) );
INV_X1 U937 ( .A(n1074), .ZN(n1232) );
NAND2_X1 U938 ( .A1(n1259), .A2(n1236), .ZN(n1074) );
NAND2_X1 U939 ( .A1(n1262), .A2(n1263), .ZN(n1221) );
NAND2_X1 U940 ( .A1(n1063), .A2(n1264), .ZN(n1263) );
NOR2_X1 U941 ( .A1(n1258), .A2(n1257), .ZN(n1063) );
INV_X1 U942 ( .A(n1265), .ZN(n1257) );
OR3_X1 U943 ( .A1(n1265), .A2(n1258), .A3(n1264), .ZN(n1262) );
INV_X1 U944 ( .A(KEYINPUT18), .ZN(n1264) );
AND3_X1 U945 ( .A1(n1226), .A2(n1266), .A3(n1062), .ZN(n1233) );
NOR2_X1 U946 ( .A1(n1267), .A2(n1082), .ZN(n1062) );
INV_X1 U947 ( .A(n1083), .ZN(n1267) );
INV_X1 U948 ( .A(n1065), .ZN(n1226) );
XOR2_X1 U949 ( .A(n1216), .B(n1268), .Z(G12) );
NAND2_X1 U950 ( .A1(KEYINPUT63), .A2(G110), .ZN(n1268) );
NAND3_X1 U951 ( .A1(n1238), .A2(n1220), .A3(n1061), .ZN(n1216) );
NOR2_X1 U952 ( .A1(n1107), .A2(n1236), .ZN(n1061) );
XNOR2_X1 U953 ( .A(n1104), .B(G475), .ZN(n1236) );
NAND2_X1 U954 ( .A1(n1111), .A2(n1153), .ZN(n1104) );
NAND3_X1 U955 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1153) );
NAND2_X1 U956 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NAND2_X1 U957 ( .A1(KEYINPUT22), .A2(n1274), .ZN(n1270) );
NAND2_X1 U958 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
XNOR2_X1 U959 ( .A(n1272), .B(KEYINPUT12), .ZN(n1275) );
NAND2_X1 U960 ( .A1(n1277), .A2(n1278), .ZN(n1269) );
INV_X1 U961 ( .A(KEYINPUT22), .ZN(n1278) );
NAND2_X1 U962 ( .A1(n1279), .A2(n1280), .ZN(n1277) );
OR3_X1 U963 ( .A1(n1272), .A2(n1273), .A3(KEYINPUT12), .ZN(n1280) );
INV_X1 U964 ( .A(n1276), .ZN(n1273) );
XOR2_X1 U965 ( .A(n1281), .B(n1282), .Z(n1276) );
XOR2_X1 U966 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U967 ( .A(n1125), .B(n1285), .Z(n1281) );
AND3_X1 U968 ( .A1(G214), .A2(n1055), .A3(n1286), .ZN(n1285) );
NAND2_X1 U969 ( .A1(KEYINPUT12), .A2(n1272), .ZN(n1279) );
XNOR2_X1 U970 ( .A(n1287), .B(G104), .ZN(n1272) );
NAND3_X1 U971 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n1287) );
NAND2_X1 U972 ( .A1(G113), .A2(n1291), .ZN(n1290) );
NAND2_X1 U973 ( .A1(KEYINPUT46), .A2(n1292), .ZN(n1289) );
NAND2_X1 U974 ( .A1(n1293), .A2(n1260), .ZN(n1292) );
XOR2_X1 U975 ( .A(KEYINPUT56), .B(n1291), .Z(n1293) );
NAND2_X1 U976 ( .A1(n1294), .A2(n1295), .ZN(n1288) );
INV_X1 U977 ( .A(KEYINPUT46), .ZN(n1295) );
NAND2_X1 U978 ( .A1(n1296), .A2(n1297), .ZN(n1294) );
OR2_X1 U979 ( .A1(n1298), .A2(KEYINPUT56), .ZN(n1297) );
NAND3_X1 U980 ( .A1(n1298), .A2(n1260), .A3(KEYINPUT56), .ZN(n1296) );
INV_X1 U981 ( .A(n1259), .ZN(n1107) );
XOR2_X1 U982 ( .A(n1299), .B(G478), .Z(n1259) );
NAND2_X1 U983 ( .A1(n1112), .A2(n1111), .ZN(n1299) );
XNOR2_X1 U984 ( .A(n1300), .B(n1301), .ZN(n1112) );
AND2_X1 U985 ( .A1(n1302), .A2(G217), .ZN(n1301) );
NAND2_X1 U986 ( .A1(n1303), .A2(KEYINPUT55), .ZN(n1300) );
XOR2_X1 U987 ( .A(n1304), .B(n1305), .Z(n1303) );
XOR2_X1 U988 ( .A(n1306), .B(n1307), .Z(n1305) );
XOR2_X1 U989 ( .A(G143), .B(n1247), .Z(n1307) );
NAND2_X1 U990 ( .A1(KEYINPUT0), .A2(n1308), .ZN(n1306) );
XOR2_X1 U991 ( .A(n1298), .B(n1309), .Z(n1304) );
XOR2_X1 U992 ( .A(n1310), .B(n1311), .Z(n1309) );
NOR2_X1 U993 ( .A1(G107), .A2(KEYINPUT62), .ZN(n1310) );
NOR3_X1 U994 ( .A1(n1080), .A2(n1228), .A3(n1065), .ZN(n1220) );
NAND2_X1 U995 ( .A1(n1248), .A2(n1070), .ZN(n1065) );
NAND2_X1 U996 ( .A1(G214), .A2(n1312), .ZN(n1070) );
INV_X1 U997 ( .A(n1068), .ZN(n1248) );
XOR2_X1 U998 ( .A(n1096), .B(n1098), .Z(n1068) );
AND2_X1 U999 ( .A1(G210), .A2(n1312), .ZN(n1098) );
NAND2_X1 U1000 ( .A1(n1286), .A2(n1111), .ZN(n1312) );
NAND2_X1 U1001 ( .A1(n1313), .A2(n1111), .ZN(n1096) );
XOR2_X1 U1002 ( .A(n1314), .B(n1197), .Z(n1313) );
XOR2_X1 U1003 ( .A(n1140), .B(n1315), .Z(n1197) );
XOR2_X1 U1004 ( .A(n1316), .B(n1138), .Z(n1315) );
XOR2_X1 U1005 ( .A(G110), .B(n1291), .Z(n1138) );
INV_X1 U1006 ( .A(n1298), .ZN(n1291) );
XNOR2_X1 U1007 ( .A(G122), .B(KEYINPUT31), .ZN(n1298) );
NOR2_X1 U1008 ( .A1(G953), .A2(n1134), .ZN(n1316) );
INV_X1 U1009 ( .A(G224), .ZN(n1134) );
XNOR2_X1 U1010 ( .A(n1317), .B(n1318), .ZN(n1140) );
XOR2_X1 U1011 ( .A(G104), .B(n1319), .Z(n1318) );
XOR2_X1 U1012 ( .A(KEYINPUT54), .B(G107), .Z(n1319) );
XOR2_X1 U1013 ( .A(n1320), .B(G101), .Z(n1317) );
NOR2_X1 U1014 ( .A1(KEYINPUT32), .A2(n1321), .ZN(n1314) );
XOR2_X1 U1015 ( .A(n1322), .B(n1323), .Z(n1321) );
NOR2_X1 U1016 ( .A1(KEYINPUT33), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1017 ( .A(n1173), .B(KEYINPUT40), .Z(n1324) );
INV_X1 U1018 ( .A(G125), .ZN(n1322) );
INV_X1 U1019 ( .A(n1266), .ZN(n1228) );
NAND2_X1 U1020 ( .A1(n1087), .A2(n1325), .ZN(n1266) );
NAND4_X1 U1021 ( .A1(G953), .A2(G902), .A3(n1256), .A4(n1135), .ZN(n1325) );
INV_X1 U1022 ( .A(G898), .ZN(n1135) );
NAND3_X1 U1023 ( .A1(n1256), .A2(n1055), .A3(G952), .ZN(n1087) );
NAND2_X1 U1024 ( .A1(G237), .A2(G234), .ZN(n1256) );
OR2_X1 U1025 ( .A1(n1083), .A2(n1082), .ZN(n1080) );
AND2_X1 U1026 ( .A1(n1326), .A2(G221), .ZN(n1082) );
XOR2_X1 U1027 ( .A(n1327), .B(KEYINPUT27), .Z(n1326) );
XOR2_X1 U1028 ( .A(n1328), .B(G469), .Z(n1083) );
NAND2_X1 U1029 ( .A1(n1329), .A2(n1111), .ZN(n1328) );
XOR2_X1 U1030 ( .A(n1330), .B(n1331), .Z(n1329) );
XOR2_X1 U1031 ( .A(n1332), .B(n1333), .Z(n1331) );
XNOR2_X1 U1032 ( .A(n1334), .B(KEYINPUT52), .ZN(n1333) );
NAND2_X1 U1033 ( .A1(KEYINPUT8), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1034 ( .A(n1336), .B(n1187), .Z(n1335) );
AND2_X1 U1035 ( .A1(n1337), .A2(n1338), .ZN(n1187) );
OR2_X1 U1036 ( .A1(n1339), .A2(G101), .ZN(n1338) );
NAND2_X1 U1037 ( .A1(n1340), .A2(n1339), .ZN(n1337) );
NAND2_X1 U1038 ( .A1(n1341), .A2(n1342), .ZN(n1339) );
OR2_X1 U1039 ( .A1(n1343), .A2(G107), .ZN(n1342) );
XOR2_X1 U1040 ( .A(n1344), .B(KEYINPUT11), .Z(n1341) );
NAND2_X1 U1041 ( .A1(G107), .A2(n1343), .ZN(n1344) );
XNOR2_X1 U1042 ( .A(n1345), .B(KEYINPUT60), .ZN(n1343) );
INV_X1 U1043 ( .A(G104), .ZN(n1345) );
XOR2_X1 U1044 ( .A(n1166), .B(KEYINPUT43), .Z(n1340) );
NAND2_X1 U1045 ( .A1(KEYINPUT21), .A2(n1173), .ZN(n1336) );
NOR2_X1 U1046 ( .A1(KEYINPUT36), .A2(n1192), .ZN(n1332) );
NAND2_X1 U1047 ( .A1(G227), .A2(n1055), .ZN(n1192) );
XOR2_X1 U1048 ( .A(n1183), .B(n1175), .Z(n1330) );
XOR2_X1 U1049 ( .A(G110), .B(n1127), .Z(n1183) );
INV_X1 U1050 ( .A(n1086), .ZN(n1238) );
NAND2_X1 U1051 ( .A1(n1265), .A2(n1258), .ZN(n1086) );
XNOR2_X1 U1052 ( .A(n1346), .B(n1146), .ZN(n1258) );
AND2_X1 U1053 ( .A1(G217), .A2(n1327), .ZN(n1146) );
NAND2_X1 U1054 ( .A1(G234), .A2(n1111), .ZN(n1327) );
NAND2_X1 U1055 ( .A1(n1144), .A2(n1111), .ZN(n1346) );
XOR2_X1 U1056 ( .A(n1347), .B(n1348), .Z(n1144) );
XOR2_X1 U1057 ( .A(n1349), .B(n1350), .Z(n1348) );
XNOR2_X1 U1058 ( .A(n1351), .B(n1352), .ZN(n1350) );
NOR2_X1 U1059 ( .A1(KEYINPUT19), .A2(n1353), .ZN(n1352) );
XOR2_X1 U1060 ( .A(G128), .B(G119), .Z(n1353) );
NAND3_X1 U1061 ( .A1(n1302), .A2(G221), .A3(KEYINPUT47), .ZN(n1351) );
AND2_X1 U1062 ( .A1(G234), .A2(n1055), .ZN(n1302) );
NOR2_X1 U1063 ( .A1(n1354), .A2(n1355), .ZN(n1349) );
NOR3_X1 U1064 ( .A1(KEYINPUT28), .A2(G125), .A3(n1127), .ZN(n1355) );
INV_X1 U1065 ( .A(G140), .ZN(n1127) );
NOR2_X1 U1066 ( .A1(n1284), .A2(n1356), .ZN(n1354) );
INV_X1 U1067 ( .A(KEYINPUT28), .ZN(n1356) );
XOR2_X1 U1068 ( .A(G125), .B(G140), .Z(n1284) );
XNOR2_X1 U1069 ( .A(G110), .B(n1357), .ZN(n1347) );
XOR2_X1 U1070 ( .A(G146), .B(G137), .Z(n1357) );
XOR2_X1 U1071 ( .A(n1358), .B(G472), .Z(n1265) );
NAND2_X1 U1072 ( .A1(n1359), .A2(n1111), .ZN(n1358) );
INV_X1 U1073 ( .A(G902), .ZN(n1111) );
XOR2_X1 U1074 ( .A(n1360), .B(n1361), .Z(n1359) );
XNOR2_X1 U1075 ( .A(n1362), .B(KEYINPUT7), .ZN(n1361) );
NAND3_X1 U1076 ( .A1(n1363), .A2(n1165), .A3(KEYINPUT38), .ZN(n1362) );
OR2_X1 U1077 ( .A1(n1167), .A2(n1166), .ZN(n1165) );
NAND2_X1 U1078 ( .A1(n1167), .A2(n1166), .ZN(n1363) );
INV_X1 U1079 ( .A(G101), .ZN(n1166) );
NAND3_X1 U1080 ( .A1(n1286), .A2(n1055), .A3(G210), .ZN(n1167) );
INV_X1 U1081 ( .A(G953), .ZN(n1055) );
INV_X1 U1082 ( .A(G237), .ZN(n1286) );
XOR2_X1 U1083 ( .A(n1364), .B(n1365), .Z(n1360) );
INV_X1 U1084 ( .A(n1171), .ZN(n1365) );
XOR2_X1 U1085 ( .A(n1320), .B(n1366), .Z(n1171) );
XOR2_X1 U1086 ( .A(KEYINPUT25), .B(KEYINPUT10), .Z(n1366) );
XOR2_X1 U1087 ( .A(n1367), .B(n1368), .Z(n1320) );
XOR2_X1 U1088 ( .A(KEYINPUT26), .B(G119), .Z(n1368) );
XOR2_X1 U1089 ( .A(n1260), .B(n1311), .Z(n1367) );
XOR2_X1 U1090 ( .A(G116), .B(KEYINPUT50), .Z(n1311) );
INV_X1 U1091 ( .A(G113), .ZN(n1260) );
NAND2_X1 U1092 ( .A1(n1369), .A2(KEYINPUT16), .ZN(n1364) );
XOR2_X1 U1093 ( .A(n1173), .B(n1175), .Z(n1369) );
AND2_X1 U1094 ( .A1(n1370), .A2(n1371), .ZN(n1175) );
NAND2_X1 U1095 ( .A1(n1372), .A2(n1125), .ZN(n1371) );
XOR2_X1 U1096 ( .A(KEYINPUT20), .B(n1373), .Z(n1370) );
NOR2_X1 U1097 ( .A1(n1125), .A2(n1372), .ZN(n1373) );
XOR2_X1 U1098 ( .A(n1247), .B(n1374), .Z(n1372) );
NAND2_X1 U1099 ( .A1(KEYINPUT41), .A2(n1375), .ZN(n1374) );
INV_X1 U1100 ( .A(G137), .ZN(n1375) );
INV_X1 U1101 ( .A(G134), .ZN(n1247) );
INV_X1 U1102 ( .A(G131), .ZN(n1125) );
XOR2_X1 U1103 ( .A(n1376), .B(n1283), .Z(n1173) );
XOR2_X1 U1104 ( .A(G143), .B(G146), .Z(n1283) );
XOR2_X1 U1105 ( .A(n1308), .B(KEYINPUT37), .Z(n1376) );
INV_X1 U1106 ( .A(G128), .ZN(n1308) );
endmodule


