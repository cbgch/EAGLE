//Key = 1110011110010001001101100110001000001000100010001110110101010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344;

XNOR2_X1 U748 ( .A(G107), .B(n1027), .ZN(G9) );
NAND2_X1 U749 ( .A1(KEYINPUT25), .A2(n1028), .ZN(n1027) );
NOR2_X1 U750 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U751 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
NAND4_X1 U752 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1031) );
NAND4_X1 U753 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1037) );
XNOR2_X1 U754 ( .A(KEYINPUT32), .B(n1043), .ZN(n1041) );
XNOR2_X1 U755 ( .A(KEYINPUT61), .B(n1044), .ZN(n1040) );
NAND3_X1 U756 ( .A1(n1045), .A2(n1046), .A3(n1039), .ZN(n1036) );
OR2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U758 ( .A1(n1042), .A2(n1049), .ZN(n1035) );
NAND2_X1 U759 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND3_X1 U760 ( .A1(n1052), .A2(n1053), .A3(n1045), .ZN(n1051) );
NAND2_X1 U761 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NAND3_X1 U762 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
OR2_X1 U763 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND3_X1 U764 ( .A1(n1061), .A2(n1062), .A3(n1059), .ZN(n1056) );
INV_X1 U765 ( .A(n1063), .ZN(n1062) );
NAND2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1061) );
NAND2_X1 U767 ( .A1(n1060), .A2(n1066), .ZN(n1054) );
NAND2_X1 U768 ( .A1(n1039), .A2(n1067), .ZN(n1050) );
AND4_X1 U769 ( .A1(n1060), .A2(n1058), .A3(n1059), .A4(n1053), .ZN(n1039) );
NOR3_X1 U770 ( .A1(n1033), .A2(G952), .A3(n1068), .ZN(n1029) );
INV_X1 U771 ( .A(n1038), .ZN(n1068) );
NAND4_X1 U772 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1038) );
NOR3_X1 U773 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
NOR2_X1 U774 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR2_X1 U775 ( .A1(n1078), .A2(n1079), .ZN(n1074) );
NAND3_X1 U776 ( .A1(n1043), .A2(n1080), .A3(n1059), .ZN(n1073) );
NOR3_X1 U777 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1071) );
XOR2_X1 U778 ( .A(n1084), .B(KEYINPUT44), .Z(n1082) );
NAND2_X1 U779 ( .A1(n1076), .A2(n1077), .ZN(n1084) );
INV_X1 U780 ( .A(G469), .ZN(n1077) );
XOR2_X1 U781 ( .A(n1085), .B(n1086), .Z(n1070) );
XNOR2_X1 U782 ( .A(n1087), .B(n1088), .ZN(n1069) );
XOR2_X1 U783 ( .A(n1089), .B(n1090), .Z(G72) );
XOR2_X1 U784 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U785 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U786 ( .A(n1095), .B(KEYINPUT15), .Z(n1094) );
NAND2_X1 U787 ( .A1(n1096), .A2(n1097), .ZN(n1091) );
NAND2_X1 U788 ( .A1(G953), .A2(n1098), .ZN(n1097) );
XOR2_X1 U789 ( .A(n1099), .B(n1100), .Z(n1096) );
XNOR2_X1 U790 ( .A(n1101), .B(n1102), .ZN(n1100) );
XOR2_X1 U791 ( .A(n1103), .B(n1104), .Z(n1099) );
XOR2_X1 U792 ( .A(n1105), .B(KEYINPUT50), .Z(n1104) );
NAND2_X1 U793 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U794 ( .A1(G137), .A2(n1108), .ZN(n1107) );
XOR2_X1 U795 ( .A(n1109), .B(KEYINPUT58), .Z(n1106) );
NAND2_X1 U796 ( .A1(G134), .A2(n1110), .ZN(n1109) );
INV_X1 U797 ( .A(G137), .ZN(n1110) );
NAND2_X1 U798 ( .A1(KEYINPUT5), .A2(n1111), .ZN(n1103) );
NAND2_X1 U799 ( .A1(G953), .A2(n1112), .ZN(n1089) );
NAND2_X1 U800 ( .A1(G900), .A2(G227), .ZN(n1112) );
NAND3_X1 U801 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(G69) );
NAND3_X1 U802 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
OR2_X1 U803 ( .A1(n1119), .A2(KEYINPUT18), .ZN(n1117) );
NAND2_X1 U804 ( .A1(n1120), .A2(KEYINPUT18), .ZN(n1116) );
NAND2_X1 U805 ( .A1(n1121), .A2(n1095), .ZN(n1120) );
NAND3_X1 U806 ( .A1(n1122), .A2(n1123), .A3(n1095), .ZN(n1114) );
XOR2_X1 U807 ( .A(KEYINPUT18), .B(n1121), .Z(n1123) );
INV_X1 U808 ( .A(n1118), .ZN(n1122) );
NAND2_X1 U809 ( .A1(KEYINPUT52), .A2(n1034), .ZN(n1118) );
NAND2_X1 U810 ( .A1(n1124), .A2(G953), .ZN(n1113) );
NAND2_X1 U811 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U812 ( .A1(n1127), .A2(n1119), .ZN(n1126) );
NAND3_X1 U813 ( .A1(KEYINPUT18), .A2(G224), .A3(G898), .ZN(n1127) );
NAND3_X1 U814 ( .A1(KEYINPUT18), .A2(G224), .A3(n1121), .ZN(n1125) );
INV_X1 U815 ( .A(n1119), .ZN(n1121) );
NAND2_X1 U816 ( .A1(n1128), .A2(n1129), .ZN(n1119) );
NAND2_X1 U817 ( .A1(G953), .A2(n1130), .ZN(n1129) );
XOR2_X1 U818 ( .A(n1131), .B(n1132), .Z(n1128) );
NOR2_X1 U819 ( .A1(KEYINPUT54), .A2(n1133), .ZN(n1132) );
NAND3_X1 U820 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1131) );
OR2_X1 U821 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND3_X1 U822 ( .A1(n1138), .A2(n1137), .A3(KEYINPUT55), .ZN(n1135) );
NOR2_X1 U823 ( .A1(KEYINPUT56), .A2(n1139), .ZN(n1138) );
NAND2_X1 U824 ( .A1(n1139), .A2(n1140), .ZN(n1134) );
INV_X1 U825 ( .A(KEYINPUT55), .ZN(n1140) );
XOR2_X1 U826 ( .A(n1141), .B(KEYINPUT30), .Z(n1139) );
NOR2_X1 U827 ( .A1(n1142), .A2(n1143), .ZN(G66) );
NOR3_X1 U828 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1143) );
AND2_X1 U829 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U830 ( .A(KEYINPUT20), .B(n1149), .Z(n1144) );
NOR3_X1 U831 ( .A1(n1147), .A2(n1150), .A3(n1148), .ZN(n1149) );
NAND3_X1 U832 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1147) );
XOR2_X1 U833 ( .A(KEYINPUT37), .B(G217), .Z(n1153) );
NOR2_X1 U834 ( .A1(n1142), .A2(n1154), .ZN(G63) );
NOR2_X1 U835 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U836 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U837 ( .A1(n1159), .A2(G478), .ZN(n1158) );
NAND2_X1 U838 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NOR2_X1 U839 ( .A1(n1160), .A2(n1161), .ZN(n1155) );
INV_X1 U840 ( .A(KEYINPUT14), .ZN(n1161) );
NOR2_X1 U841 ( .A1(n1142), .A2(n1162), .ZN(G60) );
XOR2_X1 U842 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U843 ( .A(n1165), .B(KEYINPUT60), .Z(n1163) );
NAND2_X1 U844 ( .A1(n1159), .A2(G475), .ZN(n1165) );
XOR2_X1 U845 ( .A(G104), .B(n1166), .Z(G6) );
NOR2_X1 U846 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NOR2_X1 U847 ( .A1(n1142), .A2(n1169), .ZN(G57) );
NOR2_X1 U848 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U849 ( .A(KEYINPUT3), .B(n1172), .Z(n1171) );
NOR2_X1 U850 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U851 ( .A(n1175), .B(n1176), .Z(n1173) );
NOR2_X1 U852 ( .A1(n1177), .A2(n1178), .ZN(n1170) );
XNOR2_X1 U853 ( .A(n1175), .B(n1176), .ZN(n1178) );
NAND2_X1 U854 ( .A1(n1159), .A2(n1179), .ZN(n1175) );
XOR2_X1 U855 ( .A(KEYINPUT23), .B(G472), .Z(n1179) );
NOR2_X1 U856 ( .A1(n1142), .A2(n1180), .ZN(G54) );
XOR2_X1 U857 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U858 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND2_X1 U859 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND2_X1 U860 ( .A1(KEYINPUT42), .A2(n1187), .ZN(n1186) );
NAND2_X1 U861 ( .A1(n1188), .A2(n1189), .ZN(n1185) );
INV_X1 U862 ( .A(KEYINPUT42), .ZN(n1189) );
XOR2_X1 U863 ( .A(n1190), .B(n1191), .Z(n1181) );
NAND2_X1 U864 ( .A1(n1159), .A2(G469), .ZN(n1190) );
INV_X1 U865 ( .A(n1192), .ZN(n1159) );
NOR3_X1 U866 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(G51) );
NOR3_X1 U867 ( .A1(n1196), .A2(G953), .A3(G952), .ZN(n1195) );
AND2_X1 U868 ( .A1(n1196), .A2(n1142), .ZN(n1194) );
NOR2_X1 U869 ( .A1(n1095), .A2(G952), .ZN(n1142) );
INV_X1 U870 ( .A(KEYINPUT63), .ZN(n1196) );
XOR2_X1 U871 ( .A(n1197), .B(n1198), .Z(n1193) );
NOR2_X1 U872 ( .A1(n1088), .A2(n1192), .ZN(n1198) );
NAND2_X1 U873 ( .A1(G902), .A2(n1151), .ZN(n1192) );
NAND2_X1 U874 ( .A1(n1093), .A2(n1199), .ZN(n1151) );
INV_X1 U875 ( .A(n1034), .ZN(n1199) );
NAND4_X1 U876 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1034) );
NOR3_X1 U877 ( .A1(n1204), .A2(n1028), .A3(n1205), .ZN(n1203) );
AND4_X1 U878 ( .A1(n1067), .A2(n1047), .A3(n1060), .A4(n1206), .ZN(n1028) );
NAND2_X1 U879 ( .A1(n1066), .A2(n1207), .ZN(n1202) );
NAND3_X1 U880 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1207) );
XNOR2_X1 U881 ( .A(n1211), .B(KEYINPUT28), .ZN(n1210) );
XNOR2_X1 U882 ( .A(n1212), .B(KEYINPUT17), .ZN(n1209) );
XOR2_X1 U883 ( .A(n1168), .B(KEYINPUT47), .Z(n1208) );
NAND4_X1 U884 ( .A1(n1048), .A2(n1067), .A3(n1060), .A4(n1213), .ZN(n1168) );
INV_X1 U885 ( .A(n1032), .ZN(n1093) );
NAND4_X1 U886 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1032) );
AND4_X1 U887 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1217) );
NAND2_X1 U888 ( .A1(n1083), .A2(n1222), .ZN(n1216) );
NAND2_X1 U889 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
NAND2_X1 U890 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
NAND2_X1 U891 ( .A1(n1227), .A2(n1067), .ZN(n1223) );
NOR2_X1 U892 ( .A1(KEYINPUT43), .A2(n1228), .ZN(n1197) );
XOR2_X1 U893 ( .A(n1229), .B(n1230), .Z(n1228) );
XNOR2_X1 U894 ( .A(G146), .B(n1231), .ZN(G48) );
NAND3_X1 U895 ( .A1(n1232), .A2(n1083), .A3(n1227), .ZN(n1231) );
XOR2_X1 U896 ( .A(KEYINPUT24), .B(n1067), .Z(n1232) );
XNOR2_X1 U897 ( .A(G143), .B(n1215), .ZN(G45) );
NAND4_X1 U898 ( .A1(n1233), .A2(n1234), .A3(n1063), .A4(n1235), .ZN(n1215) );
NOR3_X1 U899 ( .A1(n1236), .A2(n1167), .A3(n1237), .ZN(n1235) );
OR2_X1 U900 ( .A1(n1047), .A2(KEYINPUT6), .ZN(n1234) );
NAND2_X1 U901 ( .A1(KEYINPUT6), .A2(n1238), .ZN(n1233) );
NAND2_X1 U902 ( .A1(n1081), .A2(n1239), .ZN(n1238) );
XNOR2_X1 U903 ( .A(n1221), .B(n1240), .ZN(G42) );
NOR2_X1 U904 ( .A1(KEYINPUT12), .A2(n1241), .ZN(n1240) );
NAND4_X1 U905 ( .A1(n1226), .A2(n1048), .A3(n1064), .A4(n1065), .ZN(n1221) );
XOR2_X1 U906 ( .A(n1242), .B(n1243), .Z(G39) );
NAND2_X1 U907 ( .A1(KEYINPUT59), .A2(n1244), .ZN(n1243) );
XOR2_X1 U908 ( .A(KEYINPUT62), .B(G137), .Z(n1244) );
NAND4_X1 U909 ( .A1(n1245), .A2(n1225), .A3(n1246), .A4(n1083), .ZN(n1242) );
XOR2_X1 U910 ( .A(n1237), .B(KEYINPUT40), .Z(n1245) );
XOR2_X1 U911 ( .A(n1108), .B(n1220), .Z(G36) );
NAND3_X1 U912 ( .A1(n1226), .A2(n1047), .A3(n1063), .ZN(n1220) );
XNOR2_X1 U913 ( .A(G131), .B(n1219), .ZN(G33) );
NAND3_X1 U914 ( .A1(n1226), .A2(n1048), .A3(n1063), .ZN(n1219) );
AND2_X1 U915 ( .A1(n1246), .A2(n1067), .ZN(n1226) );
AND3_X1 U916 ( .A1(n1058), .A2(n1059), .A3(n1247), .ZN(n1246) );
INV_X1 U917 ( .A(n1248), .ZN(n1058) );
XNOR2_X1 U918 ( .A(G128), .B(n1214), .ZN(G30) );
NAND4_X1 U919 ( .A1(n1249), .A2(n1067), .A3(n1047), .A4(n1083), .ZN(n1214) );
XOR2_X1 U920 ( .A(n1250), .B(n1251), .Z(G3) );
XOR2_X1 U921 ( .A(n1252), .B(KEYINPUT27), .Z(n1251) );
NAND3_X1 U922 ( .A1(n1211), .A2(n1066), .A3(KEYINPUT2), .ZN(n1250) );
AND4_X1 U923 ( .A1(n1063), .A2(n1067), .A3(n1213), .A4(n1042), .ZN(n1211) );
XNOR2_X1 U924 ( .A(G125), .B(n1218), .ZN(G27) );
NAND3_X1 U925 ( .A1(n1064), .A2(n1227), .A3(n1045), .ZN(n1218) );
AND2_X1 U926 ( .A1(n1048), .A2(n1249), .ZN(n1227) );
AND3_X1 U927 ( .A1(n1066), .A2(n1065), .A3(n1247), .ZN(n1249) );
INV_X1 U928 ( .A(n1236), .ZN(n1247) );
NAND2_X1 U929 ( .A1(n1253), .A2(n1053), .ZN(n1236) );
NAND2_X1 U930 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND3_X1 U931 ( .A1(G902), .A2(n1098), .A3(G953), .ZN(n1255) );
INV_X1 U932 ( .A(G900), .ZN(n1098) );
XNOR2_X1 U933 ( .A(G122), .B(n1200), .ZN(G24) );
NAND4_X1 U934 ( .A1(n1256), .A2(n1060), .A3(n1257), .A4(n1081), .ZN(n1200) );
XNOR2_X1 U935 ( .A(KEYINPUT6), .B(n1239), .ZN(n1257) );
NOR2_X1 U936 ( .A1(n1083), .A2(n1065), .ZN(n1060) );
XOR2_X1 U937 ( .A(n1258), .B(n1201), .Z(G21) );
NAND3_X1 U938 ( .A1(n1225), .A2(n1083), .A3(n1256), .ZN(n1201) );
INV_X1 U939 ( .A(n1064), .ZN(n1083) );
XNOR2_X1 U940 ( .A(G116), .B(n1259), .ZN(G18) );
NAND3_X1 U941 ( .A1(n1212), .A2(n1066), .A3(KEYINPUT19), .ZN(n1259) );
AND4_X1 U942 ( .A1(n1063), .A2(n1045), .A3(n1047), .A4(n1213), .ZN(n1212) );
XOR2_X1 U943 ( .A(G113), .B(n1204), .Z(G15) );
AND3_X1 U944 ( .A1(n1063), .A2(n1048), .A3(n1256), .ZN(n1204) );
AND2_X1 U945 ( .A1(n1045), .A2(n1206), .ZN(n1256) );
NOR2_X1 U946 ( .A1(n1044), .A2(n1260), .ZN(n1045) );
INV_X1 U947 ( .A(n1043), .ZN(n1260) );
AND2_X1 U948 ( .A1(n1261), .A2(n1239), .ZN(n1048) );
NOR2_X1 U949 ( .A1(n1065), .A2(n1064), .ZN(n1063) );
XNOR2_X1 U950 ( .A(n1205), .B(n1262), .ZN(G12) );
NAND2_X1 U951 ( .A1(KEYINPUT36), .A2(G110), .ZN(n1262) );
AND4_X1 U952 ( .A1(n1225), .A2(n1067), .A3(n1064), .A4(n1206), .ZN(n1205) );
AND2_X1 U953 ( .A1(n1213), .A2(n1066), .ZN(n1206) );
INV_X1 U954 ( .A(n1167), .ZN(n1066) );
NAND2_X1 U955 ( .A1(n1248), .A2(n1059), .ZN(n1167) );
NAND2_X1 U956 ( .A1(G214), .A2(n1263), .ZN(n1059) );
XNOR2_X1 U957 ( .A(n1264), .B(n1088), .ZN(n1248) );
NAND2_X1 U958 ( .A1(G210), .A2(n1263), .ZN(n1088) );
NAND2_X1 U959 ( .A1(n1265), .A2(n1150), .ZN(n1263) );
NAND2_X1 U960 ( .A1(KEYINPUT26), .A2(n1087), .ZN(n1264) );
NAND2_X1 U961 ( .A1(n1266), .A2(n1150), .ZN(n1087) );
XNOR2_X1 U962 ( .A(n1267), .B(n1229), .ZN(n1266) );
XNOR2_X1 U963 ( .A(n1268), .B(n1269), .ZN(n1229) );
XOR2_X1 U964 ( .A(n1133), .B(n1137), .Z(n1269) );
XNOR2_X1 U965 ( .A(n1270), .B(KEYINPUT10), .ZN(n1137) );
XOR2_X1 U966 ( .A(G110), .B(n1271), .Z(n1133) );
XOR2_X1 U967 ( .A(KEYINPUT45), .B(G122), .Z(n1271) );
XOR2_X1 U968 ( .A(n1141), .B(n1272), .Z(n1268) );
AND2_X1 U969 ( .A1(n1095), .A2(G224), .ZN(n1272) );
NAND2_X1 U970 ( .A1(n1273), .A2(n1274), .ZN(n1141) );
NAND2_X1 U971 ( .A1(KEYINPUT21), .A2(n1230), .ZN(n1267) );
XNOR2_X1 U972 ( .A(n1275), .B(G125), .ZN(n1230) );
AND2_X1 U973 ( .A1(n1276), .A2(n1053), .ZN(n1213) );
NAND2_X1 U974 ( .A1(G237), .A2(G234), .ZN(n1053) );
NAND2_X1 U975 ( .A1(n1254), .A2(n1277), .ZN(n1276) );
NAND3_X1 U976 ( .A1(n1278), .A2(n1130), .A3(G953), .ZN(n1277) );
INV_X1 U977 ( .A(G898), .ZN(n1130) );
XOR2_X1 U978 ( .A(KEYINPUT34), .B(G902), .Z(n1278) );
NAND2_X1 U979 ( .A1(G952), .A2(n1279), .ZN(n1254) );
XNOR2_X1 U980 ( .A(KEYINPUT4), .B(n1033), .ZN(n1279) );
XNOR2_X1 U981 ( .A(G953), .B(KEYINPUT0), .ZN(n1033) );
XOR2_X1 U982 ( .A(n1280), .B(G472), .Z(n1064) );
NAND2_X1 U983 ( .A1(n1281), .A2(n1150), .ZN(n1280) );
XOR2_X1 U984 ( .A(n1176), .B(n1174), .Z(n1281) );
INV_X1 U985 ( .A(n1177), .ZN(n1174) );
XOR2_X1 U986 ( .A(n1282), .B(G101), .Z(n1177) );
NAND3_X1 U987 ( .A1(n1283), .A2(n1265), .A3(G210), .ZN(n1282) );
XOR2_X1 U988 ( .A(KEYINPUT53), .B(G953), .Z(n1283) );
XNOR2_X1 U989 ( .A(n1284), .B(n1285), .ZN(n1176) );
XNOR2_X1 U990 ( .A(n1286), .B(n1275), .ZN(n1284) );
XOR2_X1 U991 ( .A(G128), .B(n1287), .Z(n1275) );
NAND3_X1 U992 ( .A1(n1288), .A2(n1289), .A3(n1274), .ZN(n1286) );
NAND2_X1 U993 ( .A1(n1290), .A2(n1258), .ZN(n1274) );
INV_X1 U994 ( .A(n1291), .ZN(n1290) );
NAND2_X1 U995 ( .A1(KEYINPUT41), .A2(n1292), .ZN(n1289) );
NAND3_X1 U996 ( .A1(n1293), .A2(n1294), .A3(n1291), .ZN(n1292) );
NAND2_X1 U997 ( .A1(n1295), .A2(G113), .ZN(n1291) );
NAND3_X1 U998 ( .A1(G119), .A2(n1296), .A3(n1297), .ZN(n1294) );
NAND2_X1 U999 ( .A1(G113), .A2(n1258), .ZN(n1293) );
OR2_X1 U1000 ( .A1(n1273), .A2(KEYINPUT41), .ZN(n1288) );
AND2_X1 U1001 ( .A1(n1298), .A2(n1299), .ZN(n1273) );
NAND2_X1 U1002 ( .A1(n1300), .A2(G119), .ZN(n1299) );
XOR2_X1 U1003 ( .A(n1297), .B(n1296), .Z(n1300) );
NAND3_X1 U1004 ( .A1(n1296), .A2(n1297), .A3(n1258), .ZN(n1298) );
INV_X1 U1005 ( .A(G113), .ZN(n1297) );
INV_X1 U1006 ( .A(n1295), .ZN(n1296) );
INV_X1 U1007 ( .A(n1237), .ZN(n1067) );
NAND2_X1 U1008 ( .A1(n1044), .A2(n1043), .ZN(n1237) );
NAND2_X1 U1009 ( .A1(G221), .A2(n1152), .ZN(n1043) );
XNOR2_X1 U1010 ( .A(n1076), .B(n1301), .ZN(n1044) );
XOR2_X1 U1011 ( .A(KEYINPUT57), .B(G469), .Z(n1301) );
AND2_X1 U1012 ( .A1(n1302), .A2(n1150), .ZN(n1076) );
XOR2_X1 U1013 ( .A(n1183), .B(n1303), .Z(n1302) );
XOR2_X1 U1014 ( .A(n1188), .B(n1304), .Z(n1303) );
NOR2_X1 U1015 ( .A1(KEYINPUT31), .A2(n1285), .ZN(n1304) );
INV_X1 U1016 ( .A(n1191), .ZN(n1285) );
XOR2_X1 U1017 ( .A(n1305), .B(n1306), .Z(n1191) );
XOR2_X1 U1018 ( .A(KEYINPUT7), .B(G137), .Z(n1306) );
XOR2_X1 U1019 ( .A(n1108), .B(n1101), .Z(n1305) );
XOR2_X1 U1020 ( .A(G131), .B(KEYINPUT8), .Z(n1101) );
XNOR2_X1 U1021 ( .A(n1307), .B(n1187), .ZN(n1188) );
XOR2_X1 U1022 ( .A(G110), .B(n1241), .Z(n1187) );
NAND2_X1 U1023 ( .A1(G227), .A2(n1095), .ZN(n1307) );
XOR2_X1 U1024 ( .A(n1308), .B(n1111), .Z(n1183) );
XOR2_X1 U1025 ( .A(G128), .B(n1309), .Z(n1111) );
NOR2_X1 U1026 ( .A1(KEYINPUT33), .A2(n1287), .ZN(n1309) );
XOR2_X1 U1027 ( .A(n1270), .B(KEYINPUT48), .Z(n1308) );
XOR2_X1 U1028 ( .A(n1252), .B(n1310), .Z(n1270) );
XOR2_X1 U1029 ( .A(G107), .B(G104), .Z(n1310) );
INV_X1 U1030 ( .A(G101), .ZN(n1252) );
AND2_X1 U1031 ( .A1(n1042), .A2(n1065), .ZN(n1225) );
XNOR2_X1 U1032 ( .A(n1311), .B(n1145), .ZN(n1065) );
INV_X1 U1033 ( .A(n1085), .ZN(n1145) );
NAND2_X1 U1034 ( .A1(n1148), .A2(n1150), .ZN(n1085) );
XNOR2_X1 U1035 ( .A(n1312), .B(n1313), .ZN(n1148) );
XOR2_X1 U1036 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1037 ( .A(G110), .B(n1316), .Z(n1315) );
NOR2_X1 U1038 ( .A1(KEYINPUT46), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1039 ( .A(G146), .B(n1318), .ZN(n1317) );
NOR2_X1 U1040 ( .A1(KEYINPUT9), .A2(n1319), .ZN(n1318) );
XOR2_X1 U1041 ( .A(G140), .B(n1320), .Z(n1319) );
NOR2_X1 U1042 ( .A1(G125), .A2(KEYINPUT16), .ZN(n1320) );
NOR4_X1 U1043 ( .A1(KEYINPUT51), .A2(G953), .A3(n1321), .A4(n1322), .ZN(n1314) );
XOR2_X1 U1044 ( .A(KEYINPUT49), .B(G221), .Z(n1322) );
INV_X1 U1045 ( .A(G234), .ZN(n1321) );
XOR2_X1 U1046 ( .A(n1258), .B(n1323), .Z(n1312) );
XOR2_X1 U1047 ( .A(G137), .B(G128), .Z(n1323) );
INV_X1 U1048 ( .A(G119), .ZN(n1258) );
NAND2_X1 U1049 ( .A1(KEYINPUT1), .A2(n1086), .ZN(n1311) );
AND2_X1 U1050 ( .A1(G217), .A2(n1152), .ZN(n1086) );
NAND2_X1 U1051 ( .A1(G234), .A2(n1324), .ZN(n1152) );
XOR2_X1 U1052 ( .A(KEYINPUT11), .B(G902), .Z(n1324) );
NAND2_X1 U1053 ( .A1(n1325), .A2(n1326), .ZN(n1042) );
OR3_X1 U1054 ( .A1(n1239), .A2(n1081), .A3(KEYINPUT35), .ZN(n1326) );
INV_X1 U1055 ( .A(n1261), .ZN(n1081) );
NAND2_X1 U1056 ( .A1(KEYINPUT35), .A2(n1047), .ZN(n1325) );
NOR2_X1 U1057 ( .A1(n1239), .A2(n1261), .ZN(n1047) );
XOR2_X1 U1058 ( .A(n1327), .B(G478), .Z(n1261) );
NAND2_X1 U1059 ( .A1(n1160), .A2(n1150), .ZN(n1327) );
XOR2_X1 U1060 ( .A(n1328), .B(n1329), .Z(n1160) );
XOR2_X1 U1061 ( .A(n1330), .B(n1331), .Z(n1329) );
XOR2_X1 U1062 ( .A(G107), .B(n1332), .Z(n1331) );
AND3_X1 U1063 ( .A1(G217), .A2(n1095), .A3(G234), .ZN(n1332) );
NOR2_X1 U1064 ( .A1(KEYINPUT29), .A2(n1295), .ZN(n1330) );
XNOR2_X1 U1065 ( .A(G116), .B(KEYINPUT22), .ZN(n1295) );
XOR2_X1 U1066 ( .A(n1333), .B(n1334), .Z(n1328) );
XOR2_X1 U1067 ( .A(G128), .B(G122), .Z(n1334) );
XOR2_X1 U1068 ( .A(G143), .B(n1108), .Z(n1333) );
INV_X1 U1069 ( .A(G134), .ZN(n1108) );
NAND3_X1 U1070 ( .A1(n1335), .A2(n1336), .A3(n1080), .ZN(n1239) );
NAND2_X1 U1071 ( .A1(n1078), .A2(n1079), .ZN(n1080) );
OR3_X1 U1072 ( .A1(n1079), .A2(n1078), .A3(KEYINPUT38), .ZN(n1336) );
INV_X1 U1073 ( .A(G475), .ZN(n1079) );
NAND2_X1 U1074 ( .A1(KEYINPUT38), .A2(n1078), .ZN(n1335) );
AND2_X1 U1075 ( .A1(n1164), .A2(n1150), .ZN(n1078) );
INV_X1 U1076 ( .A(G902), .ZN(n1150) );
XNOR2_X1 U1077 ( .A(n1337), .B(n1338), .ZN(n1164) );
XOR2_X1 U1078 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1079 ( .A(G122), .B(G113), .Z(n1340) );
XOR2_X1 U1080 ( .A(KEYINPUT13), .B(G131), .Z(n1339) );
XOR2_X1 U1081 ( .A(n1341), .B(n1342), .Z(n1337) );
XNOR2_X1 U1082 ( .A(n1343), .B(n1287), .ZN(n1342) );
XNOR2_X1 U1083 ( .A(G143), .B(G146), .ZN(n1287) );
NOR2_X1 U1084 ( .A1(KEYINPUT39), .A2(n1102), .ZN(n1343) );
XOR2_X1 U1085 ( .A(G125), .B(n1241), .Z(n1102) );
INV_X1 U1086 ( .A(G140), .ZN(n1241) );
XNOR2_X1 U1087 ( .A(G104), .B(n1344), .ZN(n1341) );
AND3_X1 U1088 ( .A1(G214), .A2(n1095), .A3(n1265), .ZN(n1344) );
INV_X1 U1089 ( .A(G237), .ZN(n1265) );
INV_X1 U1090 ( .A(G953), .ZN(n1095) );
endmodule


