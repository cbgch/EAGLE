//Key = 1001110111011000100011010000000001101010111110110010101001001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
n1519, n1520;

XNOR2_X1 U828 ( .A(n1149), .B(n1150), .ZN(G9) );
NOR3_X1 U829 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
XNOR2_X1 U830 ( .A(n1154), .B(KEYINPUT56), .ZN(n1152) );
NOR2_X1 U831 ( .A1(n1155), .A2(n1156), .ZN(G75) );
NOR3_X1 U832 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1156) );
NOR2_X1 U833 ( .A1(KEYINPUT9), .A2(n1160), .ZN(n1158) );
AND4_X1 U834 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1154), .ZN(n1160) );
NOR2_X1 U835 ( .A1(n1164), .A2(n1165), .ZN(n1161) );
NAND3_X1 U836 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1157) );
NAND2_X1 U837 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND2_X1 U838 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND3_X1 U839 ( .A1(n1163), .A2(n1173), .A3(n1162), .ZN(n1172) );
NAND3_X1 U840 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1173) );
NAND2_X1 U841 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NAND2_X1 U842 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NAND3_X1 U843 ( .A1(G221), .A2(n1181), .A3(n1182), .ZN(n1180) );
NAND2_X1 U844 ( .A1(KEYINPUT9), .A2(n1154), .ZN(n1179) );
NAND2_X1 U845 ( .A1(n1183), .A2(n1184), .ZN(n1175) );
NAND2_X1 U846 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND2_X1 U847 ( .A1(KEYINPUT41), .A2(n1187), .ZN(n1186) );
NAND2_X1 U848 ( .A1(n1188), .A2(n1189), .ZN(n1185) );
NAND3_X1 U849 ( .A1(n1187), .A2(n1190), .A3(n1191), .ZN(n1174) );
INV_X1 U850 ( .A(KEYINPUT41), .ZN(n1190) );
XOR2_X1 U851 ( .A(n1192), .B(KEYINPUT20), .Z(n1187) );
NAND3_X1 U852 ( .A1(n1183), .A2(n1193), .A3(n1177), .ZN(n1171) );
NAND2_X1 U853 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NAND2_X1 U854 ( .A1(n1163), .A2(n1196), .ZN(n1195) );
NAND2_X1 U855 ( .A1(n1197), .A2(n1151), .ZN(n1196) );
NAND2_X1 U856 ( .A1(n1162), .A2(n1198), .ZN(n1194) );
NAND2_X1 U857 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND2_X1 U858 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
INV_X1 U859 ( .A(n1203), .ZN(n1199) );
INV_X1 U860 ( .A(n1164), .ZN(n1169) );
NOR3_X1 U861 ( .A1(n1204), .A2(G953), .A3(G952), .ZN(n1155) );
INV_X1 U862 ( .A(n1166), .ZN(n1204) );
NAND4_X1 U863 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1166) );
NOR4_X1 U864 ( .A1(n1209), .A2(n1191), .A3(n1210), .A4(n1211), .ZN(n1208) );
XNOR2_X1 U865 ( .A(G472), .B(n1212), .ZN(n1211) );
XOR2_X1 U866 ( .A(KEYINPUT12), .B(n1213), .Z(n1210) );
NOR2_X1 U867 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U868 ( .A(KEYINPUT18), .B(n1216), .Z(n1215) );
XOR2_X1 U869 ( .A(n1217), .B(KEYINPUT8), .Z(n1209) );
NOR3_X1 U870 ( .A1(n1218), .A2(n1219), .A3(n1188), .ZN(n1207) );
INV_X1 U871 ( .A(n1220), .ZN(n1218) );
NAND2_X1 U872 ( .A1(n1221), .A2(n1222), .ZN(n1206) );
XNOR2_X1 U873 ( .A(G478), .B(KEYINPUT42), .ZN(n1221) );
XNOR2_X1 U874 ( .A(n1223), .B(n1224), .ZN(n1205) );
XNOR2_X1 U875 ( .A(G475), .B(KEYINPUT23), .ZN(n1224) );
NAND2_X1 U876 ( .A1(n1225), .A2(n1226), .ZN(G72) );
NAND2_X1 U877 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
XOR2_X1 U878 ( .A(n1229), .B(KEYINPUT10), .Z(n1227) );
NAND2_X1 U879 ( .A1(n1230), .A2(n1231), .ZN(n1225) );
XOR2_X1 U880 ( .A(n1229), .B(n1232), .Z(n1231) );
NOR2_X1 U881 ( .A1(n1233), .A2(KEYINPUT10), .ZN(n1232) );
NOR2_X1 U882 ( .A1(G953), .A2(n1234), .ZN(n1233) );
NAND2_X1 U883 ( .A1(n1235), .A2(n1236), .ZN(n1229) );
XOR2_X1 U884 ( .A(n1237), .B(n1238), .Z(n1235) );
XNOR2_X1 U885 ( .A(n1239), .B(n1240), .ZN(n1237) );
XOR2_X1 U886 ( .A(n1228), .B(KEYINPUT52), .Z(n1230) );
NAND2_X1 U887 ( .A1(n1236), .A2(n1241), .ZN(n1228) );
NAND2_X1 U888 ( .A1(G953), .A2(n1242), .ZN(n1241) );
INV_X1 U889 ( .A(n1243), .ZN(n1236) );
XOR2_X1 U890 ( .A(n1244), .B(n1245), .Z(G69) );
NOR2_X1 U891 ( .A1(n1246), .A2(n1167), .ZN(n1245) );
NOR2_X1 U892 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND2_X1 U893 ( .A1(n1249), .A2(n1250), .ZN(n1244) );
NAND2_X1 U894 ( .A1(n1251), .A2(n1167), .ZN(n1250) );
XOR2_X1 U895 ( .A(n1252), .B(n1253), .Z(n1251) );
OR3_X1 U896 ( .A1(n1248), .A2(n1253), .A3(n1167), .ZN(n1249) );
XNOR2_X1 U897 ( .A(n1254), .B(n1255), .ZN(n1253) );
NOR2_X1 U898 ( .A1(n1256), .A2(n1257), .ZN(G66) );
XNOR2_X1 U899 ( .A(n1258), .B(n1259), .ZN(n1257) );
NOR2_X1 U900 ( .A1(n1260), .A2(n1261), .ZN(n1258) );
NOR2_X1 U901 ( .A1(n1262), .A2(n1167), .ZN(n1256) );
XNOR2_X1 U902 ( .A(G952), .B(KEYINPUT0), .ZN(n1262) );
NOR2_X1 U903 ( .A1(n1263), .A2(n1264), .ZN(G63) );
XOR2_X1 U904 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U905 ( .A(KEYINPUT63), .B(n1267), .Z(n1266) );
AND2_X1 U906 ( .A1(G478), .A2(n1268), .ZN(n1267) );
NAND2_X1 U907 ( .A1(KEYINPUT54), .A2(n1269), .ZN(n1265) );
NOR2_X1 U908 ( .A1(n1263), .A2(n1270), .ZN(G60) );
NOR3_X1 U909 ( .A1(n1223), .A2(n1271), .A3(n1272), .ZN(n1270) );
AND3_X1 U910 ( .A1(n1273), .A2(G475), .A3(n1268), .ZN(n1272) );
NOR2_X1 U911 ( .A1(n1274), .A2(n1273), .ZN(n1271) );
AND2_X1 U912 ( .A1(n1159), .A2(G475), .ZN(n1274) );
XNOR2_X1 U913 ( .A(n1275), .B(n1276), .ZN(G6) );
NOR2_X1 U914 ( .A1(n1263), .A2(n1277), .ZN(G57) );
NOR2_X1 U915 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NOR2_X1 U916 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NOR2_X1 U917 ( .A1(n1282), .A2(n1283), .ZN(n1278) );
XNOR2_X1 U918 ( .A(n1280), .B(KEYINPUT61), .ZN(n1283) );
AND2_X1 U919 ( .A1(n1284), .A2(n1285), .ZN(n1280) );
NAND2_X1 U920 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND3_X1 U921 ( .A1(G472), .A2(n1159), .A3(n1288), .ZN(n1286) );
XNOR2_X1 U922 ( .A(KEYINPUT38), .B(G902), .ZN(n1288) );
NAND4_X1 U923 ( .A1(n1289), .A2(n1290), .A3(G472), .A4(n1291), .ZN(n1284) );
INV_X1 U924 ( .A(n1287), .ZN(n1291) );
NAND3_X1 U925 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n1287) );
INV_X1 U926 ( .A(n1295), .ZN(n1294) );
NAND2_X1 U927 ( .A1(n1296), .A2(n1297), .ZN(n1293) );
INV_X1 U928 ( .A(KEYINPUT57), .ZN(n1297) );
XOR2_X1 U929 ( .A(n1298), .B(n1299), .Z(n1296) );
NAND2_X1 U930 ( .A1(n1240), .A2(n1300), .ZN(n1298) );
NAND2_X1 U931 ( .A1(KEYINPUT57), .A2(n1301), .ZN(n1292) );
NAND2_X1 U932 ( .A1(KEYINPUT38), .A2(n1261), .ZN(n1290) );
NAND2_X1 U933 ( .A1(n1302), .A2(n1303), .ZN(n1289) );
INV_X1 U934 ( .A(KEYINPUT38), .ZN(n1303) );
NAND2_X1 U935 ( .A1(n1159), .A2(n1304), .ZN(n1302) );
XNOR2_X1 U936 ( .A(KEYINPUT15), .B(n1281), .ZN(n1282) );
OR2_X1 U937 ( .A1(n1305), .A2(n1306), .ZN(n1281) );
XNOR2_X1 U938 ( .A(n1307), .B(KEYINPUT1), .ZN(n1305) );
NAND2_X1 U939 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NOR2_X1 U940 ( .A1(n1263), .A2(n1310), .ZN(G54) );
XOR2_X1 U941 ( .A(n1311), .B(n1312), .Z(n1310) );
NAND3_X1 U942 ( .A1(n1268), .A2(G469), .A3(KEYINPUT21), .ZN(n1312) );
NAND2_X1 U943 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
NAND2_X1 U944 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XOR2_X1 U945 ( .A(KEYINPUT4), .B(n1317), .Z(n1313) );
NOR2_X1 U946 ( .A1(n1315), .A2(n1316), .ZN(n1317) );
NAND2_X1 U947 ( .A1(n1318), .A2(n1319), .ZN(n1316) );
NAND2_X1 U948 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
INV_X1 U949 ( .A(KEYINPUT44), .ZN(n1321) );
XNOR2_X1 U950 ( .A(n1322), .B(n1323), .ZN(n1320) );
NAND2_X1 U951 ( .A1(n1324), .A2(n1325), .ZN(n1322) );
NAND2_X1 U952 ( .A1(n1326), .A2(KEYINPUT44), .ZN(n1318) );
XNOR2_X1 U953 ( .A(n1323), .B(n1327), .ZN(n1326) );
XNOR2_X1 U954 ( .A(n1328), .B(n1329), .ZN(n1315) );
XNOR2_X1 U955 ( .A(n1330), .B(G110), .ZN(n1329) );
NOR2_X1 U956 ( .A1(n1263), .A2(n1331), .ZN(G51) );
XOR2_X1 U957 ( .A(n1332), .B(n1333), .Z(n1331) );
XOR2_X1 U958 ( .A(n1334), .B(n1335), .Z(n1333) );
AND2_X1 U959 ( .A1(G210), .A2(n1268), .ZN(n1335) );
INV_X1 U960 ( .A(n1261), .ZN(n1268) );
NAND2_X1 U961 ( .A1(G902), .A2(n1159), .ZN(n1261) );
NAND2_X1 U962 ( .A1(n1252), .A2(n1234), .ZN(n1159) );
AND4_X1 U963 ( .A1(n1336), .A2(n1337), .A3(n1338), .A4(n1339), .ZN(n1234) );
NOR4_X1 U964 ( .A1(n1340), .A2(n1341), .A3(n1342), .A4(n1343), .ZN(n1339) );
NOR2_X1 U965 ( .A1(n1344), .A2(n1345), .ZN(n1338) );
NAND2_X1 U966 ( .A1(n1177), .A2(n1346), .ZN(n1337) );
NAND2_X1 U967 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
NAND2_X1 U968 ( .A1(KEYINPUT16), .A2(n1349), .ZN(n1348) );
XOR2_X1 U969 ( .A(n1350), .B(KEYINPUT30), .Z(n1347) );
NAND3_X1 U970 ( .A1(n1349), .A2(n1351), .A3(n1165), .ZN(n1336) );
INV_X1 U971 ( .A(KEYINPUT16), .ZN(n1351) );
AND4_X1 U972 ( .A1(n1352), .A2(n1353), .A3(n1354), .A4(n1355), .ZN(n1252) );
NOR4_X1 U973 ( .A1(n1356), .A2(n1276), .A3(n1357), .A4(n1358), .ZN(n1355) );
NOR2_X1 U974 ( .A1(n1192), .A2(n1359), .ZN(n1358) );
INV_X1 U975 ( .A(n1360), .ZN(n1192) );
NOR3_X1 U976 ( .A1(n1151), .A2(n1361), .A3(n1153), .ZN(n1357) );
INV_X1 U977 ( .A(n1362), .ZN(n1151) );
NOR3_X1 U978 ( .A1(n1153), .A2(n1361), .A3(n1197), .ZN(n1276) );
INV_X1 U979 ( .A(n1154), .ZN(n1361) );
NAND3_X1 U980 ( .A1(n1360), .A2(n1363), .A3(n1163), .ZN(n1153) );
INV_X1 U981 ( .A(n1364), .ZN(n1356) );
AND2_X1 U982 ( .A1(n1365), .A2(n1366), .ZN(n1354) );
NOR2_X1 U983 ( .A1(KEYINPUT58), .A2(n1367), .ZN(n1334) );
XNOR2_X1 U984 ( .A(n1368), .B(n1300), .ZN(n1367) );
NOR2_X1 U985 ( .A1(G125), .A2(KEYINPUT51), .ZN(n1368) );
NOR2_X1 U986 ( .A1(n1167), .A2(G952), .ZN(n1263) );
XNOR2_X1 U987 ( .A(n1369), .B(n1344), .ZN(G48) );
AND3_X1 U988 ( .A1(n1370), .A2(n1360), .A3(n1371), .ZN(n1344) );
NAND2_X1 U989 ( .A1(n1372), .A2(n1373), .ZN(G45) );
NAND2_X1 U990 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
NAND2_X1 U991 ( .A1(G143), .A2(n1376), .ZN(n1372) );
NAND2_X1 U992 ( .A1(n1377), .A2(n1378), .ZN(n1376) );
NAND2_X1 U993 ( .A1(KEYINPUT26), .A2(n1345), .ZN(n1378) );
INV_X1 U994 ( .A(n1379), .ZN(n1345) );
OR2_X1 U995 ( .A1(n1374), .A2(KEYINPUT26), .ZN(n1377) );
NOR2_X1 U996 ( .A1(KEYINPUT13), .A2(n1379), .ZN(n1374) );
NAND4_X1 U997 ( .A1(n1380), .A2(n1360), .A3(n1381), .A4(n1382), .ZN(n1379) );
XNOR2_X1 U998 ( .A(G140), .B(n1383), .ZN(G42) );
NAND2_X1 U999 ( .A1(n1349), .A2(n1177), .ZN(n1383) );
AND2_X1 U1000 ( .A1(n1384), .A2(n1154), .ZN(n1349) );
XNOR2_X1 U1001 ( .A(n1343), .B(n1385), .ZN(G39) );
XNOR2_X1 U1002 ( .A(G137), .B(KEYINPUT6), .ZN(n1385) );
AND3_X1 U1003 ( .A1(n1371), .A2(n1162), .A3(n1177), .ZN(n1343) );
XOR2_X1 U1004 ( .A(G134), .B(n1342), .Z(G36) );
AND3_X1 U1005 ( .A1(n1380), .A2(n1362), .A3(n1177), .ZN(n1342) );
INV_X1 U1006 ( .A(n1165), .ZN(n1177) );
XOR2_X1 U1007 ( .A(G131), .B(n1386), .Z(G33) );
NOR2_X1 U1008 ( .A1(n1165), .A2(n1350), .ZN(n1386) );
NAND2_X1 U1009 ( .A1(n1380), .A2(n1370), .ZN(n1350) );
AND3_X1 U1010 ( .A1(n1203), .A2(n1387), .A3(n1154), .ZN(n1380) );
NAND2_X1 U1011 ( .A1(n1189), .A2(n1388), .ZN(n1165) );
XOR2_X1 U1012 ( .A(G128), .B(n1341), .Z(G30) );
AND3_X1 U1013 ( .A1(n1362), .A2(n1360), .A3(n1371), .ZN(n1341) );
AND4_X1 U1014 ( .A1(n1389), .A2(n1154), .A3(n1387), .A4(n1202), .ZN(n1371) );
XNOR2_X1 U1015 ( .A(G101), .B(n1364), .ZN(G3) );
NAND3_X1 U1016 ( .A1(n1360), .A2(n1203), .A3(n1390), .ZN(n1364) );
XOR2_X1 U1017 ( .A(G125), .B(n1340), .Z(G27) );
AND3_X1 U1018 ( .A1(n1183), .A2(n1360), .A3(n1384), .ZN(n1340) );
AND4_X1 U1019 ( .A1(n1370), .A2(n1201), .A3(n1387), .A4(n1202), .ZN(n1384) );
NAND2_X1 U1020 ( .A1(n1164), .A2(n1391), .ZN(n1387) );
NAND3_X1 U1021 ( .A1(G902), .A2(n1392), .A3(n1243), .ZN(n1391) );
NOR2_X1 U1022 ( .A1(G900), .A2(n1167), .ZN(n1243) );
NAND2_X1 U1023 ( .A1(n1393), .A2(n1394), .ZN(G24) );
OR2_X1 U1024 ( .A1(n1352), .A2(G122), .ZN(n1394) );
XOR2_X1 U1025 ( .A(n1395), .B(KEYINPUT48), .Z(n1393) );
NAND2_X1 U1026 ( .A1(G122), .A2(n1352), .ZN(n1395) );
NAND4_X1 U1027 ( .A1(n1396), .A2(n1163), .A3(n1381), .A4(n1382), .ZN(n1352) );
XNOR2_X1 U1028 ( .A(n1397), .B(n1353), .ZN(G21) );
NAND4_X1 U1029 ( .A1(n1162), .A2(n1396), .A3(n1389), .A4(n1202), .ZN(n1353) );
NAND2_X1 U1030 ( .A1(KEYINPUT60), .A2(n1398), .ZN(n1397) );
XNOR2_X1 U1031 ( .A(G116), .B(n1366), .ZN(G18) );
NAND3_X1 U1032 ( .A1(n1362), .A2(n1203), .A3(n1396), .ZN(n1366) );
NOR2_X1 U1033 ( .A1(n1381), .A2(n1399), .ZN(n1362) );
XNOR2_X1 U1034 ( .A(G113), .B(n1365), .ZN(G15) );
NAND3_X1 U1035 ( .A1(n1396), .A2(n1203), .A3(n1370), .ZN(n1365) );
INV_X1 U1036 ( .A(n1197), .ZN(n1370) );
NAND2_X1 U1037 ( .A1(n1399), .A2(n1381), .ZN(n1197) );
NAND2_X1 U1038 ( .A1(n1400), .A2(n1401), .ZN(n1203) );
OR3_X1 U1039 ( .A1(n1202), .A2(n1201), .A3(KEYINPUT62), .ZN(n1401) );
NAND2_X1 U1040 ( .A1(KEYINPUT62), .A2(n1163), .ZN(n1400) );
NOR2_X1 U1041 ( .A1(n1202), .A2(n1389), .ZN(n1163) );
INV_X1 U1042 ( .A(n1201), .ZN(n1389) );
AND3_X1 U1043 ( .A1(n1360), .A2(n1363), .A3(n1183), .ZN(n1396) );
INV_X1 U1044 ( .A(n1191), .ZN(n1183) );
NAND2_X1 U1045 ( .A1(n1182), .A2(n1402), .ZN(n1191) );
NAND2_X1 U1046 ( .A1(G221), .A2(n1181), .ZN(n1402) );
XOR2_X1 U1047 ( .A(n1403), .B(n1404), .Z(G12) );
NOR2_X1 U1048 ( .A1(G110), .A2(KEYINPUT17), .ZN(n1404) );
NAND2_X1 U1049 ( .A1(n1360), .A2(n1405), .ZN(n1403) );
XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n1359), .ZN(n1405) );
NAND3_X1 U1051 ( .A1(n1201), .A2(n1202), .A3(n1390), .ZN(n1359) );
AND3_X1 U1052 ( .A1(n1154), .A2(n1363), .A3(n1162), .ZN(n1390) );
NOR2_X1 U1053 ( .A1(n1382), .A2(n1381), .ZN(n1162) );
NAND2_X1 U1054 ( .A1(n1406), .A2(n1407), .ZN(n1381) );
NAND2_X1 U1055 ( .A1(n1223), .A2(n1408), .ZN(n1407) );
XOR2_X1 U1056 ( .A(n1409), .B(KEYINPUT59), .Z(n1406) );
OR2_X1 U1057 ( .A1(n1408), .A2(n1223), .ZN(n1409) );
NOR2_X1 U1058 ( .A1(n1273), .A2(G902), .ZN(n1223) );
XNOR2_X1 U1059 ( .A(n1410), .B(n1411), .ZN(n1273) );
XNOR2_X1 U1060 ( .A(n1275), .B(n1412), .ZN(n1411) );
XNOR2_X1 U1061 ( .A(n1375), .B(G131), .ZN(n1412) );
INV_X1 U1062 ( .A(G104), .ZN(n1275) );
XOR2_X1 U1063 ( .A(n1413), .B(n1414), .Z(n1410) );
NOR2_X1 U1064 ( .A1(n1415), .A2(n1416), .ZN(n1414) );
XOR2_X1 U1065 ( .A(KEYINPUT45), .B(n1417), .Z(n1416) );
AND2_X1 U1066 ( .A1(n1238), .A2(G146), .ZN(n1417) );
NOR2_X1 U1067 ( .A1(G146), .A2(n1238), .ZN(n1415) );
XOR2_X1 U1068 ( .A(n1418), .B(n1419), .Z(n1413) );
AND2_X1 U1069 ( .A1(n1420), .A2(G214), .ZN(n1419) );
NAND2_X1 U1070 ( .A1(n1421), .A2(n1422), .ZN(n1418) );
NAND2_X1 U1071 ( .A1(n1423), .A2(n1424), .ZN(n1422) );
XOR2_X1 U1072 ( .A(KEYINPUT46), .B(n1425), .Z(n1421) );
NOR2_X1 U1073 ( .A1(n1423), .A2(n1424), .ZN(n1425) );
INV_X1 U1074 ( .A(G475), .ZN(n1408) );
INV_X1 U1075 ( .A(n1399), .ZN(n1382) );
NOR2_X1 U1076 ( .A1(n1426), .A2(n1219), .ZN(n1399) );
NOR2_X1 U1077 ( .A1(n1222), .A2(G478), .ZN(n1219) );
AND2_X1 U1078 ( .A1(G478), .A2(n1222), .ZN(n1426) );
NAND2_X1 U1079 ( .A1(n1269), .A2(n1304), .ZN(n1222) );
XOR2_X1 U1080 ( .A(n1427), .B(n1428), .Z(n1269) );
XOR2_X1 U1081 ( .A(n1424), .B(n1429), .Z(n1428) );
XOR2_X1 U1082 ( .A(n1430), .B(n1431), .Z(n1429) );
NOR2_X1 U1083 ( .A1(G143), .A2(KEYINPUT27), .ZN(n1431) );
AND2_X1 U1084 ( .A1(n1432), .A2(G217), .ZN(n1430) );
XOR2_X1 U1085 ( .A(n1433), .B(n1434), .Z(n1427) );
XOR2_X1 U1086 ( .A(G134), .B(G128), .Z(n1434) );
XNOR2_X1 U1087 ( .A(G116), .B(G107), .ZN(n1433) );
NAND2_X1 U1088 ( .A1(n1164), .A2(n1435), .ZN(n1363) );
NAND4_X1 U1089 ( .A1(G953), .A2(G902), .A3(n1392), .A4(n1248), .ZN(n1435) );
INV_X1 U1090 ( .A(G898), .ZN(n1248) );
NAND3_X1 U1091 ( .A1(n1392), .A2(n1167), .A3(G952), .ZN(n1164) );
NAND2_X1 U1092 ( .A1(G237), .A2(n1436), .ZN(n1392) );
NOR2_X1 U1093 ( .A1(n1182), .A2(n1437), .ZN(n1154) );
AND2_X1 U1094 ( .A1(G221), .A2(n1181), .ZN(n1437) );
XOR2_X1 U1095 ( .A(n1438), .B(G469), .Z(n1182) );
NAND2_X1 U1096 ( .A1(n1439), .A2(n1304), .ZN(n1438) );
XOR2_X1 U1097 ( .A(n1440), .B(n1441), .Z(n1439) );
XOR2_X1 U1098 ( .A(n1442), .B(n1443), .Z(n1441) );
NAND3_X1 U1099 ( .A1(n1444), .A2(n1445), .A3(n1446), .ZN(n1443) );
NAND2_X1 U1100 ( .A1(KEYINPUT28), .A2(G140), .ZN(n1446) );
NAND3_X1 U1101 ( .A1(n1330), .A2(n1447), .A3(G110), .ZN(n1445) );
NAND2_X1 U1102 ( .A1(n1448), .A2(n1449), .ZN(n1444) );
NAND2_X1 U1103 ( .A1(n1450), .A2(n1447), .ZN(n1448) );
INV_X1 U1104 ( .A(KEYINPUT28), .ZN(n1447) );
XNOR2_X1 U1105 ( .A(KEYINPUT36), .B(n1330), .ZN(n1450) );
NAND2_X1 U1106 ( .A1(n1451), .A2(n1452), .ZN(n1442) );
OR2_X1 U1107 ( .A1(n1327), .A2(n1240), .ZN(n1452) );
XOR2_X1 U1108 ( .A(n1453), .B(KEYINPUT55), .Z(n1451) );
NAND2_X1 U1109 ( .A1(n1327), .A2(n1240), .ZN(n1453) );
XNOR2_X1 U1110 ( .A(n1325), .B(n1324), .ZN(n1327) );
XOR2_X1 U1111 ( .A(n1454), .B(n1455), .Z(n1324) );
XNOR2_X1 U1112 ( .A(n1308), .B(n1456), .ZN(n1455) );
NOR2_X1 U1113 ( .A1(KEYINPUT2), .A2(n1149), .ZN(n1456) );
XNOR2_X1 U1114 ( .A(G104), .B(KEYINPUT49), .ZN(n1454) );
XOR2_X1 U1115 ( .A(n1239), .B(KEYINPUT39), .Z(n1325) );
XNOR2_X1 U1116 ( .A(G146), .B(n1457), .ZN(n1239) );
NAND2_X1 U1117 ( .A1(KEYINPUT43), .A2(n1328), .ZN(n1440) );
NOR2_X1 U1118 ( .A1(n1242), .A2(G953), .ZN(n1328) );
INV_X1 U1119 ( .A(G227), .ZN(n1242) );
NAND2_X1 U1120 ( .A1(n1217), .A2(n1220), .ZN(n1202) );
NAND3_X1 U1121 ( .A1(n1458), .A2(n1304), .A3(n1259), .ZN(n1220) );
NAND2_X1 U1122 ( .A1(G217), .A2(n1459), .ZN(n1458) );
NAND2_X1 U1123 ( .A1(n1460), .A2(n1461), .ZN(n1217) );
NAND2_X1 U1124 ( .A1(n1259), .A2(n1304), .ZN(n1461) );
XOR2_X1 U1125 ( .A(n1462), .B(n1463), .Z(n1259) );
XOR2_X1 U1126 ( .A(n1464), .B(n1465), .Z(n1463) );
NOR2_X1 U1127 ( .A1(G146), .A2(KEYINPUT25), .ZN(n1465) );
NOR3_X1 U1128 ( .A1(n1466), .A2(n1467), .A3(n1468), .ZN(n1464) );
NOR2_X1 U1129 ( .A1(n1469), .A2(n1470), .ZN(n1468) );
AND3_X1 U1130 ( .A1(n1470), .A2(n1469), .A3(KEYINPUT47), .ZN(n1467) );
AND2_X1 U1131 ( .A1(KEYINPUT40), .A2(n1449), .ZN(n1469) );
XNOR2_X1 U1132 ( .A(G128), .B(n1471), .ZN(n1470) );
NOR2_X1 U1133 ( .A1(G119), .A2(KEYINPUT32), .ZN(n1471) );
NOR2_X1 U1134 ( .A1(KEYINPUT47), .A2(n1449), .ZN(n1466) );
INV_X1 U1135 ( .A(G110), .ZN(n1449) );
XOR2_X1 U1136 ( .A(n1472), .B(n1238), .Z(n1462) );
XNOR2_X1 U1137 ( .A(G125), .B(n1330), .ZN(n1238) );
INV_X1 U1138 ( .A(G140), .ZN(n1330) );
NAND2_X1 U1139 ( .A1(n1473), .A2(n1474), .ZN(n1472) );
NAND2_X1 U1140 ( .A1(n1475), .A2(n1476), .ZN(n1474) );
XOR2_X1 U1141 ( .A(n1477), .B(KEYINPUT34), .Z(n1475) );
NAND2_X1 U1142 ( .A1(G137), .A2(n1478), .ZN(n1473) );
XOR2_X1 U1143 ( .A(n1477), .B(KEYINPUT19), .Z(n1478) );
NAND2_X1 U1144 ( .A1(G221), .A2(n1432), .ZN(n1477) );
AND2_X1 U1145 ( .A1(n1479), .A2(n1167), .ZN(n1432) );
INV_X1 U1146 ( .A(G953), .ZN(n1167) );
XNOR2_X1 U1147 ( .A(G234), .B(KEYINPUT7), .ZN(n1479) );
INV_X1 U1148 ( .A(n1260), .ZN(n1460) );
NAND2_X1 U1149 ( .A1(G217), .A2(n1181), .ZN(n1260) );
NAND2_X1 U1150 ( .A1(n1436), .A2(n1304), .ZN(n1181) );
INV_X1 U1151 ( .A(n1459), .ZN(n1436) );
XOR2_X1 U1152 ( .A(G234), .B(KEYINPUT11), .Z(n1459) );
XOR2_X1 U1153 ( .A(n1480), .B(n1212), .Z(n1201) );
NAND2_X1 U1154 ( .A1(n1481), .A2(n1304), .ZN(n1212) );
XOR2_X1 U1155 ( .A(n1482), .B(n1483), .Z(n1481) );
NOR2_X1 U1156 ( .A1(n1295), .A2(n1301), .ZN(n1483) );
NAND2_X1 U1157 ( .A1(n1484), .A2(n1485), .ZN(n1301) );
NAND2_X1 U1158 ( .A1(n1300), .A2(n1486), .ZN(n1485) );
XNOR2_X1 U1159 ( .A(n1299), .B(n1323), .ZN(n1486) );
NAND3_X1 U1160 ( .A1(n1299), .A2(n1240), .A3(n1487), .ZN(n1484) );
NOR3_X1 U1161 ( .A1(n1240), .A2(n1299), .A3(n1300), .ZN(n1295) );
NOR2_X1 U1162 ( .A1(n1488), .A2(n1489), .ZN(n1299) );
AND2_X1 U1163 ( .A1(n1490), .A2(n1491), .ZN(n1488) );
XNOR2_X1 U1164 ( .A(KEYINPUT14), .B(n1423), .ZN(n1490) );
INV_X1 U1165 ( .A(n1492), .ZN(n1423) );
INV_X1 U1166 ( .A(n1323), .ZN(n1240) );
XOR2_X1 U1167 ( .A(G131), .B(n1493), .Z(n1323) );
XNOR2_X1 U1168 ( .A(n1476), .B(G134), .ZN(n1493) );
INV_X1 U1169 ( .A(G137), .ZN(n1476) );
NOR2_X1 U1170 ( .A1(n1306), .A2(n1494), .ZN(n1482) );
NOR2_X1 U1171 ( .A1(n1495), .A2(n1496), .ZN(n1494) );
XNOR2_X1 U1172 ( .A(KEYINPUT37), .B(n1308), .ZN(n1496) );
INV_X1 U1173 ( .A(n1309), .ZN(n1495) );
NOR2_X1 U1174 ( .A1(n1308), .A2(n1309), .ZN(n1306) );
NAND2_X1 U1175 ( .A1(G210), .A2(n1420), .ZN(n1309) );
NOR2_X1 U1176 ( .A1(G953), .A2(G237), .ZN(n1420) );
NAND2_X1 U1177 ( .A1(KEYINPUT5), .A2(n1497), .ZN(n1480) );
INV_X1 U1178 ( .A(G472), .ZN(n1497) );
NOR2_X1 U1179 ( .A1(n1189), .A2(n1188), .ZN(n1360) );
INV_X1 U1180 ( .A(n1388), .ZN(n1188) );
NAND2_X1 U1181 ( .A1(G214), .A2(n1498), .ZN(n1388) );
NOR2_X1 U1182 ( .A1(n1216), .A2(n1214), .ZN(n1189) );
AND2_X1 U1183 ( .A1(n1499), .A2(n1500), .ZN(n1214) );
NOR2_X1 U1184 ( .A1(n1499), .A2(n1500), .ZN(n1216) );
AND2_X1 U1185 ( .A1(n1501), .A2(n1304), .ZN(n1500) );
XOR2_X1 U1186 ( .A(n1502), .B(n1503), .Z(n1501) );
XOR2_X1 U1187 ( .A(KEYINPUT24), .B(G125), .Z(n1503) );
XNOR2_X1 U1188 ( .A(n1332), .B(n1487), .ZN(n1502) );
INV_X1 U1189 ( .A(n1300), .ZN(n1487) );
NAND2_X1 U1190 ( .A1(n1504), .A2(n1505), .ZN(n1300) );
NAND2_X1 U1191 ( .A1(n1457), .A2(G146), .ZN(n1505) );
NAND2_X1 U1192 ( .A1(n1506), .A2(n1369), .ZN(n1504) );
INV_X1 U1193 ( .A(G146), .ZN(n1369) );
XNOR2_X1 U1194 ( .A(n1457), .B(KEYINPUT22), .ZN(n1506) );
XNOR2_X1 U1195 ( .A(G128), .B(n1375), .ZN(n1457) );
INV_X1 U1196 ( .A(G143), .ZN(n1375) );
XNOR2_X1 U1197 ( .A(n1507), .B(n1255), .ZN(n1332) );
XNOR2_X1 U1198 ( .A(n1508), .B(n1509), .ZN(n1255) );
NOR2_X1 U1199 ( .A1(n1510), .A2(n1489), .ZN(n1509) );
NOR2_X1 U1200 ( .A1(n1491), .A2(n1492), .ZN(n1489) );
AND2_X1 U1201 ( .A1(n1492), .A2(n1491), .ZN(n1510) );
XNOR2_X1 U1202 ( .A(G116), .B(n1398), .ZN(n1491) );
INV_X1 U1203 ( .A(G119), .ZN(n1398) );
XOR2_X1 U1204 ( .A(G113), .B(KEYINPUT31), .Z(n1492) );
NAND3_X1 U1205 ( .A1(n1511), .A2(n1512), .A3(n1513), .ZN(n1508) );
NAND2_X1 U1206 ( .A1(G101), .A2(n1514), .ZN(n1513) );
OR3_X1 U1207 ( .A1(n1514), .A2(G101), .A3(n1515), .ZN(n1512) );
INV_X1 U1208 ( .A(KEYINPUT3), .ZN(n1514) );
NAND2_X1 U1209 ( .A1(n1515), .A2(n1516), .ZN(n1511) );
NAND2_X1 U1210 ( .A1(KEYINPUT3), .A2(n1517), .ZN(n1516) );
XNOR2_X1 U1211 ( .A(KEYINPUT33), .B(n1308), .ZN(n1517) );
INV_X1 U1212 ( .A(G101), .ZN(n1308) );
XNOR2_X1 U1213 ( .A(G104), .B(n1149), .ZN(n1515) );
INV_X1 U1214 ( .A(G107), .ZN(n1149) );
XOR2_X1 U1215 ( .A(n1518), .B(n1519), .Z(n1507) );
NOR2_X1 U1216 ( .A1(G953), .A2(n1247), .ZN(n1519) );
INV_X1 U1217 ( .A(G224), .ZN(n1247) );
NAND2_X1 U1218 ( .A1(KEYINPUT50), .A2(n1254), .ZN(n1518) );
XNOR2_X1 U1219 ( .A(G110), .B(n1424), .ZN(n1254) );
XOR2_X1 U1220 ( .A(G122), .B(KEYINPUT29), .Z(n1424) );
NAND2_X1 U1221 ( .A1(G210), .A2(n1498), .ZN(n1499) );
NAND2_X1 U1222 ( .A1(n1520), .A2(n1304), .ZN(n1498) );
INV_X1 U1223 ( .A(G902), .ZN(n1304) );
XNOR2_X1 U1224 ( .A(G237), .B(KEYINPUT35), .ZN(n1520) );
endmodule


