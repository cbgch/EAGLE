//Key = 0010110111100101110111101100000101011101001111000101011101111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344;

XOR2_X1 U729 ( .A(G107), .B(n1020), .Z(G9) );
AND3_X1 U730 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NOR2_X1 U731 ( .A1(n1024), .A2(n1025), .ZN(G75) );
NOR4_X1 U732 ( .A1(G953), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1025) );
NOR2_X1 U733 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U734 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U735 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR2_X1 U736 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U737 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U738 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR2_X1 U739 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR3_X1 U740 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1041) );
NOR2_X1 U741 ( .A1(KEYINPUT59), .A2(n1046), .ZN(n1045) );
NOR2_X1 U742 ( .A1(n1047), .A2(n1048), .ZN(n1043) );
NOR2_X1 U743 ( .A1(n1049), .A2(n1046), .ZN(n1039) );
NOR2_X1 U744 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR3_X1 U745 ( .A1(n1046), .A2(n1052), .A3(n1042), .ZN(n1035) );
NOR2_X1 U746 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR3_X1 U747 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1053) );
INV_X1 U748 ( .A(KEYINPUT59), .ZN(n1055) );
NOR4_X1 U749 ( .A1(n1058), .A2(n1042), .A3(n1038), .A4(n1046), .ZN(n1031) );
INV_X1 U750 ( .A(n1023), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1021), .A2(n1059), .ZN(n1058) );
NOR3_X1 U752 ( .A1(n1026), .A2(G953), .A3(G952), .ZN(n1024) );
AND4_X1 U753 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1026) );
NOR3_X1 U754 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
NAND3_X1 U755 ( .A1(n1048), .A2(n1067), .A3(n1068), .ZN(n1064) );
OR2_X1 U756 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NOR3_X1 U757 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1062) );
AND2_X1 U758 ( .A1(n1074), .A2(KEYINPUT23), .ZN(n1073) );
NOR3_X1 U759 ( .A1(KEYINPUT23), .A2(n1075), .A3(n1074), .ZN(n1072) );
XNOR2_X1 U760 ( .A(G475), .B(n1076), .ZN(n1071) );
XOR2_X1 U761 ( .A(n1077), .B(KEYINPUT0), .Z(n1060) );
NAND2_X1 U762 ( .A1(n1070), .A2(n1069), .ZN(n1077) );
XOR2_X1 U763 ( .A(n1078), .B(n1079), .Z(G72) );
XOR2_X1 U764 ( .A(n1080), .B(n1081), .Z(n1079) );
NAND2_X1 U765 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U766 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U767 ( .A1(n1086), .A2(n1087), .ZN(n1080) );
NAND2_X1 U768 ( .A1(G953), .A2(n1088), .ZN(n1087) );
XNOR2_X1 U769 ( .A(KEYINPUT15), .B(n1089), .ZN(n1088) );
XOR2_X1 U770 ( .A(n1090), .B(n1091), .Z(n1086) );
XOR2_X1 U771 ( .A(n1092), .B(n1093), .Z(n1091) );
XNOR2_X1 U772 ( .A(n1094), .B(n1095), .ZN(n1090) );
NAND2_X1 U773 ( .A1(KEYINPUT55), .A2(n1096), .ZN(n1094) );
NOR2_X1 U774 ( .A1(n1097), .A2(n1082), .ZN(n1078) );
AND2_X1 U775 ( .A1(G227), .A2(G900), .ZN(n1097) );
XOR2_X1 U776 ( .A(n1098), .B(n1099), .Z(G69) );
NOR2_X1 U777 ( .A1(n1100), .A2(n1082), .ZN(n1099) );
NOR2_X1 U778 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U779 ( .A1(n1103), .A2(n1104), .ZN(n1098) );
NAND2_X1 U780 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U781 ( .A(n1107), .B(n1108), .Z(n1103) );
NOR2_X1 U782 ( .A1(n1109), .A2(G953), .ZN(n1108) );
OR2_X1 U783 ( .A1(n1105), .A2(n1106), .ZN(n1107) );
NAND2_X1 U784 ( .A1(n1110), .A2(n1111), .ZN(n1106) );
NAND2_X1 U785 ( .A1(G953), .A2(n1112), .ZN(n1111) );
XNOR2_X1 U786 ( .A(KEYINPUT43), .B(n1102), .ZN(n1112) );
INV_X1 U787 ( .A(KEYINPUT7), .ZN(n1105) );
NOR3_X1 U788 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(G66) );
AND2_X1 U789 ( .A1(KEYINPUT37), .A2(n1116), .ZN(n1115) );
NOR3_X1 U790 ( .A1(KEYINPUT37), .A2(n1082), .A3(n1117), .ZN(n1114) );
INV_X1 U791 ( .A(G952), .ZN(n1117) );
XOR2_X1 U792 ( .A(n1118), .B(n1119), .Z(n1113) );
NAND2_X1 U793 ( .A1(KEYINPUT44), .A2(n1120), .ZN(n1119) );
NAND2_X1 U794 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
XOR2_X1 U795 ( .A(KEYINPUT29), .B(G217), .Z(n1122) );
NOR2_X1 U796 ( .A1(n1116), .A2(n1123), .ZN(G63) );
XOR2_X1 U797 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND3_X1 U798 ( .A1(n1121), .A2(G478), .A3(KEYINPUT20), .ZN(n1124) );
NOR2_X1 U799 ( .A1(n1116), .A2(n1126), .ZN(G60) );
XOR2_X1 U800 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U801 ( .A1(KEYINPUT47), .A2(n1129), .ZN(n1128) );
XNOR2_X1 U802 ( .A(n1130), .B(n1131), .ZN(n1129) );
NAND2_X1 U803 ( .A1(n1121), .A2(G475), .ZN(n1127) );
XOR2_X1 U804 ( .A(G104), .B(n1132), .Z(G6) );
NOR2_X1 U805 ( .A1(n1133), .A2(n1134), .ZN(G57) );
XNOR2_X1 U806 ( .A(n1116), .B(KEYINPUT31), .ZN(n1134) );
XNOR2_X1 U807 ( .A(n1135), .B(n1136), .ZN(n1133) );
XOR2_X1 U808 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U809 ( .A1(KEYINPUT50), .A2(n1139), .ZN(n1138) );
AND2_X1 U810 ( .A1(G472), .A2(n1121), .ZN(n1137) );
NOR2_X1 U811 ( .A1(n1116), .A2(n1140), .ZN(G54) );
XNOR2_X1 U812 ( .A(n1141), .B(n1142), .ZN(n1140) );
XOR2_X1 U813 ( .A(n1143), .B(n1144), .Z(n1142) );
AND2_X1 U814 ( .A1(G469), .A2(n1121), .ZN(n1144) );
INV_X1 U815 ( .A(n1145), .ZN(n1121) );
NAND3_X1 U816 ( .A1(n1146), .A2(n1147), .A3(KEYINPUT58), .ZN(n1143) );
NAND2_X1 U817 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U818 ( .A(KEYINPUT24), .B(n1150), .Z(n1146) );
NOR2_X1 U819 ( .A1(n1149), .A2(n1151), .ZN(n1150) );
XOR2_X1 U820 ( .A(KEYINPUT28), .B(n1148), .Z(n1151) );
XNOR2_X1 U821 ( .A(n1152), .B(G140), .ZN(n1148) );
NOR3_X1 U822 ( .A1(n1116), .A2(n1153), .A3(n1154), .ZN(G51) );
NOR2_X1 U823 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U824 ( .A(KEYINPUT61), .B(n1157), .Z(n1156) );
NOR2_X1 U825 ( .A1(n1110), .A2(n1158), .ZN(n1153) );
XNOR2_X1 U826 ( .A(n1157), .B(KEYINPUT27), .ZN(n1158) );
XOR2_X1 U827 ( .A(n1159), .B(n1160), .Z(n1157) );
NOR2_X1 U828 ( .A1(n1069), .A2(n1145), .ZN(n1160) );
NAND2_X1 U829 ( .A1(G902), .A2(n1028), .ZN(n1145) );
NAND3_X1 U830 ( .A1(n1084), .A2(n1161), .A3(n1109), .ZN(n1028) );
AND4_X1 U831 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1109) );
NOR4_X1 U832 ( .A1(n1166), .A2(n1167), .A3(n1132), .A4(n1168), .ZN(n1165) );
INV_X1 U833 ( .A(n1169), .ZN(n1168) );
AND3_X1 U834 ( .A1(n1023), .A2(n1022), .A3(n1059), .ZN(n1132) );
AND2_X1 U835 ( .A1(n1170), .A2(n1171), .ZN(n1164) );
NAND3_X1 U836 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1163) );
NAND2_X1 U837 ( .A1(n1175), .A2(n1176), .ZN(n1173) );
INV_X1 U838 ( .A(KEYINPUT60), .ZN(n1176) );
NAND2_X1 U839 ( .A1(KEYINPUT60), .A2(n1177), .ZN(n1172) );
NAND4_X1 U840 ( .A1(n1021), .A2(n1023), .A3(n1178), .A4(n1179), .ZN(n1162) );
NAND2_X1 U841 ( .A1(n1175), .A2(n1180), .ZN(n1179) );
INV_X1 U842 ( .A(KEYINPUT53), .ZN(n1180) );
NAND3_X1 U843 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1175) );
NAND2_X1 U844 ( .A1(KEYINPUT53), .A2(n1177), .ZN(n1178) );
XNOR2_X1 U845 ( .A(KEYINPUT57), .B(n1085), .ZN(n1161) );
OR3_X1 U846 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1085) );
XNOR2_X1 U847 ( .A(KEYINPUT62), .B(n1187), .ZN(n1185) );
AND4_X1 U848 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1084) );
NOR4_X1 U849 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
INV_X1 U850 ( .A(n1196), .ZN(n1192) );
NAND2_X1 U851 ( .A1(n1197), .A2(n1198), .ZN(n1190) );
INV_X1 U852 ( .A(n1199), .ZN(n1198) );
XOR2_X1 U853 ( .A(n1046), .B(KEYINPUT13), .Z(n1197) );
NOR2_X1 U854 ( .A1(n1082), .A2(G952), .ZN(n1116) );
XNOR2_X1 U855 ( .A(n1200), .B(n1201), .ZN(G48) );
NOR2_X1 U856 ( .A1(n1202), .A2(n1186), .ZN(n1201) );
NAND3_X1 U857 ( .A1(n1044), .A2(n1203), .A3(n1059), .ZN(n1186) );
NAND2_X1 U858 ( .A1(n1204), .A2(n1205), .ZN(G45) );
NAND2_X1 U859 ( .A1(G143), .A2(n1188), .ZN(n1205) );
XOR2_X1 U860 ( .A(KEYINPUT21), .B(n1206), .Z(n1204) );
NOR2_X1 U861 ( .A1(G143), .A2(n1188), .ZN(n1206) );
NAND3_X1 U862 ( .A1(n1207), .A2(n1050), .A3(n1208), .ZN(n1188) );
NOR3_X1 U863 ( .A1(n1182), .A2(n1209), .A3(n1210), .ZN(n1208) );
XOR2_X1 U864 ( .A(G140), .B(n1211), .Z(G42) );
NOR2_X1 U865 ( .A1(n1046), .A2(n1199), .ZN(n1211) );
NAND3_X1 U866 ( .A1(n1059), .A2(n1051), .A3(n1207), .ZN(n1199) );
XOR2_X1 U867 ( .A(n1212), .B(G137), .Z(G39) );
NAND2_X1 U868 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND4_X1 U869 ( .A1(n1215), .A2(n1054), .A3(n1187), .A4(n1216), .ZN(n1214) );
OR2_X1 U870 ( .A1(n1189), .A2(n1216), .ZN(n1213) );
INV_X1 U871 ( .A(KEYINPUT2), .ZN(n1216) );
NAND2_X1 U872 ( .A1(n1215), .A2(n1207), .ZN(n1189) );
NOR3_X1 U873 ( .A1(n1034), .A2(n1217), .A3(n1046), .ZN(n1215) );
XOR2_X1 U874 ( .A(G134), .B(n1194), .Z(G36) );
AND2_X1 U875 ( .A1(n1218), .A2(n1021), .ZN(n1194) );
XOR2_X1 U876 ( .A(n1219), .B(n1193), .Z(G33) );
AND2_X1 U877 ( .A1(n1218), .A2(n1059), .ZN(n1193) );
NOR3_X1 U878 ( .A1(n1046), .A2(n1220), .A3(n1202), .ZN(n1218) );
INV_X1 U879 ( .A(n1207), .ZN(n1202) );
NOR2_X1 U880 ( .A1(n1184), .A2(n1187), .ZN(n1207) );
NAND2_X1 U881 ( .A1(n1221), .A2(n1048), .ZN(n1046) );
XNOR2_X1 U882 ( .A(G131), .B(KEYINPUT35), .ZN(n1219) );
NAND2_X1 U883 ( .A1(n1222), .A2(n1223), .ZN(G30) );
NAND2_X1 U884 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NAND2_X1 U885 ( .A1(G128), .A2(n1226), .ZN(n1222) );
NAND2_X1 U886 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NAND2_X1 U887 ( .A1(KEYINPUT56), .A2(n1195), .ZN(n1228) );
INV_X1 U888 ( .A(n1229), .ZN(n1195) );
OR2_X1 U889 ( .A1(n1224), .A2(KEYINPUT56), .ZN(n1227) );
NOR2_X1 U890 ( .A1(KEYINPUT6), .A2(n1229), .ZN(n1224) );
NAND4_X1 U891 ( .A1(n1021), .A2(n1044), .A3(n1230), .A4(n1183), .ZN(n1229) );
NOR2_X1 U892 ( .A1(n1187), .A2(n1217), .ZN(n1230) );
INV_X1 U893 ( .A(n1203), .ZN(n1217) );
INV_X1 U894 ( .A(n1231), .ZN(n1187) );
XOR2_X1 U895 ( .A(G101), .B(n1232), .Z(G3) );
AND2_X1 U896 ( .A1(n1022), .A2(n1174), .ZN(n1232) );
NOR2_X1 U897 ( .A1(n1220), .A2(n1034), .ZN(n1174) );
INV_X1 U898 ( .A(n1233), .ZN(n1034) );
INV_X1 U899 ( .A(n1050), .ZN(n1220) );
XNOR2_X1 U900 ( .A(G125), .B(n1196), .ZN(G27) );
NAND4_X1 U901 ( .A1(n1051), .A2(n1231), .A3(n1044), .A4(n1234), .ZN(n1196) );
AND2_X1 U902 ( .A1(n1061), .A2(n1059), .ZN(n1234) );
NAND2_X1 U903 ( .A1(n1030), .A2(n1235), .ZN(n1231) );
NAND4_X1 U904 ( .A1(G902), .A2(G953), .A3(n1236), .A4(n1089), .ZN(n1235) );
INV_X1 U905 ( .A(G900), .ZN(n1089) );
XNOR2_X1 U906 ( .A(G122), .B(n1237), .ZN(G24) );
NAND2_X1 U907 ( .A1(KEYINPUT39), .A2(n1167), .ZN(n1237) );
AND4_X1 U908 ( .A1(n1238), .A2(n1023), .A3(n1239), .A4(n1240), .ZN(n1167) );
XNOR2_X1 U909 ( .A(n1241), .B(n1242), .ZN(G21) );
NOR2_X1 U910 ( .A1(KEYINPUT3), .A2(n1171), .ZN(n1242) );
NAND3_X1 U911 ( .A1(n1233), .A2(n1203), .A3(n1238), .ZN(n1171) );
NAND2_X1 U912 ( .A1(n1243), .A2(n1244), .ZN(n1203) );
NAND3_X1 U913 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1244) );
NAND2_X1 U914 ( .A1(KEYINPUT48), .A2(n1050), .ZN(n1243) );
XNOR2_X1 U915 ( .A(G116), .B(n1170), .ZN(G18) );
NAND3_X1 U916 ( .A1(n1238), .A2(n1021), .A3(n1050), .ZN(n1170) );
NOR2_X1 U917 ( .A1(n1240), .A2(n1210), .ZN(n1021) );
XNOR2_X1 U918 ( .A(G113), .B(n1169), .ZN(G15) );
NAND3_X1 U919 ( .A1(n1059), .A2(n1238), .A3(n1050), .ZN(n1169) );
NOR2_X1 U920 ( .A1(n1248), .A2(n1246), .ZN(n1050) );
AND3_X1 U921 ( .A1(n1044), .A2(n1181), .A3(n1061), .ZN(n1238) );
INV_X1 U922 ( .A(n1038), .ZN(n1061) );
NAND2_X1 U923 ( .A1(n1249), .A2(n1056), .ZN(n1038) );
INV_X1 U924 ( .A(n1057), .ZN(n1249) );
NOR2_X1 U925 ( .A1(n1239), .A2(n1209), .ZN(n1059) );
INV_X1 U926 ( .A(n1240), .ZN(n1209) );
XNOR2_X1 U927 ( .A(n1166), .B(n1250), .ZN(G12) );
NAND2_X1 U928 ( .A1(KEYINPUT36), .A2(G110), .ZN(n1250) );
AND3_X1 U929 ( .A1(n1022), .A2(n1051), .A3(n1233), .ZN(n1166) );
NOR2_X1 U930 ( .A1(n1240), .A2(n1239), .ZN(n1233) );
INV_X1 U931 ( .A(n1210), .ZN(n1239) );
XOR2_X1 U932 ( .A(n1066), .B(KEYINPUT4), .Z(n1210) );
XNOR2_X1 U933 ( .A(n1251), .B(G478), .ZN(n1066) );
NAND2_X1 U934 ( .A1(n1125), .A2(n1252), .ZN(n1251) );
XNOR2_X1 U935 ( .A(n1253), .B(n1254), .ZN(n1125) );
AND3_X1 U936 ( .A1(G234), .A2(n1082), .A3(G217), .ZN(n1254) );
NAND2_X1 U937 ( .A1(n1255), .A2(KEYINPUT10), .ZN(n1253) );
XOR2_X1 U938 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U939 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U940 ( .A(G134), .B(G122), .Z(n1259) );
XOR2_X1 U941 ( .A(KEYINPUT32), .B(KEYINPUT19), .Z(n1258) );
XOR2_X1 U942 ( .A(n1260), .B(n1261), .Z(n1256) );
XNOR2_X1 U943 ( .A(G107), .B(G116), .ZN(n1260) );
NAND2_X1 U944 ( .A1(n1262), .A2(n1263), .ZN(n1240) );
NAND2_X1 U945 ( .A1(G475), .A2(n1076), .ZN(n1263) );
XOR2_X1 U946 ( .A(n1264), .B(KEYINPUT40), .Z(n1262) );
OR2_X1 U947 ( .A1(n1076), .A2(G475), .ZN(n1264) );
NAND2_X1 U948 ( .A1(n1265), .A2(n1252), .ZN(n1076) );
XNOR2_X1 U949 ( .A(n1130), .B(n1266), .ZN(n1265) );
INV_X1 U950 ( .A(n1131), .ZN(n1266) );
XNOR2_X1 U951 ( .A(n1267), .B(n1268), .ZN(n1131) );
XNOR2_X1 U952 ( .A(KEYINPUT1), .B(n1200), .ZN(n1268) );
XNOR2_X1 U953 ( .A(G122), .B(G125), .ZN(n1267) );
XOR2_X1 U954 ( .A(n1269), .B(n1270), .Z(n1130) );
XNOR2_X1 U955 ( .A(n1271), .B(n1272), .ZN(n1270) );
NOR2_X1 U956 ( .A1(G140), .A2(KEYINPUT12), .ZN(n1272) );
NAND2_X1 U957 ( .A1(KEYINPUT17), .A2(n1273), .ZN(n1271) );
XOR2_X1 U958 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U959 ( .A(G131), .B(G143), .ZN(n1275) );
NAND2_X1 U960 ( .A1(G214), .A2(n1276), .ZN(n1274) );
XNOR2_X1 U961 ( .A(G104), .B(G113), .ZN(n1269) );
NAND2_X1 U962 ( .A1(n1277), .A2(n1278), .ZN(n1051) );
NAND3_X1 U963 ( .A1(n1248), .A2(n1246), .A3(n1247), .ZN(n1278) );
INV_X1 U964 ( .A(KEYINPUT48), .ZN(n1247) );
NAND2_X1 U965 ( .A1(KEYINPUT48), .A2(n1023), .ZN(n1277) );
NOR2_X1 U966 ( .A1(n1246), .A2(n1245), .ZN(n1023) );
INV_X1 U967 ( .A(n1248), .ZN(n1245) );
XOR2_X1 U968 ( .A(n1065), .B(KEYINPUT22), .Z(n1248) );
XNOR2_X1 U969 ( .A(n1279), .B(G472), .ZN(n1065) );
NAND2_X1 U970 ( .A1(n1280), .A2(n1252), .ZN(n1279) );
XNOR2_X1 U971 ( .A(n1139), .B(n1135), .ZN(n1280) );
XNOR2_X1 U972 ( .A(n1281), .B(n1282), .ZN(n1135) );
XOR2_X1 U973 ( .A(n1283), .B(n1284), .Z(n1282) );
NAND2_X1 U974 ( .A1(KEYINPUT25), .A2(n1241), .ZN(n1284) );
NAND2_X1 U975 ( .A1(G210), .A2(n1276), .ZN(n1283) );
NOR2_X1 U976 ( .A1(G953), .A2(G237), .ZN(n1276) );
XNOR2_X1 U977 ( .A(G101), .B(n1285), .ZN(n1281) );
XNOR2_X1 U978 ( .A(n1286), .B(G113), .ZN(n1285) );
XNOR2_X1 U979 ( .A(n1287), .B(n1288), .ZN(n1139) );
NAND2_X1 U980 ( .A1(n1067), .A2(n1289), .ZN(n1246) );
OR2_X1 U981 ( .A1(n1074), .A2(n1075), .ZN(n1289) );
NAND2_X1 U982 ( .A1(n1075), .A2(n1074), .ZN(n1067) );
NAND2_X1 U983 ( .A1(G217), .A2(n1290), .ZN(n1074) );
NOR2_X1 U984 ( .A1(n1120), .A2(G902), .ZN(n1075) );
XNOR2_X1 U985 ( .A(n1291), .B(n1292), .ZN(n1120) );
XOR2_X1 U986 ( .A(n1093), .B(n1293), .Z(n1292) );
XOR2_X1 U987 ( .A(n1294), .B(n1295), .Z(n1293) );
NAND2_X1 U988 ( .A1(KEYINPUT9), .A2(n1200), .ZN(n1295) );
INV_X1 U989 ( .A(G146), .ZN(n1200) );
NAND3_X1 U990 ( .A1(G234), .A2(n1296), .A3(G221), .ZN(n1294) );
XNOR2_X1 U991 ( .A(KEYINPUT49), .B(n1082), .ZN(n1296) );
XNOR2_X1 U992 ( .A(n1297), .B(G140), .ZN(n1093) );
XOR2_X1 U993 ( .A(n1298), .B(n1299), .Z(n1291) );
XOR2_X1 U994 ( .A(G137), .B(n1300), .Z(n1299) );
NOR2_X1 U995 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
XOR2_X1 U996 ( .A(n1303), .B(KEYINPUT42), .Z(n1302) );
NAND2_X1 U997 ( .A1(G110), .A2(n1304), .ZN(n1303) );
NOR2_X1 U998 ( .A1(G110), .A2(n1304), .ZN(n1301) );
XNOR2_X1 U999 ( .A(n1241), .B(n1305), .ZN(n1304) );
XNOR2_X1 U1000 ( .A(KEYINPUT11), .B(n1225), .ZN(n1305) );
INV_X1 U1001 ( .A(G119), .ZN(n1241) );
XNOR2_X1 U1002 ( .A(KEYINPUT18), .B(KEYINPUT14), .ZN(n1298) );
INV_X1 U1003 ( .A(n1177), .ZN(n1022) );
NAND3_X1 U1004 ( .A1(n1183), .A2(n1181), .A3(n1044), .ZN(n1177) );
INV_X1 U1005 ( .A(n1182), .ZN(n1044) );
NAND2_X1 U1006 ( .A1(n1047), .A2(n1048), .ZN(n1182) );
NAND2_X1 U1007 ( .A1(G214), .A2(n1306), .ZN(n1048) );
INV_X1 U1008 ( .A(n1221), .ZN(n1047) );
XNOR2_X1 U1009 ( .A(n1307), .B(n1069), .ZN(n1221) );
NAND2_X1 U1010 ( .A1(G210), .A2(n1306), .ZN(n1069) );
NAND2_X1 U1011 ( .A1(n1308), .A2(n1252), .ZN(n1306) );
INV_X1 U1012 ( .A(G237), .ZN(n1308) );
XNOR2_X1 U1013 ( .A(n1070), .B(KEYINPUT52), .ZN(n1307) );
AND2_X1 U1014 ( .A1(n1309), .A2(n1252), .ZN(n1070) );
XNOR2_X1 U1015 ( .A(n1310), .B(n1155), .ZN(n1309) );
INV_X1 U1016 ( .A(n1110), .ZN(n1155) );
XNOR2_X1 U1017 ( .A(n1311), .B(n1312), .ZN(n1110) );
XOR2_X1 U1018 ( .A(n1313), .B(n1314), .Z(n1312) );
XNOR2_X1 U1019 ( .A(G119), .B(G122), .ZN(n1314) );
NAND2_X1 U1020 ( .A1(KEYINPUT5), .A2(n1315), .ZN(n1313) );
INV_X1 U1021 ( .A(G113), .ZN(n1315) );
XOR2_X1 U1022 ( .A(n1316), .B(n1317), .Z(n1311) );
XNOR2_X1 U1023 ( .A(n1318), .B(n1319), .ZN(n1317) );
NOR2_X1 U1024 ( .A1(G110), .A2(KEYINPUT34), .ZN(n1319) );
NAND2_X1 U1025 ( .A1(KEYINPUT8), .A2(n1286), .ZN(n1318) );
INV_X1 U1026 ( .A(G116), .ZN(n1286) );
NOR2_X1 U1027 ( .A1(KEYINPUT30), .A2(n1159), .ZN(n1310) );
XNOR2_X1 U1028 ( .A(n1320), .B(n1321), .ZN(n1159) );
XNOR2_X1 U1029 ( .A(KEYINPUT46), .B(n1297), .ZN(n1321) );
INV_X1 U1030 ( .A(G125), .ZN(n1297) );
XOR2_X1 U1031 ( .A(n1287), .B(n1322), .Z(n1320) );
NOR2_X1 U1032 ( .A1(G953), .A2(n1101), .ZN(n1322) );
INV_X1 U1033 ( .A(G224), .ZN(n1101) );
XNOR2_X1 U1034 ( .A(G146), .B(n1261), .ZN(n1287) );
XNOR2_X1 U1035 ( .A(n1225), .B(G143), .ZN(n1261) );
INV_X1 U1036 ( .A(G128), .ZN(n1225) );
NAND2_X1 U1037 ( .A1(n1030), .A2(n1323), .ZN(n1181) );
NAND4_X1 U1038 ( .A1(G902), .A2(G953), .A3(n1236), .A4(n1102), .ZN(n1323) );
INV_X1 U1039 ( .A(G898), .ZN(n1102) );
NAND3_X1 U1040 ( .A1(n1236), .A2(n1082), .A3(n1324), .ZN(n1030) );
XNOR2_X1 U1041 ( .A(G952), .B(KEYINPUT63), .ZN(n1324) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1236) );
XNOR2_X1 U1043 ( .A(n1054), .B(KEYINPUT54), .ZN(n1183) );
INV_X1 U1044 ( .A(n1184), .ZN(n1054) );
NAND2_X1 U1045 ( .A1(n1057), .A2(n1056), .ZN(n1184) );
NAND2_X1 U1046 ( .A1(G221), .A2(n1290), .ZN(n1056) );
NAND2_X1 U1047 ( .A1(G234), .A2(n1252), .ZN(n1290) );
XNOR2_X1 U1048 ( .A(n1325), .B(G469), .ZN(n1057) );
NAND3_X1 U1049 ( .A1(n1326), .A2(n1327), .A3(n1252), .ZN(n1325) );
INV_X1 U1050 ( .A(G902), .ZN(n1252) );
OR3_X1 U1051 ( .A1(n1328), .A2(n1329), .A3(KEYINPUT33), .ZN(n1327) );
INV_X1 U1052 ( .A(n1141), .ZN(n1328) );
NAND2_X1 U1053 ( .A1(n1330), .A2(KEYINPUT33), .ZN(n1326) );
XOR2_X1 U1054 ( .A(n1331), .B(n1329), .Z(n1330) );
XOR2_X1 U1055 ( .A(n1332), .B(n1149), .Z(n1329) );
NAND2_X1 U1056 ( .A1(G227), .A2(n1082), .ZN(n1149) );
INV_X1 U1057 ( .A(G953), .ZN(n1082) );
NAND3_X1 U1058 ( .A1(n1333), .A2(n1334), .A3(n1335), .ZN(n1332) );
NAND2_X1 U1059 ( .A1(G140), .A2(n1336), .ZN(n1335) );
OR3_X1 U1060 ( .A1(n1336), .A2(G140), .A3(n1337), .ZN(n1334) );
NAND2_X1 U1061 ( .A1(KEYINPUT51), .A2(n1152), .ZN(n1336) );
INV_X1 U1062 ( .A(G110), .ZN(n1152) );
NAND2_X1 U1063 ( .A1(G110), .A2(n1337), .ZN(n1333) );
INV_X1 U1064 ( .A(KEYINPUT45), .ZN(n1337) );
NOR2_X1 U1065 ( .A1(KEYINPUT38), .A2(n1141), .ZN(n1331) );
XNOR2_X1 U1066 ( .A(n1316), .B(n1338), .ZN(n1141) );
XNOR2_X1 U1067 ( .A(n1339), .B(n1288), .ZN(n1338) );
XNOR2_X1 U1068 ( .A(n1096), .B(n1092), .ZN(n1288) );
XOR2_X1 U1069 ( .A(G134), .B(G137), .Z(n1092) );
INV_X1 U1070 ( .A(G131), .ZN(n1096) );
INV_X1 U1071 ( .A(n1095), .ZN(n1339) );
XOR2_X1 U1072 ( .A(G128), .B(n1340), .Z(n1095) );
NOR2_X1 U1073 ( .A1(KEYINPUT26), .A2(n1341), .ZN(n1340) );
XNOR2_X1 U1074 ( .A(G146), .B(n1342), .ZN(n1341) );
NAND2_X1 U1075 ( .A1(n1343), .A2(KEYINPUT16), .ZN(n1342) );
XNOR2_X1 U1076 ( .A(G143), .B(KEYINPUT41), .ZN(n1343) );
XNOR2_X1 U1077 ( .A(G101), .B(n1344), .ZN(n1316) );
XOR2_X1 U1078 ( .A(G107), .B(G104), .Z(n1344) );
endmodule


