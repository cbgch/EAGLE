//Key = 1001110001110100001100110101101101101010000100110111101110110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369;

XOR2_X1 U759 ( .A(G107), .B(n1045), .Z(G9) );
AND2_X1 U760 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U761 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR3_X1 U762 ( .A1(n1050), .A2(G953), .A3(n1051), .ZN(n1049) );
XOR2_X1 U763 ( .A(KEYINPUT56), .B(n1052), .Z(n1050) );
NOR3_X1 U764 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NOR2_X1 U765 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U766 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U767 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U768 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U769 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U770 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U771 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U772 ( .A1(n1047), .A2(n1070), .ZN(n1068) );
NOR2_X1 U773 ( .A1(n1071), .A2(n1072), .ZN(n1066) );
NOR3_X1 U774 ( .A1(n1073), .A2(n1069), .A3(n1072), .ZN(n1062) );
NOR2_X1 U775 ( .A1(n1074), .A2(n1072), .ZN(n1058) );
NOR2_X1 U776 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U777 ( .A1(n1077), .A2(n1065), .ZN(n1076) );
NOR2_X1 U778 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U779 ( .A1(n1080), .A2(n1069), .ZN(n1079) );
NOR2_X1 U780 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U781 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NOR3_X1 U782 ( .A1(n1085), .A2(n1061), .A3(n1086), .ZN(n1078) );
NOR4_X1 U783 ( .A1(n1087), .A2(n1088), .A3(n1069), .A4(n1061), .ZN(n1075) );
NOR3_X1 U784 ( .A1(n1051), .A2(G953), .A3(G952), .ZN(n1048) );
AND4_X1 U785 ( .A1(n1089), .A2(n1083), .A3(n1090), .A4(n1091), .ZN(n1051) );
NOR4_X1 U786 ( .A1(n1092), .A2(n1093), .A3(n1069), .A4(n1088), .ZN(n1091) );
XNOR2_X1 U787 ( .A(n1084), .B(KEYINPUT22), .ZN(n1093) );
NOR3_X1 U788 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1092) );
AND2_X1 U789 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR3_X1 U790 ( .A1(n1098), .A2(KEYINPUT26), .A3(n1097), .ZN(n1095) );
OR2_X1 U791 ( .A1(n1099), .A2(KEYINPUT57), .ZN(n1097) );
AND2_X1 U792 ( .A1(n1099), .A2(KEYINPUT26), .ZN(n1094) );
NOR3_X1 U793 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1090) );
NOR2_X1 U794 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U795 ( .A(G478), .B(KEYINPUT51), .ZN(n1103) );
NAND2_X1 U796 ( .A1(n1105), .A2(n1106), .ZN(n1089) );
XOR2_X1 U797 ( .A(KEYINPUT20), .B(G475), .Z(n1106) );
XOR2_X1 U798 ( .A(n1107), .B(KEYINPUT60), .Z(n1105) );
XOR2_X1 U799 ( .A(n1108), .B(n1109), .Z(G72) );
XOR2_X1 U800 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U801 ( .A1(n1112), .A2(n1055), .ZN(n1111) );
XNOR2_X1 U802 ( .A(G953), .B(KEYINPUT15), .ZN(n1112) );
NAND2_X1 U803 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
NAND2_X1 U804 ( .A1(n1115), .A2(G900), .ZN(n1114) );
XNOR2_X1 U805 ( .A(G227), .B(KEYINPUT58), .ZN(n1115) );
XNOR2_X1 U806 ( .A(G953), .B(KEYINPUT62), .ZN(n1113) );
NOR3_X1 U807 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1108) );
NOR2_X1 U808 ( .A1(G900), .A2(n1119), .ZN(n1118) );
NOR2_X1 U809 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
XOR2_X1 U810 ( .A(KEYINPUT1), .B(n1122), .Z(n1116) );
AND2_X1 U811 ( .A1(n1121), .A2(n1120), .ZN(n1122) );
XNOR2_X1 U812 ( .A(n1123), .B(n1124), .ZN(n1120) );
XNOR2_X1 U813 ( .A(n1125), .B(n1126), .ZN(n1123) );
XNOR2_X1 U814 ( .A(G140), .B(n1127), .ZN(n1121) );
XOR2_X1 U815 ( .A(n1128), .B(n1129), .Z(G69) );
XOR2_X1 U816 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U817 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NOR2_X1 U818 ( .A1(G898), .A2(n1119), .ZN(n1132) );
NAND3_X1 U819 ( .A1(n1053), .A2(n1119), .A3(KEYINPUT28), .ZN(n1130) );
NAND2_X1 U820 ( .A1(G953), .A2(n1134), .ZN(n1128) );
NAND2_X1 U821 ( .A1(G898), .A2(G224), .ZN(n1134) );
NOR2_X1 U822 ( .A1(n1135), .A2(n1136), .ZN(G66) );
NOR3_X1 U823 ( .A1(n1137), .A2(n1098), .A3(n1138), .ZN(n1136) );
NOR2_X1 U824 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR2_X1 U825 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
NOR2_X1 U826 ( .A1(n1055), .A2(n1053), .ZN(n1141) );
XOR2_X1 U827 ( .A(KEYINPUT41), .B(n1143), .Z(n1137) );
NOR3_X1 U828 ( .A1(n1144), .A2(n1145), .A3(n1142), .ZN(n1143) );
XOR2_X1 U829 ( .A(G217), .B(KEYINPUT9), .Z(n1142) );
XNOR2_X1 U830 ( .A(KEYINPUT8), .B(n1140), .ZN(n1144) );
NOR2_X1 U831 ( .A1(n1135), .A2(n1146), .ZN(G63) );
XOR2_X1 U832 ( .A(n1147), .B(n1148), .Z(n1146) );
NAND2_X1 U833 ( .A1(n1149), .A2(G478), .ZN(n1147) );
NOR2_X1 U834 ( .A1(n1135), .A2(n1150), .ZN(G60) );
XOR2_X1 U835 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U836 ( .A1(n1149), .A2(G475), .ZN(n1151) );
XOR2_X1 U837 ( .A(G104), .B(n1153), .Z(G6) );
NOR2_X1 U838 ( .A1(n1135), .A2(n1154), .ZN(G57) );
NOR2_X1 U839 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U840 ( .A(n1157), .B(KEYINPUT38), .Z(n1156) );
NAND2_X1 U841 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NOR2_X1 U842 ( .A1(n1158), .A2(n1159), .ZN(n1155) );
AND2_X1 U843 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
NAND3_X1 U844 ( .A1(n1149), .A2(G472), .A3(n1162), .ZN(n1161) );
XNOR2_X1 U845 ( .A(n1163), .B(n1164), .ZN(n1162) );
NAND2_X1 U846 ( .A1(n1165), .A2(n1166), .ZN(n1160) );
NAND2_X1 U847 ( .A1(n1149), .A2(G472), .ZN(n1166) );
XOR2_X1 U848 ( .A(n1164), .B(n1163), .Z(n1165) );
NAND2_X1 U849 ( .A1(KEYINPUT0), .A2(n1167), .ZN(n1164) );
NOR2_X1 U850 ( .A1(n1135), .A2(n1168), .ZN(G54) );
XOR2_X1 U851 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U852 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U853 ( .A(n1173), .B(n1174), .Z(n1169) );
XOR2_X1 U854 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U855 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
INV_X1 U856 ( .A(n1179), .ZN(n1178) );
XOR2_X1 U857 ( .A(KEYINPUT27), .B(n1180), .Z(n1177) );
NAND2_X1 U858 ( .A1(n1149), .A2(G469), .ZN(n1173) );
NOR2_X1 U859 ( .A1(n1135), .A2(n1181), .ZN(G51) );
XOR2_X1 U860 ( .A(n1182), .B(n1183), .Z(n1181) );
XNOR2_X1 U861 ( .A(n1184), .B(n1133), .ZN(n1183) );
NAND2_X1 U862 ( .A1(n1149), .A2(n1185), .ZN(n1184) );
INV_X1 U863 ( .A(n1145), .ZN(n1149) );
NAND2_X1 U864 ( .A1(G902), .A2(n1186), .ZN(n1145) );
OR2_X1 U865 ( .A1(n1053), .A2(n1055), .ZN(n1186) );
NAND4_X1 U866 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1055) );
NOR4_X1 U867 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1190) );
NAND2_X1 U868 ( .A1(n1195), .A2(n1196), .ZN(n1189) );
NAND2_X1 U869 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
XNOR2_X1 U870 ( .A(KEYINPUT33), .B(n1199), .ZN(n1197) );
NAND3_X1 U871 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1187) );
NAND2_X1 U872 ( .A1(KEYINPUT31), .A2(n1203), .ZN(n1201) );
NAND2_X1 U873 ( .A1(n1204), .A2(n1205), .ZN(n1200) );
INV_X1 U874 ( .A(KEYINPUT31), .ZN(n1205) );
NAND3_X1 U875 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1204) );
NAND4_X1 U876 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1053) );
NOR4_X1 U877 ( .A1(n1153), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1212) );
NOR3_X1 U878 ( .A1(n1216), .A2(n1073), .A3(n1217), .ZN(n1215) );
NOR4_X1 U879 ( .A1(n1218), .A2(n1219), .A3(n1065), .A4(n1220), .ZN(n1214) );
XNOR2_X1 U880 ( .A(n1082), .B(KEYINPUT6), .ZN(n1218) );
AND2_X1 U881 ( .A1(n1070), .A2(n1046), .ZN(n1153) );
NOR3_X1 U882 ( .A1(n1206), .A2(n1219), .A3(n1065), .ZN(n1046) );
NOR2_X1 U883 ( .A1(n1221), .A2(n1222), .ZN(n1211) );
XOR2_X1 U884 ( .A(n1223), .B(n1224), .Z(n1182) );
NOR2_X1 U885 ( .A1(KEYINPUT63), .A2(n1225), .ZN(n1224) );
NAND3_X1 U886 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1223) );
NAND2_X1 U887 ( .A1(KEYINPUT35), .A2(n1229), .ZN(n1228) );
NAND3_X1 U888 ( .A1(n1230), .A2(n1231), .A3(n1127), .ZN(n1227) );
INV_X1 U889 ( .A(KEYINPUT35), .ZN(n1231) );
OR2_X1 U890 ( .A1(n1127), .A2(n1230), .ZN(n1226) );
NOR2_X1 U891 ( .A1(KEYINPUT48), .A2(n1229), .ZN(n1230) );
NOR2_X1 U892 ( .A1(n1119), .A2(G952), .ZN(n1135) );
XNOR2_X1 U893 ( .A(G146), .B(n1232), .ZN(G48) );
NAND2_X1 U894 ( .A1(n1195), .A2(n1233), .ZN(n1232) );
XNOR2_X1 U895 ( .A(KEYINPUT16), .B(n1198), .ZN(n1233) );
NAND3_X1 U896 ( .A1(n1234), .A2(n1088), .A3(n1235), .ZN(n1198) );
XNOR2_X1 U897 ( .A(G143), .B(n1188), .ZN(G45) );
NAND3_X1 U898 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1188) );
NOR3_X1 U899 ( .A1(n1071), .A2(n1238), .A3(n1239), .ZN(n1237) );
XNOR2_X1 U900 ( .A(n1240), .B(n1194), .ZN(G42) );
NOR3_X1 U901 ( .A1(n1088), .A2(n1241), .A3(n1203), .ZN(n1194) );
XNOR2_X1 U902 ( .A(n1242), .B(n1243), .ZN(G39) );
NOR2_X1 U903 ( .A1(n1244), .A2(n1203), .ZN(n1243) );
XOR2_X1 U904 ( .A(G134), .B(n1193), .Z(G36) );
NOR3_X1 U905 ( .A1(n1073), .A2(n1220), .A3(n1203), .ZN(n1193) );
XOR2_X1 U906 ( .A(G131), .B(n1192), .Z(G33) );
NOR3_X1 U907 ( .A1(n1216), .A2(n1073), .A3(n1203), .ZN(n1192) );
NAND2_X1 U908 ( .A1(n1235), .A2(n1208), .ZN(n1203) );
INV_X1 U909 ( .A(n1069), .ZN(n1208) );
NAND2_X1 U910 ( .A1(n1245), .A2(n1085), .ZN(n1069) );
INV_X1 U911 ( .A(n1086), .ZN(n1245) );
XOR2_X1 U912 ( .A(G128), .B(n1246), .Z(G30) );
NOR2_X1 U913 ( .A1(n1071), .A2(n1199), .ZN(n1246) );
NAND4_X1 U914 ( .A1(n1235), .A2(n1047), .A3(n1088), .A4(n1247), .ZN(n1199) );
INV_X1 U915 ( .A(n1220), .ZN(n1047) );
AND2_X1 U916 ( .A1(n1082), .A2(n1207), .ZN(n1235) );
INV_X1 U917 ( .A(n1206), .ZN(n1082) );
XNOR2_X1 U918 ( .A(G101), .B(n1210), .ZN(G3) );
NAND2_X1 U919 ( .A1(n1236), .A2(n1248), .ZN(n1210) );
XNOR2_X1 U920 ( .A(n1127), .B(n1191), .ZN(G27) );
AND4_X1 U921 ( .A1(n1249), .A2(n1207), .A3(n1195), .A4(n1250), .ZN(n1191) );
NOR2_X1 U922 ( .A1(n1061), .A2(n1241), .ZN(n1250) );
INV_X1 U923 ( .A(n1234), .ZN(n1241) );
NOR2_X1 U924 ( .A1(n1216), .A2(n1087), .ZN(n1234) );
INV_X1 U925 ( .A(n1070), .ZN(n1216) );
NAND2_X1 U926 ( .A1(n1251), .A2(n1057), .ZN(n1207) );
NAND2_X1 U927 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
INV_X1 U928 ( .A(G900), .ZN(n1253) );
XNOR2_X1 U929 ( .A(G122), .B(n1209), .ZN(G24) );
OR4_X1 U930 ( .A1(n1217), .A2(n1065), .A3(n1239), .A4(n1238), .ZN(n1209) );
NAND2_X1 U931 ( .A1(n1087), .A2(n1249), .ZN(n1065) );
XOR2_X1 U932 ( .A(n1213), .B(n1254), .Z(G21) );
NOR2_X1 U933 ( .A1(KEYINPUT2), .A2(n1255), .ZN(n1254) );
INV_X1 U934 ( .A(G119), .ZN(n1255) );
NOR2_X1 U935 ( .A1(n1244), .A2(n1217), .ZN(n1213) );
INV_X1 U936 ( .A(n1202), .ZN(n1244) );
NOR3_X1 U937 ( .A1(n1249), .A2(n1087), .A3(n1072), .ZN(n1202) );
XNOR2_X1 U938 ( .A(n1222), .B(n1256), .ZN(G18) );
NAND2_X1 U939 ( .A1(KEYINPUT52), .A2(G116), .ZN(n1256) );
NOR3_X1 U940 ( .A1(n1073), .A2(n1220), .A3(n1217), .ZN(n1222) );
INV_X1 U941 ( .A(n1257), .ZN(n1217) );
NAND2_X1 U942 ( .A1(n1258), .A2(n1259), .ZN(n1220) );
INV_X1 U943 ( .A(n1236), .ZN(n1073) );
XNOR2_X1 U944 ( .A(G113), .B(n1260), .ZN(G15) );
NAND3_X1 U945 ( .A1(n1070), .A2(n1257), .A3(n1261), .ZN(n1260) );
XNOR2_X1 U946 ( .A(n1236), .B(KEYINPUT3), .ZN(n1261) );
NOR2_X1 U947 ( .A1(n1247), .A2(n1249), .ZN(n1236) );
NOR2_X1 U948 ( .A1(n1061), .A2(n1219), .ZN(n1257) );
NAND2_X1 U949 ( .A1(n1262), .A2(n1263), .ZN(n1061) );
XNOR2_X1 U950 ( .A(n1084), .B(KEYINPUT12), .ZN(n1262) );
NOR2_X1 U951 ( .A1(n1259), .A2(n1239), .ZN(n1070) );
XNOR2_X1 U952 ( .A(n1258), .B(KEYINPUT4), .ZN(n1239) );
INV_X1 U953 ( .A(n1238), .ZN(n1259) );
XNOR2_X1 U954 ( .A(G110), .B(n1264), .ZN(G12) );
NAND2_X1 U955 ( .A1(KEYINPUT50), .A2(n1221), .ZN(n1264) );
AND3_X1 U956 ( .A1(n1249), .A2(n1247), .A3(n1248), .ZN(n1221) );
NOR3_X1 U957 ( .A1(n1206), .A2(n1219), .A3(n1072), .ZN(n1248) );
NAND2_X1 U958 ( .A1(n1238), .A2(n1258), .ZN(n1072) );
NOR2_X1 U959 ( .A1(n1265), .A2(n1101), .ZN(n1258) );
NOR2_X1 U960 ( .A1(n1107), .A2(G475), .ZN(n1101) );
AND2_X1 U961 ( .A1(n1266), .A2(n1107), .ZN(n1265) );
NAND2_X1 U962 ( .A1(n1152), .A2(n1267), .ZN(n1107) );
XNOR2_X1 U963 ( .A(n1268), .B(n1269), .ZN(n1152) );
XOR2_X1 U964 ( .A(G104), .B(n1270), .Z(n1269) );
XOR2_X1 U965 ( .A(KEYINPUT14), .B(G131), .Z(n1270) );
XOR2_X1 U966 ( .A(n1271), .B(n1272), .Z(n1268) );
XOR2_X1 U967 ( .A(n1273), .B(n1274), .Z(n1271) );
NOR2_X1 U968 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
XOR2_X1 U969 ( .A(KEYINPUT32), .B(n1277), .Z(n1276) );
NOR2_X1 U970 ( .A1(G143), .A2(n1278), .ZN(n1277) );
XOR2_X1 U971 ( .A(n1279), .B(KEYINPUT23), .Z(n1278) );
NOR2_X1 U972 ( .A1(n1279), .A2(n1280), .ZN(n1275) );
NAND2_X1 U973 ( .A1(G214), .A2(n1281), .ZN(n1279) );
NAND2_X1 U974 ( .A1(n1282), .A2(KEYINPUT54), .ZN(n1273) );
XOR2_X1 U975 ( .A(n1283), .B(n1284), .Z(n1282) );
NAND2_X1 U976 ( .A1(KEYINPUT46), .A2(n1285), .ZN(n1283) );
XNOR2_X1 U977 ( .A(n1127), .B(n1286), .ZN(n1285) );
NOR2_X1 U978 ( .A1(KEYINPUT39), .A2(n1240), .ZN(n1286) );
XOR2_X1 U979 ( .A(KEYINPUT61), .B(G475), .Z(n1266) );
NOR2_X1 U980 ( .A1(n1100), .A2(n1287), .ZN(n1238) );
NOR2_X1 U981 ( .A1(n1104), .A2(G478), .ZN(n1287) );
AND2_X1 U982 ( .A1(G478), .A2(n1104), .ZN(n1100) );
NAND2_X1 U983 ( .A1(n1148), .A2(n1267), .ZN(n1104) );
XNOR2_X1 U984 ( .A(n1288), .B(n1289), .ZN(n1148) );
XOR2_X1 U985 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U986 ( .A(G128), .B(G122), .Z(n1291) );
XNOR2_X1 U987 ( .A(n1280), .B(G134), .ZN(n1290) );
INV_X1 U988 ( .A(G143), .ZN(n1280) );
XOR2_X1 U989 ( .A(n1292), .B(n1293), .Z(n1288) );
XOR2_X1 U990 ( .A(G116), .B(G107), .Z(n1293) );
NAND2_X1 U991 ( .A1(G217), .A2(n1294), .ZN(n1292) );
NAND2_X1 U992 ( .A1(n1195), .A2(n1295), .ZN(n1219) );
NAND2_X1 U993 ( .A1(n1296), .A2(n1057), .ZN(n1295) );
NAND3_X1 U994 ( .A1(n1297), .A2(n1119), .A3(G952), .ZN(n1057) );
NAND2_X1 U995 ( .A1(n1252), .A2(n1298), .ZN(n1296) );
INV_X1 U996 ( .A(G898), .ZN(n1298) );
AND3_X1 U997 ( .A1(G902), .A2(n1297), .A3(G953), .ZN(n1252) );
NAND2_X1 U998 ( .A1(n1299), .A2(G237), .ZN(n1297) );
XNOR2_X1 U999 ( .A(G234), .B(KEYINPUT25), .ZN(n1299) );
INV_X1 U1000 ( .A(n1071), .ZN(n1195) );
NAND2_X1 U1001 ( .A1(n1086), .A2(n1085), .ZN(n1071) );
NAND2_X1 U1002 ( .A1(G214), .A2(n1300), .ZN(n1085) );
XNOR2_X1 U1003 ( .A(n1301), .B(n1185), .ZN(n1086) );
AND2_X1 U1004 ( .A1(G210), .A2(n1300), .ZN(n1185) );
NAND2_X1 U1005 ( .A1(n1302), .A2(n1267), .ZN(n1300) );
XNOR2_X1 U1006 ( .A(G237), .B(KEYINPUT44), .ZN(n1302) );
NAND2_X1 U1007 ( .A1(n1303), .A2(n1267), .ZN(n1301) );
XOR2_X1 U1008 ( .A(n1304), .B(n1305), .Z(n1303) );
XNOR2_X1 U1009 ( .A(G125), .B(n1225), .ZN(n1305) );
NAND2_X1 U1010 ( .A1(G224), .A2(n1119), .ZN(n1225) );
XOR2_X1 U1011 ( .A(n1133), .B(n1229), .Z(n1304) );
XNOR2_X1 U1012 ( .A(n1306), .B(n1307), .ZN(n1133) );
XOR2_X1 U1013 ( .A(n1308), .B(n1272), .Z(n1307) );
XOR2_X1 U1014 ( .A(G113), .B(G122), .Z(n1272) );
NOR2_X1 U1015 ( .A1(KEYINPUT21), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1016 ( .A(n1310), .B(n1311), .Z(n1306) );
XNOR2_X1 U1017 ( .A(KEYINPUT42), .B(n1312), .ZN(n1311) );
NAND2_X1 U1018 ( .A1(n1313), .A2(n1314), .ZN(n1310) );
OR2_X1 U1019 ( .A1(n1315), .A2(G101), .ZN(n1314) );
XOR2_X1 U1020 ( .A(n1316), .B(KEYINPUT24), .Z(n1313) );
NAND2_X1 U1021 ( .A1(G101), .A2(n1315), .ZN(n1316) );
NAND2_X1 U1022 ( .A1(n1084), .A2(n1263), .ZN(n1206) );
XNOR2_X1 U1023 ( .A(n1083), .B(KEYINPUT5), .ZN(n1263) );
NAND2_X1 U1024 ( .A1(G221), .A2(n1317), .ZN(n1083) );
XNOR2_X1 U1025 ( .A(n1318), .B(n1319), .ZN(n1084) );
XOR2_X1 U1026 ( .A(KEYINPUT29), .B(G469), .Z(n1319) );
NAND3_X1 U1027 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1318) );
XNOR2_X1 U1028 ( .A(KEYINPUT34), .B(n1267), .ZN(n1322) );
NAND2_X1 U1029 ( .A1(n1323), .A2(n1324), .ZN(n1321) );
INV_X1 U1030 ( .A(KEYINPUT53), .ZN(n1324) );
XOR2_X1 U1031 ( .A(n1325), .B(n1326), .Z(n1323) );
NAND2_X1 U1032 ( .A1(KEYINPUT55), .A2(n1327), .ZN(n1325) );
INV_X1 U1033 ( .A(n1328), .ZN(n1327) );
NAND3_X1 U1034 ( .A1(n1326), .A2(n1328), .A3(KEYINPUT53), .ZN(n1320) );
XNOR2_X1 U1035 ( .A(n1329), .B(n1330), .ZN(n1328) );
NOR2_X1 U1036 ( .A1(n1179), .A2(n1180), .ZN(n1330) );
AND2_X1 U1037 ( .A1(n1126), .A2(n1331), .ZN(n1180) );
NOR2_X1 U1038 ( .A1(n1331), .A2(n1126), .ZN(n1179) );
XNOR2_X1 U1039 ( .A(n1332), .B(n1333), .ZN(n1126) );
XNOR2_X1 U1040 ( .A(G128), .B(KEYINPUT7), .ZN(n1332) );
XOR2_X1 U1041 ( .A(G101), .B(n1334), .Z(n1331) );
NOR2_X1 U1042 ( .A1(KEYINPUT17), .A2(n1335), .ZN(n1334) );
INV_X1 U1043 ( .A(n1315), .ZN(n1335) );
XOR2_X1 U1044 ( .A(G104), .B(G107), .Z(n1315) );
NAND2_X1 U1045 ( .A1(KEYINPUT36), .A2(n1336), .ZN(n1329) );
XOR2_X1 U1046 ( .A(KEYINPUT40), .B(n1171), .Z(n1336) );
XOR2_X1 U1047 ( .A(n1176), .B(n1337), .Z(n1326) );
NOR2_X1 U1048 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
NOR3_X1 U1049 ( .A1(KEYINPUT49), .A2(G110), .A3(n1240), .ZN(n1339) );
INV_X1 U1050 ( .A(G140), .ZN(n1240) );
NOR2_X1 U1051 ( .A1(n1172), .A2(n1340), .ZN(n1338) );
INV_X1 U1052 ( .A(KEYINPUT49), .ZN(n1340) );
XNOR2_X1 U1053 ( .A(n1312), .B(G140), .ZN(n1172) );
AND2_X1 U1054 ( .A1(G227), .A2(n1119), .ZN(n1176) );
INV_X1 U1055 ( .A(n1087), .ZN(n1247) );
XNOR2_X1 U1056 ( .A(n1098), .B(n1099), .ZN(n1087) );
AND2_X1 U1057 ( .A1(G217), .A2(n1317), .ZN(n1099) );
NAND2_X1 U1058 ( .A1(G234), .A2(n1267), .ZN(n1317) );
NOR2_X1 U1059 ( .A1(n1140), .A2(G902), .ZN(n1098) );
XOR2_X1 U1060 ( .A(n1341), .B(n1342), .Z(n1140) );
XOR2_X1 U1061 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1062 ( .A(G137), .B(n1345), .ZN(n1344) );
NAND3_X1 U1063 ( .A1(n1346), .A2(n1347), .A3(KEYINPUT10), .ZN(n1345) );
NAND2_X1 U1064 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
NAND2_X1 U1065 ( .A1(G110), .A2(n1350), .ZN(n1349) );
NAND2_X1 U1066 ( .A1(KEYINPUT18), .A2(n1351), .ZN(n1350) );
INV_X1 U1067 ( .A(KEYINPUT43), .ZN(n1351) );
NAND3_X1 U1068 ( .A1(n1352), .A2(n1353), .A3(KEYINPUT43), .ZN(n1346) );
OR2_X1 U1069 ( .A1(n1312), .A2(KEYINPUT18), .ZN(n1353) );
NAND2_X1 U1070 ( .A1(KEYINPUT18), .A2(n1354), .ZN(n1352) );
OR2_X1 U1071 ( .A1(n1348), .A2(n1312), .ZN(n1354) );
INV_X1 U1072 ( .A(G110), .ZN(n1312) );
XOR2_X1 U1073 ( .A(G119), .B(n1355), .Z(n1348) );
NOR2_X1 U1074 ( .A1(KEYINPUT45), .A2(G128), .ZN(n1355) );
AND2_X1 U1075 ( .A1(n1294), .A2(G221), .ZN(n1343) );
AND2_X1 U1076 ( .A1(G234), .A2(n1119), .ZN(n1294) );
INV_X1 U1077 ( .A(G953), .ZN(n1119) );
XOR2_X1 U1078 ( .A(n1356), .B(n1284), .Z(n1341) );
XNOR2_X1 U1079 ( .A(n1357), .B(KEYINPUT59), .ZN(n1284) );
INV_X1 U1080 ( .A(G146), .ZN(n1357) );
NAND2_X1 U1081 ( .A1(n1358), .A2(n1359), .ZN(n1356) );
NAND2_X1 U1082 ( .A1(G140), .A2(n1127), .ZN(n1359) );
XOR2_X1 U1083 ( .A(KEYINPUT47), .B(n1360), .Z(n1358) );
NOR2_X1 U1084 ( .A1(G140), .A2(n1127), .ZN(n1360) );
INV_X1 U1085 ( .A(G125), .ZN(n1127) );
INV_X1 U1086 ( .A(n1088), .ZN(n1249) );
XNOR2_X1 U1087 ( .A(n1361), .B(G472), .ZN(n1088) );
NAND2_X1 U1088 ( .A1(n1362), .A2(n1267), .ZN(n1361) );
INV_X1 U1089 ( .A(G902), .ZN(n1267) );
XNOR2_X1 U1090 ( .A(n1363), .B(n1167), .ZN(n1362) );
XNOR2_X1 U1091 ( .A(n1364), .B(n1309), .ZN(n1167) );
XNOR2_X1 U1092 ( .A(G116), .B(G119), .ZN(n1309) );
XNOR2_X1 U1093 ( .A(G113), .B(KEYINPUT42), .ZN(n1364) );
XNOR2_X1 U1094 ( .A(n1365), .B(n1159), .ZN(n1363) );
XOR2_X1 U1095 ( .A(n1366), .B(G101), .Z(n1159) );
NAND2_X1 U1096 ( .A1(G210), .A2(n1281), .ZN(n1366) );
NOR2_X1 U1097 ( .A1(G953), .A2(G237), .ZN(n1281) );
NAND2_X1 U1098 ( .A1(KEYINPUT11), .A2(n1163), .ZN(n1365) );
XOR2_X1 U1099 ( .A(n1171), .B(n1229), .Z(n1163) );
XNOR2_X1 U1100 ( .A(n1333), .B(n1367), .ZN(n1229) );
NOR2_X1 U1101 ( .A1(G128), .A2(KEYINPUT37), .ZN(n1367) );
XOR2_X1 U1102 ( .A(G146), .B(G143), .Z(n1333) );
XNOR2_X1 U1103 ( .A(n1368), .B(n1125), .ZN(n1171) );
XOR2_X1 U1104 ( .A(G131), .B(n1369), .Z(n1125) );
XNOR2_X1 U1105 ( .A(KEYINPUT30), .B(n1242), .ZN(n1369) );
INV_X1 U1106 ( .A(G137), .ZN(n1242) );
NAND2_X1 U1107 ( .A1(KEYINPUT13), .A2(n1124), .ZN(n1368) );
XNOR2_X1 U1108 ( .A(G134), .B(KEYINPUT19), .ZN(n1124) );
endmodule


