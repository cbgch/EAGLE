//Key = 1011010010000010001010010001101001101110000011100000100011010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400;

XNOR2_X1 U781 ( .A(n1073), .B(n1074), .ZN(G9) );
NOR2_X1 U782 ( .A1(n1075), .A2(n1076), .ZN(G75) );
NOR4_X1 U783 ( .A1(n1077), .A2(n1078), .A3(G953), .A4(n1079), .ZN(n1076) );
AND4_X1 U784 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1078) );
NAND3_X1 U785 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1077) );
XOR2_X1 U786 ( .A(n1087), .B(KEYINPUT28), .Z(n1086) );
NAND2_X1 U787 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U788 ( .A1(n1082), .A2(n1090), .A3(n1091), .ZN(n1089) );
NAND2_X1 U789 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NAND4_X1 U790 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1081), .ZN(n1093) );
NAND2_X1 U791 ( .A1(n1097), .A2(n1098), .ZN(n1092) );
NAND2_X1 U792 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND4_X1 U793 ( .A1(KEYINPUT59), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1100) );
NAND2_X1 U794 ( .A1(n1095), .A2(n1104), .ZN(n1099) );
NAND2_X1 U795 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U796 ( .A1(n1102), .A2(n1107), .ZN(n1106) );
INV_X1 U797 ( .A(KEYINPUT59), .ZN(n1107) );
XNOR2_X1 U798 ( .A(n1081), .B(KEYINPUT8), .ZN(n1102) );
NAND4_X1 U799 ( .A1(n1083), .A2(n1095), .A3(n1108), .A4(n1081), .ZN(n1088) );
NAND2_X1 U800 ( .A1(n1095), .A2(n1109), .ZN(n1085) );
NAND3_X1 U801 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
NAND2_X1 U802 ( .A1(KEYINPUT29), .A2(n1113), .ZN(n1112) );
NAND2_X1 U803 ( .A1(n1083), .A2(n1114), .ZN(n1113) );
NAND3_X1 U804 ( .A1(n1115), .A2(n1081), .A3(n1083), .ZN(n1111) );
NOR2_X1 U805 ( .A1(n1116), .A2(n1117), .ZN(n1083) );
NAND3_X1 U806 ( .A1(n1082), .A2(n1118), .A3(n1091), .ZN(n1110) );
INV_X1 U807 ( .A(n1116), .ZN(n1091) );
NAND2_X1 U808 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
OR3_X1 U809 ( .A1(n1117), .A2(KEYINPUT29), .A3(n1121), .ZN(n1120) );
NAND2_X1 U810 ( .A1(n1081), .A2(n1122), .ZN(n1119) );
NOR3_X1 U811 ( .A1(n1079), .A2(G953), .A3(G952), .ZN(n1075) );
AND4_X1 U812 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n1079) );
NOR4_X1 U813 ( .A1(n1101), .A2(n1127), .A3(n1117), .A4(n1128), .ZN(n1126) );
XNOR2_X1 U814 ( .A(n1129), .B(KEYINPUT52), .ZN(n1127) );
XOR2_X1 U815 ( .A(n1130), .B(G472), .Z(n1125) );
XOR2_X1 U816 ( .A(n1131), .B(n1132), .Z(n1124) );
XNOR2_X1 U817 ( .A(G475), .B(n1133), .ZN(n1123) );
NOR2_X1 U818 ( .A1(KEYINPUT48), .A2(n1134), .ZN(n1133) );
XOR2_X1 U819 ( .A(n1135), .B(n1136), .Z(G72) );
XOR2_X1 U820 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U821 ( .A1(n1139), .A2(KEYINPUT6), .ZN(n1138) );
NOR4_X1 U822 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1139) );
NOR2_X1 U823 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NOR2_X1 U824 ( .A1(KEYINPUT35), .A2(n1146), .ZN(n1144) );
XNOR2_X1 U825 ( .A(n1147), .B(KEYINPUT60), .ZN(n1146) );
NOR2_X1 U826 ( .A1(n1148), .A2(n1149), .ZN(n1142) );
XOR2_X1 U827 ( .A(KEYINPUT49), .B(G900), .Z(n1149) );
NOR2_X1 U828 ( .A1(n1147), .A2(n1150), .ZN(n1141) );
AND3_X1 U829 ( .A1(n1150), .A2(n1145), .A3(n1147), .ZN(n1140) );
XNOR2_X1 U830 ( .A(n1151), .B(n1152), .ZN(n1147) );
XNOR2_X1 U831 ( .A(n1153), .B(n1154), .ZN(n1151) );
NAND2_X1 U832 ( .A1(KEYINPUT36), .A2(n1155), .ZN(n1153) );
NAND2_X1 U833 ( .A1(n1156), .A2(n1157), .ZN(n1145) );
NAND2_X1 U834 ( .A1(G125), .A2(n1158), .ZN(n1157) );
XOR2_X1 U835 ( .A(KEYINPUT56), .B(n1159), .Z(n1156) );
NOR2_X1 U836 ( .A1(G125), .A2(n1158), .ZN(n1159) );
INV_X1 U837 ( .A(KEYINPUT35), .ZN(n1150) );
NOR2_X1 U838 ( .A1(n1160), .A2(G953), .ZN(n1137) );
NOR2_X1 U839 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XNOR2_X1 U840 ( .A(n1163), .B(KEYINPUT57), .ZN(n1161) );
NAND2_X1 U841 ( .A1(G953), .A2(n1164), .ZN(n1135) );
NAND2_X1 U842 ( .A1(G900), .A2(G227), .ZN(n1164) );
XOR2_X1 U843 ( .A(n1165), .B(n1166), .Z(G69) );
XOR2_X1 U844 ( .A(n1167), .B(n1168), .Z(n1166) );
NAND2_X1 U845 ( .A1(G953), .A2(n1169), .ZN(n1168) );
NAND2_X1 U846 ( .A1(G898), .A2(G224), .ZN(n1169) );
NAND2_X1 U847 ( .A1(n1170), .A2(n1171), .ZN(n1167) );
NAND2_X1 U848 ( .A1(G953), .A2(n1172), .ZN(n1171) );
XOR2_X1 U849 ( .A(n1173), .B(n1174), .Z(n1170) );
NAND2_X1 U850 ( .A1(KEYINPUT34), .A2(n1175), .ZN(n1174) );
NAND2_X1 U851 ( .A1(n1176), .A2(n1177), .ZN(n1173) );
NAND2_X1 U852 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XOR2_X1 U853 ( .A(n1180), .B(KEYINPUT39), .Z(n1176) );
OR2_X1 U854 ( .A1(n1179), .A2(n1178), .ZN(n1180) );
AND2_X1 U855 ( .A1(n1181), .A2(n1148), .ZN(n1165) );
NOR2_X1 U856 ( .A1(n1182), .A2(n1183), .ZN(G66) );
XOR2_X1 U857 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U858 ( .A1(n1186), .A2(KEYINPUT9), .ZN(n1185) );
NOR2_X1 U859 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
INV_X1 U860 ( .A(n1189), .ZN(n1188) );
NOR2_X1 U861 ( .A1(n1182), .A2(n1190), .ZN(G63) );
NOR2_X1 U862 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U863 ( .A(KEYINPUT24), .B(n1193), .Z(n1192) );
AND2_X1 U864 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NOR2_X1 U865 ( .A1(n1195), .A2(n1194), .ZN(n1191) );
NAND3_X1 U866 ( .A1(n1196), .A2(n1197), .A3(G478), .ZN(n1194) );
INV_X1 U867 ( .A(n1084), .ZN(n1197) );
XNOR2_X1 U868 ( .A(KEYINPUT53), .B(n1198), .ZN(n1196) );
NOR2_X1 U869 ( .A1(n1182), .A2(n1199), .ZN(G60) );
XOR2_X1 U870 ( .A(n1200), .B(n1201), .Z(n1199) );
NAND2_X1 U871 ( .A1(n1189), .A2(G475), .ZN(n1200) );
XNOR2_X1 U872 ( .A(n1202), .B(n1203), .ZN(G6) );
NOR2_X1 U873 ( .A1(n1182), .A2(n1204), .ZN(G57) );
XOR2_X1 U874 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U875 ( .A(n1207), .B(n1208), .Z(n1206) );
NAND2_X1 U876 ( .A1(n1189), .A2(G472), .ZN(n1207) );
XOR2_X1 U877 ( .A(n1209), .B(n1210), .Z(n1205) );
NOR2_X1 U878 ( .A1(KEYINPUT42), .A2(n1211), .ZN(n1210) );
NOR2_X1 U879 ( .A1(KEYINPUT16), .A2(n1212), .ZN(n1209) );
NOR3_X1 U880 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(G54) );
AND2_X1 U881 ( .A1(KEYINPUT62), .A2(n1182), .ZN(n1215) );
NOR3_X1 U882 ( .A1(KEYINPUT62), .A2(n1148), .A3(n1216), .ZN(n1214) );
INV_X1 U883 ( .A(G952), .ZN(n1216) );
XOR2_X1 U884 ( .A(n1217), .B(n1218), .Z(n1213) );
NOR2_X1 U885 ( .A1(KEYINPUT19), .A2(n1219), .ZN(n1218) );
XOR2_X1 U886 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U887 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR2_X1 U888 ( .A1(KEYINPUT12), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U889 ( .A(n1225), .B(n1226), .ZN(n1220) );
NAND2_X1 U890 ( .A1(n1227), .A2(n1228), .ZN(n1225) );
NAND2_X1 U891 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NAND2_X1 U892 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
OR2_X1 U893 ( .A1(KEYINPUT10), .A2(KEYINPUT45), .ZN(n1232) );
NAND3_X1 U894 ( .A1(n1233), .A2(n1234), .A3(KEYINPUT45), .ZN(n1227) );
NAND2_X1 U895 ( .A1(n1231), .A2(n1235), .ZN(n1234) );
OR2_X1 U896 ( .A1(n1229), .A2(KEYINPUT10), .ZN(n1235) );
OR2_X1 U897 ( .A1(n1231), .A2(KEYINPUT10), .ZN(n1233) );
NAND2_X1 U898 ( .A1(n1189), .A2(G469), .ZN(n1217) );
NOR2_X1 U899 ( .A1(n1182), .A2(n1236), .ZN(G51) );
XOR2_X1 U900 ( .A(n1237), .B(n1238), .Z(n1236) );
NOR2_X1 U901 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
NAND2_X1 U902 ( .A1(n1189), .A2(n1132), .ZN(n1237) );
NOR2_X1 U903 ( .A1(n1198), .A2(n1084), .ZN(n1189) );
NOR3_X1 U904 ( .A1(n1162), .A2(n1163), .A3(n1181), .ZN(n1084) );
NAND4_X1 U905 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1181) );
NOR4_X1 U906 ( .A1(n1245), .A2(n1074), .A3(n1246), .A4(n1203), .ZN(n1244) );
AND3_X1 U907 ( .A1(n1247), .A2(n1081), .A3(n1115), .ZN(n1203) );
NOR4_X1 U908 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1246) );
XOR2_X1 U909 ( .A(KEYINPUT18), .B(n1122), .Z(n1251) );
XNOR2_X1 U910 ( .A(n1080), .B(KEYINPUT26), .ZN(n1249) );
INV_X1 U911 ( .A(n1252), .ZN(n1248) );
AND3_X1 U912 ( .A1(n1247), .A2(n1081), .A3(n1108), .ZN(n1074) );
NOR3_X1 U913 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1243) );
NOR4_X1 U914 ( .A1(n1256), .A2(n1105), .A3(n1082), .A4(n1257), .ZN(n1255) );
AND2_X1 U915 ( .A1(n1256), .A2(n1258), .ZN(n1254) );
INV_X1 U916 ( .A(KEYINPUT50), .ZN(n1256) );
INV_X1 U917 ( .A(n1259), .ZN(n1163) );
NAND4_X1 U918 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(n1162) );
NOR3_X1 U919 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1263) );
INV_X1 U920 ( .A(n1267), .ZN(n1266) );
NAND2_X1 U921 ( .A1(n1268), .A2(n1269), .ZN(n1262) );
NAND2_X1 U922 ( .A1(n1270), .A2(n1105), .ZN(n1269) );
XNOR2_X1 U923 ( .A(n1271), .B(KEYINPUT55), .ZN(n1270) );
INV_X1 U924 ( .A(n1272), .ZN(n1268) );
NAND2_X1 U925 ( .A1(n1095), .A2(n1273), .ZN(n1260) );
XNOR2_X1 U926 ( .A(KEYINPUT4), .B(n1274), .ZN(n1273) );
NOR2_X1 U927 ( .A1(n1148), .A2(G952), .ZN(n1182) );
XOR2_X1 U928 ( .A(G146), .B(n1265), .Z(G48) );
AND3_X1 U929 ( .A1(n1115), .A2(n1080), .A3(n1275), .ZN(n1265) );
XNOR2_X1 U930 ( .A(G143), .B(n1261), .ZN(G45) );
NAND4_X1 U931 ( .A1(n1276), .A2(n1080), .A3(n1129), .A4(n1277), .ZN(n1261) );
XNOR2_X1 U932 ( .A(n1158), .B(n1278), .ZN(G42) );
NOR2_X1 U933 ( .A1(n1105), .A2(n1272), .ZN(n1278) );
XNOR2_X1 U934 ( .A(n1259), .B(n1279), .ZN(G39) );
NOR2_X1 U935 ( .A1(KEYINPUT63), .A2(n1280), .ZN(n1279) );
INV_X1 U936 ( .A(G137), .ZN(n1280) );
NAND3_X1 U937 ( .A1(n1095), .A2(n1082), .A3(n1275), .ZN(n1259) );
XNOR2_X1 U938 ( .A(n1281), .B(n1282), .ZN(G36) );
NOR2_X1 U939 ( .A1(n1283), .A2(n1274), .ZN(n1282) );
NAND2_X1 U940 ( .A1(n1276), .A2(n1108), .ZN(n1274) );
AND3_X1 U941 ( .A1(n1122), .A2(n1284), .A3(n1271), .ZN(n1276) );
XOR2_X1 U942 ( .A(G131), .B(n1285), .Z(G33) );
NOR2_X1 U943 ( .A1(n1121), .A2(n1272), .ZN(n1285) );
NAND4_X1 U944 ( .A1(n1095), .A2(n1115), .A3(n1122), .A4(n1284), .ZN(n1272) );
INV_X1 U945 ( .A(n1283), .ZN(n1095) );
NAND2_X1 U946 ( .A1(n1103), .A2(n1286), .ZN(n1283) );
INV_X1 U947 ( .A(n1271), .ZN(n1121) );
XOR2_X1 U948 ( .A(G128), .B(n1264), .Z(G30) );
AND3_X1 U949 ( .A1(n1108), .A2(n1080), .A3(n1275), .ZN(n1264) );
AND4_X1 U950 ( .A1(n1287), .A2(n1122), .A3(n1128), .A4(n1284), .ZN(n1275) );
XNOR2_X1 U951 ( .A(G101), .B(n1288), .ZN(G3) );
NAND2_X1 U952 ( .A1(n1114), .A2(n1247), .ZN(n1288) );
INV_X1 U953 ( .A(n1250), .ZN(n1114) );
NAND2_X1 U954 ( .A1(n1082), .A2(n1271), .ZN(n1250) );
XNOR2_X1 U955 ( .A(G125), .B(n1267), .ZN(G27) );
NAND3_X1 U956 ( .A1(n1289), .A2(n1115), .A3(n1290), .ZN(n1267) );
AND3_X1 U957 ( .A1(n1097), .A2(n1284), .A3(n1080), .ZN(n1290) );
NAND2_X1 U958 ( .A1(n1116), .A2(n1291), .ZN(n1284) );
NAND4_X1 U959 ( .A1(n1292), .A2(G953), .A3(G902), .A4(n1293), .ZN(n1291) );
XNOR2_X1 U960 ( .A(G900), .B(KEYINPUT49), .ZN(n1292) );
XOR2_X1 U961 ( .A(G122), .B(n1245), .Z(G24) );
AND4_X1 U962 ( .A1(n1294), .A2(n1081), .A3(n1129), .A4(n1277), .ZN(n1245) );
NOR2_X1 U963 ( .A1(n1128), .A2(n1287), .ZN(n1081) );
XOR2_X1 U964 ( .A(n1241), .B(n1295), .Z(G21) );
XNOR2_X1 U965 ( .A(KEYINPUT14), .B(n1296), .ZN(n1295) );
NAND4_X1 U966 ( .A1(n1287), .A2(n1082), .A3(n1294), .A4(n1128), .ZN(n1241) );
INV_X1 U967 ( .A(n1297), .ZN(n1287) );
NAND2_X1 U968 ( .A1(n1298), .A2(n1299), .ZN(G18) );
NAND2_X1 U969 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
XOR2_X1 U970 ( .A(KEYINPUT37), .B(n1302), .Z(n1298) );
NOR2_X1 U971 ( .A1(n1301), .A2(n1300), .ZN(n1302) );
NAND2_X1 U972 ( .A1(n1303), .A2(n1304), .ZN(n1300) );
NAND2_X1 U973 ( .A1(n1253), .A2(n1305), .ZN(n1304) );
INV_X1 U974 ( .A(KEYINPUT15), .ZN(n1305) );
AND2_X1 U975 ( .A1(n1306), .A2(n1108), .ZN(n1253) );
NAND3_X1 U976 ( .A1(n1306), .A2(n1307), .A3(KEYINPUT15), .ZN(n1303) );
INV_X1 U977 ( .A(n1108), .ZN(n1307) );
NOR2_X1 U978 ( .A1(n1277), .A2(n1308), .ZN(n1108) );
XOR2_X1 U979 ( .A(n1242), .B(n1309), .Z(G15) );
NAND2_X1 U980 ( .A1(KEYINPUT38), .A2(G113), .ZN(n1309) );
NAND2_X1 U981 ( .A1(n1306), .A2(n1115), .ZN(n1242) );
AND2_X1 U982 ( .A1(n1308), .A2(n1277), .ZN(n1115) );
INV_X1 U983 ( .A(n1129), .ZN(n1308) );
AND2_X1 U984 ( .A1(n1271), .A2(n1294), .ZN(n1306) );
AND3_X1 U985 ( .A1(n1080), .A2(n1252), .A3(n1097), .ZN(n1294) );
INV_X1 U986 ( .A(n1117), .ZN(n1097) );
NAND2_X1 U987 ( .A1(n1096), .A2(n1310), .ZN(n1117) );
NOR2_X1 U988 ( .A1(n1297), .A2(n1128), .ZN(n1271) );
XOR2_X1 U989 ( .A(n1311), .B(n1258), .Z(G12) );
AND3_X1 U990 ( .A1(n1082), .A2(n1247), .A3(n1289), .ZN(n1258) );
INV_X1 U991 ( .A(n1105), .ZN(n1289) );
NAND2_X1 U992 ( .A1(n1128), .A2(n1297), .ZN(n1105) );
XNOR2_X1 U993 ( .A(n1312), .B(G472), .ZN(n1297) );
NAND2_X1 U994 ( .A1(n1313), .A2(KEYINPUT2), .ZN(n1312) );
XOR2_X1 U995 ( .A(n1130), .B(KEYINPUT43), .Z(n1313) );
NAND2_X1 U996 ( .A1(n1314), .A2(n1198), .ZN(n1130) );
XOR2_X1 U997 ( .A(n1315), .B(n1212), .Z(n1314) );
AND2_X1 U998 ( .A1(n1316), .A2(n1317), .ZN(n1212) );
NAND2_X1 U999 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
INV_X1 U1000 ( .A(G101), .ZN(n1319) );
NAND3_X1 U1001 ( .A1(n1320), .A2(n1148), .A3(G210), .ZN(n1318) );
NAND4_X1 U1002 ( .A1(n1320), .A2(n1148), .A3(G210), .A4(G101), .ZN(n1316) );
XOR2_X1 U1003 ( .A(n1208), .B(n1211), .Z(n1315) );
XOR2_X1 U1004 ( .A(n1321), .B(n1322), .Z(n1208) );
XNOR2_X1 U1005 ( .A(n1301), .B(n1323), .ZN(n1322) );
NOR2_X1 U1006 ( .A1(KEYINPUT40), .A2(n1296), .ZN(n1323) );
XNOR2_X1 U1007 ( .A(n1222), .B(n1324), .ZN(n1321) );
XOR2_X1 U1008 ( .A(n1325), .B(n1187), .Z(n1128) );
NAND2_X1 U1009 ( .A1(G217), .A2(n1326), .ZN(n1187) );
NAND2_X1 U1010 ( .A1(n1184), .A2(n1198), .ZN(n1325) );
XOR2_X1 U1011 ( .A(n1327), .B(n1328), .Z(n1184) );
XOR2_X1 U1012 ( .A(n1329), .B(n1330), .Z(n1328) );
NAND3_X1 U1013 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(n1329) );
NAND2_X1 U1014 ( .A1(KEYINPUT47), .A2(n1334), .ZN(n1333) );
OR4_X1 U1015 ( .A1(n1335), .A2(KEYINPUT47), .A3(n1334), .A4(n1336), .ZN(n1332) );
NAND2_X1 U1016 ( .A1(G221), .A2(n1337), .ZN(n1334) );
INV_X1 U1017 ( .A(KEYINPUT0), .ZN(n1335) );
NAND2_X1 U1018 ( .A1(n1336), .A2(n1338), .ZN(n1331) );
NAND3_X1 U1019 ( .A1(G221), .A2(n1337), .A3(KEYINPUT0), .ZN(n1338) );
XNOR2_X1 U1020 ( .A(n1155), .B(KEYINPUT25), .ZN(n1336) );
XNOR2_X1 U1021 ( .A(n1339), .B(n1340), .ZN(n1327) );
NOR2_X1 U1022 ( .A1(G125), .A2(KEYINPUT54), .ZN(n1340) );
NOR2_X1 U1023 ( .A1(KEYINPUT7), .A2(n1341), .ZN(n1339) );
XNOR2_X1 U1024 ( .A(n1342), .B(n1343), .ZN(n1341) );
XNOR2_X1 U1025 ( .A(G128), .B(n1296), .ZN(n1343) );
INV_X1 U1026 ( .A(n1257), .ZN(n1247) );
NAND3_X1 U1027 ( .A1(n1080), .A2(n1252), .A3(n1122), .ZN(n1257) );
NOR2_X1 U1028 ( .A1(n1096), .A2(n1094), .ZN(n1122) );
INV_X1 U1029 ( .A(n1310), .ZN(n1094) );
NAND2_X1 U1030 ( .A1(G221), .A2(n1326), .ZN(n1310) );
NAND2_X1 U1031 ( .A1(G234), .A2(n1198), .ZN(n1326) );
XOR2_X1 U1032 ( .A(n1344), .B(G469), .Z(n1096) );
NAND2_X1 U1033 ( .A1(n1345), .A2(n1198), .ZN(n1344) );
XOR2_X1 U1034 ( .A(n1346), .B(n1347), .Z(n1345) );
XOR2_X1 U1035 ( .A(n1222), .B(n1348), .Z(n1347) );
XNOR2_X1 U1036 ( .A(KEYINPUT23), .B(n1349), .ZN(n1348) );
NOR2_X1 U1037 ( .A1(KEYINPUT17), .A2(n1350), .ZN(n1349) );
XNOR2_X1 U1038 ( .A(n1226), .B(n1224), .ZN(n1350) );
XNOR2_X1 U1039 ( .A(n1342), .B(n1158), .ZN(n1224) );
INV_X1 U1040 ( .A(G140), .ZN(n1158) );
NAND2_X1 U1041 ( .A1(G227), .A2(n1148), .ZN(n1226) );
XNOR2_X1 U1042 ( .A(n1155), .B(n1351), .ZN(n1222) );
XOR2_X1 U1043 ( .A(KEYINPUT31), .B(n1152), .Z(n1351) );
XNOR2_X1 U1044 ( .A(n1281), .B(G131), .ZN(n1152) );
INV_X1 U1045 ( .A(G134), .ZN(n1281) );
XOR2_X1 U1046 ( .A(G137), .B(KEYINPUT20), .Z(n1155) );
XNOR2_X1 U1047 ( .A(n1229), .B(n1231), .ZN(n1346) );
XOR2_X1 U1048 ( .A(n1352), .B(KEYINPUT3), .Z(n1231) );
XOR2_X1 U1049 ( .A(G107), .B(n1353), .Z(n1229) );
NAND2_X1 U1050 ( .A1(n1116), .A2(n1354), .ZN(n1252) );
NAND4_X1 U1051 ( .A1(G953), .A2(G902), .A3(n1293), .A4(n1172), .ZN(n1354) );
INV_X1 U1052 ( .A(G898), .ZN(n1172) );
NAND3_X1 U1053 ( .A1(n1293), .A2(n1148), .A3(G952), .ZN(n1116) );
NAND2_X1 U1054 ( .A1(G237), .A2(G234), .ZN(n1293) );
NOR2_X1 U1055 ( .A1(n1103), .A2(n1101), .ZN(n1080) );
INV_X1 U1056 ( .A(n1286), .ZN(n1101) );
NAND2_X1 U1057 ( .A1(G214), .A2(n1355), .ZN(n1286) );
XNOR2_X1 U1058 ( .A(n1356), .B(n1132), .ZN(n1103) );
AND2_X1 U1059 ( .A1(G210), .A2(n1355), .ZN(n1132) );
NAND2_X1 U1060 ( .A1(n1320), .A2(n1198), .ZN(n1355) );
INV_X1 U1061 ( .A(G237), .ZN(n1320) );
NAND2_X1 U1062 ( .A1(KEYINPUT27), .A2(n1131), .ZN(n1356) );
NAND3_X1 U1063 ( .A1(n1357), .A2(n1198), .A3(n1358), .ZN(n1131) );
XNOR2_X1 U1064 ( .A(n1239), .B(KEYINPUT51), .ZN(n1358) );
AND2_X1 U1065 ( .A1(n1359), .A2(n1360), .ZN(n1239) );
INV_X1 U1066 ( .A(n1240), .ZN(n1357) );
NOR2_X1 U1067 ( .A1(n1360), .A2(n1359), .ZN(n1240) );
XOR2_X1 U1068 ( .A(n1361), .B(n1179), .Z(n1359) );
NAND2_X1 U1069 ( .A1(n1362), .A2(n1363), .ZN(n1179) );
NAND2_X1 U1070 ( .A1(n1364), .A2(n1073), .ZN(n1363) );
INV_X1 U1071 ( .A(G107), .ZN(n1073) );
XOR2_X1 U1072 ( .A(KEYINPUT46), .B(n1353), .Z(n1364) );
NAND2_X1 U1073 ( .A1(n1353), .A2(G107), .ZN(n1362) );
XNOR2_X1 U1074 ( .A(n1202), .B(G101), .ZN(n1353) );
INV_X1 U1075 ( .A(G104), .ZN(n1202) );
XNOR2_X1 U1076 ( .A(n1178), .B(n1175), .ZN(n1361) );
XNOR2_X1 U1077 ( .A(n1342), .B(n1365), .ZN(n1175) );
NOR2_X1 U1078 ( .A1(G122), .A2(KEYINPUT58), .ZN(n1365) );
XNOR2_X1 U1079 ( .A(n1366), .B(n1367), .ZN(n1178) );
XNOR2_X1 U1080 ( .A(n1296), .B(G116), .ZN(n1367) );
INV_X1 U1081 ( .A(G119), .ZN(n1296) );
NAND2_X1 U1082 ( .A1(KEYINPUT30), .A2(n1324), .ZN(n1366) );
XOR2_X1 U1083 ( .A(n1211), .B(n1368), .Z(n1360) );
XOR2_X1 U1084 ( .A(G125), .B(n1369), .Z(n1368) );
AND2_X1 U1085 ( .A1(n1148), .A2(G224), .ZN(n1369) );
XNOR2_X1 U1086 ( .A(n1154), .B(KEYINPUT61), .ZN(n1211) );
INV_X1 U1087 ( .A(n1352), .ZN(n1154) );
XNOR2_X1 U1088 ( .A(n1370), .B(n1371), .ZN(n1352) );
XOR2_X1 U1089 ( .A(G143), .B(G128), .Z(n1371) );
XNOR2_X1 U1090 ( .A(G146), .B(KEYINPUT22), .ZN(n1370) );
NOR2_X1 U1091 ( .A1(n1129), .A2(n1277), .ZN(n1082) );
XNOR2_X1 U1092 ( .A(n1134), .B(G475), .ZN(n1277) );
NAND2_X1 U1093 ( .A1(n1201), .A2(n1198), .ZN(n1134) );
INV_X1 U1094 ( .A(G902), .ZN(n1198) );
XOR2_X1 U1095 ( .A(n1372), .B(n1373), .Z(n1201) );
XNOR2_X1 U1096 ( .A(n1374), .B(n1375), .ZN(n1373) );
NOR2_X1 U1097 ( .A1(KEYINPUT21), .A2(n1324), .ZN(n1375) );
XNOR2_X1 U1098 ( .A(G113), .B(KEYINPUT1), .ZN(n1324) );
NAND2_X1 U1099 ( .A1(KEYINPUT44), .A2(n1376), .ZN(n1374) );
XOR2_X1 U1100 ( .A(n1330), .B(n1377), .Z(n1376) );
XNOR2_X1 U1101 ( .A(n1378), .B(n1379), .ZN(n1377) );
INV_X1 U1102 ( .A(G125), .ZN(n1379) );
NAND3_X1 U1103 ( .A1(n1380), .A2(n1381), .A3(n1382), .ZN(n1378) );
OR2_X1 U1104 ( .A1(n1383), .A2(G131), .ZN(n1382) );
NAND2_X1 U1105 ( .A1(KEYINPUT32), .A2(n1384), .ZN(n1381) );
NAND2_X1 U1106 ( .A1(n1385), .A2(n1383), .ZN(n1384) );
XNOR2_X1 U1107 ( .A(KEYINPUT5), .B(G131), .ZN(n1385) );
NAND2_X1 U1108 ( .A1(n1386), .A2(n1387), .ZN(n1380) );
INV_X1 U1109 ( .A(KEYINPUT32), .ZN(n1387) );
NAND2_X1 U1110 ( .A1(n1388), .A2(n1389), .ZN(n1386) );
OR2_X1 U1111 ( .A1(G131), .A2(KEYINPUT5), .ZN(n1389) );
NAND3_X1 U1112 ( .A1(G131), .A2(n1383), .A3(KEYINPUT5), .ZN(n1388) );
XNOR2_X1 U1113 ( .A(G143), .B(n1390), .ZN(n1383) );
NOR4_X1 U1114 ( .A1(KEYINPUT13), .A2(G953), .A3(G237), .A4(n1391), .ZN(n1390) );
INV_X1 U1115 ( .A(G214), .ZN(n1391) );
XNOR2_X1 U1116 ( .A(G146), .B(G140), .ZN(n1330) );
XNOR2_X1 U1117 ( .A(G104), .B(G122), .ZN(n1372) );
XNOR2_X1 U1118 ( .A(n1392), .B(G478), .ZN(n1129) );
NAND2_X1 U1119 ( .A1(n1393), .A2(n1195), .ZN(n1392) );
XOR2_X1 U1120 ( .A(n1394), .B(n1395), .Z(n1195) );
XOR2_X1 U1121 ( .A(n1396), .B(n1397), .Z(n1395) );
XNOR2_X1 U1122 ( .A(G107), .B(n1398), .ZN(n1397) );
NOR2_X1 U1123 ( .A1(G143), .A2(KEYINPUT41), .ZN(n1398) );
NAND2_X1 U1124 ( .A1(G217), .A2(n1337), .ZN(n1396) );
AND2_X1 U1125 ( .A1(G234), .A2(n1148), .ZN(n1337) );
INV_X1 U1126 ( .A(G953), .ZN(n1148) );
XOR2_X1 U1127 ( .A(n1399), .B(n1400), .Z(n1394) );
XNOR2_X1 U1128 ( .A(G122), .B(n1301), .ZN(n1400) );
INV_X1 U1129 ( .A(G116), .ZN(n1301) );
XNOR2_X1 U1130 ( .A(G134), .B(G128), .ZN(n1399) );
XNOR2_X1 U1131 ( .A(G902), .B(KEYINPUT11), .ZN(n1393) );
NAND2_X1 U1132 ( .A1(KEYINPUT33), .A2(n1342), .ZN(n1311) );
INV_X1 U1133 ( .A(G110), .ZN(n1342) );
endmodule


