//Key = 0011010010011101100000101001101011100110011100000111001110111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351;

XNOR2_X1 U731 ( .A(G107), .B(n1022), .ZN(G9) );
NOR2_X1 U732 ( .A1(n1023), .A2(n1024), .ZN(G75) );
NOR4_X1 U733 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
NOR2_X1 U734 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U735 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U736 ( .A1(KEYINPUT11), .A2(n1033), .ZN(n1032) );
NOR4_X1 U737 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1033) );
NOR2_X1 U738 ( .A1(n1038), .A2(n1037), .ZN(n1031) );
NOR2_X1 U739 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U740 ( .A1(n1041), .A2(n1036), .ZN(n1040) );
NOR2_X1 U741 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR2_X1 U742 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U743 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U744 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
AND3_X1 U745 ( .A1(KEYINPUT11), .A2(n1050), .A3(n1051), .ZN(n1042) );
NOR3_X1 U746 ( .A1(n1035), .A2(n1045), .A3(n1052), .ZN(n1039) );
INV_X1 U747 ( .A(n1053), .ZN(n1045) );
INV_X1 U748 ( .A(n1051), .ZN(n1035) );
NAND3_X1 U749 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1025) );
NAND3_X1 U750 ( .A1(n1051), .A2(n1057), .A3(n1058), .ZN(n1056) );
INV_X1 U751 ( .A(n1037), .ZN(n1058) );
NAND2_X1 U752 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND3_X1 U753 ( .A1(n1061), .A2(n1053), .A3(n1062), .ZN(n1060) );
NAND2_X1 U754 ( .A1(n1063), .A2(n1064), .ZN(n1059) );
NAND2_X1 U755 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U756 ( .A1(n1053), .A2(n1067), .ZN(n1066) );
NAND3_X1 U757 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
OR3_X1 U758 ( .A1(n1071), .A2(n1072), .A3(KEYINPUT45), .ZN(n1069) );
NAND2_X1 U759 ( .A1(KEYINPUT45), .A2(n1062), .ZN(n1068) );
NAND2_X1 U760 ( .A1(n1073), .A2(n1062), .ZN(n1065) );
NOR3_X1 U761 ( .A1(n1074), .A2(G953), .A3(G952), .ZN(n1023) );
INV_X1 U762 ( .A(n1054), .ZN(n1074) );
NAND4_X1 U763 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1054) );
NOR4_X1 U764 ( .A1(n1079), .A2(n1080), .A3(n1030), .A4(n1081), .ZN(n1078) );
XNOR2_X1 U765 ( .A(G469), .B(n1082), .ZN(n1081) );
XNOR2_X1 U766 ( .A(n1083), .B(KEYINPUT60), .ZN(n1080) );
XOR2_X1 U767 ( .A(n1084), .B(n1085), .Z(n1079) );
NAND2_X1 U768 ( .A1(KEYINPUT22), .A2(n1086), .ZN(n1084) );
NOR3_X1 U769 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1077) );
OR2_X1 U770 ( .A1(n1090), .A2(n1091), .ZN(n1075) );
XOR2_X1 U771 ( .A(n1092), .B(n1093), .Z(G72) );
NOR2_X1 U772 ( .A1(n1094), .A2(n1055), .ZN(n1093) );
NOR2_X1 U773 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XNOR2_X1 U774 ( .A(G900), .B(KEYINPUT10), .ZN(n1095) );
NAND2_X1 U775 ( .A1(n1097), .A2(n1098), .ZN(n1092) );
NAND2_X1 U776 ( .A1(n1099), .A2(n1055), .ZN(n1098) );
XNOR2_X1 U777 ( .A(n1100), .B(n1101), .ZN(n1099) );
NAND3_X1 U778 ( .A1(G900), .A2(n1101), .A3(G953), .ZN(n1097) );
XNOR2_X1 U779 ( .A(n1102), .B(n1103), .ZN(n1101) );
XNOR2_X1 U780 ( .A(n1104), .B(KEYINPUT59), .ZN(n1102) );
NAND3_X1 U781 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(G69) );
XOR2_X1 U782 ( .A(n1108), .B(KEYINPUT14), .Z(n1107) );
NAND3_X1 U783 ( .A1(n1109), .A2(n1110), .A3(G953), .ZN(n1108) );
NAND2_X1 U784 ( .A1(G898), .A2(G224), .ZN(n1109) );
NAND2_X1 U785 ( .A1(n1111), .A2(n1055), .ZN(n1106) );
XNOR2_X1 U786 ( .A(n1110), .B(n1028), .ZN(n1111) );
NAND4_X1 U787 ( .A1(G898), .A2(G224), .A3(n1112), .A4(G953), .ZN(n1105) );
INV_X1 U788 ( .A(n1110), .ZN(n1112) );
NAND2_X1 U789 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
XOR2_X1 U790 ( .A(n1115), .B(KEYINPUT31), .Z(n1113) );
NAND2_X1 U791 ( .A1(G953), .A2(n1116), .ZN(n1115) );
NOR2_X1 U792 ( .A1(n1117), .A2(n1118), .ZN(G66) );
XOR2_X1 U793 ( .A(n1119), .B(n1120), .Z(n1118) );
NOR2_X1 U794 ( .A1(n1090), .A2(n1121), .ZN(n1120) );
NOR2_X1 U795 ( .A1(n1117), .A2(n1122), .ZN(G63) );
NOR2_X1 U796 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U797 ( .A(KEYINPUT29), .B(n1125), .Z(n1124) );
NOR3_X1 U798 ( .A1(n1121), .A2(n1126), .A3(n1127), .ZN(n1125) );
XNOR2_X1 U799 ( .A(n1128), .B(KEYINPUT61), .ZN(n1126) );
NOR2_X1 U800 ( .A1(n1129), .A2(n1128), .ZN(n1123) );
XOR2_X1 U801 ( .A(n1130), .B(KEYINPUT15), .Z(n1128) );
NOR2_X1 U802 ( .A1(n1127), .A2(n1121), .ZN(n1129) );
INV_X1 U803 ( .A(G478), .ZN(n1127) );
NOR2_X1 U804 ( .A1(n1117), .A2(n1131), .ZN(G60) );
NOR3_X1 U805 ( .A1(n1085), .A2(n1132), .A3(n1133), .ZN(n1131) );
NOR3_X1 U806 ( .A1(n1134), .A2(n1086), .A3(n1121), .ZN(n1133) );
INV_X1 U807 ( .A(n1135), .ZN(n1134) );
NOR2_X1 U808 ( .A1(n1136), .A2(n1135), .ZN(n1132) );
AND2_X1 U809 ( .A1(n1137), .A2(G475), .ZN(n1136) );
XNOR2_X1 U810 ( .A(n1138), .B(n1139), .ZN(G6) );
NOR2_X1 U811 ( .A1(KEYINPUT53), .A2(n1140), .ZN(n1139) );
NOR2_X1 U812 ( .A1(n1117), .A2(n1141), .ZN(G57) );
XOR2_X1 U813 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U814 ( .A(n1144), .B(n1145), .Z(n1143) );
NOR2_X1 U815 ( .A1(n1146), .A2(n1121), .ZN(n1144) );
XOR2_X1 U816 ( .A(n1147), .B(n1148), .Z(n1142) );
XNOR2_X1 U817 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR2_X1 U818 ( .A1(KEYINPUT6), .A2(n1151), .ZN(n1150) );
NOR2_X1 U819 ( .A1(n1152), .A2(n1153), .ZN(n1147) );
XOR2_X1 U820 ( .A(n1154), .B(KEYINPUT41), .Z(n1153) );
NAND2_X1 U821 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U822 ( .A1(n1155), .A2(n1156), .ZN(n1152) );
NOR2_X1 U823 ( .A1(n1117), .A2(n1157), .ZN(G54) );
XOR2_X1 U824 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U825 ( .A1(n1160), .A2(n1121), .ZN(n1159) );
NOR3_X1 U826 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1158) );
NOR2_X1 U827 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NOR2_X1 U828 ( .A1(KEYINPUT4), .A2(n1166), .ZN(n1164) );
XNOR2_X1 U829 ( .A(n1167), .B(KEYINPUT30), .ZN(n1166) );
NOR3_X1 U830 ( .A1(n1168), .A2(KEYINPUT4), .A3(n1167), .ZN(n1162) );
INV_X1 U831 ( .A(n1165), .ZN(n1168) );
XNOR2_X1 U832 ( .A(n1169), .B(n1170), .ZN(n1165) );
XNOR2_X1 U833 ( .A(n1171), .B(n1172), .ZN(n1169) );
NOR2_X1 U834 ( .A1(KEYINPUT46), .A2(n1173), .ZN(n1172) );
XOR2_X1 U835 ( .A(KEYINPUT27), .B(n1155), .Z(n1173) );
AND2_X1 U836 ( .A1(n1167), .A2(KEYINPUT4), .ZN(n1161) );
XOR2_X1 U837 ( .A(n1174), .B(n1175), .Z(n1167) );
NOR2_X1 U838 ( .A1(KEYINPUT26), .A2(n1176), .ZN(n1175) );
XOR2_X1 U839 ( .A(n1177), .B(KEYINPUT9), .Z(n1176) );
NOR2_X1 U840 ( .A1(n1117), .A2(n1178), .ZN(G51) );
XOR2_X1 U841 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U842 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U843 ( .A(KEYINPUT18), .B(n1183), .Z(n1182) );
NOR2_X1 U844 ( .A1(KEYINPUT7), .A2(n1184), .ZN(n1183) );
NOR2_X1 U845 ( .A1(n1185), .A2(n1121), .ZN(n1181) );
NAND2_X1 U846 ( .A1(G902), .A2(n1137), .ZN(n1121) );
NAND2_X1 U847 ( .A1(n1100), .A2(n1186), .ZN(n1137) );
XNOR2_X1 U848 ( .A(KEYINPUT23), .B(n1028), .ZN(n1186) );
NAND4_X1 U849 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1028) );
AND4_X1 U850 ( .A1(n1022), .A2(n1191), .A3(n1192), .A4(n1138), .ZN(n1190) );
NAND3_X1 U851 ( .A1(n1053), .A2(n1193), .A3(n1194), .ZN(n1138) );
NAND3_X1 U852 ( .A1(n1053), .A2(n1193), .A3(n1061), .ZN(n1022) );
NAND2_X1 U853 ( .A1(n1195), .A2(n1196), .ZN(n1188) );
OR2_X1 U854 ( .A1(n1073), .A2(n1050), .ZN(n1196) );
OR2_X1 U855 ( .A1(n1197), .A2(n1070), .ZN(n1187) );
INV_X1 U856 ( .A(n1026), .ZN(n1100) );
NAND4_X1 U857 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1026) );
NOR4_X1 U858 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
INV_X1 U859 ( .A(n1206), .ZN(n1202) );
NOR2_X1 U860 ( .A1(n1207), .A2(n1208), .ZN(n1200) );
NOR2_X1 U861 ( .A1(n1070), .A2(n1209), .ZN(n1208) );
XNOR2_X1 U862 ( .A(KEYINPUT3), .B(n1210), .ZN(n1209) );
NOR2_X1 U863 ( .A1(n1211), .A2(n1212), .ZN(n1207) );
XNOR2_X1 U864 ( .A(KEYINPUT52), .B(n1213), .ZN(n1212) );
NAND3_X1 U865 ( .A1(n1214), .A2(n1062), .A3(n1063), .ZN(n1198) );
XOR2_X1 U866 ( .A(n1215), .B(n1216), .Z(n1179) );
NOR2_X1 U867 ( .A1(KEYINPUT57), .A2(n1156), .ZN(n1216) );
NOR2_X1 U868 ( .A1(n1055), .A2(G952), .ZN(n1117) );
XNOR2_X1 U869 ( .A(G146), .B(n1217), .ZN(G48) );
NAND2_X1 U870 ( .A1(KEYINPUT2), .A2(n1203), .ZN(n1217) );
NOR3_X1 U871 ( .A1(n1052), .A2(n1070), .A3(n1218), .ZN(n1203) );
XOR2_X1 U872 ( .A(n1199), .B(n1219), .Z(G45) );
XNOR2_X1 U873 ( .A(KEYINPUT63), .B(n1220), .ZN(n1219) );
NAND4_X1 U874 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1199) );
XOR2_X1 U875 ( .A(G140), .B(n1225), .Z(G42) );
NOR2_X1 U876 ( .A1(n1211), .A2(n1226), .ZN(n1225) );
XNOR2_X1 U877 ( .A(KEYINPUT39), .B(n1213), .ZN(n1226) );
NAND4_X1 U878 ( .A1(n1073), .A2(n1194), .A3(n1062), .A4(n1047), .ZN(n1211) );
XOR2_X1 U879 ( .A(G137), .B(n1227), .Z(G39) );
NOR3_X1 U880 ( .A1(n1228), .A2(n1030), .A3(n1218), .ZN(n1227) );
XNOR2_X1 U881 ( .A(KEYINPUT8), .B(n1036), .ZN(n1228) );
INV_X1 U882 ( .A(n1063), .ZN(n1036) );
XOR2_X1 U883 ( .A(G134), .B(n1205), .Z(G36) );
AND3_X1 U884 ( .A1(n1062), .A2(n1061), .A3(n1221), .ZN(n1205) );
XNOR2_X1 U885 ( .A(G131), .B(n1206), .ZN(G33) );
NAND3_X1 U886 ( .A1(n1221), .A2(n1062), .A3(n1194), .ZN(n1206) );
INV_X1 U887 ( .A(n1030), .ZN(n1062) );
NAND2_X1 U888 ( .A1(n1229), .A2(n1071), .ZN(n1030) );
AND3_X1 U889 ( .A1(n1047), .A2(n1213), .A3(n1050), .ZN(n1221) );
XOR2_X1 U890 ( .A(G128), .B(n1230), .Z(G30) );
NOR3_X1 U891 ( .A1(n1210), .A2(KEYINPUT20), .A3(n1070), .ZN(n1230) );
NAND2_X1 U892 ( .A1(n1214), .A2(n1061), .ZN(n1210) );
INV_X1 U893 ( .A(n1218), .ZN(n1214) );
NAND4_X1 U894 ( .A1(n1047), .A2(n1083), .A3(n1213), .A4(n1231), .ZN(n1218) );
XNOR2_X1 U895 ( .A(G101), .B(n1232), .ZN(G3) );
NAND2_X1 U896 ( .A1(n1195), .A2(n1050), .ZN(n1232) );
XOR2_X1 U897 ( .A(G125), .B(n1204), .Z(G27) );
AND4_X1 U898 ( .A1(n1073), .A2(n1051), .A3(n1233), .A4(n1194), .ZN(n1204) );
NOR2_X1 U899 ( .A1(n1234), .A2(n1070), .ZN(n1233) );
INV_X1 U900 ( .A(n1213), .ZN(n1234) );
NAND2_X1 U901 ( .A1(n1037), .A2(n1235), .ZN(n1213) );
NAND4_X1 U902 ( .A1(G953), .A2(G902), .A3(n1236), .A4(n1237), .ZN(n1235) );
INV_X1 U903 ( .A(G900), .ZN(n1237) );
XOR2_X1 U904 ( .A(n1238), .B(n1239), .Z(G24) );
XNOR2_X1 U905 ( .A(KEYINPUT51), .B(n1240), .ZN(n1239) );
NAND2_X1 U906 ( .A1(KEYINPUT38), .A2(n1241), .ZN(n1238) );
INV_X1 U907 ( .A(n1189), .ZN(n1241) );
NAND4_X1 U908 ( .A1(n1242), .A2(n1053), .A3(n1223), .A4(n1224), .ZN(n1189) );
NOR2_X1 U909 ( .A1(n1231), .A2(n1083), .ZN(n1053) );
XNOR2_X1 U910 ( .A(G119), .B(n1192), .ZN(G21) );
NAND4_X1 U911 ( .A1(n1242), .A2(n1063), .A3(n1083), .A4(n1231), .ZN(n1192) );
XNOR2_X1 U912 ( .A(G116), .B(n1243), .ZN(G18) );
NAND2_X1 U913 ( .A1(n1244), .A2(n1222), .ZN(n1243) );
XOR2_X1 U914 ( .A(n1197), .B(KEYINPUT54), .Z(n1244) );
NAND4_X1 U915 ( .A1(n1051), .A2(n1050), .A3(n1061), .A4(n1245), .ZN(n1197) );
NOR2_X1 U916 ( .A1(n1223), .A2(n1246), .ZN(n1061) );
XOR2_X1 U917 ( .A(G113), .B(n1247), .Z(G15) );
NOR2_X1 U918 ( .A1(KEYINPUT40), .A2(n1191), .ZN(n1247) );
NAND3_X1 U919 ( .A1(n1194), .A2(n1050), .A3(n1242), .ZN(n1191) );
AND3_X1 U920 ( .A1(n1222), .A2(n1245), .A3(n1051), .ZN(n1242) );
NOR2_X1 U921 ( .A1(n1048), .A2(n1088), .ZN(n1051) );
INV_X1 U922 ( .A(n1049), .ZN(n1088) );
INV_X1 U923 ( .A(n1034), .ZN(n1050) );
NAND2_X1 U924 ( .A1(n1248), .A2(n1083), .ZN(n1034) );
INV_X1 U925 ( .A(n1052), .ZN(n1194) );
NAND2_X1 U926 ( .A1(n1246), .A2(n1223), .ZN(n1052) );
NAND2_X1 U927 ( .A1(n1249), .A2(n1250), .ZN(G12) );
NAND2_X1 U928 ( .A1(G110), .A2(n1251), .ZN(n1250) );
XOR2_X1 U929 ( .A(KEYINPUT28), .B(n1252), .Z(n1249) );
NOR2_X1 U930 ( .A1(G110), .A2(n1251), .ZN(n1252) );
NAND2_X1 U931 ( .A1(n1195), .A2(n1253), .ZN(n1251) );
XOR2_X1 U932 ( .A(KEYINPUT21), .B(n1073), .Z(n1253) );
NOR2_X1 U933 ( .A1(n1083), .A2(n1248), .ZN(n1073) );
INV_X1 U934 ( .A(n1231), .ZN(n1248) );
NAND3_X1 U935 ( .A1(n1254), .A2(n1255), .A3(n1076), .ZN(n1231) );
NAND2_X1 U936 ( .A1(n1091), .A2(n1090), .ZN(n1076) );
NAND2_X1 U937 ( .A1(KEYINPUT1), .A2(n1090), .ZN(n1255) );
OR3_X1 U938 ( .A1(n1091), .A2(KEYINPUT1), .A3(n1090), .ZN(n1254) );
NAND2_X1 U939 ( .A1(G217), .A2(n1256), .ZN(n1090) );
NOR2_X1 U940 ( .A1(n1119), .A2(G902), .ZN(n1091) );
XOR2_X1 U941 ( .A(n1257), .B(n1258), .Z(n1119) );
XOR2_X1 U942 ( .A(G110), .B(n1259), .Z(n1258) );
XOR2_X1 U943 ( .A(KEYINPUT37), .B(G137), .Z(n1259) );
XOR2_X1 U944 ( .A(n1260), .B(n1261), .Z(n1257) );
XOR2_X1 U945 ( .A(n1262), .B(n1263), .Z(n1260) );
AND2_X1 U946 ( .A1(n1264), .A2(G221), .ZN(n1263) );
NAND2_X1 U947 ( .A1(n1265), .A2(n1266), .ZN(n1262) );
NAND2_X1 U948 ( .A1(G128), .A2(n1267), .ZN(n1266) );
XOR2_X1 U949 ( .A(KEYINPUT5), .B(n1268), .Z(n1265) );
NOR2_X1 U950 ( .A1(G128), .A2(n1267), .ZN(n1268) );
XOR2_X1 U951 ( .A(n1269), .B(n1146), .Z(n1083) );
INV_X1 U952 ( .A(G472), .ZN(n1146) );
NAND2_X1 U953 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XOR2_X1 U954 ( .A(n1272), .B(n1273), .Z(n1270) );
XNOR2_X1 U955 ( .A(n1274), .B(n1156), .ZN(n1273) );
XOR2_X1 U956 ( .A(n1275), .B(n1155), .Z(n1274) );
NAND2_X1 U957 ( .A1(KEYINPUT13), .A2(n1276), .ZN(n1275) );
XOR2_X1 U958 ( .A(KEYINPUT62), .B(n1145), .Z(n1276) );
XNOR2_X1 U959 ( .A(n1277), .B(G113), .ZN(n1145) );
NAND2_X1 U960 ( .A1(KEYINPUT42), .A2(n1278), .ZN(n1277) );
XOR2_X1 U961 ( .A(n1279), .B(n1280), .Z(n1272) );
NOR2_X1 U962 ( .A1(G101), .A2(KEYINPUT47), .ZN(n1280) );
XOR2_X1 U963 ( .A(n1149), .B(KEYINPUT0), .Z(n1279) );
NAND3_X1 U964 ( .A1(n1281), .A2(n1055), .A3(G210), .ZN(n1149) );
AND2_X1 U965 ( .A1(n1063), .A2(n1193), .ZN(n1195) );
AND3_X1 U966 ( .A1(n1222), .A2(n1245), .A3(n1047), .ZN(n1193) );
AND2_X1 U967 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U968 ( .A1(G221), .A2(n1256), .ZN(n1049) );
NAND2_X1 U969 ( .A1(G234), .A2(n1271), .ZN(n1256) );
NAND3_X1 U970 ( .A1(n1282), .A2(n1283), .A3(n1284), .ZN(n1048) );
OR2_X1 U971 ( .A1(n1082), .A2(KEYINPUT49), .ZN(n1284) );
NAND3_X1 U972 ( .A1(KEYINPUT49), .A2(n1082), .A3(G469), .ZN(n1283) );
NAND2_X1 U973 ( .A1(n1285), .A2(n1160), .ZN(n1282) );
INV_X1 U974 ( .A(G469), .ZN(n1160) );
NAND2_X1 U975 ( .A1(n1286), .A2(KEYINPUT49), .ZN(n1285) );
XOR2_X1 U976 ( .A(n1082), .B(KEYINPUT17), .Z(n1286) );
NAND2_X1 U977 ( .A1(n1287), .A2(n1271), .ZN(n1082) );
XOR2_X1 U978 ( .A(n1288), .B(n1289), .Z(n1287) );
XNOR2_X1 U979 ( .A(n1290), .B(n1291), .ZN(n1289) );
XOR2_X1 U980 ( .A(n1292), .B(n1177), .Z(n1291) );
XNOR2_X1 U981 ( .A(G140), .B(G110), .ZN(n1177) );
NAND2_X1 U982 ( .A1(KEYINPUT34), .A2(n1170), .ZN(n1292) );
INV_X1 U983 ( .A(n1104), .ZN(n1290) );
XOR2_X1 U984 ( .A(n1171), .B(n1155), .Z(n1104) );
XOR2_X1 U985 ( .A(n1293), .B(n1294), .Z(n1155) );
XNOR2_X1 U986 ( .A(G131), .B(G137), .ZN(n1293) );
XNOR2_X1 U987 ( .A(n1295), .B(n1296), .ZN(n1288) );
XOR2_X1 U988 ( .A(KEYINPUT43), .B(KEYINPUT27), .Z(n1296) );
INV_X1 U989 ( .A(n1174), .ZN(n1295) );
NOR2_X1 U990 ( .A1(n1096), .A2(G953), .ZN(n1174) );
INV_X1 U991 ( .A(G227), .ZN(n1096) );
NAND2_X1 U992 ( .A1(n1037), .A2(n1297), .ZN(n1245) );
NAND4_X1 U993 ( .A1(G953), .A2(G902), .A3(n1236), .A4(n1116), .ZN(n1297) );
INV_X1 U994 ( .A(G898), .ZN(n1116) );
NAND3_X1 U995 ( .A1(n1236), .A2(n1055), .A3(G952), .ZN(n1037) );
NAND2_X1 U996 ( .A1(G237), .A2(G234), .ZN(n1236) );
INV_X1 U997 ( .A(n1070), .ZN(n1222) );
NAND2_X1 U998 ( .A1(n1072), .A2(n1071), .ZN(n1070) );
NAND2_X1 U999 ( .A1(G214), .A2(n1298), .ZN(n1071) );
INV_X1 U1000 ( .A(n1229), .ZN(n1072) );
XNOR2_X1 U1001 ( .A(n1299), .B(n1185), .ZN(n1229) );
NAND2_X1 U1002 ( .A1(G210), .A2(n1298), .ZN(n1185) );
NAND2_X1 U1003 ( .A1(n1300), .A2(n1271), .ZN(n1298) );
INV_X1 U1004 ( .A(G237), .ZN(n1300) );
NAND2_X1 U1005 ( .A1(n1301), .A2(n1271), .ZN(n1299) );
XOR2_X1 U1006 ( .A(n1156), .B(n1302), .Z(n1301) );
XNOR2_X1 U1007 ( .A(n1215), .B(n1184), .ZN(n1302) );
NAND2_X1 U1008 ( .A1(G224), .A2(n1055), .ZN(n1184) );
XNOR2_X1 U1009 ( .A(n1114), .B(G125), .ZN(n1215) );
XNOR2_X1 U1010 ( .A(n1303), .B(n1304), .ZN(n1114) );
XOR2_X1 U1011 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1012 ( .A(G110), .B(G122), .ZN(n1306) );
NAND2_X1 U1013 ( .A1(KEYINPUT55), .A2(G113), .ZN(n1305) );
XNOR2_X1 U1014 ( .A(n1278), .B(n1170), .ZN(n1303) );
XNOR2_X1 U1015 ( .A(n1151), .B(n1307), .ZN(n1170) );
XNOR2_X1 U1016 ( .A(G107), .B(n1140), .ZN(n1307) );
INV_X1 U1017 ( .A(G104), .ZN(n1140) );
INV_X1 U1018 ( .A(G101), .ZN(n1151) );
XOR2_X1 U1019 ( .A(G116), .B(n1308), .Z(n1278) );
XNOR2_X1 U1020 ( .A(KEYINPUT12), .B(n1267), .ZN(n1308) );
INV_X1 U1021 ( .A(G119), .ZN(n1267) );
NAND2_X1 U1022 ( .A1(n1309), .A2(n1310), .ZN(n1156) );
NAND3_X1 U1023 ( .A1(G128), .A2(n1311), .A3(n1312), .ZN(n1310) );
INV_X1 U1024 ( .A(KEYINPUT50), .ZN(n1312) );
NAND2_X1 U1025 ( .A1(n1171), .A2(KEYINPUT50), .ZN(n1309) );
XOR2_X1 U1026 ( .A(G128), .B(n1311), .Z(n1171) );
XNOR2_X1 U1027 ( .A(G146), .B(n1220), .ZN(n1311) );
NOR2_X1 U1028 ( .A1(n1224), .A2(n1223), .ZN(n1063) );
XNOR2_X1 U1029 ( .A(n1085), .B(n1086), .ZN(n1223) );
INV_X1 U1030 ( .A(G475), .ZN(n1086) );
NOR2_X1 U1031 ( .A1(n1135), .A2(G902), .ZN(n1085) );
XNOR2_X1 U1032 ( .A(n1313), .B(n1314), .ZN(n1135) );
XOR2_X1 U1033 ( .A(n1261), .B(n1315), .Z(n1314) );
XOR2_X1 U1034 ( .A(n1316), .B(n1317), .Z(n1315) );
NAND2_X1 U1035 ( .A1(n1318), .A2(KEYINPUT56), .ZN(n1317) );
XNOR2_X1 U1036 ( .A(G104), .B(n1319), .ZN(n1318) );
XNOR2_X1 U1037 ( .A(n1240), .B(G113), .ZN(n1319) );
NAND3_X1 U1038 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1316) );
OR2_X1 U1039 ( .A1(n1323), .A2(n1220), .ZN(n1322) );
NAND2_X1 U1040 ( .A1(KEYINPUT35), .A2(n1324), .ZN(n1321) );
NAND2_X1 U1041 ( .A1(n1325), .A2(n1220), .ZN(n1324) );
XNOR2_X1 U1042 ( .A(KEYINPUT58), .B(n1323), .ZN(n1325) );
NAND2_X1 U1043 ( .A1(n1326), .A2(n1327), .ZN(n1320) );
INV_X1 U1044 ( .A(KEYINPUT35), .ZN(n1327) );
NAND2_X1 U1045 ( .A1(n1328), .A2(n1329), .ZN(n1326) );
OR2_X1 U1046 ( .A1(n1323), .A2(KEYINPUT58), .ZN(n1329) );
NAND3_X1 U1047 ( .A1(n1323), .A2(n1220), .A3(KEYINPUT58), .ZN(n1328) );
INV_X1 U1048 ( .A(G143), .ZN(n1220) );
NAND3_X1 U1049 ( .A1(n1281), .A2(n1055), .A3(G214), .ZN(n1323) );
XNOR2_X1 U1050 ( .A(G237), .B(KEYINPUT25), .ZN(n1281) );
XOR2_X1 U1051 ( .A(G146), .B(n1103), .Z(n1261) );
XOR2_X1 U1052 ( .A(G125), .B(G140), .Z(n1103) );
XNOR2_X1 U1053 ( .A(n1330), .B(n1331), .ZN(n1313) );
INV_X1 U1054 ( .A(G131), .ZN(n1331) );
XNOR2_X1 U1055 ( .A(KEYINPUT33), .B(KEYINPUT24), .ZN(n1330) );
INV_X1 U1056 ( .A(n1246), .ZN(n1224) );
NOR2_X1 U1057 ( .A1(n1332), .A2(n1087), .ZN(n1246) );
NOR3_X1 U1058 ( .A1(G478), .A2(G902), .A3(n1333), .ZN(n1087) );
INV_X1 U1059 ( .A(n1130), .ZN(n1333) );
XNOR2_X1 U1060 ( .A(KEYINPUT32), .B(n1089), .ZN(n1332) );
AND2_X1 U1061 ( .A1(G478), .A2(n1334), .ZN(n1089) );
NAND2_X1 U1062 ( .A1(n1130), .A2(n1271), .ZN(n1334) );
INV_X1 U1063 ( .A(G902), .ZN(n1271) );
XNOR2_X1 U1064 ( .A(n1335), .B(n1336), .ZN(n1130) );
XOR2_X1 U1065 ( .A(n1337), .B(n1338), .Z(n1336) );
NAND3_X1 U1066 ( .A1(n1339), .A2(n1340), .A3(n1341), .ZN(n1338) );
OR2_X1 U1067 ( .A1(n1342), .A2(KEYINPUT16), .ZN(n1341) );
NAND3_X1 U1068 ( .A1(KEYINPUT16), .A2(n1342), .A3(G122), .ZN(n1340) );
INV_X1 U1069 ( .A(G116), .ZN(n1342) );
NAND2_X1 U1070 ( .A1(n1343), .A2(n1240), .ZN(n1339) );
INV_X1 U1071 ( .A(G122), .ZN(n1240) );
NAND2_X1 U1072 ( .A1(n1344), .A2(KEYINPUT16), .ZN(n1343) );
XNOR2_X1 U1073 ( .A(G116), .B(KEYINPUT36), .ZN(n1344) );
NAND3_X1 U1074 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1337) );
NAND2_X1 U1075 ( .A1(KEYINPUT19), .A2(n1348), .ZN(n1347) );
NAND3_X1 U1076 ( .A1(n1349), .A2(n1350), .A3(n1294), .ZN(n1346) );
INV_X1 U1077 ( .A(KEYINPUT19), .ZN(n1350) );
OR2_X1 U1078 ( .A1(n1294), .A2(n1349), .ZN(n1345) );
NOR2_X1 U1079 ( .A1(KEYINPUT44), .A2(n1348), .ZN(n1349) );
XNOR2_X1 U1080 ( .A(G128), .B(G143), .ZN(n1348) );
XNOR2_X1 U1081 ( .A(G134), .B(KEYINPUT48), .ZN(n1294) );
XOR2_X1 U1082 ( .A(n1351), .B(G107), .Z(n1335) );
NAND2_X1 U1083 ( .A1(G217), .A2(n1264), .ZN(n1351) );
AND2_X1 U1084 ( .A1(G234), .A2(n1055), .ZN(n1264) );
INV_X1 U1085 ( .A(G953), .ZN(n1055) );
endmodule


