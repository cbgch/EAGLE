//Key = 1010110111100011000011000001000001111010110011111111111010010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325;

XOR2_X1 U737 ( .A(G107), .B(n1010), .Z(G9) );
NOR2_X1 U738 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NOR2_X1 U739 ( .A1(n1013), .A2(n1014), .ZN(G75) );
NOR4_X1 U740 ( .A1(G953), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1014) );
NOR2_X1 U741 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NOR2_X1 U742 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR2_X1 U743 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
INV_X1 U744 ( .A(n1024), .ZN(n1023) );
NOR2_X1 U745 ( .A1(n1025), .A2(n1026), .ZN(n1022) );
NOR2_X1 U746 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NOR2_X1 U747 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U748 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U749 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U750 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U751 ( .A1(n1037), .A2(n1038), .ZN(n1029) );
NOR2_X1 U752 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR3_X1 U753 ( .A1(n1038), .A2(n1041), .A3(n1032), .ZN(n1025) );
NOR2_X1 U754 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR2_X1 U755 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR4_X1 U756 ( .A1(n1046), .A2(n1032), .A3(n1038), .A4(n1028), .ZN(n1020) );
INV_X1 U757 ( .A(n1047), .ZN(n1032) );
NOR2_X1 U758 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR3_X1 U759 ( .A1(n1015), .A2(G953), .A3(G952), .ZN(n1013) );
AND4_X1 U760 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1015) );
NOR3_X1 U761 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NAND3_X1 U762 ( .A1(n1057), .A2(n1058), .A3(n1036), .ZN(n1054) );
NOR3_X1 U763 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1052) );
XNOR2_X1 U764 ( .A(n1062), .B(KEYINPUT11), .ZN(n1061) );
NOR2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(n1060) );
XNOR2_X1 U766 ( .A(KEYINPUT53), .B(n1065), .ZN(n1064) );
XNOR2_X1 U767 ( .A(n1066), .B(n1067), .ZN(n1051) );
XOR2_X1 U768 ( .A(n1068), .B(KEYINPUT55), .Z(n1066) );
XNOR2_X1 U769 ( .A(n1069), .B(KEYINPUT19), .ZN(n1050) );
XOR2_X1 U770 ( .A(n1070), .B(n1071), .Z(G72) );
XOR2_X1 U771 ( .A(n1072), .B(n1073), .Z(n1071) );
NOR2_X1 U772 ( .A1(n1074), .A2(G953), .ZN(n1073) );
NOR2_X1 U773 ( .A1(n1075), .A2(n1076), .ZN(n1072) );
XOR2_X1 U774 ( .A(n1077), .B(n1078), .Z(n1076) );
XOR2_X1 U775 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND2_X1 U776 ( .A1(KEYINPUT52), .A2(n1081), .ZN(n1080) );
NAND2_X1 U777 ( .A1(n1082), .A2(n1083), .ZN(n1079) );
NAND2_X1 U778 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U779 ( .A1(KEYINPUT49), .A2(n1086), .ZN(n1085) );
NAND2_X1 U780 ( .A1(KEYINPUT50), .A2(n1087), .ZN(n1086) );
NAND2_X1 U781 ( .A1(n1088), .A2(n1089), .ZN(n1082) );
NAND2_X1 U782 ( .A1(KEYINPUT50), .A2(n1090), .ZN(n1089) );
NAND2_X1 U783 ( .A1(n1091), .A2(KEYINPUT49), .ZN(n1090) );
INV_X1 U784 ( .A(n1084), .ZN(n1091) );
XNOR2_X1 U785 ( .A(n1092), .B(n1093), .ZN(n1084) );
XNOR2_X1 U786 ( .A(G131), .B(G134), .ZN(n1092) );
XOR2_X1 U787 ( .A(KEYINPUT13), .B(G140), .Z(n1077) );
NOR2_X1 U788 ( .A1(n1094), .A2(n1095), .ZN(n1070) );
AND2_X1 U789 ( .A1(G227), .A2(G900), .ZN(n1094) );
XOR2_X1 U790 ( .A(n1096), .B(n1097), .Z(G69) );
NOR3_X1 U791 ( .A1(n1098), .A2(KEYINPUT61), .A3(n1099), .ZN(n1097) );
AND2_X1 U792 ( .A1(G224), .A2(G898), .ZN(n1099) );
XNOR2_X1 U793 ( .A(G953), .B(KEYINPUT43), .ZN(n1098) );
NAND2_X1 U794 ( .A1(n1100), .A2(n1101), .ZN(n1096) );
NAND3_X1 U795 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
NAND2_X1 U796 ( .A1(G953), .A2(n1105), .ZN(n1103) );
XOR2_X1 U797 ( .A(n1106), .B(KEYINPUT22), .Z(n1102) );
OR2_X1 U798 ( .A1(n1106), .A2(n1104), .ZN(n1100) );
XOR2_X1 U799 ( .A(n1107), .B(n1108), .Z(n1104) );
XNOR2_X1 U800 ( .A(n1109), .B(G110), .ZN(n1108) );
NAND2_X1 U801 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
NAND2_X1 U802 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XOR2_X1 U803 ( .A(n1114), .B(KEYINPUT6), .Z(n1110) );
OR2_X1 U804 ( .A1(n1112), .A2(n1113), .ZN(n1114) );
NAND2_X1 U805 ( .A1(n1095), .A2(n1115), .ZN(n1106) );
NAND2_X1 U806 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NOR2_X1 U807 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XOR2_X1 U808 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR3_X1 U809 ( .A1(n1122), .A2(KEYINPUT24), .A3(n1123), .ZN(n1120) );
NOR2_X1 U810 ( .A1(n1118), .A2(n1124), .ZN(G63) );
XOR2_X1 U811 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND2_X1 U812 ( .A1(n1127), .A2(G478), .ZN(n1125) );
NOR2_X1 U813 ( .A1(n1118), .A2(n1128), .ZN(G60) );
XOR2_X1 U814 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR3_X1 U815 ( .A1(n1122), .A2(KEYINPUT25), .A3(n1065), .ZN(n1129) );
XNOR2_X1 U816 ( .A(G104), .B(n1131), .ZN(G6) );
NOR2_X1 U817 ( .A1(n1118), .A2(n1132), .ZN(G57) );
XOR2_X1 U818 ( .A(n1133), .B(n1134), .Z(n1132) );
XNOR2_X1 U819 ( .A(n1135), .B(n1136), .ZN(n1134) );
XOR2_X1 U820 ( .A(n1137), .B(n1138), .Z(n1133) );
XOR2_X1 U821 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR3_X1 U822 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1140) );
NOR2_X1 U823 ( .A1(KEYINPUT48), .A2(n1144), .ZN(n1143) );
AND2_X1 U824 ( .A1(n1145), .A2(n1017), .ZN(n1144) );
AND2_X1 U825 ( .A1(n1122), .A2(KEYINPUT48), .ZN(n1142) );
NAND2_X1 U826 ( .A1(KEYINPUT0), .A2(n1146), .ZN(n1139) );
NAND2_X1 U827 ( .A1(KEYINPUT41), .A2(n1147), .ZN(n1137) );
NOR2_X1 U828 ( .A1(n1118), .A2(n1148), .ZN(G54) );
XOR2_X1 U829 ( .A(n1149), .B(n1150), .Z(n1148) );
XNOR2_X1 U830 ( .A(n1151), .B(n1152), .ZN(n1150) );
NAND2_X1 U831 ( .A1(n1127), .A2(G469), .ZN(n1151) );
INV_X1 U832 ( .A(n1122), .ZN(n1127) );
XNOR2_X1 U833 ( .A(n1153), .B(n1154), .ZN(n1149) );
NOR2_X1 U834 ( .A1(KEYINPUT12), .A2(n1155), .ZN(n1154) );
NOR2_X1 U835 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U836 ( .A(KEYINPUT26), .B(n1158), .Z(n1157) );
NOR2_X1 U837 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
AND2_X1 U838 ( .A1(n1160), .A2(n1159), .ZN(n1156) );
XOR2_X1 U839 ( .A(G110), .B(n1161), .Z(n1160) );
NOR2_X1 U840 ( .A1(G140), .A2(KEYINPUT16), .ZN(n1161) );
NOR2_X1 U841 ( .A1(KEYINPUT30), .A2(n1162), .ZN(n1153) );
XOR2_X1 U842 ( .A(n1163), .B(n1164), .Z(n1162) );
XNOR2_X1 U843 ( .A(n1088), .B(n1165), .ZN(n1164) );
XOR2_X1 U844 ( .A(KEYINPUT58), .B(KEYINPUT10), .Z(n1163) );
NOR2_X1 U845 ( .A1(n1118), .A2(n1166), .ZN(G51) );
NOR2_X1 U846 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U847 ( .A(n1169), .B(n1170), .Z(n1168) );
NAND2_X1 U848 ( .A1(KEYINPUT38), .A2(n1171), .ZN(n1170) );
OR2_X1 U849 ( .A1(n1122), .A2(n1067), .ZN(n1169) );
NAND2_X1 U850 ( .A1(G902), .A2(n1017), .ZN(n1122) );
NAND3_X1 U851 ( .A1(n1116), .A2(n1172), .A3(n1074), .ZN(n1017) );
AND4_X1 U852 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1074) );
AND4_X1 U853 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
NOR2_X1 U854 ( .A1(n1181), .A2(n1182), .ZN(n1175) );
NOR2_X1 U855 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
INV_X1 U856 ( .A(KEYINPUT14), .ZN(n1183) );
NOR4_X1 U857 ( .A1(KEYINPUT14), .A2(n1185), .A3(n1028), .A4(n1186), .ZN(n1181) );
INV_X1 U858 ( .A(n1187), .ZN(n1028) );
NAND3_X1 U859 ( .A1(n1049), .A2(n1034), .A3(n1040), .ZN(n1185) );
NAND2_X1 U860 ( .A1(n1188), .A2(n1189), .ZN(n1173) );
NAND2_X1 U861 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
XNOR2_X1 U862 ( .A(n1192), .B(KEYINPUT37), .ZN(n1190) );
XOR2_X1 U863 ( .A(KEYINPUT17), .B(n1117), .Z(n1172) );
AND4_X1 U864 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1117) );
NAND2_X1 U865 ( .A1(n1197), .A2(n1034), .ZN(n1193) );
XOR2_X1 U866 ( .A(n1198), .B(KEYINPUT2), .Z(n1197) );
AND4_X1 U867 ( .A1(n1131), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1116) );
NAND2_X1 U868 ( .A1(n1202), .A2(n1034), .ZN(n1201) );
XOR2_X1 U869 ( .A(n1011), .B(KEYINPUT62), .Z(n1202) );
NAND4_X1 U870 ( .A1(n1043), .A2(n1048), .A3(n1047), .A4(n1203), .ZN(n1011) );
NAND2_X1 U871 ( .A1(n1204), .A2(n1205), .ZN(n1199) );
XNOR2_X1 U872 ( .A(n1039), .B(KEYINPUT59), .ZN(n1204) );
NAND4_X1 U873 ( .A1(n1049), .A2(n1206), .A3(n1047), .A4(n1203), .ZN(n1131) );
NOR2_X1 U874 ( .A1(KEYINPUT38), .A2(n1171), .ZN(n1167) );
XOR2_X1 U875 ( .A(n1207), .B(n1208), .Z(n1171) );
XNOR2_X1 U876 ( .A(n1209), .B(n1210), .ZN(n1208) );
NAND2_X1 U877 ( .A1(n1211), .A2(KEYINPUT21), .ZN(n1210) );
XNOR2_X1 U878 ( .A(G125), .B(KEYINPUT35), .ZN(n1211) );
XNOR2_X1 U879 ( .A(n1212), .B(n1135), .ZN(n1207) );
NOR2_X1 U880 ( .A1(n1095), .A2(G952), .ZN(n1118) );
XNOR2_X1 U881 ( .A(G146), .B(n1174), .ZN(G48) );
NAND3_X1 U882 ( .A1(n1206), .A2(n1213), .A3(n1049), .ZN(n1174) );
XNOR2_X1 U883 ( .A(G143), .B(n1180), .ZN(G45) );
NAND4_X1 U884 ( .A1(n1214), .A2(n1206), .A3(n1059), .A4(n1215), .ZN(n1180) );
XNOR2_X1 U885 ( .A(G140), .B(n1216), .ZN(G42) );
NAND2_X1 U886 ( .A1(n1217), .A2(n1192), .ZN(n1216) );
AND2_X1 U887 ( .A1(n1218), .A2(n1043), .ZN(n1192) );
XNOR2_X1 U888 ( .A(n1188), .B(KEYINPUT34), .ZN(n1217) );
XNOR2_X1 U889 ( .A(G137), .B(n1179), .ZN(G39) );
NAND4_X1 U890 ( .A1(n1024), .A2(n1188), .A3(n1213), .A4(n1043), .ZN(n1179) );
XNOR2_X1 U891 ( .A(G134), .B(n1178), .ZN(G36) );
NAND4_X1 U892 ( .A1(n1188), .A2(n1214), .A3(n1043), .A4(n1048), .ZN(n1178) );
NAND2_X1 U893 ( .A1(n1219), .A2(n1220), .ZN(G33) );
NAND2_X1 U894 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
XOR2_X1 U895 ( .A(KEYINPUT46), .B(n1223), .Z(n1219) );
NOR2_X1 U896 ( .A1(n1221), .A2(n1222), .ZN(n1223) );
AND2_X1 U897 ( .A1(n1188), .A2(n1224), .ZN(n1221) );
XNOR2_X1 U898 ( .A(KEYINPUT63), .B(n1191), .ZN(n1224) );
NAND3_X1 U899 ( .A1(n1214), .A2(n1043), .A3(n1049), .ZN(n1191) );
AND2_X1 U900 ( .A1(n1039), .A2(n1186), .ZN(n1214) );
INV_X1 U901 ( .A(n1038), .ZN(n1188) );
NAND2_X1 U902 ( .A1(n1225), .A2(n1036), .ZN(n1038) );
XNOR2_X1 U903 ( .A(G128), .B(n1177), .ZN(G30) );
NAND3_X1 U904 ( .A1(n1213), .A2(n1048), .A3(n1206), .ZN(n1177) );
AND3_X1 U905 ( .A1(n1186), .A2(n1226), .A3(n1069), .ZN(n1213) );
XOR2_X1 U906 ( .A(G101), .B(n1227), .Z(G3) );
AND2_X1 U907 ( .A1(n1039), .A2(n1205), .ZN(n1227) );
XOR2_X1 U908 ( .A(n1184), .B(n1228), .Z(G27) );
XNOR2_X1 U909 ( .A(G125), .B(KEYINPUT42), .ZN(n1228) );
NAND3_X1 U910 ( .A1(n1218), .A2(n1034), .A3(n1187), .ZN(n1184) );
AND3_X1 U911 ( .A1(n1049), .A2(n1186), .A3(n1040), .ZN(n1218) );
NAND2_X1 U912 ( .A1(n1019), .A2(n1229), .ZN(n1186) );
NAND3_X1 U913 ( .A1(G902), .A2(n1230), .A3(n1075), .ZN(n1229) );
AND2_X1 U914 ( .A1(G953), .A2(n1231), .ZN(n1075) );
XOR2_X1 U915 ( .A(KEYINPUT7), .B(G900), .Z(n1231) );
XNOR2_X1 U916 ( .A(G122), .B(n1194), .ZN(G24) );
NAND4_X1 U917 ( .A1(n1232), .A2(n1047), .A3(n1059), .A4(n1215), .ZN(n1194) );
NOR2_X1 U918 ( .A1(n1226), .A2(n1069), .ZN(n1047) );
XOR2_X1 U919 ( .A(G119), .B(n1233), .Z(G21) );
NOR2_X1 U920 ( .A1(n1012), .A2(n1198), .ZN(n1233) );
NAND3_X1 U921 ( .A1(n1187), .A2(n1024), .A3(n1234), .ZN(n1198) );
AND3_X1 U922 ( .A1(n1069), .A2(n1203), .A3(n1226), .ZN(n1234) );
XNOR2_X1 U923 ( .A(G116), .B(n1195), .ZN(G18) );
NAND3_X1 U924 ( .A1(n1039), .A2(n1048), .A3(n1232), .ZN(n1195) );
NOR2_X1 U925 ( .A1(n1215), .A2(n1235), .ZN(n1048) );
XNOR2_X1 U926 ( .A(G113), .B(n1196), .ZN(G15) );
NAND3_X1 U927 ( .A1(n1049), .A2(n1039), .A3(n1232), .ZN(n1196) );
AND3_X1 U928 ( .A1(n1034), .A2(n1203), .A3(n1187), .ZN(n1232) );
NOR2_X1 U929 ( .A1(n1044), .A2(n1055), .ZN(n1187) );
INV_X1 U930 ( .A(n1045), .ZN(n1055) );
AND2_X1 U931 ( .A1(n1062), .A2(n1069), .ZN(n1039) );
AND2_X1 U932 ( .A1(n1235), .A2(n1215), .ZN(n1049) );
INV_X1 U933 ( .A(n1059), .ZN(n1235) );
XNOR2_X1 U934 ( .A(G110), .B(n1200), .ZN(G12) );
NAND2_X1 U935 ( .A1(n1205), .A2(n1040), .ZN(n1200) );
NOR2_X1 U936 ( .A1(n1069), .A2(n1062), .ZN(n1040) );
INV_X1 U937 ( .A(n1226), .ZN(n1062) );
NAND3_X1 U938 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1226) );
NAND2_X1 U939 ( .A1(n1239), .A2(n1121), .ZN(n1238) );
OR3_X1 U940 ( .A1(n1121), .A2(n1239), .A3(G902), .ZN(n1237) );
NOR2_X1 U941 ( .A1(n1123), .A2(G234), .ZN(n1239) );
INV_X1 U942 ( .A(G217), .ZN(n1123) );
XNOR2_X1 U943 ( .A(n1240), .B(n1241), .ZN(n1121) );
XOR2_X1 U944 ( .A(n1093), .B(n1242), .Z(n1241) );
XOR2_X1 U945 ( .A(n1243), .B(n1244), .Z(n1240) );
NOR3_X1 U946 ( .A1(n1245), .A2(G953), .A3(n1246), .ZN(n1244) );
XNOR2_X1 U947 ( .A(G234), .B(KEYINPUT3), .ZN(n1246) );
INV_X1 U948 ( .A(G221), .ZN(n1245) );
XOR2_X1 U949 ( .A(n1247), .B(G146), .Z(n1243) );
NAND2_X1 U950 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
OR2_X1 U951 ( .A1(n1250), .A2(G110), .ZN(n1249) );
XOR2_X1 U952 ( .A(n1251), .B(KEYINPUT60), .Z(n1248) );
NAND2_X1 U953 ( .A1(G110), .A2(n1250), .ZN(n1251) );
XNOR2_X1 U954 ( .A(G119), .B(n1252), .ZN(n1250) );
NAND2_X1 U955 ( .A1(G902), .A2(G217), .ZN(n1236) );
XOR2_X1 U956 ( .A(n1253), .B(n1141), .Z(n1069) );
INV_X1 U957 ( .A(G472), .ZN(n1141) );
NAND2_X1 U958 ( .A1(n1254), .A2(n1145), .ZN(n1253) );
XOR2_X1 U959 ( .A(n1255), .B(n1256), .Z(n1254) );
XNOR2_X1 U960 ( .A(n1147), .B(n1136), .ZN(n1256) );
XNOR2_X1 U961 ( .A(n1112), .B(KEYINPUT36), .ZN(n1147) );
XOR2_X1 U962 ( .A(n1257), .B(n1258), .Z(n1255) );
XNOR2_X1 U963 ( .A(n1259), .B(KEYINPUT32), .ZN(n1258) );
NAND2_X1 U964 ( .A1(KEYINPUT20), .A2(n1146), .ZN(n1259) );
XOR2_X1 U965 ( .A(n1260), .B(n1261), .Z(n1146) );
NAND2_X1 U966 ( .A1(n1262), .A2(G210), .ZN(n1260) );
NAND2_X1 U967 ( .A1(KEYINPUT40), .A2(n1135), .ZN(n1257) );
INV_X1 U968 ( .A(n1263), .ZN(n1135) );
AND3_X1 U969 ( .A1(n1206), .A2(n1203), .A3(n1024), .ZN(n1205) );
NOR2_X1 U970 ( .A1(n1059), .A2(n1215), .ZN(n1024) );
NAND2_X1 U971 ( .A1(n1264), .A2(n1058), .ZN(n1215) );
NAND2_X1 U972 ( .A1(n1063), .A2(n1065), .ZN(n1058) );
OR2_X1 U973 ( .A1(n1065), .A2(n1063), .ZN(n1264) );
NOR2_X1 U974 ( .A1(n1130), .A2(G902), .ZN(n1063) );
XNOR2_X1 U975 ( .A(n1265), .B(n1266), .ZN(n1130) );
XOR2_X1 U976 ( .A(n1267), .B(n1268), .Z(n1266) );
XNOR2_X1 U977 ( .A(n1109), .B(G113), .ZN(n1268) );
XNOR2_X1 U978 ( .A(KEYINPUT51), .B(n1222), .ZN(n1267) );
INV_X1 U979 ( .A(G131), .ZN(n1222) );
XOR2_X1 U980 ( .A(n1269), .B(n1270), .Z(n1265) );
XOR2_X1 U981 ( .A(n1271), .B(n1242), .Z(n1270) );
XNOR2_X1 U982 ( .A(G140), .B(n1081), .ZN(n1242) );
INV_X1 U983 ( .A(G125), .ZN(n1081) );
XNOR2_X1 U984 ( .A(n1272), .B(n1273), .ZN(n1269) );
INV_X1 U985 ( .A(G104), .ZN(n1273) );
NAND2_X1 U986 ( .A1(n1262), .A2(G214), .ZN(n1272) );
NOR2_X1 U987 ( .A1(G953), .A2(G237), .ZN(n1262) );
INV_X1 U988 ( .A(G475), .ZN(n1065) );
XNOR2_X1 U989 ( .A(n1274), .B(G478), .ZN(n1059) );
NAND2_X1 U990 ( .A1(n1126), .A2(n1275), .ZN(n1274) );
XNOR2_X1 U991 ( .A(KEYINPUT56), .B(n1145), .ZN(n1275) );
XOR2_X1 U992 ( .A(n1276), .B(n1277), .Z(n1126) );
XOR2_X1 U993 ( .A(n1278), .B(n1279), .Z(n1277) );
AND3_X1 U994 ( .A1(G217), .A2(n1095), .A3(G234), .ZN(n1279) );
NOR2_X1 U995 ( .A1(KEYINPUT1), .A2(n1280), .ZN(n1278) );
NOR2_X1 U996 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XOR2_X1 U997 ( .A(n1283), .B(KEYINPUT45), .Z(n1282) );
NAND2_X1 U998 ( .A1(G107), .A2(n1284), .ZN(n1283) );
NOR2_X1 U999 ( .A1(G107), .A2(n1284), .ZN(n1281) );
XOR2_X1 U1000 ( .A(G116), .B(G122), .Z(n1284) );
XNOR2_X1 U1001 ( .A(G128), .B(n1285), .ZN(n1276) );
XNOR2_X1 U1002 ( .A(G143), .B(n1286), .ZN(n1285) );
NAND2_X1 U1003 ( .A1(n1019), .A2(n1287), .ZN(n1203) );
NAND4_X1 U1004 ( .A1(G902), .A2(G953), .A3(n1230), .A4(n1105), .ZN(n1287) );
INV_X1 U1005 ( .A(G898), .ZN(n1105) );
NAND3_X1 U1006 ( .A1(n1230), .A2(n1095), .A3(G952), .ZN(n1019) );
NAND2_X1 U1007 ( .A1(G237), .A2(G234), .ZN(n1230) );
AND2_X1 U1008 ( .A1(n1034), .A2(n1043), .ZN(n1206) );
AND2_X1 U1009 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U1010 ( .A1(G221), .A2(n1288), .ZN(n1045) );
NAND2_X1 U1011 ( .A1(G234), .A2(n1145), .ZN(n1288) );
NAND3_X1 U1012 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1044) );
INV_X1 U1013 ( .A(n1056), .ZN(n1291) );
NOR2_X1 U1014 ( .A1(n1292), .A2(G469), .ZN(n1056) );
OR2_X1 U1015 ( .A1(G469), .A2(KEYINPUT44), .ZN(n1290) );
NAND2_X1 U1016 ( .A1(n1293), .A2(KEYINPUT44), .ZN(n1289) );
INV_X1 U1017 ( .A(n1057), .ZN(n1293) );
NAND2_X1 U1018 ( .A1(G469), .A2(n1292), .ZN(n1057) );
NAND2_X1 U1019 ( .A1(n1294), .A2(n1145), .ZN(n1292) );
XOR2_X1 U1020 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U1021 ( .A(n1297), .B(n1298), .ZN(n1296) );
XNOR2_X1 U1022 ( .A(n1299), .B(n1300), .ZN(n1298) );
INV_X1 U1023 ( .A(n1152), .ZN(n1300) );
XOR2_X1 U1024 ( .A(n1136), .B(KEYINPUT47), .Z(n1152) );
XOR2_X1 U1025 ( .A(G131), .B(n1301), .Z(n1136) );
NOR3_X1 U1026 ( .A1(KEYINPUT28), .A2(n1302), .A3(n1303), .ZN(n1301) );
NOR2_X1 U1027 ( .A1(n1286), .A2(n1304), .ZN(n1303) );
XNOR2_X1 U1028 ( .A(n1093), .B(KEYINPUT39), .ZN(n1304) );
INV_X1 U1029 ( .A(G134), .ZN(n1286) );
NOR2_X1 U1030 ( .A1(G134), .A2(n1305), .ZN(n1302) );
XNOR2_X1 U1031 ( .A(n1093), .B(KEYINPUT27), .ZN(n1305) );
XOR2_X1 U1032 ( .A(G137), .B(KEYINPUT9), .Z(n1093) );
NAND2_X1 U1033 ( .A1(n1306), .A2(KEYINPUT15), .ZN(n1299) );
XNOR2_X1 U1034 ( .A(n1159), .B(KEYINPUT57), .ZN(n1306) );
AND2_X1 U1035 ( .A1(G227), .A2(n1307), .ZN(n1159) );
XNOR2_X1 U1036 ( .A(KEYINPUT54), .B(n1095), .ZN(n1307) );
XOR2_X1 U1037 ( .A(n1308), .B(n1309), .Z(n1295) );
XOR2_X1 U1038 ( .A(KEYINPUT10), .B(G140), .Z(n1309) );
NOR2_X1 U1039 ( .A1(KEYINPUT31), .A2(n1088), .ZN(n1308) );
INV_X1 U1040 ( .A(n1087), .ZN(n1088) );
XOR2_X1 U1041 ( .A(G128), .B(n1271), .Z(n1087) );
INV_X1 U1042 ( .A(n1012), .ZN(n1034) );
NAND2_X1 U1043 ( .A1(n1310), .A2(n1036), .ZN(n1012) );
NAND2_X1 U1044 ( .A1(G214), .A2(n1311), .ZN(n1036) );
XNOR2_X1 U1045 ( .A(KEYINPUT23), .B(n1225), .ZN(n1310) );
INV_X1 U1046 ( .A(n1035), .ZN(n1225) );
XNOR2_X1 U1047 ( .A(n1068), .B(n1312), .ZN(n1035) );
NOR2_X1 U1048 ( .A1(KEYINPUT29), .A2(n1067), .ZN(n1312) );
NAND2_X1 U1049 ( .A1(G210), .A2(n1311), .ZN(n1067) );
NAND2_X1 U1050 ( .A1(n1313), .A2(n1145), .ZN(n1311) );
INV_X1 U1051 ( .A(G237), .ZN(n1313) );
NAND2_X1 U1052 ( .A1(n1314), .A2(n1145), .ZN(n1068) );
INV_X1 U1053 ( .A(G902), .ZN(n1145) );
XOR2_X1 U1054 ( .A(n1315), .B(n1212), .Z(n1314) );
XOR2_X1 U1055 ( .A(n1316), .B(n1297), .Z(n1212) );
XNOR2_X1 U1056 ( .A(G110), .B(n1113), .ZN(n1297) );
INV_X1 U1057 ( .A(n1165), .ZN(n1113) );
XNOR2_X1 U1058 ( .A(n1317), .B(n1261), .ZN(n1165) );
XOR2_X1 U1059 ( .A(G101), .B(KEYINPUT18), .Z(n1261) );
XNOR2_X1 U1060 ( .A(G104), .B(G107), .ZN(n1317) );
XNOR2_X1 U1061 ( .A(n1318), .B(n1109), .ZN(n1316) );
INV_X1 U1062 ( .A(G122), .ZN(n1109) );
NAND2_X1 U1063 ( .A1(KEYINPUT5), .A2(n1112), .ZN(n1318) );
XNOR2_X1 U1064 ( .A(G113), .B(n1319), .ZN(n1112) );
XOR2_X1 U1065 ( .A(G119), .B(G116), .Z(n1319) );
NAND2_X1 U1066 ( .A1(n1320), .A2(n1321), .ZN(n1315) );
NAND2_X1 U1067 ( .A1(n1322), .A2(n1209), .ZN(n1321) );
XOR2_X1 U1068 ( .A(KEYINPUT8), .B(n1323), .Z(n1320) );
NOR2_X1 U1069 ( .A1(n1209), .A2(n1322), .ZN(n1323) );
XNOR2_X1 U1070 ( .A(G125), .B(n1263), .ZN(n1322) );
XOR2_X1 U1071 ( .A(n1324), .B(n1252), .Z(n1263) );
INV_X1 U1072 ( .A(G128), .ZN(n1252) );
NAND2_X1 U1073 ( .A1(KEYINPUT4), .A2(n1271), .ZN(n1324) );
XOR2_X1 U1074 ( .A(G143), .B(G146), .Z(n1271) );
AND2_X1 U1075 ( .A1(G224), .A2(n1325), .ZN(n1209) );
XNOR2_X1 U1076 ( .A(KEYINPUT33), .B(n1095), .ZN(n1325) );
INV_X1 U1077 ( .A(G953), .ZN(n1095) );
endmodule


