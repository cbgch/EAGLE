//Key = 0110111000110100010100110111000111000011111100111101100100011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
n1436, n1437, n1438, n1439, n1440;

NAND2_X1 U793 ( .A1(n1096), .A2(n1097), .ZN(G9) );
NAND2_X1 U794 ( .A1(G107), .A2(n1098), .ZN(n1097) );
XOR2_X1 U795 ( .A(n1099), .B(KEYINPUT63), .Z(n1096) );
OR2_X1 U796 ( .A1(n1098), .A2(G107), .ZN(n1099) );
NAND3_X1 U797 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1098) );
XNOR2_X1 U798 ( .A(n1103), .B(KEYINPUT5), .ZN(n1102) );
NOR2_X1 U799 ( .A1(n1104), .A2(n1105), .ZN(G75) );
NOR4_X1 U800 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1105) );
NOR3_X1 U801 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1108) );
NOR2_X1 U802 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR2_X1 U803 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR3_X1 U804 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1115) );
NOR2_X1 U805 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U806 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
XNOR2_X1 U807 ( .A(n1124), .B(KEYINPUT49), .ZN(n1123) );
NOR2_X1 U808 ( .A1(n1125), .A2(n1126), .ZN(n1122) );
XOR2_X1 U809 ( .A(n1127), .B(KEYINPUT12), .Z(n1125) );
NOR3_X1 U810 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1118) );
XNOR2_X1 U811 ( .A(KEYINPUT21), .B(n1131), .ZN(n1130) );
NOR2_X1 U812 ( .A1(n1132), .A2(n1133), .ZN(n1117) );
NOR3_X1 U813 ( .A1(n1121), .A2(n1134), .A3(n1132), .ZN(n1113) );
NOR2_X1 U814 ( .A1(n1101), .A2(n1135), .ZN(n1134) );
NAND4_X1 U815 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1106) );
NAND4_X1 U816 ( .A1(n1140), .A2(n1131), .A3(n1103), .A4(n1141), .ZN(n1137) );
NOR2_X1 U817 ( .A1(n1116), .A2(n1110), .ZN(n1141) );
INV_X1 U818 ( .A(n1142), .ZN(n1116) );
XOR2_X1 U819 ( .A(KEYINPUT0), .B(n1143), .Z(n1140) );
NOR2_X1 U820 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND4_X1 U821 ( .A1(n1146), .A2(n1147), .A3(n1142), .A4(n1148), .ZN(n1136) );
NOR2_X1 U822 ( .A1(n1110), .A2(n1149), .ZN(n1148) );
XNOR2_X1 U823 ( .A(KEYINPUT46), .B(n1121), .ZN(n1149) );
XNOR2_X1 U824 ( .A(n1132), .B(KEYINPUT53), .ZN(n1146) );
INV_X1 U825 ( .A(n1131), .ZN(n1132) );
NOR3_X1 U826 ( .A1(n1150), .A2(G953), .A3(G952), .ZN(n1104) );
INV_X1 U827 ( .A(n1138), .ZN(n1150) );
NAND4_X1 U828 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1138) );
NOR4_X1 U829 ( .A1(n1112), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1154) );
XNOR2_X1 U830 ( .A(G472), .B(n1158), .ZN(n1157) );
XNOR2_X1 U831 ( .A(n1159), .B(n1160), .ZN(n1156) );
NAND2_X1 U832 ( .A1(KEYINPUT39), .A2(n1161), .ZN(n1160) );
NOR2_X1 U833 ( .A1(n1162), .A2(n1163), .ZN(n1153) );
NAND2_X1 U834 ( .A1(G475), .A2(n1164), .ZN(n1152) );
XOR2_X1 U835 ( .A(n1165), .B(n1166), .Z(n1151) );
NAND2_X1 U836 ( .A1(KEYINPUT59), .A2(n1167), .ZN(n1166) );
NAND2_X1 U837 ( .A1(n1168), .A2(n1169), .ZN(G72) );
NAND2_X1 U838 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U839 ( .A(KEYINPUT60), .B(n1172), .Z(n1168) );
NOR2_X1 U840 ( .A1(n1170), .A2(n1173), .ZN(n1172) );
XNOR2_X1 U841 ( .A(n1174), .B(n1171), .ZN(n1173) );
NAND2_X1 U842 ( .A1(n1175), .A2(n1176), .ZN(n1171) );
NAND2_X1 U843 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XNOR2_X1 U844 ( .A(KEYINPUT30), .B(n1139), .ZN(n1177) );
XOR2_X1 U845 ( .A(n1179), .B(n1180), .Z(n1175) );
XNOR2_X1 U846 ( .A(n1181), .B(n1182), .ZN(n1180) );
NAND2_X1 U847 ( .A1(KEYINPUT23), .A2(n1183), .ZN(n1182) );
NAND2_X1 U848 ( .A1(KEYINPUT47), .A2(n1184), .ZN(n1181) );
XNOR2_X1 U849 ( .A(n1185), .B(n1186), .ZN(n1179) );
NAND2_X1 U850 ( .A1(n1187), .A2(n1188), .ZN(n1185) );
NAND2_X1 U851 ( .A1(G140), .A2(n1189), .ZN(n1188) );
XOR2_X1 U852 ( .A(KEYINPUT17), .B(n1190), .Z(n1187) );
NOR2_X1 U853 ( .A1(G140), .A2(n1189), .ZN(n1190) );
NAND2_X1 U854 ( .A1(KEYINPUT10), .A2(n1109), .ZN(n1174) );
AND2_X1 U855 ( .A1(G953), .A2(n1191), .ZN(n1170) );
NAND2_X1 U856 ( .A1(G900), .A2(G227), .ZN(n1191) );
XOR2_X1 U857 ( .A(n1192), .B(n1193), .Z(G69) );
NAND2_X1 U858 ( .A1(G953), .A2(n1194), .ZN(n1193) );
NAND2_X1 U859 ( .A1(G898), .A2(G224), .ZN(n1194) );
NAND2_X1 U860 ( .A1(KEYINPUT42), .A2(n1195), .ZN(n1192) );
XOR2_X1 U861 ( .A(n1196), .B(n1197), .Z(n1195) );
NAND2_X1 U862 ( .A1(n1139), .A2(n1198), .ZN(n1197) );
NAND2_X1 U863 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND2_X1 U864 ( .A1(n1201), .A2(n1202), .ZN(n1196) );
NAND2_X1 U865 ( .A1(G953), .A2(n1203), .ZN(n1202) );
XOR2_X1 U866 ( .A(n1204), .B(n1205), .Z(n1201) );
NAND2_X1 U867 ( .A1(n1206), .A2(n1207), .ZN(n1204) );
NAND2_X1 U868 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XOR2_X1 U869 ( .A(n1210), .B(KEYINPUT3), .Z(n1206) );
NAND2_X1 U870 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NOR2_X1 U871 ( .A1(n1213), .A2(n1214), .ZN(G66) );
NOR3_X1 U872 ( .A1(n1159), .A2(n1215), .A3(n1216), .ZN(n1214) );
AND3_X1 U873 ( .A1(n1217), .A2(n1161), .A3(n1218), .ZN(n1216) );
NOR2_X1 U874 ( .A1(n1219), .A2(n1217), .ZN(n1215) );
NOR2_X1 U875 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NOR2_X1 U876 ( .A1(n1213), .A2(n1222), .ZN(G63) );
XOR2_X1 U877 ( .A(n1223), .B(n1224), .Z(n1222) );
NAND2_X1 U878 ( .A1(n1218), .A2(G478), .ZN(n1223) );
NOR2_X1 U879 ( .A1(n1213), .A2(n1225), .ZN(G60) );
XOR2_X1 U880 ( .A(n1226), .B(n1227), .Z(n1225) );
NAND2_X1 U881 ( .A1(n1218), .A2(G475), .ZN(n1226) );
XNOR2_X1 U882 ( .A(G104), .B(n1228), .ZN(G6) );
NAND4_X1 U883 ( .A1(n1229), .A2(n1135), .A3(n1230), .A4(n1103), .ZN(n1228) );
NOR2_X1 U884 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XNOR2_X1 U885 ( .A(n1233), .B(KEYINPUT35), .ZN(n1229) );
NOR2_X1 U886 ( .A1(n1213), .A2(n1234), .ZN(G57) );
XOR2_X1 U887 ( .A(n1235), .B(n1236), .Z(n1234) );
XNOR2_X1 U888 ( .A(n1237), .B(n1238), .ZN(n1235) );
NAND2_X1 U889 ( .A1(n1218), .A2(G472), .ZN(n1237) );
NOR2_X1 U890 ( .A1(n1239), .A2(n1240), .ZN(G54) );
XOR2_X1 U891 ( .A(n1241), .B(n1242), .Z(n1240) );
XNOR2_X1 U892 ( .A(n1243), .B(n1244), .ZN(n1242) );
NAND2_X1 U893 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND3_X1 U894 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(n1246) );
INV_X1 U895 ( .A(KEYINPUT61), .ZN(n1249) );
NAND2_X1 U896 ( .A1(n1250), .A2(KEYINPUT61), .ZN(n1245) );
XOR2_X1 U897 ( .A(n1251), .B(n1252), .Z(n1241) );
NOR2_X1 U898 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NOR4_X1 U899 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1254) );
NOR2_X1 U900 ( .A1(KEYINPUT57), .A2(G110), .ZN(n1258) );
NOR2_X1 U901 ( .A1(KEYINPUT22), .A2(n1259), .ZN(n1256) );
NOR2_X1 U902 ( .A1(n1260), .A2(n1261), .ZN(n1255) );
NOR3_X1 U903 ( .A1(n1262), .A2(KEYINPUT57), .A3(G110), .ZN(n1253) );
NOR3_X1 U904 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1262) );
NOR2_X1 U905 ( .A1(n1260), .A2(n1266), .ZN(n1265) );
INV_X1 U906 ( .A(KEYINPUT22), .ZN(n1260) );
NOR2_X1 U907 ( .A1(KEYINPUT22), .A2(n1267), .ZN(n1264) );
XOR2_X1 U908 ( .A(n1268), .B(KEYINPUT50), .Z(n1251) );
NAND2_X1 U909 ( .A1(n1218), .A2(G469), .ZN(n1268) );
NOR2_X1 U910 ( .A1(n1269), .A2(n1139), .ZN(n1239) );
XNOR2_X1 U911 ( .A(G952), .B(KEYINPUT13), .ZN(n1269) );
NOR2_X1 U912 ( .A1(n1213), .A2(n1270), .ZN(G51) );
XOR2_X1 U913 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U914 ( .A(n1273), .B(n1274), .Z(n1272) );
NAND2_X1 U915 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NAND2_X1 U916 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
XOR2_X1 U917 ( .A(KEYINPUT6), .B(n1279), .Z(n1275) );
NOR2_X1 U918 ( .A1(n1277), .A2(n1278), .ZN(n1279) );
NAND2_X1 U919 ( .A1(n1218), .A2(n1280), .ZN(n1273) );
INV_X1 U920 ( .A(n1167), .ZN(n1280) );
NOR2_X1 U921 ( .A1(n1281), .A2(n1220), .ZN(n1218) );
NOR2_X1 U922 ( .A1(n1107), .A2(n1282), .ZN(n1220) );
XOR2_X1 U923 ( .A(KEYINPUT44), .B(n1109), .Z(n1282) );
NAND4_X1 U924 ( .A1(n1283), .A2(n1284), .A3(n1285), .A4(n1286), .ZN(n1109) );
AND4_X1 U925 ( .A1(n1287), .A2(n1288), .A3(n1289), .A4(n1290), .ZN(n1286) );
NOR2_X1 U926 ( .A1(n1291), .A2(n1292), .ZN(n1285) );
NAND2_X1 U927 ( .A1(n1199), .A2(n1293), .ZN(n1107) );
XNOR2_X1 U928 ( .A(KEYINPUT41), .B(n1200), .ZN(n1293) );
NAND3_X1 U929 ( .A1(n1100), .A2(n1103), .A3(n1135), .ZN(n1200) );
AND4_X1 U930 ( .A1(n1294), .A2(n1295), .A3(n1296), .A4(n1297), .ZN(n1199) );
NOR4_X1 U931 ( .A1(n1298), .A2(n1299), .A3(n1300), .A4(n1301), .ZN(n1297) );
INV_X1 U932 ( .A(n1302), .ZN(n1298) );
OR2_X1 U933 ( .A1(n1303), .A2(KEYINPUT45), .ZN(n1296) );
NAND2_X1 U934 ( .A1(n1103), .A2(n1304), .ZN(n1294) );
NAND2_X1 U935 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND4_X1 U936 ( .A1(KEYINPUT45), .A2(n1233), .A3(n1307), .A4(n1308), .ZN(n1306) );
NAND2_X1 U937 ( .A1(n1100), .A2(n1101), .ZN(n1305) );
NOR2_X1 U938 ( .A1(n1139), .A2(G952), .ZN(n1213) );
XNOR2_X1 U939 ( .A(G146), .B(n1289), .ZN(G48) );
NAND3_X1 U940 ( .A1(n1309), .A2(n1135), .A3(n1310), .ZN(n1289) );
XNOR2_X1 U941 ( .A(G143), .B(n1288), .ZN(G45) );
NAND3_X1 U942 ( .A1(n1307), .A2(n1311), .A3(n1310), .ZN(n1288) );
NAND3_X1 U943 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(G42) );
NAND2_X1 U944 ( .A1(KEYINPUT24), .A2(n1315), .ZN(n1314) );
NAND3_X1 U945 ( .A1(G140), .A2(n1316), .A3(n1283), .ZN(n1313) );
NAND2_X1 U946 ( .A1(n1317), .A2(n1318), .ZN(n1312) );
NAND2_X1 U947 ( .A1(n1319), .A2(n1316), .ZN(n1318) );
INV_X1 U948 ( .A(KEYINPUT24), .ZN(n1316) );
XNOR2_X1 U949 ( .A(G140), .B(KEYINPUT51), .ZN(n1319) );
INV_X1 U950 ( .A(n1283), .ZN(n1317) );
NAND2_X1 U951 ( .A1(n1320), .A2(n1321), .ZN(n1283) );
XNOR2_X1 U952 ( .A(G137), .B(n1284), .ZN(G39) );
NAND4_X1 U953 ( .A1(n1129), .A2(n1320), .A3(n1322), .A4(n1142), .ZN(n1284) );
XOR2_X1 U954 ( .A(n1323), .B(n1292), .Z(G36) );
AND3_X1 U955 ( .A1(n1311), .A2(n1101), .A3(n1320), .ZN(n1292) );
NAND2_X1 U956 ( .A1(KEYINPUT2), .A2(n1324), .ZN(n1323) );
NAND3_X1 U957 ( .A1(n1325), .A2(n1326), .A3(n1327), .ZN(G33) );
NAND2_X1 U958 ( .A1(n1291), .A2(n1186), .ZN(n1327) );
NAND2_X1 U959 ( .A1(n1328), .A2(n1329), .ZN(n1326) );
INV_X1 U960 ( .A(KEYINPUT11), .ZN(n1329) );
NAND2_X1 U961 ( .A1(n1330), .A2(G131), .ZN(n1328) );
XNOR2_X1 U962 ( .A(n1291), .B(KEYINPUT20), .ZN(n1330) );
NAND2_X1 U963 ( .A1(KEYINPUT11), .A2(n1331), .ZN(n1325) );
NAND2_X1 U964 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
OR3_X1 U965 ( .A1(n1186), .A2(n1291), .A3(KEYINPUT20), .ZN(n1333) );
INV_X1 U966 ( .A(G131), .ZN(n1186) );
NAND2_X1 U967 ( .A1(KEYINPUT20), .A2(n1291), .ZN(n1332) );
AND3_X1 U968 ( .A1(n1135), .A2(n1311), .A3(n1320), .ZN(n1291) );
AND2_X1 U969 ( .A1(n1310), .A2(n1131), .ZN(n1320) );
NAND2_X1 U970 ( .A1(n1334), .A2(n1335), .ZN(n1131) );
OR3_X1 U971 ( .A1(n1127), .A2(n1163), .A3(KEYINPUT12), .ZN(n1335) );
INV_X1 U972 ( .A(n1126), .ZN(n1163) );
NAND2_X1 U973 ( .A1(KEYINPUT12), .A2(n1124), .ZN(n1334) );
XNOR2_X1 U974 ( .A(G128), .B(n1287), .ZN(G30) );
NAND3_X1 U975 ( .A1(n1309), .A2(n1101), .A3(n1310), .ZN(n1287) );
AND2_X1 U976 ( .A1(n1147), .A2(n1336), .ZN(n1310) );
INV_X1 U977 ( .A(n1232), .ZN(n1147) );
XNOR2_X1 U978 ( .A(G101), .B(n1295), .ZN(G3) );
NAND3_X1 U979 ( .A1(n1142), .A2(n1100), .A3(n1311), .ZN(n1295) );
INV_X1 U980 ( .A(n1133), .ZN(n1311) );
XNOR2_X1 U981 ( .A(G125), .B(n1290), .ZN(G27) );
NAND4_X1 U982 ( .A1(n1321), .A2(n1308), .A3(n1124), .A4(n1336), .ZN(n1290) );
NAND2_X1 U983 ( .A1(n1110), .A2(n1337), .ZN(n1336) );
NAND4_X1 U984 ( .A1(G953), .A2(G902), .A3(n1338), .A4(n1178), .ZN(n1337) );
INV_X1 U985 ( .A(G900), .ZN(n1178) );
AND3_X1 U986 ( .A1(n1322), .A2(n1339), .A3(n1135), .ZN(n1321) );
XNOR2_X1 U987 ( .A(G122), .B(n1303), .ZN(G24) );
NAND4_X1 U988 ( .A1(n1307), .A2(n1308), .A3(n1103), .A4(n1340), .ZN(n1303) );
INV_X1 U989 ( .A(n1121), .ZN(n1103) );
NAND2_X1 U990 ( .A1(n1341), .A2(n1339), .ZN(n1121) );
AND3_X1 U991 ( .A1(n1155), .A2(n1342), .A3(n1124), .ZN(n1307) );
XOR2_X1 U992 ( .A(n1343), .B(n1344), .Z(G21) );
XNOR2_X1 U993 ( .A(G119), .B(KEYINPUT34), .ZN(n1344) );
NAND2_X1 U994 ( .A1(KEYINPUT26), .A2(n1301), .ZN(n1343) );
AND4_X1 U995 ( .A1(n1309), .A2(n1142), .A3(n1308), .A4(n1340), .ZN(n1301) );
INV_X1 U996 ( .A(n1112), .ZN(n1308) );
NOR3_X1 U997 ( .A1(n1128), .A2(n1345), .A3(n1339), .ZN(n1309) );
XOR2_X1 U998 ( .A(G116), .B(n1300), .Z(G18) );
AND3_X1 U999 ( .A1(n1101), .A2(n1124), .A3(n1346), .ZN(n1300) );
NOR2_X1 U1000 ( .A1(n1342), .A2(n1347), .ZN(n1101) );
XOR2_X1 U1001 ( .A(n1299), .B(n1348), .Z(G15) );
NOR2_X1 U1002 ( .A1(KEYINPUT28), .A2(n1349), .ZN(n1348) );
INV_X1 U1003 ( .A(G113), .ZN(n1349) );
AND3_X1 U1004 ( .A1(n1135), .A2(n1350), .A3(n1346), .ZN(n1299) );
NOR3_X1 U1005 ( .A1(n1112), .A2(n1233), .A3(n1133), .ZN(n1346) );
NAND2_X1 U1006 ( .A1(n1129), .A2(n1341), .ZN(n1133) );
XNOR2_X1 U1007 ( .A(n1351), .B(KEYINPUT62), .ZN(n1341) );
INV_X1 U1008 ( .A(n1339), .ZN(n1129) );
NAND2_X1 U1009 ( .A1(n1352), .A2(n1145), .ZN(n1112) );
INV_X1 U1010 ( .A(n1144), .ZN(n1352) );
AND2_X1 U1011 ( .A1(n1347), .A2(n1342), .ZN(n1135) );
INV_X1 U1012 ( .A(n1155), .ZN(n1347) );
XNOR2_X1 U1013 ( .A(G110), .B(n1302), .ZN(G12) );
NAND4_X1 U1014 ( .A1(n1322), .A2(n1142), .A3(n1100), .A4(n1339), .ZN(n1302) );
XNOR2_X1 U1015 ( .A(n1353), .B(G472), .ZN(n1339) );
NAND2_X1 U1016 ( .A1(n1354), .A2(n1158), .ZN(n1353) );
NAND2_X1 U1017 ( .A1(n1355), .A2(n1281), .ZN(n1158) );
XOR2_X1 U1018 ( .A(n1356), .B(n1236), .Z(n1355) );
XNOR2_X1 U1019 ( .A(n1357), .B(n1358), .ZN(n1236) );
XOR2_X1 U1020 ( .A(G101), .B(n1277), .Z(n1358) );
XNOR2_X1 U1021 ( .A(n1209), .B(n1243), .ZN(n1357) );
NOR2_X1 U1022 ( .A1(KEYINPUT16), .A2(n1238), .ZN(n1356) );
NAND2_X1 U1023 ( .A1(n1359), .A2(G210), .ZN(n1238) );
XOR2_X1 U1024 ( .A(KEYINPUT40), .B(KEYINPUT18), .Z(n1354) );
NOR3_X1 U1025 ( .A1(n1231), .A2(n1233), .A3(n1232), .ZN(n1100) );
NAND2_X1 U1026 ( .A1(n1144), .A2(n1145), .ZN(n1232) );
NAND2_X1 U1027 ( .A1(G221), .A2(n1360), .ZN(n1145) );
XNOR2_X1 U1028 ( .A(n1361), .B(G469), .ZN(n1144) );
NAND2_X1 U1029 ( .A1(n1362), .A2(n1281), .ZN(n1361) );
XOR2_X1 U1030 ( .A(n1363), .B(n1364), .Z(n1362) );
XNOR2_X1 U1031 ( .A(n1250), .B(n1243), .ZN(n1364) );
XNOR2_X1 U1032 ( .A(n1365), .B(n1366), .ZN(n1243) );
NOR2_X1 U1033 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
NOR3_X1 U1034 ( .A1(KEYINPUT31), .A2(G137), .A3(n1324), .ZN(n1368) );
NOR2_X1 U1035 ( .A1(n1183), .A2(n1369), .ZN(n1367) );
INV_X1 U1036 ( .A(KEYINPUT31), .ZN(n1369) );
XNOR2_X1 U1037 ( .A(n1324), .B(G137), .ZN(n1183) );
XNOR2_X1 U1038 ( .A(G131), .B(KEYINPUT8), .ZN(n1365) );
XOR2_X1 U1039 ( .A(n1248), .B(n1247), .Z(n1250) );
INV_X1 U1040 ( .A(n1184), .ZN(n1247) );
XNOR2_X1 U1041 ( .A(n1370), .B(n1371), .ZN(n1184) );
NAND2_X1 U1042 ( .A1(KEYINPUT55), .A2(n1372), .ZN(n1370) );
NAND2_X1 U1043 ( .A1(n1373), .A2(n1374), .ZN(n1248) );
OR2_X1 U1044 ( .A1(n1375), .A2(G101), .ZN(n1374) );
XOR2_X1 U1045 ( .A(n1376), .B(KEYINPUT56), .Z(n1373) );
NAND2_X1 U1046 ( .A1(G101), .A2(n1375), .ZN(n1376) );
XNOR2_X1 U1047 ( .A(G104), .B(n1377), .ZN(n1375) );
NAND2_X1 U1048 ( .A1(n1378), .A2(n1379), .ZN(n1363) );
NAND2_X1 U1049 ( .A1(G110), .A2(n1380), .ZN(n1379) );
NAND2_X1 U1050 ( .A1(n1266), .A2(n1261), .ZN(n1380) );
INV_X1 U1051 ( .A(n1263), .ZN(n1261) );
NOR2_X1 U1052 ( .A1(n1267), .A2(G140), .ZN(n1263) );
INV_X1 U1053 ( .A(n1257), .ZN(n1266) );
NOR2_X1 U1054 ( .A1(n1315), .A2(n1259), .ZN(n1257) );
NAND2_X1 U1055 ( .A1(n1381), .A2(n1382), .ZN(n1378) );
XNOR2_X1 U1056 ( .A(G140), .B(n1259), .ZN(n1381) );
INV_X1 U1057 ( .A(n1267), .ZN(n1259) );
NAND2_X1 U1058 ( .A1(G227), .A2(n1139), .ZN(n1267) );
INV_X1 U1059 ( .A(n1340), .ZN(n1233) );
NAND2_X1 U1060 ( .A1(n1110), .A2(n1383), .ZN(n1340) );
NAND4_X1 U1061 ( .A1(G953), .A2(G902), .A3(n1338), .A4(n1203), .ZN(n1383) );
INV_X1 U1062 ( .A(G898), .ZN(n1203) );
NAND3_X1 U1063 ( .A1(n1338), .A2(n1139), .A3(G952), .ZN(n1110) );
NAND2_X1 U1064 ( .A1(G237), .A2(G234), .ZN(n1338) );
INV_X1 U1065 ( .A(n1350), .ZN(n1231) );
XOR2_X1 U1066 ( .A(n1124), .B(KEYINPUT36), .Z(n1350) );
INV_X1 U1067 ( .A(n1345), .ZN(n1124) );
NAND2_X1 U1068 ( .A1(n1127), .A2(n1126), .ZN(n1345) );
NAND2_X1 U1069 ( .A1(G214), .A2(n1384), .ZN(n1126) );
XNOR2_X1 U1070 ( .A(n1385), .B(n1167), .ZN(n1127) );
NAND2_X1 U1071 ( .A1(G210), .A2(n1384), .ZN(n1167) );
NAND2_X1 U1072 ( .A1(n1386), .A2(n1281), .ZN(n1384) );
INV_X1 U1073 ( .A(G237), .ZN(n1386) );
XOR2_X1 U1074 ( .A(n1165), .B(KEYINPUT48), .Z(n1385) );
NAND2_X1 U1075 ( .A1(n1387), .A2(n1281), .ZN(n1165) );
XNOR2_X1 U1076 ( .A(n1388), .B(n1278), .ZN(n1387) );
XOR2_X1 U1077 ( .A(n1189), .B(KEYINPUT15), .Z(n1278) );
XNOR2_X1 U1078 ( .A(n1271), .B(n1389), .ZN(n1388) );
NOR2_X1 U1079 ( .A1(n1277), .A2(KEYINPUT14), .ZN(n1389) );
AND2_X1 U1080 ( .A1(n1390), .A2(n1391), .ZN(n1277) );
NAND2_X1 U1081 ( .A1(n1372), .A2(n1371), .ZN(n1391) );
XOR2_X1 U1082 ( .A(KEYINPUT4), .B(n1392), .Z(n1390) );
NOR2_X1 U1083 ( .A1(n1372), .A2(n1371), .ZN(n1392) );
XNOR2_X1 U1084 ( .A(n1393), .B(n1205), .ZN(n1271) );
XNOR2_X1 U1085 ( .A(n1382), .B(n1394), .ZN(n1205) );
NOR2_X1 U1086 ( .A1(KEYINPUT7), .A2(n1395), .ZN(n1394) );
XOR2_X1 U1087 ( .A(n1396), .B(n1397), .Z(n1393) );
NOR2_X1 U1088 ( .A1(n1398), .A2(n1399), .ZN(n1397) );
XOR2_X1 U1089 ( .A(n1400), .B(KEYINPUT25), .Z(n1399) );
NAND2_X1 U1090 ( .A1(n1401), .A2(n1402), .ZN(n1400) );
NOR2_X1 U1091 ( .A1(n1402), .A2(n1401), .ZN(n1398) );
XNOR2_X1 U1092 ( .A(KEYINPUT9), .B(n1208), .ZN(n1401) );
INV_X1 U1093 ( .A(n1212), .ZN(n1208) );
XNOR2_X1 U1094 ( .A(n1403), .B(n1404), .ZN(n1212) );
XNOR2_X1 U1095 ( .A(G104), .B(n1405), .ZN(n1404) );
NAND2_X1 U1096 ( .A1(KEYINPUT1), .A2(n1377), .ZN(n1405) );
NAND2_X1 U1097 ( .A1(KEYINPUT43), .A2(G101), .ZN(n1403) );
XNOR2_X1 U1098 ( .A(KEYINPUT27), .B(n1211), .ZN(n1402) );
INV_X1 U1099 ( .A(n1209), .ZN(n1211) );
XOR2_X1 U1100 ( .A(G113), .B(n1406), .Z(n1209) );
XOR2_X1 U1101 ( .A(G119), .B(G116), .Z(n1406) );
NAND2_X1 U1102 ( .A1(G224), .A2(n1139), .ZN(n1396) );
NOR2_X1 U1103 ( .A1(n1155), .A2(n1342), .ZN(n1142) );
NAND3_X1 U1104 ( .A1(n1407), .A2(n1408), .A3(n1409), .ZN(n1342) );
INV_X1 U1105 ( .A(n1162), .ZN(n1409) );
NOR2_X1 U1106 ( .A1(n1164), .A2(G475), .ZN(n1162) );
OR2_X1 U1107 ( .A1(n1410), .A2(G475), .ZN(n1408) );
NAND3_X1 U1108 ( .A1(n1164), .A2(n1410), .A3(G475), .ZN(n1407) );
INV_X1 U1109 ( .A(KEYINPUT54), .ZN(n1410) );
NAND2_X1 U1110 ( .A1(n1227), .A2(n1281), .ZN(n1164) );
XNOR2_X1 U1111 ( .A(n1411), .B(n1412), .ZN(n1227) );
XOR2_X1 U1112 ( .A(n1413), .B(n1414), .Z(n1412) );
XNOR2_X1 U1113 ( .A(n1395), .B(G113), .ZN(n1414) );
INV_X1 U1114 ( .A(G122), .ZN(n1395) );
XNOR2_X1 U1115 ( .A(n1315), .B(G131), .ZN(n1413) );
XOR2_X1 U1116 ( .A(n1415), .B(n1416), .Z(n1411) );
XOR2_X1 U1117 ( .A(n1417), .B(n1371), .Z(n1416) );
XOR2_X1 U1118 ( .A(G143), .B(G146), .Z(n1371) );
NOR2_X1 U1119 ( .A1(KEYINPUT37), .A2(n1189), .ZN(n1417) );
XNOR2_X1 U1120 ( .A(n1418), .B(n1419), .ZN(n1415) );
INV_X1 U1121 ( .A(G104), .ZN(n1419) );
NAND2_X1 U1122 ( .A1(n1359), .A2(G214), .ZN(n1418) );
NOR2_X1 U1123 ( .A1(G953), .A2(G237), .ZN(n1359) );
XNOR2_X1 U1124 ( .A(n1420), .B(G478), .ZN(n1155) );
NAND2_X1 U1125 ( .A1(n1421), .A2(n1281), .ZN(n1420) );
XNOR2_X1 U1126 ( .A(n1224), .B(KEYINPUT38), .ZN(n1421) );
XNOR2_X1 U1127 ( .A(n1422), .B(n1423), .ZN(n1224) );
XOR2_X1 U1128 ( .A(n1424), .B(n1425), .Z(n1423) );
XNOR2_X1 U1129 ( .A(n1377), .B(n1426), .ZN(n1425) );
NOR2_X1 U1130 ( .A1(KEYINPUT29), .A2(n1427), .ZN(n1426) );
XOR2_X1 U1131 ( .A(n1428), .B(n1429), .Z(n1427) );
XOR2_X1 U1132 ( .A(KEYINPUT19), .B(G143), .Z(n1429) );
NAND2_X1 U1133 ( .A1(KEYINPUT33), .A2(n1430), .ZN(n1428) );
INV_X1 U1134 ( .A(G107), .ZN(n1377) );
AND2_X1 U1135 ( .A1(n1431), .A2(G217), .ZN(n1424) );
XOR2_X1 U1136 ( .A(n1432), .B(n1433), .Z(n1422) );
XNOR2_X1 U1137 ( .A(KEYINPUT58), .B(n1324), .ZN(n1433) );
INV_X1 U1138 ( .A(G134), .ZN(n1324) );
XNOR2_X1 U1139 ( .A(G116), .B(G122), .ZN(n1432) );
INV_X1 U1140 ( .A(n1128), .ZN(n1322) );
XNOR2_X1 U1141 ( .A(n1351), .B(KEYINPUT32), .ZN(n1128) );
XNOR2_X1 U1142 ( .A(n1159), .B(n1161), .ZN(n1351) );
INV_X1 U1143 ( .A(n1221), .ZN(n1161) );
NAND2_X1 U1144 ( .A1(G217), .A2(n1360), .ZN(n1221) );
NAND2_X1 U1145 ( .A1(G234), .A2(n1281), .ZN(n1360) );
INV_X1 U1146 ( .A(G902), .ZN(n1281) );
NOR2_X1 U1147 ( .A1(n1217), .A2(G902), .ZN(n1159) );
XNOR2_X1 U1148 ( .A(n1434), .B(n1435), .ZN(n1217) );
XOR2_X1 U1149 ( .A(n1436), .B(n1437), .Z(n1435) );
XNOR2_X1 U1150 ( .A(G137), .B(n1189), .ZN(n1437) );
INV_X1 U1151 ( .A(G125), .ZN(n1189) );
XNOR2_X1 U1152 ( .A(G146), .B(n1315), .ZN(n1436) );
INV_X1 U1153 ( .A(G140), .ZN(n1315) );
XOR2_X1 U1154 ( .A(n1438), .B(n1439), .Z(n1434) );
XNOR2_X1 U1155 ( .A(G119), .B(n1382), .ZN(n1439) );
INV_X1 U1156 ( .A(G110), .ZN(n1382) );
XNOR2_X1 U1157 ( .A(n1440), .B(n1372), .ZN(n1438) );
INV_X1 U1158 ( .A(n1430), .ZN(n1372) );
XOR2_X1 U1159 ( .A(G128), .B(KEYINPUT52), .Z(n1430) );
NAND2_X1 U1160 ( .A1(n1431), .A2(G221), .ZN(n1440) );
AND2_X1 U1161 ( .A1(G234), .A2(n1139), .ZN(n1431) );
INV_X1 U1162 ( .A(G953), .ZN(n1139) );
endmodule


