//Key = 1111000010011100111100101011100001010000000101100101010001010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348;

XNOR2_X1 U730 ( .A(G107), .B(n1016), .ZN(G9) );
NOR2_X1 U731 ( .A1(n1017), .A2(n1018), .ZN(G75) );
XOR2_X1 U732 ( .A(n1019), .B(KEYINPUT35), .Z(n1018) );
OR3_X1 U733 ( .A1(G952), .A2(G953), .A3(n1020), .ZN(n1019) );
NOR4_X1 U734 ( .A1(n1021), .A2(n1022), .A3(G953), .A4(n1020), .ZN(n1017) );
AND4_X1 U735 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1020) );
NOR4_X1 U736 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
XOR2_X1 U737 ( .A(KEYINPUT61), .B(n1031), .Z(n1030) );
NOR2_X1 U738 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U739 ( .A1(G472), .A2(n1034), .ZN(n1033) );
XOR2_X1 U740 ( .A(n1035), .B(KEYINPUT32), .Z(n1034) );
XNOR2_X1 U741 ( .A(G469), .B(n1036), .ZN(n1029) );
NOR3_X1 U742 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1025) );
INV_X1 U743 ( .A(n1040), .ZN(n1039) );
XOR2_X1 U744 ( .A(n1041), .B(n1042), .Z(n1023) );
NOR2_X1 U745 ( .A1(G475), .A2(KEYINPUT38), .ZN(n1042) );
NOR2_X1 U746 ( .A1(n1043), .A2(n1044), .ZN(n1022) );
NOR2_X1 U747 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U748 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U749 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U751 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1051) );
NOR2_X1 U752 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U753 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U754 ( .A1(n1060), .A2(n1027), .ZN(n1058) );
NOR3_X1 U755 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1054) );
XOR2_X1 U756 ( .A(n1064), .B(KEYINPUT47), .Z(n1062) );
NOR2_X1 U757 ( .A1(n1065), .A2(n1064), .ZN(n1053) );
NOR3_X1 U758 ( .A1(n1057), .A2(n1066), .A3(n1064), .ZN(n1049) );
NOR2_X1 U759 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U760 ( .A1(n1069), .A2(n1024), .ZN(n1067) );
NOR4_X1 U761 ( .A1(n1070), .A2(n1064), .A3(n1057), .A4(n1052), .ZN(n1045) );
NOR2_X1 U762 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XOR2_X1 U763 ( .A(n1073), .B(KEYINPUT19), .Z(n1072) );
NAND3_X1 U764 ( .A1(n1074), .A2(G952), .A3(n1075), .ZN(n1021) );
XOR2_X1 U765 ( .A(n1076), .B(n1077), .Z(G72) );
XOR2_X1 U766 ( .A(n1078), .B(n1079), .Z(n1077) );
NAND2_X1 U767 ( .A1(G953), .A2(n1080), .ZN(n1079) );
NAND2_X1 U768 ( .A1(G900), .A2(G227), .ZN(n1080) );
NAND2_X1 U769 ( .A1(n1081), .A2(n1082), .ZN(n1078) );
NAND2_X1 U770 ( .A1(G953), .A2(n1083), .ZN(n1082) );
XOR2_X1 U771 ( .A(n1084), .B(n1085), .Z(n1081) );
XOR2_X1 U772 ( .A(n1086), .B(n1087), .Z(n1085) );
XOR2_X1 U773 ( .A(n1088), .B(G134), .Z(n1086) );
XOR2_X1 U774 ( .A(n1089), .B(KEYINPUT29), .Z(n1084) );
XNOR2_X1 U775 ( .A(KEYINPUT59), .B(KEYINPUT40), .ZN(n1089) );
NOR2_X1 U776 ( .A1(n1075), .A2(G953), .ZN(n1076) );
NAND2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(G69) );
NAND2_X1 U778 ( .A1(G953), .A2(n1092), .ZN(n1091) );
NAND2_X1 U779 ( .A1(n1093), .A2(G898), .ZN(n1092) );
XOR2_X1 U780 ( .A(n1094), .B(G224), .Z(n1093) );
NAND2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1090) );
XOR2_X1 U782 ( .A(n1097), .B(n1098), .Z(n1095) );
INV_X1 U783 ( .A(n1094), .ZN(n1098) );
XNOR2_X1 U784 ( .A(n1099), .B(n1100), .ZN(n1094) );
XOR2_X1 U785 ( .A(n1101), .B(n1102), .Z(n1099) );
NOR2_X1 U786 ( .A1(KEYINPUT37), .A2(n1103), .ZN(n1102) );
NAND2_X1 U787 ( .A1(KEYINPUT24), .A2(n1104), .ZN(n1097) );
NOR2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(G66) );
XOR2_X1 U789 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U790 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U791 ( .A1(n1105), .A2(n1111), .ZN(G63) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XOR2_X1 U793 ( .A(KEYINPUT62), .B(n1114), .Z(n1113) );
NOR2_X1 U794 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
AND2_X1 U795 ( .A1(n1116), .A2(n1115), .ZN(n1112) );
NAND2_X1 U796 ( .A1(n1117), .A2(G478), .ZN(n1116) );
NOR2_X1 U797 ( .A1(n1105), .A2(n1118), .ZN(G60) );
NOR3_X1 U798 ( .A1(n1041), .A2(n1119), .A3(n1120), .ZN(n1118) );
AND3_X1 U799 ( .A1(n1121), .A2(G475), .A3(n1117), .ZN(n1120) );
NOR2_X1 U800 ( .A1(n1122), .A2(n1121), .ZN(n1119) );
NOR2_X1 U801 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
INV_X1 U802 ( .A(G475), .ZN(n1124) );
NOR2_X1 U803 ( .A1(n1104), .A2(n1125), .ZN(n1123) );
XNOR2_X1 U804 ( .A(G104), .B(n1126), .ZN(G6) );
NAND4_X1 U805 ( .A1(n1127), .A2(n1128), .A3(KEYINPUT22), .A4(n1129), .ZN(n1126) );
NOR2_X1 U806 ( .A1(n1064), .A2(n1073), .ZN(n1129) );
NAND2_X1 U807 ( .A1(KEYINPUT46), .A2(n1130), .ZN(n1128) );
NAND2_X1 U808 ( .A1(n1131), .A2(n1132), .ZN(n1127) );
INV_X1 U809 ( .A(KEYINPUT46), .ZN(n1132) );
NAND3_X1 U810 ( .A1(n1133), .A2(n1065), .A3(n1068), .ZN(n1131) );
NOR2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(G57) );
XOR2_X1 U812 ( .A(KEYINPUT25), .B(n1105), .Z(n1135) );
NOR3_X1 U813 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1134) );
NOR2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR2_X1 U815 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
XOR2_X1 U816 ( .A(KEYINPUT7), .B(n1143), .Z(n1142) );
NOR3_X1 U817 ( .A1(n1144), .A2(n1143), .A3(n1141), .ZN(n1137) );
INV_X1 U818 ( .A(n1140), .ZN(n1144) );
XOR2_X1 U819 ( .A(n1145), .B(n1146), .Z(n1140) );
AND2_X1 U820 ( .A1(n1141), .A2(n1143), .ZN(n1136) );
XNOR2_X1 U821 ( .A(n1147), .B(n1148), .ZN(n1143) );
XOR2_X1 U822 ( .A(n1103), .B(n1149), .Z(n1147) );
NOR2_X1 U823 ( .A1(n1150), .A2(n1110), .ZN(n1149) );
INV_X1 U824 ( .A(KEYINPUT16), .ZN(n1141) );
NOR2_X1 U825 ( .A1(n1105), .A2(n1151), .ZN(G54) );
NOR2_X1 U826 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U827 ( .A(KEYINPUT4), .B(n1154), .Z(n1153) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
AND2_X1 U829 ( .A1(n1156), .A2(n1155), .ZN(n1152) );
XOR2_X1 U830 ( .A(n1157), .B(n1158), .Z(n1155) );
XOR2_X1 U831 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U832 ( .A(n1161), .B(n1162), .Z(n1160) );
NAND2_X1 U833 ( .A1(n1163), .A2(KEYINPUT49), .ZN(n1161) );
XNOR2_X1 U834 ( .A(n1164), .B(n1165), .ZN(n1163) );
NAND2_X1 U835 ( .A1(KEYINPUT63), .A2(n1166), .ZN(n1159) );
XOR2_X1 U836 ( .A(n1167), .B(n1168), .Z(n1157) );
XOR2_X1 U837 ( .A(n1169), .B(n1170), .Z(n1167) );
NOR2_X1 U838 ( .A1(KEYINPUT23), .A2(n1171), .ZN(n1170) );
NAND2_X1 U839 ( .A1(n1117), .A2(G469), .ZN(n1156) );
INV_X1 U840 ( .A(n1110), .ZN(n1117) );
NOR2_X1 U841 ( .A1(n1105), .A2(n1172), .ZN(G51) );
XOR2_X1 U842 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U843 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U844 ( .A(n1177), .B(n1178), .Z(n1173) );
NOR2_X1 U845 ( .A1(n1179), .A2(n1110), .ZN(n1178) );
NAND2_X1 U846 ( .A1(G902), .A2(n1180), .ZN(n1110) );
NAND2_X1 U847 ( .A1(n1075), .A2(n1074), .ZN(n1180) );
INV_X1 U848 ( .A(n1104), .ZN(n1074) );
NAND4_X1 U849 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1104) );
AND4_X1 U850 ( .A1(n1016), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1184) );
NAND3_X1 U851 ( .A1(n1071), .A2(n1188), .A3(n1189), .ZN(n1016) );
NOR2_X1 U852 ( .A1(n1190), .A2(n1191), .ZN(n1183) );
NOR2_X1 U853 ( .A1(n1065), .A2(n1192), .ZN(n1191) );
NOR3_X1 U854 ( .A1(n1073), .A2(n1064), .A3(n1130), .ZN(n1190) );
NAND4_X1 U855 ( .A1(n1059), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1181) );
NAND2_X1 U856 ( .A1(KEYINPUT57), .A2(n1130), .ZN(n1195) );
NAND2_X1 U857 ( .A1(n1196), .A2(n1197), .ZN(n1194) );
INV_X1 U858 ( .A(KEYINPUT57), .ZN(n1197) );
NAND3_X1 U859 ( .A1(n1133), .A2(n1198), .A3(n1199), .ZN(n1196) );
INV_X1 U860 ( .A(n1125), .ZN(n1075) );
NAND4_X1 U861 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1125) );
NOR4_X1 U862 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203) );
NOR3_X1 U863 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1202) );
NOR4_X1 U864 ( .A1(n1211), .A2(n1052), .A3(n1199), .A4(n1212), .ZN(n1210) );
AND2_X1 U865 ( .A1(n1211), .A2(n1213), .ZN(n1209) );
INV_X1 U866 ( .A(KEYINPUT10), .ZN(n1211) );
NOR3_X1 U867 ( .A1(n1214), .A2(n1215), .A3(n1057), .ZN(n1208) );
NOR2_X1 U868 ( .A1(n1096), .A2(G952), .ZN(n1105) );
XNOR2_X1 U869 ( .A(G146), .B(n1200), .ZN(G48) );
NAND3_X1 U870 ( .A1(n1216), .A2(n1199), .A3(n1217), .ZN(n1200) );
XNOR2_X1 U871 ( .A(n1201), .B(n1218), .ZN(G45) );
NOR2_X1 U872 ( .A1(KEYINPUT34), .A2(n1219), .ZN(n1218) );
OR4_X1 U873 ( .A1(n1220), .A2(n1214), .A3(n1065), .A4(n1221), .ZN(n1201) );
XOR2_X1 U874 ( .A(G140), .B(n1207), .Z(G42) );
NOR3_X1 U875 ( .A1(n1057), .A2(n1198), .A3(n1212), .ZN(n1207) );
XOR2_X1 U876 ( .A(n1206), .B(n1222), .Z(G39) );
NOR2_X1 U877 ( .A1(KEYINPUT54), .A2(n1223), .ZN(n1222) );
AND3_X1 U878 ( .A1(n1224), .A2(n1216), .A3(n1193), .ZN(n1206) );
XOR2_X1 U879 ( .A(G134), .B(n1225), .Z(G36) );
NOR3_X1 U880 ( .A1(n1226), .A2(n1215), .A3(n1214), .ZN(n1225) );
INV_X1 U881 ( .A(n1071), .ZN(n1215) );
XOR2_X1 U882 ( .A(KEYINPUT27), .B(n1224), .Z(n1226) );
XOR2_X1 U883 ( .A(G131), .B(n1205), .Z(G33) );
NOR3_X1 U884 ( .A1(n1214), .A2(n1057), .A3(n1073), .ZN(n1205) );
INV_X1 U885 ( .A(n1217), .ZN(n1073) );
INV_X1 U886 ( .A(n1224), .ZN(n1057) );
NOR2_X1 U887 ( .A1(n1063), .A2(n1037), .ZN(n1224) );
INV_X1 U888 ( .A(n1061), .ZN(n1037) );
NAND4_X1 U889 ( .A1(n1227), .A2(n1068), .A3(n1228), .A4(n1229), .ZN(n1214) );
XOR2_X1 U890 ( .A(G128), .B(n1204), .Z(G30) );
AND3_X1 U891 ( .A1(n1071), .A2(n1199), .A3(n1216), .ZN(n1204) );
AND4_X1 U892 ( .A1(n1068), .A2(n1027), .A3(n1228), .A4(n1229), .ZN(n1216) );
XOR2_X1 U893 ( .A(n1145), .B(n1182), .Z(G3) );
NAND4_X1 U894 ( .A1(n1193), .A2(n1189), .A3(n1227), .A4(n1229), .ZN(n1182) );
INV_X1 U895 ( .A(n1130), .ZN(n1189) );
XOR2_X1 U896 ( .A(G125), .B(n1213), .Z(G27) );
NOR3_X1 U897 ( .A1(n1212), .A2(n1065), .A3(n1052), .ZN(n1213) );
NAND3_X1 U898 ( .A1(n1217), .A2(n1228), .A3(n1059), .ZN(n1212) );
INV_X1 U899 ( .A(n1230), .ZN(n1059) );
NAND2_X1 U900 ( .A1(n1044), .A2(n1231), .ZN(n1228) );
NAND4_X1 U901 ( .A1(G902), .A2(G953), .A3(n1232), .A4(n1083), .ZN(n1231) );
INV_X1 U902 ( .A(G900), .ZN(n1083) );
XOR2_X1 U903 ( .A(G122), .B(n1233), .Z(G24) );
NOR2_X1 U904 ( .A1(n1065), .A2(n1234), .ZN(n1233) );
XNOR2_X1 U905 ( .A(KEYINPUT8), .B(n1192), .ZN(n1234) );
NAND3_X1 U906 ( .A1(n1235), .A2(n1188), .A3(n1236), .ZN(n1192) );
NOR3_X1 U907 ( .A1(n1220), .A2(n1237), .A3(n1221), .ZN(n1236) );
INV_X1 U908 ( .A(n1064), .ZN(n1188) );
NAND2_X1 U909 ( .A1(n1060), .A2(n1227), .ZN(n1064) );
INV_X1 U910 ( .A(n1052), .ZN(n1235) );
XNOR2_X1 U911 ( .A(G119), .B(n1187), .ZN(G21) );
NAND3_X1 U912 ( .A1(n1193), .A2(n1027), .A3(n1238), .ZN(n1187) );
XNOR2_X1 U913 ( .A(G116), .B(n1186), .ZN(G18) );
NAND3_X1 U914 ( .A1(n1227), .A2(n1071), .A3(n1238), .ZN(n1186) );
NOR2_X1 U915 ( .A1(n1220), .A2(n1239), .ZN(n1071) );
XOR2_X1 U916 ( .A(n1028), .B(KEYINPUT43), .Z(n1220) );
XNOR2_X1 U917 ( .A(G113), .B(n1185), .ZN(G15) );
NAND3_X1 U918 ( .A1(n1227), .A2(n1217), .A3(n1238), .ZN(n1185) );
NOR4_X1 U919 ( .A1(n1052), .A2(n1065), .A3(n1060), .A4(n1237), .ZN(n1238) );
INV_X1 U920 ( .A(n1133), .ZN(n1237) );
NAND2_X1 U921 ( .A1(n1024), .A2(n1240), .ZN(n1052) );
NOR2_X1 U922 ( .A1(n1028), .A2(n1221), .ZN(n1217) );
XOR2_X1 U923 ( .A(n1241), .B(n1242), .Z(G12) );
XOR2_X1 U924 ( .A(KEYINPUT42), .B(G110), .Z(n1242) );
NOR4_X1 U925 ( .A1(KEYINPUT44), .A2(n1130), .A3(n1048), .A4(n1230), .ZN(n1241) );
NAND2_X1 U926 ( .A1(n1060), .A2(n1027), .ZN(n1230) );
INV_X1 U927 ( .A(n1227), .ZN(n1027) );
XOR2_X1 U928 ( .A(n1109), .B(n1243), .Z(n1227) );
NOR2_X1 U929 ( .A1(n1107), .A2(n1244), .ZN(n1243) );
XOR2_X1 U930 ( .A(KEYINPUT39), .B(G902), .Z(n1244) );
NAND2_X1 U931 ( .A1(n1245), .A2(n1246), .ZN(n1107) );
NAND2_X1 U932 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND2_X1 U933 ( .A1(KEYINPUT53), .A2(n1249), .ZN(n1248) );
NAND2_X1 U934 ( .A1(KEYINPUT33), .A2(n1250), .ZN(n1249) );
INV_X1 U935 ( .A(n1251), .ZN(n1247) );
NAND2_X1 U936 ( .A1(n1252), .A2(n1253), .ZN(n1245) );
NAND2_X1 U937 ( .A1(KEYINPUT33), .A2(n1254), .ZN(n1253) );
NAND2_X1 U938 ( .A1(n1251), .A2(KEYINPUT53), .ZN(n1254) );
XOR2_X1 U939 ( .A(n1223), .B(n1255), .Z(n1251) );
NOR2_X1 U940 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
INV_X1 U941 ( .A(G221), .ZN(n1256) );
INV_X1 U942 ( .A(n1250), .ZN(n1252) );
XOR2_X1 U943 ( .A(n1258), .B(n1259), .Z(n1250) );
XOR2_X1 U944 ( .A(G119), .B(n1260), .Z(n1259) );
NOR2_X1 U945 ( .A1(KEYINPUT48), .A2(n1261), .ZN(n1260) );
XOR2_X1 U946 ( .A(n1262), .B(G125), .Z(n1261) );
NAND2_X1 U947 ( .A1(KEYINPUT12), .A2(G140), .ZN(n1262) );
XNOR2_X1 U948 ( .A(n1263), .B(n1166), .ZN(n1258) );
NAND2_X1 U949 ( .A1(G217), .A2(n1264), .ZN(n1109) );
INV_X1 U950 ( .A(n1229), .ZN(n1060) );
NAND2_X1 U951 ( .A1(n1265), .A2(n1266), .ZN(n1229) );
NAND2_X1 U952 ( .A1(n1267), .A2(n1150), .ZN(n1266) );
INV_X1 U953 ( .A(G472), .ZN(n1150) );
NAND2_X1 U954 ( .A1(KEYINPUT11), .A2(n1035), .ZN(n1267) );
NAND2_X1 U955 ( .A1(n1032), .A2(KEYINPUT11), .ZN(n1265) );
AND2_X1 U956 ( .A1(G472), .A2(n1035), .ZN(n1032) );
NAND2_X1 U957 ( .A1(n1268), .A2(n1269), .ZN(n1035) );
XOR2_X1 U958 ( .A(n1270), .B(n1271), .Z(n1268) );
XOR2_X1 U959 ( .A(n1272), .B(n1148), .Z(n1271) );
NAND2_X1 U960 ( .A1(KEYINPUT26), .A2(n1145), .ZN(n1272) );
XOR2_X1 U961 ( .A(n1146), .B(n1273), .Z(n1270) );
NOR2_X1 U962 ( .A1(KEYINPUT30), .A2(n1274), .ZN(n1273) );
NAND2_X1 U963 ( .A1(n1275), .A2(G210), .ZN(n1146) );
INV_X1 U964 ( .A(n1193), .ZN(n1048) );
NOR2_X1 U965 ( .A1(n1239), .A2(n1028), .ZN(n1193) );
XNOR2_X1 U966 ( .A(n1276), .B(G478), .ZN(n1028) );
NAND2_X1 U967 ( .A1(n1115), .A2(n1269), .ZN(n1276) );
XNOR2_X1 U968 ( .A(n1277), .B(n1278), .ZN(n1115) );
XOR2_X1 U969 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U970 ( .A(G107), .B(n1281), .Z(n1280) );
NOR2_X1 U971 ( .A1(n1257), .A2(n1282), .ZN(n1281) );
INV_X1 U972 ( .A(G217), .ZN(n1282) );
NAND2_X1 U973 ( .A1(G234), .A2(n1283), .ZN(n1257) );
XOR2_X1 U974 ( .A(G122), .B(G116), .Z(n1279) );
XOR2_X1 U975 ( .A(n1284), .B(n1285), .Z(n1277) );
XOR2_X1 U976 ( .A(KEYINPUT52), .B(G143), .Z(n1285) );
XNOR2_X1 U977 ( .A(G128), .B(G134), .ZN(n1284) );
INV_X1 U978 ( .A(n1221), .ZN(n1239) );
XNOR2_X1 U979 ( .A(n1041), .B(n1286), .ZN(n1221) );
XOR2_X1 U980 ( .A(KEYINPUT60), .B(G475), .Z(n1286) );
NOR2_X1 U981 ( .A1(n1121), .A2(G902), .ZN(n1041) );
XNOR2_X1 U982 ( .A(n1287), .B(n1288), .ZN(n1121) );
XOR2_X1 U983 ( .A(n1289), .B(n1290), .Z(n1288) );
XOR2_X1 U984 ( .A(G143), .B(G131), .Z(n1290) );
XOR2_X1 U985 ( .A(KEYINPUT41), .B(G146), .Z(n1289) );
XOR2_X1 U986 ( .A(n1291), .B(n1087), .Z(n1287) );
XOR2_X1 U987 ( .A(G125), .B(G140), .Z(n1087) );
XOR2_X1 U988 ( .A(n1292), .B(n1293), .Z(n1291) );
AND2_X1 U989 ( .A1(G214), .A2(n1275), .ZN(n1293) );
AND2_X1 U990 ( .A1(n1283), .A2(n1294), .ZN(n1275) );
NAND2_X1 U991 ( .A1(KEYINPUT51), .A2(n1295), .ZN(n1292) );
XOR2_X1 U992 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U993 ( .A(G122), .B(G113), .Z(n1297) );
NAND3_X1 U994 ( .A1(n1068), .A2(n1133), .A3(n1199), .ZN(n1130) );
INV_X1 U995 ( .A(n1065), .ZN(n1199) );
NAND2_X1 U996 ( .A1(n1063), .A2(n1061), .ZN(n1065) );
NAND2_X1 U997 ( .A1(G214), .A2(n1298), .ZN(n1061) );
NAND3_X1 U998 ( .A1(n1299), .A2(n1300), .A3(n1040), .ZN(n1063) );
NAND2_X1 U999 ( .A1(n1301), .A2(n1302), .ZN(n1040) );
NAND2_X1 U1000 ( .A1(n1038), .A2(n1303), .ZN(n1300) );
NOR2_X1 U1001 ( .A1(n1302), .A2(n1301), .ZN(n1038) );
INV_X1 U1002 ( .A(n1179), .ZN(n1301) );
NAND2_X1 U1003 ( .A1(G210), .A2(n1298), .ZN(n1179) );
NAND2_X1 U1004 ( .A1(n1294), .A2(n1269), .ZN(n1298) );
INV_X1 U1005 ( .A(G237), .ZN(n1294) );
NAND2_X1 U1006 ( .A1(n1304), .A2(n1302), .ZN(n1299) );
NAND3_X1 U1007 ( .A1(n1305), .A2(n1306), .A3(n1269), .ZN(n1302) );
NAND2_X1 U1008 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NAND2_X1 U1009 ( .A1(n1309), .A2(n1310), .ZN(n1305) );
INV_X1 U1010 ( .A(n1308), .ZN(n1310) );
XOR2_X1 U1011 ( .A(n1175), .B(KEYINPUT14), .Z(n1308) );
XOR2_X1 U1012 ( .A(n1311), .B(n1274), .Z(n1175) );
INV_X1 U1013 ( .A(n1103), .ZN(n1274) );
XOR2_X1 U1014 ( .A(n1312), .B(n1313), .Z(n1103) );
XOR2_X1 U1015 ( .A(KEYINPUT45), .B(G119), .Z(n1313) );
XNOR2_X1 U1016 ( .A(G113), .B(G116), .ZN(n1312) );
XOR2_X1 U1017 ( .A(n1101), .B(n1314), .Z(n1311) );
NOR2_X1 U1018 ( .A1(KEYINPUT5), .A2(n1100), .ZN(n1314) );
XNOR2_X1 U1019 ( .A(G122), .B(n1166), .ZN(n1100) );
NAND2_X1 U1020 ( .A1(n1315), .A2(n1316), .ZN(n1101) );
NAND2_X1 U1021 ( .A1(n1317), .A2(n1145), .ZN(n1316) );
XOR2_X1 U1022 ( .A(n1318), .B(KEYINPUT9), .Z(n1315) );
OR2_X1 U1023 ( .A1(n1145), .A2(n1317), .ZN(n1318) );
XNOR2_X1 U1024 ( .A(n1319), .B(KEYINPUT36), .ZN(n1317) );
INV_X1 U1025 ( .A(G101), .ZN(n1145) );
XNOR2_X1 U1026 ( .A(n1307), .B(KEYINPUT20), .ZN(n1309) );
XNOR2_X1 U1027 ( .A(n1320), .B(n1321), .ZN(n1307) );
XNOR2_X1 U1028 ( .A(KEYINPUT13), .B(n1177), .ZN(n1321) );
NAND2_X1 U1029 ( .A1(G224), .A2(n1283), .ZN(n1177) );
NAND2_X1 U1030 ( .A1(n1322), .A2(n1323), .ZN(n1320) );
NAND2_X1 U1031 ( .A1(KEYINPUT2), .A2(n1176), .ZN(n1323) );
XOR2_X1 U1032 ( .A(n1324), .B(n1165), .Z(n1176) );
OR3_X1 U1033 ( .A1(n1324), .A2(n1165), .A3(KEYINPUT2), .ZN(n1322) );
INV_X1 U1034 ( .A(G125), .ZN(n1324) );
INV_X1 U1035 ( .A(n1303), .ZN(n1304) );
XNOR2_X1 U1036 ( .A(KEYINPUT21), .B(KEYINPUT15), .ZN(n1303) );
NAND2_X1 U1037 ( .A1(n1044), .A2(n1325), .ZN(n1133) );
NAND4_X1 U1038 ( .A1(G902), .A2(G953), .A3(n1232), .A4(n1326), .ZN(n1325) );
INV_X1 U1039 ( .A(G898), .ZN(n1326) );
NAND3_X1 U1040 ( .A1(n1232), .A2(n1096), .A3(G952), .ZN(n1044) );
INV_X1 U1041 ( .A(G953), .ZN(n1096) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1232) );
INV_X1 U1043 ( .A(n1198), .ZN(n1068) );
NAND2_X1 U1044 ( .A1(n1069), .A2(n1024), .ZN(n1198) );
NAND2_X1 U1045 ( .A1(G221), .A2(n1264), .ZN(n1024) );
NAND2_X1 U1046 ( .A1(G234), .A2(n1269), .ZN(n1264) );
INV_X1 U1047 ( .A(n1240), .ZN(n1069) );
NAND2_X1 U1048 ( .A1(n1327), .A2(n1328), .ZN(n1240) );
NAND2_X1 U1049 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XNOR2_X1 U1050 ( .A(KEYINPUT58), .B(n1036), .ZN(n1330) );
XNOR2_X1 U1051 ( .A(G469), .B(KEYINPUT0), .ZN(n1329) );
NAND2_X1 U1052 ( .A1(n1331), .A2(n1332), .ZN(n1327) );
XOR2_X1 U1053 ( .A(n1036), .B(KEYINPUT58), .Z(n1332) );
NAND2_X1 U1054 ( .A1(n1333), .A2(n1269), .ZN(n1036) );
INV_X1 U1055 ( .A(G902), .ZN(n1269) );
XOR2_X1 U1056 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1057 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1058 ( .A(n1338), .B(KEYINPUT50), .Z(n1337) );
NAND3_X1 U1059 ( .A1(n1339), .A2(n1340), .A3(n1341), .ZN(n1338) );
NAND2_X1 U1060 ( .A1(KEYINPUT55), .A2(n1168), .ZN(n1341) );
NAND3_X1 U1061 ( .A1(n1342), .A2(n1343), .A3(n1166), .ZN(n1340) );
INV_X1 U1062 ( .A(KEYINPUT55), .ZN(n1343) );
OR2_X1 U1063 ( .A1(n1166), .A2(n1342), .ZN(n1339) );
NOR2_X1 U1064 ( .A1(KEYINPUT56), .A2(n1168), .ZN(n1342) );
XOR2_X1 U1065 ( .A(G140), .B(KEYINPUT31), .Z(n1168) );
XOR2_X1 U1066 ( .A(G110), .B(KEYINPUT28), .Z(n1166) );
NAND2_X1 U1067 ( .A1(KEYINPUT18), .A2(n1344), .ZN(n1336) );
INV_X1 U1068 ( .A(n1171), .ZN(n1344) );
NAND2_X1 U1069 ( .A1(G227), .A2(n1283), .ZN(n1171) );
XOR2_X1 U1070 ( .A(G953), .B(KEYINPUT17), .Z(n1283) );
XOR2_X1 U1071 ( .A(n1345), .B(n1164), .Z(n1334) );
XNOR2_X1 U1072 ( .A(n1319), .B(n1346), .ZN(n1164) );
XOR2_X1 U1073 ( .A(KEYINPUT59), .B(G101), .Z(n1346) );
XNOR2_X1 U1074 ( .A(G107), .B(n1296), .ZN(n1319) );
XOR2_X1 U1075 ( .A(G104), .B(KEYINPUT1), .Z(n1296) );
INV_X1 U1076 ( .A(n1148), .ZN(n1345) );
XOR2_X1 U1077 ( .A(n1162), .B(n1347), .Z(n1148) );
INV_X1 U1078 ( .A(n1088), .ZN(n1347) );
XOR2_X1 U1079 ( .A(n1169), .B(n1165), .Z(n1088) );
XNOR2_X1 U1080 ( .A(n1219), .B(n1263), .ZN(n1165) );
XOR2_X1 U1081 ( .A(G128), .B(G146), .Z(n1263) );
INV_X1 U1082 ( .A(G143), .ZN(n1219) );
XOR2_X1 U1083 ( .A(G131), .B(n1223), .Z(n1169) );
INV_X1 U1084 ( .A(G137), .ZN(n1223) );
NOR2_X1 U1085 ( .A1(n1348), .A2(G134), .ZN(n1162) );
INV_X1 U1086 ( .A(KEYINPUT3), .ZN(n1348) );
XNOR2_X1 U1087 ( .A(G469), .B(KEYINPUT6), .ZN(n1331) );
endmodule


