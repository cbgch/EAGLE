//Key = 1100010111101101110001001001111100010110111110111011100101010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314;

XOR2_X1 U725 ( .A(G107), .B(n1003), .Z(G9) );
NOR2_X1 U726 ( .A1(n1004), .A2(n1005), .ZN(G75) );
NOR4_X1 U727 ( .A1(G953), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1005) );
NOR2_X1 U728 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U729 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR4_X1 U730 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
NOR2_X1 U731 ( .A1(n1017), .A2(n1018), .ZN(n1014) );
NOR2_X1 U732 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR3_X1 U733 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NOR2_X1 U734 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U735 ( .A1(n1026), .A2(n1027), .ZN(n1019) );
NOR2_X1 U736 ( .A1(n1028), .A2(n1029), .ZN(n1013) );
NOR2_X1 U737 ( .A1(n1030), .A2(n1021), .ZN(n1028) );
NOR4_X1 U738 ( .A1(n1017), .A2(n1031), .A3(n1030), .A4(n1021), .ZN(n1011) );
NOR2_X1 U739 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U740 ( .A1(n1034), .A2(n1015), .ZN(n1033) );
NOR2_X1 U741 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U742 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U743 ( .A1(n1039), .A2(n1016), .ZN(n1032) );
NOR2_X1 U744 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR3_X1 U745 ( .A1(n1006), .A2(G953), .A3(G952), .ZN(n1004) );
AND4_X1 U746 ( .A1(n1042), .A2(n1027), .A3(n1043), .A4(n1044), .ZN(n1006) );
NOR4_X1 U747 ( .A1(n1045), .A2(n1017), .A3(n1046), .A4(n1047), .ZN(n1044) );
XNOR2_X1 U748 ( .A(n1048), .B(n1049), .ZN(n1047) );
NAND2_X1 U749 ( .A1(KEYINPUT28), .A2(n1050), .ZN(n1048) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1046) );
XNOR2_X1 U751 ( .A(KEYINPUT11), .B(n1053), .ZN(n1052) );
NOR2_X1 U752 ( .A1(n1054), .A2(n1055), .ZN(n1043) );
XOR2_X1 U753 ( .A(n1056), .B(n1057), .Z(n1054) );
NAND2_X1 U754 ( .A1(KEYINPUT43), .A2(n1058), .ZN(n1056) );
XOR2_X1 U755 ( .A(n1059), .B(n1060), .Z(G72) );
XNOR2_X1 U756 ( .A(n1061), .B(n1062), .ZN(n1060) );
NAND3_X1 U757 ( .A1(G953), .A2(n1063), .A3(KEYINPUT21), .ZN(n1062) );
NAND2_X1 U758 ( .A1(G900), .A2(G227), .ZN(n1063) );
NAND3_X1 U759 ( .A1(n1064), .A2(n1065), .A3(KEYINPUT7), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
XOR2_X1 U761 ( .A(n1068), .B(KEYINPUT58), .Z(n1066) );
XOR2_X1 U762 ( .A(KEYINPUT30), .B(G953), .Z(n1064) );
NAND2_X1 U763 ( .A1(n1069), .A2(n1070), .ZN(n1059) );
INV_X1 U764 ( .A(n1071), .ZN(n1070) );
XOR2_X1 U765 ( .A(n1072), .B(n1073), .Z(n1069) );
XOR2_X1 U766 ( .A(n1074), .B(n1075), .Z(n1073) );
XOR2_X1 U767 ( .A(n1076), .B(n1077), .Z(n1072) );
XOR2_X1 U768 ( .A(n1078), .B(n1079), .Z(G69) );
NAND2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U770 ( .A(n1082), .B(n1083), .Z(n1081) );
NAND2_X1 U771 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U772 ( .A1(n1086), .A2(n1087), .ZN(n1082) );
NAND2_X1 U773 ( .A1(G953), .A2(n1088), .ZN(n1087) );
XOR2_X1 U774 ( .A(n1089), .B(n1090), .Z(n1086) );
XOR2_X1 U775 ( .A(KEYINPUT44), .B(KEYINPUT4), .Z(n1080) );
NAND2_X1 U776 ( .A1(n1091), .A2(n1092), .ZN(n1078) );
NAND2_X1 U777 ( .A1(G898), .A2(G224), .ZN(n1092) );
XOR2_X1 U778 ( .A(KEYINPUT56), .B(G953), .Z(n1091) );
NOR2_X1 U779 ( .A1(n1093), .A2(n1094), .ZN(G66) );
XOR2_X1 U780 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U781 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
NOR2_X1 U782 ( .A1(n1093), .A2(n1099), .ZN(G63) );
XNOR2_X1 U783 ( .A(n1100), .B(n1101), .ZN(n1099) );
NOR2_X1 U784 ( .A1(n1102), .A2(n1098), .ZN(n1101) );
INV_X1 U785 ( .A(G478), .ZN(n1102) );
NOR2_X1 U786 ( .A1(n1093), .A2(n1103), .ZN(G60) );
NOR3_X1 U787 ( .A1(n1057), .A2(n1104), .A3(n1105), .ZN(n1103) );
NOR3_X1 U788 ( .A1(n1106), .A2(n1058), .A3(n1098), .ZN(n1105) );
INV_X1 U789 ( .A(n1107), .ZN(n1106) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1107), .ZN(n1104) );
AND2_X1 U791 ( .A1(n1008), .A2(G475), .ZN(n1108) );
XNOR2_X1 U792 ( .A(G104), .B(n1109), .ZN(G6) );
NAND4_X1 U793 ( .A1(KEYINPUT38), .A2(n1040), .A3(n1110), .A4(n1111), .ZN(n1109) );
NOR2_X1 U794 ( .A1(n1093), .A2(n1112), .ZN(G57) );
XOR2_X1 U795 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U796 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U797 ( .A(n1117), .B(n1118), .Z(n1113) );
XNOR2_X1 U798 ( .A(n1119), .B(KEYINPUT42), .ZN(n1118) );
NAND2_X1 U799 ( .A1(n1120), .A2(KEYINPUT10), .ZN(n1119) );
XNOR2_X1 U800 ( .A(n1121), .B(KEYINPUT13), .ZN(n1120) );
NOR2_X1 U801 ( .A1(n1050), .A2(n1098), .ZN(n1117) );
INV_X1 U802 ( .A(G472), .ZN(n1050) );
NOR2_X1 U803 ( .A1(n1093), .A2(n1122), .ZN(G54) );
XOR2_X1 U804 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U805 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U806 ( .A1(n1051), .A2(n1098), .ZN(n1126) );
INV_X1 U807 ( .A(G469), .ZN(n1051) );
NOR2_X1 U808 ( .A1(KEYINPUT39), .A2(n1127), .ZN(n1125) );
XOR2_X1 U809 ( .A(n1128), .B(KEYINPUT62), .Z(n1127) );
XNOR2_X1 U810 ( .A(n1129), .B(n1130), .ZN(n1123) );
NOR2_X1 U811 ( .A1(KEYINPUT23), .A2(n1131), .ZN(n1130) );
NOR2_X1 U812 ( .A1(n1093), .A2(n1132), .ZN(G51) );
XOR2_X1 U813 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U814 ( .A1(n1135), .A2(n1098), .ZN(n1134) );
NAND2_X1 U815 ( .A1(G902), .A2(n1008), .ZN(n1098) );
NAND3_X1 U816 ( .A1(n1136), .A2(n1068), .A3(n1067), .ZN(n1008) );
AND4_X1 U817 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1067) );
AND4_X1 U818 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1140) );
NAND2_X1 U819 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
INV_X1 U820 ( .A(n1147), .ZN(n1146) );
XOR2_X1 U821 ( .A(n1148), .B(KEYINPUT46), .Z(n1145) );
INV_X1 U822 ( .A(n1085), .ZN(n1136) );
NAND4_X1 U823 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1085) );
NOR4_X1 U824 ( .A1(n1153), .A2(n1003), .A3(n1154), .A4(n1155), .ZN(n1152) );
AND3_X1 U825 ( .A1(n1111), .A2(n1041), .A3(n1110), .ZN(n1003) );
NOR2_X1 U826 ( .A1(n1156), .A2(n1157), .ZN(n1151) );
AND3_X1 U827 ( .A1(n1040), .A2(n1111), .A3(n1110), .ZN(n1157) );
INV_X1 U828 ( .A(n1158), .ZN(n1110) );
INV_X1 U829 ( .A(n1159), .ZN(n1156) );
NAND2_X1 U830 ( .A1(n1160), .A2(n1161), .ZN(n1150) );
NAND2_X1 U831 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND3_X1 U832 ( .A1(n1164), .A2(n1111), .A3(KEYINPUT60), .ZN(n1163) );
INV_X1 U833 ( .A(n1165), .ZN(n1164) );
NAND2_X1 U834 ( .A1(n1166), .A2(n1167), .ZN(n1162) );
OR2_X1 U835 ( .A1(n1168), .A2(KEYINPUT60), .ZN(n1149) );
NOR2_X1 U836 ( .A1(KEYINPUT49), .A2(n1169), .ZN(n1133) );
XOR2_X1 U837 ( .A(n1170), .B(n1171), .Z(n1169) );
XNOR2_X1 U838 ( .A(n1172), .B(n1173), .ZN(n1171) );
NOR2_X1 U839 ( .A1(G125), .A2(KEYINPUT45), .ZN(n1172) );
NOR2_X1 U840 ( .A1(n1084), .A2(G952), .ZN(n1093) );
XOR2_X1 U841 ( .A(n1174), .B(n1141), .Z(G48) );
NAND3_X1 U842 ( .A1(n1175), .A2(n1040), .A3(n1166), .ZN(n1141) );
XOR2_X1 U843 ( .A(n1176), .B(n1137), .Z(G45) );
NAND3_X1 U844 ( .A1(n1165), .A2(n1036), .A3(n1175), .ZN(n1137) );
XOR2_X1 U845 ( .A(n1138), .B(n1177), .Z(G42) );
XNOR2_X1 U846 ( .A(G140), .B(KEYINPUT19), .ZN(n1177) );
NAND2_X1 U847 ( .A1(n1178), .A2(n1179), .ZN(n1138) );
XOR2_X1 U848 ( .A(n1180), .B(n1144), .Z(G39) );
NAND3_X1 U849 ( .A1(n1166), .A2(n1167), .A3(n1178), .ZN(n1144) );
XOR2_X1 U850 ( .A(G134), .B(n1181), .Z(G36) );
NOR2_X1 U851 ( .A1(KEYINPUT33), .A2(n1068), .ZN(n1181) );
NAND3_X1 U852 ( .A1(n1036), .A2(n1041), .A3(n1178), .ZN(n1068) );
XOR2_X1 U853 ( .A(n1143), .B(n1182), .Z(G33) );
XNOR2_X1 U854 ( .A(G131), .B(KEYINPUT2), .ZN(n1182) );
NAND3_X1 U855 ( .A1(n1040), .A2(n1036), .A3(n1178), .ZN(n1143) );
AND3_X1 U856 ( .A1(n1183), .A2(n1184), .A3(n1027), .ZN(n1178) );
INV_X1 U857 ( .A(n1030), .ZN(n1027) );
NAND2_X1 U858 ( .A1(n1185), .A2(n1025), .ZN(n1030) );
XOR2_X1 U859 ( .A(G128), .B(n1186), .Z(G30) );
NOR2_X1 U860 ( .A1(n1148), .A2(n1147), .ZN(n1186) );
NAND2_X1 U861 ( .A1(n1175), .A2(n1041), .ZN(n1147) );
AND3_X1 U862 ( .A1(n1023), .A2(n1184), .A3(n1183), .ZN(n1175) );
XOR2_X1 U863 ( .A(G101), .B(n1153), .Z(G3) );
NOR3_X1 U864 ( .A1(n1015), .A2(n1187), .A3(n1158), .ZN(n1153) );
XOR2_X1 U865 ( .A(n1188), .B(n1142), .Z(G27) );
NAND4_X1 U866 ( .A1(n1179), .A2(n1189), .A3(n1023), .A4(n1184), .ZN(n1142) );
NAND2_X1 U867 ( .A1(n1010), .A2(n1190), .ZN(n1184) );
NAND3_X1 U868 ( .A1(G902), .A2(n1191), .A3(n1071), .ZN(n1190) );
NOR2_X1 U869 ( .A1(n1084), .A2(G900), .ZN(n1071) );
XNOR2_X1 U870 ( .A(KEYINPUT47), .B(n1192), .ZN(n1191) );
AND3_X1 U871 ( .A1(n1193), .A2(n1055), .A3(n1040), .ZN(n1179) );
XOR2_X1 U872 ( .A(n1194), .B(n1168), .Z(G24) );
NAND3_X1 U873 ( .A1(n1111), .A2(n1165), .A3(n1160), .ZN(n1168) );
NAND2_X1 U874 ( .A1(n1195), .A2(n1196), .ZN(n1165) );
NAND2_X1 U875 ( .A1(n1040), .A2(n1197), .ZN(n1196) );
OR3_X1 U876 ( .A1(n1198), .A2(n1042), .A3(n1197), .ZN(n1195) );
INV_X1 U877 ( .A(n1016), .ZN(n1111) );
NAND2_X1 U878 ( .A1(n1199), .A2(n1193), .ZN(n1016) );
XOR2_X1 U879 ( .A(n1037), .B(KEYINPUT22), .Z(n1199) );
XNOR2_X1 U880 ( .A(G119), .B(n1200), .ZN(G21) );
NAND3_X1 U881 ( .A1(n1201), .A2(n1189), .A3(n1202), .ZN(n1200) );
NOR3_X1 U882 ( .A1(n1148), .A2(n1203), .A3(n1015), .ZN(n1202) );
XNOR2_X1 U883 ( .A(n1023), .B(KEYINPUT16), .ZN(n1201) );
XOR2_X1 U884 ( .A(n1204), .B(n1159), .Z(G18) );
NAND3_X1 U885 ( .A1(n1036), .A2(n1041), .A3(n1160), .ZN(n1159) );
AND3_X1 U886 ( .A1(n1023), .A2(n1205), .A3(n1189), .ZN(n1160) );
XOR2_X1 U887 ( .A(n1206), .B(KEYINPUT14), .Z(n1023) );
NAND2_X1 U888 ( .A1(n1207), .A2(n1208), .ZN(n1041) );
NAND2_X1 U889 ( .A1(n1167), .A2(n1197), .ZN(n1208) );
INV_X1 U890 ( .A(KEYINPUT52), .ZN(n1197) );
INV_X1 U891 ( .A(n1015), .ZN(n1167) );
NAND3_X1 U892 ( .A1(n1209), .A2(n1198), .A3(KEYINPUT52), .ZN(n1207) );
XOR2_X1 U893 ( .A(n1210), .B(n1211), .Z(G15) );
NAND2_X1 U894 ( .A1(KEYINPUT37), .A2(n1155), .ZN(n1211) );
AND4_X1 U895 ( .A1(n1189), .A2(n1040), .A3(n1212), .A4(n1206), .ZN(n1155) );
NOR2_X1 U896 ( .A1(n1203), .A2(n1187), .ZN(n1212) );
INV_X1 U897 ( .A(n1036), .ZN(n1187) );
NAND2_X1 U898 ( .A1(n1213), .A2(n1214), .ZN(n1036) );
OR3_X1 U899 ( .A1(n1193), .A2(n1055), .A3(KEYINPUT22), .ZN(n1214) );
NAND2_X1 U900 ( .A1(KEYINPUT22), .A2(n1166), .ZN(n1213) );
INV_X1 U901 ( .A(n1148), .ZN(n1166) );
NAND2_X1 U902 ( .A1(n1055), .A2(n1038), .ZN(n1148) );
INV_X1 U903 ( .A(n1037), .ZN(n1055) );
INV_X1 U904 ( .A(n1205), .ZN(n1203) );
NOR2_X1 U905 ( .A1(n1209), .A2(n1198), .ZN(n1040) );
INV_X1 U906 ( .A(n1042), .ZN(n1209) );
NOR2_X1 U907 ( .A1(n1021), .A2(n1017), .ZN(n1189) );
INV_X1 U908 ( .A(n1026), .ZN(n1021) );
XOR2_X1 U909 ( .A(G110), .B(n1154), .Z(G12) );
NOR4_X1 U910 ( .A1(n1158), .A2(n1015), .A3(n1038), .A4(n1037), .ZN(n1154) );
XNOR2_X1 U911 ( .A(n1215), .B(n1097), .ZN(n1037) );
NAND2_X1 U912 ( .A1(G217), .A2(n1216), .ZN(n1097) );
OR2_X1 U913 ( .A1(n1096), .A2(G902), .ZN(n1215) );
XNOR2_X1 U914 ( .A(n1217), .B(n1218), .ZN(n1096) );
XOR2_X1 U915 ( .A(n1219), .B(n1220), .Z(n1218) );
XOR2_X1 U916 ( .A(n1221), .B(G110), .Z(n1220) );
NAND2_X1 U917 ( .A1(KEYINPUT48), .A2(n1222), .ZN(n1221) );
XOR2_X1 U918 ( .A(G128), .B(G119), .Z(n1222) );
NAND2_X1 U919 ( .A1(KEYINPUT9), .A2(n1223), .ZN(n1219) );
XOR2_X1 U920 ( .A(n1180), .B(n1224), .Z(n1223) );
NAND2_X1 U921 ( .A1(n1225), .A2(G221), .ZN(n1224) );
INV_X1 U922 ( .A(G137), .ZN(n1180) );
XOR2_X1 U923 ( .A(n1226), .B(n1074), .Z(n1217) );
NAND2_X1 U924 ( .A1(KEYINPUT57), .A2(n1174), .ZN(n1226) );
INV_X1 U925 ( .A(n1193), .ZN(n1038) );
XOR2_X1 U926 ( .A(n1049), .B(G472), .Z(n1193) );
NAND2_X1 U927 ( .A1(n1227), .A2(n1228), .ZN(n1049) );
XOR2_X1 U928 ( .A(n1229), .B(n1230), .Z(n1228) );
XNOR2_X1 U929 ( .A(n1231), .B(n1115), .ZN(n1230) );
XNOR2_X1 U930 ( .A(n1232), .B(n1233), .ZN(n1115) );
NAND2_X1 U931 ( .A1(n1234), .A2(G210), .ZN(n1232) );
NAND2_X1 U932 ( .A1(KEYINPUT12), .A2(n1121), .ZN(n1231) );
AND3_X1 U933 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1121) );
INV_X1 U934 ( .A(n1238), .ZN(n1235) );
XOR2_X1 U935 ( .A(n1239), .B(G101), .Z(n1229) );
NAND2_X1 U936 ( .A1(KEYINPUT5), .A2(n1240), .ZN(n1239) );
XOR2_X1 U937 ( .A(n1241), .B(KEYINPUT25), .Z(n1227) );
NAND2_X1 U938 ( .A1(n1042), .A2(n1198), .ZN(n1015) );
XOR2_X1 U939 ( .A(n1058), .B(n1057), .Z(n1198) );
NOR2_X1 U940 ( .A1(n1107), .A2(G902), .ZN(n1057) );
NAND3_X1 U941 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1107) );
NAND2_X1 U942 ( .A1(KEYINPUT6), .A2(n1245), .ZN(n1244) );
OR3_X1 U943 ( .A1(n1246), .A2(KEYINPUT6), .A3(n1247), .ZN(n1243) );
NAND2_X1 U944 ( .A1(n1247), .A2(n1246), .ZN(n1242) );
NAND2_X1 U945 ( .A1(n1248), .A2(n1249), .ZN(n1246) );
INV_X1 U946 ( .A(n1245), .ZN(n1249) );
XOR2_X1 U947 ( .A(n1250), .B(n1251), .Z(n1245) );
XOR2_X1 U948 ( .A(n1252), .B(n1253), .Z(n1251) );
NAND2_X1 U949 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U950 ( .A1(n1256), .A2(n1174), .ZN(n1255) );
XOR2_X1 U951 ( .A(KEYINPUT20), .B(n1074), .Z(n1256) );
INV_X1 U952 ( .A(n1257), .ZN(n1074) );
NAND2_X1 U953 ( .A1(G146), .A2(n1258), .ZN(n1254) );
XOR2_X1 U954 ( .A(n1257), .B(KEYINPUT32), .Z(n1258) );
XOR2_X1 U955 ( .A(n1188), .B(G140), .Z(n1257) );
INV_X1 U956 ( .A(G125), .ZN(n1188) );
NAND2_X1 U957 ( .A1(n1234), .A2(G214), .ZN(n1252) );
NOR2_X1 U958 ( .A1(G953), .A2(G237), .ZN(n1234) );
XOR2_X1 U959 ( .A(G131), .B(n1176), .Z(n1250) );
XNOR2_X1 U960 ( .A(KEYINPUT50), .B(KEYINPUT31), .ZN(n1248) );
XNOR2_X1 U961 ( .A(n1259), .B(n1260), .ZN(n1247) );
XOR2_X1 U962 ( .A(G113), .B(G104), .Z(n1260) );
NAND2_X1 U963 ( .A1(KEYINPUT41), .A2(G122), .ZN(n1259) );
INV_X1 U964 ( .A(G475), .ZN(n1058) );
XOR2_X1 U965 ( .A(n1261), .B(G478), .Z(n1042) );
NAND2_X1 U966 ( .A1(n1100), .A2(n1241), .ZN(n1261) );
XNOR2_X1 U967 ( .A(n1262), .B(n1263), .ZN(n1100) );
XOR2_X1 U968 ( .A(n1264), .B(n1265), .Z(n1263) );
XNOR2_X1 U969 ( .A(n1266), .B(n1267), .ZN(n1265) );
NOR2_X1 U970 ( .A1(G143), .A2(KEYINPUT53), .ZN(n1267) );
NAND2_X1 U971 ( .A1(KEYINPUT17), .A2(n1268), .ZN(n1266) );
XOR2_X1 U972 ( .A(n1204), .B(n1269), .Z(n1268) );
NAND2_X1 U973 ( .A1(KEYINPUT1), .A2(n1194), .ZN(n1269) );
INV_X1 U974 ( .A(G122), .ZN(n1194) );
XOR2_X1 U975 ( .A(n1270), .B(n1271), .Z(n1262) );
XOR2_X1 U976 ( .A(G134), .B(G128), .Z(n1271) );
NAND3_X1 U977 ( .A1(KEYINPUT63), .A2(n1225), .A3(n1272), .ZN(n1270) );
XNOR2_X1 U978 ( .A(G217), .B(KEYINPUT35), .ZN(n1272) );
AND2_X1 U979 ( .A1(G234), .A2(n1084), .ZN(n1225) );
NAND3_X1 U980 ( .A1(n1206), .A2(n1205), .A3(n1183), .ZN(n1158) );
NOR2_X1 U981 ( .A1(n1017), .A2(n1026), .ZN(n1183) );
NOR2_X1 U982 ( .A1(n1273), .A2(n1045), .ZN(n1026) );
NOR2_X1 U983 ( .A1(n1053), .A2(G469), .ZN(n1045) );
AND2_X1 U984 ( .A1(G469), .A2(n1053), .ZN(n1273) );
NAND2_X1 U985 ( .A1(n1274), .A2(n1241), .ZN(n1053) );
XOR2_X1 U986 ( .A(n1128), .B(n1275), .Z(n1274) );
NOR2_X1 U987 ( .A1(KEYINPUT61), .A2(n1276), .ZN(n1275) );
XOR2_X1 U988 ( .A(n1131), .B(n1277), .Z(n1276) );
NOR2_X1 U989 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
AND3_X1 U990 ( .A1(KEYINPUT3), .A2(n1280), .A3(G140), .ZN(n1279) );
NOR2_X1 U991 ( .A1(KEYINPUT3), .A2(n1129), .ZN(n1278) );
XOR2_X1 U992 ( .A(G110), .B(G140), .Z(n1129) );
NAND2_X1 U993 ( .A1(G227), .A2(n1084), .ZN(n1131) );
XOR2_X1 U994 ( .A(n1281), .B(n1116), .Z(n1128) );
XOR2_X1 U995 ( .A(n1282), .B(n1240), .Z(n1116) );
XOR2_X1 U996 ( .A(n1283), .B(n1075), .Z(n1240) );
XOR2_X1 U997 ( .A(G131), .B(KEYINPUT24), .Z(n1075) );
NAND2_X1 U998 ( .A1(KEYINPUT59), .A2(n1077), .ZN(n1283) );
XNOR2_X1 U999 ( .A(G134), .B(n1284), .ZN(n1077) );
XOR2_X1 U1000 ( .A(KEYINPUT51), .B(G137), .Z(n1284) );
XOR2_X1 U1001 ( .A(n1285), .B(n1076), .Z(n1281) );
XOR2_X1 U1002 ( .A(G128), .B(n1286), .Z(n1076) );
XOR2_X1 U1003 ( .A(G146), .B(G143), .Z(n1286) );
NAND2_X1 U1004 ( .A1(KEYINPUT40), .A2(n1287), .ZN(n1285) );
INV_X1 U1005 ( .A(n1029), .ZN(n1017) );
NAND2_X1 U1006 ( .A1(G221), .A2(n1216), .ZN(n1029) );
NAND2_X1 U1007 ( .A1(G234), .A2(n1241), .ZN(n1216) );
NAND2_X1 U1008 ( .A1(n1288), .A2(n1289), .ZN(n1205) );
NAND4_X1 U1009 ( .A1(G953), .A2(G902), .A3(n1192), .A4(n1088), .ZN(n1289) );
INV_X1 U1010 ( .A(G898), .ZN(n1088) );
XOR2_X1 U1011 ( .A(n1010), .B(KEYINPUT18), .Z(n1288) );
NAND3_X1 U1012 ( .A1(n1192), .A2(n1084), .A3(G952), .ZN(n1010) );
NAND2_X1 U1013 ( .A1(G237), .A2(G234), .ZN(n1192) );
AND2_X1 U1014 ( .A1(n1024), .A2(n1025), .ZN(n1206) );
NAND2_X1 U1015 ( .A1(G214), .A2(n1290), .ZN(n1025) );
INV_X1 U1016 ( .A(n1185), .ZN(n1024) );
XNOR2_X1 U1017 ( .A(n1291), .B(n1135), .ZN(n1185) );
NAND2_X1 U1018 ( .A1(G210), .A2(n1290), .ZN(n1135) );
NAND2_X1 U1019 ( .A1(n1292), .A2(n1241), .ZN(n1290) );
INV_X1 U1020 ( .A(G237), .ZN(n1292) );
NAND4_X1 U1021 ( .A1(n1293), .A2(n1294), .A3(n1295), .A4(n1296), .ZN(n1291) );
OR3_X1 U1022 ( .A1(n1173), .A2(KEYINPUT34), .A3(n1297), .ZN(n1296) );
NAND2_X1 U1023 ( .A1(n1297), .A2(n1298), .ZN(n1295) );
NAND2_X1 U1024 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
INV_X1 U1025 ( .A(KEYINPUT34), .ZN(n1300) );
XOR2_X1 U1026 ( .A(n1173), .B(KEYINPUT8), .Z(n1299) );
XOR2_X1 U1027 ( .A(n1170), .B(G125), .Z(n1297) );
XNOR2_X1 U1028 ( .A(n1301), .B(n1233), .ZN(n1170) );
XNOR2_X1 U1029 ( .A(n1302), .B(n1303), .ZN(n1233) );
XOR2_X1 U1030 ( .A(n1174), .B(n1304), .Z(n1303) );
NAND2_X1 U1031 ( .A1(KEYINPUT55), .A2(n1176), .ZN(n1304) );
INV_X1 U1032 ( .A(G143), .ZN(n1176) );
INV_X1 U1033 ( .A(G146), .ZN(n1174) );
NAND2_X1 U1034 ( .A1(KEYINPUT29), .A2(G128), .ZN(n1302) );
NAND2_X1 U1035 ( .A1(G224), .A2(n1084), .ZN(n1301) );
INV_X1 U1036 ( .A(G953), .ZN(n1084) );
NAND2_X1 U1037 ( .A1(KEYINPUT34), .A2(n1173), .ZN(n1294) );
XOR2_X1 U1038 ( .A(n1305), .B(n1306), .Z(n1173) );
INV_X1 U1039 ( .A(n1089), .ZN(n1306) );
XOR2_X1 U1040 ( .A(n1307), .B(n1308), .Z(n1089) );
XOR2_X1 U1041 ( .A(n1280), .B(n1309), .Z(n1308) );
NAND4_X1 U1042 ( .A1(n1237), .A2(n1236), .A3(n1310), .A4(n1311), .ZN(n1309) );
NAND2_X1 U1043 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
INV_X1 U1044 ( .A(KEYINPUT0), .ZN(n1313) );
NAND2_X1 U1045 ( .A1(n1238), .A2(KEYINPUT0), .ZN(n1310) );
NOR2_X1 U1046 ( .A1(n1312), .A2(G119), .ZN(n1238) );
XOR2_X1 U1047 ( .A(n1210), .B(n1204), .Z(n1312) );
NAND3_X1 U1048 ( .A1(G116), .A2(n1210), .A3(G119), .ZN(n1236) );
INV_X1 U1049 ( .A(G113), .ZN(n1210) );
NAND3_X1 U1050 ( .A1(G119), .A2(n1204), .A3(G113), .ZN(n1237) );
INV_X1 U1051 ( .A(G116), .ZN(n1204) );
INV_X1 U1052 ( .A(G110), .ZN(n1280) );
NAND2_X1 U1053 ( .A1(KEYINPUT15), .A2(G122), .ZN(n1307) );
NAND2_X1 U1054 ( .A1(KEYINPUT27), .A2(n1314), .ZN(n1305) );
XOR2_X1 U1055 ( .A(KEYINPUT26), .B(n1090), .Z(n1314) );
XNOR2_X1 U1056 ( .A(n1287), .B(n1282), .ZN(n1090) );
INV_X1 U1057 ( .A(G101), .ZN(n1282) );
XOR2_X1 U1058 ( .A(G104), .B(n1264), .Z(n1287) );
XOR2_X1 U1059 ( .A(G107), .B(KEYINPUT54), .Z(n1264) );
XOR2_X1 U1060 ( .A(n1241), .B(KEYINPUT36), .Z(n1293) );
INV_X1 U1061 ( .A(G902), .ZN(n1241) );
endmodule


