//Key = 1001111000000111001100101111010001011100010101011011001000100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383;

XOR2_X1 U758 ( .A(n1045), .B(G107), .Z(G9) );
NAND2_X1 U759 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
OR3_X1 U760 ( .A1(n1048), .A2(n1049), .A3(KEYINPUT3), .ZN(n1047) );
NAND2_X1 U761 ( .A1(n1050), .A2(KEYINPUT3), .ZN(n1046) );
NOR2_X1 U762 ( .A1(n1051), .A2(n1052), .ZN(G75) );
NOR4_X1 U763 ( .A1(n1053), .A2(n1054), .A3(G953), .A4(n1055), .ZN(n1052) );
NOR3_X1 U764 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1054) );
NOR2_X1 U765 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U766 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
XNOR2_X1 U767 ( .A(n1063), .B(KEYINPUT0), .ZN(n1061) );
NAND4_X1 U768 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1053) );
NAND2_X1 U769 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND3_X1 U770 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
XOR2_X1 U771 ( .A(n1073), .B(KEYINPUT20), .Z(n1072) );
NAND2_X1 U772 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1071) );
NAND2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U776 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U777 ( .A1(KEYINPUT48), .A2(n1084), .ZN(n1078) );
NAND2_X1 U778 ( .A1(n1074), .A2(n1085), .ZN(n1070) );
INV_X1 U779 ( .A(n1056), .ZN(n1074) );
NAND3_X1 U780 ( .A1(n1086), .A2(n1080), .A3(n1087), .ZN(n1056) );
INV_X1 U781 ( .A(n1088), .ZN(n1087) );
INV_X1 U782 ( .A(n1089), .ZN(n1068) );
NAND4_X1 U783 ( .A1(n1084), .A2(n1090), .A3(n1076), .A4(n1089), .ZN(n1066) );
INV_X1 U784 ( .A(KEYINPUT48), .ZN(n1090) );
XOR2_X1 U785 ( .A(n1091), .B(KEYINPUT1), .Z(n1064) );
NAND4_X1 U786 ( .A1(n1092), .A2(n1076), .A3(n1093), .A4(n1086), .ZN(n1091) );
NOR2_X1 U787 ( .A1(n1089), .A2(n1094), .ZN(n1093) );
NOR2_X1 U788 ( .A1(n1088), .A2(n1058), .ZN(n1076) );
INV_X1 U789 ( .A(n1095), .ZN(n1058) );
NOR3_X1 U790 ( .A1(n1055), .A2(G953), .A3(G952), .ZN(n1051) );
AND4_X1 U791 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1055) );
NOR4_X1 U792 ( .A1(n1100), .A2(n1101), .A3(n1089), .A4(n1102), .ZN(n1099) );
XNOR2_X1 U793 ( .A(G469), .B(n1103), .ZN(n1102) );
AND2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(n1098) );
XNOR2_X1 U795 ( .A(n1106), .B(n1107), .ZN(n1097) );
NOR2_X1 U796 ( .A1(n1108), .A2(KEYINPUT23), .ZN(n1107) );
XOR2_X1 U797 ( .A(KEYINPUT24), .B(n1109), .Z(n1096) );
XOR2_X1 U798 ( .A(n1110), .B(n1111), .Z(G72) );
XOR2_X1 U799 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U800 ( .A1(n1114), .A2(G953), .ZN(n1113) );
NOR2_X1 U801 ( .A1(n1115), .A2(n1116), .ZN(n1112) );
XNOR2_X1 U802 ( .A(n1117), .B(n1118), .ZN(n1116) );
XOR2_X1 U803 ( .A(n1119), .B(n1120), .Z(n1118) );
NOR3_X1 U804 ( .A1(KEYINPUT60), .A2(n1121), .A3(n1122), .ZN(n1120) );
NOR3_X1 U805 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1122) );
NOR2_X1 U806 ( .A1(n1126), .A2(n1127), .ZN(n1121) );
INV_X1 U807 ( .A(n1123), .ZN(n1127) );
XOR2_X1 U808 ( .A(G131), .B(KEYINPUT28), .Z(n1123) );
NOR2_X1 U809 ( .A1(n1124), .A2(n1125), .ZN(n1126) );
NAND2_X1 U810 ( .A1(n1128), .A2(n1129), .ZN(n1125) );
OR2_X1 U811 ( .A1(G134), .A2(KEYINPUT43), .ZN(n1129) );
NAND3_X1 U812 ( .A1(G134), .A2(n1130), .A3(KEYINPUT43), .ZN(n1128) );
NOR2_X1 U813 ( .A1(G900), .A2(n1131), .ZN(n1115) );
NOR2_X1 U814 ( .A1(n1132), .A2(n1133), .ZN(n1110) );
NOR2_X1 U815 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
XOR2_X1 U816 ( .A(n1136), .B(n1137), .Z(G69) );
XOR2_X1 U817 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U818 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U819 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U820 ( .A(n1144), .B(KEYINPUT46), .Z(n1143) );
NAND2_X1 U821 ( .A1(n1145), .A2(n1146), .ZN(n1138) );
NAND2_X1 U822 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XNOR2_X1 U823 ( .A(n1050), .B(KEYINPUT32), .ZN(n1147) );
XNOR2_X1 U824 ( .A(G953), .B(KEYINPUT38), .ZN(n1145) );
NAND2_X1 U825 ( .A1(G953), .A2(n1149), .ZN(n1136) );
NAND2_X1 U826 ( .A1(G898), .A2(G224), .ZN(n1149) );
NOR2_X1 U827 ( .A1(n1150), .A2(n1151), .ZN(G66) );
XNOR2_X1 U828 ( .A(n1152), .B(n1153), .ZN(n1151) );
NOR2_X1 U829 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NOR2_X1 U830 ( .A1(n1150), .A2(n1156), .ZN(G63) );
XOR2_X1 U831 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U832 ( .A1(KEYINPUT30), .A2(n1159), .ZN(n1158) );
AND2_X1 U833 ( .A1(G478), .A2(n1160), .ZN(n1159) );
NOR2_X1 U834 ( .A1(n1150), .A2(n1161), .ZN(G60) );
NOR3_X1 U835 ( .A1(n1162), .A2(n1108), .A3(n1163), .ZN(n1161) );
NOR2_X1 U836 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NOR2_X1 U837 ( .A1(n1065), .A2(n1106), .ZN(n1165) );
XOR2_X1 U838 ( .A(n1166), .B(KEYINPUT14), .Z(n1162) );
NAND3_X1 U839 ( .A1(n1160), .A2(G475), .A3(n1164), .ZN(n1166) );
XOR2_X1 U840 ( .A(n1167), .B(n1168), .Z(G6) );
XOR2_X1 U841 ( .A(KEYINPUT63), .B(G104), .Z(n1168) );
NOR2_X1 U842 ( .A1(n1048), .A2(n1082), .ZN(n1167) );
NOR2_X1 U843 ( .A1(n1169), .A2(n1170), .ZN(G57) );
XOR2_X1 U844 ( .A(KEYINPUT7), .B(n1150), .Z(n1170) );
XOR2_X1 U845 ( .A(n1171), .B(n1172), .Z(n1169) );
XNOR2_X1 U846 ( .A(n1173), .B(n1174), .ZN(n1172) );
XOR2_X1 U847 ( .A(n1175), .B(n1176), .Z(n1171) );
XOR2_X1 U848 ( .A(n1177), .B(n1178), .Z(n1176) );
AND2_X1 U849 ( .A1(G472), .A2(n1160), .ZN(n1178) );
NAND2_X1 U850 ( .A1(KEYINPUT5), .A2(n1179), .ZN(n1175) );
NOR2_X1 U851 ( .A1(n1150), .A2(n1180), .ZN(G54) );
XOR2_X1 U852 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U853 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U854 ( .A1(KEYINPUT57), .A2(n1185), .ZN(n1184) );
NOR2_X1 U855 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
XOR2_X1 U856 ( .A(KEYINPUT56), .B(n1188), .Z(n1187) );
NOR2_X1 U857 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XNOR2_X1 U858 ( .A(KEYINPUT50), .B(G110), .ZN(n1189) );
NOR2_X1 U859 ( .A1(G140), .A2(n1191), .ZN(n1186) );
XNOR2_X1 U860 ( .A(KEYINPUT50), .B(n1192), .ZN(n1191) );
XOR2_X1 U861 ( .A(n1193), .B(n1194), .Z(n1181) );
NOR2_X1 U862 ( .A1(n1195), .A2(n1155), .ZN(n1194) );
NAND3_X1 U863 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1193) );
NAND2_X1 U864 ( .A1(KEYINPUT59), .A2(n1199), .ZN(n1198) );
NAND3_X1 U865 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1197) );
NAND2_X1 U866 ( .A1(n1203), .A2(n1204), .ZN(n1196) );
NAND2_X1 U867 ( .A1(n1205), .A2(n1201), .ZN(n1204) );
INV_X1 U868 ( .A(KEYINPUT59), .ZN(n1201) );
XNOR2_X1 U869 ( .A(n1200), .B(KEYINPUT13), .ZN(n1205) );
NOR3_X1 U870 ( .A1(n1150), .A2(n1206), .A3(n1207), .ZN(G51) );
NOR4_X1 U871 ( .A1(n1208), .A2(n1155), .A3(KEYINPUT17), .A4(n1209), .ZN(n1207) );
INV_X1 U872 ( .A(n1210), .ZN(n1208) );
NOR2_X1 U873 ( .A1(n1210), .A2(n1211), .ZN(n1206) );
NOR3_X1 U874 ( .A1(n1155), .A2(n1212), .A3(n1209), .ZN(n1211) );
AND2_X1 U875 ( .A1(n1213), .A2(KEYINPUT17), .ZN(n1212) );
INV_X1 U876 ( .A(n1160), .ZN(n1155) );
NOR2_X1 U877 ( .A1(n1214), .A2(n1065), .ZN(n1160) );
AND3_X1 U878 ( .A1(n1148), .A2(n1215), .A3(n1114), .ZN(n1065) );
AND2_X1 U879 ( .A1(n1216), .A2(n1217), .ZN(n1114) );
NOR4_X1 U880 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1217) );
NOR4_X1 U881 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1216) );
NOR2_X1 U882 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
NOR2_X1 U883 ( .A1(n1089), .A2(n1228), .ZN(n1224) );
INV_X1 U884 ( .A(n1050), .ZN(n1215) );
NOR2_X1 U885 ( .A1(n1083), .A2(n1048), .ZN(n1050) );
INV_X1 U886 ( .A(n1049), .ZN(n1083) );
AND4_X1 U887 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1148) );
NOR4_X1 U888 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1232) );
NOR3_X1 U889 ( .A1(n1082), .A2(KEYINPUT8), .A3(n1048), .ZN(n1235) );
NAND4_X1 U890 ( .A1(n1060), .A2(n1237), .A3(n1095), .A4(n1238), .ZN(n1048) );
NOR3_X1 U891 ( .A1(n1226), .A2(KEYINPUT11), .A3(n1239), .ZN(n1234) );
NOR2_X1 U892 ( .A1(n1060), .A2(n1240), .ZN(n1233) );
NOR2_X1 U893 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
NOR2_X1 U894 ( .A1(n1239), .A2(n1243), .ZN(n1242) );
INV_X1 U895 ( .A(KEYINPUT11), .ZN(n1243) );
NOR3_X1 U896 ( .A1(n1244), .A2(n1082), .A3(n1245), .ZN(n1241) );
INV_X1 U897 ( .A(KEYINPUT8), .ZN(n1245) );
INV_X1 U898 ( .A(n1246), .ZN(n1082) );
NAND3_X1 U899 ( .A1(n1095), .A2(n1238), .A3(n1237), .ZN(n1244) );
NOR2_X1 U900 ( .A1(n1247), .A2(n1248), .ZN(n1231) );
NOR2_X1 U901 ( .A1(KEYINPUT12), .A2(n1213), .ZN(n1210) );
XOR2_X1 U902 ( .A(n1249), .B(n1250), .Z(n1213) );
NAND4_X1 U903 ( .A1(KEYINPUT18), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1249) );
OR2_X1 U904 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND3_X1 U905 ( .A1(KEYINPUT25), .A2(n1255), .A3(n1254), .ZN(n1252) );
AND2_X1 U906 ( .A1(KEYINPUT15), .A2(n1256), .ZN(n1255) );
OR2_X1 U907 ( .A1(n1256), .A2(KEYINPUT25), .ZN(n1251) );
NOR2_X1 U908 ( .A1(n1133), .A2(G952), .ZN(n1150) );
XOR2_X1 U909 ( .A(G146), .B(n1223), .Z(G48) );
AND3_X1 U910 ( .A1(n1246), .A2(n1060), .A3(n1257), .ZN(n1223) );
XNOR2_X1 U911 ( .A(G143), .B(n1258), .ZN(G45) );
NAND2_X1 U912 ( .A1(n1259), .A2(n1060), .ZN(n1258) );
XOR2_X1 U913 ( .A(n1227), .B(KEYINPUT4), .Z(n1259) );
NAND3_X1 U914 ( .A1(n1260), .A2(n1085), .A3(n1261), .ZN(n1227) );
NOR3_X1 U915 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1261) );
XNOR2_X1 U916 ( .A(G140), .B(n1265), .ZN(G42) );
NAND2_X1 U917 ( .A1(KEYINPUT33), .A2(n1222), .ZN(n1265) );
AND3_X1 U918 ( .A1(n1246), .A2(n1075), .A3(n1266), .ZN(n1222) );
XNOR2_X1 U919 ( .A(n1130), .B(n1267), .ZN(G39) );
NOR2_X1 U920 ( .A1(n1089), .A2(n1268), .ZN(n1267) );
XNOR2_X1 U921 ( .A(KEYINPUT54), .B(n1228), .ZN(n1268) );
NAND2_X1 U922 ( .A1(n1086), .A2(n1257), .ZN(n1228) );
XNOR2_X1 U923 ( .A(n1221), .B(n1269), .ZN(G36) );
XNOR2_X1 U924 ( .A(G134), .B(KEYINPUT39), .ZN(n1269) );
AND3_X1 U925 ( .A1(n1085), .A2(n1049), .A3(n1266), .ZN(n1221) );
XNOR2_X1 U926 ( .A(n1270), .B(n1220), .ZN(G33) );
AND3_X1 U927 ( .A1(n1085), .A2(n1246), .A3(n1266), .ZN(n1220) );
NOR3_X1 U928 ( .A1(n1262), .A2(n1263), .A3(n1089), .ZN(n1266) );
NAND2_X1 U929 ( .A1(n1271), .A2(n1062), .ZN(n1089) );
INV_X1 U930 ( .A(n1063), .ZN(n1271) );
XOR2_X1 U931 ( .A(n1272), .B(n1219), .Z(G30) );
AND3_X1 U932 ( .A1(n1049), .A2(n1060), .A3(n1257), .ZN(n1219) );
AND4_X1 U933 ( .A1(n1237), .A2(n1100), .A3(n1273), .A4(n1274), .ZN(n1257) );
NAND2_X1 U934 ( .A1(KEYINPUT37), .A2(n1275), .ZN(n1272) );
XNOR2_X1 U935 ( .A(n1179), .B(n1276), .ZN(G3) );
NOR2_X1 U936 ( .A1(n1277), .A2(n1226), .ZN(n1276) );
XOR2_X1 U937 ( .A(n1239), .B(KEYINPUT31), .Z(n1277) );
NAND3_X1 U938 ( .A1(n1085), .A2(n1238), .A3(n1084), .ZN(n1239) );
XOR2_X1 U939 ( .A(G125), .B(n1218), .Z(G27) );
AND3_X1 U940 ( .A1(n1246), .A2(n1080), .A3(n1278), .ZN(n1218) );
NOR3_X1 U941 ( .A1(n1279), .A2(n1263), .A3(n1226), .ZN(n1278) );
INV_X1 U942 ( .A(n1273), .ZN(n1263) );
NAND2_X1 U943 ( .A1(n1088), .A2(n1280), .ZN(n1273) );
NAND4_X1 U944 ( .A1(G902), .A2(n1281), .A3(n1282), .A4(n1135), .ZN(n1280) );
INV_X1 U945 ( .A(G900), .ZN(n1135) );
XNOR2_X1 U946 ( .A(G122), .B(n1283), .ZN(G24) );
NAND2_X1 U947 ( .A1(KEYINPUT19), .A2(n1236), .ZN(n1283) );
AND4_X1 U948 ( .A1(n1260), .A2(n1284), .A3(n1095), .A4(n1101), .ZN(n1236) );
NOR2_X1 U949 ( .A1(n1274), .A2(n1100), .ZN(n1095) );
XOR2_X1 U950 ( .A(G119), .B(n1248), .Z(G21) );
AND4_X1 U951 ( .A1(n1284), .A2(n1086), .A3(n1100), .A4(n1274), .ZN(n1248) );
XOR2_X1 U952 ( .A(G116), .B(n1247), .Z(G18) );
AND3_X1 U953 ( .A1(n1085), .A2(n1049), .A3(n1284), .ZN(n1247) );
NOR2_X1 U954 ( .A1(n1260), .A2(n1264), .ZN(n1049) );
INV_X1 U955 ( .A(n1101), .ZN(n1264) );
XNOR2_X1 U956 ( .A(G113), .B(n1229), .ZN(G15) );
NAND3_X1 U957 ( .A1(n1085), .A2(n1246), .A3(n1284), .ZN(n1229) );
AND3_X1 U958 ( .A1(n1060), .A2(n1238), .A3(n1080), .ZN(n1284) );
NOR2_X1 U959 ( .A1(n1094), .A2(n1092), .ZN(n1080) );
INV_X1 U960 ( .A(n1105), .ZN(n1092) );
NOR2_X1 U961 ( .A1(n1285), .A2(n1101), .ZN(n1246) );
NOR2_X1 U962 ( .A1(n1274), .A2(n1286), .ZN(n1085) );
XNOR2_X1 U963 ( .A(G110), .B(n1230), .ZN(G12) );
NAND4_X1 U964 ( .A1(n1084), .A2(n1075), .A3(n1060), .A4(n1238), .ZN(n1230) );
NAND2_X1 U965 ( .A1(n1287), .A2(n1088), .ZN(n1238) );
NAND3_X1 U966 ( .A1(n1282), .A2(n1133), .A3(G952), .ZN(n1088) );
NAND3_X1 U967 ( .A1(n1140), .A2(n1282), .A3(G902), .ZN(n1287) );
NAND2_X1 U968 ( .A1(G237), .A2(G234), .ZN(n1282) );
NOR2_X1 U969 ( .A1(n1131), .A2(G898), .ZN(n1140) );
INV_X1 U970 ( .A(n1281), .ZN(n1131) );
XOR2_X1 U971 ( .A(G953), .B(KEYINPUT52), .Z(n1281) );
INV_X1 U972 ( .A(n1226), .ZN(n1060) );
NAND2_X1 U973 ( .A1(n1063), .A2(n1062), .ZN(n1226) );
NAND2_X1 U974 ( .A1(G214), .A2(n1288), .ZN(n1062) );
XOR2_X1 U975 ( .A(n1289), .B(n1209), .Z(n1063) );
NAND2_X1 U976 ( .A1(G210), .A2(n1288), .ZN(n1209) );
NAND2_X1 U977 ( .A1(n1290), .A2(n1214), .ZN(n1288) );
NAND2_X1 U978 ( .A1(n1291), .A2(n1214), .ZN(n1289) );
XNOR2_X1 U979 ( .A(n1250), .B(n1292), .ZN(n1291) );
XOR2_X1 U980 ( .A(n1293), .B(n1256), .Z(n1292) );
AND2_X1 U981 ( .A1(G224), .A2(n1133), .ZN(n1256) );
NAND2_X1 U982 ( .A1(KEYINPUT45), .A2(n1254), .ZN(n1293) );
XNOR2_X1 U983 ( .A(n1294), .B(G125), .ZN(n1254) );
XNOR2_X1 U984 ( .A(n1142), .B(n1295), .ZN(n1250) );
NOR2_X1 U985 ( .A1(KEYINPUT49), .A2(n1144), .ZN(n1295) );
XOR2_X1 U986 ( .A(n1296), .B(n1297), .Z(n1142) );
XNOR2_X1 U987 ( .A(n1298), .B(G110), .ZN(n1297) );
NAND2_X1 U988 ( .A1(n1299), .A2(n1300), .ZN(n1296) );
NAND3_X1 U989 ( .A1(G101), .A2(n1301), .A3(n1302), .ZN(n1300) );
INV_X1 U990 ( .A(KEYINPUT6), .ZN(n1302) );
NAND2_X1 U991 ( .A1(n1303), .A2(KEYINPUT6), .ZN(n1299) );
INV_X1 U992 ( .A(n1279), .ZN(n1075) );
NAND2_X1 U993 ( .A1(n1286), .A2(n1274), .ZN(n1279) );
NAND2_X1 U994 ( .A1(n1304), .A2(n1104), .ZN(n1274) );
NAND3_X1 U995 ( .A1(n1154), .A2(n1214), .A3(n1152), .ZN(n1104) );
XOR2_X1 U996 ( .A(KEYINPUT58), .B(n1109), .Z(n1304) );
NOR2_X1 U997 ( .A1(n1154), .A2(n1305), .ZN(n1109) );
AND2_X1 U998 ( .A1(n1152), .A2(n1214), .ZN(n1305) );
XNOR2_X1 U999 ( .A(n1306), .B(n1307), .ZN(n1152) );
XOR2_X1 U1000 ( .A(n1308), .B(n1309), .Z(n1307) );
XNOR2_X1 U1001 ( .A(n1310), .B(n1311), .ZN(n1309) );
NOR2_X1 U1002 ( .A1(KEYINPUT2), .A2(n1130), .ZN(n1311) );
NOR2_X1 U1003 ( .A1(KEYINPUT16), .A2(n1192), .ZN(n1310) );
INV_X1 U1004 ( .A(G110), .ZN(n1192) );
XNOR2_X1 U1005 ( .A(G119), .B(KEYINPUT55), .ZN(n1308) );
XNOR2_X1 U1006 ( .A(n1312), .B(n1313), .ZN(n1306) );
XOR2_X1 U1007 ( .A(n1314), .B(n1315), .Z(n1312) );
NAND2_X1 U1008 ( .A1(G221), .A2(n1316), .ZN(n1314) );
NAND2_X1 U1009 ( .A1(G217), .A2(n1317), .ZN(n1154) );
INV_X1 U1010 ( .A(n1100), .ZN(n1286) );
XNOR2_X1 U1011 ( .A(n1318), .B(G472), .ZN(n1100) );
NAND2_X1 U1012 ( .A1(n1319), .A2(n1214), .ZN(n1318) );
XOR2_X1 U1013 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1014 ( .A(n1177), .B(n1322), .Z(n1321) );
NOR2_X1 U1015 ( .A1(KEYINPUT40), .A2(n1173), .ZN(n1322) );
XOR2_X1 U1016 ( .A(n1294), .B(n1199), .Z(n1173) );
XNOR2_X1 U1017 ( .A(G128), .B(n1323), .ZN(n1294) );
NOR2_X1 U1018 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
NOR3_X1 U1019 ( .A1(KEYINPUT41), .A2(G146), .A3(n1326), .ZN(n1325) );
NOR2_X1 U1020 ( .A1(n1327), .A2(n1328), .ZN(n1324) );
INV_X1 U1021 ( .A(KEYINPUT41), .ZN(n1328) );
XNOR2_X1 U1022 ( .A(G146), .B(n1326), .ZN(n1327) );
AND3_X1 U1023 ( .A1(n1290), .A2(n1133), .A3(G210), .ZN(n1177) );
INV_X1 U1024 ( .A(G237), .ZN(n1290) );
XNOR2_X1 U1025 ( .A(n1329), .B(n1174), .ZN(n1320) );
XOR2_X1 U1026 ( .A(n1144), .B(KEYINPUT53), .Z(n1174) );
XOR2_X1 U1027 ( .A(n1330), .B(n1331), .Z(n1144) );
XOR2_X1 U1028 ( .A(KEYINPUT47), .B(G119), .Z(n1331) );
XNOR2_X1 U1029 ( .A(G116), .B(G113), .ZN(n1330) );
NAND2_X1 U1030 ( .A1(KEYINPUT51), .A2(n1179), .ZN(n1329) );
INV_X1 U1031 ( .A(G101), .ZN(n1179) );
AND2_X1 U1032 ( .A1(n1086), .A2(n1237), .ZN(n1084) );
INV_X1 U1033 ( .A(n1262), .ZN(n1237) );
NAND2_X1 U1034 ( .A1(n1105), .A2(n1094), .ZN(n1262) );
NAND3_X1 U1035 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1094) );
NAND2_X1 U1036 ( .A1(G469), .A2(n1103), .ZN(n1334) );
NAND2_X1 U1037 ( .A1(KEYINPUT42), .A2(n1335), .ZN(n1333) );
NAND2_X1 U1038 ( .A1(n1336), .A2(n1195), .ZN(n1335) );
INV_X1 U1039 ( .A(G469), .ZN(n1195) );
XNOR2_X1 U1040 ( .A(KEYINPUT9), .B(n1103), .ZN(n1336) );
NAND2_X1 U1041 ( .A1(n1337), .A2(n1338), .ZN(n1332) );
INV_X1 U1042 ( .A(KEYINPUT42), .ZN(n1338) );
NAND2_X1 U1043 ( .A1(n1339), .A2(n1340), .ZN(n1337) );
NAND2_X1 U1044 ( .A1(KEYINPUT9), .A2(n1103), .ZN(n1340) );
OR3_X1 U1045 ( .A1(G469), .A2(KEYINPUT9), .A3(n1103), .ZN(n1339) );
NAND2_X1 U1046 ( .A1(n1341), .A2(n1214), .ZN(n1103) );
XOR2_X1 U1047 ( .A(n1342), .B(n1343), .Z(n1341) );
XNOR2_X1 U1048 ( .A(n1202), .B(n1200), .ZN(n1343) );
INV_X1 U1049 ( .A(n1199), .ZN(n1200) );
NAND3_X1 U1050 ( .A1(n1344), .A2(n1345), .A3(n1346), .ZN(n1199) );
NAND2_X1 U1051 ( .A1(n1124), .A2(G131), .ZN(n1346) );
NOR2_X1 U1052 ( .A1(n1130), .A2(G134), .ZN(n1124) );
NAND3_X1 U1053 ( .A1(G134), .A2(n1270), .A3(G137), .ZN(n1345) );
INV_X1 U1054 ( .A(G131), .ZN(n1270) );
NAND2_X1 U1055 ( .A1(n1347), .A2(n1130), .ZN(n1344) );
INV_X1 U1056 ( .A(G137), .ZN(n1130) );
XNOR2_X1 U1057 ( .A(G131), .B(G134), .ZN(n1347) );
INV_X1 U1058 ( .A(n1203), .ZN(n1202) );
XOR2_X1 U1059 ( .A(n1303), .B(n1348), .Z(n1203) );
INV_X1 U1060 ( .A(n1117), .ZN(n1348) );
XOR2_X1 U1061 ( .A(G143), .B(n1315), .Z(n1117) );
XNOR2_X1 U1062 ( .A(n1275), .B(G146), .ZN(n1315) );
INV_X1 U1063 ( .A(G128), .ZN(n1275) );
XOR2_X1 U1064 ( .A(G101), .B(n1301), .Z(n1303) );
XOR2_X1 U1065 ( .A(G104), .B(G107), .Z(n1301) );
XNOR2_X1 U1066 ( .A(n1183), .B(n1349), .ZN(n1342) );
XNOR2_X1 U1067 ( .A(n1190), .B(G110), .ZN(n1349) );
INV_X1 U1068 ( .A(G140), .ZN(n1190) );
NOR2_X1 U1069 ( .A1(n1134), .A2(G953), .ZN(n1183) );
INV_X1 U1070 ( .A(G227), .ZN(n1134) );
NAND2_X1 U1071 ( .A1(G221), .A2(n1317), .ZN(n1105) );
NAND2_X1 U1072 ( .A1(G234), .A2(n1214), .ZN(n1317) );
NOR2_X1 U1073 ( .A1(n1101), .A2(n1260), .ZN(n1086) );
INV_X1 U1074 ( .A(n1285), .ZN(n1260) );
XOR2_X1 U1075 ( .A(n1108), .B(n1350), .Z(n1285) );
XNOR2_X1 U1076 ( .A(KEYINPUT35), .B(n1106), .ZN(n1350) );
INV_X1 U1077 ( .A(G475), .ZN(n1106) );
NOR2_X1 U1078 ( .A1(n1164), .A2(G902), .ZN(n1108) );
AND2_X1 U1079 ( .A1(n1351), .A2(n1352), .ZN(n1164) );
NAND2_X1 U1080 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
XOR2_X1 U1081 ( .A(KEYINPUT29), .B(n1355), .Z(n1351) );
NOR2_X1 U1082 ( .A1(n1353), .A2(n1354), .ZN(n1355) );
XOR2_X1 U1083 ( .A(n1356), .B(n1357), .Z(n1354) );
XOR2_X1 U1084 ( .A(KEYINPUT62), .B(G104), .Z(n1357) );
NAND2_X1 U1085 ( .A1(n1358), .A2(n1359), .ZN(n1356) );
NAND2_X1 U1086 ( .A1(G113), .A2(n1298), .ZN(n1359) );
XOR2_X1 U1087 ( .A(KEYINPUT26), .B(n1360), .Z(n1358) );
NOR2_X1 U1088 ( .A1(G113), .A2(n1298), .ZN(n1360) );
XOR2_X1 U1089 ( .A(n1361), .B(n1362), .Z(n1353) );
XOR2_X1 U1090 ( .A(KEYINPUT55), .B(G146), .Z(n1362) );
XNOR2_X1 U1091 ( .A(n1363), .B(n1364), .ZN(n1361) );
NOR2_X1 U1092 ( .A1(KEYINPUT21), .A2(n1313), .ZN(n1364) );
XOR2_X1 U1093 ( .A(n1119), .B(KEYINPUT34), .Z(n1313) );
XNOR2_X1 U1094 ( .A(G125), .B(G140), .ZN(n1119) );
NOR2_X1 U1095 ( .A1(KEYINPUT61), .A2(n1365), .ZN(n1363) );
XOR2_X1 U1096 ( .A(n1366), .B(n1367), .Z(n1365) );
XOR2_X1 U1097 ( .A(n1368), .B(n1369), .Z(n1367) );
NAND2_X1 U1098 ( .A1(KEYINPUT22), .A2(G131), .ZN(n1369) );
NAND3_X1 U1099 ( .A1(G214), .A2(n1133), .A3(n1370), .ZN(n1368) );
XNOR2_X1 U1100 ( .A(G237), .B(KEYINPUT10), .ZN(n1370) );
XNOR2_X1 U1101 ( .A(G143), .B(KEYINPUT44), .ZN(n1366) );
XNOR2_X1 U1102 ( .A(n1371), .B(G478), .ZN(n1101) );
NAND2_X1 U1103 ( .A1(n1214), .A2(n1157), .ZN(n1371) );
NAND2_X1 U1104 ( .A1(n1372), .A2(n1373), .ZN(n1157) );
NAND4_X1 U1105 ( .A1(n1374), .A2(n1316), .A3(n1375), .A4(n1376), .ZN(n1373) );
NAND2_X1 U1106 ( .A1(n1377), .A2(n1378), .ZN(n1372) );
NAND2_X1 U1107 ( .A1(n1375), .A2(n1376), .ZN(n1378) );
NAND2_X1 U1108 ( .A1(n1379), .A2(n1380), .ZN(n1376) );
XNOR2_X1 U1109 ( .A(n1381), .B(KEYINPUT27), .ZN(n1375) );
OR2_X1 U1110 ( .A1(n1380), .A2(n1379), .ZN(n1381) );
XNOR2_X1 U1111 ( .A(G107), .B(n1382), .ZN(n1379) );
XNOR2_X1 U1112 ( .A(n1298), .B(G116), .ZN(n1382) );
INV_X1 U1113 ( .A(G122), .ZN(n1298) );
XOR2_X1 U1114 ( .A(G128), .B(n1383), .Z(n1380) );
XNOR2_X1 U1115 ( .A(n1326), .B(G134), .ZN(n1383) );
INV_X1 U1116 ( .A(G143), .ZN(n1326) );
NAND2_X1 U1117 ( .A1(n1316), .A2(n1374), .ZN(n1377) );
XNOR2_X1 U1118 ( .A(G217), .B(KEYINPUT36), .ZN(n1374) );
AND2_X1 U1119 ( .A1(G234), .A2(n1133), .ZN(n1316) );
INV_X1 U1120 ( .A(G953), .ZN(n1133) );
INV_X1 U1121 ( .A(G902), .ZN(n1214) );
endmodule


