//Key = 1110010111001011100100001001100111011111101000001001111010001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328;

XOR2_X1 U729 ( .A(G107), .B(n1005), .Z(G9) );
NOR3_X1 U730 ( .A1(n1006), .A2(KEYINPUT59), .A3(n1007), .ZN(n1005) );
NOR2_X1 U731 ( .A1(n1008), .A2(n1009), .ZN(G75) );
XOR2_X1 U732 ( .A(n1010), .B(KEYINPUT12), .Z(n1009) );
NAND3_X1 U733 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1010) );
NOR3_X1 U734 ( .A1(n1014), .A2(n1011), .A3(n1015), .ZN(n1008) );
INV_X1 U735 ( .A(G952), .ZN(n1011) );
NAND3_X1 U736 ( .A1(n1013), .A2(n1012), .A3(n1016), .ZN(n1014) );
NAND2_X1 U737 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND2_X1 U738 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND4_X1 U739 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1020) );
NAND2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U741 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND3_X1 U742 ( .A1(n1027), .A2(n1029), .A3(n1030), .ZN(n1019) );
NAND2_X1 U743 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NAND3_X1 U744 ( .A1(n1022), .A2(n1033), .A3(n1021), .ZN(n1032) );
NAND2_X1 U745 ( .A1(n1034), .A2(n1006), .ZN(n1033) );
NAND2_X1 U746 ( .A1(n1023), .A2(n1035), .ZN(n1031) );
NAND2_X1 U747 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U748 ( .A1(n1021), .A2(n1038), .ZN(n1037) );
NAND2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U750 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U751 ( .A1(n1022), .A2(n1043), .ZN(n1036) );
NAND2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U753 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
INV_X1 U754 ( .A(n1048), .ZN(n1017) );
NAND4_X1 U755 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1013) );
NOR3_X1 U756 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
XOR2_X1 U757 ( .A(n1042), .B(KEYINPUT2), .Z(n1055) );
XOR2_X1 U758 ( .A(n1056), .B(n1057), .Z(n1054) );
NAND2_X1 U759 ( .A1(n1058), .A2(KEYINPUT61), .ZN(n1056) );
XNOR2_X1 U760 ( .A(G478), .B(KEYINPUT23), .ZN(n1058) );
NAND3_X1 U761 ( .A1(n1059), .A2(n1060), .A3(n1030), .ZN(n1053) );
OR2_X1 U762 ( .A1(G475), .A2(KEYINPUT8), .ZN(n1060) );
NAND3_X1 U763 ( .A1(G475), .A2(n1061), .A3(KEYINPUT8), .ZN(n1059) );
NOR3_X1 U764 ( .A1(n1046), .A2(n1062), .A3(n1041), .ZN(n1051) );
XOR2_X1 U765 ( .A(n1063), .B(n1064), .Z(n1050) );
NOR2_X1 U766 ( .A1(n1065), .A2(KEYINPUT11), .ZN(n1064) );
INV_X1 U767 ( .A(n1066), .ZN(n1065) );
XOR2_X1 U768 ( .A(G472), .B(n1067), .Z(n1049) );
NOR2_X1 U769 ( .A1(n1068), .A2(KEYINPUT34), .ZN(n1067) );
XOR2_X1 U770 ( .A(n1069), .B(n1070), .Z(G72) );
NOR2_X1 U771 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U772 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XNOR2_X1 U773 ( .A(KEYINPUT17), .B(n1075), .ZN(n1074) );
NOR2_X1 U774 ( .A1(n1076), .A2(n1075), .ZN(n1071) );
NAND2_X1 U775 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NAND2_X1 U776 ( .A1(G953), .A2(n1079), .ZN(n1078) );
XOR2_X1 U777 ( .A(n1080), .B(n1081), .Z(n1077) );
XOR2_X1 U778 ( .A(G125), .B(n1082), .Z(n1081) );
NOR2_X1 U779 ( .A1(KEYINPUT44), .A2(n1083), .ZN(n1082) );
XOR2_X1 U780 ( .A(n1084), .B(n1085), .Z(n1083) );
NAND3_X1 U781 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1084) );
NAND2_X1 U782 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
OR3_X1 U783 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1087) );
INV_X1 U784 ( .A(KEYINPUT5), .ZN(n1090) );
NAND2_X1 U785 ( .A1(n1092), .A2(n1091), .ZN(n1086) );
NAND2_X1 U786 ( .A1(KEYINPUT16), .A2(G131), .ZN(n1091) );
XNOR2_X1 U787 ( .A(n1093), .B(KEYINPUT63), .ZN(n1092) );
XOR2_X1 U788 ( .A(KEYINPUT58), .B(G140), .Z(n1080) );
XOR2_X1 U789 ( .A(n1073), .B(KEYINPUT35), .Z(n1076) );
NAND2_X1 U790 ( .A1(n1012), .A2(n1094), .ZN(n1073) );
NAND3_X1 U791 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1094) );
INV_X1 U792 ( .A(n1098), .ZN(n1097) );
XOR2_X1 U793 ( .A(KEYINPUT42), .B(n1099), .Z(n1095) );
NAND2_X1 U794 ( .A1(G953), .A2(n1100), .ZN(n1069) );
NAND2_X1 U795 ( .A1(G900), .A2(G227), .ZN(n1100) );
NAND2_X1 U796 ( .A1(n1101), .A2(n1102), .ZN(G69) );
NAND2_X1 U797 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
INV_X1 U798 ( .A(n1105), .ZN(n1103) );
NAND2_X1 U799 ( .A1(n1105), .A2(n1106), .ZN(n1101) );
NAND2_X1 U800 ( .A1(n1107), .A2(n1104), .ZN(n1106) );
NAND2_X1 U801 ( .A1(G953), .A2(n1108), .ZN(n1104) );
INV_X1 U802 ( .A(G224), .ZN(n1108) );
INV_X1 U803 ( .A(n1109), .ZN(n1107) );
XOR2_X1 U804 ( .A(n1110), .B(n1111), .Z(n1105) );
NOR2_X1 U805 ( .A1(n1109), .A2(n1112), .ZN(n1111) );
XOR2_X1 U806 ( .A(KEYINPUT54), .B(n1113), .Z(n1112) );
NOR2_X1 U807 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U808 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XNOR2_X1 U809 ( .A(n1118), .B(KEYINPUT47), .ZN(n1117) );
NOR2_X1 U810 ( .A1(n1119), .A2(n1118), .ZN(n1114) );
XOR2_X1 U811 ( .A(n1120), .B(n1121), .Z(n1118) );
NAND2_X1 U812 ( .A1(KEYINPUT14), .A2(n1122), .ZN(n1120) );
NAND2_X1 U813 ( .A1(n1123), .A2(n1012), .ZN(n1110) );
NAND2_X1 U814 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U815 ( .A(n1126), .B(KEYINPUT30), .Z(n1124) );
NOR2_X1 U816 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XNOR2_X1 U817 ( .A(n1129), .B(n1130), .ZN(n1128) );
NOR2_X1 U818 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U819 ( .A(KEYINPUT33), .B(G217), .Z(n1132) );
NOR2_X1 U820 ( .A1(n1127), .A2(n1133), .ZN(G63) );
NOR3_X1 U821 ( .A1(n1057), .A2(n1134), .A3(n1135), .ZN(n1133) );
AND3_X1 U822 ( .A1(n1136), .A2(G478), .A3(n1137), .ZN(n1135) );
NOR2_X1 U823 ( .A1(n1138), .A2(n1136), .ZN(n1134) );
AND2_X1 U824 ( .A1(n1015), .A2(G478), .ZN(n1138) );
NOR2_X1 U825 ( .A1(n1127), .A2(n1139), .ZN(G60) );
XOR2_X1 U826 ( .A(n1140), .B(n1141), .Z(n1139) );
AND2_X1 U827 ( .A1(G475), .A2(n1137), .ZN(n1140) );
XOR2_X1 U828 ( .A(n1142), .B(n1143), .Z(G6) );
XOR2_X1 U829 ( .A(KEYINPUT28), .B(G104), .Z(n1143) );
NOR2_X1 U830 ( .A1(n1127), .A2(n1144), .ZN(G57) );
XOR2_X1 U831 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U832 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U833 ( .A(n1149), .B(n1150), .Z(n1145) );
AND2_X1 U834 ( .A1(G472), .A2(n1137), .ZN(n1150) );
NOR2_X1 U835 ( .A1(KEYINPUT18), .A2(n1151), .ZN(n1149) );
XOR2_X1 U836 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U837 ( .A1(n1127), .A2(n1154), .ZN(G54) );
XNOR2_X1 U838 ( .A(n1155), .B(n1156), .ZN(n1154) );
XOR2_X1 U839 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND3_X1 U840 ( .A1(n1137), .A2(G469), .A3(KEYINPUT56), .ZN(n1158) );
INV_X1 U841 ( .A(n1131), .ZN(n1137) );
NAND2_X1 U842 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NAND2_X1 U843 ( .A1(n1161), .A2(n1152), .ZN(n1160) );
XOR2_X1 U844 ( .A(KEYINPUT15), .B(n1162), .Z(n1159) );
NOR2_X1 U845 ( .A1(n1152), .A2(n1163), .ZN(n1162) );
XOR2_X1 U846 ( .A(KEYINPUT50), .B(n1161), .Z(n1163) );
XOR2_X1 U847 ( .A(n1164), .B(n1165), .Z(n1161) );
XOR2_X1 U848 ( .A(n1153), .B(KEYINPUT48), .Z(n1164) );
NOR2_X1 U849 ( .A1(n1127), .A2(n1166), .ZN(G51) );
NOR2_X1 U850 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U851 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U852 ( .A1(n1066), .A2(n1131), .ZN(n1170) );
NAND2_X1 U853 ( .A1(G902), .A2(n1015), .ZN(n1131) );
NAND3_X1 U854 ( .A1(n1171), .A2(n1125), .A3(n1172), .ZN(n1015) );
NOR3_X1 U855 ( .A1(n1098), .A2(n1173), .A3(n1099), .ZN(n1172) );
NAND4_X1 U856 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1098) );
NOR3_X1 U857 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1177) );
AND4_X1 U858 ( .A1(n1181), .A2(n1182), .A3(n1021), .A4(n1183), .ZN(n1180) );
AND3_X1 U859 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1178) );
AND4_X1 U860 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1125) );
AND4_X1 U861 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1142), .ZN(n1190) );
OR2_X1 U862 ( .A1(n1034), .A2(n1007), .ZN(n1142) );
OR2_X1 U863 ( .A1(n1006), .A2(n1007), .ZN(n1189) );
NAND2_X1 U864 ( .A1(n1194), .A2(n1030), .ZN(n1007) );
XOR2_X1 U865 ( .A(n1096), .B(KEYINPUT13), .Z(n1171) );
AND2_X1 U866 ( .A1(n1195), .A2(KEYINPUT36), .ZN(n1169) );
NOR2_X1 U867 ( .A1(KEYINPUT36), .A2(n1195), .ZN(n1167) );
XNOR2_X1 U868 ( .A(n1196), .B(n1197), .ZN(n1195) );
NOR2_X1 U869 ( .A1(KEYINPUT10), .A2(n1198), .ZN(n1197) );
XOR2_X1 U870 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U871 ( .A1(KEYINPUT49), .A2(n1201), .ZN(n1200) );
AND2_X1 U872 ( .A1(G953), .A2(n1202), .ZN(n1127) );
XOR2_X1 U873 ( .A(KEYINPUT40), .B(G952), .Z(n1202) );
XOR2_X1 U874 ( .A(n1203), .B(n1204), .Z(G48) );
NAND4_X1 U875 ( .A1(KEYINPUT19), .A2(n1184), .A3(n1186), .A4(n1185), .ZN(n1204) );
XOR2_X1 U876 ( .A(n1205), .B(G143), .Z(G45) );
NAND2_X1 U877 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND4_X1 U878 ( .A1(n1039), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1207) );
INV_X1 U879 ( .A(KEYINPUT32), .ZN(n1210) );
NAND2_X1 U880 ( .A1(n1099), .A2(KEYINPUT32), .ZN(n1206) );
AND3_X1 U881 ( .A1(n1182), .A2(n1208), .A3(n1209), .ZN(n1099) );
NOR4_X1 U882 ( .A1(n1025), .A2(n1044), .A3(n1211), .A4(n1212), .ZN(n1209) );
INV_X1 U883 ( .A(n1185), .ZN(n1044) );
XNOR2_X1 U884 ( .A(G140), .B(n1213), .ZN(G42) );
NAND4_X1 U885 ( .A1(n1214), .A2(n1183), .A3(n1021), .A4(n1182), .ZN(n1213) );
XOR2_X1 U886 ( .A(n1181), .B(KEYINPUT43), .Z(n1214) );
XNOR2_X1 U887 ( .A(G137), .B(n1175), .ZN(G39) );
NAND3_X1 U888 ( .A1(n1184), .A2(n1023), .A3(n1021), .ZN(n1175) );
INV_X1 U889 ( .A(n1215), .ZN(n1021) );
XNOR2_X1 U890 ( .A(G134), .B(n1096), .ZN(G36) );
NAND2_X1 U891 ( .A1(n1216), .A2(n1217), .ZN(n1096) );
XOR2_X1 U892 ( .A(G131), .B(n1179), .Z(G33) );
AND2_X1 U893 ( .A1(n1216), .A2(n1186), .ZN(n1179) );
NOR4_X1 U894 ( .A1(n1215), .A2(n1025), .A3(n1039), .A4(n1212), .ZN(n1216) );
NAND2_X1 U895 ( .A1(n1047), .A2(n1218), .ZN(n1215) );
XOR2_X1 U896 ( .A(n1219), .B(n1176), .Z(G30) );
NAND3_X1 U897 ( .A1(n1217), .A2(n1185), .A3(n1184), .ZN(n1176) );
NOR4_X1 U898 ( .A1(n1039), .A2(n1030), .A3(n1027), .A4(n1212), .ZN(n1184) );
INV_X1 U899 ( .A(n1181), .ZN(n1212) );
XOR2_X1 U900 ( .A(n1220), .B(n1173), .Z(G3) );
INV_X1 U901 ( .A(n1126), .ZN(n1173) );
NAND3_X1 U902 ( .A1(n1023), .A2(n1182), .A3(n1221), .ZN(n1126) );
NAND2_X1 U903 ( .A1(KEYINPUT9), .A2(n1222), .ZN(n1220) );
XOR2_X1 U904 ( .A(n1223), .B(n1174), .Z(G27) );
NAND4_X1 U905 ( .A1(n1183), .A2(n1022), .A3(n1185), .A4(n1181), .ZN(n1174) );
NAND2_X1 U906 ( .A1(n1048), .A2(n1224), .ZN(n1181) );
NAND4_X1 U907 ( .A1(G902), .A2(G953), .A3(n1225), .A4(n1079), .ZN(n1224) );
INV_X1 U908 ( .A(G900), .ZN(n1079) );
NOR3_X1 U909 ( .A1(n1226), .A2(n1030), .A3(n1034), .ZN(n1183) );
XNOR2_X1 U910 ( .A(G122), .B(n1187), .ZN(G24) );
NAND4_X1 U911 ( .A1(n1030), .A2(n1227), .A3(n1022), .A4(n1228), .ZN(n1187) );
NOR3_X1 U912 ( .A1(n1226), .A2(n1229), .A3(n1211), .ZN(n1228) );
XOR2_X1 U913 ( .A(n1230), .B(n1188), .Z(G21) );
NAND4_X1 U914 ( .A1(n1022), .A2(n1023), .A3(n1231), .A4(n1227), .ZN(n1188) );
INV_X1 U915 ( .A(n1232), .ZN(n1227) );
NOR2_X1 U916 ( .A1(n1027), .A2(n1030), .ZN(n1231) );
INV_X1 U917 ( .A(n1226), .ZN(n1027) );
XNOR2_X1 U918 ( .A(G116), .B(n1193), .ZN(G18) );
NAND3_X1 U919 ( .A1(n1221), .A2(n1217), .A3(n1022), .ZN(n1193) );
INV_X1 U920 ( .A(n1006), .ZN(n1217) );
NAND2_X1 U921 ( .A1(n1229), .A2(n1233), .ZN(n1006) );
XNOR2_X1 U922 ( .A(KEYINPUT26), .B(n1211), .ZN(n1233) );
XOR2_X1 U923 ( .A(n1234), .B(n1192), .Z(G15) );
NAND3_X1 U924 ( .A1(n1186), .A2(n1221), .A3(n1022), .ZN(n1192) );
NOR2_X1 U925 ( .A1(n1235), .A2(n1041), .ZN(n1022) );
INV_X1 U926 ( .A(n1042), .ZN(n1235) );
NOR2_X1 U927 ( .A1(n1025), .A2(n1232), .ZN(n1221) );
NAND2_X1 U928 ( .A1(n1030), .A2(n1226), .ZN(n1025) );
INV_X1 U929 ( .A(n1034), .ZN(n1186) );
NAND2_X1 U930 ( .A1(n1236), .A2(n1208), .ZN(n1034) );
INV_X1 U931 ( .A(n1229), .ZN(n1208) );
XNOR2_X1 U932 ( .A(G110), .B(n1191), .ZN(G12) );
NAND3_X1 U933 ( .A1(n1194), .A2(n1028), .A3(n1023), .ZN(n1191) );
AND2_X1 U934 ( .A1(n1236), .A2(n1229), .ZN(n1023) );
NOR2_X1 U935 ( .A1(n1237), .A2(n1062), .ZN(n1229) );
NOR2_X1 U936 ( .A1(n1061), .A2(G475), .ZN(n1062) );
AND2_X1 U937 ( .A1(G475), .A2(n1061), .ZN(n1237) );
OR2_X1 U938 ( .A1(n1141), .A2(G902), .ZN(n1061) );
XNOR2_X1 U939 ( .A(n1203), .B(n1238), .ZN(n1141) );
XOR2_X1 U940 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U941 ( .A(n1241), .B(n1242), .Z(n1240) );
XOR2_X1 U942 ( .A(G104), .B(n1243), .Z(n1242) );
AND3_X1 U943 ( .A1(G214), .A2(n1012), .A3(n1244), .ZN(n1243) );
XOR2_X1 U944 ( .A(n1245), .B(n1246), .Z(n1241) );
NOR2_X1 U945 ( .A1(G125), .A2(KEYINPUT3), .ZN(n1246) );
NAND2_X1 U946 ( .A1(KEYINPUT7), .A2(G143), .ZN(n1245) );
XOR2_X1 U947 ( .A(n1247), .B(n1248), .Z(n1239) );
XOR2_X1 U948 ( .A(G140), .B(G131), .Z(n1248) );
XOR2_X1 U949 ( .A(n1234), .B(G122), .Z(n1247) );
INV_X1 U950 ( .A(G113), .ZN(n1234) );
INV_X1 U951 ( .A(G146), .ZN(n1203) );
XOR2_X1 U952 ( .A(n1211), .B(KEYINPUT6), .Z(n1236) );
XNOR2_X1 U953 ( .A(n1057), .B(G478), .ZN(n1211) );
NOR2_X1 U954 ( .A1(n1136), .A2(G902), .ZN(n1057) );
XNOR2_X1 U955 ( .A(n1249), .B(n1250), .ZN(n1136) );
XOR2_X1 U956 ( .A(n1251), .B(n1252), .Z(n1250) );
XOR2_X1 U957 ( .A(G122), .B(G116), .Z(n1252) );
XOR2_X1 U958 ( .A(G134), .B(G128), .Z(n1251) );
XOR2_X1 U959 ( .A(n1253), .B(n1254), .Z(n1249) );
AND3_X1 U960 ( .A1(G234), .A2(n1012), .A3(G217), .ZN(n1254) );
XOR2_X1 U961 ( .A(n1255), .B(G107), .Z(n1253) );
NAND2_X1 U962 ( .A1(KEYINPUT51), .A2(n1256), .ZN(n1255) );
INV_X1 U963 ( .A(G143), .ZN(n1256) );
INV_X1 U964 ( .A(n1030), .ZN(n1028) );
XOR2_X1 U965 ( .A(n1257), .B(n1258), .Z(n1030) );
NOR2_X1 U966 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
INV_X1 U967 ( .A(G217), .ZN(n1260) );
XOR2_X1 U968 ( .A(n1261), .B(KEYINPUT0), .Z(n1259) );
NAND2_X1 U969 ( .A1(n1129), .A2(n1262), .ZN(n1257) );
XNOR2_X1 U970 ( .A(n1263), .B(n1264), .ZN(n1129) );
XOR2_X1 U971 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U972 ( .A(G128), .B(G125), .Z(n1266) );
XOR2_X1 U973 ( .A(G146), .B(G137), .Z(n1265) );
XOR2_X1 U974 ( .A(n1267), .B(n1268), .Z(n1263) );
XOR2_X1 U975 ( .A(n1269), .B(G119), .Z(n1267) );
NAND3_X1 U976 ( .A1(n1270), .A2(n1012), .A3(G221), .ZN(n1269) );
XOR2_X1 U977 ( .A(KEYINPUT20), .B(G234), .Z(n1270) );
NOR3_X1 U978 ( .A1(n1226), .A2(n1039), .A3(n1232), .ZN(n1194) );
NAND2_X1 U979 ( .A1(n1185), .A2(n1271), .ZN(n1232) );
NAND2_X1 U980 ( .A1(n1048), .A2(n1272), .ZN(n1271) );
NAND3_X1 U981 ( .A1(n1109), .A2(n1225), .A3(G902), .ZN(n1272) );
NOR2_X1 U982 ( .A1(G898), .A2(n1012), .ZN(n1109) );
NAND3_X1 U983 ( .A1(n1225), .A2(n1012), .A3(G952), .ZN(n1048) );
NAND2_X1 U984 ( .A1(G237), .A2(G234), .ZN(n1225) );
NOR2_X1 U985 ( .A1(n1047), .A2(n1046), .ZN(n1185) );
INV_X1 U986 ( .A(n1218), .ZN(n1046) );
NAND2_X1 U987 ( .A1(G214), .A2(n1273), .ZN(n1218) );
XOR2_X1 U988 ( .A(n1066), .B(n1063), .Z(n1047) );
AND3_X1 U989 ( .A1(n1274), .A2(n1262), .A3(n1275), .ZN(n1063) );
XOR2_X1 U990 ( .A(n1276), .B(KEYINPUT57), .Z(n1275) );
OR2_X1 U991 ( .A1(n1196), .A2(n1277), .ZN(n1276) );
NAND2_X1 U992 ( .A1(n1277), .A2(n1196), .ZN(n1274) );
NAND3_X1 U993 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1196) );
NAND2_X1 U994 ( .A1(KEYINPUT45), .A2(n1281), .ZN(n1280) );
NAND3_X1 U995 ( .A1(n1282), .A2(n1283), .A3(n1116), .ZN(n1279) );
INV_X1 U996 ( .A(KEYINPUT45), .ZN(n1283) );
OR2_X1 U997 ( .A1(n1116), .A2(n1282), .ZN(n1278) );
NOR2_X1 U998 ( .A1(KEYINPUT4), .A2(n1281), .ZN(n1282) );
XNOR2_X1 U999 ( .A(n1122), .B(n1284), .ZN(n1281) );
NOR2_X1 U1000 ( .A1(n1121), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U1001 ( .A(KEYINPUT55), .B(KEYINPUT24), .ZN(n1285) );
XOR2_X1 U1002 ( .A(n1286), .B(n1287), .Z(n1121) );
XOR2_X1 U1003 ( .A(G116), .B(G113), .Z(n1287) );
NAND2_X1 U1004 ( .A1(KEYINPUT39), .A2(n1230), .ZN(n1286) );
XOR2_X1 U1005 ( .A(n1165), .B(KEYINPUT31), .Z(n1122) );
INV_X1 U1006 ( .A(n1119), .ZN(n1116) );
XOR2_X1 U1007 ( .A(G110), .B(G122), .Z(n1119) );
NAND2_X1 U1008 ( .A1(n1288), .A2(n1289), .ZN(n1277) );
NAND2_X1 U1009 ( .A1(n1201), .A2(n1290), .ZN(n1289) );
NAND2_X1 U1010 ( .A1(n1291), .A2(n1292), .ZN(n1288) );
XNOR2_X1 U1011 ( .A(n1201), .B(n1293), .ZN(n1292) );
XOR2_X1 U1012 ( .A(KEYINPUT46), .B(KEYINPUT25), .Z(n1293) );
XNOR2_X1 U1013 ( .A(n1294), .B(n1085), .ZN(n1201) );
XOR2_X1 U1014 ( .A(n1223), .B(KEYINPUT53), .Z(n1294) );
INV_X1 U1015 ( .A(G125), .ZN(n1223) );
INV_X1 U1016 ( .A(n1290), .ZN(n1291) );
XOR2_X1 U1017 ( .A(n1199), .B(KEYINPUT29), .Z(n1290) );
NAND2_X1 U1018 ( .A1(G224), .A2(n1012), .ZN(n1199) );
NAND2_X1 U1019 ( .A1(G210), .A2(n1273), .ZN(n1066) );
NAND2_X1 U1020 ( .A1(n1244), .A2(n1262), .ZN(n1273) );
INV_X1 U1021 ( .A(n1182), .ZN(n1039) );
NOR2_X1 U1022 ( .A1(n1042), .A2(n1041), .ZN(n1182) );
AND2_X1 U1023 ( .A1(G221), .A2(n1261), .ZN(n1041) );
NAND2_X1 U1024 ( .A1(G234), .A2(n1262), .ZN(n1261) );
XOR2_X1 U1025 ( .A(n1295), .B(G469), .Z(n1042) );
NAND2_X1 U1026 ( .A1(n1296), .A2(n1262), .ZN(n1295) );
XOR2_X1 U1027 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U1028 ( .A(n1152), .B(n1299), .Z(n1298) );
NAND2_X1 U1029 ( .A1(KEYINPUT27), .A2(n1153), .ZN(n1299) );
XOR2_X1 U1030 ( .A(n1300), .B(n1301), .Z(n1297) );
INV_X1 U1031 ( .A(n1165), .ZN(n1301) );
XOR2_X1 U1032 ( .A(n1222), .B(n1302), .Z(n1165) );
XOR2_X1 U1033 ( .A(G107), .B(G104), .Z(n1302) );
NAND2_X1 U1034 ( .A1(KEYINPUT1), .A2(n1155), .ZN(n1300) );
XNOR2_X1 U1035 ( .A(n1303), .B(n1268), .ZN(n1155) );
XOR2_X1 U1036 ( .A(G110), .B(G140), .Z(n1268) );
NAND2_X1 U1037 ( .A1(G227), .A2(n1012), .ZN(n1303) );
XOR2_X1 U1038 ( .A(n1068), .B(G472), .Z(n1226) );
AND3_X1 U1039 ( .A1(n1304), .A2(n1305), .A3(n1262), .ZN(n1068) );
INV_X1 U1040 ( .A(G902), .ZN(n1262) );
NAND2_X1 U1041 ( .A1(n1306), .A2(n1152), .ZN(n1305) );
NAND2_X1 U1042 ( .A1(n1307), .A2(n1308), .ZN(n1304) );
INV_X1 U1043 ( .A(n1152), .ZN(n1308) );
NAND3_X1 U1044 ( .A1(n1309), .A2(n1310), .A3(n1311), .ZN(n1152) );
OR2_X1 U1045 ( .A1(n1089), .A2(KEYINPUT38), .ZN(n1311) );
NAND3_X1 U1046 ( .A1(KEYINPUT38), .A2(n1089), .A3(n1093), .ZN(n1310) );
INV_X1 U1047 ( .A(G131), .ZN(n1089) );
NAND2_X1 U1048 ( .A1(n1312), .A2(n1313), .ZN(n1309) );
NAND2_X1 U1049 ( .A1(KEYINPUT38), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1050 ( .A(KEYINPUT52), .B(G131), .Z(n1314) );
INV_X1 U1051 ( .A(n1093), .ZN(n1312) );
XNOR2_X1 U1052 ( .A(G134), .B(G137), .ZN(n1093) );
XOR2_X1 U1053 ( .A(n1315), .B(n1306), .Z(n1307) );
XOR2_X1 U1054 ( .A(n1085), .B(n1316), .Z(n1306) );
XNOR2_X1 U1055 ( .A(n1317), .B(n1318), .ZN(n1316) );
NOR2_X1 U1056 ( .A1(KEYINPUT22), .A2(n1148), .ZN(n1318) );
AND2_X1 U1057 ( .A1(n1319), .A2(n1320), .ZN(n1148) );
NAND2_X1 U1058 ( .A1(n1321), .A2(n1222), .ZN(n1320) );
INV_X1 U1059 ( .A(G101), .ZN(n1222) );
NAND3_X1 U1060 ( .A1(n1244), .A2(n1012), .A3(G210), .ZN(n1321) );
NAND4_X1 U1061 ( .A1(n1244), .A2(n1012), .A3(G210), .A4(G101), .ZN(n1319) );
INV_X1 U1062 ( .A(G953), .ZN(n1012) );
INV_X1 U1063 ( .A(G237), .ZN(n1244) );
NAND2_X1 U1064 ( .A1(KEYINPUT60), .A2(n1147), .ZN(n1317) );
XNOR2_X1 U1065 ( .A(n1322), .B(G113), .ZN(n1147) );
NAND3_X1 U1066 ( .A1(n1323), .A2(n1324), .A3(n1325), .ZN(n1322) );
NAND2_X1 U1067 ( .A1(KEYINPUT21), .A2(G116), .ZN(n1325) );
NAND3_X1 U1068 ( .A1(n1326), .A2(n1327), .A3(n1230), .ZN(n1324) );
INV_X1 U1069 ( .A(KEYINPUT21), .ZN(n1327) );
OR2_X1 U1070 ( .A1(n1230), .A2(n1326), .ZN(n1323) );
NOR2_X1 U1071 ( .A1(G116), .A2(KEYINPUT41), .ZN(n1326) );
INV_X1 U1072 ( .A(G119), .ZN(n1230) );
INV_X1 U1073 ( .A(n1153), .ZN(n1085) );
XOR2_X1 U1074 ( .A(n1219), .B(n1328), .Z(n1153) );
XOR2_X1 U1075 ( .A(G146), .B(G143), .Z(n1328) );
INV_X1 U1076 ( .A(G128), .ZN(n1219) );
XNOR2_X1 U1077 ( .A(KEYINPUT62), .B(KEYINPUT37), .ZN(n1315) );
endmodule


