//Key = 0000001010000010010111001110100010000000110000101100010001110000


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140;

XOR2_X2 U1214 ( .A(n1889), .B(KEYINPUT13), .Z(n1927) );
INV_X2 U1215 ( .A(n1830), .ZN(n1756) );
INV_X2 U1216 ( .A(U280), .ZN(n1757) );
INV_X1 U1217 ( .A(n1611), .ZN(U375) );
NAND2_X1 U1218 ( .A1(n1612), .A2(n1613), .ZN(U344) );
NAND2_X1 U1219 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1614), .ZN(n1613) );
NAND2_X1 U1220 ( .A1(DATA_IN_7_), .A2(n1615), .ZN(n1612) );
NAND2_X1 U1221 ( .A1(n1616), .A2(n1617), .ZN(U343) );
NAND2_X1 U1222 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1614), .ZN(n1617) );
NAND2_X1 U1223 ( .A1(DATA_IN_6_), .A2(n1615), .ZN(n1616) );
NAND2_X1 U1224 ( .A1(n1618), .A2(n1619), .ZN(U342) );
NAND2_X1 U1225 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1614), .ZN(n1619) );
NAND2_X1 U1226 ( .A1(DATA_IN_5_), .A2(n1615), .ZN(n1618) );
NAND2_X1 U1227 ( .A1(n1620), .A2(n1621), .ZN(U341) );
NAND2_X1 U1228 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1614), .ZN(n1621) );
NAND2_X1 U1229 ( .A1(DATA_IN_4_), .A2(n1615), .ZN(n1620) );
NAND2_X1 U1230 ( .A1(n1622), .A2(n1623), .ZN(U340) );
NAND2_X1 U1231 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1614), .ZN(n1623) );
NAND2_X1 U1232 ( .A1(DATA_IN_3_), .A2(n1615), .ZN(n1622) );
NAND2_X1 U1233 ( .A1(n1624), .A2(n1625), .ZN(U339) );
NAND2_X1 U1234 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1614), .ZN(n1625) );
NAND2_X1 U1235 ( .A1(DATA_IN_2_), .A2(n1615), .ZN(n1624) );
NAND2_X1 U1236 ( .A1(n1626), .A2(n1627), .ZN(U338) );
NAND2_X1 U1237 ( .A1(n1628), .A2(RMAX_REG_1__SCAN_IN), .ZN(n1627) );
XOR2_X1 U1238 ( .A(n1614), .B(KEYINPUT45), .Z(n1628) );
NAND2_X1 U1239 ( .A1(DATA_IN_1_), .A2(n1615), .ZN(n1626) );
NAND2_X1 U1240 ( .A1(n1629), .A2(n1630), .ZN(U337) );
NAND2_X1 U1241 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1614), .ZN(n1630) );
NAND2_X1 U1242 ( .A1(n1611), .A2(n1631), .ZN(n1614) );
NAND2_X1 U1243 ( .A1(n1632), .A2(n1633), .ZN(n1631) );
NAND2_X1 U1244 ( .A1(DATA_IN_0_), .A2(n1615), .ZN(n1629) );
NAND2_X1 U1245 ( .A1(n1634), .A2(n1635), .ZN(n1615) );
NAND2_X1 U1246 ( .A1(n1636), .A2(n1637), .ZN(n1635) );
XOR2_X1 U1247 ( .A(STATO_REG_1__SCAN_IN), .B(KEYINPUT16), .Z(n1636) );
NAND2_X1 U1248 ( .A1(n1638), .A2(n1639), .ZN(U336) );
NAND2_X1 U1249 ( .A1(DATA_IN_7_), .A2(n1640), .ZN(n1639) );
NAND2_X1 U1250 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1641), .ZN(n1638) );
NAND2_X1 U1251 ( .A1(n1642), .A2(n1643), .ZN(U335) );
NAND2_X1 U1252 ( .A1(DATA_IN_6_), .A2(n1640), .ZN(n1643) );
NAND2_X1 U1253 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1641), .ZN(n1642) );
NAND2_X1 U1254 ( .A1(n1644), .A2(n1645), .ZN(U334) );
NAND2_X1 U1255 ( .A1(DATA_IN_5_), .A2(n1640), .ZN(n1645) );
NAND2_X1 U1256 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1641), .ZN(n1644) );
NAND2_X1 U1257 ( .A1(n1646), .A2(n1647), .ZN(U333) );
NAND2_X1 U1258 ( .A1(DATA_IN_4_), .A2(n1640), .ZN(n1647) );
NAND2_X1 U1259 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1641), .ZN(n1646) );
NAND2_X1 U1260 ( .A1(n1648), .A2(n1649), .ZN(U332) );
NAND2_X1 U1261 ( .A1(DATA_IN_3_), .A2(n1640), .ZN(n1649) );
NAND2_X1 U1262 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1641), .ZN(n1648) );
NAND2_X1 U1263 ( .A1(n1650), .A2(n1651), .ZN(U331) );
NAND2_X1 U1264 ( .A1(DATA_IN_2_), .A2(n1640), .ZN(n1651) );
NAND2_X1 U1265 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1641), .ZN(n1650) );
NAND2_X1 U1266 ( .A1(n1652), .A2(n1653), .ZN(U330) );
NAND2_X1 U1267 ( .A1(DATA_IN_1_), .A2(n1640), .ZN(n1653) );
NAND2_X1 U1268 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1641), .ZN(n1652) );
NAND2_X1 U1269 ( .A1(n1654), .A2(n1655), .ZN(U329) );
NAND2_X1 U1270 ( .A1(DATA_IN_0_), .A2(n1640), .ZN(n1655) );
NAND2_X1 U1271 ( .A1(n1634), .A2(n1656), .ZN(n1640) );
OR2_X1 U1272 ( .A1(n1657), .A2(n1658), .ZN(n1656) );
NAND2_X1 U1273 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1641), .ZN(n1654) );
NAND2_X1 U1274 ( .A1(n1611), .A2(n1659), .ZN(n1641) );
NAND2_X1 U1275 ( .A1(n1634), .A2(n1657), .ZN(n1659) );
NAND2_X1 U1276 ( .A1(n1632), .A2(n1660), .ZN(n1657) );
NAND2_X1 U1277 ( .A1(n1661), .A2(n1662), .ZN(n1660) );
NAND3_X1 U1278 ( .A1(n1663), .A2(n1664), .A3(n1665), .ZN(n1662) );
NAND2_X1 U1279 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1666), .ZN(n1665) );
NAND3_X1 U1280 ( .A1(n1667), .A2(n1668), .A3(n1669), .ZN(n1664) );
NAND2_X1 U1281 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1670), .ZN(n1669) );
NAND3_X1 U1282 ( .A1(n1671), .A2(n1672), .A3(n1673), .ZN(n1668) );
NAND2_X1 U1283 ( .A1(DATA_IN_5_), .A2(n1674), .ZN(n1673) );
NAND3_X1 U1284 ( .A1(n1675), .A2(n1676), .A3(n1677), .ZN(n1672) );
XOR2_X1 U1285 ( .A(n1678), .B(KEYINPUT9), .Z(n1677) );
NAND3_X1 U1286 ( .A1(n1679), .A2(n1680), .A3(n1681), .ZN(n1678) );
NAND2_X1 U1287 ( .A1(DATA_IN_3_), .A2(n1682), .ZN(n1681) );
NAND3_X1 U1288 ( .A1(n1683), .A2(n1684), .A3(n1685), .ZN(n1680) );
NAND2_X1 U1289 ( .A1(n1686), .A2(RMIN_REG_2__SCAN_IN), .ZN(n1685) );
XNOR2_X1 U1290 ( .A(DATA_IN_2_), .B(KEYINPUT63), .ZN(n1686) );
NAND3_X1 U1291 ( .A1(n1687), .A2(n1688), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1684) );
INV_X1 U1292 ( .A(DATA_IN_0_), .ZN(n1688) );
NAND2_X1 U1293 ( .A1(DATA_IN_1_), .A2(n1689), .ZN(n1687) );
NAND2_X1 U1294 ( .A1(n1690), .A2(n1691), .ZN(n1683) );
XOR2_X1 U1295 ( .A(RMIN_REG_1__SCAN_IN), .B(KEYINPUT56), .Z(n1690) );
NAND2_X1 U1296 ( .A1(DATA_IN_2_), .A2(n1692), .ZN(n1679) );
NAND2_X1 U1297 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1693), .ZN(n1676) );
NAND2_X1 U1298 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1694), .ZN(n1675) );
NAND2_X1 U1299 ( .A1(DATA_IN_4_), .A2(n1695), .ZN(n1671) );
NAND2_X1 U1300 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1696), .ZN(n1667) );
NAND2_X1 U1301 ( .A1(DATA_IN_6_), .A2(n1697), .ZN(n1663) );
NAND2_X1 U1302 ( .A1(DATA_IN_7_), .A2(n1698), .ZN(n1661) );
INV_X1 U1303 ( .A(n1637), .ZN(n1632) );
NAND2_X1 U1304 ( .A1(n1699), .A2(n1700), .ZN(n1637) );
NAND2_X1 U1305 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1666), .ZN(n1700) );
INV_X1 U1306 ( .A(DATA_IN_7_), .ZN(n1666) );
NAND3_X1 U1307 ( .A1(n1701), .A2(n1702), .A3(n1703), .ZN(n1699) );
NAND2_X1 U1308 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1670), .ZN(n1703) );
NAND3_X1 U1309 ( .A1(n1704), .A2(n1705), .A3(n1706), .ZN(n1702) );
XOR2_X1 U1310 ( .A(n1707), .B(KEYINPUT37), .Z(n1706) );
NAND3_X1 U1311 ( .A1(n1708), .A2(n1709), .A3(n1710), .ZN(n1707) );
NAND2_X1 U1312 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1696), .ZN(n1710) );
INV_X1 U1313 ( .A(DATA_IN_5_), .ZN(n1696) );
NAND3_X1 U1314 ( .A1(n1711), .A2(n1712), .A3(n1713), .ZN(n1709) );
NAND2_X1 U1315 ( .A1(DATA_IN_4_), .A2(n1714), .ZN(n1713) );
NAND3_X1 U1316 ( .A1(n1715), .A2(n1716), .A3(n1717), .ZN(n1712) );
NAND2_X1 U1317 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1693), .ZN(n1717) );
NAND3_X1 U1318 ( .A1(n1718), .A2(n1719), .A3(n1720), .ZN(n1716) );
NAND2_X1 U1319 ( .A1(DATA_IN_2_), .A2(n1721), .ZN(n1720) );
NAND3_X1 U1320 ( .A1(n1722), .A2(n1723), .A3(DATA_IN_0_), .ZN(n1719) );
INV_X1 U1321 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1723) );
NAND2_X1 U1322 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1691), .ZN(n1722) );
NAND2_X1 U1323 ( .A1(DATA_IN_1_), .A2(n1724), .ZN(n1718) );
NAND2_X1 U1324 ( .A1(n1725), .A2(RMAX_REG_2__SCAN_IN), .ZN(n1715) );
XNOR2_X1 U1325 ( .A(DATA_IN_2_), .B(KEYINPUT1), .ZN(n1725) );
NAND2_X1 U1326 ( .A1(DATA_IN_3_), .A2(n1726), .ZN(n1711) );
NAND2_X1 U1327 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1694), .ZN(n1708) );
INV_X1 U1328 ( .A(DATA_IN_4_), .ZN(n1694) );
NAND2_X1 U1329 ( .A1(DATA_IN_5_), .A2(n1727), .ZN(n1705) );
XOR2_X1 U1330 ( .A(RMAX_REG_5__SCAN_IN), .B(KEYINPUT53), .Z(n1727) );
NAND2_X1 U1331 ( .A1(DATA_IN_6_), .A2(n1728), .ZN(n1704) );
NAND2_X1 U1332 ( .A1(n1729), .A2(DATA_IN_7_), .ZN(n1701) );
XNOR2_X1 U1333 ( .A(RMAX_REG_7__SCAN_IN), .B(KEYINPUT5), .ZN(n1729) );
NAND2_X1 U1334 ( .A1(n1730), .A2(n1731), .ZN(U328) );
NAND2_X1 U1335 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1732), .ZN(n1731) );
XNOR2_X1 U1336 ( .A(KEYINPUT6), .B(n1733), .ZN(n1732) );
NAND2_X1 U1337 ( .A1(n1734), .A2(DATA_IN_7_), .ZN(n1730) );
NAND2_X1 U1338 ( .A1(n1735), .A2(n1736), .ZN(U327) );
NAND2_X1 U1339 ( .A1(DATA_IN_6_), .A2(n1737), .ZN(n1736) );
XOR2_X1 U1340 ( .A(KEYINPUT60), .B(n1734), .Z(n1737) );
NAND2_X1 U1341 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1733), .ZN(n1735) );
NAND2_X1 U1342 ( .A1(n1738), .A2(n1739), .ZN(U326) );
NAND2_X1 U1343 ( .A1(n1734), .A2(DATA_IN_5_), .ZN(n1739) );
XOR2_X1 U1344 ( .A(KEYINPUT20), .B(n1740), .Z(n1738) );
AND2_X1 U1345 ( .A1(n1733), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1740) );
NAND2_X1 U1346 ( .A1(n1741), .A2(n1742), .ZN(U325) );
NAND2_X1 U1347 ( .A1(n1734), .A2(DATA_IN_4_), .ZN(n1742) );
NAND2_X1 U1348 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1733), .ZN(n1741) );
NAND2_X1 U1349 ( .A1(n1743), .A2(n1744), .ZN(U324) );
NAND2_X1 U1350 ( .A1(n1745), .A2(RLAST_REG_3__SCAN_IN), .ZN(n1744) );
XOR2_X1 U1351 ( .A(n1733), .B(KEYINPUT47), .Z(n1745) );
NAND2_X1 U1352 ( .A1(n1734), .A2(DATA_IN_3_), .ZN(n1743) );
NAND2_X1 U1353 ( .A1(n1746), .A2(n1747), .ZN(U323) );
NAND2_X1 U1354 ( .A1(n1734), .A2(DATA_IN_2_), .ZN(n1747) );
NAND2_X1 U1355 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1733), .ZN(n1746) );
NAND2_X1 U1356 ( .A1(n1748), .A2(n1749), .ZN(U322) );
NAND2_X1 U1357 ( .A1(n1734), .A2(DATA_IN_1_), .ZN(n1749) );
NAND2_X1 U1358 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1733), .ZN(n1748) );
NAND2_X1 U1359 ( .A1(n1750), .A2(n1751), .ZN(U321) );
NAND2_X1 U1360 ( .A1(n1734), .A2(DATA_IN_0_), .ZN(n1751) );
AND2_X1 U1361 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1752), .ZN(n1734) );
NAND2_X1 U1362 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1733), .ZN(n1750) );
NAND2_X1 U1363 ( .A1(n1611), .A2(n1752), .ZN(n1733) );
NAND2_X1 U1364 ( .A1(n1753), .A2(n1633), .ZN(n1752) );
NAND2_X1 U1365 ( .A1(n1633), .A2(n1658), .ZN(n1611) );
NAND2_X1 U1366 ( .A1(n1754), .A2(n1755), .ZN(U320) );
NAND2_X1 U1367 ( .A1(n1756), .A2(DATA_IN_7_), .ZN(n1755) );
NAND2_X1 U1368 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1757), .ZN(n1754) );
NAND2_X1 U1369 ( .A1(n1758), .A2(n1759), .ZN(U319) );
NAND2_X1 U1370 ( .A1(n1756), .A2(DATA_IN_6_), .ZN(n1759) );
NAND2_X1 U1371 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1757), .ZN(n1758) );
NAND2_X1 U1372 ( .A1(n1760), .A2(n1761), .ZN(U318) );
NAND2_X1 U1373 ( .A1(n1756), .A2(DATA_IN_5_), .ZN(n1761) );
NAND2_X1 U1374 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1757), .ZN(n1760) );
NAND2_X1 U1375 ( .A1(n1762), .A2(n1763), .ZN(U317) );
NAND2_X1 U1376 ( .A1(n1756), .A2(DATA_IN_4_), .ZN(n1763) );
NAND2_X1 U1377 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1757), .ZN(n1762) );
NAND2_X1 U1378 ( .A1(n1764), .A2(n1765), .ZN(U316) );
NAND2_X1 U1379 ( .A1(n1756), .A2(DATA_IN_3_), .ZN(n1765) );
NAND2_X1 U1380 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1757), .ZN(n1764) );
NAND2_X1 U1381 ( .A1(n1766), .A2(n1767), .ZN(U315) );
NAND2_X1 U1382 ( .A1(n1756), .A2(DATA_IN_2_), .ZN(n1767) );
NAND2_X1 U1383 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1757), .ZN(n1766) );
NAND2_X1 U1384 ( .A1(n1768), .A2(n1769), .ZN(U314) );
NAND2_X1 U1385 ( .A1(DATA_IN_1_), .A2(n1770), .ZN(n1769) );
XOR2_X1 U1386 ( .A(KEYINPUT7), .B(n1756), .Z(n1770) );
NAND2_X1 U1387 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1757), .ZN(n1768) );
NAND2_X1 U1388 ( .A1(n1771), .A2(n1772), .ZN(U313) );
NAND2_X1 U1389 ( .A1(n1756), .A2(DATA_IN_0_), .ZN(n1772) );
NAND2_X1 U1390 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1757), .ZN(n1771) );
NAND2_X1 U1391 ( .A1(n1773), .A2(n1774), .ZN(U312) );
NAND2_X1 U1392 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1756), .ZN(n1774) );
NAND2_X1 U1393 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1757), .ZN(n1773) );
NAND2_X1 U1394 ( .A1(n1775), .A2(n1776), .ZN(U311) );
NAND2_X1 U1395 ( .A1(n1756), .A2(n1777), .ZN(n1776) );
XOR2_X1 U1396 ( .A(REG1_REG_6__SCAN_IN), .B(KEYINPUT35), .Z(n1777) );
NAND2_X1 U1397 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1757), .ZN(n1775) );
NAND2_X1 U1398 ( .A1(n1778), .A2(n1779), .ZN(U310) );
NAND2_X1 U1399 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1756), .ZN(n1779) );
NAND2_X1 U1400 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1757), .ZN(n1778) );
NAND2_X1 U1401 ( .A1(n1780), .A2(n1781), .ZN(U309) );
NAND2_X1 U1402 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1756), .ZN(n1781) );
NAND2_X1 U1403 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1757), .ZN(n1780) );
NAND2_X1 U1404 ( .A1(n1782), .A2(n1783), .ZN(U308) );
NAND2_X1 U1405 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1756), .ZN(n1783) );
NAND2_X1 U1406 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1757), .ZN(n1782) );
NAND2_X1 U1407 ( .A1(n1784), .A2(n1785), .ZN(U307) );
NAND2_X1 U1408 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1756), .ZN(n1785) );
NAND2_X1 U1409 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1757), .ZN(n1784) );
NAND2_X1 U1410 ( .A1(n1786), .A2(n1787), .ZN(U306) );
NAND2_X1 U1411 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1756), .ZN(n1787) );
NAND2_X1 U1412 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1757), .ZN(n1786) );
NAND2_X1 U1413 ( .A1(n1788), .A2(n1789), .ZN(U305) );
NAND2_X1 U1414 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1756), .ZN(n1789) );
NAND2_X1 U1415 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1757), .ZN(n1788) );
NAND2_X1 U1416 ( .A1(n1790), .A2(n1791), .ZN(U304) );
NAND2_X1 U1417 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1756), .ZN(n1791) );
NAND2_X1 U1418 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1757), .ZN(n1790) );
NAND2_X1 U1419 ( .A1(n1792), .A2(n1793), .ZN(U303) );
NAND2_X1 U1420 ( .A1(n1794), .A2(n1756), .ZN(n1793) );
XNOR2_X1 U1421 ( .A(REG2_REG_6__SCAN_IN), .B(KEYINPUT21), .ZN(n1794) );
NAND2_X1 U1422 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1757), .ZN(n1792) );
NAND2_X1 U1423 ( .A1(n1795), .A2(n1796), .ZN(U302) );
NAND2_X1 U1424 ( .A1(n1797), .A2(n1757), .ZN(n1796) );
XOR2_X1 U1425 ( .A(REG3_REG_5__SCAN_IN), .B(KEYINPUT44), .Z(n1797) );
NAND2_X1 U1426 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1756), .ZN(n1795) );
NAND2_X1 U1427 ( .A1(n1798), .A2(n1799), .ZN(U301) );
NAND2_X1 U1428 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1757), .ZN(n1799) );
XOR2_X1 U1429 ( .A(KEYINPUT19), .B(n1800), .Z(n1798) );
AND2_X1 U1430 ( .A1(n1756), .A2(REG2_REG_4__SCAN_IN), .ZN(n1800) );
NAND2_X1 U1431 ( .A1(n1801), .A2(n1802), .ZN(U300) );
NAND2_X1 U1432 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1756), .ZN(n1802) );
NAND2_X1 U1433 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1757), .ZN(n1801) );
NAND2_X1 U1434 ( .A1(n1803), .A2(n1804), .ZN(U299) );
NAND2_X1 U1435 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1756), .ZN(n1804) );
NAND2_X1 U1436 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1757), .ZN(n1803) );
NAND2_X1 U1437 ( .A1(n1805), .A2(n1806), .ZN(U298) );
NAND2_X1 U1438 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1756), .ZN(n1806) );
NAND2_X1 U1439 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1757), .ZN(n1805) );
NAND2_X1 U1440 ( .A1(n1807), .A2(n1808), .ZN(U297) );
NAND2_X1 U1441 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1809), .ZN(n1808) );
XOR2_X1 U1442 ( .A(KEYINPUT43), .B(n1757), .Z(n1809) );
NAND2_X1 U1443 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1756), .ZN(n1807) );
NAND2_X1 U1444 ( .A1(n1810), .A2(n1811), .ZN(U296) );
NAND2_X1 U1445 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1756), .ZN(n1811) );
NAND2_X1 U1446 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1757), .ZN(n1810) );
NAND2_X1 U1447 ( .A1(n1812), .A2(n1813), .ZN(U295) );
NAND2_X1 U1448 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1756), .ZN(n1813) );
NAND2_X1 U1449 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1757), .ZN(n1812) );
NAND2_X1 U1450 ( .A1(n1814), .A2(n1815), .ZN(U294) );
NAND2_X1 U1451 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1756), .ZN(n1815) );
NAND2_X1 U1452 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1757), .ZN(n1814) );
NAND2_X1 U1453 ( .A1(n1816), .A2(n1817), .ZN(U293) );
NAND2_X1 U1454 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1818), .ZN(n1817) );
XOR2_X1 U1455 ( .A(KEYINPUT36), .B(n1756), .Z(n1818) );
NAND2_X1 U1456 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1757), .ZN(n1816) );
NAND2_X1 U1457 ( .A1(n1819), .A2(n1820), .ZN(U292) );
NAND2_X1 U1458 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1756), .ZN(n1820) );
NAND2_X1 U1459 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1757), .ZN(n1819) );
NAND2_X1 U1460 ( .A1(n1821), .A2(n1822), .ZN(U291) );
NAND2_X1 U1461 ( .A1(n1756), .A2(n1823), .ZN(n1822) );
XOR2_X1 U1462 ( .A(REG3_REG_2__SCAN_IN), .B(KEYINPUT11), .Z(n1823) );
NAND2_X1 U1463 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1757), .ZN(n1821) );
NAND2_X1 U1464 ( .A1(n1824), .A2(n1825), .ZN(U290) );
NAND2_X1 U1465 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1757), .ZN(n1825) );
XOR2_X1 U1466 ( .A(n1826), .B(KEYINPUT0), .Z(n1824) );
NAND2_X1 U1467 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1756), .ZN(n1826) );
NAND2_X1 U1468 ( .A1(n1827), .A2(n1828), .ZN(U289) );
NAND2_X1 U1469 ( .A1(n1829), .A2(REG4_REG_0__SCAN_IN), .ZN(n1828) );
XOR2_X1 U1470 ( .A(U280), .B(KEYINPUT57), .Z(n1829) );
NAND2_X1 U1471 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1756), .ZN(n1827) );
NAND4_X1 U1472 ( .A1(n1831), .A2(n1832), .A3(n1833), .A4(n1834), .ZN(U288));
NAND2_X1 U1473 ( .A1(n1835), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1834) );
NOR2_X1 U1474 ( .A1(n1836), .A2(n1837), .ZN(n1833) );
NOR2_X1 U1475 ( .A1(n1838), .A2(n1839), .ZN(n1837) );
XNOR2_X1 U1476 ( .A(n1840), .B(KEYINPUT15), .ZN(n1838) );
NAND2_X1 U1477 ( .A1(n1841), .A2(REG4_REG_7__SCAN_IN), .ZN(n1832) );
NAND2_X1 U1478 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1757), .ZN(n1831) );
NAND4_X1 U1479 ( .A1(n1842), .A2(n1843), .A3(n1844), .A4(n1845), .ZN(U287));
NOR3_X1 U1480 ( .A1(n1846), .A2(n1836), .A3(n1847), .ZN(n1845) );
NOR3_X1 U1481 ( .A1(n1848), .A2(n1849), .A3(n1850), .ZN(n1847) );
XNOR2_X1 U1482 ( .A(n1851), .B(n1852), .ZN(n1850) );
XOR2_X1 U1483 ( .A(KEYINPUT39), .B(KEYINPUT3), .Z(n1852) );
AND3_X1 U1484 ( .A1(n1853), .A2(n1849), .A3(n1854), .ZN(n1836) );
XNOR2_X1 U1485 ( .A(n1851), .B(KEYINPUT30), .ZN(n1854) );
NOR2_X1 U1486 ( .A1(n1855), .A2(n1839), .ZN(n1846) );
NOR2_X1 U1487 ( .A1(n1856), .A2(n1840), .ZN(n1855) );
AND3_X1 U1488 ( .A1(n1857), .A2(n1858), .A3(n1859), .ZN(n1840) );
XOR2_X1 U1489 ( .A(n1860), .B(KEYINPUT62), .Z(n1859) );
NOR2_X1 U1490 ( .A1(n1857), .A2(n1860), .ZN(n1856) );
NAND2_X1 U1491 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1757), .ZN(n1844) );
NAND2_X1 U1492 ( .A1(n1835), .A2(RLAST_REG_6__SCAN_IN), .ZN(n1843) );
NAND2_X1 U1493 ( .A1(n1841), .A2(REG4_REG_6__SCAN_IN), .ZN(n1842) );
NAND4_X1 U1494 ( .A1(n1861), .A2(n1862), .A3(n1863), .A4(n1864), .ZN(U286));
NOR3_X1 U1495 ( .A1(n1865), .A2(n1866), .A3(n1867), .ZN(n1864) );
NOR3_X1 U1496 ( .A1(n1848), .A2(n1851), .A3(n1868), .ZN(n1867) );
NOR2_X1 U1497 ( .A1(n1869), .A2(n1870), .ZN(n1868) );
AND2_X1 U1498 ( .A1(n1871), .A2(n1870), .ZN(n1851) );
NAND2_X1 U1499 ( .A1(n1872), .A2(n1873), .ZN(n1870) );
OR2_X1 U1500 ( .A1(n1857), .A2(n1858), .ZN(n1873) );
XOR2_X1 U1501 ( .A(KEYINPUT48), .B(n1849), .Z(n1872) );
AND2_X1 U1502 ( .A1(n1874), .A2(n1875), .ZN(n1849) );
XOR2_X1 U1503 ( .A(KEYINPUT38), .B(n1858), .Z(n1875) );
XOR2_X1 U1504 ( .A(n1857), .B(KEYINPUT33), .Z(n1874) );
XNOR2_X1 U1505 ( .A(n1869), .B(n1876), .ZN(n1871) );
XOR2_X1 U1506 ( .A(KEYINPUT58), .B(KEYINPUT52), .Z(n1876) );
NOR3_X1 U1507 ( .A1(n1839), .A2(n1877), .A3(n1878), .ZN(n1866) );
NOR2_X1 U1508 ( .A1(n1879), .A2(n1880), .ZN(n1878) );
INV_X1 U1509 ( .A(n1860), .ZN(n1877) );
NAND2_X1 U1510 ( .A1(n1879), .A2(n1880), .ZN(n1860) );
XOR2_X1 U1511 ( .A(n1881), .B(n1857), .Z(n1880) );
NOR2_X1 U1512 ( .A1(n1857), .A2(n1882), .ZN(n1865) );
XOR2_X1 U1513 ( .A(n1883), .B(n1884), .Z(n1857) );
XOR2_X1 U1514 ( .A(n1885), .B(n1886), .Z(n1884) );
NOR2_X1 U1515 ( .A1(n1887), .A2(n1888), .ZN(n1886) );
NOR2_X1 U1516 ( .A1(n1728), .A2(n1889), .ZN(n1888) );
NOR2_X1 U1517 ( .A1(n1670), .A2(n1890), .ZN(n1887) );
NOR2_X1 U1518 ( .A1(n1891), .A2(n1892), .ZN(n1885) );
NOR2_X1 U1519 ( .A1(n1697), .A2(n1889), .ZN(n1892) );
NOR2_X1 U1520 ( .A1(n1893), .A2(n1890), .ZN(n1891) );
NAND2_X1 U1521 ( .A1(n1894), .A2(n1895), .ZN(n1883) );
NAND2_X1 U1522 ( .A1(n1896), .A2(n1897), .ZN(n1895) );
NAND2_X1 U1523 ( .A1(n1898), .A2(n1899), .ZN(n1896) );
OR2_X1 U1524 ( .A1(n1899), .A2(n1898), .ZN(n1894) );
NAND2_X1 U1525 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1757), .ZN(n1863) );
NAND2_X1 U1526 ( .A1(n1835), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1862) );
NAND2_X1 U1527 ( .A1(n1841), .A2(REG4_REG_5__SCAN_IN), .ZN(n1861) );
NAND4_X1 U1528 ( .A1(n1900), .A2(n1901), .A3(n1902), .A4(n1903), .ZN(U285));
NOR3_X1 U1529 ( .A1(n1904), .A2(n1905), .A3(n1906), .ZN(n1903) );
NOR3_X1 U1530 ( .A1(n1839), .A2(n1879), .A3(n1907), .ZN(n1906) );
NOR2_X1 U1531 ( .A1(n1908), .A2(n1909), .ZN(n1907) );
NOR2_X1 U1532 ( .A1(n1910), .A2(n1911), .ZN(n1908) );
NOR3_X1 U1533 ( .A1(n1912), .A2(n1910), .A3(n1911), .ZN(n1879) );
XOR2_X1 U1534 ( .A(KEYINPUT14), .B(n1909), .Z(n1912) );
NAND3_X1 U1535 ( .A1(n1913), .A2(n1914), .A3(n1881), .ZN(n1909) );
NAND2_X1 U1536 ( .A1(n1915), .A2(n1916), .ZN(n1914) );
INV_X1 U1537 ( .A(KEYINPUT2), .ZN(n1916) );
NAND2_X1 U1538 ( .A1(KEYINPUT2), .A2(n1917), .ZN(n1913) );
NOR3_X1 U1539 ( .A1(n1918), .A2(n1869), .A3(n1919), .ZN(n1905) );
NOR3_X1 U1540 ( .A1(n1915), .A2(n1858), .A3(n1920), .ZN(n1919) );
AND2_X1 U1541 ( .A1(n1920), .A2(n1921), .ZN(n1869) );
OR2_X1 U1542 ( .A1(n1858), .A2(n1915), .ZN(n1921) );
NOR2_X1 U1543 ( .A1(n1922), .A2(n1917), .ZN(n1915) );
INV_X1 U1544 ( .A(n1881), .ZN(n1858) );
NAND2_X1 U1545 ( .A1(n1917), .A2(n1922), .ZN(n1881) );
NOR2_X1 U1546 ( .A1(n1923), .A2(n1910), .ZN(n1920) );
XOR2_X1 U1547 ( .A(KEYINPUT28), .B(n1853), .Z(n1918) );
NOR2_X1 U1548 ( .A1(n1922), .A2(n1882), .ZN(n1904) );
XOR2_X1 U1549 ( .A(n1897), .B(n1924), .Z(n1922) );
XOR2_X1 U1550 ( .A(n1898), .B(n1899), .Z(n1924) );
NAND2_X1 U1551 ( .A1(n1925), .A2(n1926), .ZN(n1899) );
NAND2_X1 U1552 ( .A1(n1927), .A2(REG4_REG_5__SCAN_IN), .ZN(n1926) );
NAND2_X1 U1553 ( .A1(RESTART), .A2(RMIN_REG_5__SCAN_IN), .ZN(n1925) );
NAND2_X1 U1554 ( .A1(n1928), .A2(n1929), .ZN(n1898) );
NAND2_X1 U1555 ( .A1(n1927), .A2(DATA_IN_5_), .ZN(n1929) );
NAND2_X1 U1556 ( .A1(RESTART), .A2(RMAX_REG_5__SCAN_IN), .ZN(n1928) );
NAND2_X1 U1557 ( .A1(n1930), .A2(n1931), .ZN(n1897) );
NAND2_X1 U1558 ( .A1(n1932), .A2(n1933), .ZN(n1931) );
XOR2_X1 U1559 ( .A(n1934), .B(KEYINPUT51), .Z(n1932) );
NAND2_X1 U1560 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1757), .ZN(n1902) );
NAND2_X1 U1561 ( .A1(n1835), .A2(RLAST_REG_4__SCAN_IN), .ZN(n1901) );
NAND2_X1 U1562 ( .A1(n1841), .A2(REG4_REG_4__SCAN_IN), .ZN(n1900) );
NAND4_X1 U1563 ( .A1(n1935), .A2(n1936), .A3(n1937), .A4(n1938), .ZN(U284));
NOR3_X1 U1564 ( .A1(n1939), .A2(n1940), .A3(n1941), .ZN(n1938) );
NOR2_X1 U1565 ( .A1(n1942), .A2(n1943), .ZN(n1941) );
AND2_X1 U1566 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1835), .ZN(n1940) );
XNOR2_X1 U1567 ( .A(n1944), .B(KEYINPUT4), .ZN(n1939) );
NAND2_X1 U1568 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1757), .ZN(n1944) );
NAND2_X1 U1569 ( .A1(n1945), .A2(n1946), .ZN(n1937) );
NAND2_X1 U1570 ( .A1(n1947), .A2(n1948), .ZN(n1936) );
XOR2_X1 U1571 ( .A(n1911), .B(n1910), .Z(n1947) );
INV_X1 U1572 ( .A(n1949), .ZN(n1911) );
NAND2_X1 U1573 ( .A1(n1950), .A2(n1853), .ZN(n1935) );
XOR2_X1 U1574 ( .A(n1923), .B(n1910), .Z(n1950) );
NOR2_X1 U1575 ( .A1(n1917), .A2(n1951), .ZN(n1910) );
AND2_X1 U1576 ( .A1(n1946), .A2(n1952), .ZN(n1951) );
NOR2_X1 U1577 ( .A1(n1952), .A2(n1946), .ZN(n1917) );
NAND2_X1 U1578 ( .A1(n1953), .A2(n1954), .ZN(n1946) );
NAND2_X1 U1579 ( .A1(n1955), .A2(n1956), .ZN(n1954) );
NAND2_X1 U1580 ( .A1(n1933), .A2(n1930), .ZN(n1956) );
NAND2_X1 U1581 ( .A1(n1957), .A2(n1958), .ZN(n1930) );
NAND2_X1 U1582 ( .A1(n1959), .A2(n1960), .ZN(n1933) );
INV_X1 U1583 ( .A(n1934), .ZN(n1955) );
NAND2_X1 U1584 ( .A1(n1961), .A2(n1934), .ZN(n1953) );
NAND2_X1 U1585 ( .A1(n1962), .A2(n1963), .ZN(n1934) );
NAND2_X1 U1586 ( .A1(n1964), .A2(n1965), .ZN(n1963) );
NAND2_X1 U1587 ( .A1(n1966), .A2(n1967), .ZN(n1964) );
OR2_X1 U1588 ( .A1(n1967), .A2(n1966), .ZN(n1962) );
XOR2_X1 U1589 ( .A(n1958), .B(n1957), .Z(n1961) );
INV_X1 U1590 ( .A(n1960), .ZN(n1957) );
NAND2_X1 U1591 ( .A1(n1968), .A2(n1969), .ZN(n1960) );
NAND2_X1 U1592 ( .A1(n1927), .A2(REG4_REG_4__SCAN_IN), .ZN(n1969) );
NAND2_X1 U1593 ( .A1(RESTART), .A2(RMIN_REG_4__SCAN_IN), .ZN(n1968) );
INV_X1 U1594 ( .A(n1959), .ZN(n1958) );
NAND2_X1 U1595 ( .A1(n1970), .A2(n1971), .ZN(n1959) );
NAND2_X1 U1596 ( .A1(RESTART), .A2(n1972), .ZN(n1971) );
XOR2_X1 U1597 ( .A(RMAX_REG_4__SCAN_IN), .B(KEYINPUT42), .Z(n1972) );
NAND2_X1 U1598 ( .A1(n1927), .A2(DATA_IN_4_), .ZN(n1970) );
NAND4_X1 U1599 ( .A1(n1973), .A2(n1974), .A3(n1975), .A4(n1976), .ZN(U283));
NOR3_X1 U1600 ( .A1(n1977), .A2(n1978), .A3(n1979), .ZN(n1976) );
NOR2_X1 U1601 ( .A1(n1980), .A2(n1848), .ZN(n1979) );
XOR2_X1 U1602 ( .A(n1981), .B(KEYINPUT10), .Z(n1980) );
NAND2_X1 U1603 ( .A1(n1923), .A2(n1982), .ZN(n1981) );
NAND2_X1 U1604 ( .A1(n1983), .A2(n1984), .ZN(n1982) );
NAND2_X1 U1605 ( .A1(n1985), .A2(n1986), .ZN(n1984) );
NAND3_X1 U1606 ( .A1(n1986), .A2(n1987), .A3(n1985), .ZN(n1923) );
NOR3_X1 U1607 ( .A1(n1839), .A2(n1949), .A3(n1988), .ZN(n1978) );
AND2_X1 U1608 ( .A1(n1989), .A2(n1983), .ZN(n1988) );
NOR2_X1 U1609 ( .A1(n1989), .A2(n1983), .ZN(n1949) );
INV_X1 U1610 ( .A(n1987), .ZN(n1983) );
NAND2_X1 U1611 ( .A1(n1990), .A2(n1952), .ZN(n1987) );
OR2_X1 U1612 ( .A1(n1991), .A2(n1992), .ZN(n1952) );
NAND2_X1 U1613 ( .A1(n1992), .A2(n1991), .ZN(n1990) );
AND2_X1 U1614 ( .A1(n1992), .A2(n1945), .ZN(n1977) );
XNOR2_X1 U1615 ( .A(n1965), .B(n1993), .ZN(n1992) );
XOR2_X1 U1616 ( .A(n1966), .B(n1967), .Z(n1993) );
NAND2_X1 U1617 ( .A1(n1994), .A2(n1995), .ZN(n1967) );
NAND2_X1 U1618 ( .A1(n1927), .A2(DATA_IN_3_), .ZN(n1995) );
NAND2_X1 U1619 ( .A1(RESTART), .A2(RMAX_REG_3__SCAN_IN), .ZN(n1994) );
NAND2_X1 U1620 ( .A1(n1996), .A2(n1997), .ZN(n1966) );
NAND2_X1 U1621 ( .A1(n1927), .A2(REG4_REG_3__SCAN_IN), .ZN(n1997) );
NAND2_X1 U1622 ( .A1(RESTART), .A2(RMIN_REG_3__SCAN_IN), .ZN(n1996) );
NAND2_X1 U1623 ( .A1(n1998), .A2(n1999), .ZN(n1965) );
NAND2_X1 U1624 ( .A1(n2000), .A2(n2001), .ZN(n1999) );
NAND2_X1 U1625 ( .A1(n2002), .A2(n2003), .ZN(n2001) );
INV_X1 U1626 ( .A(n2004), .ZN(n2000) );
OR2_X1 U1627 ( .A1(n2002), .A2(n2003), .ZN(n1998) );
NAND2_X1 U1628 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1757), .ZN(n1975) );
NAND2_X1 U1629 ( .A1(n1835), .A2(RLAST_REG_2__SCAN_IN), .ZN(n1974) );
NAND2_X1 U1630 ( .A1(n1841), .A2(REG4_REG_2__SCAN_IN), .ZN(n1973) );
NAND4_X1 U1631 ( .A1(n2005), .A2(n2006), .A3(n2007), .A4(n2008), .ZN(U282));
NOR3_X1 U1632 ( .A1(n2009), .A2(n2010), .A3(n2011), .ZN(n2008) );
NOR2_X1 U1633 ( .A1(n1848), .A2(n2012), .ZN(n2011) );
XNOR2_X1 U1634 ( .A(n1986), .B(n1985), .ZN(n2012) );
NOR3_X1 U1635 ( .A1(n2013), .A2(n2014), .A3(n2015), .ZN(n2010) );
NOR2_X1 U1636 ( .A1(n2016), .A2(n2017), .ZN(n2015) );
NOR2_X1 U1637 ( .A1(KEYINPUT61), .A2(n2018), .ZN(n2016) );
NOR2_X1 U1638 ( .A1(KEYINPUT61), .A2(n1989), .ZN(n2014) );
NAND2_X1 U1639 ( .A1(n2017), .A2(n2019), .ZN(n1989) );
AND2_X1 U1640 ( .A1(n2020), .A2(n2021), .ZN(n2017) );
OR2_X1 U1641 ( .A1(n1986), .A2(KEYINPUT54), .ZN(n2021) );
NAND2_X1 U1642 ( .A1(n1991), .A2(n2022), .ZN(n1986) );
NAND2_X1 U1643 ( .A1(n2023), .A2(n2024), .ZN(n2022) );
OR2_X1 U1644 ( .A1(n2024), .A2(n2023), .ZN(n1991) );
NAND3_X1 U1645 ( .A1(n2023), .A2(n2024), .A3(KEYINPUT54), .ZN(n2020) );
XOR2_X1 U1646 ( .A(KEYINPUT17), .B(n1948), .Z(n2013) );
AND2_X1 U1647 ( .A1(n2023), .A2(n1945), .ZN(n2009) );
INV_X1 U1648 ( .A(n1882), .ZN(n1945) );
XNOR2_X1 U1649 ( .A(n2025), .B(n2026), .ZN(n2023) );
XOR2_X1 U1650 ( .A(n2003), .B(n2002), .Z(n2026) );
NAND2_X1 U1651 ( .A1(n2027), .A2(n2028), .ZN(n2002) );
NAND2_X1 U1652 ( .A1(n1927), .A2(DATA_IN_2_), .ZN(n2028) );
NAND2_X1 U1653 ( .A1(RESTART), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2027) );
NAND2_X1 U1654 ( .A1(n2029), .A2(n2030), .ZN(n2003) );
XOR2_X1 U1655 ( .A(n2031), .B(KEYINPUT31), .Z(n2029) );
NAND2_X1 U1656 ( .A1(n2032), .A2(n2033), .ZN(n2031) );
NAND2_X1 U1657 ( .A1(KEYINPUT41), .A2(n2004), .ZN(n2025) );
NAND2_X1 U1658 ( .A1(n2034), .A2(n2035), .ZN(n2004) );
NAND2_X1 U1659 ( .A1(n1927), .A2(REG4_REG_2__SCAN_IN), .ZN(n2035) );
XOR2_X1 U1660 ( .A(KEYINPUT25), .B(n2036), .Z(n2034) );
NOR2_X1 U1661 ( .A1(n1692), .A2(n1889), .ZN(n2036) );
NAND2_X1 U1662 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1757), .ZN(n2007) );
NAND2_X1 U1663 ( .A1(n1835), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2006) );
NAND2_X1 U1664 ( .A1(n1841), .A2(REG4_REG_1__SCAN_IN), .ZN(n2005) );
NAND4_X1 U1665 ( .A1(n2037), .A2(n2038), .A3(n2039), .A4(n2040), .ZN(U281));
NOR3_X1 U1666 ( .A1(n2041), .A2(n2042), .A3(n2043), .ZN(n2040) );
NOR2_X1 U1667 ( .A1(n2044), .A2(n1882), .ZN(n2043) );
NAND4_X1 U1668 ( .A1(STATO_REG_1__SCAN_IN), .A2(n2045), .A3(n2046), .A4(U280), .ZN(n1882) );
NAND2_X1 U1669 ( .A1(n1927), .A2(n2047), .ZN(n2045) );
NAND3_X1 U1670 ( .A1(n2048), .A2(n2049), .A3(ENABLE), .ZN(n2047) );
INV_X1 U1671 ( .A(AVERAGE), .ZN(n2049) );
NOR2_X1 U1672 ( .A1(n1839), .A2(n2019), .ZN(n2042) );
INV_X1 U1673 ( .A(n1948), .ZN(n1839) );
NOR3_X1 U1674 ( .A1(n1658), .A2(n1757), .A3(n2046), .ZN(n1948) );
NAND3_X1 U1675 ( .A1(n2050), .A2(n2051), .A3(RESTART), .ZN(n2046) );
NAND2_X1 U1676 ( .A1(n2052), .A2(n1698), .ZN(n2051) );
INV_X1 U1677 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1698) );
NAND2_X1 U1678 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n2053), .ZN(n2052) );
OR2_X1 U1679 ( .A1(n2053), .A2(RMAX_REG_7__SCAN_IN), .ZN(n2050) );
NAND2_X1 U1680 ( .A1(n2054), .A2(n2055), .ZN(n2053) );
NAND2_X1 U1681 ( .A1(n2056), .A2(n1697), .ZN(n2055) );
INV_X1 U1682 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1697) );
NAND3_X1 U1683 ( .A1(n2057), .A2(n2058), .A3(RMAX_REG_6__SCAN_IN), .ZN(n2056) );
XOR2_X1 U1684 ( .A(n2059), .B(KEYINPUT22), .Z(n2054) );
NAND2_X1 U1685 ( .A1(n1728), .A2(n2060), .ZN(n2059) );
NAND2_X1 U1686 ( .A1(n2057), .A2(n2058), .ZN(n2060) );
NAND3_X1 U1687 ( .A1(n2061), .A2(n2062), .A3(n2063), .ZN(n2058) );
NAND2_X1 U1688 ( .A1(RMIN_REG_5__SCAN_IN), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2063) );
NAND3_X1 U1689 ( .A1(n2064), .A2(n2065), .A3(n2066), .ZN(n2062) );
NAND2_X1 U1690 ( .A1(n1714), .A2(n1695), .ZN(n2066) );
INV_X1 U1691 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1695) );
INV_X1 U1692 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1714) );
NAND3_X1 U1693 ( .A1(n2067), .A2(n2068), .A3(n2069), .ZN(n2065) );
NAND2_X1 U1694 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2069) );
NAND3_X1 U1695 ( .A1(n2070), .A2(n2071), .A3(n2072), .ZN(n2068) );
NAND2_X1 U1696 ( .A1(n1721), .A2(n1692), .ZN(n2072) );
INV_X1 U1697 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1692) );
INV_X1 U1698 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1721) );
NAND2_X1 U1699 ( .A1(n2073), .A2(n2074), .ZN(n2071) );
NAND2_X1 U1700 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2074) );
XOR2_X1 U1701 ( .A(n2075), .B(KEYINPUT12), .Z(n2073) );
NAND2_X1 U1702 ( .A1(RMIN_REG_1__SCAN_IN), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2075) );
NAND2_X1 U1703 ( .A1(n1724), .A2(n1689), .ZN(n2070) );
INV_X1 U1704 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1689) );
NAND2_X1 U1705 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2067) );
NAND2_X1 U1706 ( .A1(n1726), .A2(n1682), .ZN(n2064) );
INV_X1 U1707 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1682) );
INV_X1 U1708 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1726) );
NAND2_X1 U1709 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2061) );
NAND2_X1 U1710 ( .A1(n2076), .A2(n1674), .ZN(n2057) );
INV_X1 U1711 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1674) );
INV_X1 U1712 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n2076) );
INV_X1 U1713 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1728) );
XOR2_X1 U1714 ( .A(n2077), .B(KEYINPUT32), .Z(n2041) );
OR2_X1 U1715 ( .A1(n1985), .A2(n1848), .ZN(n2077) );
INV_X1 U1716 ( .A(n1853), .ZN(n1848) );
NOR4_X1 U1717 ( .A1(n1753), .A2(n2048), .A3(n2078), .A4(AVERAGE), .ZN(n1853));
XNOR2_X1 U1718 ( .A(KEYINPUT23), .B(n2079), .ZN(n2078) );
NAND2_X1 U1719 ( .A1(n2080), .A2(n2081), .ZN(n2048) );
OR2_X1 U1720 ( .A1(DATA_IN_7_), .A2(REG4_REG_7__SCAN_IN), .ZN(n2081) );
NAND3_X1 U1721 ( .A1(n2082), .A2(n2083), .A3(n2084), .ZN(n2080) );
NAND2_X1 U1722 ( .A1(n1670), .A2(n1893), .ZN(n2084) );
INV_X1 U1723 ( .A(REG4_REG_6__SCAN_IN), .ZN(n1893) );
INV_X1 U1724 ( .A(DATA_IN_6_), .ZN(n1670) );
NAND2_X1 U1725 ( .A1(n2085), .A2(n2086), .ZN(n2083) );
NAND2_X1 U1726 ( .A1(REG4_REG_6__SCAN_IN), .A2(DATA_IN_6_), .ZN(n2086) );
NAND2_X1 U1727 ( .A1(n2087), .A2(n2088), .ZN(n2085) );
OR2_X1 U1728 ( .A1(DATA_IN_5_), .A2(REG4_REG_5__SCAN_IN), .ZN(n2088) );
NAND3_X1 U1729 ( .A1(n2089), .A2(n2090), .A3(n2091), .ZN(n2087) );
NAND2_X1 U1730 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2091) );
NAND3_X1 U1731 ( .A1(n2092), .A2(n2093), .A3(n2094), .ZN(n2090) );
OR2_X1 U1732 ( .A1(DATA_IN_4_), .A2(REG4_REG_4__SCAN_IN), .ZN(n2094) );
NAND3_X1 U1733 ( .A1(n2095), .A2(n2096), .A3(n2097), .ZN(n2093) );
NAND2_X1 U1734 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2097) );
NAND3_X1 U1735 ( .A1(n2098), .A2(n2099), .A3(n2100), .ZN(n2096) );
OR2_X1 U1736 ( .A1(DATA_IN_2_), .A2(REG4_REG_2__SCAN_IN), .ZN(n2100) );
NAND2_X1 U1737 ( .A1(n2101), .A2(n2102), .ZN(n2099) );
INV_X1 U1738 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2102) );
OR2_X1 U1739 ( .A1(n2103), .A2(n1691), .ZN(n2101) );
NAND2_X1 U1740 ( .A1(n2103), .A2(n1691), .ZN(n2098) );
INV_X1 U1741 ( .A(DATA_IN_1_), .ZN(n1691) );
NAND2_X1 U1742 ( .A1(n2104), .A2(DATA_IN_0_), .ZN(n2103) );
XNOR2_X1 U1743 ( .A(REG4_REG_0__SCAN_IN), .B(KEYINPUT24), .ZN(n2104) );
NAND2_X1 U1744 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2095) );
NAND2_X1 U1745 ( .A1(n1693), .A2(n1942), .ZN(n2092) );
INV_X1 U1746 ( .A(REG4_REG_3__SCAN_IN), .ZN(n1942) );
INV_X1 U1747 ( .A(DATA_IN_3_), .ZN(n1693) );
NAND2_X1 U1748 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2089) );
NAND2_X1 U1749 ( .A1(n2105), .A2(DATA_IN_7_), .ZN(n2082) );
XNOR2_X1 U1750 ( .A(REG4_REG_7__SCAN_IN), .B(KEYINPUT8), .ZN(n2105) );
NAND2_X1 U1751 ( .A1(n2106), .A2(n2107), .ZN(n1985) );
OR2_X1 U1752 ( .A1(n2018), .A2(KEYINPUT18), .ZN(n2107) );
INV_X1 U1753 ( .A(n2019), .ZN(n2018) );
NAND2_X1 U1754 ( .A1(n2024), .A2(n2108), .ZN(n2019) );
NAND2_X1 U1755 ( .A1(n2109), .A2(n2110), .ZN(n2108) );
OR2_X1 U1756 ( .A1(n2110), .A2(n2109), .ZN(n2024) );
NAND3_X1 U1757 ( .A1(n2109), .A2(n2044), .A3(KEYINPUT18), .ZN(n2106) );
INV_X1 U1758 ( .A(n2110), .ZN(n2044) );
NAND2_X1 U1759 ( .A1(n2111), .A2(n2112), .ZN(n2110) );
NAND2_X1 U1760 ( .A1(n2113), .A2(n2032), .ZN(n2112) );
NAND2_X1 U1761 ( .A1(n2030), .A2(n2033), .ZN(n2113) );
OR2_X1 U1762 ( .A1(n2114), .A2(n2115), .ZN(n2033) );
NAND2_X1 U1763 ( .A1(n2116), .A2(n2114), .ZN(n2030) );
XOR2_X1 U1764 ( .A(n2117), .B(KEYINPUT59), .Z(n2116) );
NAND2_X1 U1765 ( .A1(n2118), .A2(n2119), .ZN(n2111) );
XOR2_X1 U1766 ( .A(n2114), .B(n2115), .Z(n2119) );
INV_X1 U1767 ( .A(n2117), .ZN(n2115) );
NAND2_X1 U1768 ( .A1(n2120), .A2(n2121), .ZN(n2114) );
NAND2_X1 U1769 ( .A1(n1927), .A2(DATA_IN_1_), .ZN(n2121) );
XOR2_X1 U1770 ( .A(KEYINPUT46), .B(n2122), .Z(n2120) );
NOR2_X1 U1771 ( .A1(n2123), .A2(n1889), .ZN(n2122) );
XOR2_X1 U1772 ( .A(n1724), .B(KEYINPUT29), .Z(n2123) );
INV_X1 U1773 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1724) );
INV_X1 U1774 ( .A(n2032), .ZN(n2118) );
NAND2_X1 U1775 ( .A1(n2124), .A2(n2125), .ZN(n2032) );
NAND2_X1 U1776 ( .A1(n1927), .A2(REG4_REG_1__SCAN_IN), .ZN(n2125) );
NAND2_X1 U1777 ( .A1(RESTART), .A2(RMIN_REG_1__SCAN_IN), .ZN(n2124) );
AND3_X1 U1778 ( .A1(n2126), .A2(n2127), .A3(n2117), .ZN(n2109) );
NAND2_X1 U1779 ( .A1(n2128), .A2(n2129), .ZN(n2117) );
NAND2_X1 U1780 ( .A1(n2130), .A2(n2131), .ZN(n2129) );
OR2_X1 U1781 ( .A1(n2132), .A2(KEYINPUT26), .ZN(n2127) );
NAND4_X1 U1782 ( .A1(n2130), .A2(n2131), .A3(n2132), .A4(KEYINPUT26), .ZN(n2126) );
INV_X1 U1783 ( .A(n2128), .ZN(n2132) );
NAND2_X1 U1784 ( .A1(n2133), .A2(n2134), .ZN(n2128) );
NAND2_X1 U1785 ( .A1(n2135), .A2(RMIN_REG_0__SCAN_IN), .ZN(n2134) );
XOR2_X1 U1786 ( .A(n1889), .B(KEYINPUT49), .Z(n2135) );
NAND2_X1 U1787 ( .A1(n1927), .A2(REG4_REG_0__SCAN_IN), .ZN(n2133) );
NAND2_X1 U1788 ( .A1(n2136), .A2(DATA_IN_0_), .ZN(n2131) );
XOR2_X1 U1789 ( .A(n1927), .B(KEYINPUT50), .Z(n2136) );
NAND2_X1 U1790 ( .A1(RESTART), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2130) );
NAND2_X1 U1791 ( .A1(n2137), .A2(RLAST_REG_0__SCAN_IN), .ZN(n2039) );
XNOR2_X1 U1792 ( .A(n1835), .B(KEYINPUT40), .ZN(n2137) );
AND2_X1 U1793 ( .A1(n2079), .A2(n1753), .ZN(n1835) );
INV_X1 U1794 ( .A(ENABLE), .ZN(n1753) );
NAND2_X1 U1795 ( .A1(n1841), .A2(n2138), .ZN(n2038) );
XOR2_X1 U1796 ( .A(REG4_REG_0__SCAN_IN), .B(KEYINPUT27), .Z(n2138) );
INV_X1 U1797 ( .A(n1943), .ZN(n1841) );
NAND3_X1 U1798 ( .A1(ENABLE), .A2(n2079), .A3(AVERAGE), .ZN(n1943) );
NOR3_X1 U1799 ( .A1(n1658), .A2(n1757), .A3(n1890), .ZN(n2079) );
INV_X1 U1800 ( .A(n1927), .ZN(n1890) );
INV_X1 U1801 ( .A(RESTART), .ZN(n1889) );
NAND2_X1 U1802 ( .A1(n2139), .A2(n1757), .ZN(n2037) );
XOR2_X1 U1803 ( .A(KEYINPUT55), .B(DATA_OUT_REG_0__SCAN_IN), .Z(n2139) );
NAND2_X1 U1804 ( .A1(n1830), .A2(n2140), .ZN(U280) );
NAND2_X1 U1805 ( .A1(STATO_REG_0__SCAN_IN), .A2(n1658), .ZN(n2140) );
INV_X1 U1806 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1658) );
NAND2_X1 U1807 ( .A1(n1634), .A2(STATO_REG_1__SCAN_IN), .ZN(n1830) );
XOR2_X1 U1808 ( .A(n1633), .B(KEYINPUT34), .Z(n1634) );
INV_X1 U1809 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1633) );
endmodule


