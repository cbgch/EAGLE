//Key = 1110110000011101010101011110000100101110111001010000111010100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310;

XNOR2_X1 U729 ( .A(G107), .B(n1008), .ZN(G9) );
NOR2_X1 U730 ( .A1(n1009), .A2(n1010), .ZN(G75) );
NOR4_X1 U731 ( .A1(G953), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1010) );
NOR2_X1 U732 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR2_X1 U733 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR3_X1 U734 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1017) );
NOR2_X1 U735 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
AND2_X1 U736 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR3_X1 U737 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1021) );
NOR3_X1 U738 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
NOR2_X1 U739 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U740 ( .A1(n1024), .A2(n1033), .ZN(n1026) );
NOR4_X1 U741 ( .A1(n1034), .A2(n1035), .A3(n1025), .A4(n1028), .ZN(n1016) );
NOR3_X1 U742 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NOR2_X1 U743 ( .A1(n1039), .A2(n1018), .ZN(n1038) );
NOR2_X1 U744 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U745 ( .A1(KEYINPUT6), .A2(n1042), .ZN(n1041) );
NOR2_X1 U746 ( .A1(n1043), .A2(n1020), .ZN(n1037) );
NOR2_X1 U747 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
XOR2_X1 U748 ( .A(KEYINPUT23), .B(n1046), .Z(n1045) );
NOR2_X1 U749 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
AND3_X1 U750 ( .A1(KEYINPUT0), .A2(n1049), .A3(n1050), .ZN(n1048) );
NOR2_X1 U751 ( .A1(KEYINPUT0), .A2(n1018), .ZN(n1047) );
NOR2_X1 U752 ( .A1(n1024), .A2(n1051), .ZN(n1034) );
AND3_X1 U753 ( .A1(KEYINPUT6), .A2(n1052), .A3(n1053), .ZN(n1051) );
NOR3_X1 U754 ( .A1(n1011), .A2(G953), .A3(G952), .ZN(n1009) );
AND4_X1 U755 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1011) );
NOR4_X1 U756 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1057) );
XNOR2_X1 U757 ( .A(G469), .B(n1062), .ZN(n1061) );
XOR2_X1 U758 ( .A(KEYINPUT46), .B(n1025), .Z(n1060) );
XNOR2_X1 U759 ( .A(n1063), .B(n1064), .ZN(n1059) );
NAND2_X1 U760 ( .A1(KEYINPUT41), .A2(G478), .ZN(n1064) );
NOR3_X1 U761 ( .A1(n1065), .A2(n1066), .A3(n1050), .ZN(n1056) );
NAND2_X1 U762 ( .A1(G475), .A2(n1067), .ZN(n1055) );
XOR2_X1 U763 ( .A(n1068), .B(n1069), .Z(n1054) );
XOR2_X1 U764 ( .A(n1070), .B(KEYINPUT57), .Z(n1069) );
NAND2_X1 U765 ( .A1(KEYINPUT21), .A2(n1071), .ZN(n1068) );
XOR2_X1 U766 ( .A(n1072), .B(n1073), .Z(G72) );
XOR2_X1 U767 ( .A(n1074), .B(n1075), .Z(n1073) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
AND2_X1 U769 ( .A1(G227), .A2(G900), .ZN(n1076) );
NAND2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1074) );
NAND2_X1 U771 ( .A1(G953), .A2(n1080), .ZN(n1079) );
XOR2_X1 U772 ( .A(n1081), .B(n1082), .Z(n1078) );
XOR2_X1 U773 ( .A(KEYINPUT27), .B(n1083), .Z(n1082) );
XOR2_X1 U774 ( .A(n1084), .B(n1085), .Z(n1081) );
NAND2_X1 U775 ( .A1(n1077), .A2(n1086), .ZN(n1072) );
XOR2_X1 U776 ( .A(n1087), .B(n1088), .Z(G69) );
XOR2_X1 U777 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U778 ( .A1(n1091), .A2(n1077), .ZN(n1090) );
AND2_X1 U779 ( .A1(G224), .A2(G898), .ZN(n1091) );
NAND2_X1 U780 ( .A1(n1092), .A2(n1093), .ZN(n1089) );
NAND2_X1 U781 ( .A1(G953), .A2(n1094), .ZN(n1093) );
XOR2_X1 U782 ( .A(n1095), .B(n1096), .Z(n1092) );
XNOR2_X1 U783 ( .A(n1097), .B(n1098), .ZN(n1096) );
NAND2_X1 U784 ( .A1(KEYINPUT56), .A2(n1099), .ZN(n1097) );
XOR2_X1 U785 ( .A(n1100), .B(n1101), .Z(n1095) );
NAND2_X1 U786 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
XOR2_X1 U787 ( .A(KEYINPUT49), .B(KEYINPUT36), .Z(n1103) );
XNOR2_X1 U788 ( .A(n1104), .B(G101), .ZN(n1102) );
NAND2_X1 U789 ( .A1(n1077), .A2(n1105), .ZN(n1087) );
NAND2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR2_X1 U791 ( .A1(n1108), .A2(n1109), .ZN(G66) );
XOR2_X1 U792 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U793 ( .A1(KEYINPUT30), .A2(n1112), .ZN(n1111) );
NAND2_X1 U794 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
NOR2_X1 U795 ( .A1(n1108), .A2(n1115), .ZN(G63) );
NOR3_X1 U796 ( .A1(n1063), .A2(n1116), .A3(n1117), .ZN(n1115) );
AND3_X1 U797 ( .A1(n1118), .A2(G478), .A3(n1113), .ZN(n1117) );
NOR2_X1 U798 ( .A1(n1119), .A2(n1118), .ZN(n1116) );
AND2_X1 U799 ( .A1(n1013), .A2(G478), .ZN(n1119) );
NOR2_X1 U800 ( .A1(n1108), .A2(n1120), .ZN(G60) );
XOR2_X1 U801 ( .A(n1121), .B(n1122), .Z(n1120) );
AND2_X1 U802 ( .A1(G475), .A2(n1113), .ZN(n1122) );
XNOR2_X1 U803 ( .A(G104), .B(n1107), .ZN(G6) );
NOR2_X1 U804 ( .A1(n1108), .A2(n1123), .ZN(G57) );
XOR2_X1 U805 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U806 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U807 ( .A(n1128), .B(n1129), .Z(n1124) );
XOR2_X1 U808 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U809 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XNOR2_X1 U810 ( .A(G472), .B(KEYINPUT20), .ZN(n1132) );
NOR2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(n1130) );
XOR2_X1 U812 ( .A(KEYINPUT54), .B(KEYINPUT38), .Z(n1135) );
XOR2_X1 U813 ( .A(KEYINPUT26), .B(n1136), .Z(n1134) );
NAND2_X1 U814 ( .A1(KEYINPUT15), .A2(n1137), .ZN(n1128) );
INV_X1 U815 ( .A(n1138), .ZN(n1137) );
NOR2_X1 U816 ( .A1(n1108), .A2(n1139), .ZN(G54) );
XOR2_X1 U817 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U818 ( .A(n1142), .B(n1143), .ZN(n1141) );
NAND2_X1 U819 ( .A1(n1144), .A2(n1145), .ZN(n1142) );
NAND2_X1 U820 ( .A1(n1084), .A2(n1146), .ZN(n1145) );
NAND2_X1 U821 ( .A1(KEYINPUT2), .A2(n1147), .ZN(n1146) );
NAND2_X1 U822 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND2_X1 U823 ( .A1(n1150), .A2(n1151), .ZN(n1144) );
NAND2_X1 U824 ( .A1(n1149), .A2(n1152), .ZN(n1151) );
NAND2_X1 U825 ( .A1(KEYINPUT2), .A2(n1153), .ZN(n1152) );
INV_X1 U826 ( .A(KEYINPUT63), .ZN(n1149) );
INV_X1 U827 ( .A(n1148), .ZN(n1150) );
XOR2_X1 U828 ( .A(n1154), .B(n1155), .Z(n1140) );
XOR2_X1 U829 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U830 ( .A1(KEYINPUT12), .A2(n1158), .ZN(n1157) );
AND2_X1 U831 ( .A1(G469), .A2(n1113), .ZN(n1154) );
INV_X1 U832 ( .A(n1133), .ZN(n1113) );
NOR2_X1 U833 ( .A1(n1108), .A2(n1159), .ZN(G51) );
XOR2_X1 U834 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U835 ( .A(KEYINPUT10), .B(n1162), .Z(n1161) );
NOR2_X1 U836 ( .A1(n1163), .A2(n1133), .ZN(n1162) );
NAND2_X1 U837 ( .A1(G902), .A2(n1013), .ZN(n1133) );
NAND3_X1 U838 ( .A1(n1164), .A2(n1165), .A3(n1106), .ZN(n1013) );
AND4_X1 U839 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1106) );
AND4_X1 U840 ( .A1(n1008), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1169) );
NAND4_X1 U841 ( .A1(n1173), .A2(n1052), .A3(n1033), .A4(n1174), .ZN(n1008) );
XNOR2_X1 U842 ( .A(KEYINPUT61), .B(n1107), .ZN(n1165) );
NAND3_X1 U843 ( .A1(n1033), .A2(n1173), .A3(n1175), .ZN(n1107) );
INV_X1 U844 ( .A(n1086), .ZN(n1164) );
NAND4_X1 U845 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1086) );
AND3_X1 U846 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1179) );
NAND3_X1 U847 ( .A1(n1023), .A2(n1040), .A3(n1183), .ZN(n1178) );
NAND3_X1 U848 ( .A1(n1028), .A2(n1184), .A3(n1025), .ZN(n1176) );
NAND2_X1 U849 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND3_X1 U850 ( .A1(n1187), .A2(n1188), .A3(n1044), .ZN(n1186) );
NAND2_X1 U851 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
OR3_X1 U852 ( .A1(n1191), .A2(KEYINPUT58), .A3(n1042), .ZN(n1189) );
NAND3_X1 U853 ( .A1(n1192), .A2(n1193), .A3(n1029), .ZN(n1187) );
NAND3_X1 U854 ( .A1(n1052), .A2(n1194), .A3(KEYINPUT58), .ZN(n1193) );
NAND2_X1 U855 ( .A1(n1040), .A2(n1195), .ZN(n1192) );
XOR2_X1 U856 ( .A(KEYINPUT19), .B(n1191), .Z(n1195) );
NAND2_X1 U857 ( .A1(n1183), .A2(n1196), .ZN(n1185) );
XNOR2_X1 U858 ( .A(G210), .B(KEYINPUT33), .ZN(n1163) );
XOR2_X1 U859 ( .A(n1197), .B(n1198), .Z(n1160) );
NOR2_X1 U860 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U861 ( .A(n1201), .B(KEYINPUT37), .Z(n1200) );
NAND2_X1 U862 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NOR2_X1 U863 ( .A1(n1204), .A2(G952), .ZN(n1108) );
XOR2_X1 U864 ( .A(KEYINPUT35), .B(n1077), .Z(n1204) );
XOR2_X1 U865 ( .A(n1205), .B(n1206), .Z(G48) );
NAND4_X1 U866 ( .A1(n1207), .A2(n1040), .A3(n1208), .A4(n1194), .ZN(n1206) );
XOR2_X1 U867 ( .A(KEYINPUT43), .B(n1044), .Z(n1208) );
XNOR2_X1 U868 ( .A(G143), .B(n1177), .ZN(G45) );
NAND3_X1 U869 ( .A1(n1209), .A2(n1023), .A3(n1210), .ZN(n1177) );
XNOR2_X1 U870 ( .A(G140), .B(n1180), .ZN(G42) );
NAND3_X1 U871 ( .A1(n1175), .A2(n1028), .A3(n1183), .ZN(n1180) );
XNOR2_X1 U872 ( .A(G137), .B(n1211), .ZN(G39) );
NAND4_X1 U873 ( .A1(n1025), .A2(n1028), .A3(n1044), .A4(n1212), .ZN(n1211) );
NOR3_X1 U874 ( .A1(n1213), .A2(n1020), .A3(n1036), .ZN(n1212) );
XOR2_X1 U875 ( .A(KEYINPUT60), .B(n1191), .Z(n1213) );
INV_X1 U876 ( .A(n1174), .ZN(n1025) );
XOR2_X1 U877 ( .A(n1182), .B(n1214), .Z(G36) );
XOR2_X1 U878 ( .A(KEYINPUT31), .B(G134), .Z(n1214) );
NAND3_X1 U879 ( .A1(n1023), .A2(n1052), .A3(n1183), .ZN(n1182) );
XNOR2_X1 U880 ( .A(G131), .B(n1215), .ZN(G33) );
NAND4_X1 U881 ( .A1(KEYINPUT13), .A2(n1183), .A3(n1023), .A4(n1040), .ZN(n1215) );
NOR2_X1 U882 ( .A1(n1036), .A2(n1216), .ZN(n1183) );
INV_X1 U883 ( .A(n1024), .ZN(n1036) );
NOR2_X1 U884 ( .A1(n1031), .A2(n1065), .ZN(n1024) );
INV_X1 U885 ( .A(n1032), .ZN(n1065) );
XOR2_X1 U886 ( .A(n1217), .B(n1218), .Z(G30) );
NOR2_X1 U887 ( .A1(KEYINPUT3), .A2(n1219), .ZN(n1218) );
AND3_X1 U888 ( .A1(n1210), .A2(n1052), .A3(n1207), .ZN(n1219) );
INV_X1 U889 ( .A(n1216), .ZN(n1210) );
NAND2_X1 U890 ( .A1(n1044), .A2(n1194), .ZN(n1216) );
XOR2_X1 U891 ( .A(n1168), .B(n1220), .Z(G3) );
NAND2_X1 U892 ( .A1(KEYINPUT34), .A2(G101), .ZN(n1220) );
NAND3_X1 U893 ( .A1(n1196), .A2(n1173), .A3(n1023), .ZN(n1168) );
XOR2_X1 U894 ( .A(n1203), .B(n1181), .Z(G27) );
NAND3_X1 U895 ( .A1(n1175), .A2(n1053), .A3(n1221), .ZN(n1181) );
NOR3_X1 U896 ( .A1(n1190), .A2(n1191), .A3(n1033), .ZN(n1221) );
INV_X1 U897 ( .A(n1194), .ZN(n1191) );
NAND2_X1 U898 ( .A1(n1015), .A2(n1222), .ZN(n1194) );
NAND4_X1 U899 ( .A1(G953), .A2(G902), .A3(n1223), .A4(n1080), .ZN(n1222) );
INV_X1 U900 ( .A(G900), .ZN(n1080) );
AND2_X1 U901 ( .A1(n1040), .A2(n1174), .ZN(n1175) );
XNOR2_X1 U902 ( .A(G122), .B(n1166), .ZN(G24) );
NAND4_X1 U903 ( .A1(n1209), .A2(n1224), .A3(n1033), .A4(n1174), .ZN(n1166) );
NOR3_X1 U904 ( .A1(n1190), .A2(n1225), .A3(n1226), .ZN(n1209) );
XNOR2_X1 U905 ( .A(G119), .B(n1167), .ZN(G21) );
NAND3_X1 U906 ( .A1(n1224), .A2(n1196), .A3(n1207), .ZN(n1167) );
NOR3_X1 U907 ( .A1(n1174), .A2(n1033), .A3(n1190), .ZN(n1207) );
XOR2_X1 U908 ( .A(n1172), .B(n1227), .Z(G18) );
NAND2_X1 U909 ( .A1(KEYINPUT11), .A2(G116), .ZN(n1227) );
NAND4_X1 U910 ( .A1(n1023), .A2(n1224), .A3(n1052), .A4(n1029), .ZN(n1172) );
INV_X1 U911 ( .A(n1042), .ZN(n1052) );
NAND2_X1 U912 ( .A1(n1225), .A2(n1228), .ZN(n1042) );
XNOR2_X1 U913 ( .A(G113), .B(n1171), .ZN(G15) );
NAND4_X1 U914 ( .A1(n1023), .A2(n1040), .A3(n1224), .A4(n1229), .ZN(n1171) );
AND2_X1 U915 ( .A1(n1053), .A2(n1230), .ZN(n1224) );
INV_X1 U916 ( .A(n1018), .ZN(n1053) );
NAND2_X1 U917 ( .A1(n1049), .A2(n1231), .ZN(n1018) );
NOR2_X1 U918 ( .A1(n1228), .A2(n1225), .ZN(n1040) );
NOR2_X1 U919 ( .A1(n1028), .A2(n1174), .ZN(n1023) );
XNOR2_X1 U920 ( .A(G110), .B(n1170), .ZN(G12) );
NAND4_X1 U921 ( .A1(n1196), .A2(n1173), .A3(n1174), .A4(n1028), .ZN(n1170) );
INV_X1 U922 ( .A(n1033), .ZN(n1028) );
XNOR2_X1 U923 ( .A(n1058), .B(KEYINPUT14), .ZN(n1033) );
XNOR2_X1 U924 ( .A(n1232), .B(n1114), .ZN(n1058) );
AND2_X1 U925 ( .A1(G217), .A2(n1233), .ZN(n1114) );
OR2_X1 U926 ( .A1(n1112), .A2(G902), .ZN(n1232) );
XOR2_X1 U927 ( .A(n1234), .B(n1235), .Z(n1112) );
XNOR2_X1 U928 ( .A(n1236), .B(n1237), .ZN(n1235) );
XOR2_X1 U929 ( .A(n1238), .B(n1239), .Z(n1237) );
NOR2_X1 U930 ( .A1(KEYINPUT44), .A2(n1085), .ZN(n1239) );
NAND2_X1 U931 ( .A1(n1240), .A2(G221), .ZN(n1238) );
XOR2_X1 U932 ( .A(n1241), .B(n1242), .Z(n1234) );
XOR2_X1 U933 ( .A(G128), .B(G110), .Z(n1242) );
XOR2_X1 U934 ( .A(G137), .B(n1205), .Z(n1241) );
XOR2_X1 U935 ( .A(n1243), .B(G472), .Z(n1174) );
NAND2_X1 U936 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XOR2_X1 U937 ( .A(n1246), .B(n1247), .Z(n1244) );
XOR2_X1 U938 ( .A(n1136), .B(n1248), .Z(n1247) );
XOR2_X1 U939 ( .A(n1126), .B(n1098), .Z(n1248) );
XOR2_X1 U940 ( .A(n1236), .B(KEYINPUT51), .Z(n1126) );
XOR2_X1 U941 ( .A(n1202), .B(n1083), .Z(n1136) );
XOR2_X1 U942 ( .A(n1249), .B(n1250), .Z(n1246) );
NOR2_X1 U943 ( .A1(KEYINPUT32), .A2(n1251), .ZN(n1250) );
NOR3_X1 U944 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1251) );
AND2_X1 U945 ( .A1(n1255), .A2(G101), .ZN(n1254) );
NOR3_X1 U946 ( .A1(G101), .A2(KEYINPUT8), .A3(n1255), .ZN(n1253) );
OR2_X1 U947 ( .A1(KEYINPUT39), .A2(n1138), .ZN(n1255) );
AND2_X1 U948 ( .A1(n1138), .A2(KEYINPUT8), .ZN(n1252) );
NAND2_X1 U949 ( .A1(n1256), .A2(G210), .ZN(n1138) );
XNOR2_X1 U950 ( .A(KEYINPUT55), .B(KEYINPUT17), .ZN(n1249) );
AND3_X1 U951 ( .A1(n1229), .A2(n1230), .A3(n1044), .ZN(n1173) );
NOR2_X1 U952 ( .A1(n1049), .A2(n1050), .ZN(n1044) );
INV_X1 U953 ( .A(n1231), .ZN(n1050) );
NAND2_X1 U954 ( .A1(G221), .A2(n1233), .ZN(n1231) );
NAND2_X1 U955 ( .A1(G234), .A2(n1245), .ZN(n1233) );
XNOR2_X1 U956 ( .A(n1062), .B(n1257), .ZN(n1049) );
NOR2_X1 U957 ( .A1(KEYINPUT16), .A2(n1258), .ZN(n1257) );
XNOR2_X1 U958 ( .A(G469), .B(KEYINPUT24), .ZN(n1258) );
NAND2_X1 U959 ( .A1(n1259), .A2(n1245), .ZN(n1062) );
XNOR2_X1 U960 ( .A(n1158), .B(n1260), .ZN(n1259) );
XNOR2_X1 U961 ( .A(n1261), .B(n1156), .ZN(n1260) );
NAND2_X1 U962 ( .A1(G227), .A2(n1077), .ZN(n1156) );
NAND2_X1 U963 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NAND2_X1 U964 ( .A1(n1264), .A2(n1143), .ZN(n1263) );
XOR2_X1 U965 ( .A(n1265), .B(KEYINPUT59), .Z(n1262) );
OR2_X1 U966 ( .A1(n1143), .A2(n1264), .ZN(n1265) );
XNOR2_X1 U967 ( .A(n1266), .B(n1153), .ZN(n1264) );
INV_X1 U968 ( .A(n1084), .ZN(n1153) );
XOR2_X1 U969 ( .A(n1267), .B(G128), .Z(n1084) );
NAND2_X1 U970 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND2_X1 U971 ( .A1(G143), .A2(n1205), .ZN(n1269) );
XOR2_X1 U972 ( .A(KEYINPUT42), .B(n1270), .Z(n1268) );
NOR2_X1 U973 ( .A1(G143), .A2(n1205), .ZN(n1270) );
INV_X1 U974 ( .A(G146), .ZN(n1205) );
NAND2_X1 U975 ( .A1(KEYINPUT47), .A2(n1148), .ZN(n1266) );
XNOR2_X1 U976 ( .A(G101), .B(n1271), .ZN(n1148) );
NOR2_X1 U977 ( .A1(KEYINPUT9), .A2(n1104), .ZN(n1271) );
XOR2_X1 U978 ( .A(n1083), .B(KEYINPUT52), .Z(n1143) );
XNOR2_X1 U979 ( .A(n1272), .B(n1273), .ZN(n1083) );
XOR2_X1 U980 ( .A(KEYINPUT53), .B(G137), .Z(n1273) );
XNOR2_X1 U981 ( .A(G131), .B(G134), .ZN(n1272) );
XOR2_X1 U982 ( .A(G140), .B(G110), .Z(n1158) );
NAND2_X1 U983 ( .A1(n1274), .A2(n1015), .ZN(n1230) );
NAND3_X1 U984 ( .A1(n1223), .A2(n1077), .A3(G952), .ZN(n1015) );
XOR2_X1 U985 ( .A(KEYINPUT1), .B(n1275), .Z(n1274) );
AND4_X1 U986 ( .A1(n1094), .A2(n1223), .A3(G902), .A4(G953), .ZN(n1275) );
NAND2_X1 U987 ( .A1(G237), .A2(G234), .ZN(n1223) );
INV_X1 U988 ( .A(G898), .ZN(n1094) );
XOR2_X1 U989 ( .A(n1029), .B(KEYINPUT28), .Z(n1229) );
INV_X1 U990 ( .A(n1190), .ZN(n1029) );
NAND2_X1 U991 ( .A1(n1031), .A2(n1032), .ZN(n1190) );
NAND2_X1 U992 ( .A1(G214), .A2(n1276), .ZN(n1032) );
XNOR2_X1 U993 ( .A(n1277), .B(n1070), .ZN(n1031) );
NAND2_X1 U994 ( .A1(n1278), .A2(n1245), .ZN(n1070) );
XOR2_X1 U995 ( .A(n1279), .B(n1280), .Z(n1278) );
INV_X1 U996 ( .A(n1197), .ZN(n1280) );
XOR2_X1 U997 ( .A(n1281), .B(n1282), .Z(n1197) );
XNOR2_X1 U998 ( .A(n1104), .B(n1283), .ZN(n1282) );
XOR2_X1 U999 ( .A(n1284), .B(n1101), .Z(n1283) );
NOR2_X1 U1000 ( .A1(KEYINPUT50), .A2(n1236), .ZN(n1101) );
XOR2_X1 U1001 ( .A(G119), .B(KEYINPUT4), .Z(n1236) );
NAND2_X1 U1002 ( .A1(G224), .A2(n1077), .ZN(n1284) );
XOR2_X1 U1003 ( .A(G107), .B(n1285), .Z(n1104) );
INV_X1 U1004 ( .A(n1286), .ZN(n1285) );
XNOR2_X1 U1005 ( .A(n1127), .B(n1099), .ZN(n1281) );
XOR2_X1 U1006 ( .A(G110), .B(n1287), .Z(n1099) );
XOR2_X1 U1007 ( .A(KEYINPUT18), .B(G122), .Z(n1287) );
XOR2_X1 U1008 ( .A(G101), .B(n1098), .Z(n1127) );
XOR2_X1 U1009 ( .A(G113), .B(G116), .Z(n1098) );
NOR2_X1 U1010 ( .A1(n1199), .A2(n1288), .ZN(n1279) );
XOR2_X1 U1011 ( .A(n1289), .B(KEYINPUT5), .Z(n1288) );
NAND2_X1 U1012 ( .A1(n1290), .A2(n1203), .ZN(n1289) );
XNOR2_X1 U1013 ( .A(n1202), .B(KEYINPUT45), .ZN(n1290) );
NOR2_X1 U1014 ( .A1(n1203), .A2(n1202), .ZN(n1199) );
XNOR2_X1 U1015 ( .A(n1217), .B(n1291), .ZN(n1202) );
INV_X1 U1016 ( .A(G128), .ZN(n1217) );
INV_X1 U1017 ( .A(G125), .ZN(n1203) );
NAND2_X1 U1018 ( .A1(KEYINPUT40), .A2(n1071), .ZN(n1277) );
NAND2_X1 U1019 ( .A1(G210), .A2(n1276), .ZN(n1071) );
OR2_X1 U1020 ( .A1(G902), .A2(G237), .ZN(n1276) );
INV_X1 U1021 ( .A(n1020), .ZN(n1196) );
NAND2_X1 U1022 ( .A1(n1225), .A2(n1226), .ZN(n1020) );
INV_X1 U1023 ( .A(n1228), .ZN(n1226) );
XNOR2_X1 U1024 ( .A(n1063), .B(n1292), .ZN(n1228) );
NOR2_X1 U1025 ( .A1(G478), .A2(KEYINPUT48), .ZN(n1292) );
NOR2_X1 U1026 ( .A1(n1118), .A2(G902), .ZN(n1063) );
XNOR2_X1 U1027 ( .A(n1293), .B(n1294), .ZN(n1118) );
XOR2_X1 U1028 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U1029 ( .A(G107), .B(n1297), .ZN(n1296) );
NOR2_X1 U1030 ( .A1(G134), .A2(KEYINPUT22), .ZN(n1297) );
NAND2_X1 U1031 ( .A1(G217), .A2(n1240), .ZN(n1295) );
AND2_X1 U1032 ( .A1(G234), .A2(n1077), .ZN(n1240) );
INV_X1 U1033 ( .A(G953), .ZN(n1077) );
XOR2_X1 U1034 ( .A(n1298), .B(n1299), .Z(n1293) );
XOR2_X1 U1035 ( .A(G143), .B(G128), .Z(n1299) );
XNOR2_X1 U1036 ( .A(G116), .B(G122), .ZN(n1298) );
NOR2_X1 U1037 ( .A1(n1300), .A2(n1066), .ZN(n1225) );
NOR3_X1 U1038 ( .A1(G475), .A2(G902), .A3(n1121), .ZN(n1066) );
AND2_X1 U1039 ( .A1(n1301), .A2(n1067), .ZN(n1300) );
NAND2_X1 U1040 ( .A1(n1302), .A2(n1245), .ZN(n1067) );
INV_X1 U1041 ( .A(G902), .ZN(n1245) );
INV_X1 U1042 ( .A(n1121), .ZN(n1302) );
XOR2_X1 U1043 ( .A(n1303), .B(n1304), .Z(n1121) );
XOR2_X1 U1044 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U1045 ( .A(n1307), .B(n1308), .Z(n1306) );
NOR2_X1 U1046 ( .A1(KEYINPUT7), .A2(n1309), .ZN(n1308) );
XNOR2_X1 U1047 ( .A(G113), .B(G122), .ZN(n1309) );
NAND2_X1 U1048 ( .A1(n1256), .A2(G214), .ZN(n1307) );
NOR2_X1 U1049 ( .A1(G953), .A2(G237), .ZN(n1256) );
XNOR2_X1 U1050 ( .A(G131), .B(KEYINPUT62), .ZN(n1305) );
XOR2_X1 U1051 ( .A(n1286), .B(n1310), .Z(n1303) );
XOR2_X1 U1052 ( .A(n1291), .B(n1085), .Z(n1310) );
XOR2_X1 U1053 ( .A(G140), .B(G125), .Z(n1085) );
XOR2_X1 U1054 ( .A(G143), .B(G146), .Z(n1291) );
XNOR2_X1 U1055 ( .A(G104), .B(KEYINPUT25), .ZN(n1286) );
XOR2_X1 U1056 ( .A(KEYINPUT29), .B(G475), .Z(n1301) );
endmodule


