//Key = 0100011000010000101101001101010111010111100110000010110101110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310;

XOR2_X1 U720 ( .A(G107), .B(n987), .Z(G9) );
NOR2_X1 U721 ( .A1(n988), .A2(n989), .ZN(G75) );
XOR2_X1 U722 ( .A(KEYINPUT0), .B(n990), .Z(n989) );
NOR3_X1 U723 ( .A1(n991), .A2(n992), .A3(n993), .ZN(n990) );
NOR3_X1 U724 ( .A1(n994), .A2(n995), .A3(n996), .ZN(n992) );
NOR2_X1 U725 ( .A1(n997), .A2(n998), .ZN(n995) );
NOR2_X1 U726 ( .A1(n999), .A2(n1000), .ZN(n998) );
NOR2_X1 U727 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NOR2_X1 U728 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NOR3_X1 U729 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n1001) );
XNOR2_X1 U730 ( .A(KEYINPUT19), .B(n1004), .ZN(n1005) );
NOR3_X1 U731 ( .A1(n1004), .A2(n1008), .A3(n1009), .ZN(n997) );
NAND3_X1 U732 ( .A1(n1010), .A2(n1011), .A3(n1012), .ZN(n991) );
NAND4_X1 U733 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
NOR3_X1 U734 ( .A1(n1009), .A2(n1017), .A3(n1000), .ZN(n1016) );
NOR2_X1 U735 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
INV_X1 U736 ( .A(n1020), .ZN(n1009) );
INV_X1 U737 ( .A(n1004), .ZN(n1015) );
NAND2_X1 U738 ( .A1(KEYINPUT38), .A2(n1021), .ZN(n1004) );
NAND4_X1 U739 ( .A1(n1022), .A2(n1023), .A3(n1019), .A4(n1024), .ZN(n1014) );
NAND2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(n1022) );
NAND2_X1 U741 ( .A1(n996), .A2(n994), .ZN(n1013) );
INV_X1 U742 ( .A(n1027), .ZN(n994) );
NOR3_X1 U743 ( .A1(n1028), .A2(G953), .A3(G952), .ZN(n988) );
INV_X1 U744 ( .A(n1010), .ZN(n1028) );
NAND4_X1 U745 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1010) );
NOR4_X1 U746 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1032) );
XOR2_X1 U747 ( .A(n1037), .B(n1038), .Z(n1036) );
NOR2_X1 U748 ( .A1(KEYINPUT34), .A2(n1039), .ZN(n1038) );
XOR2_X1 U749 ( .A(KEYINPUT28), .B(n1040), .Z(n1035) );
XOR2_X1 U750 ( .A(KEYINPUT62), .B(n1041), .Z(n1034) );
NOR3_X1 U751 ( .A1(n1042), .A2(n1025), .A3(n1043), .ZN(n1031) );
XNOR2_X1 U752 ( .A(n1044), .B(n1045), .ZN(n1030) );
XNOR2_X1 U753 ( .A(G475), .B(KEYINPUT39), .ZN(n1045) );
XOR2_X1 U754 ( .A(n1046), .B(n1047), .Z(n1029) );
NAND2_X1 U755 ( .A1(KEYINPUT5), .A2(n1048), .ZN(n1047) );
XOR2_X1 U756 ( .A(n1049), .B(n1050), .Z(G72) );
NAND2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U758 ( .A1(G900), .A2(G227), .ZN(n1052) );
NAND2_X1 U759 ( .A1(KEYINPUT6), .A2(n1053), .ZN(n1049) );
XOR2_X1 U760 ( .A(n1054), .B(n1055), .Z(n1053) );
NAND2_X1 U761 ( .A1(n1011), .A2(n1056), .ZN(n1055) );
NAND2_X1 U762 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U763 ( .A1(n1059), .A2(n1060), .ZN(n1054) );
INV_X1 U764 ( .A(n1061), .ZN(n1060) );
XNOR2_X1 U765 ( .A(n1062), .B(n1063), .ZN(n1059) );
NAND3_X1 U766 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1062) );
NAND2_X1 U767 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U768 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
INV_X1 U769 ( .A(KEYINPUT43), .ZN(n1070) );
NAND2_X1 U770 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
XNOR2_X1 U771 ( .A(KEYINPUT7), .B(n1067), .ZN(n1072) );
INV_X1 U772 ( .A(n1068), .ZN(n1071) );
NAND2_X1 U773 ( .A1(KEYINPUT43), .A2(n1073), .ZN(n1064) );
NAND2_X1 U774 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U775 ( .A1(KEYINPUT7), .A2(n1067), .ZN(n1075) );
OR3_X1 U776 ( .A1(n1068), .A2(KEYINPUT7), .A3(n1067), .ZN(n1074) );
XNOR2_X1 U777 ( .A(G131), .B(n1076), .ZN(n1067) );
NOR2_X1 U778 ( .A1(KEYINPUT51), .A2(n1077), .ZN(n1076) );
XNOR2_X1 U779 ( .A(n1078), .B(KEYINPUT48), .ZN(n1068) );
XOR2_X1 U780 ( .A(n1079), .B(n1080), .Z(G69) );
XOR2_X1 U781 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND2_X1 U782 ( .A1(n1051), .A2(n1083), .ZN(n1082) );
NAND2_X1 U783 ( .A1(G898), .A2(G224), .ZN(n1083) );
XNOR2_X1 U784 ( .A(G953), .B(KEYINPUT44), .ZN(n1051) );
NAND2_X1 U785 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
XOR2_X1 U786 ( .A(n1086), .B(n1087), .Z(n1084) );
XOR2_X1 U787 ( .A(KEYINPUT29), .B(n1088), .Z(n1087) );
NOR2_X1 U788 ( .A1(n1089), .A2(G953), .ZN(n1079) );
NOR2_X1 U789 ( .A1(n1090), .A2(n1091), .ZN(G66) );
NOR3_X1 U790 ( .A1(n1037), .A2(n1092), .A3(n1093), .ZN(n1091) );
NOR4_X1 U791 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1093) );
INV_X1 U792 ( .A(n1098), .ZN(n1094) );
NOR2_X1 U793 ( .A1(n1099), .A2(n1098), .ZN(n1092) );
NOR3_X1 U794 ( .A1(n1095), .A2(n1100), .A3(n1096), .ZN(n1099) );
INV_X1 U795 ( .A(G217), .ZN(n1096) );
INV_X1 U796 ( .A(KEYINPUT52), .ZN(n1095) );
NOR2_X1 U797 ( .A1(n1090), .A2(n1101), .ZN(G63) );
NOR2_X1 U798 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U799 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U800 ( .A1(KEYINPUT41), .A2(n1106), .ZN(n1105) );
NOR2_X1 U801 ( .A1(n1107), .A2(n1097), .ZN(n1104) );
AND2_X1 U802 ( .A1(n1106), .A2(KEYINPUT41), .ZN(n1102) );
NOR2_X1 U803 ( .A1(n1090), .A2(n1108), .ZN(G60) );
NOR3_X1 U804 ( .A1(n1044), .A2(n1109), .A3(n1110), .ZN(n1108) );
NOR2_X1 U805 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U806 ( .A1(n1100), .A2(n1113), .ZN(n1111) );
INV_X1 U807 ( .A(n993), .ZN(n1100) );
NOR3_X1 U808 ( .A1(n1114), .A2(n1113), .A3(n1097), .ZN(n1109) );
INV_X1 U809 ( .A(n1112), .ZN(n1114) );
NAND2_X1 U810 ( .A1(n1115), .A2(n1116), .ZN(G6) );
NAND2_X1 U811 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
INV_X1 U812 ( .A(G104), .ZN(n1118) );
NAND2_X1 U813 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NAND2_X1 U814 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
OR2_X1 U815 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
INV_X1 U816 ( .A(KEYINPUT40), .ZN(n1122) );
NAND2_X1 U817 ( .A1(G104), .A2(n1123), .ZN(n1115) );
NOR2_X1 U818 ( .A1(n1124), .A2(KEYINPUT23), .ZN(n1123) );
INV_X1 U819 ( .A(n1121), .ZN(n1124) );
NOR2_X1 U820 ( .A1(n1090), .A2(n1125), .ZN(G57) );
XOR2_X1 U821 ( .A(n1126), .B(n1127), .Z(n1125) );
XNOR2_X1 U822 ( .A(n1128), .B(n1129), .ZN(n1127) );
NOR2_X1 U823 ( .A1(KEYINPUT49), .A2(n1130), .ZN(n1129) );
XNOR2_X1 U824 ( .A(n1131), .B(n1132), .ZN(n1126) );
NOR2_X1 U825 ( .A1(n1133), .A2(n1097), .ZN(n1132) );
NOR2_X1 U826 ( .A1(n1090), .A2(n1134), .ZN(G54) );
XOR2_X1 U827 ( .A(n1135), .B(n1136), .Z(n1134) );
XNOR2_X1 U828 ( .A(n1137), .B(n1078), .ZN(n1136) );
XNOR2_X1 U829 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR2_X1 U830 ( .A1(KEYINPUT20), .A2(n1140), .ZN(n1139) );
XOR2_X1 U831 ( .A(n1141), .B(n1142), .Z(n1135) );
NOR2_X1 U832 ( .A1(n1048), .A2(n1097), .ZN(n1142) );
XNOR2_X1 U833 ( .A(G110), .B(n1143), .ZN(n1141) );
NOR2_X1 U834 ( .A1(n1090), .A2(n1144), .ZN(G51) );
XOR2_X1 U835 ( .A(n1145), .B(n1146), .Z(n1144) );
XNOR2_X1 U836 ( .A(n1147), .B(n1148), .ZN(n1146) );
NOR3_X1 U837 ( .A1(n1097), .A2(KEYINPUT10), .A3(n1149), .ZN(n1148) );
INV_X1 U838 ( .A(G210), .ZN(n1149) );
NAND2_X1 U839 ( .A1(G902), .A2(n993), .ZN(n1097) );
NAND3_X1 U840 ( .A1(n1057), .A2(n1150), .A3(n1089), .ZN(n993) );
AND4_X1 U841 ( .A1(n1121), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1089) );
NOR4_X1 U842 ( .A1(n1154), .A2(n1155), .A3(n987), .A4(n1156), .ZN(n1153) );
INV_X1 U843 ( .A(n1157), .ZN(n1156) );
AND4_X1 U844 ( .A1(n1158), .A2(n1159), .A3(n1019), .A4(n1160), .ZN(n987) );
NAND2_X1 U845 ( .A1(n1161), .A2(n1162), .ZN(n1152) );
INV_X1 U846 ( .A(n1008), .ZN(n1162) );
NOR2_X1 U847 ( .A1(n1163), .A2(n1159), .ZN(n1008) );
NAND2_X1 U848 ( .A1(n1164), .A2(n1160), .ZN(n1121) );
XNOR2_X1 U849 ( .A(KEYINPUT58), .B(n1058), .ZN(n1150) );
AND4_X1 U850 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1057) );
NOR4_X1 U851 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1168) );
XOR2_X1 U852 ( .A(n1173), .B(n1174), .Z(n1145) );
XNOR2_X1 U853 ( .A(G125), .B(n1175), .ZN(n1174) );
NAND2_X1 U854 ( .A1(n1176), .A2(KEYINPUT16), .ZN(n1173) );
XNOR2_X1 U855 ( .A(n1177), .B(KEYINPUT30), .ZN(n1176) );
NOR2_X1 U856 ( .A1(n1011), .A2(G952), .ZN(n1090) );
XNOR2_X1 U857 ( .A(n1178), .B(n1169), .ZN(G48) );
AND3_X1 U858 ( .A1(n1163), .A2(n1179), .A3(n1180), .ZN(n1169) );
XNOR2_X1 U859 ( .A(G143), .B(n1167), .ZN(G45) );
NAND4_X1 U860 ( .A1(n1181), .A2(n1182), .A3(n1179), .A4(n1183), .ZN(n1167) );
XOR2_X1 U861 ( .A(n1165), .B(n1184), .Z(G42) );
XNOR2_X1 U862 ( .A(G140), .B(KEYINPUT56), .ZN(n1184) );
NAND4_X1 U863 ( .A1(n1020), .A2(n1164), .A3(n996), .A4(n1185), .ZN(n1165) );
NOR3_X1 U864 ( .A1(n1033), .A2(n1023), .A3(n1186), .ZN(n1164) );
INV_X1 U865 ( .A(n1163), .ZN(n1186) );
XNOR2_X1 U866 ( .A(G137), .B(n1166), .ZN(G39) );
NAND3_X1 U867 ( .A1(n1180), .A2(n1187), .A3(n1020), .ZN(n1166) );
XOR2_X1 U868 ( .A(G134), .B(n1172), .Z(G36) );
AND3_X1 U869 ( .A1(n1182), .A2(n1159), .A3(n1020), .ZN(n1172) );
XOR2_X1 U870 ( .A(G131), .B(n1171), .Z(G33) );
AND3_X1 U871 ( .A1(n1182), .A2(n1163), .A3(n1020), .ZN(n1171) );
NOR2_X1 U872 ( .A1(n1007), .A2(n1043), .ZN(n1020) );
NOR4_X1 U873 ( .A1(n1023), .A2(n1019), .A3(n996), .A4(n1188), .ZN(n1182) );
XNOR2_X1 U874 ( .A(n1058), .B(n1189), .ZN(G30) );
NOR2_X1 U875 ( .A1(KEYINPUT13), .A2(n1190), .ZN(n1189) );
NAND3_X1 U876 ( .A1(n1159), .A2(n1179), .A3(n1180), .ZN(n1058) );
NOR4_X1 U877 ( .A1(n1024), .A2(n1023), .A3(n1019), .A4(n1188), .ZN(n1180) );
INV_X1 U878 ( .A(n1158), .ZN(n1023) );
XNOR2_X1 U879 ( .A(n1128), .B(n1191), .ZN(G3) );
NOR2_X1 U880 ( .A1(KEYINPUT42), .A2(n1151), .ZN(n1191) );
NAND4_X1 U881 ( .A1(n1187), .A2(n1158), .A3(n1160), .A4(n1033), .ZN(n1151) );
XOR2_X1 U882 ( .A(G125), .B(n1170), .Z(G27) );
AND4_X1 U883 ( .A1(n1163), .A2(n1027), .A3(n1192), .A4(n996), .ZN(n1170) );
NOR2_X1 U884 ( .A1(n1188), .A2(n1003), .ZN(n1192) );
INV_X1 U885 ( .A(n1179), .ZN(n1003) );
INV_X1 U886 ( .A(n1185), .ZN(n1188) );
NAND2_X1 U887 ( .A1(n1193), .A2(n1194), .ZN(n1185) );
NAND3_X1 U888 ( .A1(G902), .A2(n1021), .A3(n1061), .ZN(n1194) );
NOR2_X1 U889 ( .A1(n1011), .A2(G900), .ZN(n1061) );
XNOR2_X1 U890 ( .A(G122), .B(n1157), .ZN(G24) );
NAND4_X1 U891 ( .A1(n1181), .A2(n1027), .A3(n1160), .A4(n1183), .ZN(n1157) );
NOR2_X1 U892 ( .A1(n1195), .A2(n1033), .ZN(n1027) );
XOR2_X1 U893 ( .A(G119), .B(n1155), .Z(G21) );
AND4_X1 U894 ( .A1(n1196), .A2(n1033), .A3(n996), .A4(n1197), .ZN(n1155) );
NOR2_X1 U895 ( .A1(n1000), .A2(n1195), .ZN(n1197) );
INV_X1 U896 ( .A(n1024), .ZN(n996) );
XNOR2_X1 U897 ( .A(G116), .B(n1198), .ZN(G18) );
NAND2_X1 U898 ( .A1(n1161), .A2(n1159), .ZN(n1198) );
NOR2_X1 U899 ( .A1(n1181), .A2(n1199), .ZN(n1159) );
XOR2_X1 U900 ( .A(n1200), .B(n1201), .Z(G15) );
NAND2_X1 U901 ( .A1(KEYINPUT1), .A2(G113), .ZN(n1201) );
NAND2_X1 U902 ( .A1(n1202), .A2(n1161), .ZN(n1200) );
AND3_X1 U903 ( .A1(n1160), .A2(n1033), .A3(n1018), .ZN(n1161) );
INV_X1 U904 ( .A(n1195), .ZN(n1018) );
NAND2_X1 U905 ( .A1(n1026), .A2(n1203), .ZN(n1195) );
AND2_X1 U906 ( .A1(n1196), .A2(n1024), .ZN(n1160) );
XNOR2_X1 U907 ( .A(n1163), .B(KEYINPUT24), .ZN(n1202) );
NOR2_X1 U908 ( .A1(n1204), .A2(n1183), .ZN(n1163) );
XOR2_X1 U909 ( .A(n1154), .B(n1205), .Z(G12) );
NOR2_X1 U910 ( .A1(KEYINPUT17), .A2(n1206), .ZN(n1205) );
INV_X1 U911 ( .A(G110), .ZN(n1206) );
AND4_X1 U912 ( .A1(n1019), .A2(n1196), .A3(n1158), .A4(n1207), .ZN(n1154) );
NOR2_X1 U913 ( .A1(n1000), .A2(n1024), .ZN(n1207) );
XOR2_X1 U914 ( .A(n1208), .B(n1039), .Z(n1024) );
NAND2_X1 U915 ( .A1(G217), .A2(n1209), .ZN(n1039) );
XNOR2_X1 U916 ( .A(n1037), .B(KEYINPUT37), .ZN(n1208) );
NOR2_X1 U917 ( .A1(n1098), .A2(G902), .ZN(n1037) );
XNOR2_X1 U918 ( .A(n1210), .B(n1211), .ZN(n1098) );
XOR2_X1 U919 ( .A(n1212), .B(n1213), .Z(n1211) );
NAND2_X1 U920 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND2_X1 U921 ( .A1(G110), .A2(n1216), .ZN(n1215) );
XOR2_X1 U922 ( .A(KEYINPUT31), .B(n1217), .Z(n1214) );
NOR2_X1 U923 ( .A1(G110), .A2(n1216), .ZN(n1217) );
XNOR2_X1 U924 ( .A(n1190), .B(G119), .ZN(n1216) );
NAND3_X1 U925 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1212) );
NAND2_X1 U926 ( .A1(KEYINPUT54), .A2(n1063), .ZN(n1220) );
NAND3_X1 U927 ( .A1(n1221), .A2(n1222), .A3(n1178), .ZN(n1219) );
INV_X1 U928 ( .A(KEYINPUT54), .ZN(n1222) );
OR2_X1 U929 ( .A1(n1178), .A2(n1221), .ZN(n1218) );
NOR2_X1 U930 ( .A1(KEYINPUT46), .A2(n1063), .ZN(n1221) );
XNOR2_X1 U931 ( .A(G125), .B(G140), .ZN(n1063) );
INV_X1 U932 ( .A(G146), .ZN(n1178) );
NAND2_X1 U933 ( .A1(n1223), .A2(n1224), .ZN(n1210) );
NAND2_X1 U934 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U935 ( .A(n1227), .B(KEYINPUT26), .Z(n1223) );
OR2_X1 U936 ( .A1(n1226), .A2(n1225), .ZN(n1227) );
AND3_X1 U937 ( .A1(G234), .A2(n1011), .A3(G221), .ZN(n1225) );
XOR2_X1 U938 ( .A(G137), .B(KEYINPUT47), .Z(n1226) );
INV_X1 U939 ( .A(n1187), .ZN(n1000) );
NOR2_X1 U940 ( .A1(n1183), .A2(n1181), .ZN(n1187) );
INV_X1 U941 ( .A(n1204), .ZN(n1181) );
XOR2_X1 U942 ( .A(n1228), .B(n1229), .Z(n1204) );
INV_X1 U943 ( .A(n1044), .ZN(n1229) );
NOR2_X1 U944 ( .A1(n1112), .A2(G902), .ZN(n1044) );
XNOR2_X1 U945 ( .A(n1230), .B(n1231), .ZN(n1112) );
XOR2_X1 U946 ( .A(n1232), .B(n1233), .Z(n1231) );
NAND2_X1 U947 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U948 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U949 ( .A1(n1238), .A2(G122), .ZN(n1234) );
XNOR2_X1 U950 ( .A(KEYINPUT3), .B(n1236), .ZN(n1238) );
XOR2_X1 U951 ( .A(n1239), .B(n1240), .Z(n1236) );
NOR2_X1 U952 ( .A1(G140), .A2(KEYINPUT60), .ZN(n1240) );
XNOR2_X1 U953 ( .A(G113), .B(G125), .ZN(n1239) );
NAND2_X1 U954 ( .A1(n1241), .A2(KEYINPUT11), .ZN(n1232) );
XOR2_X1 U955 ( .A(n1242), .B(G131), .Z(n1241) );
NAND2_X1 U956 ( .A1(n1243), .A2(KEYINPUT63), .ZN(n1242) );
XOR2_X1 U957 ( .A(n1244), .B(G143), .Z(n1243) );
NAND4_X1 U958 ( .A1(KEYINPUT57), .A2(G214), .A3(n1245), .A4(n1011), .ZN(n1244) );
XNOR2_X1 U959 ( .A(G104), .B(G146), .ZN(n1230) );
NAND2_X1 U960 ( .A1(KEYINPUT35), .A2(n1113), .ZN(n1228) );
INV_X1 U961 ( .A(G475), .ZN(n1113) );
INV_X1 U962 ( .A(n1199), .ZN(n1183) );
NOR2_X1 U963 ( .A1(n1246), .A2(n1040), .ZN(n1199) );
NOR2_X1 U964 ( .A1(n1247), .A2(n1248), .ZN(n1040) );
XNOR2_X1 U965 ( .A(KEYINPUT32), .B(n1042), .ZN(n1246) );
AND2_X1 U966 ( .A1(n1248), .A2(n1247), .ZN(n1042) );
XNOR2_X1 U967 ( .A(n1107), .B(KEYINPUT55), .ZN(n1247) );
INV_X1 U968 ( .A(G478), .ZN(n1107) );
NOR2_X1 U969 ( .A1(n1106), .A2(G902), .ZN(n1248) );
XNOR2_X1 U970 ( .A(n1249), .B(n1250), .ZN(n1106) );
XNOR2_X1 U971 ( .A(n1251), .B(n1252), .ZN(n1250) );
NAND2_X1 U972 ( .A1(KEYINPUT53), .A2(n1253), .ZN(n1251) );
XOR2_X1 U973 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U974 ( .A(G116), .B(G107), .Z(n1255) );
XNOR2_X1 U975 ( .A(KEYINPUT27), .B(n1237), .ZN(n1254) );
XOR2_X1 U976 ( .A(n1256), .B(G134), .Z(n1249) );
NAND3_X1 U977 ( .A1(G234), .A2(n1011), .A3(G217), .ZN(n1256) );
NOR2_X1 U978 ( .A1(n1026), .A2(n1025), .ZN(n1158) );
INV_X1 U979 ( .A(n1203), .ZN(n1025) );
NAND2_X1 U980 ( .A1(G221), .A2(n1209), .ZN(n1203) );
NAND2_X1 U981 ( .A1(G234), .A2(n1257), .ZN(n1209) );
XNOR2_X1 U982 ( .A(n1046), .B(n1048), .ZN(n1026) );
INV_X1 U983 ( .A(G469), .ZN(n1048) );
NAND2_X1 U984 ( .A1(n1258), .A2(n1257), .ZN(n1046) );
XOR2_X1 U985 ( .A(n1259), .B(n1260), .Z(n1258) );
XNOR2_X1 U986 ( .A(n1261), .B(n1262), .ZN(n1260) );
INV_X1 U987 ( .A(n1138), .ZN(n1262) );
XNOR2_X1 U988 ( .A(n1263), .B(G140), .ZN(n1138) );
XOR2_X1 U989 ( .A(n1140), .B(n1264), .Z(n1261) );
NOR2_X1 U990 ( .A1(KEYINPUT22), .A2(n1078), .ZN(n1264) );
XNOR2_X1 U991 ( .A(n1265), .B(n1190), .ZN(n1078) );
NAND2_X1 U992 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
OR2_X1 U993 ( .A1(n1268), .A2(G143), .ZN(n1267) );
XOR2_X1 U994 ( .A(n1269), .B(KEYINPUT45), .Z(n1266) );
NAND2_X1 U995 ( .A1(G143), .A2(n1268), .ZN(n1269) );
XOR2_X1 U996 ( .A(G146), .B(KEYINPUT21), .Z(n1268) );
XNOR2_X1 U997 ( .A(G101), .B(n1270), .ZN(n1140) );
XOR2_X1 U998 ( .A(n1271), .B(n1272), .Z(n1259) );
NOR2_X1 U999 ( .A1(KEYINPUT8), .A2(G110), .ZN(n1272) );
XNOR2_X1 U1000 ( .A(KEYINPUT15), .B(n1273), .ZN(n1271) );
NOR2_X1 U1001 ( .A1(KEYINPUT4), .A2(n1274), .ZN(n1273) );
XNOR2_X1 U1002 ( .A(n1143), .B(KEYINPUT14), .ZN(n1274) );
AND2_X1 U1003 ( .A1(G227), .A2(n1011), .ZN(n1143) );
AND2_X1 U1004 ( .A1(n1179), .A2(n1275), .ZN(n1196) );
NAND2_X1 U1005 ( .A1(n1193), .A2(n1276), .ZN(n1275) );
NAND3_X1 U1006 ( .A1(n1277), .A2(n1021), .A3(G902), .ZN(n1276) );
INV_X1 U1007 ( .A(n1085), .ZN(n1277) );
NAND2_X1 U1008 ( .A1(G953), .A2(n1278), .ZN(n1085) );
XOR2_X1 U1009 ( .A(KEYINPUT25), .B(G898), .Z(n1278) );
NAND3_X1 U1010 ( .A1(n1021), .A2(n1011), .A3(G952), .ZN(n1193) );
NAND2_X1 U1011 ( .A1(G237), .A2(G234), .ZN(n1021) );
NOR2_X1 U1012 ( .A1(n1279), .A2(n1043), .ZN(n1179) );
INV_X1 U1013 ( .A(n1006), .ZN(n1043) );
NAND2_X1 U1014 ( .A1(G214), .A2(n1280), .ZN(n1006) );
INV_X1 U1015 ( .A(n1007), .ZN(n1279) );
XOR2_X1 U1016 ( .A(n1041), .B(KEYINPUT61), .Z(n1007) );
XNOR2_X1 U1017 ( .A(n1281), .B(n1282), .ZN(n1041) );
AND2_X1 U1018 ( .A1(n1280), .A2(G210), .ZN(n1282) );
NAND2_X1 U1019 ( .A1(n1257), .A2(n1245), .ZN(n1280) );
NAND2_X1 U1020 ( .A1(n1283), .A2(n1257), .ZN(n1281) );
XNOR2_X1 U1021 ( .A(n1284), .B(n1285), .ZN(n1283) );
INV_X1 U1022 ( .A(n1147), .ZN(n1285) );
XNOR2_X1 U1023 ( .A(n1286), .B(n1088), .ZN(n1147) );
XNOR2_X1 U1024 ( .A(n1237), .B(G110), .ZN(n1088) );
INV_X1 U1025 ( .A(G122), .ZN(n1237) );
NAND2_X1 U1026 ( .A1(KEYINPUT18), .A2(n1086), .ZN(n1286) );
XOR2_X1 U1027 ( .A(n1287), .B(n1288), .Z(n1086) );
XNOR2_X1 U1028 ( .A(G101), .B(n1289), .ZN(n1288) );
NAND3_X1 U1029 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1289) );
OR2_X1 U1030 ( .A1(n1293), .A2(KEYINPUT59), .ZN(n1292) );
NAND3_X1 U1031 ( .A1(KEYINPUT59), .A2(n1294), .A3(n1295), .ZN(n1291) );
INV_X1 U1032 ( .A(n1296), .ZN(n1294) );
NAND2_X1 U1033 ( .A1(G113), .A2(n1296), .ZN(n1290) );
NAND2_X1 U1034 ( .A1(KEYINPUT50), .A2(n1293), .ZN(n1296) );
NAND2_X1 U1035 ( .A1(KEYINPUT33), .A2(n1270), .ZN(n1287) );
XOR2_X1 U1036 ( .A(G107), .B(G104), .Z(n1270) );
NAND2_X1 U1037 ( .A1(n1297), .A2(n1298), .ZN(n1284) );
NAND2_X1 U1038 ( .A1(n1299), .A2(n1175), .ZN(n1298) );
XOR2_X1 U1039 ( .A(n1300), .B(KEYINPUT36), .Z(n1297) );
OR2_X1 U1040 ( .A1(n1175), .A2(n1299), .ZN(n1300) );
XOR2_X1 U1041 ( .A(n1177), .B(n1301), .Z(n1299) );
XOR2_X1 U1042 ( .A(KEYINPUT9), .B(G125), .Z(n1301) );
NAND2_X1 U1043 ( .A1(G224), .A2(n1011), .ZN(n1175) );
INV_X1 U1044 ( .A(n1033), .ZN(n1019) );
XOR2_X1 U1045 ( .A(n1302), .B(n1133), .Z(n1033) );
INV_X1 U1046 ( .A(G472), .ZN(n1133) );
NAND2_X1 U1047 ( .A1(n1303), .A2(n1257), .ZN(n1302) );
INV_X1 U1048 ( .A(G902), .ZN(n1257) );
XNOR2_X1 U1049 ( .A(n1304), .B(n1305), .ZN(n1303) );
INV_X1 U1050 ( .A(n1131), .ZN(n1305) );
XNOR2_X1 U1051 ( .A(n1306), .B(n1307), .ZN(n1131) );
XNOR2_X1 U1052 ( .A(n1295), .B(n1293), .ZN(n1307) );
XOR2_X1 U1053 ( .A(G116), .B(G119), .Z(n1293) );
INV_X1 U1054 ( .A(G113), .ZN(n1295) );
XNOR2_X1 U1055 ( .A(n1263), .B(n1308), .ZN(n1306) );
INV_X1 U1056 ( .A(n1177), .ZN(n1308) );
XOR2_X1 U1057 ( .A(G146), .B(n1252), .Z(n1177) );
XNOR2_X1 U1058 ( .A(n1190), .B(G143), .ZN(n1252) );
INV_X1 U1059 ( .A(G128), .ZN(n1190) );
XOR2_X1 U1060 ( .A(n1077), .B(G131), .Z(n1263) );
XNOR2_X1 U1061 ( .A(G134), .B(n1309), .ZN(n1077) );
XOR2_X1 U1062 ( .A(KEYINPUT12), .B(G137), .Z(n1309) );
NOR2_X1 U1063 ( .A1(KEYINPUT2), .A2(n1310), .ZN(n1304) );
XNOR2_X1 U1064 ( .A(n1130), .B(n1128), .ZN(n1310) );
INV_X1 U1065 ( .A(G101), .ZN(n1128) );
NAND3_X1 U1066 ( .A1(n1245), .A2(n1011), .A3(G210), .ZN(n1130) );
INV_X1 U1067 ( .A(G953), .ZN(n1011) );
INV_X1 U1068 ( .A(G237), .ZN(n1245) );
endmodule


