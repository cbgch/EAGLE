//Key = 0001111100111101101111010010010000001010001100000111001100100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367;

XNOR2_X1 U741 ( .A(G107), .B(n1029), .ZN(G9) );
NOR2_X1 U742 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U743 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
NOR2_X1 U744 ( .A1(KEYINPUT23), .A2(n1036), .ZN(n1035) );
NOR3_X1 U745 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NOR2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1034) );
NOR2_X1 U747 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U748 ( .A1(n1044), .A2(n1037), .ZN(n1043) );
NOR3_X1 U749 ( .A1(n1045), .A2(n1046), .A3(n1038), .ZN(n1042) );
NOR2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U751 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1047) );
NOR2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
AND2_X1 U754 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U755 ( .A1(n1057), .A2(n1058), .ZN(n1053) );
NOR2_X1 U756 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U757 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NAND4_X1 U758 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1032) );
NAND3_X1 U759 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1064) );
XOR2_X1 U760 ( .A(n1070), .B(KEYINPUT44), .Z(n1069) );
XOR2_X1 U761 ( .A(KEYINPUT56), .B(n1071), .Z(n1068) );
NOR2_X1 U762 ( .A1(n1041), .A2(n1037), .ZN(n1071) );
INV_X1 U763 ( .A(n1072), .ZN(n1037) );
NAND3_X1 U764 ( .A1(n1073), .A2(n1074), .A3(n1072), .ZN(n1063) );
NOR4_X1 U765 ( .A1(n1045), .A2(n1049), .A3(n1058), .A4(n1052), .ZN(n1072) );
NAND2_X1 U766 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U767 ( .A1(KEYINPUT23), .A2(n1077), .ZN(n1076) );
NOR3_X1 U768 ( .A1(n1078), .A2(G953), .A3(G952), .ZN(n1030) );
INV_X1 U769 ( .A(n1065), .ZN(n1078) );
NAND4_X1 U770 ( .A1(n1079), .A2(n1073), .A3(n1080), .A4(n1081), .ZN(n1065) );
NOR4_X1 U771 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1081) );
XOR2_X1 U772 ( .A(n1086), .B(n1087), .Z(n1085) );
XOR2_X1 U773 ( .A(KEYINPUT55), .B(G478), .Z(n1087) );
NOR3_X1 U774 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1084) );
NOR2_X1 U775 ( .A1(KEYINPUT31), .A2(n1091), .ZN(n1090) );
INV_X1 U776 ( .A(n1092), .ZN(n1091) );
NOR2_X1 U777 ( .A1(n1093), .A2(n1092), .ZN(n1089) );
NOR2_X1 U778 ( .A1(KEYINPUT31), .A2(G472), .ZN(n1093) );
INV_X1 U779 ( .A(KEYINPUT58), .ZN(n1088) );
NOR2_X1 U780 ( .A1(n1094), .A2(n1095), .ZN(n1083) );
NOR2_X1 U781 ( .A1(n1096), .A2(n1092), .ZN(n1094) );
XOR2_X1 U782 ( .A(n1097), .B(KEYINPUT0), .Z(n1092) );
NOR2_X1 U783 ( .A1(KEYINPUT58), .A2(KEYINPUT31), .ZN(n1096) );
NOR2_X1 U784 ( .A1(n1058), .A2(n1098), .ZN(n1080) );
INV_X1 U785 ( .A(n1099), .ZN(n1058) );
XOR2_X1 U786 ( .A(n1100), .B(G469), .Z(n1079) );
XOR2_X1 U787 ( .A(n1101), .B(n1102), .Z(G72) );
XOR2_X1 U788 ( .A(n1103), .B(n1104), .Z(n1102) );
NAND2_X1 U789 ( .A1(n1066), .A2(n1105), .ZN(n1104) );
NAND2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1103) );
NAND2_X1 U791 ( .A1(G953), .A2(n1108), .ZN(n1107) );
XNOR2_X1 U792 ( .A(n1109), .B(n1110), .ZN(n1106) );
XOR2_X1 U793 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U794 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U795 ( .A(KEYINPUT25), .B(n1115), .Z(n1114) );
NOR2_X1 U796 ( .A1(G125), .A2(n1116), .ZN(n1115) );
INV_X1 U797 ( .A(n1117), .ZN(n1113) );
NOR3_X1 U798 ( .A1(n1066), .A2(KEYINPUT1), .A3(n1118), .ZN(n1101) );
NOR2_X1 U799 ( .A1(n1119), .A2(n1108), .ZN(n1118) );
XOR2_X1 U800 ( .A(n1120), .B(n1121), .Z(G69) );
NOR2_X1 U801 ( .A1(n1122), .A2(n1066), .ZN(n1121) );
XOR2_X1 U802 ( .A(n1123), .B(KEYINPUT16), .Z(n1122) );
NAND2_X1 U803 ( .A1(G224), .A2(n1124), .ZN(n1123) );
XOR2_X1 U804 ( .A(KEYINPUT17), .B(G898), .Z(n1124) );
NAND2_X1 U805 ( .A1(n1125), .A2(n1126), .ZN(n1120) );
NAND2_X1 U806 ( .A1(n1127), .A2(n1066), .ZN(n1126) );
XOR2_X1 U807 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND2_X1 U808 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
XOR2_X1 U809 ( .A(n1132), .B(KEYINPUT28), .Z(n1130) );
NAND3_X1 U810 ( .A1(G898), .A2(n1129), .A3(G953), .ZN(n1125) );
XOR2_X1 U811 ( .A(n1133), .B(KEYINPUT9), .Z(n1129) );
NOR2_X1 U812 ( .A1(n1134), .A2(n1135), .ZN(G66) );
XNOR2_X1 U813 ( .A(n1136), .B(n1137), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR2_X1 U815 ( .A1(n1134), .A2(n1140), .ZN(G63) );
NOR3_X1 U816 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1140) );
NOR3_X1 U817 ( .A1(n1144), .A2(n1145), .A3(n1139), .ZN(n1143) );
INV_X1 U818 ( .A(G478), .ZN(n1145) );
NOR2_X1 U819 ( .A1(n1146), .A2(n1147), .ZN(n1142) );
AND2_X1 U820 ( .A1(n1033), .A2(G478), .ZN(n1146) );
NOR2_X1 U821 ( .A1(n1134), .A2(n1148), .ZN(G60) );
XNOR2_X1 U822 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR2_X1 U823 ( .A1(n1151), .A2(n1139), .ZN(n1150) );
INV_X1 U824 ( .A(G475), .ZN(n1151) );
XOR2_X1 U825 ( .A(n1152), .B(n1153), .Z(G6) );
NOR2_X1 U826 ( .A1(n1154), .A2(n1044), .ZN(n1153) );
XOR2_X1 U827 ( .A(n1155), .B(KEYINPUT40), .Z(n1154) );
XNOR2_X1 U828 ( .A(G104), .B(KEYINPUT12), .ZN(n1152) );
NOR2_X1 U829 ( .A1(n1134), .A2(n1156), .ZN(G57) );
XOR2_X1 U830 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U831 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U832 ( .A(n1161), .B(n1162), .Z(n1159) );
NOR2_X1 U833 ( .A1(n1095), .A2(n1139), .ZN(n1162) );
INV_X1 U834 ( .A(G472), .ZN(n1095) );
XOR2_X1 U835 ( .A(n1163), .B(n1164), .Z(n1157) );
XOR2_X1 U836 ( .A(G101), .B(n1165), .Z(n1164) );
NOR2_X1 U837 ( .A1(n1134), .A2(n1166), .ZN(G54) );
XOR2_X1 U838 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U839 ( .A(n1169), .B(n1170), .Z(n1168) );
NAND2_X1 U840 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND2_X1 U841 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
INV_X1 U842 ( .A(KEYINPUT57), .ZN(n1174) );
NAND3_X1 U843 ( .A1(G140), .A2(n1175), .A3(KEYINPUT57), .ZN(n1171) );
XOR2_X1 U844 ( .A(n1176), .B(n1177), .Z(n1167) );
NOR2_X1 U845 ( .A1(n1178), .A2(n1139), .ZN(n1176) );
INV_X1 U846 ( .A(G469), .ZN(n1178) );
NOR2_X1 U847 ( .A1(n1134), .A2(n1179), .ZN(G51) );
XOR2_X1 U848 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U849 ( .A(n1182), .B(n1183), .Z(n1181) );
NAND3_X1 U850 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1182) );
OR2_X1 U851 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND3_X1 U852 ( .A1(n1188), .A2(n1187), .A3(KEYINPUT5), .ZN(n1185) );
NOR2_X1 U853 ( .A1(KEYINPUT59), .A2(n1189), .ZN(n1188) );
NAND2_X1 U854 ( .A1(n1189), .A2(n1190), .ZN(n1184) );
INV_X1 U855 ( .A(KEYINPUT5), .ZN(n1190) );
XNOR2_X1 U856 ( .A(KEYINPUT33), .B(n1191), .ZN(n1180) );
NOR2_X1 U857 ( .A1(KEYINPUT24), .A2(n1192), .ZN(n1191) );
NOR3_X1 U858 ( .A1(n1193), .A2(n1194), .A3(n1139), .ZN(n1192) );
NAND2_X1 U859 ( .A1(G902), .A2(n1033), .ZN(n1139) );
NAND3_X1 U860 ( .A1(n1131), .A2(n1132), .A3(n1195), .ZN(n1033) );
INV_X1 U861 ( .A(n1105), .ZN(n1195) );
NAND4_X1 U862 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1105) );
NOR4_X1 U863 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
NAND2_X1 U864 ( .A1(n1204), .A2(n1205), .ZN(n1198) );
NAND2_X1 U865 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND3_X1 U866 ( .A1(n1098), .A2(n1208), .A3(n1209), .ZN(n1207) );
NAND2_X1 U867 ( .A1(n1077), .A2(n1073), .ZN(n1206) );
AND4_X1 U868 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1131) );
AND3_X1 U869 ( .A1(n1214), .A2(n1029), .A3(n1215), .ZN(n1213) );
NAND3_X1 U870 ( .A1(n1099), .A2(n1216), .A3(n1217), .ZN(n1029) );
NAND2_X1 U871 ( .A1(n1209), .A2(n1218), .ZN(n1212) );
NAND2_X1 U872 ( .A1(n1155), .A2(n1219), .ZN(n1218) );
NAND3_X1 U873 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1219) );
XOR2_X1 U874 ( .A(KEYINPUT42), .B(n1223), .Z(n1221) );
NAND4_X1 U875 ( .A1(n1077), .A2(n1217), .A3(n1099), .A4(n1224), .ZN(n1155) );
NAND2_X1 U876 ( .A1(n1055), .A2(n1225), .ZN(n1211) );
NAND2_X1 U877 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
OR2_X1 U878 ( .A1(n1228), .A2(KEYINPUT47), .ZN(n1227) );
NAND2_X1 U879 ( .A1(n1229), .A2(n1216), .ZN(n1226) );
NAND3_X1 U880 ( .A1(KEYINPUT47), .A2(n1230), .A3(n1049), .ZN(n1210) );
INV_X1 U881 ( .A(n1228), .ZN(n1230) );
XOR2_X1 U882 ( .A(KEYINPUT53), .B(n1231), .Z(n1193) );
NOR2_X1 U883 ( .A1(n1066), .A2(G952), .ZN(n1134) );
XOR2_X1 U884 ( .A(n1232), .B(n1203), .Z(G48) );
NOR3_X1 U885 ( .A1(n1039), .A2(n1044), .A3(n1233), .ZN(n1203) );
INV_X1 U886 ( .A(n1077), .ZN(n1039) );
NAND2_X1 U887 ( .A1(KEYINPUT63), .A2(n1234), .ZN(n1232) );
XOR2_X1 U888 ( .A(n1235), .B(n1236), .Z(G45) );
NAND2_X1 U889 ( .A1(KEYINPUT15), .A2(G143), .ZN(n1236) );
NAND4_X1 U890 ( .A1(n1237), .A2(n1204), .A3(n1098), .A4(n1208), .ZN(n1235) );
INV_X1 U891 ( .A(n1238), .ZN(n1204) );
XOR2_X1 U892 ( .A(n1044), .B(KEYINPUT19), .Z(n1237) );
XOR2_X1 U893 ( .A(n1116), .B(n1196), .Z(G42) );
NAND3_X1 U894 ( .A1(n1073), .A2(n1217), .A3(n1239), .ZN(n1196) );
XOR2_X1 U895 ( .A(G137), .B(n1202), .Z(G39) );
NOR3_X1 U896 ( .A1(n1233), .A2(n1038), .A3(n1041), .ZN(n1202) );
XOR2_X1 U897 ( .A(G134), .B(n1201), .Z(G36) );
NOR3_X1 U898 ( .A1(n1038), .A2(n1075), .A3(n1238), .ZN(n1201) );
XOR2_X1 U899 ( .A(n1240), .B(n1241), .Z(G33) );
NOR3_X1 U900 ( .A1(n1242), .A2(n1038), .A3(n1238), .ZN(n1241) );
NAND2_X1 U901 ( .A1(n1220), .A2(n1243), .ZN(n1238) );
INV_X1 U902 ( .A(n1073), .ZN(n1038) );
NOR2_X1 U903 ( .A1(n1244), .A2(n1067), .ZN(n1073) );
INV_X1 U904 ( .A(n1070), .ZN(n1244) );
XOR2_X1 U905 ( .A(KEYINPUT49), .B(n1077), .Z(n1242) );
XNOR2_X1 U906 ( .A(G131), .B(KEYINPUT50), .ZN(n1240) );
XOR2_X1 U907 ( .A(G128), .B(n1200), .Z(G30) );
NOR3_X1 U908 ( .A1(n1044), .A2(n1075), .A3(n1233), .ZN(n1200) );
NAND4_X1 U909 ( .A1(n1056), .A2(n1060), .A3(n1245), .A4(n1243), .ZN(n1233) );
XNOR2_X1 U910 ( .A(G101), .B(n1246), .ZN(G3) );
NAND2_X1 U911 ( .A1(n1247), .A2(n1220), .ZN(n1246) );
AND2_X1 U912 ( .A1(n1229), .A2(n1060), .ZN(n1220) );
XOR2_X1 U913 ( .A(G125), .B(n1248), .Z(G27) );
NOR2_X1 U914 ( .A1(KEYINPUT37), .A2(n1197), .ZN(n1248) );
NAND3_X1 U915 ( .A1(n1249), .A2(n1250), .A3(n1239), .ZN(n1197) );
AND3_X1 U916 ( .A1(n1077), .A2(n1243), .A3(n1056), .ZN(n1239) );
NAND2_X1 U917 ( .A1(n1045), .A2(n1251), .ZN(n1243) );
NAND4_X1 U918 ( .A1(n1252), .A2(G953), .A3(n1253), .A4(n1108), .ZN(n1251) );
INV_X1 U919 ( .A(G900), .ZN(n1108) );
XOR2_X1 U920 ( .A(n1254), .B(KEYINPUT21), .Z(n1252) );
XOR2_X1 U921 ( .A(n1255), .B(n1214), .Z(G24) );
NAND4_X1 U922 ( .A1(n1099), .A2(n1098), .A3(n1249), .A4(n1256), .ZN(n1214) );
AND3_X1 U923 ( .A1(n1208), .A2(n1224), .A3(n1250), .ZN(n1256) );
XOR2_X1 U924 ( .A(G119), .B(n1257), .Z(G21) );
NOR2_X1 U925 ( .A1(n1049), .A2(n1228), .ZN(n1257) );
NAND3_X1 U926 ( .A1(n1056), .A2(n1245), .A3(n1247), .ZN(n1228) );
XOR2_X1 U927 ( .A(n1258), .B(n1259), .Z(G18) );
NAND3_X1 U928 ( .A1(n1229), .A2(n1216), .A3(n1260), .ZN(n1259) );
XOR2_X1 U929 ( .A(n1049), .B(KEYINPUT26), .Z(n1260) );
NOR3_X1 U930 ( .A1(n1075), .A2(n1223), .A3(n1044), .ZN(n1216) );
NAND2_X1 U931 ( .A1(n1261), .A2(n1208), .ZN(n1075) );
XNOR2_X1 U932 ( .A(G113), .B(n1132), .ZN(G15) );
NAND4_X1 U933 ( .A1(n1229), .A2(n1077), .A3(n1249), .A4(n1224), .ZN(n1132) );
NOR2_X1 U934 ( .A1(n1049), .A2(n1044), .ZN(n1249) );
INV_X1 U935 ( .A(n1055), .ZN(n1049) );
NOR2_X1 U936 ( .A1(n1061), .A2(n1082), .ZN(n1055) );
INV_X1 U937 ( .A(n1062), .ZN(n1082) );
NOR2_X1 U938 ( .A1(n1208), .A2(n1261), .ZN(n1077) );
INV_X1 U939 ( .A(n1050), .ZN(n1229) );
NAND2_X1 U940 ( .A1(n1099), .A2(n1245), .ZN(n1050) );
XOR2_X1 U941 ( .A(n1250), .B(KEYINPUT20), .Z(n1245) );
XOR2_X1 U942 ( .A(n1175), .B(n1215), .Z(G12) );
NAND3_X1 U943 ( .A1(n1056), .A2(n1217), .A3(n1247), .ZN(n1215) );
NOR3_X1 U944 ( .A1(n1044), .A2(n1223), .A3(n1041), .ZN(n1247) );
INV_X1 U945 ( .A(n1222), .ZN(n1041) );
NOR2_X1 U946 ( .A1(n1208), .A2(n1098), .ZN(n1222) );
INV_X1 U947 ( .A(n1261), .ZN(n1098) );
XOR2_X1 U948 ( .A(n1262), .B(G475), .Z(n1261) );
NAND2_X1 U949 ( .A1(n1149), .A2(n1254), .ZN(n1262) );
XOR2_X1 U950 ( .A(n1263), .B(n1264), .Z(n1149) );
XNOR2_X1 U951 ( .A(n1265), .B(n1266), .ZN(n1264) );
NOR2_X1 U952 ( .A1(KEYINPUT32), .A2(n1267), .ZN(n1266) );
XOR2_X1 U953 ( .A(n1268), .B(n1269), .Z(n1267) );
XNOR2_X1 U954 ( .A(n1270), .B(n1271), .ZN(n1269) );
NOR2_X1 U955 ( .A1(G131), .A2(KEYINPUT27), .ZN(n1271) );
NAND2_X1 U956 ( .A1(n1272), .A2(KEYINPUT10), .ZN(n1270) );
XOR2_X1 U957 ( .A(n1234), .B(n1273), .Z(n1272) );
XOR2_X1 U958 ( .A(n1274), .B(n1275), .Z(n1268) );
NAND4_X1 U959 ( .A1(KEYINPUT62), .A2(G214), .A3(n1276), .A4(n1277), .ZN(n1275) );
NAND2_X1 U960 ( .A1(KEYINPUT4), .A2(n1255), .ZN(n1265) );
XNOR2_X1 U961 ( .A(n1278), .B(n1141), .ZN(n1208) );
INV_X1 U962 ( .A(n1086), .ZN(n1141) );
NAND2_X1 U963 ( .A1(n1144), .A2(n1254), .ZN(n1086) );
INV_X1 U964 ( .A(n1147), .ZN(n1144) );
XOR2_X1 U965 ( .A(n1279), .B(n1280), .Z(n1147) );
XOR2_X1 U966 ( .A(n1281), .B(n1282), .Z(n1280) );
XOR2_X1 U967 ( .A(n1283), .B(n1284), .Z(n1282) );
NAND2_X1 U968 ( .A1(KEYINPUT18), .A2(G128), .ZN(n1284) );
NAND2_X1 U969 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
NAND2_X1 U970 ( .A1(G116), .A2(n1255), .ZN(n1286) );
INV_X1 U971 ( .A(G122), .ZN(n1255) );
XOR2_X1 U972 ( .A(n1287), .B(KEYINPUT35), .Z(n1285) );
NAND2_X1 U973 ( .A1(G122), .A2(n1258), .ZN(n1287) );
INV_X1 U974 ( .A(G116), .ZN(n1258) );
NOR2_X1 U975 ( .A1(KEYINPUT14), .A2(n1288), .ZN(n1281) );
XOR2_X1 U976 ( .A(n1289), .B(n1290), .Z(n1279) );
XOR2_X1 U977 ( .A(G143), .B(G134), .Z(n1290) );
NAND2_X1 U978 ( .A1(n1291), .A2(n1292), .ZN(n1289) );
XOR2_X1 U979 ( .A(KEYINPUT8), .B(G217), .Z(n1292) );
NAND2_X1 U980 ( .A1(KEYINPUT38), .A2(G478), .ZN(n1278) );
INV_X1 U981 ( .A(n1224), .ZN(n1223) );
NAND2_X1 U982 ( .A1(n1045), .A2(n1293), .ZN(n1224) );
NAND4_X1 U983 ( .A1(G953), .A2(G902), .A3(n1253), .A4(n1294), .ZN(n1293) );
INV_X1 U984 ( .A(G898), .ZN(n1294) );
NAND3_X1 U985 ( .A1(n1253), .A2(n1066), .A3(G952), .ZN(n1045) );
NAND2_X1 U986 ( .A1(G237), .A2(G234), .ZN(n1253) );
INV_X1 U987 ( .A(n1209), .ZN(n1044) );
NOR2_X1 U988 ( .A1(n1070), .A2(n1067), .ZN(n1209) );
AND2_X1 U989 ( .A1(G214), .A2(n1295), .ZN(n1067) );
XOR2_X1 U990 ( .A(n1296), .B(n1297), .Z(n1070) );
NOR2_X1 U991 ( .A1(n1231), .A2(n1298), .ZN(n1297) );
XOR2_X1 U992 ( .A(n1194), .B(KEYINPUT46), .Z(n1298) );
INV_X1 U993 ( .A(n1295), .ZN(n1231) );
NAND2_X1 U994 ( .A1(n1299), .A2(n1277), .ZN(n1295) );
INV_X1 U995 ( .A(G237), .ZN(n1277) );
NAND2_X1 U996 ( .A1(n1300), .A2(n1254), .ZN(n1296) );
XOR2_X1 U997 ( .A(n1133), .B(n1301), .Z(n1300) );
XNOR2_X1 U998 ( .A(n1187), .B(n1302), .ZN(n1301) );
NOR2_X1 U999 ( .A1(KEYINPUT48), .A2(n1189), .ZN(n1302) );
XOR2_X1 U1000 ( .A(n1163), .B(G125), .Z(n1189) );
NAND2_X1 U1001 ( .A1(G224), .A2(n1276), .ZN(n1187) );
INV_X1 U1002 ( .A(n1183), .ZN(n1133) );
XOR2_X1 U1003 ( .A(n1303), .B(n1304), .Z(n1183) );
XOR2_X1 U1004 ( .A(n1263), .B(n1305), .Z(n1304) );
XOR2_X1 U1005 ( .A(G122), .B(G110), .Z(n1305) );
XOR2_X1 U1006 ( .A(G104), .B(G113), .Z(n1263) );
XOR2_X1 U1007 ( .A(n1306), .B(n1307), .Z(n1303) );
AND2_X1 U1008 ( .A1(n1060), .A2(n1250), .ZN(n1217) );
INV_X1 U1009 ( .A(n1052), .ZN(n1250) );
XOR2_X1 U1010 ( .A(n1097), .B(n1308), .Z(n1052) );
XOR2_X1 U1011 ( .A(KEYINPUT51), .B(G472), .Z(n1308) );
NAND2_X1 U1012 ( .A1(n1309), .A2(n1254), .ZN(n1097) );
XOR2_X1 U1013 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1014 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U1015 ( .A(KEYINPUT34), .B(G101), .Z(n1313) );
NOR2_X1 U1016 ( .A1(KEYINPUT2), .A2(n1163), .ZN(n1312) );
NAND4_X1 U1017 ( .A1(n1314), .A2(n1315), .A3(n1316), .A4(n1317), .ZN(n1163) );
NAND3_X1 U1018 ( .A1(KEYINPUT13), .A2(n1318), .A3(n1319), .ZN(n1317) );
XOR2_X1 U1019 ( .A(KEYINPUT30), .B(G128), .Z(n1318) );
OR2_X1 U1020 ( .A1(n1319), .A2(KEYINPUT13), .ZN(n1316) );
NAND3_X1 U1021 ( .A1(G128), .A2(n1320), .A3(n1321), .ZN(n1315) );
INV_X1 U1022 ( .A(KEYINPUT61), .ZN(n1321) );
NAND2_X1 U1023 ( .A1(KEYINPUT30), .A2(n1319), .ZN(n1320) );
INV_X1 U1024 ( .A(n1322), .ZN(n1319) );
NAND3_X1 U1025 ( .A1(n1323), .A2(n1324), .A3(KEYINPUT61), .ZN(n1314) );
OR2_X1 U1026 ( .A1(n1322), .A2(KEYINPUT30), .ZN(n1323) );
XOR2_X1 U1027 ( .A(n1325), .B(n1160), .Z(n1310) );
INV_X1 U1028 ( .A(n1111), .ZN(n1160) );
XNOR2_X1 U1029 ( .A(n1326), .B(n1161), .ZN(n1325) );
NAND2_X1 U1030 ( .A1(n1327), .A2(n1328), .ZN(n1161) );
NAND2_X1 U1031 ( .A1(G113), .A2(n1307), .ZN(n1328) );
XOR2_X1 U1032 ( .A(n1329), .B(KEYINPUT45), .Z(n1327) );
OR2_X1 U1033 ( .A1(n1307), .A2(G113), .ZN(n1329) );
XOR2_X1 U1034 ( .A(G119), .B(G116), .Z(n1307) );
NAND2_X1 U1035 ( .A1(KEYINPUT3), .A2(n1165), .ZN(n1326) );
NOR3_X1 U1036 ( .A1(n1330), .A2(G237), .A3(n1194), .ZN(n1165) );
INV_X1 U1037 ( .A(G210), .ZN(n1194) );
AND2_X1 U1038 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U1039 ( .A1(G221), .A2(n1331), .ZN(n1062) );
NAND2_X1 U1040 ( .A1(n1332), .A2(n1333), .ZN(n1061) );
NAND2_X1 U1041 ( .A1(G469), .A2(n1100), .ZN(n1333) );
XOR2_X1 U1042 ( .A(KEYINPUT7), .B(n1334), .Z(n1332) );
NOR2_X1 U1043 ( .A1(G469), .A2(n1100), .ZN(n1334) );
NAND2_X1 U1044 ( .A1(n1335), .A2(n1254), .ZN(n1100) );
XNOR2_X1 U1045 ( .A(n1177), .B(n1336), .ZN(n1335) );
XOR2_X1 U1046 ( .A(n1173), .B(n1337), .Z(n1336) );
NOR2_X1 U1047 ( .A1(KEYINPUT60), .A2(n1338), .ZN(n1337) );
XOR2_X1 U1048 ( .A(n1169), .B(KEYINPUT6), .Z(n1338) );
XOR2_X1 U1049 ( .A(n1339), .B(n1109), .Z(n1169) );
XNOR2_X1 U1050 ( .A(n1324), .B(n1322), .ZN(n1109) );
XNOR2_X1 U1051 ( .A(n1274), .B(G146), .ZN(n1322) );
INV_X1 U1052 ( .A(G143), .ZN(n1274) );
INV_X1 U1053 ( .A(G128), .ZN(n1324) );
XOR2_X1 U1054 ( .A(n1306), .B(G104), .Z(n1339) );
XOR2_X1 U1055 ( .A(G101), .B(n1288), .Z(n1306) );
XNOR2_X1 U1056 ( .A(G107), .B(KEYINPUT36), .ZN(n1288) );
XOR2_X1 U1057 ( .A(n1175), .B(G140), .Z(n1173) );
XNOR2_X1 U1058 ( .A(n1111), .B(n1340), .ZN(n1177) );
NOR2_X1 U1059 ( .A1(n1330), .A2(n1119), .ZN(n1340) );
INV_X1 U1060 ( .A(G227), .ZN(n1119) );
INV_X1 U1061 ( .A(n1276), .ZN(n1330) );
XNOR2_X1 U1062 ( .A(G131), .B(n1341), .ZN(n1111) );
XOR2_X1 U1063 ( .A(G137), .B(G134), .Z(n1341) );
XOR2_X1 U1064 ( .A(n1099), .B(KEYINPUT54), .Z(n1056) );
XNOR2_X1 U1065 ( .A(n1342), .B(n1138), .ZN(n1099) );
NAND2_X1 U1066 ( .A1(G217), .A2(n1331), .ZN(n1138) );
NAND2_X1 U1067 ( .A1(G234), .A2(n1299), .ZN(n1331) );
XOR2_X1 U1068 ( .A(G902), .B(KEYINPUT43), .Z(n1299) );
NAND2_X1 U1069 ( .A1(n1136), .A2(n1254), .ZN(n1342) );
INV_X1 U1070 ( .A(G902), .ZN(n1254) );
XNOR2_X1 U1071 ( .A(n1343), .B(n1344), .ZN(n1136) );
XOR2_X1 U1072 ( .A(n1345), .B(n1346), .Z(n1344) );
XOR2_X1 U1073 ( .A(G128), .B(G119), .Z(n1346) );
NOR2_X1 U1074 ( .A1(KEYINPUT39), .A2(G137), .ZN(n1345) );
XOR2_X1 U1075 ( .A(n1347), .B(n1348), .Z(n1343) );
XOR2_X1 U1076 ( .A(n1349), .B(n1350), .Z(n1348) );
NAND2_X1 U1077 ( .A1(KEYINPUT11), .A2(n1175), .ZN(n1350) );
NAND2_X1 U1078 ( .A1(n1291), .A2(G221), .ZN(n1349) );
AND2_X1 U1079 ( .A1(n1276), .A2(G234), .ZN(n1291) );
XOR2_X1 U1080 ( .A(n1066), .B(KEYINPUT22), .Z(n1276) );
INV_X1 U1081 ( .A(G953), .ZN(n1066) );
NAND3_X1 U1082 ( .A1(n1351), .A2(n1352), .A3(n1353), .ZN(n1347) );
NAND2_X1 U1083 ( .A1(G146), .A2(n1273), .ZN(n1353) );
NAND2_X1 U1084 ( .A1(KEYINPUT41), .A2(n1354), .ZN(n1352) );
NAND2_X1 U1085 ( .A1(n1355), .A2(n1234), .ZN(n1354) );
XOR2_X1 U1086 ( .A(n1273), .B(KEYINPUT29), .Z(n1355) );
NAND2_X1 U1087 ( .A1(n1356), .A2(n1357), .ZN(n1351) );
INV_X1 U1088 ( .A(KEYINPUT41), .ZN(n1357) );
NAND2_X1 U1089 ( .A1(n1358), .A2(n1359), .ZN(n1356) );
NAND3_X1 U1090 ( .A1(KEYINPUT29), .A2(n1234), .A3(n1360), .ZN(n1359) );
INV_X1 U1091 ( .A(G146), .ZN(n1234) );
OR2_X1 U1092 ( .A1(n1360), .A2(KEYINPUT29), .ZN(n1358) );
INV_X1 U1093 ( .A(n1273), .ZN(n1360) );
NAND2_X1 U1094 ( .A1(n1361), .A2(n1362), .ZN(n1273) );
NAND2_X1 U1095 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
INV_X1 U1096 ( .A(KEYINPUT52), .ZN(n1364) );
NAND2_X1 U1097 ( .A1(n1117), .A2(n1365), .ZN(n1363) );
NAND2_X1 U1098 ( .A1(G140), .A2(n1366), .ZN(n1365) );
NAND2_X1 U1099 ( .A1(G125), .A2(n1116), .ZN(n1117) );
INV_X1 U1100 ( .A(G140), .ZN(n1116) );
NAND2_X1 U1101 ( .A1(KEYINPUT52), .A2(n1367), .ZN(n1361) );
XOR2_X1 U1102 ( .A(n1366), .B(G140), .Z(n1367) );
INV_X1 U1103 ( .A(G125), .ZN(n1366) );
INV_X1 U1104 ( .A(G110), .ZN(n1175) );
endmodule


