//Key = 1101110011110101110010100100001001111101111010110010010010001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266;

XOR2_X1 U697 ( .A(G107), .B(n957), .Z(G9) );
NAND4_X1 U698 ( .A1(n958), .A2(n959), .A3(n960), .A4(n961), .ZN(G75) );
NAND4_X1 U699 ( .A1(n962), .A2(n963), .A3(n964), .A4(n965), .ZN(n960) );
NOR4_X1 U700 ( .A1(n966), .A2(n967), .A3(n968), .A4(n969), .ZN(n965) );
XNOR2_X1 U701 ( .A(KEYINPUT2), .B(n970), .ZN(n969) );
XNOR2_X1 U702 ( .A(n971), .B(n972), .ZN(n967) );
NOR2_X1 U703 ( .A1(G475), .A2(KEYINPUT59), .ZN(n972) );
XNOR2_X1 U704 ( .A(n973), .B(n974), .ZN(n966) );
NAND2_X1 U705 ( .A1(KEYINPUT40), .A2(n975), .ZN(n973) );
NOR3_X1 U706 ( .A1(n976), .A2(n977), .A3(n978), .ZN(n964) );
NAND2_X1 U707 ( .A1(n979), .A2(n980), .ZN(n963) );
NAND2_X1 U708 ( .A1(n981), .A2(n982), .ZN(n962) );
NAND2_X1 U709 ( .A1(n983), .A2(n984), .ZN(n959) );
NAND2_X1 U710 ( .A1(n985), .A2(n986), .ZN(n984) );
NAND4_X1 U711 ( .A1(n970), .A2(n987), .A3(n988), .A4(n989), .ZN(n986) );
NAND3_X1 U712 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n988) );
NAND2_X1 U713 ( .A1(n993), .A2(n994), .ZN(n992) );
NAND3_X1 U714 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n994) );
NAND2_X1 U715 ( .A1(n998), .A2(n999), .ZN(n996) );
OR3_X1 U716 ( .A1(n1000), .A2(n1001), .A3(n999), .ZN(n995) );
INV_X1 U717 ( .A(KEYINPUT13), .ZN(n999) );
NAND3_X1 U718 ( .A1(n1002), .A2(n1003), .A3(n998), .ZN(n991) );
NAND2_X1 U719 ( .A1(n1004), .A2(n1005), .ZN(n990) );
XNOR2_X1 U720 ( .A(KEYINPUT21), .B(n968), .ZN(n1005) );
NAND4_X1 U721 ( .A1(n998), .A2(n993), .A3(n1006), .A4(n1007), .ZN(n985) );
NAND2_X1 U722 ( .A1(n978), .A2(n1008), .ZN(n1007) );
NAND3_X1 U723 ( .A1(n987), .A2(n1009), .A3(n970), .ZN(n1008) );
INV_X1 U724 ( .A(n989), .ZN(n978) );
NAND2_X1 U725 ( .A1(n1010), .A2(n989), .ZN(n1006) );
NAND2_X1 U726 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND3_X1 U727 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NAND2_X1 U728 ( .A1(n987), .A2(n1016), .ZN(n1015) );
NAND2_X1 U729 ( .A1(n970), .A2(n1009), .ZN(n1016) );
INV_X1 U730 ( .A(KEYINPUT14), .ZN(n1009) );
NAND2_X1 U731 ( .A1(n1017), .A2(n1018), .ZN(n1011) );
INV_X1 U732 ( .A(n1019), .ZN(n983) );
XOR2_X1 U733 ( .A(n1020), .B(n1021), .Z(G72) );
NOR2_X1 U734 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
XNOR2_X1 U735 ( .A(n1024), .B(n1025), .ZN(n1023) );
XNOR2_X1 U736 ( .A(KEYINPUT58), .B(n1026), .ZN(n1025) );
NOR2_X1 U737 ( .A1(KEYINPUT61), .A2(n1027), .ZN(n1026) );
XNOR2_X1 U738 ( .A(n1028), .B(n1029), .ZN(n1027) );
NAND2_X1 U739 ( .A1(KEYINPUT60), .A2(n1030), .ZN(n1028) );
XOR2_X1 U740 ( .A(n1031), .B(n1032), .Z(n1030) );
XNOR2_X1 U741 ( .A(G131), .B(G137), .ZN(n1032) );
NAND2_X1 U742 ( .A1(KEYINPUT53), .A2(n1033), .ZN(n1031) );
NAND3_X1 U743 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1020) );
INV_X1 U744 ( .A(n1022), .ZN(n1035) );
OR2_X1 U745 ( .A1(n961), .A2(G227), .ZN(n1034) );
XOR2_X1 U746 ( .A(n1037), .B(n1038), .Z(G69) );
XOR2_X1 U747 ( .A(n1039), .B(n1040), .Z(n1038) );
NAND2_X1 U748 ( .A1(G953), .A2(n1041), .ZN(n1040) );
NAND2_X1 U749 ( .A1(G224), .A2(G898), .ZN(n1041) );
NAND3_X1 U750 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1039) );
NAND2_X1 U751 ( .A1(n1045), .A2(G953), .ZN(n1044) );
NAND2_X1 U752 ( .A1(KEYINPUT55), .A2(n1046), .ZN(n1043) );
NAND2_X1 U753 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
OR2_X1 U754 ( .A1(n1049), .A2(KEYINPUT55), .ZN(n1042) );
NOR2_X1 U755 ( .A1(n1050), .A2(G953), .ZN(n1037) );
NOR2_X1 U756 ( .A1(n1051), .A2(n1052), .ZN(G66) );
XNOR2_X1 U757 ( .A(n1053), .B(n1054), .ZN(n1052) );
NOR2_X1 U758 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U759 ( .A1(n1051), .A2(n1057), .ZN(G63) );
XOR2_X1 U760 ( .A(n1058), .B(n1059), .Z(n1057) );
NOR2_X1 U761 ( .A1(n1060), .A2(n1056), .ZN(n1058) );
NOR2_X1 U762 ( .A1(n1051), .A2(n1061), .ZN(G60) );
NOR3_X1 U763 ( .A1(n971), .A2(n1062), .A3(n1063), .ZN(n1061) );
NOR3_X1 U764 ( .A1(n1064), .A2(n1056), .A3(n1065), .ZN(n1063) );
NOR2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1062) );
NOR2_X1 U766 ( .A1(n958), .A2(n1065), .ZN(n1067) );
INV_X1 U767 ( .A(G475), .ZN(n1065) );
XNOR2_X1 U768 ( .A(G104), .B(n1068), .ZN(G6) );
NAND2_X1 U769 ( .A1(KEYINPUT1), .A2(n1069), .ZN(n1068) );
NOR2_X1 U770 ( .A1(n1051), .A2(n1070), .ZN(G57) );
XOR2_X1 U771 ( .A(n1071), .B(n1072), .Z(n1070) );
XOR2_X1 U772 ( .A(n1073), .B(n1074), .Z(n1072) );
XOR2_X1 U773 ( .A(n1075), .B(n1076), .Z(n1073) );
NOR2_X1 U774 ( .A1(KEYINPUT62), .A2(n1077), .ZN(n1076) );
INV_X1 U775 ( .A(G101), .ZN(n1077) );
XOR2_X1 U776 ( .A(n1078), .B(n1079), .Z(n1071) );
NOR2_X1 U777 ( .A1(n975), .A2(n1056), .ZN(n1079) );
XOR2_X1 U778 ( .A(n1080), .B(KEYINPUT18), .Z(n1078) );
NOR2_X1 U779 ( .A1(n1051), .A2(n1081), .ZN(G54) );
XOR2_X1 U780 ( .A(n1082), .B(n1083), .Z(n1081) );
XOR2_X1 U781 ( .A(n1084), .B(n1085), .Z(n1083) );
NOR3_X1 U782 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1085) );
AND2_X1 U783 ( .A1(KEYINPUT11), .A2(n1089), .ZN(n1088) );
NOR2_X1 U784 ( .A1(KEYINPUT11), .A2(n1090), .ZN(n1087) );
NAND3_X1 U785 ( .A1(n1091), .A2(n1092), .A3(G469), .ZN(n1084) );
NAND2_X1 U786 ( .A1(KEYINPUT36), .A2(n1056), .ZN(n1092) );
NAND2_X1 U787 ( .A1(G902), .A2(n1093), .ZN(n1056) );
NAND2_X1 U788 ( .A1(n1094), .A2(n1095), .ZN(n1091) );
INV_X1 U789 ( .A(KEYINPUT36), .ZN(n1095) );
NAND2_X1 U790 ( .A1(n958), .A2(G902), .ZN(n1094) );
INV_X1 U791 ( .A(n1093), .ZN(n958) );
NOR2_X1 U792 ( .A1(n1051), .A2(n1096), .ZN(G51) );
XOR2_X1 U793 ( .A(n1097), .B(n1098), .Z(n1096) );
XNOR2_X1 U794 ( .A(n1099), .B(n1049), .ZN(n1098) );
NOR3_X1 U795 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
NOR2_X1 U796 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U797 ( .A1(KEYINPUT45), .A2(n1105), .ZN(n1103) );
XOR2_X1 U798 ( .A(n1106), .B(KEYINPUT57), .Z(n1105) );
NOR3_X1 U799 ( .A1(G125), .A2(KEYINPUT45), .A3(n1106), .ZN(n1101) );
AND2_X1 U800 ( .A1(n1106), .A2(KEYINPUT45), .ZN(n1100) );
XOR2_X1 U801 ( .A(n1107), .B(n1108), .Z(n1097) );
XOR2_X1 U802 ( .A(KEYINPUT22), .B(n1109), .Z(n1108) );
NAND4_X1 U803 ( .A1(n1110), .A2(KEYINPUT5), .A3(n1111), .A4(n1093), .ZN(n1107) );
NAND2_X1 U804 ( .A1(n1050), .A2(n1036), .ZN(n1093) );
AND4_X1 U805 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1036) );
NOR4_X1 U806 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1115) );
INV_X1 U807 ( .A(n1120), .ZN(n1119) );
AND2_X1 U808 ( .A1(n1121), .A2(n1122), .ZN(n1114) );
NAND3_X1 U809 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1112) );
XNOR2_X1 U810 ( .A(KEYINPUT28), .B(n997), .ZN(n1124) );
AND2_X1 U811 ( .A1(n1126), .A2(n1127), .ZN(n1050) );
NOR4_X1 U812 ( .A1(n1128), .A2(n1129), .A3(n1069), .A4(n957), .ZN(n1127) );
AND3_X1 U813 ( .A1(n1123), .A2(n993), .A3(n1130), .ZN(n957) );
AND3_X1 U814 ( .A1(n1130), .A2(n993), .A3(n1131), .ZN(n1069) );
AND4_X1 U815 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1126) );
XNOR2_X1 U816 ( .A(G902), .B(KEYINPUT47), .ZN(n1110) );
NOR2_X1 U817 ( .A1(n961), .A2(G952), .ZN(n1051) );
XNOR2_X1 U818 ( .A(G146), .B(n1113), .ZN(G48) );
NAND3_X1 U819 ( .A1(n1131), .A2(n1136), .A3(n1125), .ZN(n1113) );
INV_X1 U820 ( .A(n1137), .ZN(n1125) );
XNOR2_X1 U821 ( .A(G143), .B(n1122), .ZN(G45) );
NAND4_X1 U822 ( .A1(n1138), .A2(n1139), .A3(n1136), .A4(n1140), .ZN(n1122) );
XOR2_X1 U823 ( .A(n1141), .B(G140), .Z(G42) );
NAND2_X1 U824 ( .A1(KEYINPUT35), .A2(n1121), .ZN(n1141) );
NAND3_X1 U825 ( .A1(n998), .A2(n1017), .A3(n1142), .ZN(n1121) );
XOR2_X1 U826 ( .A(G137), .B(n1118), .Z(G39) );
NOR3_X1 U827 ( .A1(n968), .A2(n1018), .A3(n1137), .ZN(n1118) );
INV_X1 U828 ( .A(n987), .ZN(n1018) );
XNOR2_X1 U829 ( .A(n1033), .B(n1117), .ZN(G36) );
AND3_X1 U830 ( .A1(n1139), .A2(n1123), .A3(n998), .ZN(n1117) );
XNOR2_X1 U831 ( .A(n1116), .B(n1143), .ZN(G33) );
NAND2_X1 U832 ( .A1(n1144), .A2(KEYINPUT9), .ZN(n1143) );
XNOR2_X1 U833 ( .A(G131), .B(KEYINPUT56), .ZN(n1144) );
AND3_X1 U834 ( .A1(n1139), .A2(n1131), .A3(n998), .ZN(n1116) );
INV_X1 U835 ( .A(n968), .ZN(n998) );
NAND2_X1 U836 ( .A1(n1145), .A2(n1000), .ZN(n968) );
INV_X1 U837 ( .A(n1001), .ZN(n1145) );
AND4_X1 U838 ( .A1(n1004), .A2(n1017), .A3(n1146), .A4(n989), .ZN(n1139) );
XNOR2_X1 U839 ( .A(n1147), .B(n1148), .ZN(G30) );
NOR4_X1 U840 ( .A1(KEYINPUT24), .A2(n997), .A3(n1013), .A4(n1137), .ZN(n1148) );
NAND3_X1 U841 ( .A1(n1149), .A2(n1017), .A3(n1150), .ZN(n1137) );
AND3_X1 U842 ( .A1(n1146), .A2(n989), .A3(n1151), .ZN(n1150) );
INV_X1 U843 ( .A(n1123), .ZN(n1013) );
INV_X1 U844 ( .A(n1136), .ZN(n997) );
NAND2_X1 U845 ( .A1(n1152), .A2(n1153), .ZN(G3) );
OR2_X1 U846 ( .A1(n1135), .A2(G101), .ZN(n1153) );
XOR2_X1 U847 ( .A(n1154), .B(KEYINPUT48), .Z(n1152) );
NAND2_X1 U848 ( .A1(G101), .A2(n1135), .ZN(n1154) );
NAND3_X1 U849 ( .A1(n987), .A2(n1130), .A3(n1004), .ZN(n1135) );
XOR2_X1 U850 ( .A(n1155), .B(n1156), .Z(G27) );
XNOR2_X1 U851 ( .A(KEYINPUT32), .B(n1104), .ZN(n1156) );
NOR2_X1 U852 ( .A1(KEYINPUT6), .A2(n1120), .ZN(n1155) );
NAND3_X1 U853 ( .A1(n970), .A2(n1136), .A3(n1142), .ZN(n1120) );
AND3_X1 U854 ( .A1(n1002), .A2(n1131), .A3(n1157), .ZN(n1142) );
AND3_X1 U855 ( .A1(n1003), .A2(n989), .A3(n1146), .ZN(n1157) );
NAND2_X1 U856 ( .A1(n1019), .A2(n1158), .ZN(n1146) );
NAND3_X1 U857 ( .A1(G902), .A2(n1159), .A3(n1022), .ZN(n1158) );
NOR2_X1 U858 ( .A1(G900), .A2(n961), .ZN(n1022) );
XNOR2_X1 U859 ( .A(G122), .B(n1134), .ZN(G24) );
NAND4_X1 U860 ( .A1(n1138), .A2(n1160), .A3(n993), .A4(n1140), .ZN(n1134) );
AND2_X1 U861 ( .A1(n1002), .A2(n1161), .ZN(n993) );
XNOR2_X1 U862 ( .A(KEYINPUT54), .B(n1151), .ZN(n1161) );
XOR2_X1 U863 ( .A(n1133), .B(n1162), .Z(G21) );
XOR2_X1 U864 ( .A(KEYINPUT39), .B(G119), .Z(n1162) );
NAND4_X1 U865 ( .A1(n1160), .A2(n987), .A3(n1149), .A4(n1151), .ZN(n1133) );
XNOR2_X1 U866 ( .A(n1132), .B(n1163), .ZN(G18) );
NOR2_X1 U867 ( .A1(KEYINPUT7), .A2(n1164), .ZN(n1163) );
NAND3_X1 U868 ( .A1(n1004), .A2(n1123), .A3(n1160), .ZN(n1132) );
AND4_X1 U869 ( .A1(n970), .A2(n1136), .A3(n1165), .A4(n989), .ZN(n1160) );
XNOR2_X1 U870 ( .A(n1166), .B(KEYINPUT38), .ZN(n1136) );
NAND2_X1 U871 ( .A1(n1001), .A2(n1000), .ZN(n1166) );
NOR2_X1 U872 ( .A1(n1138), .A2(n1167), .ZN(n1123) );
INV_X1 U873 ( .A(n1140), .ZN(n1167) );
XOR2_X1 U874 ( .A(G113), .B(n1129), .Z(G15) );
AND4_X1 U875 ( .A1(n1004), .A2(n1131), .A3(n970), .A4(n1168), .ZN(n1129) );
INV_X1 U876 ( .A(n1017), .ZN(n970) );
INV_X1 U877 ( .A(n1014), .ZN(n1131) );
NAND2_X1 U878 ( .A1(n1138), .A2(n1169), .ZN(n1014) );
XNOR2_X1 U879 ( .A(KEYINPUT12), .B(n1140), .ZN(n1169) );
NOR2_X1 U880 ( .A1(n1151), .A2(n1002), .ZN(n1004) );
NAND2_X1 U881 ( .A1(n1170), .A2(n1171), .ZN(G12) );
NAND2_X1 U882 ( .A1(n1128), .A2(n1172), .ZN(n1171) );
XOR2_X1 U883 ( .A(KEYINPUT50), .B(n1173), .Z(n1170) );
NOR2_X1 U884 ( .A1(n1128), .A2(n1172), .ZN(n1173) );
AND4_X1 U885 ( .A1(n987), .A2(n1130), .A3(n1002), .A4(n1003), .ZN(n1128) );
XNOR2_X1 U886 ( .A(n1151), .B(KEYINPUT16), .ZN(n1003) );
NAND3_X1 U887 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1151) );
INV_X1 U888 ( .A(n977), .ZN(n1176) );
NOR2_X1 U889 ( .A1(n982), .A2(n981), .ZN(n977) );
NAND2_X1 U890 ( .A1(KEYINPUT27), .A2(n1055), .ZN(n1175) );
NAND3_X1 U891 ( .A1(n982), .A2(n1177), .A3(n981), .ZN(n1174) );
INV_X1 U892 ( .A(n1055), .ZN(n981) );
NAND2_X1 U893 ( .A1(G217), .A2(n1178), .ZN(n1055) );
INV_X1 U894 ( .A(KEYINPUT27), .ZN(n1177) );
NAND2_X1 U895 ( .A1(n1053), .A2(n1179), .ZN(n982) );
XNOR2_X1 U896 ( .A(n1180), .B(n1181), .ZN(n1053) );
XOR2_X1 U897 ( .A(n1182), .B(n1183), .Z(n1181) );
XNOR2_X1 U898 ( .A(n1147), .B(G119), .ZN(n1183) );
XOR2_X1 U899 ( .A(G146), .B(G137), .Z(n1182) );
XOR2_X1 U900 ( .A(n1184), .B(n1185), .Z(n1180) );
XNOR2_X1 U901 ( .A(G110), .B(n1186), .ZN(n1185) );
NAND3_X1 U902 ( .A1(G234), .A2(n961), .A3(G221), .ZN(n1186) );
NAND2_X1 U903 ( .A1(KEYINPUT42), .A2(n1024), .ZN(n1184) );
INV_X1 U904 ( .A(n1149), .ZN(n1002) );
XOR2_X1 U905 ( .A(n974), .B(n975), .Z(n1149) );
INV_X1 U906 ( .A(G472), .ZN(n975) );
NAND2_X1 U907 ( .A1(n1187), .A2(n1179), .ZN(n974) );
XNOR2_X1 U908 ( .A(n1188), .B(n1189), .ZN(n1187) );
INV_X1 U909 ( .A(n1190), .ZN(n1189) );
XOR2_X1 U910 ( .A(n1075), .B(n1191), .Z(n1188) );
NOR2_X1 U911 ( .A1(KEYINPUT43), .A2(n1080), .ZN(n1191) );
NAND2_X1 U912 ( .A1(n1192), .A2(n1193), .ZN(n1080) );
XNOR2_X1 U913 ( .A(G210), .B(KEYINPUT8), .ZN(n1192) );
XOR2_X1 U914 ( .A(n1194), .B(n1195), .Z(n1075) );
XNOR2_X1 U915 ( .A(n1033), .B(G116), .ZN(n1195) );
XOR2_X1 U916 ( .A(n1196), .B(n1106), .Z(n1194) );
AND2_X1 U917 ( .A1(n1168), .A2(n1017), .ZN(n1130) );
XNOR2_X1 U918 ( .A(n1197), .B(G469), .ZN(n1017) );
NAND2_X1 U919 ( .A1(n1198), .A2(n1179), .ZN(n1197) );
XOR2_X1 U920 ( .A(n1082), .B(n1199), .Z(n1198) );
NOR2_X1 U921 ( .A1(n1089), .A2(n1086), .ZN(n1199) );
AND2_X1 U922 ( .A1(n1200), .A2(n1201), .ZN(n1086) );
NOR2_X1 U923 ( .A1(n1201), .A2(n1200), .ZN(n1089) );
INV_X1 U924 ( .A(n1090), .ZN(n1200) );
XOR2_X1 U925 ( .A(G140), .B(n1172), .Z(n1090) );
NAND2_X1 U926 ( .A1(G227), .A2(n961), .ZN(n1201) );
XOR2_X1 U927 ( .A(n1202), .B(n1203), .Z(n1082) );
XNOR2_X1 U928 ( .A(n1204), .B(n1205), .ZN(n1203) );
XOR2_X1 U929 ( .A(n1196), .B(n1206), .Z(n1205) );
XOR2_X1 U930 ( .A(G137), .B(n1207), .Z(n1196) );
NOR2_X1 U931 ( .A1(G131), .A2(n1208), .ZN(n1207) );
XNOR2_X1 U932 ( .A(KEYINPUT31), .B(KEYINPUT30), .ZN(n1208) );
INV_X1 U933 ( .A(n1029), .ZN(n1204) );
XNOR2_X1 U934 ( .A(n1209), .B(n1210), .ZN(n1029) );
NOR2_X1 U935 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XOR2_X1 U936 ( .A(n1213), .B(KEYINPUT17), .Z(n1212) );
NAND2_X1 U937 ( .A1(G146), .A2(n1214), .ZN(n1213) );
NOR2_X1 U938 ( .A1(G146), .A2(n1215), .ZN(n1211) );
XOR2_X1 U939 ( .A(KEYINPUT26), .B(n1214), .Z(n1215) );
XNOR2_X1 U940 ( .A(n1216), .B(KEYINPUT25), .ZN(n1214) );
NAND2_X1 U941 ( .A1(KEYINPUT4), .A2(n1147), .ZN(n1209) );
XNOR2_X1 U942 ( .A(G101), .B(n1217), .ZN(n1202) );
XNOR2_X1 U943 ( .A(KEYINPUT10), .B(n1218), .ZN(n1217) );
INV_X1 U944 ( .A(G104), .ZN(n1218) );
AND4_X1 U945 ( .A1(n1001), .A2(n1000), .A3(n1165), .A4(n989), .ZN(n1168) );
NAND2_X1 U946 ( .A1(n1219), .A2(n1178), .ZN(n989) );
NAND2_X1 U947 ( .A1(G234), .A2(n1179), .ZN(n1178) );
XNOR2_X1 U948 ( .A(G221), .B(KEYINPUT41), .ZN(n1219) );
NAND2_X1 U949 ( .A1(n1019), .A2(n1220), .ZN(n1165) );
NAND4_X1 U950 ( .A1(n1045), .A2(G953), .A3(G902), .A4(n1159), .ZN(n1220) );
XNOR2_X1 U951 ( .A(G898), .B(KEYINPUT23), .ZN(n1045) );
NAND3_X1 U952 ( .A1(n1159), .A2(n961), .A3(G952), .ZN(n1019) );
NAND2_X1 U953 ( .A1(G237), .A2(G234), .ZN(n1159) );
NAND2_X1 U954 ( .A1(G214), .A2(n1221), .ZN(n1000) );
XNOR2_X1 U955 ( .A(n1222), .B(n1111), .ZN(n1001) );
AND2_X1 U956 ( .A1(G210), .A2(n1221), .ZN(n1111) );
NAND2_X1 U957 ( .A1(n1223), .A2(n1179), .ZN(n1221) );
INV_X1 U958 ( .A(G237), .ZN(n1223) );
NAND2_X1 U959 ( .A1(n1224), .A2(n1179), .ZN(n1222) );
INV_X1 U960 ( .A(G902), .ZN(n1179) );
XOR2_X1 U961 ( .A(n1225), .B(n1226), .Z(n1224) );
XOR2_X1 U962 ( .A(n1106), .B(n1227), .Z(n1226) );
NOR2_X1 U963 ( .A1(KEYINPUT49), .A2(n1049), .ZN(n1227) );
XOR2_X1 U964 ( .A(n1047), .B(n1048), .Z(n1049) );
XNOR2_X1 U965 ( .A(n1172), .B(G122), .ZN(n1048) );
INV_X1 U966 ( .A(G110), .ZN(n1172) );
XNOR2_X1 U967 ( .A(n1190), .B(n1228), .ZN(n1047) );
XOR2_X1 U968 ( .A(n1229), .B(n1230), .Z(n1228) );
NAND2_X1 U969 ( .A1(KEYINPUT20), .A2(n1164), .ZN(n1230) );
NAND3_X1 U970 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1229) );
OR2_X1 U971 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U972 ( .A1(n1236), .A2(n1237), .ZN(n1232) );
INV_X1 U973 ( .A(KEYINPUT34), .ZN(n1237) );
NAND2_X1 U974 ( .A1(n1238), .A2(n1235), .ZN(n1236) );
XNOR2_X1 U975 ( .A(KEYINPUT44), .B(n1234), .ZN(n1238) );
NAND2_X1 U976 ( .A1(KEYINPUT34), .A2(n1239), .ZN(n1231) );
NAND2_X1 U977 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
OR2_X1 U978 ( .A1(n1234), .A2(KEYINPUT44), .ZN(n1241) );
NAND3_X1 U979 ( .A1(n1235), .A2(n1234), .A3(KEYINPUT44), .ZN(n1240) );
XOR2_X1 U980 ( .A(G104), .B(KEYINPUT63), .Z(n1234) );
XOR2_X1 U981 ( .A(G107), .B(KEYINPUT37), .Z(n1235) );
XOR2_X1 U982 ( .A(G101), .B(n1074), .Z(n1190) );
XOR2_X1 U983 ( .A(G113), .B(G119), .Z(n1074) );
XNOR2_X1 U984 ( .A(n1242), .B(n1147), .ZN(n1106) );
NAND2_X1 U985 ( .A1(KEYINPUT3), .A2(n1243), .ZN(n1242) );
XNOR2_X1 U986 ( .A(G125), .B(n1109), .ZN(n1225) );
AND2_X1 U987 ( .A1(G224), .A2(n961), .ZN(n1109) );
NOR2_X1 U988 ( .A1(n1140), .A2(n1138), .ZN(n987) );
XNOR2_X1 U989 ( .A(n971), .B(n1244), .ZN(n1138) );
NOR2_X1 U990 ( .A1(G475), .A2(KEYINPUT52), .ZN(n1244) );
NOR2_X1 U991 ( .A1(n1066), .A2(G902), .ZN(n971) );
INV_X1 U992 ( .A(n1064), .ZN(n1066) );
NAND2_X1 U993 ( .A1(n1245), .A2(n1246), .ZN(n1064) );
NAND2_X1 U994 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
XOR2_X1 U995 ( .A(KEYINPUT46), .B(n1249), .Z(n1245) );
NOR2_X1 U996 ( .A1(n1247), .A2(n1248), .ZN(n1249) );
XNOR2_X1 U997 ( .A(n1250), .B(n1251), .ZN(n1248) );
XOR2_X1 U998 ( .A(KEYINPUT15), .B(G122), .Z(n1251) );
XNOR2_X1 U999 ( .A(G113), .B(G104), .ZN(n1250) );
XNOR2_X1 U1000 ( .A(n1252), .B(n1253), .ZN(n1247) );
XOR2_X1 U1001 ( .A(n1024), .B(n1243), .Z(n1253) );
XNOR2_X1 U1002 ( .A(n1216), .B(G146), .ZN(n1243) );
XNOR2_X1 U1003 ( .A(G140), .B(n1104), .ZN(n1024) );
INV_X1 U1004 ( .A(G125), .ZN(n1104) );
XOR2_X1 U1005 ( .A(n1254), .B(G131), .Z(n1252) );
NAND2_X1 U1006 ( .A1(n1193), .A2(G214), .ZN(n1254) );
NOR2_X1 U1007 ( .A1(G953), .A2(G237), .ZN(n1193) );
NAND2_X1 U1008 ( .A1(n1255), .A2(n1256), .ZN(n1140) );
NAND2_X1 U1009 ( .A1(n1257), .A2(n980), .ZN(n1256) );
XNOR2_X1 U1010 ( .A(KEYINPUT0), .B(n979), .ZN(n1257) );
XNOR2_X1 U1011 ( .A(n976), .B(KEYINPUT29), .ZN(n1255) );
NOR2_X1 U1012 ( .A1(n980), .A2(n979), .ZN(n976) );
XOR2_X1 U1013 ( .A(n1060), .B(KEYINPUT33), .Z(n979) );
INV_X1 U1014 ( .A(G478), .ZN(n1060) );
OR2_X1 U1015 ( .A1(n1059), .A2(G902), .ZN(n980) );
XNOR2_X1 U1016 ( .A(n1258), .B(n1259), .ZN(n1059) );
XNOR2_X1 U1017 ( .A(n1260), .B(n1206), .ZN(n1259) );
XNOR2_X1 U1018 ( .A(G107), .B(n1033), .ZN(n1206) );
INV_X1 U1019 ( .A(G134), .ZN(n1033) );
NAND2_X1 U1020 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
NAND2_X1 U1021 ( .A1(G143), .A2(n1147), .ZN(n1262) );
INV_X1 U1022 ( .A(G128), .ZN(n1147) );
XOR2_X1 U1023 ( .A(n1263), .B(KEYINPUT51), .Z(n1261) );
NAND2_X1 U1024 ( .A1(G128), .A2(n1216), .ZN(n1263) );
INV_X1 U1025 ( .A(G143), .ZN(n1216) );
XOR2_X1 U1026 ( .A(n1264), .B(n1265), .Z(n1258) );
XNOR2_X1 U1027 ( .A(G122), .B(n1164), .ZN(n1265) );
INV_X1 U1028 ( .A(G116), .ZN(n1164) );
NAND3_X1 U1029 ( .A1(n1266), .A2(n961), .A3(G217), .ZN(n1264) );
INV_X1 U1030 ( .A(G953), .ZN(n961) );
XOR2_X1 U1031 ( .A(KEYINPUT19), .B(G234), .Z(n1266) );
endmodule


