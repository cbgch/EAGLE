//Key = 0011001111010111011111010111101100001111111100010100011001101110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399, n1400, n1401, n1402;

XNOR2_X1 U771 ( .A(G107), .B(n1058), .ZN(G9) );
NAND4_X1 U772 ( .A1(KEYINPUT15), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1058) );
NOR2_X1 U773 ( .A1(n1062), .A2(n1063), .ZN(G75) );
NOR4_X1 U774 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1063) );
XOR2_X1 U775 ( .A(KEYINPUT50), .B(n1068), .Z(n1065) );
NOR4_X1 U776 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1068) );
NAND3_X1 U777 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1069) );
XOR2_X1 U778 ( .A(n1076), .B(KEYINPUT27), .Z(n1075) );
NAND4_X1 U779 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1064) );
NAND3_X1 U780 ( .A1(n1074), .A2(n1081), .A3(KEYINPUT16), .ZN(n1078) );
NAND4_X1 U781 ( .A1(n1073), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1081) );
NAND2_X1 U782 ( .A1(n1073), .A2(n1085), .ZN(n1077) );
NAND2_X1 U783 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND3_X1 U784 ( .A1(n1061), .A2(n1088), .A3(n1074), .ZN(n1087) );
NAND2_X1 U785 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U786 ( .A1(n1082), .A2(n1091), .ZN(n1090) );
NAND2_X1 U787 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U788 ( .A1(n1094), .A2(n1083), .ZN(n1089) );
XNOR2_X1 U789 ( .A(n1095), .B(KEYINPUT25), .ZN(n1094) );
NAND3_X1 U790 ( .A1(n1083), .A2(n1096), .A3(n1082), .ZN(n1086) );
NAND2_X1 U791 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U792 ( .A1(n1074), .A2(n1099), .ZN(n1098) );
NAND2_X1 U793 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U794 ( .A1(n1084), .A2(n1102), .ZN(n1101) );
INV_X1 U795 ( .A(KEYINPUT16), .ZN(n1102) );
NAND2_X1 U796 ( .A1(n1061), .A2(n1103), .ZN(n1097) );
NAND2_X1 U797 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U798 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
INV_X1 U799 ( .A(n1108), .ZN(n1104) );
INV_X1 U800 ( .A(n1109), .ZN(n1073) );
AND3_X1 U801 ( .A1(n1079), .A2(n1080), .A3(n1110), .ZN(n1062) );
NAND4_X1 U802 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1079) );
NOR4_X1 U803 ( .A1(n1115), .A2(n1116), .A3(n1117), .A4(n1118), .ZN(n1114) );
NAND3_X1 U804 ( .A1(n1119), .A2(n1076), .A3(n1120), .ZN(n1115) );
NOR3_X1 U805 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1113) );
XOR2_X1 U806 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U807 ( .A(n1126), .B(KEYINPUT11), .Z(n1125) );
NAND2_X1 U808 ( .A1(KEYINPUT57), .A2(n1127), .ZN(n1124) );
XNOR2_X1 U809 ( .A(G469), .B(n1128), .ZN(n1122) );
XOR2_X1 U810 ( .A(KEYINPUT52), .B(n1129), .Z(n1121) );
XOR2_X1 U811 ( .A(KEYINPUT2), .B(n1130), .Z(n1112) );
NOR2_X1 U812 ( .A1(n1131), .A2(n1132), .ZN(n1111) );
AND2_X1 U813 ( .A1(n1133), .A2(G478), .ZN(n1132) );
NOR2_X1 U814 ( .A1(n1134), .A2(n1135), .ZN(n1131) );
XNOR2_X1 U815 ( .A(KEYINPUT38), .B(n1136), .ZN(n1135) );
XOR2_X1 U816 ( .A(n1137), .B(n1138), .Z(G72) );
NOR2_X1 U817 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U818 ( .A(n1141), .B(KEYINPUT39), .Z(n1140) );
NAND3_X1 U819 ( .A1(n1066), .A2(n1080), .A3(n1142), .ZN(n1141) );
NOR2_X1 U820 ( .A1(n1066), .A2(n1142), .ZN(n1139) );
NAND3_X1 U821 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1142) );
NAND2_X1 U822 ( .A1(G953), .A2(n1146), .ZN(n1145) );
NAND2_X1 U823 ( .A1(n1147), .A2(n1148), .ZN(n1144) );
NAND2_X1 U824 ( .A1(KEYINPUT43), .A2(n1149), .ZN(n1148) );
XOR2_X1 U825 ( .A(n1150), .B(n1151), .Z(n1147) );
NAND2_X1 U826 ( .A1(n1152), .A2(n1153), .ZN(n1150) );
NAND2_X1 U827 ( .A1(n1154), .A2(KEYINPUT47), .ZN(n1153) );
OR2_X1 U828 ( .A1(n1154), .A2(KEYINPUT13), .ZN(n1152) );
NAND3_X1 U829 ( .A1(KEYINPUT43), .A2(n1149), .A3(n1155), .ZN(n1143) );
XNOR2_X1 U830 ( .A(n1156), .B(n1151), .ZN(n1155) );
NAND2_X1 U831 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND2_X1 U832 ( .A1(n1154), .A2(KEYINPUT13), .ZN(n1158) );
OR2_X1 U833 ( .A1(n1154), .A2(KEYINPUT47), .ZN(n1157) );
NAND2_X1 U834 ( .A1(G953), .A2(n1159), .ZN(n1137) );
NAND2_X1 U835 ( .A1(G900), .A2(G227), .ZN(n1159) );
NAND2_X1 U836 ( .A1(n1160), .A2(n1161), .ZN(G69) );
NAND2_X1 U837 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U838 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
NAND2_X1 U839 ( .A1(G953), .A2(n1166), .ZN(n1165) );
INV_X1 U840 ( .A(n1167), .ZN(n1164) );
NAND2_X1 U841 ( .A1(n1168), .A2(n1169), .ZN(n1160) );
NAND2_X1 U842 ( .A1(G953), .A2(n1170), .ZN(n1169) );
NAND2_X1 U843 ( .A1(G898), .A2(G224), .ZN(n1170) );
INV_X1 U844 ( .A(n1163), .ZN(n1168) );
NAND2_X1 U845 ( .A1(KEYINPUT6), .A2(n1171), .ZN(n1163) );
XOR2_X1 U846 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U847 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XOR2_X1 U848 ( .A(n1080), .B(KEYINPUT36), .Z(n1175) );
INV_X1 U849 ( .A(n1067), .ZN(n1174) );
NOR2_X1 U850 ( .A1(n1167), .A2(n1176), .ZN(n1172) );
XOR2_X1 U851 ( .A(n1177), .B(n1178), .Z(n1176) );
NAND2_X1 U852 ( .A1(n1179), .A2(n1180), .ZN(n1177) );
NAND2_X1 U853 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U854 ( .A(n1183), .B(KEYINPUT10), .Z(n1179) );
OR2_X1 U855 ( .A1(n1181), .A2(n1182), .ZN(n1183) );
NOR2_X1 U856 ( .A1(n1184), .A2(n1185), .ZN(G66) );
XOR2_X1 U857 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U858 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NOR2_X1 U859 ( .A1(n1184), .A2(n1190), .ZN(G63) );
XOR2_X1 U860 ( .A(n1191), .B(n1192), .Z(n1190) );
NAND2_X1 U861 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NAND2_X1 U862 ( .A1(KEYINPUT26), .A2(n1195), .ZN(n1194) );
NAND2_X1 U863 ( .A1(KEYINPUT12), .A2(n1196), .ZN(n1193) );
INV_X1 U864 ( .A(n1195), .ZN(n1196) );
NAND2_X1 U865 ( .A1(n1197), .A2(G478), .ZN(n1195) );
NOR2_X1 U866 ( .A1(n1184), .A2(n1198), .ZN(G60) );
XOR2_X1 U867 ( .A(n1199), .B(n1200), .Z(n1198) );
AND2_X1 U868 ( .A1(G475), .A2(n1197), .ZN(n1200) );
XOR2_X1 U869 ( .A(G104), .B(n1201), .Z(G6) );
NOR2_X1 U870 ( .A1(n1184), .A2(n1202), .ZN(G57) );
XOR2_X1 U871 ( .A(n1203), .B(n1204), .Z(n1202) );
XOR2_X1 U872 ( .A(n1205), .B(n1206), .Z(n1204) );
NOR2_X1 U873 ( .A1(n1207), .A2(KEYINPUT55), .ZN(n1205) );
NOR2_X1 U874 ( .A1(n1127), .A2(n1189), .ZN(n1207) );
INV_X1 U875 ( .A(G472), .ZN(n1127) );
XOR2_X1 U876 ( .A(n1208), .B(KEYINPUT59), .Z(n1203) );
NAND4_X1 U877 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1208) );
OR3_X1 U878 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1212) );
NAND3_X1 U879 ( .A1(n1214), .A2(n1216), .A3(n1215), .ZN(n1211) );
XNOR2_X1 U880 ( .A(n1217), .B(KEYINPUT21), .ZN(n1214) );
NOR4_X1 U881 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(G54) );
AND2_X1 U882 ( .A1(KEYINPUT62), .A2(n1184), .ZN(n1221) );
NOR3_X1 U883 ( .A1(KEYINPUT62), .A2(n1080), .A3(n1110), .ZN(n1220) );
INV_X1 U884 ( .A(G952), .ZN(n1110) );
NOR2_X1 U885 ( .A1(n1222), .A2(n1223), .ZN(n1219) );
NOR2_X1 U886 ( .A1(n1224), .A2(n1225), .ZN(n1222) );
AND2_X1 U887 ( .A1(KEYINPUT1), .A2(n1226), .ZN(n1225) );
NOR2_X1 U888 ( .A1(KEYINPUT1), .A2(n1227), .ZN(n1224) );
AND2_X1 U889 ( .A1(n1223), .A2(n1227), .ZN(n1218) );
OR2_X1 U890 ( .A1(KEYINPUT51), .A2(n1226), .ZN(n1227) );
XNOR2_X1 U891 ( .A(n1228), .B(n1229), .ZN(n1226) );
XNOR2_X1 U892 ( .A(n1182), .B(n1154), .ZN(n1229) );
XNOR2_X1 U893 ( .A(n1230), .B(n1231), .ZN(n1154) );
XOR2_X1 U894 ( .A(n1232), .B(G131), .Z(n1228) );
NAND2_X1 U895 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND2_X1 U896 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XOR2_X1 U897 ( .A(KEYINPUT32), .B(n1237), .Z(n1236) );
NAND2_X1 U898 ( .A1(n1197), .A2(G469), .ZN(n1223) );
INV_X1 U899 ( .A(n1189), .ZN(n1197) );
NOR2_X1 U900 ( .A1(n1238), .A2(n1239), .ZN(G51) );
XOR2_X1 U901 ( .A(n1240), .B(n1241), .Z(n1239) );
XNOR2_X1 U902 ( .A(n1242), .B(n1243), .ZN(n1241) );
XOR2_X1 U903 ( .A(n1217), .B(n1244), .Z(n1243) );
NOR2_X1 U904 ( .A1(n1136), .A2(n1189), .ZN(n1244) );
NAND2_X1 U905 ( .A1(G902), .A2(n1245), .ZN(n1189) );
OR2_X1 U906 ( .A1(n1067), .A2(n1066), .ZN(n1245) );
NAND4_X1 U907 ( .A1(n1246), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1066) );
NOR4_X1 U908 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1249) );
AND2_X1 U909 ( .A1(n1254), .A2(n1255), .ZN(n1248) );
NAND2_X1 U910 ( .A1(n1256), .A2(n1257), .ZN(n1246) );
XOR2_X1 U911 ( .A(KEYINPUT22), .B(n1074), .Z(n1257) );
NAND4_X1 U912 ( .A1(n1258), .A2(n1259), .A3(n1260), .A4(n1261), .ZN(n1067) );
NOR4_X1 U913 ( .A1(n1201), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1261) );
INV_X1 U914 ( .A(n1265), .ZN(n1264) );
INV_X1 U915 ( .A(n1266), .ZN(n1263) );
NOR3_X1 U916 ( .A1(n1267), .A2(n1093), .A3(n1268), .ZN(n1262) );
XOR2_X1 U917 ( .A(KEYINPUT30), .B(n1061), .Z(n1267) );
NOR3_X1 U918 ( .A1(n1268), .A2(n1071), .A3(n1092), .ZN(n1201) );
NOR2_X1 U919 ( .A1(n1269), .A2(n1270), .ZN(n1260) );
NAND4_X1 U920 ( .A1(n1271), .A2(n1060), .A3(n1272), .A4(n1273), .ZN(n1258) );
OR2_X1 U921 ( .A1(n1274), .A2(KEYINPUT45), .ZN(n1273) );
NAND2_X1 U922 ( .A1(KEYINPUT45), .A2(n1275), .ZN(n1272) );
NAND3_X1 U923 ( .A1(n1082), .A2(n1108), .A3(n1276), .ZN(n1275) );
INV_X1 U924 ( .A(n1277), .ZN(n1276) );
XOR2_X1 U925 ( .A(n1278), .B(n1279), .Z(n1240) );
XOR2_X1 U926 ( .A(KEYINPUT40), .B(n1280), .Z(n1279) );
NOR2_X1 U927 ( .A1(G125), .A2(KEYINPUT56), .ZN(n1278) );
XNOR2_X1 U928 ( .A(n1184), .B(KEYINPUT49), .ZN(n1238) );
NOR2_X1 U929 ( .A1(n1080), .A2(G952), .ZN(n1184) );
XNOR2_X1 U930 ( .A(G146), .B(n1247), .ZN(G48) );
NAND3_X1 U931 ( .A1(n1281), .A2(n1108), .A3(n1282), .ZN(n1247) );
XOR2_X1 U932 ( .A(n1283), .B(n1255), .Z(G45) );
NAND4_X1 U933 ( .A1(n1284), .A2(n1108), .A3(n1285), .A4(n1286), .ZN(n1255) );
XNOR2_X1 U934 ( .A(G140), .B(n1287), .ZN(G42) );
NAND2_X1 U935 ( .A1(n1288), .A2(n1074), .ZN(n1287) );
XNOR2_X1 U936 ( .A(n1256), .B(KEYINPUT17), .ZN(n1288) );
AND2_X1 U937 ( .A1(n1289), .A2(n1095), .ZN(n1256) );
XOR2_X1 U938 ( .A(n1254), .B(n1290), .Z(G39) );
NAND2_X1 U939 ( .A1(KEYINPUT54), .A2(G137), .ZN(n1290) );
NAND3_X1 U940 ( .A1(n1282), .A2(n1083), .A3(n1074), .ZN(n1254) );
XOR2_X1 U941 ( .A(G134), .B(n1253), .Z(G36) );
AND3_X1 U942 ( .A1(n1284), .A2(n1060), .A3(n1074), .ZN(n1253) );
XOR2_X1 U943 ( .A(G131), .B(n1252), .Z(G33) );
AND3_X1 U944 ( .A1(n1284), .A2(n1281), .A3(n1074), .ZN(n1252) );
AND2_X1 U945 ( .A1(n1107), .A2(n1119), .ZN(n1074) );
AND3_X1 U946 ( .A1(n1095), .A2(n1291), .A3(n1271), .ZN(n1284) );
XOR2_X1 U947 ( .A(G128), .B(n1251), .Z(G30) );
AND3_X1 U948 ( .A1(n1060), .A2(n1108), .A3(n1282), .ZN(n1251) );
AND4_X1 U949 ( .A1(n1292), .A2(n1095), .A3(n1293), .A4(n1291), .ZN(n1282) );
INV_X1 U950 ( .A(n1093), .ZN(n1060) );
XNOR2_X1 U951 ( .A(G101), .B(n1259), .ZN(G3) );
NAND3_X1 U952 ( .A1(n1083), .A2(n1059), .A3(n1271), .ZN(n1259) );
INV_X1 U953 ( .A(n1100), .ZN(n1271) );
XOR2_X1 U954 ( .A(G125), .B(n1250), .Z(G27) );
AND3_X1 U955 ( .A1(n1082), .A2(n1108), .A3(n1289), .ZN(n1250) );
AND3_X1 U956 ( .A1(n1084), .A2(n1291), .A3(n1281), .ZN(n1289) );
INV_X1 U957 ( .A(n1092), .ZN(n1281) );
NAND2_X1 U958 ( .A1(n1109), .A2(n1294), .ZN(n1291) );
NAND4_X1 U959 ( .A1(G902), .A2(G953), .A3(n1295), .A4(n1146), .ZN(n1294) );
INV_X1 U960 ( .A(G900), .ZN(n1146) );
XOR2_X1 U961 ( .A(n1296), .B(n1265), .Z(G24) );
NAND4_X1 U962 ( .A1(n1274), .A2(n1061), .A3(n1285), .A4(n1286), .ZN(n1265) );
INV_X1 U963 ( .A(n1071), .ZN(n1061) );
NAND2_X1 U964 ( .A1(n1297), .A2(n1298), .ZN(n1071) );
XOR2_X1 U965 ( .A(n1299), .B(n1266), .Z(G21) );
NAND4_X1 U966 ( .A1(n1292), .A2(n1274), .A3(n1083), .A4(n1293), .ZN(n1266) );
INV_X1 U967 ( .A(n1300), .ZN(n1274) );
XOR2_X1 U968 ( .A(G116), .B(n1301), .Z(G18) );
NOR3_X1 U969 ( .A1(n1100), .A2(n1093), .A3(n1300), .ZN(n1301) );
NAND2_X1 U970 ( .A1(n1302), .A2(n1285), .ZN(n1093) );
XOR2_X1 U971 ( .A(G113), .B(n1270), .Z(G15) );
NOR3_X1 U972 ( .A1(n1100), .A2(n1300), .A3(n1092), .ZN(n1270) );
NAND2_X1 U973 ( .A1(n1303), .A2(n1286), .ZN(n1092) );
INV_X1 U974 ( .A(n1302), .ZN(n1286) );
NAND3_X1 U975 ( .A1(n1108), .A2(n1277), .A3(n1082), .ZN(n1300) );
NOR2_X1 U976 ( .A1(n1070), .A2(n1304), .ZN(n1082) );
NAND2_X1 U977 ( .A1(n1292), .A2(n1297), .ZN(n1100) );
XOR2_X1 U978 ( .A(n1298), .B(KEYINPUT28), .Z(n1292) );
XOR2_X1 U979 ( .A(G110), .B(n1269), .Z(G12) );
AND3_X1 U980 ( .A1(n1084), .A2(n1059), .A3(n1083), .ZN(n1269) );
INV_X1 U981 ( .A(n1072), .ZN(n1083) );
NAND2_X1 U982 ( .A1(n1302), .A2(n1303), .ZN(n1072) );
XNOR2_X1 U983 ( .A(KEYINPUT5), .B(n1285), .ZN(n1303) );
NAND3_X1 U984 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1285) );
INV_X1 U985 ( .A(n1116), .ZN(n1307) );
NOR2_X1 U986 ( .A1(n1133), .A2(G478), .ZN(n1116) );
OR2_X1 U987 ( .A1(G478), .A2(KEYINPUT7), .ZN(n1306) );
NAND3_X1 U988 ( .A1(G478), .A2(n1133), .A3(KEYINPUT7), .ZN(n1305) );
NAND2_X1 U989 ( .A1(n1308), .A2(n1191), .ZN(n1133) );
NAND2_X1 U990 ( .A1(n1309), .A2(n1310), .ZN(n1191) );
NAND2_X1 U991 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U992 ( .A(KEYINPUT37), .B(n1313), .Z(n1309) );
NOR2_X1 U993 ( .A1(n1311), .A2(n1312), .ZN(n1313) );
NAND3_X1 U994 ( .A1(n1314), .A2(G234), .A3(G217), .ZN(n1312) );
XOR2_X1 U995 ( .A(n1315), .B(n1316), .Z(n1311) );
XOR2_X1 U996 ( .A(G128), .B(n1317), .Z(n1316) );
NOR2_X1 U997 ( .A1(KEYINPUT63), .A2(n1318), .ZN(n1317) );
XNOR2_X1 U998 ( .A(G107), .B(n1319), .ZN(n1318) );
NAND2_X1 U999 ( .A1(KEYINPUT19), .A2(n1320), .ZN(n1319) );
XOR2_X1 U1000 ( .A(G122), .B(G116), .Z(n1320) );
XOR2_X1 U1001 ( .A(G134), .B(n1283), .Z(n1315) );
NOR2_X1 U1002 ( .A1(n1321), .A2(n1118), .ZN(n1302) );
NOR3_X1 U1003 ( .A1(G475), .A2(G902), .A3(n1199), .ZN(n1118) );
XOR2_X1 U1004 ( .A(n1117), .B(KEYINPUT35), .Z(n1321) );
AND2_X1 U1005 ( .A1(G475), .A2(n1322), .ZN(n1117) );
NAND2_X1 U1006 ( .A1(n1323), .A2(n1308), .ZN(n1322) );
INV_X1 U1007 ( .A(n1199), .ZN(n1323) );
XOR2_X1 U1008 ( .A(n1324), .B(n1325), .Z(n1199) );
XNOR2_X1 U1009 ( .A(n1326), .B(n1151), .ZN(n1325) );
NAND2_X1 U1010 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
NAND2_X1 U1011 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XOR2_X1 U1012 ( .A(KEYINPUT20), .B(n1331), .Z(n1327) );
NOR2_X1 U1013 ( .A1(n1329), .A2(n1330), .ZN(n1331) );
XNOR2_X1 U1014 ( .A(G113), .B(n1332), .ZN(n1329) );
NOR2_X1 U1015 ( .A1(KEYINPUT48), .A2(n1296), .ZN(n1332) );
INV_X1 U1016 ( .A(G122), .ZN(n1296) );
XOR2_X1 U1017 ( .A(n1333), .B(n1334), .Z(n1324) );
NOR2_X1 U1018 ( .A1(KEYINPUT46), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1019 ( .A(n1336), .B(G143), .Z(n1335) );
NAND2_X1 U1020 ( .A1(n1337), .A2(G214), .ZN(n1336) );
XOR2_X1 U1021 ( .A(G146), .B(n1149), .Z(n1333) );
INV_X1 U1022 ( .A(n1268), .ZN(n1059) );
NAND3_X1 U1023 ( .A1(n1108), .A2(n1277), .A3(n1095), .ZN(n1268) );
NOR2_X1 U1024 ( .A1(n1304), .A2(n1338), .ZN(n1095) );
INV_X1 U1025 ( .A(n1070), .ZN(n1338) );
XOR2_X1 U1026 ( .A(G469), .B(n1339), .Z(n1070) );
NOR2_X1 U1027 ( .A1(KEYINPUT34), .A2(n1128), .ZN(n1339) );
NAND2_X1 U1028 ( .A1(n1340), .A2(n1308), .ZN(n1128) );
XOR2_X1 U1029 ( .A(n1341), .B(n1342), .Z(n1340) );
NAND2_X1 U1030 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
NAND2_X1 U1031 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
NAND2_X1 U1032 ( .A1(KEYINPUT61), .A2(n1347), .ZN(n1346) );
NAND2_X1 U1033 ( .A1(KEYINPUT41), .A2(n1213), .ZN(n1347) );
INV_X1 U1034 ( .A(n1348), .ZN(n1345) );
NAND2_X1 U1035 ( .A1(n1216), .A2(n1349), .ZN(n1343) );
NAND2_X1 U1036 ( .A1(KEYINPUT41), .A2(n1350), .ZN(n1349) );
NAND2_X1 U1037 ( .A1(n1348), .A2(KEYINPUT61), .ZN(n1350) );
XOR2_X1 U1038 ( .A(n1182), .B(n1231), .Z(n1348) );
XNOR2_X1 U1039 ( .A(n1351), .B(G128), .ZN(n1231) );
NAND2_X1 U1040 ( .A1(n1352), .A2(KEYINPUT42), .ZN(n1351) );
XOR2_X1 U1041 ( .A(n1283), .B(n1353), .Z(n1352) );
XOR2_X1 U1042 ( .A(KEYINPUT4), .B(G146), .Z(n1353) );
NAND2_X1 U1043 ( .A1(n1354), .A2(n1355), .ZN(n1341) );
NAND2_X1 U1044 ( .A1(n1237), .A2(n1235), .ZN(n1355) );
XNOR2_X1 U1045 ( .A(KEYINPUT60), .B(n1233), .ZN(n1354) );
OR2_X1 U1046 ( .A1(n1235), .A2(n1237), .ZN(n1233) );
AND2_X1 U1047 ( .A1(G227), .A2(n1314), .ZN(n1237) );
XOR2_X1 U1048 ( .A(G140), .B(n1356), .Z(n1235) );
XOR2_X1 U1049 ( .A(n1076), .B(KEYINPUT3), .Z(n1304) );
NAND2_X1 U1050 ( .A1(G221), .A2(n1357), .ZN(n1076) );
NAND2_X1 U1051 ( .A1(n1109), .A2(n1358), .ZN(n1277) );
NAND3_X1 U1052 ( .A1(n1167), .A2(n1295), .A3(G902), .ZN(n1358) );
NOR2_X1 U1053 ( .A1(n1080), .A2(G898), .ZN(n1167) );
NAND3_X1 U1054 ( .A1(n1295), .A2(n1080), .A3(G952), .ZN(n1109) );
NAND2_X1 U1055 ( .A1(G237), .A2(G234), .ZN(n1295) );
NOR2_X1 U1056 ( .A1(n1106), .A2(n1107), .ZN(n1108) );
NOR2_X1 U1057 ( .A1(n1359), .A2(n1130), .ZN(n1107) );
AND2_X1 U1058 ( .A1(n1134), .A2(n1136), .ZN(n1130) );
INV_X1 U1059 ( .A(n1360), .ZN(n1134) );
AND2_X1 U1060 ( .A1(n1361), .A2(n1360), .ZN(n1359) );
NAND3_X1 U1061 ( .A1(n1362), .A2(n1308), .A3(n1363), .ZN(n1360) );
XOR2_X1 U1062 ( .A(n1364), .B(KEYINPUT29), .Z(n1363) );
NAND2_X1 U1063 ( .A1(n1365), .A2(n1242), .ZN(n1364) );
OR2_X1 U1064 ( .A1(n1242), .A2(n1365), .ZN(n1362) );
XNOR2_X1 U1065 ( .A(n1366), .B(n1367), .ZN(n1365) );
XOR2_X1 U1066 ( .A(G125), .B(n1280), .Z(n1367) );
NOR2_X1 U1067 ( .A1(n1166), .A2(n1368), .ZN(n1280) );
INV_X1 U1068 ( .A(G224), .ZN(n1166) );
NAND2_X1 U1069 ( .A1(KEYINPUT8), .A2(n1217), .ZN(n1366) );
XNOR2_X1 U1070 ( .A(n1369), .B(n1178), .ZN(n1242) );
XOR2_X1 U1071 ( .A(G110), .B(n1370), .Z(n1178) );
XOR2_X1 U1072 ( .A(KEYINPUT58), .B(G122), .Z(n1370) );
NAND3_X1 U1073 ( .A1(n1371), .A2(n1372), .A3(n1373), .ZN(n1369) );
NAND2_X1 U1074 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
NAND2_X1 U1075 ( .A1(n1376), .A2(KEYINPUT9), .ZN(n1375) );
XOR2_X1 U1076 ( .A(n1182), .B(KEYINPUT24), .Z(n1376) );
INV_X1 U1077 ( .A(n1181), .ZN(n1374) );
NAND3_X1 U1078 ( .A1(KEYINPUT9), .A2(n1181), .A3(n1182), .ZN(n1372) );
XNOR2_X1 U1079 ( .A(G113), .B(n1377), .ZN(n1181) );
NOR2_X1 U1080 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
XOR2_X1 U1081 ( .A(n1380), .B(KEYINPUT31), .Z(n1379) );
NAND2_X1 U1082 ( .A1(n1381), .A2(n1299), .ZN(n1380) );
XOR2_X1 U1083 ( .A(KEYINPUT33), .B(G116), .Z(n1381) );
NOR2_X1 U1084 ( .A1(G116), .A2(n1299), .ZN(n1378) );
INV_X1 U1085 ( .A(G119), .ZN(n1299) );
OR2_X1 U1086 ( .A1(n1182), .A2(KEYINPUT9), .ZN(n1371) );
XOR2_X1 U1087 ( .A(n1382), .B(n1383), .Z(n1182) );
XOR2_X1 U1088 ( .A(G107), .B(n1330), .Z(n1382) );
INV_X1 U1089 ( .A(G104), .ZN(n1330) );
XOR2_X1 U1090 ( .A(n1136), .B(KEYINPUT23), .Z(n1361) );
NAND2_X1 U1091 ( .A1(G210), .A2(n1384), .ZN(n1136) );
INV_X1 U1092 ( .A(n1119), .ZN(n1106) );
NAND2_X1 U1093 ( .A1(G214), .A2(n1384), .ZN(n1119) );
NAND2_X1 U1094 ( .A1(n1385), .A2(n1308), .ZN(n1384) );
INV_X1 U1095 ( .A(G237), .ZN(n1385) );
AND2_X1 U1096 ( .A1(n1298), .A2(n1293), .ZN(n1084) );
XOR2_X1 U1097 ( .A(n1297), .B(KEYINPUT18), .Z(n1293) );
NOR2_X1 U1098 ( .A1(n1386), .A2(n1129), .ZN(n1297) );
NOR2_X1 U1099 ( .A1(n1188), .A2(n1387), .ZN(n1129) );
XOR2_X1 U1100 ( .A(KEYINPUT53), .B(n1120), .Z(n1386) );
NAND2_X1 U1101 ( .A1(n1387), .A2(n1188), .ZN(n1120) );
NAND2_X1 U1102 ( .A1(G217), .A2(n1357), .ZN(n1188) );
NAND2_X1 U1103 ( .A1(G234), .A2(n1308), .ZN(n1357) );
NOR2_X1 U1104 ( .A1(n1186), .A2(G902), .ZN(n1387) );
XOR2_X1 U1105 ( .A(n1388), .B(n1389), .Z(n1186) );
XNOR2_X1 U1106 ( .A(n1151), .B(n1390), .ZN(n1389) );
XNOR2_X1 U1107 ( .A(n1391), .B(n1392), .ZN(n1390) );
AND3_X1 U1108 ( .A1(G221), .A2(G234), .A3(n1314), .ZN(n1392) );
XOR2_X1 U1109 ( .A(G140), .B(G125), .Z(n1151) );
XOR2_X1 U1110 ( .A(n1356), .B(n1393), .Z(n1388) );
XOR2_X1 U1111 ( .A(G137), .B(G119), .Z(n1393) );
INV_X1 U1112 ( .A(G110), .ZN(n1356) );
XOR2_X1 U1113 ( .A(n1126), .B(n1394), .Z(n1298) );
XOR2_X1 U1114 ( .A(KEYINPUT44), .B(G472), .Z(n1394) );
NAND2_X1 U1115 ( .A1(n1395), .A2(n1308), .ZN(n1126) );
INV_X1 U1116 ( .A(G902), .ZN(n1308) );
XOR2_X1 U1117 ( .A(n1396), .B(n1206), .Z(n1395) );
XNOR2_X1 U1118 ( .A(n1397), .B(n1383), .ZN(n1206) );
XOR2_X1 U1119 ( .A(G101), .B(KEYINPUT14), .Z(n1383) );
NAND2_X1 U1120 ( .A1(n1337), .A2(G210), .ZN(n1397) );
NOR2_X1 U1121 ( .A1(n1368), .A2(G237), .ZN(n1337) );
INV_X1 U1122 ( .A(n1314), .ZN(n1368) );
XOR2_X1 U1123 ( .A(n1080), .B(KEYINPUT0), .Z(n1314) );
INV_X1 U1124 ( .A(G953), .ZN(n1080) );
NAND3_X1 U1125 ( .A1(n1209), .A2(n1210), .A3(n1398), .ZN(n1396) );
NAND2_X1 U1126 ( .A1(n1399), .A2(n1216), .ZN(n1398) );
XOR2_X1 U1127 ( .A(n1215), .B(n1400), .Z(n1399) );
NAND3_X1 U1128 ( .A1(n1400), .A2(n1215), .A3(n1213), .ZN(n1210) );
INV_X1 U1129 ( .A(n1216), .ZN(n1213) );
OR3_X1 U1130 ( .A1(n1216), .A2(n1400), .A3(n1215), .ZN(n1209) );
XOR2_X1 U1131 ( .A(G113), .B(n1401), .Z(n1215) );
XOR2_X1 U1132 ( .A(G119), .B(G116), .Z(n1401) );
INV_X1 U1133 ( .A(n1217), .ZN(n1400) );
XOR2_X1 U1134 ( .A(n1283), .B(n1391), .Z(n1217) );
XOR2_X1 U1135 ( .A(G128), .B(G146), .Z(n1391) );
INV_X1 U1136 ( .A(G143), .ZN(n1283) );
XNOR2_X1 U1137 ( .A(n1149), .B(n1402), .ZN(n1216) );
INV_X1 U1138 ( .A(n1230), .ZN(n1402) );
XNOR2_X1 U1139 ( .A(G134), .B(G137), .ZN(n1230) );
INV_X1 U1140 ( .A(G131), .ZN(n1149) );
endmodule


