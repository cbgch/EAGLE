//Key = 1100111000010111011001001111111111010000100110101110100011110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325;

XOR2_X1 U732 ( .A(G107), .B(n1000), .Z(G9) );
NAND4_X1 U733 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(G75) );
NAND3_X1 U734 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n1004) );
NAND2_X1 U735 ( .A1(G952), .A2(n1008), .ZN(n1003) );
NAND3_X1 U736 ( .A1(n1009), .A2(n1005), .A3(n1010), .ZN(n1008) );
NAND2_X1 U737 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NAND2_X1 U738 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND3_X1 U739 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NAND3_X1 U740 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1016) );
NAND2_X1 U741 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
XNOR2_X1 U742 ( .A(n1023), .B(KEYINPUT15), .ZN(n1021) );
NAND2_X1 U743 ( .A1(n1023), .A2(n1024), .ZN(n1019) );
NAND2_X1 U744 ( .A1(n1025), .A2(n1026), .ZN(n1018) );
NAND2_X1 U745 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U746 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND3_X1 U747 ( .A1(n1031), .A2(n1032), .A3(n1023), .ZN(n1013) );
NAND2_X1 U748 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U749 ( .A1(KEYINPUT62), .A2(n1035), .ZN(n1033) );
NAND4_X1 U750 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1025), .ZN(n1031) );
NAND2_X1 U751 ( .A1(n1015), .A2(n1039), .ZN(n1038) );
NAND2_X1 U752 ( .A1(n1017), .A2(n1040), .ZN(n1037) );
NAND2_X1 U753 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U754 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U755 ( .A1(n1035), .A2(n1045), .ZN(n1036) );
INV_X1 U756 ( .A(KEYINPUT62), .ZN(n1045) );
XOR2_X1 U757 ( .A(n1046), .B(KEYINPUT20), .Z(n1011) );
OR2_X1 U758 ( .A1(n1006), .A2(n1005), .ZN(n1001) );
NAND4_X1 U759 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1005) );
NOR4_X1 U760 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1050) );
NOR3_X1 U761 ( .A1(n1055), .A2(KEYINPUT3), .A3(n1056), .ZN(n1052) );
AND2_X1 U762 ( .A1(n1055), .A2(KEYINPUT3), .ZN(n1051) );
XOR2_X1 U763 ( .A(KEYINPUT55), .B(n1057), .Z(n1047) );
NOR3_X1 U764 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
XOR2_X1 U765 ( .A(KEYINPUT10), .B(n1061), .Z(n1060) );
NOR2_X1 U766 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
XOR2_X1 U767 ( .A(n1064), .B(KEYINPUT40), .Z(n1059) );
NAND3_X1 U768 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1058) );
NAND2_X1 U769 ( .A1(n1063), .A2(n1062), .ZN(n1067) );
XNOR2_X1 U770 ( .A(n1068), .B(KEYINPUT19), .ZN(n1063) );
INV_X1 U771 ( .A(KEYINPUT28), .ZN(n1006) );
XOR2_X1 U772 ( .A(n1069), .B(n1070), .Z(G72) );
XOR2_X1 U773 ( .A(n1071), .B(n1072), .Z(n1070) );
NOR2_X1 U774 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XNOR2_X1 U775 ( .A(G953), .B(KEYINPUT30), .ZN(n1074) );
INV_X1 U776 ( .A(n1075), .ZN(n1073) );
NOR2_X1 U777 ( .A1(n1076), .A2(n1077), .ZN(n1071) );
XOR2_X1 U778 ( .A(n1078), .B(n1079), .Z(n1077) );
XNOR2_X1 U779 ( .A(n1080), .B(n1081), .ZN(n1079) );
XNOR2_X1 U780 ( .A(n1082), .B(n1083), .ZN(n1078) );
NAND4_X1 U781 ( .A1(KEYINPUT49), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1082) );
NAND2_X1 U782 ( .A1(KEYINPUT34), .A2(n1087), .ZN(n1086) );
NAND2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XNOR2_X1 U784 ( .A(KEYINPUT12), .B(n1090), .ZN(n1088) );
NAND2_X1 U785 ( .A1(n1091), .A2(n1092), .ZN(n1085) );
INV_X1 U786 ( .A(KEYINPUT34), .ZN(n1092) );
NAND2_X1 U787 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
OR3_X1 U788 ( .A1(n1090), .A2(G134), .A3(KEYINPUT12), .ZN(n1094) );
NAND2_X1 U789 ( .A1(KEYINPUT12), .A2(n1090), .ZN(n1093) );
NAND2_X1 U790 ( .A1(G134), .A2(n1090), .ZN(n1084) );
NOR2_X1 U791 ( .A1(G900), .A2(n1095), .ZN(n1076) );
XNOR2_X1 U792 ( .A(KEYINPUT31), .B(n1002), .ZN(n1095) );
NOR2_X1 U793 ( .A1(n1096), .A2(n1002), .ZN(n1069) );
NOR2_X1 U794 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U795 ( .A1(n1099), .A2(n1100), .ZN(G69) );
NAND2_X1 U796 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U797 ( .A1(n1103), .A2(n1104), .ZN(n1099) );
NAND2_X1 U798 ( .A1(n1105), .A2(n1102), .ZN(n1104) );
NAND2_X1 U799 ( .A1(G953), .A2(n1106), .ZN(n1102) );
INV_X1 U800 ( .A(G224), .ZN(n1106) );
INV_X1 U801 ( .A(n1101), .ZN(n1103) );
XNOR2_X1 U802 ( .A(n1107), .B(n1108), .ZN(n1101) );
NOR2_X1 U803 ( .A1(G953), .A2(n1109), .ZN(n1108) );
XOR2_X1 U804 ( .A(KEYINPUT36), .B(n1110), .Z(n1109) );
NOR2_X1 U805 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XNOR2_X1 U806 ( .A(n1113), .B(KEYINPUT46), .ZN(n1111) );
NAND2_X1 U807 ( .A1(n1114), .A2(n1105), .ZN(n1107) );
INV_X1 U808 ( .A(n1115), .ZN(n1105) );
XOR2_X1 U809 ( .A(n1116), .B(n1117), .Z(n1114) );
XOR2_X1 U810 ( .A(KEYINPUT50), .B(n1118), .Z(n1117) );
NOR2_X1 U811 ( .A1(KEYINPUT38), .A2(n1119), .ZN(n1118) );
NOR2_X1 U812 ( .A1(n1120), .A2(n1121), .ZN(G66) );
XOR2_X1 U813 ( .A(n1122), .B(n1123), .Z(n1121) );
NAND2_X1 U814 ( .A1(KEYINPUT59), .A2(n1124), .ZN(n1123) );
NAND2_X1 U815 ( .A1(n1125), .A2(n1126), .ZN(n1122) );
NOR3_X1 U816 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(G63) );
NOR3_X1 U817 ( .A1(n1130), .A2(n1002), .A3(n1007), .ZN(n1129) );
INV_X1 U818 ( .A(G952), .ZN(n1007) );
AND2_X1 U819 ( .A1(n1130), .A2(n1120), .ZN(n1128) );
INV_X1 U820 ( .A(KEYINPUT45), .ZN(n1130) );
XOR2_X1 U821 ( .A(n1131), .B(n1132), .Z(n1127) );
NOR2_X1 U822 ( .A1(KEYINPUT9), .A2(n1133), .ZN(n1132) );
AND2_X1 U823 ( .A1(G478), .A2(n1125), .ZN(n1131) );
NOR2_X1 U824 ( .A1(n1120), .A2(n1134), .ZN(G60) );
XOR2_X1 U825 ( .A(n1135), .B(n1136), .Z(n1134) );
NAND3_X1 U826 ( .A1(n1125), .A2(G475), .A3(KEYINPUT21), .ZN(n1135) );
XNOR2_X1 U827 ( .A(n1137), .B(n1113), .ZN(G6) );
NOR2_X1 U828 ( .A1(n1120), .A2(n1138), .ZN(G57) );
XOR2_X1 U829 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U830 ( .A(n1141), .B(n1142), .Z(n1140) );
AND2_X1 U831 ( .A1(G472), .A2(n1125), .ZN(n1142) );
NOR2_X1 U832 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
XNOR2_X1 U833 ( .A(n1145), .B(KEYINPUT11), .ZN(n1144) );
NOR2_X1 U834 ( .A1(n1120), .A2(n1146), .ZN(G54) );
XOR2_X1 U835 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U836 ( .A(n1149), .B(n1150), .Z(n1148) );
AND2_X1 U837 ( .A1(G469), .A2(n1125), .ZN(n1149) );
XOR2_X1 U838 ( .A(n1151), .B(G146), .Z(n1147) );
NAND2_X1 U839 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND4_X1 U840 ( .A1(n1154), .A2(KEYINPUT24), .A3(n1155), .A4(n1156), .ZN(n1153) );
NAND2_X1 U841 ( .A1(n1157), .A2(n1158), .ZN(n1152) );
NAND2_X1 U842 ( .A1(n1155), .A2(n1159), .ZN(n1158) );
OR2_X1 U843 ( .A1(n1156), .A2(n1154), .ZN(n1159) );
INV_X1 U844 ( .A(KEYINPUT53), .ZN(n1156) );
NAND2_X1 U845 ( .A1(KEYINPUT24), .A2(n1154), .ZN(n1157) );
XOR2_X1 U846 ( .A(n1160), .B(G140), .Z(n1154) );
NAND2_X1 U847 ( .A1(KEYINPUT57), .A2(n1161), .ZN(n1160) );
NOR2_X1 U848 ( .A1(n1120), .A2(n1162), .ZN(G51) );
NOR2_X1 U849 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U850 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U851 ( .A1(n1068), .A2(n1167), .ZN(n1166) );
INV_X1 U852 ( .A(n1125), .ZN(n1167) );
NOR2_X1 U853 ( .A1(n1168), .A2(n1010), .ZN(n1125) );
NOR3_X1 U854 ( .A1(n1112), .A2(n1113), .A3(n1075), .ZN(n1010) );
NAND4_X1 U855 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1075) );
NOR4_X1 U856 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1172) );
INV_X1 U857 ( .A(n1177), .ZN(n1176) );
INV_X1 U858 ( .A(n1178), .ZN(n1175) );
NAND2_X1 U859 ( .A1(n1179), .A2(n1180), .ZN(n1171) );
XNOR2_X1 U860 ( .A(KEYINPUT37), .B(n1181), .ZN(n1179) );
NAND3_X1 U861 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1169) );
NAND2_X1 U862 ( .A1(n1185), .A2(n1186), .ZN(n1183) );
OR2_X1 U863 ( .A1(n1187), .A2(KEYINPUT48), .ZN(n1185) );
NAND3_X1 U864 ( .A1(n1188), .A2(n1189), .A3(n1023), .ZN(n1182) );
NAND2_X1 U865 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
XNOR2_X1 U866 ( .A(KEYINPUT35), .B(n1022), .ZN(n1190) );
NAND2_X1 U867 ( .A1(KEYINPUT48), .A2(n1192), .ZN(n1188) );
AND3_X1 U868 ( .A1(n1193), .A2(n1025), .A3(n1191), .ZN(n1113) );
NAND4_X1 U869 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1112) );
NOR4_X1 U870 ( .A1(n1198), .A2(n1199), .A3(n1000), .A4(n1200), .ZN(n1197) );
AND3_X1 U871 ( .A1(n1039), .A2(n1025), .A3(n1193), .ZN(n1000) );
NAND2_X1 U872 ( .A1(n1201), .A2(n1202), .ZN(n1196) );
XNOR2_X1 U873 ( .A(n1015), .B(KEYINPUT1), .ZN(n1201) );
NOR2_X1 U874 ( .A1(n1203), .A2(n1204), .ZN(n1165) );
AND2_X1 U875 ( .A1(n1204), .A2(n1203), .ZN(n1163) );
XNOR2_X1 U876 ( .A(n1205), .B(n1206), .ZN(n1203) );
XOR2_X1 U877 ( .A(KEYINPUT29), .B(n1207), .Z(n1206) );
NOR2_X1 U878 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XOR2_X1 U879 ( .A(n1210), .B(KEYINPUT27), .Z(n1209) );
NAND2_X1 U880 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NOR2_X1 U881 ( .A1(n1212), .A2(n1211), .ZN(n1208) );
NAND3_X1 U882 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1211) );
OR2_X1 U883 ( .A1(n1216), .A2(KEYINPUT43), .ZN(n1215) );
NAND3_X1 U884 ( .A1(KEYINPUT43), .A2(n1216), .A3(n1217), .ZN(n1214) );
NAND2_X1 U885 ( .A1(G125), .A2(n1218), .ZN(n1213) );
NAND2_X1 U886 ( .A1(KEYINPUT43), .A2(n1219), .ZN(n1218) );
XNOR2_X1 U887 ( .A(KEYINPUT39), .B(n1220), .ZN(n1219) );
INV_X1 U888 ( .A(KEYINPUT25), .ZN(n1204) );
NOR2_X1 U889 ( .A1(n1002), .A2(G952), .ZN(n1120) );
XNOR2_X1 U890 ( .A(G146), .B(n1170), .ZN(G48) );
NAND4_X1 U891 ( .A1(n1184), .A2(n1221), .A3(n1191), .A4(n1180), .ZN(n1170) );
XNOR2_X1 U892 ( .A(n1083), .B(n1174), .ZN(G45) );
AND4_X1 U893 ( .A1(n1054), .A2(n1222), .A3(n1022), .A4(n1223), .ZN(n1174) );
NOR2_X1 U894 ( .A1(n1027), .A2(n1224), .ZN(n1223) );
NAND2_X1 U895 ( .A1(n1225), .A2(n1226), .ZN(G42) );
OR2_X1 U896 ( .A1(n1177), .A2(G140), .ZN(n1226) );
XOR2_X1 U897 ( .A(n1227), .B(KEYINPUT47), .Z(n1225) );
NAND2_X1 U898 ( .A1(G140), .A2(n1177), .ZN(n1227) );
NAND4_X1 U899 ( .A1(n1023), .A2(n1184), .A3(n1024), .A4(n1191), .ZN(n1177) );
XOR2_X1 U900 ( .A(G137), .B(n1228), .Z(G39) );
NOR3_X1 U901 ( .A1(n1229), .A2(n1224), .A3(n1187), .ZN(n1228) );
XNOR2_X1 U902 ( .A(KEYINPUT4), .B(n1186), .ZN(n1229) );
XNOR2_X1 U903 ( .A(G134), .B(n1178), .ZN(G36) );
NAND2_X1 U904 ( .A1(n1230), .A2(n1039), .ZN(n1178) );
NAND2_X1 U905 ( .A1(n1231), .A2(n1232), .ZN(G33) );
NAND2_X1 U906 ( .A1(G131), .A2(n1233), .ZN(n1232) );
NAND2_X1 U907 ( .A1(n1230), .A2(n1191), .ZN(n1233) );
INV_X1 U908 ( .A(n1234), .ZN(n1230) );
XOR2_X1 U909 ( .A(KEYINPUT18), .B(n1235), .Z(n1231) );
NOR3_X1 U910 ( .A1(n1234), .A2(G131), .A3(n1236), .ZN(n1235) );
NAND3_X1 U911 ( .A1(n1184), .A2(n1022), .A3(n1023), .ZN(n1234) );
INV_X1 U912 ( .A(n1186), .ZN(n1023) );
NAND2_X1 U913 ( .A1(n1030), .A2(n1065), .ZN(n1186) );
INV_X1 U914 ( .A(n1224), .ZN(n1184) );
NAND2_X1 U915 ( .A1(n1237), .A2(n1238), .ZN(n1224) );
INV_X1 U916 ( .A(n1041), .ZN(n1237) );
XOR2_X1 U917 ( .A(n1239), .B(KEYINPUT14), .Z(n1041) );
XNOR2_X1 U918 ( .A(n1240), .B(n1241), .ZN(G30) );
NOR2_X1 U919 ( .A1(n1027), .A2(n1181), .ZN(n1241) );
NAND4_X1 U920 ( .A1(n1221), .A2(n1039), .A3(n1239), .A4(n1238), .ZN(n1181) );
INV_X1 U921 ( .A(n1180), .ZN(n1027) );
XNOR2_X1 U922 ( .A(n1242), .B(n1199), .ZN(G3) );
AND3_X1 U923 ( .A1(n1193), .A2(n1022), .A3(n1017), .ZN(n1199) );
XOR2_X1 U924 ( .A(n1173), .B(n1243), .Z(G27) );
NOR2_X1 U925 ( .A1(KEYINPUT60), .A2(n1217), .ZN(n1243) );
INV_X1 U926 ( .A(G125), .ZN(n1217) );
AND4_X1 U927 ( .A1(n1035), .A2(n1024), .A3(n1180), .A4(n1238), .ZN(n1173) );
NAND2_X1 U928 ( .A1(n1244), .A2(n1245), .ZN(n1238) );
NAND4_X1 U929 ( .A1(G902), .A2(G953), .A3(n1046), .A4(n1098), .ZN(n1245) );
INV_X1 U930 ( .A(G900), .ZN(n1098) );
NOR2_X1 U931 ( .A1(n1246), .A2(n1236), .ZN(n1035) );
XNOR2_X1 U932 ( .A(G122), .B(n1194), .ZN(G24) );
NAND4_X1 U933 ( .A1(n1247), .A2(n1025), .A3(n1054), .A4(n1222), .ZN(n1194) );
INV_X1 U934 ( .A(n1034), .ZN(n1025) );
NAND2_X1 U935 ( .A1(n1248), .A2(n1249), .ZN(n1034) );
XNOR2_X1 U936 ( .A(n1250), .B(n1049), .ZN(n1248) );
XOR2_X1 U937 ( .A(n1195), .B(n1251), .Z(G21) );
NAND2_X1 U938 ( .A1(KEYINPUT5), .A2(G119), .ZN(n1251) );
NAND2_X1 U939 ( .A1(n1247), .A2(n1192), .ZN(n1195) );
INV_X1 U940 ( .A(n1187), .ZN(n1192) );
NAND2_X1 U941 ( .A1(n1017), .A2(n1221), .ZN(n1187) );
XOR2_X1 U942 ( .A(G116), .B(n1198), .Z(G18) );
AND3_X1 U943 ( .A1(n1039), .A2(n1022), .A3(n1247), .ZN(n1198) );
AND3_X1 U944 ( .A1(n1180), .A2(n1252), .A3(n1015), .ZN(n1247) );
XOR2_X1 U945 ( .A(n1253), .B(KEYINPUT41), .Z(n1180) );
NOR2_X1 U946 ( .A1(n1222), .A2(n1254), .ZN(n1039) );
XNOR2_X1 U947 ( .A(G113), .B(n1255), .ZN(G15) );
NAND3_X1 U948 ( .A1(n1202), .A2(n1015), .A3(KEYINPUT0), .ZN(n1255) );
INV_X1 U949 ( .A(n1246), .ZN(n1015) );
NAND2_X1 U950 ( .A1(n1044), .A2(n1066), .ZN(n1246) );
AND4_X1 U951 ( .A1(n1191), .A2(n1253), .A3(n1022), .A4(n1252), .ZN(n1202) );
NAND2_X1 U952 ( .A1(n1256), .A2(n1257), .ZN(n1022) );
NAND3_X1 U953 ( .A1(n1053), .A2(n1049), .A3(n1250), .ZN(n1257) );
INV_X1 U954 ( .A(KEYINPUT7), .ZN(n1250) );
NAND2_X1 U955 ( .A1(KEYINPUT7), .A2(n1221), .ZN(n1256) );
NOR2_X1 U956 ( .A1(n1049), .A2(n1249), .ZN(n1221) );
INV_X1 U957 ( .A(n1053), .ZN(n1249) );
INV_X1 U958 ( .A(n1236), .ZN(n1191) );
NAND2_X1 U959 ( .A1(n1254), .A2(n1222), .ZN(n1236) );
INV_X1 U960 ( .A(n1054), .ZN(n1254) );
XNOR2_X1 U961 ( .A(n1161), .B(n1200), .ZN(G12) );
AND3_X1 U962 ( .A1(n1024), .A2(n1193), .A3(n1017), .ZN(n1200) );
NOR2_X1 U963 ( .A1(n1054), .A2(n1222), .ZN(n1017) );
NAND2_X1 U964 ( .A1(n1048), .A2(n1258), .ZN(n1222) );
OR2_X1 U965 ( .A1(n1055), .A2(n1056), .ZN(n1258) );
NAND2_X1 U966 ( .A1(n1056), .A2(n1055), .ZN(n1048) );
XNOR2_X1 U967 ( .A(G475), .B(KEYINPUT22), .ZN(n1055) );
AND2_X1 U968 ( .A1(n1136), .A2(n1168), .ZN(n1056) );
XOR2_X1 U969 ( .A(n1259), .B(n1260), .Z(n1136) );
XOR2_X1 U970 ( .A(n1261), .B(n1262), .Z(n1260) );
XNOR2_X1 U971 ( .A(G113), .B(G122), .ZN(n1262) );
NAND2_X1 U972 ( .A1(KEYINPUT44), .A2(n1263), .ZN(n1261) );
XNOR2_X1 U973 ( .A(KEYINPUT61), .B(n1080), .ZN(n1263) );
INV_X1 U974 ( .A(n1264), .ZN(n1080) );
XOR2_X1 U975 ( .A(n1265), .B(n1266), .Z(n1259) );
XOR2_X1 U976 ( .A(n1267), .B(n1268), .Z(n1265) );
NOR2_X1 U977 ( .A1(G131), .A2(KEYINPUT54), .ZN(n1268) );
NAND2_X1 U978 ( .A1(n1269), .A2(G214), .ZN(n1267) );
XNOR2_X1 U979 ( .A(n1270), .B(G478), .ZN(n1054) );
NAND2_X1 U980 ( .A1(n1133), .A2(n1168), .ZN(n1270) );
XNOR2_X1 U981 ( .A(n1271), .B(n1272), .ZN(n1133) );
XOR2_X1 U982 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U983 ( .A(n1240), .B(G122), .ZN(n1274) );
XNOR2_X1 U984 ( .A(n1083), .B(G134), .ZN(n1273) );
INV_X1 U985 ( .A(G143), .ZN(n1083) );
XOR2_X1 U986 ( .A(n1275), .B(n1276), .Z(n1271) );
XOR2_X1 U987 ( .A(n1277), .B(G116), .Z(n1275) );
NAND2_X1 U988 ( .A1(G217), .A2(n1278), .ZN(n1277) );
AND3_X1 U989 ( .A1(n1253), .A2(n1252), .A3(n1239), .ZN(n1193) );
NOR2_X1 U990 ( .A1(n1044), .A2(n1043), .ZN(n1239) );
INV_X1 U991 ( .A(n1066), .ZN(n1043) );
NAND2_X1 U992 ( .A1(G221), .A2(n1279), .ZN(n1066) );
XNOR2_X1 U993 ( .A(n1064), .B(KEYINPUT26), .ZN(n1044) );
XOR2_X1 U994 ( .A(n1280), .B(n1281), .Z(n1064) );
XOR2_X1 U995 ( .A(KEYINPUT23), .B(G469), .Z(n1281) );
NAND2_X1 U996 ( .A1(n1282), .A2(n1168), .ZN(n1280) );
XOR2_X1 U997 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U998 ( .A(n1155), .B(n1285), .Z(n1284) );
XNOR2_X1 U999 ( .A(KEYINPUT32), .B(n1161), .ZN(n1285) );
NOR2_X1 U1000 ( .A1(n1097), .A2(G953), .ZN(n1155) );
INV_X1 U1001 ( .A(G227), .ZN(n1097) );
XNOR2_X1 U1002 ( .A(n1150), .B(n1286), .ZN(n1283) );
XNOR2_X1 U1003 ( .A(n1287), .B(n1288), .ZN(n1150) );
XOR2_X1 U1004 ( .A(n1266), .B(n1289), .Z(n1288) );
XNOR2_X1 U1005 ( .A(n1137), .B(G143), .ZN(n1266) );
XOR2_X1 U1006 ( .A(n1290), .B(KEYINPUT6), .Z(n1287) );
NAND2_X1 U1007 ( .A1(n1244), .A2(n1291), .ZN(n1252) );
NAND3_X1 U1008 ( .A1(n1115), .A2(n1046), .A3(G902), .ZN(n1291) );
NOR2_X1 U1009 ( .A1(G898), .A2(n1002), .ZN(n1115) );
NAND3_X1 U1010 ( .A1(n1046), .A2(n1002), .A3(G952), .ZN(n1244) );
NAND2_X1 U1011 ( .A1(G237), .A2(G234), .ZN(n1046) );
NOR2_X1 U1012 ( .A1(n1030), .A2(n1029), .ZN(n1253) );
INV_X1 U1013 ( .A(n1065), .ZN(n1029) );
NAND2_X1 U1014 ( .A1(G214), .A2(n1292), .ZN(n1065) );
XNOR2_X1 U1015 ( .A(n1062), .B(n1068), .ZN(n1030) );
NAND2_X1 U1016 ( .A1(G210), .A2(n1292), .ZN(n1068) );
NAND2_X1 U1017 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U1018 ( .A(KEYINPUT63), .B(G237), .Z(n1293) );
NAND2_X1 U1019 ( .A1(n1295), .A2(n1296), .ZN(n1062) );
XOR2_X1 U1020 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U1021 ( .A(n1299), .B(n1205), .Z(n1298) );
XNOR2_X1 U1022 ( .A(n1116), .B(n1119), .ZN(n1205) );
XOR2_X1 U1023 ( .A(n1161), .B(n1300), .Z(n1119) );
NOR2_X1 U1024 ( .A1(KEYINPUT2), .A2(n1301), .ZN(n1300) );
INV_X1 U1025 ( .A(G122), .ZN(n1301) );
XOR2_X1 U1026 ( .A(n1302), .B(n1303), .Z(n1116) );
XNOR2_X1 U1027 ( .A(G113), .B(n1304), .ZN(n1303) );
NAND2_X1 U1028 ( .A1(KEYINPUT13), .A2(n1137), .ZN(n1304) );
INV_X1 U1029 ( .A(G104), .ZN(n1137) );
XNOR2_X1 U1030 ( .A(n1289), .B(n1305), .ZN(n1302) );
NOR2_X1 U1031 ( .A1(KEYINPUT42), .A2(n1306), .ZN(n1305) );
XOR2_X1 U1032 ( .A(G101), .B(n1276), .Z(n1289) );
XOR2_X1 U1033 ( .A(G107), .B(KEYINPUT51), .Z(n1276) );
NAND2_X1 U1034 ( .A1(KEYINPUT33), .A2(n1220), .ZN(n1299) );
INV_X1 U1035 ( .A(n1216), .ZN(n1220) );
XOR2_X1 U1036 ( .A(G128), .B(n1307), .Z(n1216) );
XNOR2_X1 U1037 ( .A(G125), .B(n1212), .ZN(n1297) );
NAND2_X1 U1038 ( .A1(G224), .A2(n1002), .ZN(n1212) );
XNOR2_X1 U1039 ( .A(KEYINPUT58), .B(n1168), .ZN(n1295) );
NOR2_X1 U1040 ( .A1(n1053), .A2(n1049), .ZN(n1024) );
XOR2_X1 U1041 ( .A(n1308), .B(n1126), .Z(n1049) );
AND2_X1 U1042 ( .A1(G217), .A2(n1279), .ZN(n1126) );
NAND2_X1 U1043 ( .A1(G234), .A2(n1294), .ZN(n1279) );
XNOR2_X1 U1044 ( .A(n1168), .B(KEYINPUT56), .ZN(n1294) );
OR2_X1 U1045 ( .A1(n1124), .A2(G902), .ZN(n1308) );
XNOR2_X1 U1046 ( .A(n1309), .B(n1310), .ZN(n1124) );
XNOR2_X1 U1047 ( .A(n1161), .B(n1311), .ZN(n1310) );
XNOR2_X1 U1048 ( .A(n1240), .B(G119), .ZN(n1311) );
XNOR2_X1 U1049 ( .A(n1312), .B(n1313), .ZN(n1309) );
INV_X1 U1050 ( .A(n1090), .ZN(n1313) );
XNOR2_X1 U1051 ( .A(n1264), .B(n1314), .ZN(n1312) );
AND2_X1 U1052 ( .A1(G221), .A2(n1278), .ZN(n1314) );
AND2_X1 U1053 ( .A1(G234), .A2(n1002), .ZN(n1278) );
INV_X1 U1054 ( .A(G953), .ZN(n1002) );
XOR2_X1 U1055 ( .A(G125), .B(n1286), .Z(n1264) );
XOR2_X1 U1056 ( .A(G140), .B(G146), .Z(n1286) );
XNOR2_X1 U1057 ( .A(n1315), .B(G472), .ZN(n1053) );
NAND2_X1 U1058 ( .A1(n1316), .A2(n1168), .ZN(n1315) );
INV_X1 U1059 ( .A(G902), .ZN(n1168) );
XNOR2_X1 U1060 ( .A(n1139), .B(n1317), .ZN(n1316) );
XOR2_X1 U1061 ( .A(KEYINPUT16), .B(n1318), .Z(n1317) );
NOR2_X1 U1062 ( .A1(n1143), .A2(n1145), .ZN(n1318) );
NOR2_X1 U1063 ( .A1(n1319), .A2(n1242), .ZN(n1145) );
AND2_X1 U1064 ( .A1(n1242), .A2(n1319), .ZN(n1143) );
NAND2_X1 U1065 ( .A1(n1269), .A2(G210), .ZN(n1319) );
NOR2_X1 U1066 ( .A1(G953), .A2(G237), .ZN(n1269) );
INV_X1 U1067 ( .A(G101), .ZN(n1242) );
XNOR2_X1 U1068 ( .A(n1320), .B(n1321), .ZN(n1139) );
XNOR2_X1 U1069 ( .A(n1322), .B(n1307), .ZN(n1321) );
NOR2_X1 U1070 ( .A1(KEYINPUT8), .A2(n1323), .ZN(n1307) );
XNOR2_X1 U1071 ( .A(G143), .B(G146), .ZN(n1323) );
INV_X1 U1072 ( .A(G113), .ZN(n1322) );
XNOR2_X1 U1073 ( .A(n1290), .B(n1306), .ZN(n1320) );
XNOR2_X1 U1074 ( .A(G116), .B(G119), .ZN(n1306) );
XOR2_X1 U1075 ( .A(n1324), .B(n1081), .Z(n1290) );
XNOR2_X1 U1076 ( .A(n1240), .B(G131), .ZN(n1081) );
INV_X1 U1077 ( .A(G128), .ZN(n1240) );
XNOR2_X1 U1078 ( .A(n1325), .B(n1089), .ZN(n1324) );
INV_X1 U1079 ( .A(G134), .ZN(n1089) );
NAND2_X1 U1080 ( .A1(KEYINPUT17), .A2(n1090), .ZN(n1325) );
XOR2_X1 U1081 ( .A(G137), .B(KEYINPUT52), .Z(n1090) );
INV_X1 U1082 ( .A(G110), .ZN(n1161) );
endmodule


