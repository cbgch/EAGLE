//Key = 0010011010001010000111001110111101111111101101110111101111101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320;

XNOR2_X1 U719 ( .A(n1009), .B(n1010), .ZN(G9) );
NOR2_X1 U720 ( .A1(KEYINPUT10), .A2(n1011), .ZN(n1010) );
NOR2_X1 U721 ( .A1(n1012), .A2(n1013), .ZN(G75) );
NOR3_X1 U722 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NOR2_X1 U723 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NOR2_X1 U724 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
XOR2_X1 U725 ( .A(n1021), .B(KEYINPUT36), .Z(n1020) );
NAND2_X1 U726 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NOR2_X1 U727 ( .A1(n1024), .A2(n1025), .ZN(n1019) );
NOR2_X1 U728 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR3_X1 U729 ( .A1(n1028), .A2(n1029), .A3(n1023), .ZN(n1027) );
NOR2_X1 U730 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR2_X1 U731 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U732 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U733 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U734 ( .A1(n1038), .A2(n1039), .ZN(n1030) );
NOR2_X1 U735 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR3_X1 U736 ( .A1(n1042), .A2(n1043), .A3(n1033), .ZN(n1026) );
XOR2_X1 U737 ( .A(KEYINPUT25), .B(n1044), .Z(n1042) );
NAND3_X1 U738 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1014) );
NAND3_X1 U739 ( .A1(n1048), .A2(n1049), .A3(n1022), .ZN(n1047) );
NOR4_X1 U740 ( .A1(n1033), .A2(n1039), .A3(n1028), .A4(n1024), .ZN(n1022) );
INV_X1 U741 ( .A(n1050), .ZN(n1024) );
INV_X1 U742 ( .A(n1044), .ZN(n1039) );
NAND2_X1 U743 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NAND2_X1 U744 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR3_X1 U745 ( .A1(n1055), .A2(G953), .A3(G952), .ZN(n1012) );
INV_X1 U746 ( .A(n1045), .ZN(n1055) );
NAND4_X1 U747 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1045) );
NOR4_X1 U748 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1059) );
XOR2_X1 U749 ( .A(KEYINPUT63), .B(n1064), .Z(n1063) );
XOR2_X1 U750 ( .A(n1065), .B(n1066), .Z(n1062) );
XOR2_X1 U751 ( .A(n1067), .B(n1068), .Z(n1061) );
XNOR2_X1 U752 ( .A(n1069), .B(n1070), .ZN(n1060) );
NOR2_X1 U753 ( .A1(KEYINPUT59), .A2(n1071), .ZN(n1070) );
NOR3_X1 U754 ( .A1(n1072), .A2(n1073), .A3(n1053), .ZN(n1058) );
NAND2_X1 U755 ( .A1(G478), .A2(n1074), .ZN(n1057) );
XNOR2_X1 U756 ( .A(n1075), .B(n1076), .ZN(n1056) );
NAND2_X1 U757 ( .A1(KEYINPUT61), .A2(n1077), .ZN(n1075) );
XOR2_X1 U758 ( .A(n1078), .B(n1079), .Z(G72) );
NAND2_X1 U759 ( .A1(G953), .A2(n1080), .ZN(n1079) );
NAND2_X1 U760 ( .A1(G900), .A2(G227), .ZN(n1080) );
NAND2_X1 U761 ( .A1(n1081), .A2(n1082), .ZN(n1078) );
NAND4_X1 U762 ( .A1(KEYINPUT20), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1082) );
NAND2_X1 U763 ( .A1(n1086), .A2(n1087), .ZN(n1081) );
NAND2_X1 U764 ( .A1(n1083), .A2(n1088), .ZN(n1087) );
OR2_X1 U765 ( .A1(KEYINPUT20), .A2(n1084), .ZN(n1088) );
AND2_X1 U766 ( .A1(n1089), .A2(n1046), .ZN(n1083) );
NAND2_X1 U767 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U768 ( .A1(n1084), .A2(n1085), .ZN(n1086) );
INV_X1 U769 ( .A(KEYINPUT3), .ZN(n1085) );
AND2_X1 U770 ( .A1(n1092), .A2(n1093), .ZN(n1084) );
NAND2_X1 U771 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
XOR2_X1 U772 ( .A(n1096), .B(n1097), .Z(n1092) );
XNOR2_X1 U773 ( .A(n1098), .B(n1099), .ZN(n1096) );
NAND2_X1 U774 ( .A1(KEYINPUT37), .A2(n1100), .ZN(n1099) );
XOR2_X1 U775 ( .A(n1101), .B(n1102), .Z(n1100) );
NAND2_X1 U776 ( .A1(n1103), .A2(KEYINPUT54), .ZN(n1102) );
XNOR2_X1 U777 ( .A(n1104), .B(KEYINPUT47), .ZN(n1103) );
NAND2_X1 U778 ( .A1(n1105), .A2(KEYINPUT29), .ZN(n1098) );
XNOR2_X1 U779 ( .A(G125), .B(n1106), .ZN(n1105) );
NOR2_X1 U780 ( .A1(G140), .A2(KEYINPUT17), .ZN(n1106) );
XOR2_X1 U781 ( .A(n1107), .B(n1108), .Z(G69) );
NOR2_X1 U782 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR3_X1 U783 ( .A1(n1046), .A2(n1111), .A3(n1112), .ZN(n1110) );
INV_X1 U784 ( .A(G224), .ZN(n1112) );
XOR2_X1 U785 ( .A(KEYINPUT26), .B(G898), .Z(n1111) );
AND3_X1 U786 ( .A1(n1046), .A2(n1113), .A3(n1114), .ZN(n1109) );
NOR3_X1 U787 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1107) );
NOR2_X1 U788 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
XOR2_X1 U789 ( .A(KEYINPUT32), .B(n1120), .Z(n1115) );
AND2_X1 U790 ( .A1(n1119), .A2(n1118), .ZN(n1120) );
NOR2_X1 U791 ( .A1(n1121), .A2(n1122), .ZN(G66) );
NOR3_X1 U792 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1122) );
NOR3_X1 U793 ( .A1(n1126), .A2(n1068), .A3(n1127), .ZN(n1125) );
NOR2_X1 U794 ( .A1(n1128), .A2(n1129), .ZN(n1124) );
NOR2_X1 U795 ( .A1(n1130), .A2(n1068), .ZN(n1129) );
INV_X1 U796 ( .A(n1016), .ZN(n1130) );
INV_X1 U797 ( .A(n1126), .ZN(n1128) );
NOR2_X1 U798 ( .A1(n1121), .A2(n1131), .ZN(G63) );
XNOR2_X1 U799 ( .A(n1132), .B(n1133), .ZN(n1131) );
NOR2_X1 U800 ( .A1(n1134), .A2(n1127), .ZN(n1133) );
NOR2_X1 U801 ( .A1(n1121), .A2(n1135), .ZN(G60) );
XNOR2_X1 U802 ( .A(n1136), .B(n1137), .ZN(n1135) );
NOR2_X1 U803 ( .A1(n1138), .A2(n1127), .ZN(n1136) );
INV_X1 U804 ( .A(G475), .ZN(n1138) );
XOR2_X1 U805 ( .A(n1113), .B(n1139), .Z(G6) );
XNOR2_X1 U806 ( .A(G104), .B(KEYINPUT18), .ZN(n1139) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1140), .ZN(G57) );
XOR2_X1 U808 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U809 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U810 ( .A1(n1065), .A2(n1127), .ZN(n1143) );
INV_X1 U811 ( .A(G472), .ZN(n1065) );
XOR2_X1 U812 ( .A(n1145), .B(G101), .Z(n1141) );
NOR2_X1 U813 ( .A1(n1121), .A2(n1146), .ZN(G54) );
XOR2_X1 U814 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U815 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR2_X1 U816 ( .A1(KEYINPUT1), .A2(n1151), .ZN(n1149) );
XNOR2_X1 U817 ( .A(n1152), .B(n1153), .ZN(n1151) );
NAND2_X1 U818 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NAND2_X1 U819 ( .A1(G140), .A2(n1156), .ZN(n1155) );
XOR2_X1 U820 ( .A(KEYINPUT5), .B(n1157), .Z(n1154) );
NOR2_X1 U821 ( .A1(G140), .A2(n1156), .ZN(n1157) );
XOR2_X1 U822 ( .A(n1158), .B(n1159), .Z(n1147) );
NOR2_X1 U823 ( .A1(n1071), .A2(n1127), .ZN(n1159) );
INV_X1 U824 ( .A(G469), .ZN(n1071) );
NAND3_X1 U825 ( .A1(n1160), .A2(n1161), .A3(KEYINPUT51), .ZN(n1158) );
NAND3_X1 U826 ( .A1(n1097), .A2(n1162), .A3(n1163), .ZN(n1161) );
INV_X1 U827 ( .A(KEYINPUT12), .ZN(n1163) );
NAND2_X1 U828 ( .A1(n1164), .A2(KEYINPUT12), .ZN(n1160) );
NOR2_X1 U829 ( .A1(n1121), .A2(n1165), .ZN(G51) );
XOR2_X1 U830 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U831 ( .A1(n1168), .A2(n1127), .ZN(n1167) );
NAND2_X1 U832 ( .A1(G902), .A2(n1016), .ZN(n1127) );
NAND4_X1 U833 ( .A1(n1169), .A2(n1114), .A3(n1090), .A4(n1170), .ZN(n1016) );
XNOR2_X1 U834 ( .A(KEYINPUT21), .B(n1113), .ZN(n1170) );
NAND2_X1 U835 ( .A1(n1041), .A2(n1171), .ZN(n1113) );
AND3_X1 U836 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1090) );
NAND2_X1 U837 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND2_X1 U838 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NAND2_X1 U839 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XOR2_X1 U840 ( .A(n1018), .B(KEYINPUT42), .Z(n1179) );
NAND2_X1 U841 ( .A1(n1041), .A2(n1181), .ZN(n1177) );
AND4_X1 U842 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1114) );
AND4_X1 U843 ( .A1(n1009), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1185) );
NAND2_X1 U844 ( .A1(n1040), .A2(n1171), .ZN(n1009) );
AND3_X1 U845 ( .A1(n1035), .A2(n1181), .A3(n1189), .ZN(n1171) );
AND3_X1 U846 ( .A1(n1190), .A2(n1191), .A3(n1048), .ZN(n1189) );
NAND2_X1 U847 ( .A1(n1192), .A2(n1181), .ZN(n1184) );
XNOR2_X1 U848 ( .A(n1193), .B(KEYINPUT49), .ZN(n1192) );
XNOR2_X1 U849 ( .A(n1091), .B(KEYINPUT34), .ZN(n1169) );
AND4_X1 U850 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1091) );
NAND2_X1 U851 ( .A1(n1198), .A2(n1181), .ZN(n1194) );
XOR2_X1 U852 ( .A(n1199), .B(KEYINPUT33), .Z(n1198) );
NAND4_X1 U853 ( .A1(n1200), .A2(n1040), .A3(n1035), .A4(n1201), .ZN(n1199) );
XNOR2_X1 U854 ( .A(KEYINPUT35), .B(n1202), .ZN(n1201) );
NOR2_X1 U855 ( .A1(KEYINPUT15), .A2(n1203), .ZN(n1166) );
NOR2_X1 U856 ( .A1(n1046), .A2(G952), .ZN(n1121) );
XNOR2_X1 U857 ( .A(G146), .B(n1204), .ZN(G48) );
NAND3_X1 U858 ( .A1(n1175), .A2(n1041), .A3(n1205), .ZN(n1204) );
XOR2_X1 U859 ( .A(n1051), .B(KEYINPUT39), .Z(n1205) );
INV_X1 U860 ( .A(n1181), .ZN(n1051) );
XOR2_X1 U861 ( .A(n1206), .B(G143), .Z(G45) );
NAND2_X1 U862 ( .A1(KEYINPUT31), .A2(n1172), .ZN(n1206) );
NAND3_X1 U863 ( .A1(n1207), .A2(n1202), .A3(n1208), .ZN(n1172) );
XNOR2_X1 U864 ( .A(G140), .B(n1173), .ZN(G42) );
NAND2_X1 U865 ( .A1(n1209), .A2(n1210), .ZN(n1173) );
XOR2_X1 U866 ( .A(G137), .B(n1211), .Z(G39) );
NOR3_X1 U867 ( .A1(n1212), .A2(n1033), .A3(n1018), .ZN(n1211) );
NAND2_X1 U868 ( .A1(n1213), .A2(n1214), .ZN(G36) );
NAND2_X1 U869 ( .A1(G134), .A2(n1195), .ZN(n1214) );
XOR2_X1 U870 ( .A(n1215), .B(KEYINPUT27), .Z(n1213) );
OR2_X1 U871 ( .A1(n1195), .A2(G134), .ZN(n1215) );
NAND3_X1 U872 ( .A1(n1216), .A2(n1040), .A3(n1210), .ZN(n1195) );
XNOR2_X1 U873 ( .A(n1196), .B(n1217), .ZN(G33) );
NOR2_X1 U874 ( .A1(KEYINPUT41), .A2(n1101), .ZN(n1217) );
NAND3_X1 U875 ( .A1(n1041), .A2(n1216), .A3(n1210), .ZN(n1196) );
AND3_X1 U876 ( .A1(n1035), .A2(n1202), .A3(n1218), .ZN(n1210) );
INV_X1 U877 ( .A(n1018), .ZN(n1218) );
NAND2_X1 U878 ( .A1(n1054), .A2(n1219), .ZN(n1018) );
XOR2_X1 U879 ( .A(G128), .B(n1220), .Z(G30) );
AND3_X1 U880 ( .A1(n1175), .A2(n1181), .A3(n1040), .ZN(n1220) );
INV_X1 U881 ( .A(n1212), .ZN(n1175) );
NAND3_X1 U882 ( .A1(n1035), .A2(n1202), .A3(n1200), .ZN(n1212) );
XOR2_X1 U883 ( .A(n1221), .B(n1182), .Z(G3) );
NAND3_X1 U884 ( .A1(n1180), .A2(n1191), .A3(n1208), .ZN(n1182) );
AND3_X1 U885 ( .A1(n1035), .A2(n1181), .A3(n1216), .ZN(n1208) );
XNOR2_X1 U886 ( .A(G125), .B(n1197), .ZN(G27) );
NAND4_X1 U887 ( .A1(n1209), .A2(n1044), .A3(n1181), .A4(n1202), .ZN(n1197) );
NAND2_X1 U888 ( .A1(n1222), .A2(n1223), .ZN(n1202) );
NAND4_X1 U889 ( .A1(n1094), .A2(G902), .A3(n1050), .A4(n1095), .ZN(n1223) );
INV_X1 U890 ( .A(G900), .ZN(n1095) );
XNOR2_X1 U891 ( .A(KEYINPUT43), .B(n1224), .ZN(n1222) );
AND3_X1 U892 ( .A1(n1041), .A2(n1190), .A3(n1023), .ZN(n1209) );
XNOR2_X1 U893 ( .A(G122), .B(n1183), .ZN(G24) );
NAND4_X1 U894 ( .A1(n1207), .A2(n1225), .A3(n1190), .A4(n1048), .ZN(n1183) );
AND2_X1 U895 ( .A1(n1226), .A2(n1227), .ZN(n1207) );
XOR2_X1 U896 ( .A(KEYINPUT9), .B(n1064), .Z(n1226) );
XOR2_X1 U897 ( .A(G119), .B(n1228), .Z(G21) );
NOR2_X1 U898 ( .A1(KEYINPUT11), .A2(n1188), .ZN(n1228) );
NAND3_X1 U899 ( .A1(n1200), .A2(n1225), .A3(n1180), .ZN(n1188) );
NOR2_X1 U900 ( .A1(n1048), .A2(n1190), .ZN(n1200) );
XNOR2_X1 U901 ( .A(G116), .B(n1187), .ZN(G18) );
NAND3_X1 U902 ( .A1(n1216), .A2(n1040), .A3(n1225), .ZN(n1187) );
AND2_X1 U903 ( .A1(n1229), .A2(n1227), .ZN(n1040) );
XNOR2_X1 U904 ( .A(G113), .B(n1186), .ZN(G15) );
NAND3_X1 U905 ( .A1(n1225), .A2(n1216), .A3(n1041), .ZN(n1186) );
NOR2_X1 U906 ( .A1(n1227), .A2(n1229), .ZN(n1041) );
INV_X1 U907 ( .A(n1043), .ZN(n1216) );
NAND2_X1 U908 ( .A1(n1028), .A2(n1048), .ZN(n1043) );
AND3_X1 U909 ( .A1(n1181), .A2(n1191), .A3(n1044), .ZN(n1225) );
NOR2_X1 U910 ( .A1(n1036), .A2(n1072), .ZN(n1044) );
INV_X1 U911 ( .A(n1037), .ZN(n1072) );
NAND3_X1 U912 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(G12) );
NAND3_X1 U913 ( .A1(n1181), .A2(n1233), .A3(n1193), .ZN(n1232) );
NAND2_X1 U914 ( .A1(KEYINPUT24), .A2(n1234), .ZN(n1233) );
NAND2_X1 U915 ( .A1(KEYINPUT57), .A2(n1156), .ZN(n1234) );
OR2_X1 U916 ( .A1(G110), .A2(KEYINPUT24), .ZN(n1231) );
NAND3_X1 U917 ( .A1(G110), .A2(n1235), .A3(KEYINPUT24), .ZN(n1230) );
NAND3_X1 U918 ( .A1(n1193), .A2(n1181), .A3(KEYINPUT57), .ZN(n1235) );
NOR2_X1 U919 ( .A1(n1054), .A2(n1053), .ZN(n1181) );
INV_X1 U920 ( .A(n1219), .ZN(n1053) );
NAND2_X1 U921 ( .A1(G214), .A2(n1236), .ZN(n1219) );
XOR2_X1 U922 ( .A(n1076), .B(n1077), .Z(n1054) );
INV_X1 U923 ( .A(n1168), .ZN(n1077) );
NAND2_X1 U924 ( .A1(G210), .A2(n1236), .ZN(n1168) );
NAND2_X1 U925 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NAND2_X1 U926 ( .A1(n1239), .A2(n1240), .ZN(n1076) );
XNOR2_X1 U927 ( .A(KEYINPUT45), .B(n1203), .ZN(n1239) );
XOR2_X1 U928 ( .A(n1241), .B(n1242), .Z(n1203) );
XOR2_X1 U929 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U930 ( .A(n1245), .B(G125), .Z(n1244) );
NAND2_X1 U931 ( .A1(KEYINPUT14), .A2(n1119), .ZN(n1245) );
XOR2_X1 U932 ( .A(n1156), .B(n1246), .Z(n1119) );
INV_X1 U933 ( .A(G110), .ZN(n1156) );
NAND2_X1 U934 ( .A1(G224), .A2(n1247), .ZN(n1243) );
XNOR2_X1 U935 ( .A(n1118), .B(n1097), .ZN(n1241) );
XNOR2_X1 U936 ( .A(n1248), .B(n1249), .ZN(n1118) );
XOR2_X1 U937 ( .A(KEYINPUT16), .B(n1250), .Z(n1249) );
AND4_X1 U938 ( .A1(n1190), .A2(n1191), .A3(n1035), .A4(n1251), .ZN(n1193) );
NOR2_X1 U939 ( .A1(n1033), .A2(n1048), .ZN(n1251) );
INV_X1 U940 ( .A(n1023), .ZN(n1048) );
XOR2_X1 U941 ( .A(n1252), .B(n1123), .Z(n1023) );
INV_X1 U942 ( .A(n1067), .ZN(n1123) );
NAND2_X1 U943 ( .A1(n1126), .A2(n1240), .ZN(n1067) );
NAND2_X1 U944 ( .A1(n1253), .A2(n1254), .ZN(n1126) );
OR2_X1 U945 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XOR2_X1 U946 ( .A(n1257), .B(KEYINPUT4), .Z(n1253) );
NAND2_X1 U947 ( .A1(n1256), .A2(n1255), .ZN(n1257) );
XNOR2_X1 U948 ( .A(n1258), .B(n1259), .ZN(n1255) );
XOR2_X1 U949 ( .A(KEYINPUT23), .B(G137), .Z(n1259) );
NAND2_X1 U950 ( .A1(G221), .A2(n1260), .ZN(n1258) );
XNOR2_X1 U951 ( .A(n1261), .B(n1262), .ZN(n1256) );
XOR2_X1 U952 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U953 ( .A(G119), .B(n1265), .ZN(n1261) );
XOR2_X1 U954 ( .A(KEYINPUT38), .B(G128), .Z(n1265) );
NAND2_X1 U955 ( .A1(KEYINPUT30), .A2(n1068), .ZN(n1252) );
NAND2_X1 U956 ( .A1(G217), .A2(n1266), .ZN(n1068) );
INV_X1 U957 ( .A(n1180), .ZN(n1033) );
NOR2_X1 U958 ( .A1(n1227), .A2(n1064), .ZN(n1180) );
INV_X1 U959 ( .A(n1229), .ZN(n1064) );
XOR2_X1 U960 ( .A(n1267), .B(G475), .Z(n1229) );
NAND2_X1 U961 ( .A1(n1137), .A2(n1268), .ZN(n1267) );
XOR2_X1 U962 ( .A(KEYINPUT6), .B(G902), .Z(n1268) );
XOR2_X1 U963 ( .A(n1269), .B(n1270), .Z(n1137) );
NOR2_X1 U964 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XOR2_X1 U965 ( .A(n1273), .B(KEYINPUT19), .Z(n1272) );
NAND2_X1 U966 ( .A1(G104), .A2(n1274), .ZN(n1273) );
NOR2_X1 U967 ( .A1(G104), .A2(n1274), .ZN(n1271) );
XOR2_X1 U968 ( .A(n1275), .B(n1276), .Z(n1274) );
XOR2_X1 U969 ( .A(KEYINPUT40), .B(n1277), .Z(n1276) );
INV_X1 U970 ( .A(n1246), .ZN(n1275) );
NAND2_X1 U971 ( .A1(KEYINPUT8), .A2(n1278), .ZN(n1269) );
XNOR2_X1 U972 ( .A(n1264), .B(n1279), .ZN(n1278) );
XOR2_X1 U973 ( .A(n1280), .B(G140), .Z(n1279) );
NAND2_X1 U974 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
OR2_X1 U975 ( .A1(n1101), .A2(n1283), .ZN(n1282) );
XOR2_X1 U976 ( .A(n1284), .B(KEYINPUT7), .Z(n1281) );
NAND2_X1 U977 ( .A1(n1283), .A2(n1101), .ZN(n1284) );
INV_X1 U978 ( .A(G131), .ZN(n1101) );
XNOR2_X1 U979 ( .A(n1285), .B(G143), .ZN(n1283) );
NAND2_X1 U980 ( .A1(G214), .A2(n1286), .ZN(n1285) );
XOR2_X1 U981 ( .A(G146), .B(G125), .Z(n1264) );
NAND3_X1 U982 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n1227) );
INV_X1 U983 ( .A(n1073), .ZN(n1289) );
NOR2_X1 U984 ( .A1(n1074), .A2(G478), .ZN(n1073) );
NAND2_X1 U985 ( .A1(KEYINPUT22), .A2(n1134), .ZN(n1288) );
INV_X1 U986 ( .A(G478), .ZN(n1134) );
NAND3_X1 U987 ( .A1(n1074), .A2(n1290), .A3(G478), .ZN(n1287) );
INV_X1 U988 ( .A(KEYINPUT22), .ZN(n1290) );
NAND2_X1 U989 ( .A1(n1132), .A2(n1240), .ZN(n1074) );
XNOR2_X1 U990 ( .A(n1291), .B(n1292), .ZN(n1132) );
XOR2_X1 U991 ( .A(n1293), .B(n1246), .Z(n1292) );
XNOR2_X1 U992 ( .A(G122), .B(KEYINPUT56), .ZN(n1246) );
NAND2_X1 U993 ( .A1(G217), .A2(n1260), .ZN(n1293) );
AND2_X1 U994 ( .A1(G234), .A2(n1247), .ZN(n1260) );
XOR2_X1 U995 ( .A(n1294), .B(n1295), .Z(n1291) );
NOR2_X1 U996 ( .A1(KEYINPUT53), .A2(n1296), .ZN(n1295) );
XOR2_X1 U997 ( .A(G134), .B(n1297), .Z(n1296) );
XOR2_X1 U998 ( .A(n1011), .B(G116), .Z(n1294) );
INV_X1 U999 ( .A(G107), .ZN(n1011) );
AND2_X1 U1000 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U1001 ( .A1(G221), .A2(n1266), .ZN(n1037) );
NAND2_X1 U1002 ( .A1(G234), .A2(n1237), .ZN(n1266) );
XOR2_X1 U1003 ( .A(G902), .B(KEYINPUT52), .Z(n1237) );
XNOR2_X1 U1004 ( .A(n1069), .B(G469), .ZN(n1036) );
NAND2_X1 U1005 ( .A1(n1298), .A2(n1240), .ZN(n1069) );
XOR2_X1 U1006 ( .A(n1299), .B(n1300), .Z(n1298) );
XNOR2_X1 U1007 ( .A(n1164), .B(n1263), .ZN(n1300) );
XOR2_X1 U1008 ( .A(G110), .B(G140), .Z(n1263) );
XOR2_X1 U1009 ( .A(n1097), .B(n1162), .Z(n1164) );
INV_X1 U1010 ( .A(n1248), .ZN(n1162) );
XOR2_X1 U1011 ( .A(n1301), .B(n1302), .Z(n1248) );
XOR2_X1 U1012 ( .A(G104), .B(G101), .Z(n1302) );
XOR2_X1 U1013 ( .A(n1303), .B(G107), .Z(n1301) );
XNOR2_X1 U1014 ( .A(KEYINPUT58), .B(KEYINPUT46), .ZN(n1303) );
XOR2_X1 U1015 ( .A(n1304), .B(n1305), .Z(n1299) );
NOR2_X1 U1016 ( .A1(KEYINPUT62), .A2(n1150), .ZN(n1305) );
XOR2_X1 U1017 ( .A(n1153), .B(KEYINPUT44), .Z(n1304) );
NAND2_X1 U1018 ( .A1(G227), .A2(n1247), .ZN(n1153) );
NAND2_X1 U1019 ( .A1(n1224), .A2(n1306), .ZN(n1191) );
NAND3_X1 U1020 ( .A1(G902), .A2(n1050), .A3(n1117), .ZN(n1306) );
NOR2_X1 U1021 ( .A1(n1307), .A2(G898), .ZN(n1117) );
INV_X1 U1022 ( .A(n1094), .ZN(n1307) );
XOR2_X1 U1023 ( .A(n1046), .B(KEYINPUT28), .Z(n1094) );
NAND3_X1 U1024 ( .A1(n1050), .A2(n1046), .A3(n1308), .ZN(n1224) );
XNOR2_X1 U1025 ( .A(G952), .B(KEYINPUT55), .ZN(n1308) );
NAND2_X1 U1026 ( .A1(G237), .A2(G234), .ZN(n1050) );
INV_X1 U1027 ( .A(n1028), .ZN(n1190) );
XNOR2_X1 U1028 ( .A(n1309), .B(n1066), .ZN(n1028) );
NAND2_X1 U1029 ( .A1(n1310), .A2(n1240), .ZN(n1066) );
INV_X1 U1030 ( .A(G902), .ZN(n1240) );
XNOR2_X1 U1031 ( .A(n1311), .B(n1144), .ZN(n1310) );
XNOR2_X1 U1032 ( .A(n1312), .B(n1250), .ZN(n1144) );
XNOR2_X1 U1033 ( .A(n1313), .B(n1277), .ZN(n1250) );
XOR2_X1 U1034 ( .A(G113), .B(KEYINPUT0), .Z(n1277) );
XNOR2_X1 U1035 ( .A(G116), .B(G119), .ZN(n1313) );
XOR2_X1 U1036 ( .A(n1150), .B(n1097), .Z(n1312) );
XOR2_X1 U1037 ( .A(G146), .B(n1297), .Z(n1097) );
XOR2_X1 U1038 ( .A(G128), .B(G143), .Z(n1297) );
NAND2_X1 U1039 ( .A1(n1314), .A2(n1315), .ZN(n1150) );
OR2_X1 U1040 ( .A1(n1104), .A2(G131), .ZN(n1315) );
XOR2_X1 U1041 ( .A(n1316), .B(KEYINPUT48), .Z(n1314) );
NAND2_X1 U1042 ( .A1(G131), .A2(n1104), .ZN(n1316) );
XOR2_X1 U1043 ( .A(G137), .B(G134), .Z(n1104) );
NAND2_X1 U1044 ( .A1(n1317), .A2(n1318), .ZN(n1311) );
NAND2_X1 U1045 ( .A1(n1145), .A2(n1221), .ZN(n1318) );
XOR2_X1 U1046 ( .A(KEYINPUT60), .B(n1319), .Z(n1317) );
NOR2_X1 U1047 ( .A1(n1221), .A2(n1145), .ZN(n1319) );
NAND2_X1 U1048 ( .A1(G210), .A2(n1286), .ZN(n1145) );
AND2_X1 U1049 ( .A1(n1247), .A2(n1238), .ZN(n1286) );
INV_X1 U1050 ( .A(G237), .ZN(n1238) );
XOR2_X1 U1051 ( .A(n1046), .B(KEYINPUT13), .Z(n1247) );
INV_X1 U1052 ( .A(G953), .ZN(n1046) );
INV_X1 U1053 ( .A(G101), .ZN(n1221) );
NAND2_X1 U1054 ( .A1(KEYINPUT2), .A2(n1320), .ZN(n1309) );
XOR2_X1 U1055 ( .A(KEYINPUT50), .B(G472), .Z(n1320) );
endmodule


