//Key = 1101010001111001100001000110100001110100000001011001101110111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324;

XOR2_X1 U727 ( .A(n1013), .B(G107), .Z(G9) );
NAND2_X1 U728 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND2_X1 U729 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
INV_X1 U730 ( .A(KEYINPUT39), .ZN(n1017) );
NAND3_X1 U731 ( .A1(n1018), .A2(n1019), .A3(KEYINPUT39), .ZN(n1014) );
NOR2_X1 U732 ( .A1(n1020), .A2(n1021), .ZN(G75) );
NOR4_X1 U733 ( .A1(G953), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1021) );
NOR2_X1 U734 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U735 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR2_X1 U736 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
INV_X1 U737 ( .A(n1031), .ZN(n1030) );
NOR2_X1 U738 ( .A1(n1032), .A2(n1033), .ZN(n1029) );
NOR2_X1 U739 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR3_X1 U740 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1032) );
NOR2_X1 U741 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR4_X1 U742 ( .A1(n1041), .A2(n1042), .A3(n1035), .A4(n1036), .ZN(n1027) );
INV_X1 U743 ( .A(n1043), .ZN(n1036) );
INV_X1 U744 ( .A(n1044), .ZN(n1035) );
NOR3_X1 U745 ( .A1(n1037), .A2(n1045), .A3(n1046), .ZN(n1042) );
NOR2_X1 U746 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U747 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U748 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U749 ( .A1(n1053), .A2(n1054), .ZN(n1045) );
NOR2_X1 U750 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U751 ( .A1(n1031), .A2(n1057), .ZN(n1041) );
NOR3_X1 U752 ( .A1(n1022), .A2(G953), .A3(G952), .ZN(n1020) );
AND4_X1 U753 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1022) );
NOR4_X1 U754 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1061) );
XNOR2_X1 U755 ( .A(n1066), .B(n1067), .ZN(n1065) );
XNOR2_X1 U756 ( .A(n1068), .B(n1069), .ZN(n1064) );
XOR2_X1 U757 ( .A(KEYINPUT20), .B(n1070), .Z(n1063) );
NOR3_X1 U758 ( .A1(n1071), .A2(n1072), .A3(n1037), .ZN(n1060) );
NAND2_X1 U759 ( .A1(n1073), .A2(n1074), .ZN(n1059) );
XNOR2_X1 U760 ( .A(G469), .B(KEYINPUT52), .ZN(n1073) );
NAND2_X1 U761 ( .A1(n1075), .A2(n1076), .ZN(G72) );
NAND2_X1 U762 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U763 ( .A1(G953), .A2(n1079), .ZN(n1078) );
NAND2_X1 U764 ( .A1(G900), .A2(G227), .ZN(n1079) );
NAND2_X1 U765 ( .A1(n1080), .A2(n1081), .ZN(n1075) );
NAND2_X1 U766 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U767 ( .A1(G953), .A2(n1084), .ZN(n1083) );
INV_X1 U768 ( .A(n1085), .ZN(n1082) );
INV_X1 U769 ( .A(n1077), .ZN(n1080) );
XNOR2_X1 U770 ( .A(n1086), .B(n1087), .ZN(n1077) );
NOR2_X1 U771 ( .A1(n1085), .A2(n1088), .ZN(n1087) );
XOR2_X1 U772 ( .A(n1089), .B(n1090), .Z(n1088) );
XOR2_X1 U773 ( .A(n1091), .B(n1092), .Z(n1090) );
XNOR2_X1 U774 ( .A(n1093), .B(G131), .ZN(n1092) );
NOR2_X1 U775 ( .A1(KEYINPUT50), .A2(n1094), .ZN(n1091) );
XNOR2_X1 U776 ( .A(n1095), .B(n1096), .ZN(n1094) );
NOR2_X1 U777 ( .A1(G125), .A2(KEYINPUT18), .ZN(n1096) );
XNOR2_X1 U778 ( .A(n1097), .B(n1098), .ZN(n1089) );
NAND2_X1 U779 ( .A1(KEYINPUT45), .A2(n1099), .ZN(n1098) );
NAND2_X1 U780 ( .A1(KEYINPUT12), .A2(n1100), .ZN(n1097) );
NAND2_X1 U781 ( .A1(n1101), .A2(n1102), .ZN(n1086) );
NAND2_X1 U782 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U783 ( .A(KEYINPUT54), .B(n1105), .ZN(n1101) );
XOR2_X1 U784 ( .A(n1106), .B(n1107), .Z(G69) );
XOR2_X1 U785 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U786 ( .A1(G953), .A2(n1110), .ZN(n1109) );
NAND2_X1 U787 ( .A1(G898), .A2(G224), .ZN(n1110) );
NAND3_X1 U788 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1108) );
XOR2_X1 U789 ( .A(n1114), .B(KEYINPUT41), .Z(n1113) );
NAND2_X1 U790 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U791 ( .A1(n1117), .A2(n1118), .ZN(n1112) );
XNOR2_X1 U792 ( .A(KEYINPUT40), .B(n1105), .ZN(n1117) );
OR2_X1 U793 ( .A1(n1116), .A2(n1115), .ZN(n1111) );
NOR2_X1 U794 ( .A1(n1119), .A2(G953), .ZN(n1106) );
NOR2_X1 U795 ( .A1(n1120), .A2(n1121), .ZN(G66) );
XOR2_X1 U796 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U797 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
NOR2_X1 U798 ( .A1(n1126), .A2(n1127), .ZN(G63) );
XNOR2_X1 U799 ( .A(n1120), .B(KEYINPUT1), .ZN(n1127) );
NOR3_X1 U800 ( .A1(n1067), .A2(n1128), .A3(n1129), .ZN(n1126) );
AND3_X1 U801 ( .A1(n1130), .A2(G478), .A3(n1131), .ZN(n1129) );
NOR2_X1 U802 ( .A1(n1132), .A2(n1130), .ZN(n1128) );
AND2_X1 U803 ( .A1(n1024), .A2(G478), .ZN(n1132) );
NOR2_X1 U804 ( .A1(n1120), .A2(n1133), .ZN(G60) );
XOR2_X1 U805 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND3_X1 U806 ( .A1(n1131), .A2(G475), .A3(KEYINPUT10), .ZN(n1134) );
XOR2_X1 U807 ( .A(G104), .B(n1136), .Z(G6) );
NOR2_X1 U808 ( .A1(n1120), .A2(n1137), .ZN(G57) );
XOR2_X1 U809 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U810 ( .A1(KEYINPUT30), .A2(n1140), .ZN(n1139) );
XOR2_X1 U811 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U812 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U813 ( .A1(KEYINPUT53), .A2(n1145), .ZN(n1143) );
XNOR2_X1 U814 ( .A(n1146), .B(n1147), .ZN(n1141) );
NAND3_X1 U815 ( .A1(n1131), .A2(G472), .A3(KEYINPUT63), .ZN(n1146) );
NOR2_X1 U816 ( .A1(n1148), .A2(n1149), .ZN(n1138) );
NOR2_X1 U817 ( .A1(n1120), .A2(n1150), .ZN(G54) );
XOR2_X1 U818 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U819 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U820 ( .A1(KEYINPUT7), .A2(n1155), .ZN(n1154) );
AND2_X1 U821 ( .A1(G469), .A2(n1131), .ZN(n1153) );
INV_X1 U822 ( .A(n1125), .ZN(n1131) );
XNOR2_X1 U823 ( .A(n1156), .B(n1145), .ZN(n1151) );
INV_X1 U824 ( .A(n1157), .ZN(n1145) );
NOR2_X1 U825 ( .A1(n1120), .A2(n1158), .ZN(G51) );
XOR2_X1 U826 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U827 ( .A1(n1069), .A2(n1125), .ZN(n1160) );
NAND2_X1 U828 ( .A1(G902), .A2(n1024), .ZN(n1125) );
NAND3_X1 U829 ( .A1(n1119), .A2(n1103), .A3(n1161), .ZN(n1024) );
XOR2_X1 U830 ( .A(n1104), .B(KEYINPUT46), .Z(n1161) );
AND4_X1 U831 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1103) );
NOR4_X1 U832 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
NAND2_X1 U833 ( .A1(n1170), .A2(n1171), .ZN(n1164) );
AND4_X1 U834 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1119) );
NOR4_X1 U835 ( .A1(n1176), .A2(n1136), .A3(n1016), .A4(n1177), .ZN(n1175) );
AND2_X1 U836 ( .A1(n1055), .A2(n1018), .ZN(n1016) );
AND2_X1 U837 ( .A1(n1056), .A2(n1018), .ZN(n1136) );
AND2_X1 U838 ( .A1(n1044), .A2(n1178), .ZN(n1018) );
INV_X1 U839 ( .A(n1179), .ZN(n1176) );
NOR2_X1 U840 ( .A1(n1180), .A2(n1181), .ZN(n1174) );
NAND2_X1 U841 ( .A1(n1182), .A2(n1183), .ZN(n1159) );
NAND2_X1 U842 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NAND2_X1 U843 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NAND2_X1 U844 ( .A1(KEYINPUT62), .A2(n1188), .ZN(n1187) );
INV_X1 U845 ( .A(KEYINPUT4), .ZN(n1186) );
NAND2_X1 U846 ( .A1(n1189), .A2(n1190), .ZN(n1182) );
NAND2_X1 U847 ( .A1(KEYINPUT62), .A2(n1191), .ZN(n1190) );
OR2_X1 U848 ( .A1(n1184), .A2(KEYINPUT4), .ZN(n1191) );
NOR2_X1 U849 ( .A1(n1105), .A2(G952), .ZN(n1120) );
XNOR2_X1 U850 ( .A(n1192), .B(n1162), .ZN(G48) );
NAND3_X1 U851 ( .A1(n1056), .A2(n1050), .A3(n1193), .ZN(n1162) );
XNOR2_X1 U852 ( .A(G146), .B(KEYINPUT35), .ZN(n1192) );
XOR2_X1 U853 ( .A(n1163), .B(n1194), .Z(G45) );
XNOR2_X1 U854 ( .A(G143), .B(KEYINPUT29), .ZN(n1194) );
NAND4_X1 U855 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1163) );
XNOR2_X1 U856 ( .A(G140), .B(n1199), .ZN(G42) );
NAND2_X1 U857 ( .A1(KEYINPUT11), .A2(n1168), .ZN(n1199) );
AND3_X1 U858 ( .A1(n1056), .A2(n1039), .A3(n1170), .ZN(n1168) );
XNOR2_X1 U859 ( .A(G137), .B(n1104), .ZN(G39) );
NAND2_X1 U860 ( .A1(n1031), .A2(n1193), .ZN(n1104) );
NOR2_X1 U861 ( .A1(n1054), .A2(n1048), .ZN(n1031) );
INV_X1 U862 ( .A(n1200), .ZN(n1048) );
XNOR2_X1 U863 ( .A(G134), .B(n1201), .ZN(G36) );
NAND4_X1 U864 ( .A1(n1202), .A2(n1203), .A3(n1171), .A4(n1198), .ZN(n1201) );
XNOR2_X1 U865 ( .A(n1204), .B(KEYINPUT37), .ZN(n1202) );
XOR2_X1 U866 ( .A(G131), .B(n1167), .Z(G33) );
AND3_X1 U867 ( .A1(n1056), .A2(n1040), .A3(n1170), .ZN(n1167) );
NOR3_X1 U868 ( .A1(n1034), .A2(n1205), .A3(n1054), .ZN(n1170) );
INV_X1 U869 ( .A(n1203), .ZN(n1054) );
NOR2_X1 U870 ( .A1(n1206), .A2(n1051), .ZN(n1203) );
XOR2_X1 U871 ( .A(n1207), .B(n1166), .Z(G30) );
AND3_X1 U872 ( .A1(n1055), .A2(n1050), .A3(n1193), .ZN(n1166) );
NOR4_X1 U873 ( .A1(n1208), .A2(n1034), .A3(n1058), .A4(n1205), .ZN(n1193) );
INV_X1 U874 ( .A(n1198), .ZN(n1205) );
INV_X1 U875 ( .A(n1204), .ZN(n1034) );
XNOR2_X1 U876 ( .A(G128), .B(KEYINPUT9), .ZN(n1207) );
NAND2_X1 U877 ( .A1(n1209), .A2(n1210), .ZN(G3) );
NAND2_X1 U878 ( .A1(G101), .A2(n1211), .ZN(n1210) );
XOR2_X1 U879 ( .A(n1212), .B(KEYINPUT14), .Z(n1209) );
NAND2_X1 U880 ( .A1(n1177), .A2(n1213), .ZN(n1212) );
INV_X1 U881 ( .A(n1211), .ZN(n1177) );
NAND3_X1 U882 ( .A1(n1200), .A2(n1214), .A3(n1196), .ZN(n1211) );
AND3_X1 U883 ( .A1(n1204), .A2(n1050), .A3(n1040), .ZN(n1196) );
XOR2_X1 U884 ( .A(G125), .B(n1169), .Z(G27) );
AND4_X1 U885 ( .A1(n1043), .A2(n1039), .A3(n1056), .A4(n1215), .ZN(n1169) );
AND3_X1 U886 ( .A1(n1050), .A2(n1057), .A3(n1198), .ZN(n1215) );
NAND2_X1 U887 ( .A1(n1026), .A2(n1216), .ZN(n1198) );
NAND3_X1 U888 ( .A1(G902), .A2(n1217), .A3(n1085), .ZN(n1216) );
NOR2_X1 U889 ( .A1(n1105), .A2(G900), .ZN(n1085) );
XNOR2_X1 U890 ( .A(G122), .B(n1179), .ZN(G24) );
NAND4_X1 U891 ( .A1(n1195), .A2(n1218), .A3(n1197), .A4(n1044), .ZN(n1179) );
NOR2_X1 U892 ( .A1(n1219), .A2(n1220), .ZN(n1044) );
XNOR2_X1 U893 ( .A(n1062), .B(KEYINPUT28), .ZN(n1195) );
XOR2_X1 U894 ( .A(n1172), .B(n1221), .Z(G21) );
NAND2_X1 U895 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
XNOR2_X1 U896 ( .A(G119), .B(KEYINPUT33), .ZN(n1223) );
XNOR2_X1 U897 ( .A(KEYINPUT59), .B(KEYINPUT55), .ZN(n1222) );
NAND4_X1 U898 ( .A1(n1218), .A2(n1200), .A3(n1220), .A4(n1219), .ZN(n1172) );
XNOR2_X1 U899 ( .A(G116), .B(n1173), .ZN(G18) );
NAND2_X1 U900 ( .A1(n1171), .A2(n1218), .ZN(n1173) );
AND2_X1 U901 ( .A1(n1040), .A2(n1055), .ZN(n1171) );
INV_X1 U902 ( .A(n1019), .ZN(n1055) );
NAND2_X1 U903 ( .A1(n1197), .A2(n1224), .ZN(n1019) );
XNOR2_X1 U904 ( .A(n1225), .B(n1181), .ZN(G15) );
AND3_X1 U905 ( .A1(n1040), .A2(n1218), .A3(n1056), .ZN(n1181) );
NOR2_X1 U906 ( .A1(n1224), .A2(n1197), .ZN(n1056) );
INV_X1 U907 ( .A(n1062), .ZN(n1224) );
AND4_X1 U908 ( .A1(n1043), .A2(n1050), .A3(n1214), .A4(n1057), .ZN(n1218) );
NOR2_X1 U909 ( .A1(n1058), .A2(n1220), .ZN(n1040) );
INV_X1 U910 ( .A(n1208), .ZN(n1220) );
INV_X1 U911 ( .A(n1219), .ZN(n1058) );
NAND2_X1 U912 ( .A1(n1226), .A2(n1227), .ZN(G12) );
NAND2_X1 U913 ( .A1(n1180), .A2(n1228), .ZN(n1227) );
XOR2_X1 U914 ( .A(KEYINPUT48), .B(n1229), .Z(n1226) );
NOR2_X1 U915 ( .A1(n1180), .A2(n1228), .ZN(n1229) );
INV_X1 U916 ( .A(G110), .ZN(n1228) );
AND3_X1 U917 ( .A1(n1039), .A2(n1178), .A3(n1200), .ZN(n1180) );
NOR2_X1 U918 ( .A1(n1062), .A2(n1197), .ZN(n1200) );
XOR2_X1 U919 ( .A(n1230), .B(n1067), .Z(n1197) );
NOR2_X1 U920 ( .A1(n1130), .A2(G902), .ZN(n1067) );
XNOR2_X1 U921 ( .A(n1231), .B(n1232), .ZN(n1130) );
XOR2_X1 U922 ( .A(n1233), .B(n1234), .Z(n1232) );
XNOR2_X1 U923 ( .A(G134), .B(n1235), .ZN(n1234) );
NAND2_X1 U924 ( .A1(KEYINPUT0), .A2(n1236), .ZN(n1235) );
NAND3_X1 U925 ( .A1(G234), .A2(n1105), .A3(G217), .ZN(n1236) );
NOR2_X1 U926 ( .A1(n1237), .A2(n1238), .ZN(n1233) );
XOR2_X1 U927 ( .A(KEYINPUT13), .B(n1239), .Z(n1238) );
AND2_X1 U928 ( .A1(n1240), .A2(G116), .ZN(n1239) );
NOR2_X1 U929 ( .A1(G116), .A2(n1240), .ZN(n1237) );
XNOR2_X1 U930 ( .A(n1241), .B(n1242), .ZN(n1231) );
NAND2_X1 U931 ( .A1(KEYINPUT21), .A2(n1066), .ZN(n1230) );
INV_X1 U932 ( .A(G478), .ZN(n1066) );
XNOR2_X1 U933 ( .A(n1243), .B(n1244), .ZN(n1062) );
XOR2_X1 U934 ( .A(KEYINPUT6), .B(G475), .Z(n1244) );
NAND2_X1 U935 ( .A1(n1135), .A2(n1245), .ZN(n1243) );
XOR2_X1 U936 ( .A(n1246), .B(n1247), .Z(n1135) );
XOR2_X1 U937 ( .A(n1248), .B(n1249), .Z(n1247) );
XNOR2_X1 U938 ( .A(G131), .B(n1240), .ZN(n1249) );
INV_X1 U939 ( .A(G122), .ZN(n1240) );
XNOR2_X1 U940 ( .A(KEYINPUT23), .B(n1250), .ZN(n1248) );
XOR2_X1 U941 ( .A(n1251), .B(n1252), .Z(n1246) );
XOR2_X1 U942 ( .A(n1253), .B(n1254), .Z(n1251) );
NAND3_X1 U943 ( .A1(n1255), .A2(G214), .A3(n1256), .ZN(n1253) );
XNOR2_X1 U944 ( .A(G953), .B(KEYINPUT19), .ZN(n1256) );
AND3_X1 U945 ( .A1(n1050), .A2(n1214), .A3(n1204), .ZN(n1178) );
NOR2_X1 U946 ( .A1(n1037), .A2(n1043), .ZN(n1204) );
NOR2_X1 U947 ( .A1(n1257), .A2(n1072), .ZN(n1043) );
NOR2_X1 U948 ( .A1(n1074), .A2(G469), .ZN(n1072) );
AND2_X1 U949 ( .A1(n1258), .A2(G469), .ZN(n1257) );
XOR2_X1 U950 ( .A(n1074), .B(KEYINPUT49), .Z(n1258) );
NAND2_X1 U951 ( .A1(n1259), .A2(n1245), .ZN(n1074) );
XNOR2_X1 U952 ( .A(n1155), .B(n1260), .ZN(n1259) );
XOR2_X1 U953 ( .A(n1156), .B(n1261), .Z(n1260) );
NOR2_X1 U954 ( .A1(KEYINPUT8), .A2(n1157), .ZN(n1261) );
XOR2_X1 U955 ( .A(n1262), .B(n1263), .Z(n1156) );
XNOR2_X1 U956 ( .A(n1095), .B(n1264), .ZN(n1263) );
NOR2_X1 U957 ( .A1(G953), .A2(n1084), .ZN(n1264) );
INV_X1 U958 ( .A(G227), .ZN(n1084) );
INV_X1 U959 ( .A(G140), .ZN(n1095) );
XOR2_X1 U960 ( .A(n1099), .B(n1265), .Z(n1262) );
XNOR2_X1 U961 ( .A(n1266), .B(n1267), .ZN(n1099) );
XNOR2_X1 U962 ( .A(n1268), .B(n1269), .ZN(n1267) );
NOR2_X1 U963 ( .A1(KEYINPUT17), .A2(n1270), .ZN(n1269) );
XNOR2_X1 U964 ( .A(KEYINPUT51), .B(G143), .ZN(n1270) );
XOR2_X1 U965 ( .A(G104), .B(n1271), .Z(n1155) );
INV_X1 U966 ( .A(n1057), .ZN(n1037) );
NAND2_X1 U967 ( .A1(G221), .A2(n1272), .ZN(n1057) );
NAND2_X1 U968 ( .A1(n1026), .A2(n1273), .ZN(n1214) );
NAND4_X1 U969 ( .A1(G953), .A2(G902), .A3(n1217), .A4(n1118), .ZN(n1273) );
INV_X1 U970 ( .A(G898), .ZN(n1118) );
NAND3_X1 U971 ( .A1(n1217), .A2(n1105), .A3(G952), .ZN(n1026) );
NAND2_X1 U972 ( .A1(G237), .A2(G234), .ZN(n1217) );
NOR2_X1 U973 ( .A1(n1274), .A2(n1206), .ZN(n1050) );
XOR2_X1 U974 ( .A(n1071), .B(KEYINPUT2), .Z(n1206) );
INV_X1 U975 ( .A(n1052), .ZN(n1071) );
NAND2_X1 U976 ( .A1(G214), .A2(n1275), .ZN(n1052) );
INV_X1 U977 ( .A(n1051), .ZN(n1274) );
XOR2_X1 U978 ( .A(n1276), .B(n1068), .Z(n1051) );
AND2_X1 U979 ( .A1(n1277), .A2(n1245), .ZN(n1068) );
XOR2_X1 U980 ( .A(n1278), .B(n1184), .Z(n1277) );
XOR2_X1 U981 ( .A(n1115), .B(n1279), .Z(n1184) );
NOR2_X1 U982 ( .A1(KEYINPUT24), .A2(n1116), .ZN(n1279) );
XNOR2_X1 U983 ( .A(n1280), .B(n1281), .ZN(n1116) );
XOR2_X1 U984 ( .A(G116), .B(n1282), .Z(n1281) );
XNOR2_X1 U985 ( .A(KEYINPUT57), .B(n1283), .ZN(n1282) );
INV_X1 U986 ( .A(G119), .ZN(n1283) );
XNOR2_X1 U987 ( .A(n1252), .B(n1271), .ZN(n1280) );
XNOR2_X1 U988 ( .A(n1284), .B(n1241), .ZN(n1271) );
XOR2_X1 U989 ( .A(G107), .B(KEYINPUT58), .Z(n1241) );
XNOR2_X1 U990 ( .A(G101), .B(KEYINPUT56), .ZN(n1284) );
XNOR2_X1 U991 ( .A(G104), .B(n1225), .ZN(n1252) );
XNOR2_X1 U992 ( .A(G122), .B(n1285), .ZN(n1115) );
NOR2_X1 U993 ( .A1(KEYINPUT32), .A2(n1265), .ZN(n1285) );
NAND2_X1 U994 ( .A1(KEYINPUT34), .A2(n1189), .ZN(n1278) );
INV_X1 U995 ( .A(n1188), .ZN(n1189) );
XNOR2_X1 U996 ( .A(n1286), .B(n1144), .ZN(n1188) );
XNOR2_X1 U997 ( .A(G125), .B(n1287), .ZN(n1286) );
AND2_X1 U998 ( .A1(n1105), .A2(G224), .ZN(n1287) );
NAND2_X1 U999 ( .A1(KEYINPUT60), .A2(n1069), .ZN(n1276) );
NAND2_X1 U1000 ( .A1(G210), .A2(n1275), .ZN(n1069) );
NAND2_X1 U1001 ( .A1(n1288), .A2(n1245), .ZN(n1275) );
INV_X1 U1002 ( .A(G237), .ZN(n1288) );
NOR2_X1 U1003 ( .A1(n1208), .A2(n1219), .ZN(n1039) );
XNOR2_X1 U1004 ( .A(n1289), .B(G472), .ZN(n1219) );
NAND2_X1 U1005 ( .A1(n1290), .A2(n1245), .ZN(n1289) );
XOR2_X1 U1006 ( .A(n1291), .B(n1292), .Z(n1290) );
XOR2_X1 U1007 ( .A(n1293), .B(n1294), .Z(n1292) );
NOR2_X1 U1008 ( .A1(KEYINPUT43), .A2(n1157), .ZN(n1294) );
XNOR2_X1 U1009 ( .A(n1295), .B(n1296), .ZN(n1157) );
XNOR2_X1 U1010 ( .A(n1100), .B(G131), .ZN(n1296) );
INV_X1 U1011 ( .A(G134), .ZN(n1100) );
NAND2_X1 U1012 ( .A1(KEYINPUT5), .A2(n1093), .ZN(n1295) );
INV_X1 U1013 ( .A(G137), .ZN(n1093) );
NOR2_X1 U1014 ( .A1(n1149), .A2(n1297), .ZN(n1293) );
XNOR2_X1 U1015 ( .A(n1148), .B(KEYINPUT47), .ZN(n1297) );
AND4_X1 U1016 ( .A1(G101), .A2(G210), .A3(n1255), .A4(n1105), .ZN(n1148) );
AND2_X1 U1017 ( .A1(n1213), .A2(n1298), .ZN(n1149) );
NAND3_X1 U1018 ( .A1(n1255), .A2(n1105), .A3(G210), .ZN(n1298) );
XNOR2_X1 U1019 ( .A(G237), .B(KEYINPUT44), .ZN(n1255) );
INV_X1 U1020 ( .A(G101), .ZN(n1213) );
NAND2_X1 U1021 ( .A1(n1299), .A2(n1300), .ZN(n1291) );
NAND2_X1 U1022 ( .A1(n1301), .A2(n1147), .ZN(n1300) );
XOR2_X1 U1023 ( .A(KEYINPUT27), .B(n1144), .Z(n1301) );
NAND2_X1 U1024 ( .A1(n1302), .A2(n1303), .ZN(n1299) );
INV_X1 U1025 ( .A(n1147), .ZN(n1303) );
NAND2_X1 U1026 ( .A1(n1304), .A2(n1305), .ZN(n1147) );
NAND2_X1 U1027 ( .A1(n1306), .A2(n1225), .ZN(n1305) );
XOR2_X1 U1028 ( .A(KEYINPUT16), .B(n1307), .Z(n1304) );
NOR2_X1 U1029 ( .A1(n1225), .A2(n1306), .ZN(n1307) );
XOR2_X1 U1030 ( .A(G116), .B(n1308), .Z(n1306) );
NOR2_X1 U1031 ( .A1(G119), .A2(KEYINPUT42), .ZN(n1308) );
INV_X1 U1032 ( .A(G113), .ZN(n1225) );
XOR2_X1 U1033 ( .A(KEYINPUT3), .B(n1144), .Z(n1302) );
XOR2_X1 U1034 ( .A(n1242), .B(n1309), .Z(n1144) );
XOR2_X1 U1035 ( .A(KEYINPUT51), .B(n1310), .Z(n1309) );
NOR2_X1 U1036 ( .A1(KEYINPUT22), .A2(n1266), .ZN(n1310) );
XNOR2_X1 U1037 ( .A(G128), .B(n1250), .ZN(n1242) );
INV_X1 U1038 ( .A(G143), .ZN(n1250) );
XOR2_X1 U1039 ( .A(n1070), .B(KEYINPUT25), .Z(n1208) );
XOR2_X1 U1040 ( .A(n1311), .B(n1124), .Z(n1070) );
NAND2_X1 U1041 ( .A1(G217), .A2(n1272), .ZN(n1124) );
NAND2_X1 U1042 ( .A1(G234), .A2(n1245), .ZN(n1272) );
INV_X1 U1043 ( .A(G902), .ZN(n1245) );
OR2_X1 U1044 ( .A1(n1123), .A2(G902), .ZN(n1311) );
XNOR2_X1 U1045 ( .A(n1312), .B(n1313), .ZN(n1123) );
XOR2_X1 U1046 ( .A(n1314), .B(n1315), .Z(n1313) );
XNOR2_X1 U1047 ( .A(G119), .B(n1316), .ZN(n1315) );
NAND2_X1 U1048 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND2_X1 U1049 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
XOR2_X1 U1050 ( .A(n1321), .B(KEYINPUT61), .Z(n1317) );
NAND2_X1 U1051 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
INV_X1 U1052 ( .A(n1320), .ZN(n1323) );
NAND3_X1 U1053 ( .A1(G234), .A2(n1105), .A3(G221), .ZN(n1320) );
INV_X1 U1054 ( .A(G953), .ZN(n1105) );
XNOR2_X1 U1055 ( .A(n1319), .B(KEYINPUT36), .ZN(n1322) );
XOR2_X1 U1056 ( .A(G137), .B(KEYINPUT15), .Z(n1319) );
NOR2_X1 U1057 ( .A1(KEYINPUT38), .A2(n1268), .ZN(n1314) );
INV_X1 U1058 ( .A(G128), .ZN(n1268) );
XOR2_X1 U1059 ( .A(n1265), .B(n1254), .Z(n1312) );
XOR2_X1 U1060 ( .A(n1324), .B(n1266), .Z(n1254) );
XNOR2_X1 U1061 ( .A(G146), .B(KEYINPUT26), .ZN(n1266) );
XNOR2_X1 U1062 ( .A(G125), .B(G140), .ZN(n1324) );
XNOR2_X1 U1063 ( .A(G110), .B(KEYINPUT31), .ZN(n1265) );
endmodule


