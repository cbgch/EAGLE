//Key = 0010100110100110000000111110110110101011011011000100010000101101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347;

XNOR2_X1 U745 ( .A(G107), .B(n1034), .ZN(G9) );
NAND4_X1 U746 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1034) );
XNOR2_X1 U747 ( .A(n1039), .B(KEYINPUT44), .ZN(n1035) );
NOR2_X1 U748 ( .A1(n1040), .A2(n1041), .ZN(G75) );
NOR4_X1 U749 ( .A1(n1042), .A2(n1043), .A3(G953), .A4(n1044), .ZN(n1041) );
NOR2_X1 U750 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U751 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U752 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U753 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U754 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR2_X1 U755 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U756 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
XOR2_X1 U758 ( .A(KEYINPUT33), .B(n1061), .Z(n1060) );
NOR2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1055) );
NOR2_X1 U761 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR4_X1 U762 ( .A1(n1068), .A2(n1058), .A3(n1069), .A4(n1070), .ZN(n1051) );
NOR3_X1 U763 ( .A1(n1065), .A2(n1068), .A3(n1058), .ZN(n1047) );
INV_X1 U764 ( .A(n1038), .ZN(n1058) );
AND3_X1 U765 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1068) );
NAND2_X1 U766 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
OR2_X1 U767 ( .A1(n1036), .A2(n1076), .ZN(n1075) );
NAND2_X1 U768 ( .A1(n1077), .A2(n1078), .ZN(n1071) );
NAND2_X1 U769 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND3_X1 U770 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1080) );
NAND2_X1 U771 ( .A1(n1039), .A2(n1070), .ZN(n1079) );
INV_X1 U772 ( .A(KEYINPUT52), .ZN(n1070) );
NOR3_X1 U773 ( .A1(n1044), .A2(G953), .A3(G952), .ZN(n1040) );
AND4_X1 U774 ( .A1(n1084), .A2(n1073), .A3(n1085), .A4(n1086), .ZN(n1044) );
NOR4_X1 U775 ( .A1(n1083), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1086) );
XNOR2_X1 U776 ( .A(n1090), .B(n1091), .ZN(n1088) );
NAND2_X1 U777 ( .A1(KEYINPUT45), .A2(n1092), .ZN(n1090) );
INV_X1 U778 ( .A(n1081), .ZN(n1087) );
INV_X1 U779 ( .A(n1093), .ZN(n1083) );
NOR2_X1 U780 ( .A1(n1094), .A2(n1095), .ZN(n1085) );
XNOR2_X1 U781 ( .A(KEYINPUT59), .B(n1096), .ZN(n1095) );
XNOR2_X1 U782 ( .A(KEYINPUT27), .B(n1082), .ZN(n1094) );
XNOR2_X1 U783 ( .A(n1097), .B(n1098), .ZN(n1084) );
NAND2_X1 U784 ( .A1(KEYINPUT32), .A2(n1099), .ZN(n1097) );
XOR2_X1 U785 ( .A(n1100), .B(n1101), .Z(G72) );
NOR2_X1 U786 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
AND2_X1 U787 ( .A1(G227), .A2(G900), .ZN(n1102) );
NAND2_X1 U788 ( .A1(n1104), .A2(n1105), .ZN(n1100) );
NAND2_X1 U789 ( .A1(n1106), .A2(n1103), .ZN(n1105) );
XNOR2_X1 U790 ( .A(n1107), .B(n1108), .ZN(n1106) );
NAND3_X1 U791 ( .A1(n1108), .A2(n1109), .A3(G953), .ZN(n1104) );
INV_X1 U792 ( .A(n1110), .ZN(n1109) );
XNOR2_X1 U793 ( .A(n1111), .B(n1112), .ZN(n1108) );
XNOR2_X1 U794 ( .A(n1113), .B(n1114), .ZN(n1112) );
NAND2_X1 U795 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NAND2_X1 U796 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U797 ( .A(KEYINPUT2), .B(n1119), .Z(n1115) );
NOR2_X1 U798 ( .A1(n1117), .A2(n1118), .ZN(n1119) );
INV_X1 U799 ( .A(G131), .ZN(n1118) );
XNOR2_X1 U800 ( .A(KEYINPUT13), .B(n1120), .ZN(n1111) );
NOR2_X1 U801 ( .A1(KEYINPUT57), .A2(n1121), .ZN(n1120) );
XOR2_X1 U802 ( .A(n1122), .B(n1123), .Z(G69) );
NOR2_X1 U803 ( .A1(n1124), .A2(n1103), .ZN(n1123) );
AND2_X1 U804 ( .A1(G224), .A2(G898), .ZN(n1124) );
NAND2_X1 U805 ( .A1(n1125), .A2(n1126), .ZN(n1122) );
NAND2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U807 ( .A1(n1129), .A2(n1103), .ZN(n1128) );
XOR2_X1 U808 ( .A(KEYINPUT53), .B(n1130), .Z(n1125) );
NOR3_X1 U809 ( .A1(n1131), .A2(G953), .A3(n1127), .ZN(n1130) );
AND2_X1 U810 ( .A1(n1132), .A2(n1133), .ZN(n1127) );
XNOR2_X1 U811 ( .A(n1134), .B(n1135), .ZN(n1133) );
XOR2_X1 U812 ( .A(n1136), .B(KEYINPUT15), .Z(n1132) );
NAND2_X1 U813 ( .A1(G953), .A2(n1137), .ZN(n1136) );
INV_X1 U814 ( .A(n1129), .ZN(n1131) );
NAND2_X1 U815 ( .A1(n1138), .A2(n1139), .ZN(n1129) );
NOR2_X1 U816 ( .A1(n1140), .A2(n1141), .ZN(G66) );
XOR2_X1 U817 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U818 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND2_X1 U819 ( .A1(KEYINPUT34), .A2(n1146), .ZN(n1142) );
XOR2_X1 U820 ( .A(KEYINPUT48), .B(n1147), .Z(n1146) );
NOR2_X1 U821 ( .A1(n1140), .A2(n1148), .ZN(G63) );
XOR2_X1 U822 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U823 ( .A1(n1151), .A2(n1145), .ZN(n1150) );
XNOR2_X1 U824 ( .A(G478), .B(KEYINPUT62), .ZN(n1151) );
NOR2_X1 U825 ( .A1(n1140), .A2(n1152), .ZN(G60) );
XOR2_X1 U826 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U827 ( .A1(n1098), .A2(n1145), .ZN(n1154) );
XNOR2_X1 U828 ( .A(G104), .B(n1155), .ZN(G6) );
NOR2_X1 U829 ( .A1(n1140), .A2(n1156), .ZN(G57) );
XOR2_X1 U830 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U831 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U832 ( .A(KEYINPUT3), .B(n1161), .Z(n1157) );
NOR2_X1 U833 ( .A1(n1162), .A2(n1145), .ZN(n1161) );
NOR2_X1 U834 ( .A1(n1140), .A2(n1163), .ZN(G54) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U836 ( .A(KEYINPUT50), .B(n1166), .Z(n1165) );
NOR3_X1 U837 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1166) );
NOR2_X1 U838 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
INV_X1 U839 ( .A(KEYINPUT18), .ZN(n1171) );
NOR3_X1 U840 ( .A1(KEYINPUT18), .A2(n1172), .A3(n1173), .ZN(n1168) );
AND2_X1 U841 ( .A1(n1173), .A2(n1172), .ZN(n1167) );
XNOR2_X1 U842 ( .A(n1174), .B(n1175), .ZN(n1172) );
NAND2_X1 U843 ( .A1(KEYINPUT39), .A2(n1170), .ZN(n1173) );
XNOR2_X1 U844 ( .A(n1176), .B(n1177), .ZN(n1164) );
NOR2_X1 U845 ( .A1(n1178), .A2(n1145), .ZN(n1177) );
NOR2_X1 U846 ( .A1(n1140), .A2(n1179), .ZN(G51) );
XOR2_X1 U847 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U848 ( .A(n1182), .B(n1183), .Z(n1181) );
NOR3_X1 U849 ( .A1(n1145), .A2(KEYINPUT40), .A3(n1184), .ZN(n1182) );
NAND2_X1 U850 ( .A1(G902), .A2(n1042), .ZN(n1145) );
NAND3_X1 U851 ( .A1(n1185), .A2(n1107), .A3(n1138), .ZN(n1042) );
AND4_X1 U852 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1138) );
NAND3_X1 U853 ( .A1(n1036), .A2(n1066), .A3(n1190), .ZN(n1186) );
AND4_X1 U854 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1107) );
AND4_X1 U855 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1194) );
NAND2_X1 U856 ( .A1(n1199), .A2(n1200), .ZN(n1193) );
NAND2_X1 U857 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NAND3_X1 U858 ( .A1(n1036), .A2(n1059), .A3(n1203), .ZN(n1202) );
NAND2_X1 U859 ( .A1(n1204), .A2(n1205), .ZN(n1201) );
XNOR2_X1 U860 ( .A(n1050), .B(KEYINPUT12), .ZN(n1205) );
INV_X1 U861 ( .A(n1077), .ZN(n1050) );
XNOR2_X1 U862 ( .A(n1139), .B(KEYINPUT29), .ZN(n1185) );
AND4_X1 U863 ( .A1(n1206), .A2(n1155), .A3(n1207), .A4(n1208), .ZN(n1139) );
NAND3_X1 U864 ( .A1(n1076), .A2(n1038), .A3(n1209), .ZN(n1155) );
NAND3_X1 U865 ( .A1(n1036), .A2(n1038), .A3(n1209), .ZN(n1206) );
XOR2_X1 U866 ( .A(n1210), .B(n1211), .Z(n1180) );
NOR2_X1 U867 ( .A1(KEYINPUT16), .A2(n1212), .ZN(n1211) );
XNOR2_X1 U868 ( .A(n1213), .B(G125), .ZN(n1210) );
NOR2_X1 U869 ( .A1(n1103), .A2(G952), .ZN(n1140) );
XNOR2_X1 U870 ( .A(G146), .B(n1191), .ZN(G48) );
NAND4_X1 U871 ( .A1(n1203), .A2(n1199), .A3(n1076), .A4(n1059), .ZN(n1191) );
XNOR2_X1 U872 ( .A(n1196), .B(n1214), .ZN(G45) );
NOR2_X1 U873 ( .A1(KEYINPUT35), .A2(n1215), .ZN(n1214) );
NAND4_X1 U874 ( .A1(n1203), .A2(n1066), .A3(n1216), .A4(n1059), .ZN(n1196) );
AND2_X1 U875 ( .A1(n1217), .A2(n1089), .ZN(n1216) );
NAND2_X1 U876 ( .A1(n1218), .A2(n1219), .ZN(G42) );
OR2_X1 U877 ( .A1(n1192), .A2(G140), .ZN(n1219) );
XOR2_X1 U878 ( .A(n1220), .B(KEYINPUT30), .Z(n1218) );
NAND2_X1 U879 ( .A1(G140), .A2(n1192), .ZN(n1220) );
NAND3_X1 U880 ( .A1(n1204), .A2(n1076), .A3(n1067), .ZN(n1192) );
XOR2_X1 U881 ( .A(n1221), .B(n1222), .Z(G39) );
NAND2_X1 U882 ( .A1(n1204), .A2(n1223), .ZN(n1222) );
NAND2_X1 U883 ( .A1(n1224), .A2(KEYINPUT25), .ZN(n1221) );
XNOR2_X1 U884 ( .A(G137), .B(KEYINPUT8), .ZN(n1224) );
XOR2_X1 U885 ( .A(n1195), .B(n1225), .Z(G36) );
XOR2_X1 U886 ( .A(KEYINPUT24), .B(G134), .Z(n1225) );
NAND3_X1 U887 ( .A1(n1036), .A2(n1066), .A3(n1204), .ZN(n1195) );
NAND2_X1 U888 ( .A1(n1226), .A2(n1227), .ZN(G33) );
OR2_X1 U889 ( .A1(n1198), .A2(G131), .ZN(n1227) );
XOR2_X1 U890 ( .A(n1228), .B(KEYINPUT21), .Z(n1226) );
NAND2_X1 U891 ( .A1(G131), .A2(n1198), .ZN(n1228) );
NAND3_X1 U892 ( .A1(n1076), .A2(n1066), .A3(n1204), .ZN(n1198) );
AND2_X1 U893 ( .A1(n1203), .A2(n1073), .ZN(n1204) );
INV_X1 U894 ( .A(n1065), .ZN(n1073) );
NAND2_X1 U895 ( .A1(n1229), .A2(n1063), .ZN(n1065) );
INV_X1 U896 ( .A(n1062), .ZN(n1229) );
XOR2_X1 U897 ( .A(n1230), .B(n1231), .Z(G30) );
NOR2_X1 U898 ( .A1(KEYINPUT46), .A2(n1232), .ZN(n1231) );
NOR2_X1 U899 ( .A1(n1233), .A2(n1234), .ZN(n1230) );
XOR2_X1 U900 ( .A(n1235), .B(KEYINPUT43), .Z(n1233) );
NAND3_X1 U901 ( .A1(n1199), .A2(n1036), .A3(n1203), .ZN(n1235) );
AND2_X1 U902 ( .A1(n1039), .A2(n1236), .ZN(n1203) );
XNOR2_X1 U903 ( .A(G101), .B(n1207), .ZN(G3) );
NAND3_X1 U904 ( .A1(n1066), .A2(n1077), .A3(n1209), .ZN(n1207) );
XNOR2_X1 U905 ( .A(G125), .B(n1197), .ZN(G27) );
NAND4_X1 U906 ( .A1(n1059), .A2(n1236), .A3(n1074), .A4(n1237), .ZN(n1197) );
NOR2_X1 U907 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND2_X1 U908 ( .A1(n1240), .A2(n1046), .ZN(n1236) );
NAND4_X1 U909 ( .A1(G953), .A2(G902), .A3(n1110), .A4(n1241), .ZN(n1240) );
XOR2_X1 U910 ( .A(G900), .B(KEYINPUT26), .Z(n1110) );
XNOR2_X1 U911 ( .A(G122), .B(n1187), .ZN(G24) );
NAND4_X1 U912 ( .A1(n1190), .A2(n1038), .A3(n1089), .A4(n1217), .ZN(n1187) );
NAND2_X1 U913 ( .A1(n1242), .A2(n1243), .ZN(n1038) );
NAND2_X1 U914 ( .A1(n1066), .A2(n1244), .ZN(n1243) );
OR3_X1 U915 ( .A1(n1245), .A2(n1246), .A3(n1244), .ZN(n1242) );
XNOR2_X1 U916 ( .A(G119), .B(n1188), .ZN(G21) );
NAND2_X1 U917 ( .A1(n1223), .A2(n1190), .ZN(n1188) );
AND2_X1 U918 ( .A1(n1199), .A2(n1077), .ZN(n1223) );
AND2_X1 U919 ( .A1(n1246), .A2(n1245), .ZN(n1199) );
XNOR2_X1 U920 ( .A(G116), .B(n1247), .ZN(G18) );
NAND4_X1 U921 ( .A1(n1248), .A2(n1036), .A3(n1037), .A4(n1066), .ZN(n1247) );
XNOR2_X1 U922 ( .A(n1074), .B(KEYINPUT63), .ZN(n1248) );
NAND2_X1 U923 ( .A1(n1249), .A2(n1250), .ZN(G15) );
OR2_X1 U924 ( .A1(n1189), .A2(n1251), .ZN(n1250) );
XOR2_X1 U925 ( .A(n1252), .B(KEYINPUT51), .Z(n1249) );
NAND2_X1 U926 ( .A1(n1251), .A2(n1189), .ZN(n1252) );
NAND3_X1 U927 ( .A1(n1190), .A2(n1066), .A3(n1076), .ZN(n1189) );
INV_X1 U928 ( .A(n1238), .ZN(n1076) );
NAND2_X1 U929 ( .A1(n1253), .A2(n1217), .ZN(n1238) );
XNOR2_X1 U930 ( .A(KEYINPUT37), .B(n1089), .ZN(n1253) );
NOR2_X1 U931 ( .A1(n1246), .A2(n1096), .ZN(n1066) );
INV_X1 U932 ( .A(n1245), .ZN(n1096) );
AND2_X1 U933 ( .A1(n1074), .A2(n1037), .ZN(n1190) );
INV_X1 U934 ( .A(n1054), .ZN(n1074) );
NAND3_X1 U935 ( .A1(n1082), .A2(n1093), .A3(n1081), .ZN(n1054) );
XOR2_X1 U936 ( .A(G113), .B(KEYINPUT55), .Z(n1251) );
XNOR2_X1 U937 ( .A(G110), .B(n1208), .ZN(G12) );
NAND3_X1 U938 ( .A1(n1067), .A2(n1077), .A3(n1209), .ZN(n1208) );
AND2_X1 U939 ( .A1(n1037), .A2(n1039), .ZN(n1209) );
INV_X1 U940 ( .A(n1069), .ZN(n1039) );
NAND2_X1 U941 ( .A1(n1093), .A2(n1254), .ZN(n1069) );
NAND2_X1 U942 ( .A1(n1081), .A2(n1082), .ZN(n1254) );
NAND2_X1 U943 ( .A1(G469), .A2(n1255), .ZN(n1082) );
NAND2_X1 U944 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND3_X1 U945 ( .A1(n1178), .A2(n1257), .A3(n1256), .ZN(n1081) );
XOR2_X1 U946 ( .A(n1258), .B(n1259), .Z(n1256) );
XNOR2_X1 U947 ( .A(n1260), .B(n1176), .ZN(n1259) );
XNOR2_X1 U948 ( .A(n1261), .B(n1159), .ZN(n1176) );
XNOR2_X1 U949 ( .A(n1262), .B(n1263), .ZN(n1261) );
INV_X1 U950 ( .A(n1114), .ZN(n1263) );
XOR2_X1 U951 ( .A(n1264), .B(n1232), .Z(n1114) );
NAND2_X1 U952 ( .A1(KEYINPUT58), .A2(n1265), .ZN(n1264) );
XOR2_X1 U953 ( .A(KEYINPUT61), .B(n1266), .Z(n1265) );
NAND2_X1 U954 ( .A1(n1267), .A2(n1268), .ZN(n1262) );
NAND2_X1 U955 ( .A1(KEYINPUT60), .A2(n1174), .ZN(n1260) );
XNOR2_X1 U956 ( .A(G140), .B(n1170), .ZN(n1258) );
AND2_X1 U957 ( .A1(G227), .A2(n1103), .ZN(n1170) );
INV_X1 U958 ( .A(G469), .ZN(n1178) );
NAND2_X1 U959 ( .A1(G221), .A2(n1269), .ZN(n1093) );
AND2_X1 U960 ( .A1(n1059), .A2(n1270), .ZN(n1037) );
NAND2_X1 U961 ( .A1(n1046), .A2(n1271), .ZN(n1270) );
NAND4_X1 U962 ( .A1(G953), .A2(G902), .A3(n1241), .A4(n1137), .ZN(n1271) );
INV_X1 U963 ( .A(G898), .ZN(n1137) );
NAND3_X1 U964 ( .A1(n1241), .A2(n1103), .A3(G952), .ZN(n1046) );
NAND2_X1 U965 ( .A1(G237), .A2(G234), .ZN(n1241) );
INV_X1 U966 ( .A(n1234), .ZN(n1059) );
NAND2_X1 U967 ( .A1(n1062), .A2(n1063), .ZN(n1234) );
NAND2_X1 U968 ( .A1(G214), .A2(n1272), .ZN(n1063) );
XOR2_X1 U969 ( .A(n1273), .B(n1184), .Z(n1062) );
NAND2_X1 U970 ( .A1(G210), .A2(n1272), .ZN(n1184) );
NAND2_X1 U971 ( .A1(n1257), .A2(n1274), .ZN(n1272) );
NAND2_X1 U972 ( .A1(n1275), .A2(n1257), .ZN(n1273) );
XOR2_X1 U973 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U974 ( .A(n1183), .B(n1278), .ZN(n1277) );
NOR2_X1 U975 ( .A1(n1213), .A2(KEYINPUT9), .ZN(n1278) );
XNOR2_X1 U976 ( .A(n1134), .B(n1279), .ZN(n1183) );
NOR2_X1 U977 ( .A1(KEYINPUT1), .A2(n1135), .ZN(n1279) );
XOR2_X1 U978 ( .A(n1280), .B(n1281), .Z(n1135) );
NAND2_X1 U979 ( .A1(KEYINPUT22), .A2(n1282), .ZN(n1280) );
XOR2_X1 U980 ( .A(n1283), .B(n1284), .Z(n1134) );
XNOR2_X1 U981 ( .A(n1285), .B(n1174), .ZN(n1283) );
NAND3_X1 U982 ( .A1(n1286), .A2(n1287), .A3(n1268), .ZN(n1285) );
OR3_X1 U983 ( .A1(n1288), .A2(G107), .A3(n1289), .ZN(n1268) );
NAND2_X1 U984 ( .A1(KEYINPUT19), .A2(n1290), .ZN(n1287) );
XOR2_X1 U985 ( .A(n1291), .B(n1289), .Z(n1290) );
NAND2_X1 U986 ( .A1(G107), .A2(n1288), .ZN(n1291) );
OR2_X1 U987 ( .A1(n1267), .A2(KEYINPUT19), .ZN(n1286) );
AND2_X1 U988 ( .A1(n1292), .A2(n1293), .ZN(n1267) );
NAND2_X1 U989 ( .A1(n1294), .A2(G107), .ZN(n1293) );
XNOR2_X1 U990 ( .A(G104), .B(n1289), .ZN(n1294) );
NAND3_X1 U991 ( .A1(n1289), .A2(n1288), .A3(n1295), .ZN(n1292) );
INV_X1 U992 ( .A(G107), .ZN(n1295) );
XOR2_X1 U993 ( .A(n1296), .B(KEYINPUT5), .Z(n1289) );
XOR2_X1 U994 ( .A(n1212), .B(n1297), .Z(n1276) );
XOR2_X1 U995 ( .A(KEYINPUT41), .B(G125), .Z(n1297) );
NAND2_X1 U996 ( .A1(G224), .A2(n1103), .ZN(n1212) );
NAND2_X1 U997 ( .A1(n1298), .A2(n1299), .ZN(n1077) );
OR3_X1 U998 ( .A1(n1217), .A2(n1089), .A3(KEYINPUT37), .ZN(n1299) );
NAND2_X1 U999 ( .A1(KEYINPUT37), .A2(n1036), .ZN(n1298) );
NOR2_X1 U1000 ( .A1(n1217), .A2(n1300), .ZN(n1036) );
INV_X1 U1001 ( .A(n1089), .ZN(n1300) );
XOR2_X1 U1002 ( .A(G478), .B(n1301), .Z(n1089) );
NOR2_X1 U1003 ( .A1(n1149), .A2(G902), .ZN(n1301) );
AND2_X1 U1004 ( .A1(n1302), .A2(n1303), .ZN(n1149) );
NAND2_X1 U1005 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
XOR2_X1 U1006 ( .A(KEYINPUT10), .B(n1306), .Z(n1302) );
NOR2_X1 U1007 ( .A1(n1304), .A2(n1305), .ZN(n1306) );
XNOR2_X1 U1008 ( .A(n1307), .B(n1308), .ZN(n1305) );
XOR2_X1 U1009 ( .A(n1309), .B(n1310), .Z(n1308) );
XNOR2_X1 U1010 ( .A(G134), .B(KEYINPUT6), .ZN(n1310) );
NAND2_X1 U1011 ( .A1(KEYINPUT14), .A2(n1311), .ZN(n1309) );
XNOR2_X1 U1012 ( .A(n1215), .B(G128), .ZN(n1311) );
INV_X1 U1013 ( .A(G143), .ZN(n1215) );
XNOR2_X1 U1014 ( .A(n1284), .B(n1312), .ZN(n1307) );
XOR2_X1 U1015 ( .A(n1313), .B(n1314), .Z(n1312) );
NOR2_X1 U1016 ( .A1(G107), .A2(KEYINPUT11), .ZN(n1313) );
AND3_X1 U1017 ( .A1(G217), .A2(n1103), .A3(G234), .ZN(n1304) );
XNOR2_X1 U1018 ( .A(n1099), .B(n1098), .ZN(n1217) );
INV_X1 U1019 ( .A(G475), .ZN(n1098) );
NOR2_X1 U1020 ( .A1(n1153), .A2(G902), .ZN(n1099) );
XOR2_X1 U1021 ( .A(n1315), .B(n1316), .Z(n1153) );
XNOR2_X1 U1022 ( .A(n1266), .B(n1317), .ZN(n1316) );
XOR2_X1 U1023 ( .A(n1318), .B(n1319), .Z(n1317) );
AND3_X1 U1024 ( .A1(G214), .A2(n1103), .A3(n1274), .ZN(n1319) );
NAND2_X1 U1025 ( .A1(n1320), .A2(KEYINPUT31), .ZN(n1318) );
XOR2_X1 U1026 ( .A(n1321), .B(G125), .Z(n1320) );
NAND2_X1 U1027 ( .A1(KEYINPUT36), .A2(n1175), .ZN(n1321) );
XOR2_X1 U1028 ( .A(n1322), .B(n1323), .Z(n1315) );
XNOR2_X1 U1029 ( .A(n1288), .B(n1324), .ZN(n1323) );
NOR2_X1 U1030 ( .A1(KEYINPUT0), .A2(n1284), .ZN(n1324) );
XOR2_X1 U1031 ( .A(G122), .B(KEYINPUT23), .Z(n1284) );
INV_X1 U1032 ( .A(G104), .ZN(n1288) );
XNOR2_X1 U1033 ( .A(G113), .B(G131), .ZN(n1322) );
INV_X1 U1034 ( .A(n1239), .ZN(n1067) );
NAND2_X1 U1035 ( .A1(n1325), .A2(n1246), .ZN(n1239) );
XOR2_X1 U1036 ( .A(n1091), .B(n1092), .Z(n1246) );
NAND2_X1 U1037 ( .A1(n1326), .A2(n1269), .ZN(n1092) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1257), .ZN(n1269) );
XNOR2_X1 U1039 ( .A(KEYINPUT47), .B(n1144), .ZN(n1326) );
INV_X1 U1040 ( .A(G217), .ZN(n1144) );
NAND2_X1 U1041 ( .A1(n1147), .A2(n1257), .ZN(n1091) );
INV_X1 U1042 ( .A(G902), .ZN(n1257) );
XNOR2_X1 U1043 ( .A(n1327), .B(n1328), .ZN(n1147) );
XOR2_X1 U1044 ( .A(n1329), .B(n1330), .Z(n1328) );
XNOR2_X1 U1045 ( .A(G137), .B(n1174), .ZN(n1330) );
INV_X1 U1046 ( .A(G110), .ZN(n1174) );
XOR2_X1 U1047 ( .A(KEYINPUT56), .B(G146), .Z(n1329) );
XNOR2_X1 U1048 ( .A(n1121), .B(n1331), .ZN(n1327) );
XOR2_X1 U1049 ( .A(n1332), .B(n1333), .Z(n1331) );
AND3_X1 U1050 ( .A1(G221), .A2(n1103), .A3(G234), .ZN(n1333) );
NOR2_X1 U1051 ( .A1(KEYINPUT17), .A2(n1334), .ZN(n1332) );
XNOR2_X1 U1052 ( .A(n1232), .B(n1335), .ZN(n1334) );
NOR2_X1 U1053 ( .A1(G119), .A2(KEYINPUT54), .ZN(n1335) );
INV_X1 U1054 ( .A(G128), .ZN(n1232) );
XNOR2_X1 U1055 ( .A(G125), .B(n1175), .ZN(n1121) );
INV_X1 U1056 ( .A(G140), .ZN(n1175) );
XNOR2_X1 U1057 ( .A(n1244), .B(n1245), .ZN(n1325) );
XOR2_X1 U1058 ( .A(n1336), .B(n1162), .Z(n1245) );
INV_X1 U1059 ( .A(G472), .ZN(n1162) );
NAND2_X1 U1060 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
XOR2_X1 U1061 ( .A(n1339), .B(n1160), .Z(n1338) );
XNOR2_X1 U1062 ( .A(n1340), .B(n1341), .ZN(n1160) );
XNOR2_X1 U1063 ( .A(n1296), .B(n1282), .ZN(n1341) );
XNOR2_X1 U1064 ( .A(G119), .B(n1314), .ZN(n1282) );
XOR2_X1 U1065 ( .A(G116), .B(KEYINPUT7), .Z(n1314) );
XOR2_X1 U1066 ( .A(G101), .B(KEYINPUT38), .Z(n1296) );
XNOR2_X1 U1067 ( .A(n1213), .B(n1342), .ZN(n1340) );
XNOR2_X1 U1068 ( .A(n1281), .B(n1343), .ZN(n1342) );
AND3_X1 U1069 ( .A1(G210), .A2(n1103), .A3(n1274), .ZN(n1343) );
INV_X1 U1070 ( .A(G237), .ZN(n1274) );
INV_X1 U1071 ( .A(G953), .ZN(n1103) );
INV_X1 U1072 ( .A(G113), .ZN(n1281) );
AND2_X1 U1073 ( .A1(n1344), .A2(n1345), .ZN(n1213) );
NAND2_X1 U1074 ( .A1(G128), .A2(n1266), .ZN(n1345) );
XOR2_X1 U1075 ( .A(KEYINPUT28), .B(n1346), .Z(n1344) );
NOR2_X1 U1076 ( .A1(G128), .A2(n1266), .ZN(n1346) );
XOR2_X1 U1077 ( .A(G143), .B(G146), .Z(n1266) );
NAND2_X1 U1078 ( .A1(KEYINPUT4), .A2(n1159), .ZN(n1339) );
XOR2_X1 U1079 ( .A(n1347), .B(n1117), .Z(n1159) );
XNOR2_X1 U1080 ( .A(G134), .B(G137), .ZN(n1117) );
XNOR2_X1 U1081 ( .A(G131), .B(KEYINPUT49), .ZN(n1347) );
XNOR2_X1 U1082 ( .A(G902), .B(KEYINPUT20), .ZN(n1337) );
INV_X1 U1083 ( .A(KEYINPUT42), .ZN(n1244) );
endmodule


