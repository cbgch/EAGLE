//Key = 1000000000000111001101000101011110100011010001101000011101011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273;

XNOR2_X1 U703 ( .A(G107), .B(n973), .ZN(G9) );
NAND4_X1 U704 ( .A1(n974), .A2(n975), .A3(n976), .A4(n977), .ZN(n973) );
NOR2_X1 U705 ( .A1(n978), .A2(n979), .ZN(n976) );
XOR2_X1 U706 ( .A(n980), .B(KEYINPUT37), .Z(n978) );
XOR2_X1 U707 ( .A(n981), .B(KEYINPUT12), .Z(n974) );
NOR2_X1 U708 ( .A1(n982), .A2(n983), .ZN(G75) );
XOR2_X1 U709 ( .A(n984), .B(KEYINPUT0), .Z(n983) );
NAND3_X1 U710 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n984) );
NOR3_X1 U711 ( .A1(n988), .A2(n985), .A3(n989), .ZN(n982) );
INV_X1 U712 ( .A(G952), .ZN(n985) );
NAND3_X1 U713 ( .A1(n987), .A2(n986), .A3(n990), .ZN(n988) );
NAND2_X1 U714 ( .A1(n991), .A2(n992), .ZN(n990) );
NAND2_X1 U715 ( .A1(n993), .A2(n994), .ZN(n992) );
NAND3_X1 U716 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n994) );
NAND2_X1 U717 ( .A1(n998), .A2(n999), .ZN(n996) );
NAND2_X1 U718 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NAND2_X1 U719 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NAND2_X1 U720 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
INV_X1 U721 ( .A(n975), .ZN(n1002) );
NAND2_X1 U722 ( .A1(n1006), .A2(n1007), .ZN(n998) );
NAND3_X1 U723 ( .A1(n1000), .A2(n1008), .A3(n1006), .ZN(n993) );
NAND2_X1 U724 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND2_X1 U725 ( .A1(n997), .A2(n1011), .ZN(n1010) );
XOR2_X1 U726 ( .A(n1012), .B(n1013), .Z(n1011) );
NAND2_X1 U727 ( .A1(n995), .A2(n1014), .ZN(n1009) );
NAND2_X1 U728 ( .A1(n980), .A2(n1015), .ZN(n1014) );
NAND2_X1 U729 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
INV_X1 U730 ( .A(n1018), .ZN(n1016) );
INV_X1 U731 ( .A(n1019), .ZN(n991) );
NAND4_X1 U732 ( .A1(n1020), .A2(n1018), .A3(n1021), .A4(n1022), .ZN(n987) );
NOR3_X1 U733 ( .A1(n1023), .A2(n979), .A3(n1024), .ZN(n1022) );
XOR2_X1 U734 ( .A(n1025), .B(n1026), .Z(n1021) );
XOR2_X1 U735 ( .A(G475), .B(n1027), .Z(n1026) );
NOR2_X1 U736 ( .A1(n1028), .A2(KEYINPUT42), .ZN(n1027) );
XOR2_X1 U737 ( .A(KEYINPUT55), .B(KEYINPUT41), .Z(n1025) );
XOR2_X1 U738 ( .A(n1029), .B(n1030), .Z(n1020) );
XOR2_X1 U739 ( .A(n1031), .B(KEYINPUT57), .Z(n1030) );
XOR2_X1 U740 ( .A(n1032), .B(n1033), .Z(G72) );
XOR2_X1 U741 ( .A(n1034), .B(n1035), .Z(n1033) );
NOR2_X1 U742 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
XOR2_X1 U743 ( .A(n1038), .B(n1039), .Z(n1037) );
NOR2_X1 U744 ( .A1(KEYINPUT20), .A2(n1040), .ZN(n1039) );
NOR2_X1 U745 ( .A1(n1041), .A2(n1042), .ZN(n1038) );
XOR2_X1 U746 ( .A(KEYINPUT49), .B(n1043), .Z(n1042) );
AND2_X1 U747 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U748 ( .A1(n1044), .A2(n1045), .ZN(n1041) );
XOR2_X1 U749 ( .A(G131), .B(n1046), .Z(n1045) );
INV_X1 U750 ( .A(n1047), .ZN(n1044) );
NOR2_X1 U751 ( .A1(G900), .A2(n986), .ZN(n1036) );
NAND2_X1 U752 ( .A1(n1048), .A2(n1049), .ZN(n1034) );
NAND3_X1 U753 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
XNOR2_X1 U754 ( .A(n1053), .B(KEYINPUT39), .ZN(n1052) );
XOR2_X1 U755 ( .A(KEYINPUT14), .B(G953), .Z(n1048) );
NAND2_X1 U756 ( .A1(G953), .A2(n1054), .ZN(n1032) );
NAND2_X1 U757 ( .A1(G900), .A2(G227), .ZN(n1054) );
XOR2_X1 U758 ( .A(n1055), .B(n1056), .Z(G69) );
XOR2_X1 U759 ( .A(n1057), .B(n1058), .Z(n1056) );
NOR2_X1 U760 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XOR2_X1 U761 ( .A(KEYINPUT4), .B(n1061), .Z(n1060) );
NOR2_X1 U762 ( .A1(G898), .A2(n986), .ZN(n1061) );
INV_X1 U763 ( .A(n1062), .ZN(n1059) );
NOR2_X1 U764 ( .A1(KEYINPUT22), .A2(n1063), .ZN(n1057) );
NOR2_X1 U765 ( .A1(n1064), .A2(n986), .ZN(n1063) );
NOR2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U767 ( .A1(n986), .A2(n1067), .ZN(n1055) );
NAND4_X1 U768 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1067) );
NOR2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(G66) );
XOR2_X1 U770 ( .A(n1074), .B(n1075), .Z(n1073) );
NOR2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U772 ( .A1(n1072), .A2(n1078), .ZN(G63) );
XOR2_X1 U773 ( .A(n1079), .B(n1080), .Z(n1078) );
XOR2_X1 U774 ( .A(n1081), .B(KEYINPUT16), .Z(n1079) );
NAND2_X1 U775 ( .A1(n1082), .A2(G478), .ZN(n1081) );
NOR2_X1 U776 ( .A1(n1072), .A2(n1083), .ZN(G60) );
NOR3_X1 U777 ( .A1(n1028), .A2(n1084), .A3(n1085), .ZN(n1083) );
AND3_X1 U778 ( .A1(n1086), .A2(G475), .A3(n1082), .ZN(n1085) );
NOR2_X1 U779 ( .A1(n1087), .A2(n1086), .ZN(n1084) );
AND2_X1 U780 ( .A1(n989), .A2(G475), .ZN(n1087) );
XOR2_X1 U781 ( .A(G104), .B(n1088), .Z(G6) );
NOR4_X1 U782 ( .A1(KEYINPUT28), .A2(n979), .A3(n1089), .A4(n1090), .ZN(n1088) );
NOR2_X1 U783 ( .A1(n1091), .A2(n1092), .ZN(G57) );
XOR2_X1 U784 ( .A(KEYINPUT56), .B(n1072), .Z(n1092) );
XOR2_X1 U785 ( .A(n1093), .B(n1094), .Z(n1091) );
XOR2_X1 U786 ( .A(n1095), .B(n1096), .Z(n1094) );
XOR2_X1 U787 ( .A(n1097), .B(n1098), .Z(n1093) );
XOR2_X1 U788 ( .A(n1099), .B(n1100), .Z(n1098) );
NAND2_X1 U789 ( .A1(n1082), .A2(G472), .ZN(n1100) );
NAND2_X1 U790 ( .A1(KEYINPUT62), .A2(n1047), .ZN(n1097) );
NOR3_X1 U791 ( .A1(n1072), .A2(n1101), .A3(n1102), .ZN(G54) );
NOR2_X1 U792 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U793 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NOR2_X1 U794 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U795 ( .A1(n1109), .A2(n1110), .ZN(n1105) );
NOR2_X1 U796 ( .A1(n1111), .A2(n1112), .ZN(n1101) );
NOR2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U798 ( .A1(n1109), .A2(n1108), .ZN(n1114) );
XOR2_X1 U799 ( .A(n1115), .B(n1110), .Z(n1108) );
XNOR2_X1 U800 ( .A(KEYINPUT35), .B(KEYINPUT33), .ZN(n1115) );
NOR2_X1 U801 ( .A1(n1107), .A2(n1110), .ZN(n1113) );
XOR2_X1 U802 ( .A(n1116), .B(n1117), .Z(n1110) );
AND2_X1 U803 ( .A1(G469), .A2(n1082), .ZN(n1117) );
INV_X1 U804 ( .A(n1077), .ZN(n1082) );
NAND2_X1 U805 ( .A1(G902), .A2(n989), .ZN(n1077) );
XOR2_X1 U806 ( .A(n1118), .B(n1119), .Z(n1116) );
NOR2_X1 U807 ( .A1(KEYINPUT52), .A2(n1120), .ZN(n1119) );
INV_X1 U808 ( .A(n1109), .ZN(n1107) );
INV_X1 U809 ( .A(n1104), .ZN(n1111) );
NOR2_X1 U810 ( .A1(n1072), .A2(n1121), .ZN(G51) );
XOR2_X1 U811 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U812 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND2_X1 U813 ( .A1(KEYINPUT31), .A2(n1062), .ZN(n1125) );
NAND3_X1 U814 ( .A1(G902), .A2(n1126), .A3(n1127), .ZN(n1124) );
XOR2_X1 U815 ( .A(n989), .B(KEYINPUT47), .Z(n1127) );
NAND4_X1 U816 ( .A1(n1053), .A2(n1128), .A3(n1050), .A4(n1129), .ZN(n989) );
AND4_X1 U817 ( .A1(n1071), .A2(n1070), .A3(n1051), .A4(n1069), .ZN(n1129) );
NAND3_X1 U818 ( .A1(n995), .A2(n1007), .A3(n1130), .ZN(n1069) );
OR2_X1 U819 ( .A1(n1131), .A2(n977), .ZN(n1007) );
INV_X1 U820 ( .A(n979), .ZN(n995) );
NAND2_X1 U821 ( .A1(n1132), .A2(n997), .ZN(n1051) );
XOR2_X1 U822 ( .A(n1133), .B(KEYINPUT15), .Z(n1132) );
AND3_X1 U823 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1050) );
XOR2_X1 U824 ( .A(KEYINPUT10), .B(n1068), .Z(n1128) );
AND4_X1 U825 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1068) );
AND4_X1 U826 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1053) );
NOR2_X1 U827 ( .A1(n1145), .A2(n1146), .ZN(n1141) );
NOR3_X1 U828 ( .A1(n1147), .A2(n1148), .A3(n980), .ZN(n1146) );
INV_X1 U829 ( .A(KEYINPUT58), .ZN(n1147) );
NOR2_X1 U830 ( .A1(KEYINPUT58), .A2(n1149), .ZN(n1145) );
NOR2_X1 U831 ( .A1(n986), .A2(G952), .ZN(n1072) );
XNOR2_X1 U832 ( .A(n1136), .B(n1150), .ZN(G48) );
NOR2_X1 U833 ( .A1(KEYINPUT44), .A2(n1151), .ZN(n1150) );
NAND3_X1 U834 ( .A1(n1152), .A2(n1153), .A3(n1131), .ZN(n1136) );
XNOR2_X1 U835 ( .A(G143), .B(n1134), .ZN(G45) );
NAND4_X1 U836 ( .A1(n1154), .A2(n1153), .A3(n1024), .A4(n1155), .ZN(n1134) );
XOR2_X1 U837 ( .A(n1156), .B(G140), .Z(G42) );
NAND2_X1 U838 ( .A1(KEYINPUT25), .A2(n1135), .ZN(n1156) );
NAND3_X1 U839 ( .A1(n997), .A2(n975), .A3(n1157), .ZN(n1135) );
XOR2_X1 U840 ( .A(n1158), .B(n1159), .Z(G39) );
NOR2_X1 U841 ( .A1(n1160), .A2(KEYINPUT50), .ZN(n1159) );
NOR2_X1 U842 ( .A1(n1133), .A2(n1161), .ZN(n1160) );
NAND2_X1 U843 ( .A1(n1152), .A2(n1000), .ZN(n1133) );
XNOR2_X1 U844 ( .A(G134), .B(n1142), .ZN(G36) );
NAND3_X1 U845 ( .A1(n997), .A2(n977), .A3(n1154), .ZN(n1142) );
XNOR2_X1 U846 ( .A(G131), .B(n1143), .ZN(G33) );
NAND3_X1 U847 ( .A1(n1131), .A2(n997), .A3(n1154), .ZN(n1143) );
AND2_X1 U848 ( .A1(n1162), .A2(n1163), .ZN(n1154) );
INV_X1 U849 ( .A(n1161), .ZN(n997) );
NAND2_X1 U850 ( .A1(n1017), .A2(n1018), .ZN(n1161) );
XNOR2_X1 U851 ( .A(G128), .B(n1164), .ZN(G30) );
NOR2_X1 U852 ( .A1(n1165), .A2(KEYINPUT51), .ZN(n1164) );
INV_X1 U853 ( .A(n1149), .ZN(n1165) );
NAND2_X1 U854 ( .A1(n1148), .A2(n1153), .ZN(n1149) );
AND2_X1 U855 ( .A1(n1152), .A2(n977), .ZN(n1148) );
AND2_X1 U856 ( .A1(n1162), .A2(n1013), .ZN(n1152) );
AND3_X1 U857 ( .A1(n1012), .A2(n1166), .A3(n975), .ZN(n1162) );
XOR2_X1 U858 ( .A(n1167), .B(n1070), .Z(G3) );
NAND4_X1 U859 ( .A1(n1000), .A2(n1130), .A3(n1163), .A4(n1012), .ZN(n1070) );
XNOR2_X1 U860 ( .A(n1168), .B(n1144), .ZN(G27) );
NAND3_X1 U861 ( .A1(n1157), .A2(n1153), .A3(n1006), .ZN(n1144) );
AND4_X1 U862 ( .A1(n1169), .A2(n1131), .A3(n1013), .A4(n1166), .ZN(n1157) );
NAND2_X1 U863 ( .A1(n1170), .A2(n1019), .ZN(n1166) );
NAND2_X1 U864 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
INV_X1 U865 ( .A(G900), .ZN(n1172) );
XNOR2_X1 U866 ( .A(G125), .B(KEYINPUT48), .ZN(n1168) );
XOR2_X1 U867 ( .A(n1173), .B(G122), .Z(G24) );
NAND2_X1 U868 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NAND3_X1 U869 ( .A1(n1176), .A2(n980), .A3(n1177), .ZN(n1175) );
OR2_X1 U870 ( .A1(n1138), .A2(n1177), .ZN(n1174) );
INV_X1 U871 ( .A(KEYINPUT27), .ZN(n1177) );
NAND2_X1 U872 ( .A1(n1176), .A2(n1153), .ZN(n1138) );
AND4_X1 U873 ( .A1(n1155), .A2(n981), .A3(n1024), .A4(n1178), .ZN(n1176) );
NOR2_X1 U874 ( .A1(n979), .A2(n1023), .ZN(n1178) );
NAND2_X1 U875 ( .A1(n1163), .A2(n1169), .ZN(n979) );
XOR2_X1 U876 ( .A(n1179), .B(n1180), .Z(G21) );
XOR2_X1 U877 ( .A(KEYINPUT38), .B(G119), .Z(n1180) );
NAND2_X1 U878 ( .A1(KEYINPUT13), .A2(n1181), .ZN(n1179) );
INV_X1 U879 ( .A(n1137), .ZN(n1181) );
NAND3_X1 U880 ( .A1(n1000), .A2(n1013), .A3(n1182), .ZN(n1137) );
NAND2_X1 U881 ( .A1(n1183), .A2(n1184), .ZN(G18) );
NAND2_X1 U882 ( .A1(G116), .A2(n1139), .ZN(n1184) );
XOR2_X1 U883 ( .A(KEYINPUT21), .B(n1185), .Z(n1183) );
NOR2_X1 U884 ( .A1(G116), .A2(n1139), .ZN(n1185) );
NAND3_X1 U885 ( .A1(n1163), .A2(n977), .A3(n1182), .ZN(n1139) );
NOR2_X1 U886 ( .A1(n1155), .A2(n1186), .ZN(n977) );
XNOR2_X1 U887 ( .A(G113), .B(n1140), .ZN(G15) );
NAND3_X1 U888 ( .A1(n1163), .A2(n1131), .A3(n1182), .ZN(n1140) );
AND4_X1 U889 ( .A1(n1006), .A2(n1153), .A3(n1012), .A4(n981), .ZN(n1182) );
INV_X1 U890 ( .A(n1169), .ZN(n1012) );
INV_X1 U891 ( .A(n1023), .ZN(n1006) );
NAND2_X1 U892 ( .A1(n1005), .A2(n1187), .ZN(n1023) );
INV_X1 U893 ( .A(n1090), .ZN(n1131) );
NAND2_X1 U894 ( .A1(n1186), .A2(n1155), .ZN(n1090) );
XNOR2_X1 U895 ( .A(n1071), .B(n1188), .ZN(G12) );
NOR2_X1 U896 ( .A1(KEYINPUT63), .A2(n1189), .ZN(n1188) );
NAND4_X1 U897 ( .A1(n1000), .A2(n1130), .A3(n1169), .A4(n1013), .ZN(n1071) );
INV_X1 U898 ( .A(n1163), .ZN(n1013) );
XNOR2_X1 U899 ( .A(n1190), .B(n1076), .ZN(n1163) );
NAND2_X1 U900 ( .A1(G217), .A2(n1191), .ZN(n1076) );
OR2_X1 U901 ( .A1(n1075), .A2(G902), .ZN(n1190) );
XNOR2_X1 U902 ( .A(n1192), .B(n1193), .ZN(n1075) );
NOR2_X1 U903 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
XOR2_X1 U904 ( .A(n1196), .B(KEYINPUT54), .Z(n1195) );
NAND2_X1 U905 ( .A1(n1197), .A2(G110), .ZN(n1196) );
NOR2_X1 U906 ( .A1(G110), .A2(n1197), .ZN(n1194) );
XOR2_X1 U907 ( .A(n1198), .B(n1199), .Z(n1197) );
XOR2_X1 U908 ( .A(KEYINPUT18), .B(G128), .Z(n1199) );
INV_X1 U909 ( .A(G119), .ZN(n1198) );
XNOR2_X1 U910 ( .A(n1200), .B(n1201), .ZN(n1192) );
NOR2_X1 U911 ( .A1(KEYINPUT2), .A2(n1202), .ZN(n1201) );
XOR2_X1 U912 ( .A(n1203), .B(n1040), .Z(n1202) );
NOR2_X1 U913 ( .A1(KEYINPUT43), .A2(n1204), .ZN(n1200) );
XOR2_X1 U914 ( .A(n1205), .B(G137), .Z(n1204) );
NAND4_X1 U915 ( .A1(n1206), .A2(KEYINPUT46), .A3(G221), .A4(G234), .ZN(n1205) );
XOR2_X1 U916 ( .A(n986), .B(KEYINPUT3), .Z(n1206) );
XOR2_X1 U917 ( .A(n1207), .B(G472), .Z(n1169) );
NAND4_X1 U918 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1207) );
OR3_X1 U919 ( .A1(n1212), .A2(n1213), .A3(KEYINPUT9), .ZN(n1211) );
NAND2_X1 U920 ( .A1(KEYINPUT9), .A2(n1214), .ZN(n1210) );
NAND2_X1 U921 ( .A1(n1213), .A2(n1212), .ZN(n1208) );
NAND2_X1 U922 ( .A1(KEYINPUT34), .A2(n1215), .ZN(n1212) );
INV_X1 U923 ( .A(n1214), .ZN(n1215) );
XOR2_X1 U924 ( .A(n1099), .B(G101), .Z(n1214) );
NAND2_X1 U925 ( .A1(G210), .A2(n1216), .ZN(n1099) );
XNOR2_X1 U926 ( .A(n1217), .B(n1218), .ZN(n1213) );
XOR2_X1 U927 ( .A(n1047), .B(n1095), .Z(n1218) );
XOR2_X1 U928 ( .A(n1219), .B(n1220), .Z(n1095) );
NOR2_X1 U929 ( .A1(KEYINPUT5), .A2(n1221), .ZN(n1220) );
XOR2_X1 U930 ( .A(n1222), .B(G119), .Z(n1221) );
NAND2_X1 U931 ( .A1(KEYINPUT29), .A2(n1223), .ZN(n1222) );
XNOR2_X1 U932 ( .A(G113), .B(KEYINPUT53), .ZN(n1217) );
INV_X1 U933 ( .A(n1089), .ZN(n1130) );
NAND3_X1 U934 ( .A1(n1153), .A2(n981), .A3(n975), .ZN(n1089) );
NOR2_X1 U935 ( .A1(n1005), .A2(n1004), .ZN(n975) );
INV_X1 U936 ( .A(n1187), .ZN(n1004) );
NAND2_X1 U937 ( .A1(G221), .A2(n1191), .ZN(n1187) );
NAND2_X1 U938 ( .A1(G234), .A2(n1209), .ZN(n1191) );
XOR2_X1 U939 ( .A(n1224), .B(G469), .Z(n1005) );
NAND2_X1 U940 ( .A1(n1225), .A2(n1209), .ZN(n1224) );
XOR2_X1 U941 ( .A(n1226), .B(n1227), .Z(n1225) );
XOR2_X1 U942 ( .A(KEYINPUT23), .B(n1228), .Z(n1227) );
NOR2_X1 U943 ( .A1(KEYINPUT11), .A2(n1229), .ZN(n1228) );
XNOR2_X1 U944 ( .A(n1118), .B(n1120), .ZN(n1229) );
XOR2_X1 U945 ( .A(G140), .B(n1189), .Z(n1120) );
INV_X1 U946 ( .A(G110), .ZN(n1189) );
NAND2_X1 U947 ( .A1(G227), .A2(n986), .ZN(n1118) );
XOR2_X1 U948 ( .A(n1104), .B(n1230), .Z(n1226) );
NOR2_X1 U949 ( .A1(KEYINPUT40), .A2(n1109), .ZN(n1230) );
XOR2_X1 U950 ( .A(n1047), .B(KEYINPUT7), .Z(n1109) );
XOR2_X1 U951 ( .A(n1219), .B(n1231), .Z(n1104) );
NOR2_X1 U952 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
XOR2_X1 U953 ( .A(n1234), .B(KEYINPUT19), .Z(n1233) );
NAND2_X1 U954 ( .A1(n1235), .A2(n1167), .ZN(n1234) );
INV_X1 U955 ( .A(G101), .ZN(n1167) );
XOR2_X1 U956 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U957 ( .A(KEYINPUT61), .B(KEYINPUT59), .Z(n1237) );
AND2_X1 U958 ( .A1(n1236), .A2(G101), .ZN(n1232) );
XOR2_X1 U959 ( .A(n1238), .B(n1046), .Z(n1219) );
XNOR2_X1 U960 ( .A(G134), .B(n1158), .ZN(n1046) );
INV_X1 U961 ( .A(G137), .ZN(n1158) );
XNOR2_X1 U962 ( .A(KEYINPUT36), .B(n1239), .ZN(n1238) );
NOR2_X1 U963 ( .A1(G131), .A2(KEYINPUT1), .ZN(n1239) );
NAND2_X1 U964 ( .A1(n1019), .A2(n1240), .ZN(n981) );
NAND2_X1 U965 ( .A1(n1171), .A2(n1066), .ZN(n1240) );
INV_X1 U966 ( .A(G898), .ZN(n1066) );
AND3_X1 U967 ( .A1(n1241), .A2(n1242), .A3(G953), .ZN(n1171) );
XOR2_X1 U968 ( .A(KEYINPUT17), .B(G902), .Z(n1241) );
NAND3_X1 U969 ( .A1(n1242), .A2(n986), .A3(G952), .ZN(n1019) );
NAND2_X1 U970 ( .A1(G237), .A2(G234), .ZN(n1242) );
INV_X1 U971 ( .A(n980), .ZN(n1153) );
NAND2_X1 U972 ( .A1(n1243), .A2(n1018), .ZN(n980) );
NAND2_X1 U973 ( .A1(G214), .A2(n1244), .ZN(n1018) );
XNOR2_X1 U974 ( .A(n1017), .B(KEYINPUT8), .ZN(n1243) );
XNOR2_X1 U975 ( .A(n1245), .B(n1126), .ZN(n1017) );
INV_X1 U976 ( .A(n1031), .ZN(n1126) );
NAND2_X1 U977 ( .A1(G210), .A2(n1244), .ZN(n1031) );
NAND2_X1 U978 ( .A1(n1246), .A2(n1209), .ZN(n1244) );
INV_X1 U979 ( .A(G237), .ZN(n1246) );
NAND2_X1 U980 ( .A1(KEYINPUT30), .A2(n1029), .ZN(n1245) );
NAND2_X1 U981 ( .A1(n1247), .A2(n1209), .ZN(n1029) );
XOR2_X1 U982 ( .A(n1248), .B(n1249), .Z(n1247) );
XOR2_X1 U983 ( .A(KEYINPUT32), .B(KEYINPUT26), .Z(n1249) );
XOR2_X1 U984 ( .A(n1062), .B(n1122), .Z(n1248) );
XOR2_X1 U985 ( .A(n1250), .B(n1047), .Z(n1122) );
XOR2_X1 U986 ( .A(n1151), .B(n1251), .Z(n1047) );
INV_X1 U987 ( .A(G146), .ZN(n1151) );
XNOR2_X1 U988 ( .A(G125), .B(n1252), .ZN(n1250) );
NOR2_X1 U989 ( .A1(G953), .A2(n1065), .ZN(n1252) );
INV_X1 U990 ( .A(G224), .ZN(n1065) );
XOR2_X1 U991 ( .A(n1253), .B(n1254), .Z(n1062) );
XOR2_X1 U992 ( .A(n1255), .B(n1096), .Z(n1254) );
XOR2_X1 U993 ( .A(G101), .B(G113), .Z(n1096) );
XOR2_X1 U994 ( .A(n1256), .B(n1257), .Z(n1253) );
XOR2_X1 U995 ( .A(G119), .B(G110), .Z(n1257) );
NAND2_X1 U996 ( .A1(KEYINPUT60), .A2(n1236), .ZN(n1256) );
XOR2_X1 U997 ( .A(G104), .B(G107), .Z(n1236) );
NOR2_X1 U998 ( .A1(n1024), .A2(n1155), .ZN(n1000) );
XOR2_X1 U999 ( .A(n1028), .B(G475), .Z(n1155) );
NOR2_X1 U1000 ( .A1(n1086), .A2(G902), .ZN(n1028) );
XOR2_X1 U1001 ( .A(n1258), .B(n1259), .Z(n1086) );
XOR2_X1 U1002 ( .A(n1260), .B(n1261), .Z(n1259) );
XOR2_X1 U1003 ( .A(G122), .B(G113), .Z(n1261) );
XOR2_X1 U1004 ( .A(G143), .B(G131), .Z(n1260) );
XOR2_X1 U1005 ( .A(n1262), .B(n1263), .Z(n1258) );
AND2_X1 U1006 ( .A1(n1216), .A2(G214), .ZN(n1263) );
NOR2_X1 U1007 ( .A1(G953), .A2(G237), .ZN(n1216) );
XOR2_X1 U1008 ( .A(n1264), .B(G104), .Z(n1262) );
NAND2_X1 U1009 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NAND2_X1 U1010 ( .A1(n1203), .A2(n1040), .ZN(n1266) );
XOR2_X1 U1011 ( .A(KEYINPUT45), .B(n1267), .Z(n1265) );
NOR2_X1 U1012 ( .A1(n1203), .A2(n1040), .ZN(n1267) );
XNOR2_X1 U1013 ( .A(G125), .B(G140), .ZN(n1040) );
XNOR2_X1 U1014 ( .A(G146), .B(KEYINPUT24), .ZN(n1203) );
INV_X1 U1015 ( .A(n1186), .ZN(n1024) );
XOR2_X1 U1016 ( .A(n1268), .B(G478), .Z(n1186) );
NAND2_X1 U1017 ( .A1(n1080), .A2(n1209), .ZN(n1268) );
INV_X1 U1018 ( .A(G902), .ZN(n1209) );
XNOR2_X1 U1019 ( .A(n1269), .B(n1270), .ZN(n1080) );
XOR2_X1 U1020 ( .A(G107), .B(n1271), .Z(n1270) );
XOR2_X1 U1021 ( .A(KEYINPUT6), .B(G134), .Z(n1271) );
XOR2_X1 U1022 ( .A(n1272), .B(n1251), .Z(n1269) );
XOR2_X1 U1023 ( .A(G128), .B(G143), .Z(n1251) );
XOR2_X1 U1024 ( .A(n1273), .B(n1255), .Z(n1272) );
XNOR2_X1 U1025 ( .A(G122), .B(n1223), .ZN(n1255) );
INV_X1 U1026 ( .A(G116), .ZN(n1223) );
NAND3_X1 U1027 ( .A1(G234), .A2(n986), .A3(G217), .ZN(n1273) );
INV_X1 U1028 ( .A(G953), .ZN(n986) );
endmodule


