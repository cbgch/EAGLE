//Key = 0111110011001011000100010110111111100001101011110000001100001110


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
n2385, n2386, n2387, n2388;

OR2_X1 U1328 ( .A1(n2388), .A2(n1796), .ZN(U280) );
OR2_X1 U1329 ( .A1(n1940), .A2(STATO_REG_0__SCAN_IN), .ZN(n1795) );
INV_X2 U1330 ( .A(n1795), .ZN(n1796) );
INV_X2 U1331 ( .A(U280), .ZN(n1797) );
XNOR2_X1 U1332 ( .A(KEYINPUT49), .B(n1798), .ZN(U375) );
NAND2_X1 U1333 ( .A1(n1799), .A2(n1800), .ZN(U344) );
NAND2_X1 U1334 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1801), .ZN(n1800) );
NAND2_X1 U1335 ( .A1(n1802), .A2(DATA_IN_7_), .ZN(n1799) );
NAND2_X1 U1336 ( .A1(n1803), .A2(n1804), .ZN(U343) );
NAND2_X1 U1337 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1801), .ZN(n1804) );
NAND2_X1 U1338 ( .A1(n1802), .A2(DATA_IN_6_), .ZN(n1803) );
NAND2_X1 U1339 ( .A1(n1805), .A2(n1806), .ZN(U342) );
NAND2_X1 U1340 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1801), .ZN(n1806) );
NAND2_X1 U1341 ( .A1(n1802), .A2(DATA_IN_5_), .ZN(n1805) );
NAND2_X1 U1342 ( .A1(n1807), .A2(n1808), .ZN(U341) );
NAND2_X1 U1343 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1801), .ZN(n1808) );
NAND2_X1 U1344 ( .A1(n1802), .A2(DATA_IN_4_), .ZN(n1807) );
NAND2_X1 U1345 ( .A1(n1809), .A2(n1810), .ZN(U340) );
NAND2_X1 U1346 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1801), .ZN(n1810) );
NAND2_X1 U1347 ( .A1(n1802), .A2(DATA_IN_3_), .ZN(n1809) );
NAND2_X1 U1348 ( .A1(n1811), .A2(n1812), .ZN(U339) );
NAND2_X1 U1349 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1801), .ZN(n1812) );
NAND2_X1 U1350 ( .A1(n1802), .A2(DATA_IN_2_), .ZN(n1811) );
NAND2_X1 U1351 ( .A1(n1813), .A2(n1814), .ZN(U338) );
NAND2_X1 U1352 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1801), .ZN(n1814) );
NAND2_X1 U1353 ( .A1(n1802), .A2(DATA_IN_1_), .ZN(n1813) );
NAND2_X1 U1354 ( .A1(n1815), .A2(n1816), .ZN(U337) );
NAND2_X1 U1355 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1801), .ZN(n1816) );
NAND2_X1 U1356 ( .A1(n1802), .A2(DATA_IN_0_), .ZN(n1815) );
INV_X1 U1357 ( .A(n1801), .ZN(n1802) );
NAND2_X1 U1358 ( .A1(n1798), .A2(n1817), .ZN(n1801) );
NAND3_X1 U1359 ( .A1(n1818), .A2(n1819), .A3(n1820), .ZN(n1817) );
NAND2_X1 U1360 ( .A1(n1821), .A2(n1822), .ZN(U336) );
NAND2_X1 U1361 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1823), .ZN(n1822) );
XOR2_X1 U1362 ( .A(KEYINPUT30), .B(n1824), .Z(n1821) );
NOR2_X1 U1363 ( .A1(n1825), .A2(n1826), .ZN(n1824) );
XNOR2_X1 U1364 ( .A(DATA_IN_7_), .B(KEYINPUT22), .ZN(n1826) );
INV_X1 U1365 ( .A(n1827), .ZN(n1825) );
NAND2_X1 U1366 ( .A1(n1828), .A2(n1829), .ZN(U335) );
NAND2_X1 U1367 ( .A1(DATA_IN_6_), .A2(n1827), .ZN(n1829) );
NAND2_X1 U1368 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1823), .ZN(n1828) );
NAND2_X1 U1369 ( .A1(n1830), .A2(n1831), .ZN(U334) );
NAND2_X1 U1370 ( .A1(DATA_IN_5_), .A2(n1832), .ZN(n1831) );
XNOR2_X1 U1371 ( .A(KEYINPUT42), .B(n1827), .ZN(n1832) );
NAND2_X1 U1372 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1823), .ZN(n1830) );
NAND2_X1 U1373 ( .A1(n1833), .A2(n1834), .ZN(U333) );
NAND2_X1 U1374 ( .A1(n1835), .A2(n1827), .ZN(n1834) );
XNOR2_X1 U1375 ( .A(DATA_IN_4_), .B(KEYINPUT32), .ZN(n1835) );
NAND2_X1 U1376 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1823), .ZN(n1833) );
NAND2_X1 U1377 ( .A1(n1836), .A2(n1837), .ZN(U332) );
NAND2_X1 U1378 ( .A1(DATA_IN_3_), .A2(n1827), .ZN(n1837) );
NAND2_X1 U1379 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1823), .ZN(n1836) );
NAND2_X1 U1380 ( .A1(n1838), .A2(n1839), .ZN(U331) );
NAND2_X1 U1381 ( .A1(DATA_IN_2_), .A2(n1827), .ZN(n1839) );
NAND2_X1 U1382 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1823), .ZN(n1838) );
NAND2_X1 U1383 ( .A1(n1840), .A2(n1841), .ZN(U330) );
NAND2_X1 U1384 ( .A1(DATA_IN_1_), .A2(n1827), .ZN(n1841) );
XOR2_X1 U1385 ( .A(KEYINPUT33), .B(n1842), .Z(n1840) );
AND2_X1 U1386 ( .A1(n1823), .A2(RMIN_REG_1__SCAN_IN), .ZN(n1842) );
NAND2_X1 U1387 ( .A1(n1843), .A2(n1844), .ZN(U329) );
NAND2_X1 U1388 ( .A1(DATA_IN_0_), .A2(n1827), .ZN(n1844) );
NAND2_X1 U1389 ( .A1(n1845), .A2(n1846), .ZN(n1827) );
NAND3_X1 U1390 ( .A1(n1847), .A2(n1818), .A3(STATO_REG_1__SCAN_IN), .ZN(n1846) );
NAND2_X1 U1391 ( .A1(n1848), .A2(n1849), .ZN(n1847) );
NAND2_X1 U1392 ( .A1(n1850), .A2(n1820), .ZN(n1849) );
INV_X1 U1393 ( .A(n1851), .ZN(n1850) );
XNOR2_X1 U1394 ( .A(n1819), .B(KEYINPUT5), .ZN(n1845) );
NAND2_X1 U1395 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1823), .ZN(n1843) );
NAND2_X1 U1396 ( .A1(n1798), .A2(n1852), .ZN(n1823) );
NAND2_X1 U1397 ( .A1(n1853), .A2(n1819), .ZN(n1852) );
NAND3_X1 U1398 ( .A1(n1820), .A2(n1818), .A3(n1854), .ZN(n1853) );
NAND2_X1 U1399 ( .A1(n1848), .A2(n1851), .ZN(n1854) );
NAND3_X1 U1400 ( .A1(n1855), .A2(n1856), .A3(n1857), .ZN(n1851) );
NAND2_X1 U1401 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1858), .ZN(n1857) );
NAND3_X1 U1402 ( .A1(n1859), .A2(n1860), .A3(n1861), .ZN(n1856) );
NAND2_X1 U1403 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1862), .ZN(n1861) );
NAND3_X1 U1404 ( .A1(n1863), .A2(n1864), .A3(n1865), .ZN(n1860) );
NAND2_X1 U1405 ( .A1(DATA_IN_5_), .A2(n1866), .ZN(n1865) );
NAND3_X1 U1406 ( .A1(n1867), .A2(n1868), .A3(n1869), .ZN(n1864) );
NAND2_X1 U1407 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1870), .ZN(n1869) );
NAND3_X1 U1408 ( .A1(n1871), .A2(n1872), .A3(n1873), .ZN(n1868) );
NAND2_X1 U1409 ( .A1(DATA_IN_3_), .A2(n1874), .ZN(n1873) );
NAND3_X1 U1410 ( .A1(n1875), .A2(n1876), .A3(n1877), .ZN(n1872) );
NAND2_X1 U1411 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1878), .ZN(n1877) );
NAND3_X1 U1412 ( .A1(n1879), .A2(n1880), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1876) );
NAND2_X1 U1413 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1881), .ZN(n1875) );
NAND2_X1 U1414 ( .A1(n1882), .A2(n1883), .ZN(n1881) );
NAND2_X1 U1415 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1879), .ZN(n1883) );
XNOR2_X1 U1416 ( .A(KEYINPUT10), .B(n1880), .ZN(n1882) );
NAND2_X1 U1417 ( .A1(DATA_IN_2_), .A2(n1884), .ZN(n1871) );
NAND2_X1 U1418 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1885), .ZN(n1867) );
NAND2_X1 U1419 ( .A1(DATA_IN_4_), .A2(n1886), .ZN(n1863) );
NAND2_X1 U1420 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1887), .ZN(n1859) );
NAND2_X1 U1421 ( .A1(DATA_IN_6_), .A2(n1888), .ZN(n1855) );
NAND2_X1 U1422 ( .A1(DATA_IN_7_), .A2(n1889), .ZN(n1848) );
NAND3_X1 U1423 ( .A1(n1890), .A2(n1891), .A3(n1892), .ZN(n1818) );
NAND2_X1 U1424 ( .A1(DATA_IN_7_), .A2(n1893), .ZN(n1892) );
NAND3_X1 U1425 ( .A1(n1894), .A2(n1895), .A3(n1896), .ZN(n1891) );
NAND2_X1 U1426 ( .A1(DATA_IN_6_), .A2(n1897), .ZN(n1896) );
NAND3_X1 U1427 ( .A1(n1898), .A2(n1899), .A3(n1900), .ZN(n1895) );
NAND2_X1 U1428 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1887), .ZN(n1900) );
NAND3_X1 U1429 ( .A1(n1901), .A2(n1902), .A3(n1903), .ZN(n1899) );
NAND2_X1 U1430 ( .A1(DATA_IN_4_), .A2(n1904), .ZN(n1903) );
NAND3_X1 U1431 ( .A1(n1905), .A2(n1906), .A3(n1907), .ZN(n1902) );
NAND2_X1 U1432 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1885), .ZN(n1907) );
NAND3_X1 U1433 ( .A1(n1908), .A2(n1909), .A3(n1910), .ZN(n1906) );
NAND2_X1 U1434 ( .A1(DATA_IN_2_), .A2(n1911), .ZN(n1910) );
NAND3_X1 U1435 ( .A1(n1912), .A2(n1913), .A3(DATA_IN_0_), .ZN(n1909) );
INV_X1 U1436 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1913) );
NAND2_X1 U1437 ( .A1(n1914), .A2(n1880), .ZN(n1912) );
XNOR2_X1 U1438 ( .A(RMAX_REG_1__SCAN_IN), .B(KEYINPUT29), .ZN(n1914) );
NAND2_X1 U1439 ( .A1(DATA_IN_1_), .A2(n1915), .ZN(n1908) );
NAND2_X1 U1440 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1878), .ZN(n1905) );
NAND2_X1 U1441 ( .A1(DATA_IN_3_), .A2(n1916), .ZN(n1901) );
NAND2_X1 U1442 ( .A1(n1917), .A2(RMAX_REG_4__SCAN_IN), .ZN(n1898) );
XNOR2_X1 U1443 ( .A(DATA_IN_4_), .B(KEYINPUT17), .ZN(n1917) );
NAND2_X1 U1444 ( .A1(DATA_IN_5_), .A2(n1918), .ZN(n1894) );
NAND2_X1 U1445 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1919), .ZN(n1890) );
XNOR2_X1 U1446 ( .A(KEYINPUT14), .B(n1862), .ZN(n1919) );
NAND2_X1 U1447 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1858), .ZN(n1820) );
NAND2_X1 U1448 ( .A1(n1920), .A2(n1921), .ZN(U328) );
NAND2_X1 U1449 ( .A1(n1922), .A2(DATA_IN_7_), .ZN(n1921) );
NAND2_X1 U1450 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1923), .ZN(n1920) );
NAND2_X1 U1451 ( .A1(n1924), .A2(n1925), .ZN(U327) );
NAND2_X1 U1452 ( .A1(n1922), .A2(DATA_IN_6_), .ZN(n1925) );
NAND2_X1 U1453 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1923), .ZN(n1924) );
NAND2_X1 U1454 ( .A1(n1926), .A2(n1927), .ZN(U326) );
NAND2_X1 U1455 ( .A1(n1922), .A2(DATA_IN_5_), .ZN(n1927) );
NAND2_X1 U1456 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1923), .ZN(n1926) );
NAND2_X1 U1457 ( .A1(n1928), .A2(n1929), .ZN(U325) );
NAND2_X1 U1458 ( .A1(n1922), .A2(DATA_IN_4_), .ZN(n1929) );
NAND2_X1 U1459 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1923), .ZN(n1928) );
NAND2_X1 U1460 ( .A1(n1930), .A2(n1931), .ZN(U324) );
NAND2_X1 U1461 ( .A1(n1922), .A2(DATA_IN_3_), .ZN(n1931) );
NAND2_X1 U1462 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1923), .ZN(n1930) );
NAND2_X1 U1463 ( .A1(n1932), .A2(n1933), .ZN(U323) );
NAND2_X1 U1464 ( .A1(n1922), .A2(DATA_IN_2_), .ZN(n1933) );
NAND2_X1 U1465 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1923), .ZN(n1932) );
NAND2_X1 U1466 ( .A1(n1934), .A2(n1935), .ZN(U322) );
NAND2_X1 U1467 ( .A1(n1922), .A2(DATA_IN_1_), .ZN(n1935) );
NAND2_X1 U1468 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1923), .ZN(n1934) );
NAND2_X1 U1469 ( .A1(n1936), .A2(n1937), .ZN(U321) );
NAND2_X1 U1470 ( .A1(n1922), .A2(DATA_IN_0_), .ZN(n1937) );
AND2_X1 U1471 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1938), .ZN(n1922) );
NAND2_X1 U1472 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1923), .ZN(n1936) );
NAND2_X1 U1473 ( .A1(n1798), .A2(n1938), .ZN(n1923) );
NAND2_X1 U1474 ( .A1(n1819), .A2(n1939), .ZN(n1938) );
NAND2_X1 U1475 ( .A1(n1940), .A2(n1819), .ZN(n1798) );
NAND2_X1 U1476 ( .A1(n1941), .A2(n1942), .ZN(U320) );
NAND2_X1 U1477 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1797), .ZN(n1942) );
NAND2_X1 U1478 ( .A1(n1796), .A2(DATA_IN_7_), .ZN(n1941) );
NAND2_X1 U1479 ( .A1(n1943), .A2(n1944), .ZN(U319) );
NAND2_X1 U1480 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1797), .ZN(n1944) );
NAND2_X1 U1481 ( .A1(n1796), .A2(DATA_IN_6_), .ZN(n1943) );
NAND2_X1 U1482 ( .A1(n1945), .A2(n1946), .ZN(U318) );
NAND2_X1 U1483 ( .A1(n1796), .A2(DATA_IN_5_), .ZN(n1946) );
XOR2_X1 U1484 ( .A(KEYINPUT3), .B(n1947), .Z(n1945) );
NOR2_X1 U1485 ( .A1(U280), .A2(n1948), .ZN(n1947) );
XOR2_X1 U1486 ( .A(REG1_REG_5__SCAN_IN), .B(KEYINPUT62), .Z(n1948) );
NAND2_X1 U1487 ( .A1(n1949), .A2(n1950), .ZN(U317) );
NAND2_X1 U1488 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1797), .ZN(n1950) );
NAND2_X1 U1489 ( .A1(n1796), .A2(DATA_IN_4_), .ZN(n1949) );
NAND2_X1 U1490 ( .A1(n1951), .A2(n1952), .ZN(U316) );
NAND2_X1 U1491 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1797), .ZN(n1952) );
NAND2_X1 U1492 ( .A1(n1796), .A2(DATA_IN_3_), .ZN(n1951) );
NAND2_X1 U1493 ( .A1(n1953), .A2(n1954), .ZN(U315) );
NAND2_X1 U1494 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1797), .ZN(n1954) );
NAND2_X1 U1495 ( .A1(n1796), .A2(DATA_IN_2_), .ZN(n1953) );
NAND2_X1 U1496 ( .A1(n1955), .A2(n1956), .ZN(U314) );
NAND2_X1 U1497 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1957), .ZN(n1956) );
XNOR2_X1 U1498 ( .A(KEYINPUT56), .B(U280), .ZN(n1957) );
NAND2_X1 U1499 ( .A1(n1796), .A2(DATA_IN_1_), .ZN(n1955) );
NAND2_X1 U1500 ( .A1(n1958), .A2(n1959), .ZN(U313) );
NAND2_X1 U1501 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1797), .ZN(n1959) );
NAND2_X1 U1502 ( .A1(n1796), .A2(DATA_IN_0_), .ZN(n1958) );
NAND2_X1 U1503 ( .A1(n1960), .A2(n1961), .ZN(U312) );
NAND2_X1 U1504 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1797), .ZN(n1961) );
NAND2_X1 U1505 ( .A1(n1796), .A2(REG1_REG_7__SCAN_IN), .ZN(n1960) );
NAND2_X1 U1506 ( .A1(n1962), .A2(n1963), .ZN(U311) );
NAND2_X1 U1507 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1797), .ZN(n1963) );
NAND2_X1 U1508 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1796), .ZN(n1962) );
NAND2_X1 U1509 ( .A1(n1964), .A2(n1965), .ZN(U310) );
NAND2_X1 U1510 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1797), .ZN(n1965) );
NAND2_X1 U1511 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1796), .ZN(n1964) );
NAND2_X1 U1512 ( .A1(n1966), .A2(n1967), .ZN(U309) );
NAND2_X1 U1513 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1797), .ZN(n1967) );
NAND2_X1 U1514 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1796), .ZN(n1966) );
NAND2_X1 U1515 ( .A1(n1968), .A2(n1969), .ZN(U308) );
NAND2_X1 U1516 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1797), .ZN(n1969) );
NAND2_X1 U1517 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1796), .ZN(n1968) );
NAND2_X1 U1518 ( .A1(n1970), .A2(n1971), .ZN(U307) );
NAND2_X1 U1519 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1797), .ZN(n1971) );
NAND2_X1 U1520 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1796), .ZN(n1970) );
NAND2_X1 U1521 ( .A1(n1972), .A2(n1973), .ZN(U306) );
NAND2_X1 U1522 ( .A1(n1974), .A2(n1797), .ZN(n1973) );
XOR2_X1 U1523 ( .A(REG2_REG_1__SCAN_IN), .B(KEYINPUT41), .Z(n1974) );
NAND2_X1 U1524 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1796), .ZN(n1972) );
NAND2_X1 U1525 ( .A1(n1975), .A2(n1976), .ZN(U305) );
NAND2_X1 U1526 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1797), .ZN(n1976) );
NAND2_X1 U1527 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1796), .ZN(n1975) );
NAND2_X1 U1528 ( .A1(n1977), .A2(n1978), .ZN(U304) );
NAND2_X1 U1529 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1797), .ZN(n1978) );
NAND2_X1 U1530 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1796), .ZN(n1977) );
NAND2_X1 U1531 ( .A1(n1979), .A2(n1980), .ZN(U303) );
NAND2_X1 U1532 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1981), .ZN(n1980) );
XNOR2_X1 U1533 ( .A(KEYINPUT11), .B(U280), .ZN(n1981) );
NAND2_X1 U1534 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1796), .ZN(n1979) );
NAND2_X1 U1535 ( .A1(n1982), .A2(n1983), .ZN(U302) );
NAND2_X1 U1536 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1797), .ZN(n1983) );
NAND2_X1 U1537 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1796), .ZN(n1982) );
NAND2_X1 U1538 ( .A1(n1984), .A2(n1985), .ZN(U301) );
NAND2_X1 U1539 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1797), .ZN(n1985) );
NAND2_X1 U1540 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1796), .ZN(n1984) );
NAND2_X1 U1541 ( .A1(n1986), .A2(n1987), .ZN(U300) );
NAND2_X1 U1542 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1797), .ZN(n1987) );
NAND2_X1 U1543 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1796), .ZN(n1986) );
NAND2_X1 U1544 ( .A1(n1988), .A2(n1989), .ZN(U299) );
NAND2_X1 U1545 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1797), .ZN(n1989) );
NAND2_X1 U1546 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1796), .ZN(n1988) );
NAND2_X1 U1547 ( .A1(n1990), .A2(n1991), .ZN(U298) );
NAND2_X1 U1548 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1992), .ZN(n1991) );
XNOR2_X1 U1549 ( .A(KEYINPUT51), .B(U280), .ZN(n1992) );
NAND2_X1 U1550 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1796), .ZN(n1990) );
NAND2_X1 U1551 ( .A1(n1993), .A2(n1994), .ZN(U297) );
NAND2_X1 U1552 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1797), .ZN(n1994) );
NAND2_X1 U1553 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1796), .ZN(n1993) );
NAND2_X1 U1554 ( .A1(n1995), .A2(n1996), .ZN(U296) );
NAND2_X1 U1555 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1797), .ZN(n1996) );
NAND2_X1 U1556 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1796), .ZN(n1995) );
NAND2_X1 U1557 ( .A1(n1997), .A2(n1998), .ZN(U295) );
NAND2_X1 U1558 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1797), .ZN(n1998) );
NAND2_X1 U1559 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1796), .ZN(n1997) );
NAND2_X1 U1560 ( .A1(n1999), .A2(n2000), .ZN(U294) );
NAND2_X1 U1561 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1797), .ZN(n2000) );
NAND2_X1 U1562 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1796), .ZN(n1999) );
NAND2_X1 U1563 ( .A1(n2001), .A2(n2002), .ZN(U293) );
NAND2_X1 U1564 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1797), .ZN(n2002) );
NAND2_X1 U1565 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1796), .ZN(n2001) );
NAND2_X1 U1566 ( .A1(n2003), .A2(n2004), .ZN(U292) );
NAND2_X1 U1567 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1797), .ZN(n2004) );
NAND2_X1 U1568 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1796), .ZN(n2003) );
NAND2_X1 U1569 ( .A1(n2005), .A2(n2006), .ZN(U291) );
NAND2_X1 U1570 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1797), .ZN(n2006) );
NAND2_X1 U1571 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1796), .ZN(n2005) );
NAND2_X1 U1572 ( .A1(n2007), .A2(n2008), .ZN(U290) );
NAND2_X1 U1573 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1797), .ZN(n2008) );
NAND2_X1 U1574 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1796), .ZN(n2007) );
NAND2_X1 U1575 ( .A1(n2009), .A2(n2010), .ZN(U289) );
NAND2_X1 U1576 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1797), .ZN(n2010) );
NAND2_X1 U1577 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1796), .ZN(n2009) );
NAND4_X1 U1578 ( .A1(n2011), .A2(n2012), .A3(n2013), .A4(n2014), .ZN(U288));
NAND2_X1 U1579 ( .A1(n2015), .A2(REG4_REG_7__SCAN_IN), .ZN(n2014) );
NOR2_X1 U1580 ( .A1(n2016), .A2(n2017), .ZN(n2013) );
NOR2_X1 U1581 ( .A1(n2018), .A2(n2019), .ZN(n2017) );
XNOR2_X1 U1582 ( .A(KEYINPUT45), .B(n2020), .ZN(n2019) );
NOR3_X1 U1583 ( .A1(n2021), .A2(n2022), .A3(n2023), .ZN(n2016) );
NAND2_X1 U1584 ( .A1(n2024), .A2(RLAST_REG_7__SCAN_IN), .ZN(n2012) );
NAND2_X1 U1585 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1797), .ZN(n2011) );
NAND4_X1 U1586 ( .A1(n2025), .A2(n2026), .A3(n2027), .A4(n2028), .ZN(U287));
NOR2_X1 U1587 ( .A1(n2029), .A2(n2030), .ZN(n2028) );
AND2_X1 U1588 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n2024), .ZN(n2030) );
NOR2_X1 U1589 ( .A1(n2031), .A2(n2032), .ZN(n2029) );
NAND2_X1 U1590 ( .A1(n2033), .A2(n2034), .ZN(n2027) );
NAND2_X1 U1591 ( .A1(n2035), .A2(n2036), .ZN(n2034) );
NAND2_X1 U1592 ( .A1(n2037), .A2(n2038), .ZN(n2036) );
XNOR2_X1 U1593 ( .A(n2039), .B(KEYINPUT48), .ZN(n2035) );
NAND2_X1 U1594 ( .A1(n2040), .A2(n2041), .ZN(n2026) );
INV_X1 U1595 ( .A(n2023), .ZN(n2041) );
XOR2_X1 U1596 ( .A(n2021), .B(n2042), .Z(n2040) );
XOR2_X1 U1597 ( .A(KEYINPUT39), .B(n2022), .Z(n2042) );
NAND2_X1 U1598 ( .A1(n2043), .A2(n1797), .ZN(n2025) );
XNOR2_X1 U1599 ( .A(KEYINPUT26), .B(DATA_OUT_REG_6__SCAN_IN), .ZN(n2043) );
NAND4_X1 U1600 ( .A1(n2044), .A2(n2045), .A3(n2046), .A4(n2047), .ZN(U286));
NOR3_X1 U1601 ( .A1(n2048), .A2(n2049), .A3(n2050), .ZN(n2047) );
NOR2_X1 U1602 ( .A1(n2051), .A2(n2018), .ZN(n2050) );
NOR2_X1 U1603 ( .A1(n2052), .A2(n2039), .ZN(n2051) );
INV_X1 U1604 ( .A(n2020), .ZN(n2039) );
NAND3_X1 U1605 ( .A1(n2053), .A2(n2054), .A3(n2055), .ZN(n2020) );
XNOR2_X1 U1606 ( .A(n2056), .B(KEYINPUT31), .ZN(n2055) );
NOR2_X1 U1607 ( .A1(n2037), .A2(n2057), .ZN(n2052) );
NOR2_X1 U1608 ( .A1(n2058), .A2(n2059), .ZN(n2057) );
NOR2_X1 U1609 ( .A1(n2056), .A2(n2054), .ZN(n2058) );
INV_X1 U1610 ( .A(n2053), .ZN(n2037) );
NAND2_X1 U1611 ( .A1(n2060), .A2(n2059), .ZN(n2053) );
XNOR2_X1 U1612 ( .A(n2056), .B(n2061), .ZN(n2060) );
AND2_X1 U1613 ( .A1(n2054), .A2(KEYINPUT31), .ZN(n2061) );
NOR3_X1 U1614 ( .A1(n2062), .A2(n2022), .A3(n2023), .ZN(n2049) );
AND2_X1 U1615 ( .A1(n2063), .A2(n2064), .ZN(n2022) );
XNOR2_X1 U1616 ( .A(KEYINPUT4), .B(n2065), .ZN(n2064) );
XOR2_X1 U1617 ( .A(KEYINPUT59), .B(n2066), .Z(n2062) );
NOR2_X1 U1618 ( .A1(n2063), .A2(n2065), .ZN(n2066) );
NAND2_X1 U1619 ( .A1(n2021), .A2(n2067), .ZN(n2065) );
NAND2_X1 U1620 ( .A1(n2038), .A2(n2068), .ZN(n2067) );
INV_X1 U1621 ( .A(n2054), .ZN(n2038) );
NAND2_X1 U1622 ( .A1(n2069), .A2(n2054), .ZN(n2021) );
NOR2_X1 U1623 ( .A1(n2054), .A2(n2070), .ZN(n2048) );
NAND2_X1 U1624 ( .A1(n2071), .A2(n2072), .ZN(n2054) );
NAND3_X1 U1625 ( .A1(n2073), .A2(n2074), .A3(n2075), .ZN(n2072) );
XOR2_X1 U1626 ( .A(n2076), .B(n2077), .Z(n2075) );
NAND2_X1 U1627 ( .A1(n2078), .A2(n2079), .ZN(n2074) );
NAND2_X1 U1628 ( .A1(n2080), .A2(n2081), .ZN(n2073) );
NAND3_X1 U1629 ( .A1(n2078), .A2(n2082), .A3(n2083), .ZN(n2071) );
XOR2_X1 U1630 ( .A(n2084), .B(n2076), .Z(n2083) );
NAND2_X1 U1631 ( .A1(n2085), .A2(n2086), .ZN(n2076) );
NAND2_X1 U1632 ( .A1(RESTART), .A2(n1888), .ZN(n2086) );
NAND2_X1 U1633 ( .A1(n2031), .A2(n2087), .ZN(n2085) );
INV_X1 U1634 ( .A(REG4_REG_6__SCAN_IN), .ZN(n2031) );
NAND2_X1 U1635 ( .A1(KEYINPUT44), .A2(n2077), .ZN(n2084) );
NAND2_X1 U1636 ( .A1(n2088), .A2(n2089), .ZN(n2077) );
NAND2_X1 U1637 ( .A1(RESTART), .A2(n1897), .ZN(n2089) );
INV_X1 U1638 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1897) );
NAND2_X1 U1639 ( .A1(n1862), .A2(n2087), .ZN(n2088) );
NAND2_X1 U1640 ( .A1(n2090), .A2(n2091), .ZN(n2082) );
NAND2_X1 U1641 ( .A1(n2092), .A2(n2080), .ZN(n2091) );
XNOR2_X1 U1642 ( .A(n2093), .B(KEYINPUT6), .ZN(n2092) );
INV_X1 U1643 ( .A(n2079), .ZN(n2090) );
NAND2_X1 U1644 ( .A1(n2094), .A2(n2093), .ZN(n2078) );
NAND2_X1 U1645 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1797), .ZN(n2046) );
NAND2_X1 U1646 ( .A1(n2015), .A2(REG4_REG_5__SCAN_IN), .ZN(n2045) );
NAND2_X1 U1647 ( .A1(n2024), .A2(RLAST_REG_5__SCAN_IN), .ZN(n2044) );
NAND4_X1 U1648 ( .A1(n2095), .A2(n2096), .A3(n2097), .A4(n2098), .ZN(U285));
NOR3_X1 U1649 ( .A1(n2099), .A2(n2100), .A3(n2101), .ZN(n2098) );
NOR3_X1 U1650 ( .A1(n2018), .A2(n2059), .A3(n2102), .ZN(n2101) );
NOR2_X1 U1651 ( .A1(n2103), .A2(n2104), .ZN(n2102) );
AND2_X1 U1652 ( .A1(n2105), .A2(n2106), .ZN(n2103) );
AND3_X1 U1653 ( .A1(n2105), .A2(n2104), .A3(n2106), .ZN(n2059) );
NAND2_X1 U1654 ( .A1(n2107), .A2(n2108), .ZN(n2104) );
NAND2_X1 U1655 ( .A1(n2109), .A2(n2110), .ZN(n2108) );
OR2_X1 U1656 ( .A1(n2111), .A2(n2112), .ZN(n2109) );
INV_X1 U1657 ( .A(n2056), .ZN(n2107) );
NOR3_X1 U1658 ( .A1(n2110), .A2(n2112), .A3(n2111), .ZN(n2056) );
NOR3_X1 U1659 ( .A1(n2023), .A2(n2063), .A3(n2113), .ZN(n2100) );
NOR2_X1 U1660 ( .A1(n2114), .A2(n2115), .ZN(n2113) );
AND2_X1 U1661 ( .A1(n2116), .A2(n2117), .ZN(n2114) );
AND3_X1 U1662 ( .A1(n2116), .A2(n2115), .A3(n2117), .ZN(n2063) );
NAND2_X1 U1663 ( .A1(n2068), .A2(n2118), .ZN(n2115) );
NAND2_X1 U1664 ( .A1(n2119), .A2(n2110), .ZN(n2118) );
OR2_X1 U1665 ( .A1(n2120), .A2(n2112), .ZN(n2119) );
INV_X1 U1666 ( .A(n2069), .ZN(n2068) );
NOR3_X1 U1667 ( .A1(n2120), .A2(n2112), .A3(n2110), .ZN(n2069) );
NOR2_X1 U1668 ( .A1(n2121), .A2(n2122), .ZN(n2099) );
XOR2_X1 U1669 ( .A(RLAST_REG_4__SCAN_IN), .B(KEYINPUT47), .Z(n2122) );
NAND2_X1 U1670 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1797), .ZN(n2097) );
NAND2_X1 U1671 ( .A1(n2123), .A2(n2110), .ZN(n2096) );
NAND2_X1 U1672 ( .A1(n2124), .A2(n2125), .ZN(n2110) );
NAND2_X1 U1673 ( .A1(n2126), .A2(n2079), .ZN(n2125) );
NAND2_X1 U1674 ( .A1(n2127), .A2(n2128), .ZN(n2126) );
NAND2_X1 U1675 ( .A1(n2093), .A2(n2080), .ZN(n2128) );
INV_X1 U1676 ( .A(n2081), .ZN(n2093) );
XOR2_X1 U1677 ( .A(n2129), .B(KEYINPUT27), .Z(n2127) );
NAND2_X1 U1678 ( .A1(n2130), .A2(n2081), .ZN(n2129) );
XNOR2_X1 U1679 ( .A(n2094), .B(KEYINPUT28), .ZN(n2130) );
INV_X1 U1680 ( .A(n2080), .ZN(n2094) );
XOR2_X1 U1681 ( .A(KEYINPUT1), .B(n2131), .Z(n2124) );
NOR2_X1 U1682 ( .A1(n2132), .A2(n2079), .ZN(n2131) );
NAND2_X1 U1683 ( .A1(n2133), .A2(n2134), .ZN(n2079) );
NAND2_X1 U1684 ( .A1(n2135), .A2(n2136), .ZN(n2134) );
XNOR2_X1 U1685 ( .A(n2137), .B(KEYINPUT16), .ZN(n2135) );
XNOR2_X1 U1686 ( .A(n2138), .B(n2081), .ZN(n2132) );
NAND3_X1 U1687 ( .A1(n2139), .A2(n2140), .A3(n2141), .ZN(n2081) );
NAND2_X1 U1688 ( .A1(n2142), .A2(n1918), .ZN(n2141) );
INV_X1 U1689 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1918) );
NAND2_X1 U1690 ( .A1(DATA_IN_5_), .A2(n2087), .ZN(n2142) );
OR3_X1 U1691 ( .A1(DATA_IN_5_), .A2(KEYINPUT52), .A3(RESTART), .ZN(n2140) );
NAND2_X1 U1692 ( .A1(KEYINPUT52), .A2(RESTART), .ZN(n2139) );
NAND2_X1 U1693 ( .A1(KEYINPUT19), .A2(n2080), .ZN(n2138) );
NAND2_X1 U1694 ( .A1(n2143), .A2(n2144), .ZN(n2080) );
NAND2_X1 U1695 ( .A1(RESTART), .A2(n1866), .ZN(n2144) );
NAND2_X1 U1696 ( .A1(n2145), .A2(n2087), .ZN(n2143) );
NAND2_X1 U1697 ( .A1(n2015), .A2(REG4_REG_4__SCAN_IN), .ZN(n2095) );
NAND4_X1 U1698 ( .A1(n2146), .A2(n2147), .A3(n2148), .A4(n2149), .ZN(U284));
NOR3_X1 U1699 ( .A1(n2150), .A2(n2151), .A3(n2152), .ZN(n2149) );
NOR2_X1 U1700 ( .A1(n2153), .A2(n2070), .ZN(n2152) );
NOR2_X1 U1701 ( .A1(n2018), .A2(n2154), .ZN(n2151) );
XNOR2_X1 U1702 ( .A(n2105), .B(n2155), .ZN(n2154) );
NOR2_X1 U1703 ( .A1(KEYINPUT20), .A2(n2156), .ZN(n2155) );
XNOR2_X1 U1704 ( .A(n2112), .B(n2111), .ZN(n2105) );
NOR2_X1 U1705 ( .A1(n2157), .A2(n2032), .ZN(n2150) );
XOR2_X1 U1706 ( .A(KEYINPUT9), .B(n2158), .Z(n2148) );
NOR2_X1 U1707 ( .A1(n2023), .A2(n2159), .ZN(n2158) );
XNOR2_X1 U1708 ( .A(n2117), .B(n2116), .ZN(n2159) );
XNOR2_X1 U1709 ( .A(n2120), .B(n2112), .ZN(n2116) );
INV_X1 U1710 ( .A(n2153), .ZN(n2112) );
NAND2_X1 U1711 ( .A1(n2160), .A2(n2161), .ZN(n2153) );
NAND2_X1 U1712 ( .A1(n2137), .A2(n2162), .ZN(n2161) );
NAND2_X1 U1713 ( .A1(n2163), .A2(n2164), .ZN(n2162) );
NAND2_X1 U1714 ( .A1(n2165), .A2(n2166), .ZN(n2164) );
XOR2_X1 U1715 ( .A(n2167), .B(KEYINPUT38), .Z(n2163) );
NAND2_X1 U1716 ( .A1(n2168), .A2(n2169), .ZN(n2167) );
XNOR2_X1 U1717 ( .A(KEYINPUT61), .B(n2170), .ZN(n2168) );
INV_X1 U1718 ( .A(n2171), .ZN(n2137) );
NAND2_X1 U1719 ( .A1(n2172), .A2(n2171), .ZN(n2160) );
NAND2_X1 U1720 ( .A1(n2173), .A2(n2174), .ZN(n2171) );
NAND2_X1 U1721 ( .A1(n2175), .A2(n2176), .ZN(n2174) );
NAND2_X1 U1722 ( .A1(n2177), .A2(n2178), .ZN(n2175) );
NAND2_X1 U1723 ( .A1(n2179), .A2(n2180), .ZN(n2173) );
NAND2_X1 U1724 ( .A1(n2136), .A2(n2133), .ZN(n2172) );
NAND2_X1 U1725 ( .A1(n2166), .A2(n2170), .ZN(n2133) );
NAND2_X1 U1726 ( .A1(n2165), .A2(n2169), .ZN(n2136) );
INV_X1 U1727 ( .A(n2166), .ZN(n2169) );
NAND2_X1 U1728 ( .A1(n2181), .A2(n2182), .ZN(n2166) );
NAND2_X1 U1729 ( .A1(RESTART), .A2(n1886), .ZN(n2182) );
NAND2_X1 U1730 ( .A1(n2183), .A2(n2087), .ZN(n2181) );
INV_X1 U1731 ( .A(n2170), .ZN(n2165) );
NAND2_X1 U1732 ( .A1(n2184), .A2(n2185), .ZN(n2170) );
NAND2_X1 U1733 ( .A1(RESTART), .A2(n1904), .ZN(n2185) );
NAND2_X1 U1734 ( .A1(n1870), .A2(n2087), .ZN(n2184) );
NAND2_X1 U1735 ( .A1(n2024), .A2(RLAST_REG_3__SCAN_IN), .ZN(n2147) );
NAND2_X1 U1736 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1797), .ZN(n2146) );
NAND4_X1 U1737 ( .A1(n2186), .A2(n2187), .A3(n2188), .A4(n2189), .ZN(U283));
NOR3_X1 U1738 ( .A1(n2190), .A2(n2191), .A3(n2192), .ZN(n2189) );
NOR3_X1 U1739 ( .A1(n2023), .A2(n2117), .A3(n2193), .ZN(n2192) );
NOR2_X1 U1740 ( .A1(n2194), .A2(n2195), .ZN(n2193) );
AND2_X1 U1741 ( .A1(n2196), .A2(n2197), .ZN(n2194) );
AND3_X1 U1742 ( .A1(n2195), .A2(n2196), .A3(n2197), .ZN(n2117) );
NAND2_X1 U1743 ( .A1(n2120), .A2(n2198), .ZN(n2195) );
NAND2_X1 U1744 ( .A1(n2199), .A2(n2200), .ZN(n2120) );
NOR3_X1 U1745 ( .A1(n2018), .A2(n2106), .A3(n2201), .ZN(n2191) );
NOR2_X1 U1746 ( .A1(n2202), .A2(n2203), .ZN(n2201) );
INV_X1 U1747 ( .A(n2156), .ZN(n2106) );
NAND2_X1 U1748 ( .A1(n2202), .A2(n2203), .ZN(n2156) );
NAND2_X1 U1749 ( .A1(n2111), .A2(n2198), .ZN(n2203) );
NAND2_X1 U1750 ( .A1(n2204), .A2(n2205), .ZN(n2198) );
NAND2_X1 U1751 ( .A1(n2206), .A2(n2200), .ZN(n2111) );
XNOR2_X1 U1752 ( .A(n2199), .B(KEYINPUT54), .ZN(n2206) );
NOR2_X1 U1753 ( .A1(n2200), .A2(n2070), .ZN(n2190) );
INV_X1 U1754 ( .A(n2204), .ZN(n2200) );
NAND2_X1 U1755 ( .A1(n2207), .A2(n2208), .ZN(n2204) );
NAND2_X1 U1756 ( .A1(n2209), .A2(n2210), .ZN(n2208) );
NAND2_X1 U1757 ( .A1(n2211), .A2(n2212), .ZN(n2210) );
NAND2_X1 U1758 ( .A1(KEYINPUT57), .A2(n2213), .ZN(n2212) );
XNOR2_X1 U1759 ( .A(n2177), .B(n2214), .ZN(n2211) );
OR2_X1 U1760 ( .A1(KEYINPUT7), .A2(n2179), .ZN(n2214) );
INV_X1 U1761 ( .A(n2176), .ZN(n2209) );
NAND3_X1 U1762 ( .A1(n2213), .A2(n2215), .A3(n2176), .ZN(n2207) );
NAND2_X1 U1763 ( .A1(n2216), .A2(n2217), .ZN(n2176) );
NAND2_X1 U1764 ( .A1(n2218), .A2(n2219), .ZN(n2217) );
NAND2_X1 U1765 ( .A1(n2220), .A2(n2221), .ZN(n2219) );
INV_X1 U1766 ( .A(n2222), .ZN(n2221) );
XNOR2_X1 U1767 ( .A(KEYINPUT43), .B(n2223), .ZN(n2220) );
NAND2_X1 U1768 ( .A1(n2223), .A2(n2222), .ZN(n2216) );
INV_X1 U1769 ( .A(KEYINPUT57), .ZN(n2215) );
NAND2_X1 U1770 ( .A1(n2224), .A2(n2225), .ZN(n2213) );
NAND2_X1 U1771 ( .A1(n2179), .A2(n2177), .ZN(n2225) );
INV_X1 U1772 ( .A(n2180), .ZN(n2177) );
XOR2_X1 U1773 ( .A(KEYINPUT40), .B(n2226), .Z(n2224) );
NOR2_X1 U1774 ( .A1(n2179), .A2(n2227), .ZN(n2226) );
XNOR2_X1 U1775 ( .A(KEYINPUT7), .B(n2180), .ZN(n2227) );
NAND3_X1 U1776 ( .A1(n2228), .A2(n2229), .A3(n2230), .ZN(n2180) );
NAND2_X1 U1777 ( .A1(n2231), .A2(n1874), .ZN(n2230) );
NAND2_X1 U1778 ( .A1(REG4_REG_3__SCAN_IN), .A2(n2087), .ZN(n2231) );
OR2_X1 U1779 ( .A1(n2087), .A2(KEYINPUT25), .ZN(n2229) );
NAND3_X1 U1780 ( .A1(n2157), .A2(n2087), .A3(KEYINPUT25), .ZN(n2228) );
INV_X1 U1781 ( .A(n2178), .ZN(n2179) );
NAND3_X1 U1782 ( .A1(n2232), .A2(n2233), .A3(n2234), .ZN(n2178) );
NAND2_X1 U1783 ( .A1(KEYINPUT35), .A2(n1916), .ZN(n2234) );
NAND3_X1 U1784 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n2235), .A3(RESTART), .ZN(n2233) );
NAND2_X1 U1785 ( .A1(n2236), .A2(n2087), .ZN(n2232) );
NAND2_X1 U1786 ( .A1(n2235), .A2(n1885), .ZN(n2236) );
INV_X1 U1787 ( .A(KEYINPUT35), .ZN(n2235) );
NAND2_X1 U1788 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1797), .ZN(n2188) );
NAND2_X1 U1789 ( .A1(n2015), .A2(REG4_REG_2__SCAN_IN), .ZN(n2187) );
NAND2_X1 U1790 ( .A1(n2024), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2186) );
NAND4_X1 U1791 ( .A1(n2237), .A2(n2238), .A3(n2239), .A4(n2240), .ZN(U282));
NOR3_X1 U1792 ( .A1(n2241), .A2(n2242), .A3(n2243), .ZN(n2240) );
NOR2_X1 U1793 ( .A1(n2244), .A2(n2018), .ZN(n2243) );
INV_X1 U1794 ( .A(n2033), .ZN(n2018) );
NOR3_X1 U1795 ( .A1(n2245), .A2(n2246), .A3(n2247), .ZN(n2244) );
AND3_X1 U1796 ( .A1(n2248), .A2(n2249), .A3(KEYINPUT15), .ZN(n2247) );
NOR2_X1 U1797 ( .A1(n2248), .A2(n2250), .ZN(n2246) );
NOR2_X1 U1798 ( .A1(n2251), .A2(n2252), .ZN(n2250) );
NOR2_X1 U1799 ( .A1(KEYINPUT53), .A2(n2249), .ZN(n2252) );
NOR2_X1 U1800 ( .A1(KEYINPUT15), .A2(n2253), .ZN(n2251) );
INV_X1 U1801 ( .A(n2254), .ZN(n2248) );
AND2_X1 U1802 ( .A1(n2202), .A2(KEYINPUT53), .ZN(n2245) );
NOR2_X1 U1803 ( .A1(n2254), .A2(n2249), .ZN(n2202) );
INV_X1 U1804 ( .A(n2253), .ZN(n2249) );
NAND2_X1 U1805 ( .A1(n2255), .A2(n2205), .ZN(n2253) );
NOR2_X1 U1806 ( .A1(n2023), .A2(n2256), .ZN(n2242) );
XNOR2_X1 U1807 ( .A(n2196), .B(n2197), .ZN(n2256) );
NAND2_X1 U1808 ( .A1(n2257), .A2(n2205), .ZN(n2196) );
INV_X1 U1809 ( .A(n2199), .ZN(n2205) );
NOR3_X1 U1810 ( .A1(n2258), .A2(n2259), .A3(n2260), .ZN(n2199) );
XOR2_X1 U1811 ( .A(n2255), .B(KEYINPUT36), .Z(n2257) );
NAND2_X1 U1812 ( .A1(n2260), .A2(n2261), .ZN(n2255) );
NAND2_X1 U1813 ( .A1(n2262), .A2(n2263), .ZN(n2261) );
AND2_X1 U1814 ( .A1(n2260), .A2(n2123), .ZN(n2241) );
NAND2_X1 U1815 ( .A1(n2264), .A2(n2265), .ZN(n2260) );
NAND2_X1 U1816 ( .A1(n2266), .A2(n2267), .ZN(n2265) );
NAND2_X1 U1817 ( .A1(n2222), .A2(n2268), .ZN(n2267) );
XNOR2_X1 U1818 ( .A(n2269), .B(n2270), .ZN(n2266) );
NAND3_X1 U1819 ( .A1(n2271), .A2(n2272), .A3(n2222), .ZN(n2264) );
NAND2_X1 U1820 ( .A1(n2273), .A2(n2274), .ZN(n2222) );
NAND2_X1 U1821 ( .A1(n2275), .A2(n2276), .ZN(n2274) );
NAND2_X1 U1822 ( .A1(n2277), .A2(n2278), .ZN(n2273) );
NAND2_X1 U1823 ( .A1(n2218), .A2(n2279), .ZN(n2272) );
NAND2_X1 U1824 ( .A1(n2269), .A2(n2268), .ZN(n2279) );
INV_X1 U1825 ( .A(KEYINPUT63), .ZN(n2268) );
NAND2_X1 U1826 ( .A1(n2270), .A2(n2269), .ZN(n2271) );
INV_X1 U1827 ( .A(n2223), .ZN(n2269) );
NAND2_X1 U1828 ( .A1(n2280), .A2(n2281), .ZN(n2223) );
NAND2_X1 U1829 ( .A1(n1878), .A2(n2087), .ZN(n2281) );
NAND2_X1 U1830 ( .A1(n2282), .A2(RESTART), .ZN(n2280) );
XNOR2_X1 U1831 ( .A(n1911), .B(KEYINPUT55), .ZN(n2282) );
INV_X1 U1832 ( .A(n2218), .ZN(n2270) );
NAND2_X1 U1833 ( .A1(n2283), .A2(n2284), .ZN(n2218) );
NAND2_X1 U1834 ( .A1(RESTART), .A2(n1884), .ZN(n2284) );
NAND2_X1 U1835 ( .A1(n2285), .A2(n2087), .ZN(n2283) );
NAND2_X1 U1836 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1797), .ZN(n2239) );
NAND2_X1 U1837 ( .A1(n2015), .A2(REG4_REG_1__SCAN_IN), .ZN(n2238) );
NAND2_X1 U1838 ( .A1(n2024), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2237) );
NAND4_X1 U1839 ( .A1(n2286), .A2(n2287), .A3(n2288), .A4(n2289), .ZN(U281));
NOR3_X1 U1840 ( .A1(n2290), .A2(n2291), .A3(n2292), .ZN(n2289) );
NOR2_X1 U1841 ( .A1(n2023), .A2(n2197), .ZN(n2292) );
XOR2_X1 U1842 ( .A(n2259), .B(n2293), .Z(n2197) );
NOR2_X1 U1843 ( .A1(KEYINPUT18), .A2(n2258), .ZN(n2293) );
NAND3_X1 U1844 ( .A1(RESTART), .A2(n2294), .A3(n2295), .ZN(n2023) );
XOR2_X1 U1845 ( .A(KEYINPUT24), .B(n2296), .Z(n2294) );
NOR2_X1 U1846 ( .A1(n2297), .A2(n2032), .ZN(n2291) );
INV_X1 U1847 ( .A(n2015), .ZN(n2032) );
NOR2_X1 U1848 ( .A1(n2298), .A2(n2299), .ZN(n2015) );
AND2_X1 U1849 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n2024), .ZN(n2290) );
INV_X1 U1850 ( .A(n2121), .ZN(n2024) );
NAND3_X1 U1851 ( .A1(n1939), .A2(n2087), .A3(n2296), .ZN(n2121) );
INV_X1 U1852 ( .A(ENABLE), .ZN(n1939) );
NAND2_X1 U1853 ( .A1(n2123), .A2(n2258), .ZN(n2288) );
INV_X1 U1854 ( .A(n2070), .ZN(n2123) );
NAND3_X1 U1855 ( .A1(n2300), .A2(n2301), .A3(n2296), .ZN(n2070) );
NAND2_X1 U1856 ( .A1(n2302), .A2(n2087), .ZN(n2301) );
NAND3_X1 U1857 ( .A1(n2303), .A2(n2298), .A3(ENABLE), .ZN(n2302) );
INV_X1 U1858 ( .A(AVERAGE), .ZN(n2298) );
NAND2_X1 U1859 ( .A1(n2295), .A2(RESTART), .ZN(n2300) );
XOR2_X1 U1860 ( .A(n2304), .B(KEYINPUT60), .Z(n2295) );
NAND2_X1 U1861 ( .A1(n2305), .A2(n2306), .ZN(n2304) );
NAND2_X1 U1862 ( .A1(n2307), .A2(n1889), .ZN(n2306) );
INV_X1 U1863 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1889) );
OR2_X1 U1864 ( .A1(n2308), .A2(n1893), .ZN(n2307) );
NAND2_X1 U1865 ( .A1(n2308), .A2(n1893), .ZN(n2305) );
INV_X1 U1866 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1893) );
NAND2_X1 U1867 ( .A1(n2309), .A2(n2310), .ZN(n2308) );
NAND2_X1 U1868 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n2311), .ZN(n2310) );
NAND2_X1 U1869 ( .A1(n2312), .A2(n1888), .ZN(n2311) );
XOR2_X1 U1870 ( .A(n2313), .B(KEYINPUT21), .Z(n2312) );
OR2_X1 U1871 ( .A1(n2313), .A2(n1888), .ZN(n2309) );
INV_X1 U1872 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1888) );
NAND2_X1 U1873 ( .A1(n2314), .A2(n2315), .ZN(n2313) );
NAND2_X1 U1874 ( .A1(n2316), .A2(n1866), .ZN(n2315) );
INV_X1 U1875 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1866) );
NAND2_X1 U1876 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n2317), .ZN(n2316) );
OR2_X1 U1877 ( .A1(n2317), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2314) );
XNOR2_X1 U1878 ( .A(n2318), .B(KEYINPUT34), .ZN(n2317) );
NAND2_X1 U1879 ( .A1(n2319), .A2(n2320), .ZN(n2318) );
NAND2_X1 U1880 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2320) );
NAND3_X1 U1881 ( .A1(n2321), .A2(n2322), .A3(n2323), .ZN(n2319) );
NAND2_X1 U1882 ( .A1(n1904), .A2(n1886), .ZN(n2323) );
INV_X1 U1883 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1886) );
INV_X1 U1884 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1904) );
NAND3_X1 U1885 ( .A1(n2324), .A2(n2325), .A3(n2326), .ZN(n2322) );
NAND2_X1 U1886 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2326) );
NAND3_X1 U1887 ( .A1(n2327), .A2(n2328), .A3(n2329), .ZN(n2325) );
NAND2_X1 U1888 ( .A1(n1911), .A2(n1884), .ZN(n2329) );
INV_X1 U1889 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1884) );
INV_X1 U1890 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1911) );
NAND2_X1 U1891 ( .A1(n2330), .A2(n2331), .ZN(n2328) );
NAND2_X1 U1892 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n2332), .ZN(n2331) );
XNOR2_X1 U1893 ( .A(n1915), .B(KEYINPUT13), .ZN(n2332) );
NAND2_X1 U1894 ( .A1(n1915), .A2(n2333), .ZN(n2327) );
INV_X1 U1895 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1915) );
NAND2_X1 U1896 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2324) );
NAND2_X1 U1897 ( .A1(n1916), .A2(n1874), .ZN(n2321) );
INV_X1 U1898 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1874) );
INV_X1 U1899 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1916) );
NAND2_X1 U1900 ( .A1(n2033), .A2(n2334), .ZN(n2287) );
XNOR2_X1 U1901 ( .A(KEYINPUT46), .B(n2254), .ZN(n2334) );
NAND2_X1 U1902 ( .A1(n2335), .A2(n2336), .ZN(n2254) );
NAND2_X1 U1903 ( .A1(n2258), .A2(n2263), .ZN(n2336) );
XOR2_X1 U1904 ( .A(n2337), .B(KEYINPUT0), .Z(n2335) );
NAND2_X1 U1905 ( .A1(n2259), .A2(n2262), .ZN(n2337) );
INV_X1 U1906 ( .A(n2258), .ZN(n2262) );
NAND3_X1 U1907 ( .A1(n2338), .A2(n2339), .A3(n2340), .ZN(n2258) );
NAND2_X1 U1908 ( .A1(n2278), .A2(n2341), .ZN(n2340) );
NAND2_X1 U1909 ( .A1(n2342), .A2(n2343), .ZN(n2341) );
NAND2_X1 U1910 ( .A1(n2344), .A2(n2345), .ZN(n2343) );
XNOR2_X1 U1911 ( .A(n2346), .B(KEYINPUT37), .ZN(n2345) );
NAND2_X1 U1912 ( .A1(n2346), .A2(n2277), .ZN(n2342) );
NAND3_X1 U1913 ( .A1(n2277), .A2(n2347), .A3(n2275), .ZN(n2339) );
XOR2_X1 U1914 ( .A(n2344), .B(KEYINPUT12), .Z(n2277) );
NAND2_X1 U1915 ( .A1(n2346), .A2(n2348), .ZN(n2338) );
XOR2_X1 U1916 ( .A(n2276), .B(KEYINPUT23), .Z(n2348) );
NAND2_X1 U1917 ( .A1(n2344), .A2(n2347), .ZN(n2276) );
INV_X1 U1918 ( .A(n2278), .ZN(n2347) );
AND2_X1 U1919 ( .A1(n2349), .A2(n2350), .ZN(n2344) );
NAND2_X1 U1920 ( .A1(n1880), .A2(n2087), .ZN(n2350) );
NAND2_X1 U1921 ( .A1(n2351), .A2(RESTART), .ZN(n2349) );
XNOR2_X1 U1922 ( .A(RMAX_REG_1__SCAN_IN), .B(KEYINPUT58), .ZN(n2351) );
INV_X1 U1923 ( .A(n2275), .ZN(n2346) );
NAND2_X1 U1924 ( .A1(n2352), .A2(n2353), .ZN(n2275) );
NAND2_X1 U1925 ( .A1(RESTART), .A2(n2333), .ZN(n2353) );
INV_X1 U1926 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n2333) );
NAND2_X1 U1927 ( .A1(n2354), .A2(n2087), .ZN(n2352) );
INV_X1 U1928 ( .A(n2263), .ZN(n2259) );
NAND3_X1 U1929 ( .A1(n2355), .A2(n2356), .A3(n2278), .ZN(n2263) );
NAND2_X1 U1930 ( .A1(n2357), .A2(n2358), .ZN(n2278) );
NAND2_X1 U1931 ( .A1(RESTART), .A2(n2330), .ZN(n2358) );
NAND2_X1 U1932 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2330) );
NAND2_X1 U1933 ( .A1(n2359), .A2(n2087), .ZN(n2357) );
NAND2_X1 U1934 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2359) );
NAND3_X1 U1935 ( .A1(n1879), .A2(n2297), .A3(n2087), .ZN(n2356) );
INV_X1 U1936 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2297) );
OR3_X1 U1937 ( .A1(RMAX_REG_0__SCAN_IN), .A2(RMIN_REG_0__SCAN_IN), .A3(n2087), .ZN(n2355) );
NOR3_X1 U1938 ( .A1(n2303), .A2(AVERAGE), .A3(n2299), .ZN(n2033) );
NAND3_X1 U1939 ( .A1(n2296), .A2(n2087), .A3(ENABLE), .ZN(n2299) );
INV_X1 U1940 ( .A(RESTART), .ZN(n2087) );
NOR2_X1 U1941 ( .A1(n1940), .A2(n1797), .ZN(n2296) );
NAND2_X1 U1942 ( .A1(n2360), .A2(n2361), .ZN(n2303) );
NAND2_X1 U1943 ( .A1(n2362), .A2(n2363), .ZN(n2361) );
INV_X1 U1944 ( .A(REG4_REG_7__SCAN_IN), .ZN(n2363) );
OR2_X1 U1945 ( .A1(n2364), .A2(n1858), .ZN(n2362) );
NAND2_X1 U1946 ( .A1(n2364), .A2(n1858), .ZN(n2360) );
INV_X1 U1947 ( .A(DATA_IN_7_), .ZN(n1858) );
NAND2_X1 U1948 ( .A1(n2365), .A2(n2366), .ZN(n2364) );
NAND2_X1 U1949 ( .A1(REG4_REG_6__SCAN_IN), .A2(n2367), .ZN(n2366) );
NAND2_X1 U1950 ( .A1(n2368), .A2(n2369), .ZN(n2367) );
XNOR2_X1 U1951 ( .A(KEYINPUT8), .B(n1862), .ZN(n2368) );
OR2_X1 U1952 ( .A1(n2369), .A2(n1862), .ZN(n2365) );
INV_X1 U1953 ( .A(DATA_IN_6_), .ZN(n1862) );
NAND2_X1 U1954 ( .A1(n2370), .A2(n2371), .ZN(n2369) );
NAND3_X1 U1955 ( .A1(n2372), .A2(n2373), .A3(n2374), .ZN(n2371) );
NAND2_X1 U1956 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2374) );
NAND3_X1 U1957 ( .A1(n2375), .A2(n2376), .A3(n2377), .ZN(n2373) );
NAND2_X1 U1958 ( .A1(n1870), .A2(n2183), .ZN(n2377) );
INV_X1 U1959 ( .A(REG4_REG_4__SCAN_IN), .ZN(n2183) );
INV_X1 U1960 ( .A(DATA_IN_4_), .ZN(n1870) );
NAND3_X1 U1961 ( .A1(n2378), .A2(n2379), .A3(n2380), .ZN(n2376) );
NAND2_X1 U1962 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2380) );
NAND3_X1 U1963 ( .A1(n2381), .A2(n2382), .A3(n2383), .ZN(n2379) );
NAND2_X1 U1964 ( .A1(n1878), .A2(n2285), .ZN(n2383) );
INV_X1 U1965 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2285) );
INV_X1 U1966 ( .A(DATA_IN_2_), .ZN(n1878) );
NAND2_X1 U1967 ( .A1(n2384), .A2(n2354), .ZN(n2382) );
INV_X1 U1968 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2354) );
OR2_X1 U1969 ( .A1(n2385), .A2(n1880), .ZN(n2384) );
NAND2_X1 U1970 ( .A1(n2385), .A2(n1880), .ZN(n2381) );
INV_X1 U1971 ( .A(DATA_IN_1_), .ZN(n1880) );
NAND2_X1 U1972 ( .A1(REG4_REG_0__SCAN_IN), .A2(n2386), .ZN(n2385) );
XNOR2_X1 U1973 ( .A(KEYINPUT50), .B(n1879), .ZN(n2386) );
INV_X1 U1974 ( .A(DATA_IN_0_), .ZN(n1879) );
NAND2_X1 U1975 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2378) );
NAND2_X1 U1976 ( .A1(n1885), .A2(n2157), .ZN(n2375) );
INV_X1 U1977 ( .A(REG4_REG_3__SCAN_IN), .ZN(n2157) );
INV_X1 U1978 ( .A(DATA_IN_3_), .ZN(n1885) );
NAND2_X1 U1979 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2372) );
NAND2_X1 U1980 ( .A1(n2145), .A2(n1887), .ZN(n2370) );
INV_X1 U1981 ( .A(DATA_IN_5_), .ZN(n1887) );
INV_X1 U1982 ( .A(REG4_REG_5__SCAN_IN), .ZN(n2145) );
NAND2_X1 U1983 ( .A1(n2387), .A2(n1797), .ZN(n2286) );
XNOR2_X1 U1984 ( .A(KEYINPUT2), .B(DATA_OUT_REG_0__SCAN_IN), .ZN(n2387) );
INV_X1 U1985 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1940) );
NOR2_X1 U1986 ( .A1(n1819), .A2(STATO_REG_1__SCAN_IN), .ZN(n2388) );
INV_X1 U1987 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1819) );
endmodule


