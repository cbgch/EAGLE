//Key = 0000110101001110010101000101001000010000101101000001100010001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290;

XOR2_X1 U711 ( .A(G107), .B(n970), .Z(G9) );
NAND3_X1 U712 ( .A1(n971), .A2(n972), .A3(n973), .ZN(G75) );
NAND2_X1 U713 ( .A1(G952), .A2(n974), .ZN(n973) );
NAND3_X1 U714 ( .A1(n975), .A2(n976), .A3(n977), .ZN(n974) );
NAND2_X1 U715 ( .A1(n978), .A2(n979), .ZN(n976) );
NAND2_X1 U716 ( .A1(n980), .A2(n981), .ZN(n979) );
NAND4_X1 U717 ( .A1(n982), .A2(n983), .A3(n984), .A4(n985), .ZN(n981) );
NOR2_X1 U718 ( .A1(n986), .A2(n987), .ZN(n985) );
NAND2_X1 U719 ( .A1(n988), .A2(n989), .ZN(n984) );
NAND3_X1 U720 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n983) );
NAND2_X1 U721 ( .A1(n993), .A2(n994), .ZN(n992) );
NAND2_X1 U722 ( .A1(n989), .A2(n995), .ZN(n994) );
NAND2_X1 U723 ( .A1(n996), .A2(n997), .ZN(n982) );
NAND4_X1 U724 ( .A1(n998), .A2(n999), .A3(n1000), .A4(n1001), .ZN(n980) );
NOR2_X1 U725 ( .A1(n997), .A2(n996), .ZN(n1001) );
NAND2_X1 U726 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NAND4_X1 U727 ( .A1(n1004), .A2(n1005), .A3(n1003), .A4(n1006), .ZN(n999) );
NAND2_X1 U728 ( .A1(n987), .A2(n986), .ZN(n998) );
XOR2_X1 U729 ( .A(n1007), .B(KEYINPUT38), .Z(n978) );
NAND4_X1 U730 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n971) );
NOR4_X1 U731 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1011) );
XOR2_X1 U732 ( .A(n1016), .B(n1017), .Z(n1013) );
NOR2_X1 U733 ( .A1(KEYINPUT3), .A2(n1018), .ZN(n1017) );
XOR2_X1 U734 ( .A(KEYINPUT34), .B(G478), .Z(n1018) );
XOR2_X1 U735 ( .A(n1019), .B(n1020), .Z(n1010) );
NAND2_X1 U736 ( .A1(KEYINPUT43), .A2(n1021), .ZN(n1019) );
INV_X1 U737 ( .A(n1022), .ZN(n1021) );
INV_X1 U738 ( .A(n996), .ZN(n1009) );
XNOR2_X1 U739 ( .A(n1002), .B(KEYINPUT26), .ZN(n1008) );
XOR2_X1 U740 ( .A(n1023), .B(n1024), .Z(G72) );
XOR2_X1 U741 ( .A(n1025), .B(n1026), .Z(n1024) );
NOR2_X1 U742 ( .A1(n1027), .A2(n972), .ZN(n1026) );
NOR2_X1 U743 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U744 ( .A1(n1030), .A2(n1031), .ZN(n1025) );
NAND2_X1 U745 ( .A1(n1032), .A2(n1029), .ZN(n1031) );
XNOR2_X1 U746 ( .A(KEYINPUT18), .B(n972), .ZN(n1032) );
XOR2_X1 U747 ( .A(n1033), .B(n1034), .Z(n1030) );
XOR2_X1 U748 ( .A(n1035), .B(n1036), .Z(n1034) );
XNOR2_X1 U749 ( .A(n1037), .B(KEYINPUT17), .ZN(n1033) );
NAND2_X1 U750 ( .A1(n1038), .A2(KEYINPUT4), .ZN(n1037) );
XNOR2_X1 U751 ( .A(n1039), .B(KEYINPUT5), .ZN(n1038) );
NAND2_X1 U752 ( .A1(n972), .A2(n1040), .ZN(n1023) );
XOR2_X1 U753 ( .A(n1041), .B(n1042), .Z(G69) );
NOR2_X1 U754 ( .A1(n1043), .A2(n972), .ZN(n1042) );
AND2_X1 U755 ( .A1(G224), .A2(G898), .ZN(n1043) );
NAND2_X1 U756 ( .A1(n1044), .A2(n1045), .ZN(n1041) );
NAND2_X1 U757 ( .A1(n1046), .A2(n972), .ZN(n1045) );
XOR2_X1 U758 ( .A(n975), .B(n1047), .Z(n1046) );
OR3_X1 U759 ( .A1(n1048), .A2(n1047), .A3(n972), .ZN(n1044) );
NOR2_X1 U760 ( .A1(n1049), .A2(n1050), .ZN(G66) );
XOR2_X1 U761 ( .A(n1051), .B(n1052), .Z(n1050) );
NOR3_X1 U762 ( .A1(n1053), .A2(KEYINPUT24), .A3(n1022), .ZN(n1052) );
NOR2_X1 U763 ( .A1(n1049), .A2(n1054), .ZN(G63) );
XOR2_X1 U764 ( .A(n1055), .B(n1056), .Z(n1054) );
AND2_X1 U765 ( .A1(G478), .A2(n1057), .ZN(n1055) );
NOR3_X1 U766 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(G60) );
AND3_X1 U767 ( .A1(KEYINPUT29), .A2(G953), .A3(G952), .ZN(n1060) );
NOR2_X1 U768 ( .A1(KEYINPUT29), .A2(n1061), .ZN(n1059) );
INV_X1 U769 ( .A(n1049), .ZN(n1061) );
XOR2_X1 U770 ( .A(n1062), .B(n1063), .Z(n1058) );
XOR2_X1 U771 ( .A(KEYINPUT61), .B(n1064), .Z(n1063) );
AND2_X1 U772 ( .A1(G475), .A2(n1057), .ZN(n1064) );
XOR2_X1 U773 ( .A(n1065), .B(n1066), .Z(G6) );
NOR2_X1 U774 ( .A1(n989), .A2(n1067), .ZN(n1066) );
NOR2_X1 U775 ( .A1(n1068), .A2(n1069), .ZN(n1065) );
XNOR2_X1 U776 ( .A(KEYINPUT42), .B(KEYINPUT15), .ZN(n1068) );
NOR2_X1 U777 ( .A1(n1049), .A2(n1070), .ZN(G57) );
XOR2_X1 U778 ( .A(n1071), .B(n1072), .Z(n1070) );
NAND2_X1 U779 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND3_X1 U780 ( .A1(G210), .A2(n1075), .A3(G101), .ZN(n1074) );
XOR2_X1 U781 ( .A(n1076), .B(KEYINPUT6), .Z(n1073) );
NAND2_X1 U782 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U783 ( .A1(G210), .A2(n1075), .ZN(n1078) );
NAND3_X1 U784 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1071) );
NAND2_X1 U785 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
OR3_X1 U786 ( .A1(n1083), .A2(n1082), .A3(KEYINPUT11), .ZN(n1080) );
XNOR2_X1 U787 ( .A(n1084), .B(n1085), .ZN(n1082) );
NAND2_X1 U788 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
OR2_X1 U789 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U790 ( .A(n1090), .B(KEYINPUT28), .Z(n1086) );
NAND2_X1 U791 ( .A1(n1089), .A2(n1088), .ZN(n1090) );
NAND2_X1 U792 ( .A1(KEYINPUT25), .A2(n1091), .ZN(n1083) );
NAND2_X1 U793 ( .A1(n1057), .A2(G472), .ZN(n1091) );
NAND3_X1 U794 ( .A1(n1057), .A2(G472), .A3(KEYINPUT11), .ZN(n1079) );
NOR2_X1 U795 ( .A1(n1049), .A2(n1092), .ZN(G54) );
XOR2_X1 U796 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U797 ( .A(n1088), .B(n1095), .Z(n1094) );
XOR2_X1 U798 ( .A(n1096), .B(n1097), .Z(n1093) );
XOR2_X1 U799 ( .A(n1098), .B(n1099), .Z(n1097) );
AND2_X1 U800 ( .A1(G469), .A2(n1057), .ZN(n1099) );
INV_X1 U801 ( .A(n1053), .ZN(n1057) );
NOR2_X1 U802 ( .A1(n1100), .A2(n1101), .ZN(G51) );
XOR2_X1 U803 ( .A(KEYINPUT32), .B(n1049), .Z(n1101) );
NOR2_X1 U804 ( .A1(n972), .A2(G952), .ZN(n1049) );
XOR2_X1 U805 ( .A(n1102), .B(n1103), .Z(n1100) );
XNOR2_X1 U806 ( .A(n1104), .B(n1039), .ZN(n1103) );
XOR2_X1 U807 ( .A(n1105), .B(n1106), .Z(n1102) );
NOR2_X1 U808 ( .A1(G125), .A2(KEYINPUT50), .ZN(n1106) );
NOR3_X1 U809 ( .A1(n1053), .A2(n1107), .A3(n1108), .ZN(n1105) );
NAND2_X1 U810 ( .A1(n1109), .A2(n1110), .ZN(n1053) );
NAND2_X1 U811 ( .A1(n977), .A2(n1111), .ZN(n1110) );
XOR2_X1 U812 ( .A(KEYINPUT58), .B(n975), .Z(n1111) );
AND2_X1 U813 ( .A1(n1112), .A2(n1113), .ZN(n975) );
NOR4_X1 U814 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n970), .ZN(n1113) );
AND3_X1 U815 ( .A1(n993), .A2(n1117), .A3(n1118), .ZN(n970) );
NOR2_X1 U816 ( .A1(n1119), .A2(n989), .ZN(n1116) );
XOR2_X1 U817 ( .A(n1067), .B(KEYINPUT44), .Z(n1119) );
NAND4_X1 U818 ( .A1(n1120), .A2(n993), .A3(n1121), .A4(n1122), .ZN(n1067) );
INV_X1 U819 ( .A(n1123), .ZN(n1114) );
NOR4_X1 U820 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1112) );
NOR4_X1 U821 ( .A1(n1128), .A2(n1129), .A3(n987), .A4(n1130), .ZN(n1127) );
INV_X1 U822 ( .A(n1131), .ZN(n987) );
NOR2_X1 U823 ( .A1(KEYINPUT21), .A2(n1132), .ZN(n1129) );
NOR2_X1 U824 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U825 ( .A1(n1135), .A2(n1136), .ZN(n1128) );
INV_X1 U826 ( .A(KEYINPUT21), .ZN(n1136) );
INV_X1 U827 ( .A(n1040), .ZN(n977) );
NAND4_X1 U828 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1040) );
NOR4_X1 U829 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1140) );
INV_X1 U830 ( .A(n1145), .ZN(n1143) );
NOR3_X1 U831 ( .A1(n1146), .A2(n1004), .A3(n1147), .ZN(n1142) );
XNOR2_X1 U832 ( .A(KEYINPUT47), .B(n1148), .ZN(n1146) );
NOR4_X1 U833 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1139) );
AND4_X1 U834 ( .A1(KEYINPUT22), .A2(n1153), .A3(n1005), .A4(n1154), .ZN(n1152) );
NOR2_X1 U835 ( .A1(KEYINPUT22), .A2(n1155), .ZN(n1151) );
INV_X1 U836 ( .A(n1156), .ZN(n1155) );
NOR2_X1 U837 ( .A1(n1157), .A2(n1158), .ZN(n1150) );
INV_X1 U838 ( .A(KEYINPUT27), .ZN(n1157) );
NOR3_X1 U839 ( .A1(KEYINPUT27), .A2(n1159), .A3(n1160), .ZN(n1149) );
XNOR2_X1 U840 ( .A(KEYINPUT63), .B(n1161), .ZN(n1109) );
XNOR2_X1 U841 ( .A(G146), .B(n1162), .ZN(G48) );
NAND2_X1 U842 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NAND2_X1 U843 ( .A1(KEYINPUT60), .A2(n1137), .ZN(n1164) );
NAND2_X1 U844 ( .A1(KEYINPUT46), .A2(n1165), .ZN(n1163) );
INV_X1 U845 ( .A(n1137), .ZN(n1165) );
NAND2_X1 U846 ( .A1(n1166), .A2(n1120), .ZN(n1137) );
XNOR2_X1 U847 ( .A(G143), .B(n1158), .ZN(G45) );
OR2_X1 U848 ( .A1(n1160), .A2(n990), .ZN(n1158) );
NAND3_X1 U849 ( .A1(n1121), .A2(n1134), .A3(n1167), .ZN(n1160) );
NOR3_X1 U850 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1167) );
NAND3_X1 U851 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(G42) );
OR2_X1 U852 ( .A1(n1156), .A2(KEYINPUT35), .ZN(n1173) );
NAND3_X1 U853 ( .A1(KEYINPUT35), .A2(n1156), .A3(n1174), .ZN(n1172) );
NAND2_X1 U854 ( .A1(G140), .A2(n1175), .ZN(n1171) );
NAND2_X1 U855 ( .A1(n1176), .A2(KEYINPUT35), .ZN(n1175) );
XNOR2_X1 U856 ( .A(n1156), .B(KEYINPUT45), .ZN(n1176) );
NOR3_X1 U857 ( .A1(n1005), .A2(n1177), .A3(n991), .ZN(n1156) );
XOR2_X1 U858 ( .A(G137), .B(n1141), .Z(G39) );
NOR4_X1 U859 ( .A1(n986), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1141) );
XOR2_X1 U860 ( .A(n1138), .B(n1180), .Z(G36) );
XNOR2_X1 U861 ( .A(G134), .B(KEYINPUT49), .ZN(n1180) );
NAND3_X1 U862 ( .A1(n1154), .A2(n1118), .A3(n1159), .ZN(n1138) );
XNOR2_X1 U863 ( .A(n1181), .B(n1144), .ZN(G33) );
NOR2_X1 U864 ( .A1(n1130), .A2(n1177), .ZN(n1144) );
INV_X1 U865 ( .A(n1154), .ZN(n1177) );
NOR3_X1 U866 ( .A1(n1003), .A2(n1169), .A3(n996), .ZN(n1154) );
NAND2_X1 U867 ( .A1(n1182), .A2(n995), .ZN(n996) );
INV_X1 U868 ( .A(n1121), .ZN(n1003) );
XNOR2_X1 U869 ( .A(G128), .B(n1183), .ZN(G30) );
NAND2_X1 U870 ( .A1(n1166), .A2(n1118), .ZN(n1183) );
NOR2_X1 U871 ( .A1(n1147), .A2(n1169), .ZN(n1166) );
INV_X1 U872 ( .A(n1148), .ZN(n1169) );
NAND4_X1 U873 ( .A1(n1184), .A2(n1121), .A3(n1134), .A4(n1014), .ZN(n1147) );
XNOR2_X1 U874 ( .A(G101), .B(n1185), .ZN(G3) );
NAND2_X1 U875 ( .A1(KEYINPUT7), .A2(n1115), .ZN(n1185) );
AND3_X1 U876 ( .A1(n1186), .A2(n1117), .A3(n1159), .ZN(n1115) );
NAND2_X1 U877 ( .A1(n1187), .A2(n1188), .ZN(G27) );
OR2_X1 U878 ( .A1(n1145), .A2(G125), .ZN(n1188) );
XOR2_X1 U879 ( .A(n1189), .B(KEYINPUT54), .Z(n1187) );
NAND2_X1 U880 ( .A1(G125), .A2(n1145), .ZN(n1189) );
NAND4_X1 U881 ( .A1(n1134), .A2(n1148), .A3(n1131), .A4(n1190), .ZN(n1145) );
NOR2_X1 U882 ( .A1(n1005), .A2(n991), .ZN(n1190) );
INV_X1 U883 ( .A(n1153), .ZN(n991) );
INV_X1 U884 ( .A(n1120), .ZN(n1005) );
NAND2_X1 U885 ( .A1(n1191), .A2(n1192), .ZN(n1148) );
NAND4_X1 U886 ( .A1(G953), .A2(n1193), .A3(n1007), .A4(n1029), .ZN(n1192) );
INV_X1 U887 ( .A(G900), .ZN(n1029) );
XNOR2_X1 U888 ( .A(KEYINPUT20), .B(n1161), .ZN(n1193) );
INV_X1 U889 ( .A(n989), .ZN(n1134) );
XOR2_X1 U890 ( .A(G122), .B(n1194), .Z(G24) );
NOR2_X1 U891 ( .A1(KEYINPUT53), .A2(n1195), .ZN(n1194) );
INV_X1 U892 ( .A(n1126), .ZN(n1195) );
NOR4_X1 U893 ( .A1(n1196), .A2(n997), .A3(n1168), .A4(n1170), .ZN(n1126) );
INV_X1 U894 ( .A(n993), .ZN(n997) );
NOR2_X1 U895 ( .A1(n1014), .A2(n1184), .ZN(n993) );
XNOR2_X1 U896 ( .A(n1125), .B(n1197), .ZN(G21) );
NAND2_X1 U897 ( .A1(KEYINPUT40), .A2(G119), .ZN(n1197) );
NOR4_X1 U898 ( .A1(n1196), .A2(n986), .A3(n1178), .A4(n1179), .ZN(n1125) );
INV_X1 U899 ( .A(n1186), .ZN(n986) );
NAND2_X1 U900 ( .A1(n1198), .A2(n1199), .ZN(G18) );
OR2_X1 U901 ( .A1(n1200), .A2(n1124), .ZN(n1199) );
XOR2_X1 U902 ( .A(n1201), .B(KEYINPUT2), .Z(n1198) );
NAND2_X1 U903 ( .A1(n1124), .A2(n1200), .ZN(n1201) );
NOR3_X1 U904 ( .A1(n990), .A2(n1004), .A3(n1196), .ZN(n1124) );
INV_X1 U905 ( .A(n1118), .ZN(n1004) );
NOR2_X1 U906 ( .A1(n1015), .A2(n1168), .ZN(n1118) );
INV_X1 U907 ( .A(n1202), .ZN(n1168) );
INV_X1 U908 ( .A(n1159), .ZN(n990) );
XOR2_X1 U909 ( .A(G113), .B(n1203), .Z(G15) );
NOR2_X1 U910 ( .A1(n1130), .A2(n1196), .ZN(n1203) );
NAND2_X1 U911 ( .A1(n1131), .A2(n1135), .ZN(n1196) );
NOR2_X1 U912 ( .A1(n1002), .A2(n1012), .ZN(n1131) );
NAND2_X1 U913 ( .A1(n1159), .A2(n1120), .ZN(n1130) );
NOR2_X1 U914 ( .A1(n1202), .A2(n1170), .ZN(n1120) );
INV_X1 U915 ( .A(n1015), .ZN(n1170) );
NOR2_X1 U916 ( .A1(n1179), .A2(n1184), .ZN(n1159) );
INV_X1 U917 ( .A(n1178), .ZN(n1184) );
INV_X1 U918 ( .A(n1014), .ZN(n1179) );
XNOR2_X1 U919 ( .A(G110), .B(n1123), .ZN(G12) );
NAND3_X1 U920 ( .A1(n1186), .A2(n1117), .A3(n1153), .ZN(n1123) );
NOR2_X1 U921 ( .A1(n1178), .A2(n1014), .ZN(n1153) );
XNOR2_X1 U922 ( .A(n1204), .B(G472), .ZN(n1014) );
NAND2_X1 U923 ( .A1(n1205), .A2(n1161), .ZN(n1204) );
XOR2_X1 U924 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U925 ( .A(n1208), .B(n1209), .Z(n1207) );
XNOR2_X1 U926 ( .A(n1077), .B(n1210), .ZN(n1209) );
NOR2_X1 U927 ( .A1(KEYINPUT62), .A2(n1085), .ZN(n1210) );
NOR3_X1 U928 ( .A1(n1108), .A2(KEYINPUT23), .A3(n1211), .ZN(n1208) );
XNOR2_X1 U929 ( .A(n1088), .B(n1039), .ZN(n1206) );
XNOR2_X1 U930 ( .A(n1212), .B(n1020), .ZN(n1178) );
NOR2_X1 U931 ( .A1(n1051), .A2(G902), .ZN(n1020) );
XNOR2_X1 U932 ( .A(n1213), .B(n1214), .ZN(n1051) );
XOR2_X1 U933 ( .A(n1215), .B(n1216), .Z(n1214) );
NAND2_X1 U934 ( .A1(G221), .A2(n1217), .ZN(n1216) );
INV_X1 U935 ( .A(n1218), .ZN(n1217) );
NAND2_X1 U936 ( .A1(n1219), .A2(KEYINPUT30), .ZN(n1215) );
XOR2_X1 U937 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U938 ( .A(n1222), .B(n1223), .Z(n1221) );
XNOR2_X1 U939 ( .A(n1224), .B(n1225), .ZN(n1223) );
NOR2_X1 U940 ( .A1(G146), .A2(KEYINPUT37), .ZN(n1225) );
NAND2_X1 U941 ( .A1(KEYINPUT9), .A2(n1174), .ZN(n1224) );
NOR2_X1 U942 ( .A1(G119), .A2(KEYINPUT59), .ZN(n1222) );
XNOR2_X1 U943 ( .A(G110), .B(n1226), .ZN(n1220) );
XNOR2_X1 U944 ( .A(n1227), .B(G125), .ZN(n1226) );
NAND2_X1 U945 ( .A1(KEYINPUT14), .A2(n1022), .ZN(n1212) );
NAND2_X1 U946 ( .A1(G217), .A2(n1228), .ZN(n1022) );
AND2_X1 U947 ( .A1(n1121), .A2(n1135), .ZN(n1117) );
NOR2_X1 U948 ( .A1(n989), .A2(n1133), .ZN(n1135) );
INV_X1 U949 ( .A(n1122), .ZN(n1133) );
NAND2_X1 U950 ( .A1(n1191), .A2(n1229), .ZN(n1122) );
NAND4_X1 U951 ( .A1(n1048), .A2(G953), .A3(G902), .A4(n1007), .ZN(n1229) );
XNOR2_X1 U952 ( .A(G898), .B(KEYINPUT1), .ZN(n1048) );
NAND3_X1 U953 ( .A1(n1007), .A2(n972), .A3(G952), .ZN(n1191) );
NAND2_X1 U954 ( .A1(G237), .A2(G234), .ZN(n1007) );
NAND2_X1 U955 ( .A1(n1230), .A2(n995), .ZN(n989) );
OR2_X1 U956 ( .A1(n1231), .A2(n1107), .ZN(n995) );
XNOR2_X1 U957 ( .A(KEYINPUT8), .B(n1182), .ZN(n1230) );
INV_X1 U958 ( .A(n988), .ZN(n1182) );
XNOR2_X1 U959 ( .A(n1232), .B(n1233), .ZN(n988) );
NOR2_X1 U960 ( .A1(n1107), .A2(n1108), .ZN(n1233) );
INV_X1 U961 ( .A(G210), .ZN(n1108) );
NOR2_X1 U962 ( .A1(n1234), .A2(G237), .ZN(n1107) );
NAND2_X1 U963 ( .A1(n1235), .A2(n1161), .ZN(n1232) );
INV_X1 U964 ( .A(G902), .ZN(n1161) );
XOR2_X1 U965 ( .A(n1104), .B(n1236), .Z(n1235) );
XOR2_X1 U966 ( .A(G125), .B(n1237), .Z(n1236) );
NOR2_X1 U967 ( .A1(KEYINPUT41), .A2(n1039), .ZN(n1237) );
XNOR2_X1 U968 ( .A(n1047), .B(n1238), .ZN(n1104) );
AND2_X1 U969 ( .A1(n972), .A2(G224), .ZN(n1238) );
XNOR2_X1 U970 ( .A(n1239), .B(n1240), .ZN(n1047) );
XNOR2_X1 U971 ( .A(n1069), .B(n1241), .ZN(n1240) );
XNOR2_X1 U972 ( .A(KEYINPUT48), .B(n1242), .ZN(n1241) );
INV_X1 U973 ( .A(G110), .ZN(n1242) );
XOR2_X1 U974 ( .A(n1243), .B(n1244), .Z(n1239) );
XNOR2_X1 U975 ( .A(n1085), .B(n1077), .ZN(n1243) );
XNOR2_X1 U976 ( .A(G113), .B(n1245), .ZN(n1085) );
XNOR2_X1 U977 ( .A(G119), .B(n1200), .ZN(n1245) );
NOR2_X1 U978 ( .A1(n1246), .A2(n1012), .ZN(n1121) );
INV_X1 U979 ( .A(n1006), .ZN(n1012) );
NAND2_X1 U980 ( .A1(G221), .A2(n1228), .ZN(n1006) );
NAND2_X1 U981 ( .A1(n1247), .A2(G234), .ZN(n1228) );
INV_X1 U982 ( .A(n1234), .ZN(n1247) );
XOR2_X1 U983 ( .A(G902), .B(KEYINPUT16), .Z(n1234) );
INV_X1 U984 ( .A(n1002), .ZN(n1246) );
XNOR2_X1 U985 ( .A(n1248), .B(G469), .ZN(n1002) );
NAND2_X1 U986 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
XOR2_X1 U987 ( .A(n1251), .B(n1252), .Z(n1250) );
XNOR2_X1 U988 ( .A(n1253), .B(n1088), .ZN(n1252) );
XNOR2_X1 U989 ( .A(n1254), .B(n1035), .ZN(n1088) );
XOR2_X1 U990 ( .A(G134), .B(n1213), .Z(n1035) );
XOR2_X1 U991 ( .A(G137), .B(KEYINPUT36), .Z(n1213) );
NAND2_X1 U992 ( .A1(KEYINPUT52), .A2(n1181), .ZN(n1254) );
INV_X1 U993 ( .A(G131), .ZN(n1181) );
NAND2_X1 U994 ( .A1(KEYINPUT12), .A2(n1255), .ZN(n1253) );
XNOR2_X1 U995 ( .A(n1256), .B(n1095), .ZN(n1255) );
XNOR2_X1 U996 ( .A(G110), .B(n1174), .ZN(n1095) );
NAND2_X1 U997 ( .A1(KEYINPUT19), .A2(n1098), .ZN(n1256) );
NOR2_X1 U998 ( .A1(n1028), .A2(G953), .ZN(n1098) );
INV_X1 U999 ( .A(G227), .ZN(n1028) );
XNOR2_X1 U1000 ( .A(n1257), .B(KEYINPUT0), .ZN(n1251) );
NAND2_X1 U1001 ( .A1(n1258), .A2(KEYINPUT13), .ZN(n1257) );
XNOR2_X1 U1002 ( .A(n1096), .B(KEYINPUT10), .ZN(n1258) );
XOR2_X1 U1003 ( .A(n1259), .B(n1089), .Z(n1096) );
INV_X1 U1004 ( .A(n1039), .ZN(n1089) );
XOR2_X1 U1005 ( .A(G128), .B(n1260), .Z(n1039) );
XNOR2_X1 U1006 ( .A(n1261), .B(n1077), .ZN(n1259) );
INV_X1 U1007 ( .A(G101), .ZN(n1077) );
NAND2_X1 U1008 ( .A1(KEYINPUT51), .A2(n1262), .ZN(n1261) );
XNOR2_X1 U1009 ( .A(G107), .B(n1069), .ZN(n1262) );
XNOR2_X1 U1010 ( .A(G902), .B(KEYINPUT57), .ZN(n1249) );
NOR2_X1 U1011 ( .A1(n1202), .A2(n1015), .ZN(n1186) );
XNOR2_X1 U1012 ( .A(n1263), .B(G475), .ZN(n1015) );
OR2_X1 U1013 ( .A1(n1062), .A2(G902), .ZN(n1263) );
XNOR2_X1 U1014 ( .A(n1264), .B(n1265), .ZN(n1062) );
XOR2_X1 U1015 ( .A(n1260), .B(n1036), .Z(n1265) );
XOR2_X1 U1016 ( .A(G125), .B(n1266), .Z(n1036) );
XNOR2_X1 U1017 ( .A(n1174), .B(G131), .ZN(n1266) );
INV_X1 U1018 ( .A(G140), .ZN(n1174) );
XNOR2_X1 U1019 ( .A(G146), .B(n1267), .ZN(n1260) );
XOR2_X1 U1020 ( .A(n1268), .B(n1269), .Z(n1264) );
NOR2_X1 U1021 ( .A1(n1211), .A2(n1231), .ZN(n1269) );
INV_X1 U1022 ( .A(G214), .ZN(n1231) );
INV_X1 U1023 ( .A(n1075), .ZN(n1211) );
NOR2_X1 U1024 ( .A1(G953), .A2(G237), .ZN(n1075) );
NAND3_X1 U1025 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1268) );
NAND2_X1 U1026 ( .A1(KEYINPUT39), .A2(n1273), .ZN(n1272) );
NAND3_X1 U1027 ( .A1(n1274), .A2(n1275), .A3(n1069), .ZN(n1271) );
INV_X1 U1028 ( .A(KEYINPUT39), .ZN(n1275) );
OR2_X1 U1029 ( .A1(n1069), .A2(n1274), .ZN(n1270) );
NOR2_X1 U1030 ( .A1(KEYINPUT55), .A2(n1273), .ZN(n1274) );
XNOR2_X1 U1031 ( .A(G113), .B(G122), .ZN(n1273) );
INV_X1 U1032 ( .A(G104), .ZN(n1069) );
XNOR2_X1 U1033 ( .A(n1016), .B(G478), .ZN(n1202) );
OR2_X1 U1034 ( .A1(n1056), .A2(G902), .ZN(n1016) );
XNOR2_X1 U1035 ( .A(n1276), .B(n1277), .ZN(n1056) );
XOR2_X1 U1036 ( .A(n1278), .B(n1244), .Z(n1277) );
XOR2_X1 U1037 ( .A(G107), .B(G122), .Z(n1244) );
NOR3_X1 U1038 ( .A1(n1279), .A2(KEYINPUT33), .A3(n1218), .ZN(n1278) );
NAND2_X1 U1039 ( .A1(G234), .A2(n972), .ZN(n1218) );
INV_X1 U1040 ( .A(G953), .ZN(n972) );
INV_X1 U1041 ( .A(G217), .ZN(n1279) );
XOR2_X1 U1042 ( .A(n1280), .B(n1281), .Z(n1276) );
XNOR2_X1 U1043 ( .A(G134), .B(n1200), .ZN(n1281) );
INV_X1 U1044 ( .A(G116), .ZN(n1200) );
NAND3_X1 U1045 ( .A1(n1282), .A2(n1283), .A3(n1284), .ZN(n1280) );
NAND2_X1 U1046 ( .A1(G143), .A2(n1227), .ZN(n1284) );
INV_X1 U1047 ( .A(G128), .ZN(n1227) );
NAND2_X1 U1048 ( .A1(KEYINPUT31), .A2(n1285), .ZN(n1283) );
NAND2_X1 U1049 ( .A1(n1286), .A2(n1267), .ZN(n1285) );
XNOR2_X1 U1050 ( .A(KEYINPUT56), .B(G128), .ZN(n1286) );
NAND2_X1 U1051 ( .A1(n1287), .A2(n1288), .ZN(n1282) );
INV_X1 U1052 ( .A(KEYINPUT31), .ZN(n1288) );
NAND2_X1 U1053 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
OR2_X1 U1054 ( .A1(G128), .A2(KEYINPUT56), .ZN(n1290) );
NAND3_X1 U1055 ( .A1(G128), .A2(n1267), .A3(KEYINPUT56), .ZN(n1289) );
INV_X1 U1056 ( .A(G143), .ZN(n1267) );
endmodule


