//Key = 0101100000110001111001111011111001000100001011100010111110001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363;

NAND2_X1 U746 ( .A1(n1027), .A2(n1028), .ZN(G9) );
NAND2_X1 U747 ( .A1(G107), .A2(n1029), .ZN(n1028) );
XOR2_X1 U748 ( .A(KEYINPUT55), .B(n1030), .Z(n1027) );
NOR2_X1 U749 ( .A1(G107), .A2(n1029), .ZN(n1030) );
NOR2_X1 U750 ( .A1(n1031), .A2(n1032), .ZN(G75) );
NOR3_X1 U751 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1032) );
NAND3_X1 U752 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1033) );
NAND2_X1 U753 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U754 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND4_X1 U755 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
NAND3_X1 U756 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND2_X1 U757 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U758 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND3_X1 U759 ( .A1(n1050), .A2(n1054), .A3(n1055), .ZN(n1041) );
NAND2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NAND3_X1 U761 ( .A1(n1058), .A2(n1059), .A3(n1044), .ZN(n1057) );
NAND2_X1 U762 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U763 ( .A1(n1062), .A2(n1043), .ZN(n1058) );
XNOR2_X1 U764 ( .A(n1063), .B(n1064), .ZN(n1062) );
INV_X1 U765 ( .A(n1065), .ZN(n1056) );
INV_X1 U766 ( .A(n1066), .ZN(n1039) );
NOR3_X1 U767 ( .A1(n1067), .A2(G953), .A3(G952), .ZN(n1031) );
INV_X1 U768 ( .A(n1036), .ZN(n1067) );
NAND4_X1 U769 ( .A1(n1043), .A2(n1045), .A3(n1068), .A4(n1069), .ZN(n1036) );
NOR4_X1 U770 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
XOR2_X1 U771 ( .A(KEYINPUT59), .B(n1074), .Z(n1073) );
XNOR2_X1 U772 ( .A(G472), .B(n1075), .ZN(n1072) );
XOR2_X1 U773 ( .A(KEYINPUT34), .B(n1076), .Z(n1071) );
NOR2_X1 U774 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR3_X1 U775 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1068) );
NOR2_X1 U776 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
INV_X1 U777 ( .A(n1077), .ZN(n1083) );
XOR2_X1 U778 ( .A(n1078), .B(KEYINPUT56), .Z(n1082) );
XOR2_X1 U779 ( .A(n1084), .B(KEYINPUT46), .Z(n1079) );
NAND2_X1 U780 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XNOR2_X1 U781 ( .A(n1087), .B(KEYINPUT44), .ZN(n1085) );
XOR2_X1 U782 ( .A(n1088), .B(n1089), .Z(G72) );
NOR2_X1 U783 ( .A1(n1090), .A2(n1037), .ZN(n1089) );
AND2_X1 U784 ( .A1(G227), .A2(G900), .ZN(n1090) );
NAND2_X1 U785 ( .A1(n1091), .A2(n1092), .ZN(n1088) );
NAND2_X1 U786 ( .A1(n1093), .A2(n1037), .ZN(n1092) );
XOR2_X1 U787 ( .A(n1035), .B(n1094), .Z(n1093) );
NAND3_X1 U788 ( .A1(n1094), .A2(G900), .A3(G953), .ZN(n1091) );
AND2_X1 U789 ( .A1(n1095), .A2(KEYINPUT17), .ZN(n1094) );
XOR2_X1 U790 ( .A(n1096), .B(n1097), .Z(n1095) );
XOR2_X1 U791 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U792 ( .A1(G131), .A2(KEYINPUT6), .ZN(n1098) );
XOR2_X1 U793 ( .A(n1100), .B(n1101), .Z(n1096) );
XOR2_X1 U794 ( .A(n1102), .B(n1103), .Z(G69) );
NOR2_X1 U795 ( .A1(n1104), .A2(n1037), .ZN(n1103) );
AND2_X1 U796 ( .A1(G224), .A2(G898), .ZN(n1104) );
NAND2_X1 U797 ( .A1(n1105), .A2(n1106), .ZN(n1102) );
NAND2_X1 U798 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
OR2_X1 U799 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U800 ( .A(KEYINPUT42), .B(n1111), .Z(n1105) );
NOR4_X1 U801 ( .A1(n1110), .A2(n1107), .A3(n1109), .A4(n1112), .ZN(n1111) );
NOR2_X1 U802 ( .A1(G898), .A2(n1037), .ZN(n1112) );
NOR2_X1 U803 ( .A1(n1113), .A2(n1114), .ZN(n1109) );
AND2_X1 U804 ( .A1(n1037), .A2(n1115), .ZN(n1107) );
NAND3_X1 U805 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
AND3_X1 U806 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1118) );
AND2_X1 U807 ( .A1(n1122), .A2(n1113), .ZN(n1110) );
NAND3_X1 U808 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1113) );
NAND2_X1 U809 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U810 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
INV_X1 U811 ( .A(KEYINPUT47), .ZN(n1129) );
XOR2_X1 U812 ( .A(KEYINPUT53), .B(n1130), .Z(n1128) );
OR3_X1 U813 ( .A1(n1126), .A2(n1130), .A3(KEYINPUT47), .ZN(n1124) );
NAND2_X1 U814 ( .A1(n1130), .A2(KEYINPUT47), .ZN(n1123) );
XNOR2_X1 U815 ( .A(KEYINPUT12), .B(n1131), .ZN(n1122) );
NOR2_X1 U816 ( .A1(n1132), .A2(n1133), .ZN(G66) );
NOR3_X1 U817 ( .A1(n1077), .A2(n1134), .A3(n1135), .ZN(n1133) );
NOR4_X1 U818 ( .A1(n1136), .A2(n1137), .A3(KEYINPUT51), .A4(n1078), .ZN(n1135) );
INV_X1 U819 ( .A(n1138), .ZN(n1137) );
INV_X1 U820 ( .A(n1139), .ZN(n1136) );
NOR2_X1 U821 ( .A1(n1140), .A2(n1139), .ZN(n1134) );
NOR3_X1 U822 ( .A1(n1078), .A2(KEYINPUT51), .A3(n1141), .ZN(n1140) );
NOR2_X1 U823 ( .A1(n1132), .A2(n1142), .ZN(G63) );
XOR2_X1 U824 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U825 ( .A(n1145), .B(KEYINPUT5), .Z(n1144) );
NAND2_X1 U826 ( .A1(n1138), .A2(G478), .ZN(n1143) );
NOR2_X1 U827 ( .A1(n1132), .A2(n1146), .ZN(G60) );
XOR2_X1 U828 ( .A(n1147), .B(n1148), .Z(n1146) );
NAND2_X1 U829 ( .A1(n1138), .A2(G475), .ZN(n1147) );
XOR2_X1 U830 ( .A(G104), .B(n1149), .Z(G6) );
NOR2_X1 U831 ( .A1(n1150), .A2(n1052), .ZN(n1149) );
NOR2_X1 U832 ( .A1(n1132), .A2(n1151), .ZN(G57) );
XOR2_X1 U833 ( .A(n1152), .B(n1153), .Z(n1151) );
XNOR2_X1 U834 ( .A(n1154), .B(n1155), .ZN(n1153) );
NOR2_X1 U835 ( .A1(KEYINPUT32), .A2(n1156), .ZN(n1155) );
XOR2_X1 U836 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U837 ( .A(n1159), .B(n1160), .ZN(n1158) );
NOR3_X1 U838 ( .A1(n1161), .A2(KEYINPUT62), .A3(n1162), .ZN(n1160) );
NOR2_X1 U839 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XNOR2_X1 U840 ( .A(n1165), .B(KEYINPUT31), .ZN(n1164) );
NOR2_X1 U841 ( .A1(n1166), .A2(n1167), .ZN(n1163) );
NOR2_X1 U842 ( .A1(n1168), .A2(n1169), .ZN(n1166) );
NOR2_X1 U843 ( .A1(n1170), .A2(n1171), .ZN(n1161) );
INV_X1 U844 ( .A(n1168), .ZN(n1171) );
NOR2_X1 U845 ( .A1(n1167), .A2(n1169), .ZN(n1170) );
INV_X1 U846 ( .A(KEYINPUT28), .ZN(n1169) );
NAND2_X1 U847 ( .A1(n1138), .A2(G472), .ZN(n1157) );
NAND2_X1 U848 ( .A1(KEYINPUT60), .A2(n1172), .ZN(n1152) );
NOR2_X1 U849 ( .A1(n1132), .A2(n1173), .ZN(G54) );
NOR2_X1 U850 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XOR2_X1 U851 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U852 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND2_X1 U853 ( .A1(n1138), .A2(G469), .ZN(n1176) );
NOR2_X1 U854 ( .A1(n1179), .A2(n1178), .ZN(n1174) );
INV_X1 U855 ( .A(KEYINPUT0), .ZN(n1178) );
NAND2_X1 U856 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NAND2_X1 U857 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
XNOR2_X1 U858 ( .A(n1165), .B(n1184), .ZN(n1183) );
XNOR2_X1 U859 ( .A(n1185), .B(n1186), .ZN(n1182) );
XOR2_X1 U860 ( .A(n1187), .B(KEYINPUT13), .Z(n1180) );
NAND2_X1 U861 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XNOR2_X1 U862 ( .A(n1186), .B(n1190), .ZN(n1189) );
NOR2_X1 U863 ( .A1(KEYINPUT19), .A2(n1191), .ZN(n1186) );
XNOR2_X1 U864 ( .A(n1192), .B(n1193), .ZN(n1191) );
NOR2_X1 U865 ( .A1(G140), .A2(KEYINPUT25), .ZN(n1193) );
XNOR2_X1 U866 ( .A(n1184), .B(n1167), .ZN(n1188) );
XOR2_X1 U867 ( .A(n1194), .B(n1195), .Z(n1184) );
NOR2_X1 U868 ( .A1(KEYINPUT61), .A2(n1196), .ZN(n1195) );
XNOR2_X1 U869 ( .A(G101), .B(n1197), .ZN(n1196) );
NOR2_X1 U870 ( .A1(n1132), .A2(n1198), .ZN(G51) );
XOR2_X1 U871 ( .A(n1199), .B(n1200), .Z(n1198) );
XOR2_X1 U872 ( .A(n1201), .B(n1202), .Z(n1200) );
NAND2_X1 U873 ( .A1(n1203), .A2(n1204), .ZN(n1201) );
XOR2_X1 U874 ( .A(n1205), .B(KEYINPUT35), .Z(n1203) );
NAND2_X1 U875 ( .A1(n1138), .A2(G210), .ZN(n1199) );
NOR2_X1 U876 ( .A1(n1206), .A2(n1141), .ZN(n1138) );
NOR2_X1 U877 ( .A1(n1034), .A2(n1207), .ZN(n1141) );
XOR2_X1 U878 ( .A(KEYINPUT41), .B(n1035), .Z(n1207) );
NAND4_X1 U879 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1035) );
NOR4_X1 U880 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1211) );
NOR2_X1 U881 ( .A1(n1216), .A2(n1217), .ZN(n1210) );
NOR3_X1 U882 ( .A1(n1218), .A2(n1219), .A3(n1053), .ZN(n1217) );
INV_X1 U883 ( .A(n1220), .ZN(n1053) );
XNOR2_X1 U884 ( .A(n1221), .B(KEYINPUT2), .ZN(n1219) );
NAND2_X1 U885 ( .A1(n1222), .A2(n1116), .ZN(n1034) );
AND4_X1 U886 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1029), .ZN(n1116) );
NAND2_X1 U887 ( .A1(n1220), .A2(n1226), .ZN(n1029) );
NAND2_X1 U888 ( .A1(n1227), .A2(n1226), .ZN(n1224) );
INV_X1 U889 ( .A(n1150), .ZN(n1226) );
NAND2_X1 U890 ( .A1(n1228), .A2(n1050), .ZN(n1150) );
XNOR2_X1 U891 ( .A(n1229), .B(KEYINPUT23), .ZN(n1227) );
NAND2_X1 U892 ( .A1(n1230), .A2(n1228), .ZN(n1223) );
INV_X1 U893 ( .A(n1047), .ZN(n1230) );
XOR2_X1 U894 ( .A(n1231), .B(KEYINPUT26), .Z(n1222) );
NAND4_X1 U895 ( .A1(n1232), .A2(n1117), .A3(n1119), .A4(n1120), .ZN(n1231) );
XOR2_X1 U896 ( .A(n1121), .B(KEYINPUT8), .Z(n1232) );
NOR2_X1 U897 ( .A1(n1037), .A2(G952), .ZN(n1132) );
XNOR2_X1 U898 ( .A(G146), .B(n1209), .ZN(G48) );
NAND3_X1 U899 ( .A1(n1229), .A2(n1233), .A3(n1234), .ZN(n1209) );
XOR2_X1 U900 ( .A(G143), .B(n1216), .Z(G45) );
AND3_X1 U901 ( .A1(n1221), .A2(n1233), .A3(n1235), .ZN(n1216) );
AND3_X1 U902 ( .A1(n1074), .A2(n1236), .A3(n1237), .ZN(n1235) );
XNOR2_X1 U903 ( .A(G140), .B(n1208), .ZN(G42) );
NAND4_X1 U904 ( .A1(n1238), .A2(n1229), .A3(n1239), .A4(n1240), .ZN(n1208) );
XNOR2_X1 U905 ( .A(n1241), .B(n1215), .ZN(G39) );
AND3_X1 U906 ( .A1(n1242), .A2(n1238), .A3(n1243), .ZN(n1215) );
NAND2_X1 U907 ( .A1(n1244), .A2(n1245), .ZN(G36) );
NAND2_X1 U908 ( .A1(G134), .A2(n1246), .ZN(n1245) );
XOR2_X1 U909 ( .A(KEYINPUT52), .B(n1247), .Z(n1244) );
NOR2_X1 U910 ( .A1(G134), .A2(n1246), .ZN(n1247) );
NAND3_X1 U911 ( .A1(n1220), .A2(n1221), .A3(n1238), .ZN(n1246) );
XNOR2_X1 U912 ( .A(n1248), .B(n1214), .ZN(G33) );
AND3_X1 U913 ( .A1(n1229), .A2(n1221), .A3(n1238), .ZN(n1214) );
INV_X1 U914 ( .A(n1218), .ZN(n1238) );
NAND4_X1 U915 ( .A1(n1044), .A2(n1045), .A3(n1060), .A4(n1237), .ZN(n1218) );
INV_X1 U916 ( .A(n1061), .ZN(n1045) );
XNOR2_X1 U917 ( .A(G128), .B(n1249), .ZN(G30) );
NAND2_X1 U918 ( .A1(KEYINPUT3), .A2(n1213), .ZN(n1249) );
AND3_X1 U919 ( .A1(n1220), .A2(n1233), .A3(n1234), .ZN(n1213) );
AND3_X1 U920 ( .A1(n1240), .A2(n1237), .A3(n1242), .ZN(n1234) );
XNOR2_X1 U921 ( .A(n1172), .B(n1250), .ZN(G3) );
NOR3_X1 U922 ( .A1(n1047), .A2(n1251), .A3(n1252), .ZN(n1250) );
INV_X1 U923 ( .A(n1233), .ZN(n1252) );
XOR2_X1 U924 ( .A(n1253), .B(KEYINPUT29), .Z(n1251) );
NAND2_X1 U925 ( .A1(n1055), .A2(n1221), .ZN(n1047) );
INV_X1 U926 ( .A(G101), .ZN(n1172) );
XOR2_X1 U927 ( .A(n1212), .B(n1254), .Z(G27) );
NOR2_X1 U928 ( .A1(KEYINPUT49), .A2(n1255), .ZN(n1254) );
AND3_X1 U929 ( .A1(n1065), .A2(n1229), .A3(n1256), .ZN(n1212) );
AND3_X1 U930 ( .A1(n1239), .A2(n1237), .A3(n1240), .ZN(n1256) );
NAND2_X1 U931 ( .A1(n1066), .A2(n1257), .ZN(n1237) );
NAND4_X1 U932 ( .A1(G902), .A2(G953), .A3(n1258), .A4(n1259), .ZN(n1257) );
INV_X1 U933 ( .A(G900), .ZN(n1259) );
XNOR2_X1 U934 ( .A(n1260), .B(n1117), .ZN(G24) );
NAND4_X1 U935 ( .A1(n1261), .A2(n1050), .A3(n1074), .A4(n1236), .ZN(n1117) );
NAND2_X1 U936 ( .A1(n1262), .A2(n1263), .ZN(n1050) );
OR3_X1 U937 ( .A1(n1242), .A2(n1240), .A3(KEYINPUT20), .ZN(n1263) );
NAND2_X1 U938 ( .A1(KEYINPUT20), .A2(n1221), .ZN(n1262) );
NAND2_X1 U939 ( .A1(KEYINPUT50), .A2(n1264), .ZN(n1260) );
XOR2_X1 U940 ( .A(KEYINPUT63), .B(G122), .Z(n1264) );
XOR2_X1 U941 ( .A(n1119), .B(n1265), .Z(G21) );
NAND2_X1 U942 ( .A1(KEYINPUT18), .A2(G119), .ZN(n1265) );
NAND3_X1 U943 ( .A1(n1242), .A2(n1243), .A3(n1261), .ZN(n1119) );
INV_X1 U944 ( .A(n1266), .ZN(n1242) );
XNOR2_X1 U945 ( .A(G116), .B(n1121), .ZN(G18) );
NAND3_X1 U946 ( .A1(n1220), .A2(n1221), .A3(n1261), .ZN(n1121) );
NOR2_X1 U947 ( .A1(n1074), .A2(n1267), .ZN(n1220) );
XNOR2_X1 U948 ( .A(G113), .B(n1120), .ZN(G15) );
NAND3_X1 U949 ( .A1(n1229), .A2(n1221), .A3(n1261), .ZN(n1120) );
AND2_X1 U950 ( .A1(n1065), .A2(n1253), .ZN(n1261) );
NOR3_X1 U951 ( .A1(n1061), .A2(n1044), .A3(n1060), .ZN(n1065) );
NOR2_X1 U952 ( .A1(n1240), .A2(n1266), .ZN(n1221) );
INV_X1 U953 ( .A(n1052), .ZN(n1229) );
NAND2_X1 U954 ( .A1(n1267), .A2(n1074), .ZN(n1052) );
XOR2_X1 U955 ( .A(n1225), .B(n1268), .Z(G12) );
XNOR2_X1 U956 ( .A(KEYINPUT4), .B(n1192), .ZN(n1268) );
NAND2_X1 U957 ( .A1(n1269), .A2(n1228), .ZN(n1225) );
AND2_X1 U958 ( .A1(n1233), .A2(n1253), .ZN(n1228) );
NAND2_X1 U959 ( .A1(n1066), .A2(n1270), .ZN(n1253) );
NAND4_X1 U960 ( .A1(G902), .A2(G953), .A3(n1258), .A4(n1271), .ZN(n1270) );
INV_X1 U961 ( .A(G898), .ZN(n1271) );
NAND3_X1 U962 ( .A1(n1258), .A2(n1037), .A3(G952), .ZN(n1066) );
NAND2_X1 U963 ( .A1(G237), .A2(G234), .ZN(n1258) );
NOR3_X1 U964 ( .A1(n1043), .A2(n1044), .A3(n1061), .ZN(n1233) );
NAND2_X1 U965 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NAND2_X1 U966 ( .A1(G214), .A2(n1272), .ZN(n1064) );
NAND2_X1 U967 ( .A1(G221), .A2(n1273), .ZN(n1063) );
INV_X1 U968 ( .A(n1070), .ZN(n1044) );
XNOR2_X1 U969 ( .A(n1274), .B(n1275), .ZN(n1070) );
NOR2_X1 U970 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XNOR2_X1 U971 ( .A(KEYINPUT43), .B(n1272), .ZN(n1277) );
OR2_X1 U972 ( .A1(G902), .A2(G237), .ZN(n1272) );
INV_X1 U973 ( .A(G210), .ZN(n1276) );
NAND2_X1 U974 ( .A1(n1278), .A2(n1206), .ZN(n1274) );
XOR2_X1 U975 ( .A(n1202), .B(n1279), .Z(n1278) );
NAND2_X1 U976 ( .A1(n1204), .A2(n1205), .ZN(n1279) );
NAND2_X1 U977 ( .A1(n1280), .A2(n1281), .ZN(n1205) );
OR2_X1 U978 ( .A1(n1281), .A2(n1280), .ZN(n1204) );
XNOR2_X1 U979 ( .A(n1282), .B(n1283), .ZN(n1280) );
NAND2_X1 U980 ( .A1(G224), .A2(n1284), .ZN(n1281) );
NAND2_X1 U981 ( .A1(n1285), .A2(n1286), .ZN(n1202) );
OR2_X1 U982 ( .A1(n1287), .A2(n1131), .ZN(n1286) );
XOR2_X1 U983 ( .A(n1288), .B(KEYINPUT14), .Z(n1285) );
NAND2_X1 U984 ( .A1(n1131), .A2(n1287), .ZN(n1288) );
XNOR2_X1 U985 ( .A(n1289), .B(n1130), .ZN(n1287) );
XNOR2_X1 U986 ( .A(n1290), .B(n1291), .ZN(n1130) );
NOR2_X1 U987 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XOR2_X1 U988 ( .A(n1294), .B(KEYINPUT30), .Z(n1293) );
NAND2_X1 U989 ( .A1(G119), .A2(n1295), .ZN(n1294) );
NAND2_X1 U990 ( .A1(KEYINPUT45), .A2(n1296), .ZN(n1290) );
INV_X1 U991 ( .A(G113), .ZN(n1296) );
NAND2_X1 U992 ( .A1(KEYINPUT24), .A2(n1126), .ZN(n1289) );
XOR2_X1 U993 ( .A(G101), .B(n1297), .Z(n1126) );
NOR2_X1 U994 ( .A1(KEYINPUT58), .A2(n1197), .ZN(n1297) );
XNOR2_X1 U995 ( .A(G104), .B(G107), .ZN(n1197) );
INV_X1 U996 ( .A(n1114), .ZN(n1131) );
XNOR2_X1 U997 ( .A(n1298), .B(n1299), .ZN(n1114) );
XNOR2_X1 U998 ( .A(G110), .B(KEYINPUT21), .ZN(n1298) );
INV_X1 U999 ( .A(n1060), .ZN(n1043) );
XNOR2_X1 U1000 ( .A(n1300), .B(G469), .ZN(n1060) );
NAND2_X1 U1001 ( .A1(n1301), .A2(n1206), .ZN(n1300) );
XOR2_X1 U1002 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U1003 ( .A(n1304), .B(n1305), .Z(n1303) );
XNOR2_X1 U1004 ( .A(n1306), .B(n1167), .ZN(n1304) );
NAND2_X1 U1005 ( .A1(KEYINPUT10), .A2(n1194), .ZN(n1306) );
XOR2_X1 U1006 ( .A(n1100), .B(G128), .Z(n1194) );
XOR2_X1 U1007 ( .A(n1307), .B(KEYINPUT40), .Z(n1100) );
NAND2_X1 U1008 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND2_X1 U1009 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
XOR2_X1 U1010 ( .A(KEYINPUT27), .B(n1312), .Z(n1308) );
NOR2_X1 U1011 ( .A1(n1310), .A2(n1311), .ZN(n1312) );
XOR2_X1 U1012 ( .A(n1313), .B(n1314), .Z(n1302) );
XNOR2_X1 U1013 ( .A(n1192), .B(G107), .ZN(n1314) );
XNOR2_X1 U1014 ( .A(n1185), .B(G101), .ZN(n1313) );
INV_X1 U1015 ( .A(n1190), .ZN(n1185) );
NAND2_X1 U1016 ( .A1(G227), .A2(n1284), .ZN(n1190) );
INV_X1 U1017 ( .A(n1048), .ZN(n1269) );
NAND2_X1 U1018 ( .A1(n1243), .A2(n1239), .ZN(n1048) );
XOR2_X1 U1019 ( .A(n1266), .B(KEYINPUT20), .Z(n1239) );
XNOR2_X1 U1020 ( .A(n1075), .B(n1315), .ZN(n1266) );
NOR2_X1 U1021 ( .A1(G472), .A2(KEYINPUT9), .ZN(n1315) );
NAND2_X1 U1022 ( .A1(n1316), .A2(n1206), .ZN(n1075) );
XOR2_X1 U1023 ( .A(n1317), .B(n1318), .Z(n1316) );
XNOR2_X1 U1024 ( .A(G101), .B(n1154), .ZN(n1318) );
AND2_X1 U1025 ( .A1(G210), .A2(n1319), .ZN(n1154) );
NAND3_X1 U1026 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1317) );
XOR2_X1 U1027 ( .A(KEYINPUT54), .B(n1323), .Z(n1322) );
NOR2_X1 U1028 ( .A1(n1159), .A2(n1324), .ZN(n1323) );
NAND2_X1 U1029 ( .A1(n1159), .A2(n1324), .ZN(n1321) );
XNOR2_X1 U1030 ( .A(n1167), .B(n1168), .ZN(n1324) );
XNOR2_X1 U1031 ( .A(n1282), .B(G128), .ZN(n1168) );
NAND2_X1 U1032 ( .A1(KEYINPUT11), .A2(n1325), .ZN(n1282) );
XNOR2_X1 U1033 ( .A(n1311), .B(n1310), .ZN(n1325) );
INV_X1 U1034 ( .A(G146), .ZN(n1311) );
INV_X1 U1035 ( .A(n1165), .ZN(n1167) );
XOR2_X1 U1036 ( .A(G131), .B(n1099), .Z(n1165) );
XNOR2_X1 U1037 ( .A(n1241), .B(G134), .ZN(n1099) );
INV_X1 U1038 ( .A(G137), .ZN(n1241) );
AND3_X1 U1039 ( .A1(n1326), .A2(n1327), .A3(n1328), .ZN(n1159) );
NAND2_X1 U1040 ( .A1(n1292), .A2(n1329), .ZN(n1328) );
NOR2_X1 U1041 ( .A1(n1295), .A2(G119), .ZN(n1292) );
OR3_X1 U1042 ( .A1(n1329), .A2(G116), .A3(G119), .ZN(n1327) );
INV_X1 U1043 ( .A(n1330), .ZN(n1329) );
NAND2_X1 U1044 ( .A1(n1331), .A2(G119), .ZN(n1326) );
XNOR2_X1 U1045 ( .A(G116), .B(n1330), .ZN(n1331) );
NOR2_X1 U1046 ( .A1(G113), .A2(KEYINPUT39), .ZN(n1330) );
XOR2_X1 U1047 ( .A(KEYINPUT37), .B(KEYINPUT36), .Z(n1320) );
AND2_X1 U1048 ( .A1(n1055), .A2(n1240), .ZN(n1243) );
XOR2_X1 U1049 ( .A(n1332), .B(n1078), .Z(n1240) );
NAND2_X1 U1050 ( .A1(G217), .A2(n1273), .ZN(n1078) );
NAND2_X1 U1051 ( .A1(G234), .A2(n1206), .ZN(n1273) );
XNOR2_X1 U1052 ( .A(n1077), .B(KEYINPUT57), .ZN(n1332) );
NOR2_X1 U1053 ( .A1(n1139), .A2(G902), .ZN(n1077) );
XNOR2_X1 U1054 ( .A(n1333), .B(n1334), .ZN(n1139) );
XNOR2_X1 U1055 ( .A(n1335), .B(n1336), .ZN(n1334) );
XNOR2_X1 U1056 ( .A(n1101), .B(n1337), .ZN(n1336) );
NOR3_X1 U1057 ( .A1(n1338), .A2(KEYINPUT38), .A3(n1339), .ZN(n1337) );
INV_X1 U1058 ( .A(G221), .ZN(n1338) );
XOR2_X1 U1059 ( .A(G140), .B(n1283), .Z(n1101) );
XNOR2_X1 U1060 ( .A(n1255), .B(G128), .ZN(n1283) );
XOR2_X1 U1061 ( .A(n1340), .B(n1341), .Z(n1333) );
XNOR2_X1 U1062 ( .A(G119), .B(n1192), .ZN(n1341) );
INV_X1 U1063 ( .A(G110), .ZN(n1192) );
XNOR2_X1 U1064 ( .A(G137), .B(KEYINPUT15), .ZN(n1340) );
NOR2_X1 U1065 ( .A1(n1236), .A2(n1074), .ZN(n1055) );
XNOR2_X1 U1066 ( .A(n1342), .B(G475), .ZN(n1074) );
NAND2_X1 U1067 ( .A1(n1148), .A2(n1206), .ZN(n1342) );
XOR2_X1 U1068 ( .A(n1343), .B(n1344), .Z(n1148) );
XNOR2_X1 U1069 ( .A(n1305), .B(n1345), .ZN(n1344) );
XNOR2_X1 U1070 ( .A(n1299), .B(n1335), .ZN(n1345) );
XOR2_X1 U1071 ( .A(G146), .B(KEYINPUT7), .Z(n1335) );
XOR2_X1 U1072 ( .A(G104), .B(G140), .Z(n1305) );
XOR2_X1 U1073 ( .A(n1346), .B(n1347), .Z(n1343) );
XNOR2_X1 U1074 ( .A(n1255), .B(G113), .ZN(n1347) );
INV_X1 U1075 ( .A(G125), .ZN(n1255) );
NAND2_X1 U1076 ( .A1(KEYINPUT1), .A2(n1348), .ZN(n1346) );
XOR2_X1 U1077 ( .A(n1310), .B(n1349), .Z(n1348) );
XNOR2_X1 U1078 ( .A(n1248), .B(n1350), .ZN(n1349) );
AND2_X1 U1079 ( .A1(n1319), .A2(G214), .ZN(n1350) );
NOR2_X1 U1080 ( .A1(n1351), .A2(G237), .ZN(n1319) );
INV_X1 U1081 ( .A(G131), .ZN(n1248) );
INV_X1 U1082 ( .A(n1267), .ZN(n1236) );
NOR2_X1 U1083 ( .A1(n1080), .A2(n1352), .ZN(n1267) );
AND2_X1 U1084 ( .A1(n1087), .A2(n1086), .ZN(n1352) );
NOR2_X1 U1085 ( .A1(n1086), .A2(n1087), .ZN(n1080) );
AND2_X1 U1086 ( .A1(n1206), .A2(n1145), .ZN(n1087) );
NAND2_X1 U1087 ( .A1(n1353), .A2(n1354), .ZN(n1145) );
NAND2_X1 U1088 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
XOR2_X1 U1089 ( .A(n1357), .B(n1358), .Z(n1353) );
NOR2_X1 U1090 ( .A1(n1339), .A2(n1359), .ZN(n1358) );
INV_X1 U1091 ( .A(G217), .ZN(n1359) );
NAND2_X1 U1092 ( .A1(G234), .A2(n1284), .ZN(n1339) );
INV_X1 U1093 ( .A(n1351), .ZN(n1284) );
XOR2_X1 U1094 ( .A(n1037), .B(KEYINPUT22), .Z(n1351) );
INV_X1 U1095 ( .A(G953), .ZN(n1037) );
OR2_X1 U1096 ( .A1(n1356), .A2(n1355), .ZN(n1357) );
XNOR2_X1 U1097 ( .A(n1360), .B(n1361), .ZN(n1355) );
XNOR2_X1 U1098 ( .A(n1295), .B(n1362), .ZN(n1361) );
XOR2_X1 U1099 ( .A(G134), .B(G128), .Z(n1362) );
INV_X1 U1100 ( .A(G116), .ZN(n1295) );
XOR2_X1 U1101 ( .A(n1363), .B(n1299), .Z(n1360) );
XOR2_X1 U1102 ( .A(G122), .B(KEYINPUT16), .Z(n1299) );
XNOR2_X1 U1103 ( .A(G107), .B(n1310), .ZN(n1363) );
XOR2_X1 U1104 ( .A(G143), .B(KEYINPUT48), .Z(n1310) );
INV_X1 U1105 ( .A(KEYINPUT33), .ZN(n1356) );
INV_X1 U1106 ( .A(G902), .ZN(n1206) );
INV_X1 U1107 ( .A(G478), .ZN(n1086) );
endmodule


