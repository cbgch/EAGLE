//Key = 0110011010011011011000000100000111101010100000101001111110111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345;

XNOR2_X1 U743 ( .A(G107), .B(n1023), .ZN(G9) );
NAND4_X1 U744 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1023) );
NOR3_X1 U745 ( .A1(n1028), .A2(KEYINPUT57), .A3(n1029), .ZN(n1027) );
INV_X1 U746 ( .A(n1030), .ZN(n1028) );
OR2_X1 U747 ( .A1(n1031), .A2(n1032), .ZN(n1025) );
NAND2_X1 U748 ( .A1(n1033), .A2(n1031), .ZN(n1024) );
INV_X1 U749 ( .A(KEYINPUT6), .ZN(n1031) );
NAND2_X1 U750 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR2_X1 U751 ( .A1(n1036), .A2(n1037), .ZN(G75) );
NOR4_X1 U752 ( .A1(G953), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1037) );
NOR2_X1 U753 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U754 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR3_X1 U755 ( .A1(n1045), .A2(n1046), .A3(n1029), .ZN(n1044) );
NOR2_X1 U756 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U757 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U758 ( .A1(n1051), .A2(n1026), .ZN(n1049) );
NOR2_X1 U759 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U760 ( .A1(n1054), .A2(n1055), .ZN(n1047) );
NOR2_X1 U761 ( .A1(n1030), .A2(n1056), .ZN(n1054) );
NOR3_X1 U762 ( .A1(n1050), .A2(n1057), .A3(n1055), .ZN(n1043) );
NOR2_X1 U763 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U764 ( .A1(n1060), .A2(n1029), .ZN(n1059) );
NOR2_X1 U765 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U766 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U767 ( .A1(n1065), .A2(n1045), .ZN(n1058) );
INV_X1 U768 ( .A(n1066), .ZN(n1045) );
NOR2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR3_X1 U770 ( .A1(n1038), .A2(G953), .A3(G952), .ZN(n1036) );
AND2_X1 U771 ( .A1(n1069), .A2(n1070), .ZN(n1038) );
NOR4_X1 U772 ( .A1(n1071), .A2(n1072), .A3(n1055), .A4(n1073), .ZN(n1070) );
INV_X1 U773 ( .A(n1074), .ZN(n1055) );
NOR2_X1 U774 ( .A1(n1075), .A2(n1076), .ZN(n1072) );
NOR2_X1 U775 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U776 ( .A(n1079), .B(KEYINPUT17), .Z(n1077) );
INV_X1 U777 ( .A(n1080), .ZN(n1075) );
NOR4_X1 U778 ( .A1(n1081), .A2(n1082), .A3(n1050), .A4(n1083), .ZN(n1069) );
XOR2_X1 U779 ( .A(KEYINPUT20), .B(n1084), .Z(n1083) );
INV_X1 U780 ( .A(n1085), .ZN(n1050) );
NOR2_X1 U781 ( .A1(KEYINPUT2), .A2(n1079), .ZN(n1082) );
NOR3_X1 U782 ( .A1(n1086), .A2(n1080), .A3(n1078), .ZN(n1081) );
INV_X1 U783 ( .A(KEYINPUT2), .ZN(n1078) );
NAND2_X1 U784 ( .A1(n1087), .A2(n1088), .ZN(G72) );
NAND2_X1 U785 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XOR2_X1 U786 ( .A(n1091), .B(KEYINPUT3), .Z(n1087) );
NAND2_X1 U787 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U788 ( .A(KEYINPUT8), .B(n1089), .Z(n1093) );
XNOR2_X1 U789 ( .A(n1094), .B(n1095), .ZN(n1089) );
NOR2_X1 U790 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U791 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U792 ( .A1(KEYINPUT21), .A2(n1100), .ZN(n1099) );
XNOR2_X1 U793 ( .A(n1101), .B(n1102), .ZN(n1100) );
XOR2_X1 U794 ( .A(G140), .B(n1103), .Z(n1098) );
NOR2_X1 U795 ( .A1(G900), .A2(n1104), .ZN(n1096) );
NAND2_X1 U796 ( .A1(n1104), .A2(n1105), .ZN(n1094) );
NAND2_X1 U797 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XNOR2_X1 U798 ( .A(KEYINPUT54), .B(n1108), .ZN(n1107) );
INV_X1 U799 ( .A(n1090), .ZN(n1092) );
NAND2_X1 U800 ( .A1(G953), .A2(n1109), .ZN(n1090) );
NAND2_X1 U801 ( .A1(G900), .A2(G227), .ZN(n1109) );
NAND2_X1 U802 ( .A1(n1110), .A2(n1111), .ZN(G69) );
NAND2_X1 U803 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U804 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
OR2_X1 U805 ( .A1(KEYINPUT32), .A2(KEYINPUT37), .ZN(n1115) );
NAND3_X1 U806 ( .A1(KEYINPUT32), .A2(n1116), .A3(n1117), .ZN(n1110) );
INV_X1 U807 ( .A(n1113), .ZN(n1117) );
NAND2_X1 U808 ( .A1(G953), .A2(n1118), .ZN(n1113) );
NAND2_X1 U809 ( .A1(G898), .A2(G224), .ZN(n1118) );
XOR2_X1 U810 ( .A(KEYINPUT37), .B(n1114), .Z(n1116) );
AND2_X1 U811 ( .A1(n1119), .A2(n1120), .ZN(n1114) );
NAND3_X1 U812 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1120) );
XNOR2_X1 U813 ( .A(KEYINPUT36), .B(n1124), .ZN(n1123) );
NAND2_X1 U814 ( .A1(G953), .A2(n1125), .ZN(n1122) );
NAND2_X1 U815 ( .A1(n1126), .A2(n1104), .ZN(n1121) );
NAND3_X1 U816 ( .A1(n1126), .A2(n1104), .A3(n1127), .ZN(n1119) );
XOR2_X1 U817 ( .A(KEYINPUT36), .B(n1124), .Z(n1127) );
NAND2_X1 U818 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NOR2_X1 U819 ( .A1(n1130), .A2(n1131), .ZN(G66) );
XOR2_X1 U820 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U821 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
NOR2_X1 U822 ( .A1(n1130), .A2(n1136), .ZN(G63) );
XOR2_X1 U823 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U824 ( .A1(n1134), .A2(G478), .ZN(n1137) );
NOR2_X1 U825 ( .A1(n1130), .A2(n1139), .ZN(G60) );
XOR2_X1 U826 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U827 ( .A1(n1134), .A2(G475), .ZN(n1140) );
XOR2_X1 U828 ( .A(n1142), .B(n1143), .Z(G6) );
NOR2_X1 U829 ( .A1(n1144), .A2(n1145), .ZN(G57) );
XOR2_X1 U830 ( .A(KEYINPUT35), .B(n1130), .Z(n1145) );
XNOR2_X1 U831 ( .A(n1146), .B(n1147), .ZN(n1144) );
XOR2_X1 U832 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U833 ( .A1(n1134), .A2(G472), .ZN(n1149) );
NAND2_X1 U834 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
NOR2_X1 U835 ( .A1(n1130), .A2(n1152), .ZN(G54) );
XOR2_X1 U836 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U837 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND2_X1 U838 ( .A1(KEYINPUT59), .A2(n1157), .ZN(n1156) );
NAND2_X1 U839 ( .A1(n1134), .A2(G469), .ZN(n1155) );
XOR2_X1 U840 ( .A(n1158), .B(n1159), .Z(n1153) );
NOR2_X1 U841 ( .A1(n1130), .A2(n1160), .ZN(G51) );
XOR2_X1 U842 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U843 ( .A(n1163), .B(n1164), .Z(n1162) );
NAND2_X1 U844 ( .A1(n1134), .A2(n1086), .ZN(n1164) );
AND2_X1 U845 ( .A1(n1165), .A2(n1040), .ZN(n1134) );
NAND4_X1 U846 ( .A1(n1166), .A2(n1128), .A3(n1106), .A4(n1108), .ZN(n1040) );
AND4_X1 U847 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1106) );
AND4_X1 U848 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1170) );
NAND2_X1 U849 ( .A1(n1175), .A2(n1176), .ZN(n1169) );
NAND2_X1 U850 ( .A1(n1177), .A2(n1062), .ZN(n1167) );
AND4_X1 U851 ( .A1(n1143), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1128) );
AND4_X1 U852 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1180) );
NAND2_X1 U853 ( .A1(n1185), .A2(n1062), .ZN(n1179) );
XOR2_X1 U854 ( .A(n1186), .B(KEYINPUT40), .Z(n1185) );
NAND4_X1 U855 ( .A1(n1187), .A2(n1026), .A3(n1188), .A4(n1030), .ZN(n1178) );
NOR2_X1 U856 ( .A1(n1189), .A2(n1029), .ZN(n1188) );
XOR2_X1 U857 ( .A(n1035), .B(KEYINPUT11), .Z(n1187) );
NAND4_X1 U858 ( .A1(n1032), .A2(n1056), .A3(n1026), .A4(n1190), .ZN(n1143) );
XOR2_X1 U859 ( .A(n1129), .B(KEYINPUT28), .Z(n1166) );
XOR2_X1 U860 ( .A(n1191), .B(KEYINPUT46), .Z(n1165) );
NOR2_X1 U861 ( .A1(n1192), .A2(n1193), .ZN(n1161) );
NOR2_X1 U862 ( .A1(n1103), .A2(n1194), .ZN(n1193) );
XOR2_X1 U863 ( .A(KEYINPUT27), .B(n1195), .Z(n1194) );
AND2_X1 U864 ( .A1(n1103), .A2(n1195), .ZN(n1192) );
XNOR2_X1 U865 ( .A(n1196), .B(n1197), .ZN(n1195) );
NOR2_X1 U866 ( .A1(KEYINPUT7), .A2(n1124), .ZN(n1197) );
NOR2_X1 U867 ( .A1(n1104), .A2(G952), .ZN(n1130) );
XNOR2_X1 U868 ( .A(n1168), .B(n1198), .ZN(G48) );
XOR2_X1 U869 ( .A(KEYINPUT29), .B(G146), .Z(n1198) );
NAND3_X1 U870 ( .A1(n1056), .A2(n1062), .A3(n1199), .ZN(n1168) );
XNOR2_X1 U871 ( .A(G143), .B(n1174), .ZN(G45) );
NAND4_X1 U872 ( .A1(n1176), .A2(n1200), .A3(n1062), .A4(n1201), .ZN(n1174) );
XNOR2_X1 U873 ( .A(G140), .B(n1173), .ZN(G42) );
NAND3_X1 U874 ( .A1(n1068), .A2(n1026), .A3(n1175), .ZN(n1173) );
INV_X1 U875 ( .A(n1202), .ZN(n1175) );
XOR2_X1 U876 ( .A(n1203), .B(n1172), .Z(G39) );
NAND3_X1 U877 ( .A1(n1066), .A2(n1085), .A3(n1199), .ZN(n1172) );
XNOR2_X1 U878 ( .A(G134), .B(n1171), .ZN(G36) );
NAND4_X1 U879 ( .A1(n1066), .A2(n1176), .A3(n1030), .A4(n1201), .ZN(n1171) );
XOR2_X1 U880 ( .A(G131), .B(n1204), .Z(G33) );
NOR3_X1 U881 ( .A1(n1202), .A2(n1205), .A3(n1206), .ZN(n1204) );
XOR2_X1 U882 ( .A(n1207), .B(KEYINPUT30), .Z(n1205) );
NAND3_X1 U883 ( .A1(n1056), .A2(n1201), .A3(n1066), .ZN(n1202) );
NOR2_X1 U884 ( .A1(n1063), .A2(n1071), .ZN(n1066) );
INV_X1 U885 ( .A(n1064), .ZN(n1071) );
XOR2_X1 U886 ( .A(G128), .B(n1208), .Z(G30) );
NOR2_X1 U887 ( .A1(n1035), .A2(n1209), .ZN(n1208) );
XOR2_X1 U888 ( .A(KEYINPUT58), .B(n1177), .Z(n1209) );
AND2_X1 U889 ( .A1(n1199), .A2(n1030), .ZN(n1177) );
NOR4_X1 U890 ( .A1(n1207), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1199) );
XOR2_X1 U891 ( .A(n1213), .B(n1129), .Z(G3) );
NAND2_X1 U892 ( .A1(n1176), .A2(n1214), .ZN(n1129) );
NOR2_X1 U893 ( .A1(n1206), .A2(n1207), .ZN(n1176) );
XOR2_X1 U894 ( .A(n1215), .B(G125), .Z(G27) );
NAND2_X1 U895 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND3_X1 U896 ( .A1(n1212), .A2(n1218), .A3(n1219), .ZN(n1217) );
INV_X1 U897 ( .A(n1201), .ZN(n1212) );
OR2_X1 U898 ( .A1(n1108), .A2(n1219), .ZN(n1216) );
INV_X1 U899 ( .A(KEYINPUT34), .ZN(n1219) );
NAND2_X1 U900 ( .A1(n1218), .A2(n1201), .ZN(n1108) );
NAND2_X1 U901 ( .A1(n1042), .A2(n1220), .ZN(n1201) );
NAND4_X1 U902 ( .A1(G953), .A2(G902), .A3(n1221), .A4(n1222), .ZN(n1220) );
INV_X1 U903 ( .A(G900), .ZN(n1222) );
AND4_X1 U904 ( .A1(n1068), .A2(n1056), .A3(n1074), .A4(n1062), .ZN(n1218) );
INV_X1 U905 ( .A(n1035), .ZN(n1062) );
XOR2_X1 U906 ( .A(G122), .B(n1223), .Z(G24) );
NOR2_X1 U907 ( .A1(n1035), .A2(n1186), .ZN(n1223) );
NAND4_X1 U908 ( .A1(n1200), .A2(n1074), .A3(n1190), .A4(n1034), .ZN(n1186) );
INV_X1 U909 ( .A(n1029), .ZN(n1190) );
NAND2_X1 U910 ( .A1(n1211), .A2(n1210), .ZN(n1029) );
AND2_X1 U911 ( .A1(n1224), .A2(n1225), .ZN(n1200) );
XOR2_X1 U912 ( .A(n1226), .B(KEYINPUT53), .Z(n1224) );
XOR2_X1 U913 ( .A(n1227), .B(n1184), .Z(G21) );
NAND4_X1 U914 ( .A1(n1214), .A2(n1074), .A3(n1073), .A4(n1084), .ZN(n1184) );
INV_X1 U915 ( .A(n1211), .ZN(n1084) );
XOR2_X1 U916 ( .A(n1183), .B(n1228), .Z(G18) );
NAND2_X1 U917 ( .A1(KEYINPUT52), .A2(G116), .ZN(n1228) );
NAND4_X1 U918 ( .A1(n1032), .A2(n1067), .A3(n1074), .A4(n1030), .ZN(n1183) );
NOR2_X1 U919 ( .A1(n1225), .A2(n1226), .ZN(n1030) );
XOR2_X1 U920 ( .A(n1229), .B(n1230), .Z(G15) );
XOR2_X1 U921 ( .A(KEYINPUT16), .B(G113), .Z(n1230) );
NOR2_X1 U922 ( .A1(KEYINPUT62), .A2(n1181), .ZN(n1229) );
NAND4_X1 U923 ( .A1(n1032), .A2(n1067), .A3(n1056), .A4(n1074), .ZN(n1181) );
NOR2_X1 U924 ( .A1(n1052), .A2(n1231), .ZN(n1074) );
INV_X1 U925 ( .A(n1053), .ZN(n1231) );
AND2_X1 U926 ( .A1(n1226), .A2(n1225), .ZN(n1056) );
INV_X1 U927 ( .A(n1206), .ZN(n1067) );
NAND2_X1 U928 ( .A1(n1211), .A2(n1073), .ZN(n1206) );
XNOR2_X1 U929 ( .A(G110), .B(n1182), .ZN(G12) );
NAND3_X1 U930 ( .A1(n1068), .A2(n1026), .A3(n1214), .ZN(n1182) );
AND2_X1 U931 ( .A1(n1032), .A2(n1085), .ZN(n1214) );
NOR2_X1 U932 ( .A1(n1232), .A2(n1225), .ZN(n1085) );
XNOR2_X1 U933 ( .A(n1233), .B(G475), .ZN(n1225) );
NAND2_X1 U934 ( .A1(n1141), .A2(n1191), .ZN(n1233) );
XOR2_X1 U935 ( .A(n1234), .B(n1235), .Z(n1141) );
XOR2_X1 U936 ( .A(n1236), .B(n1237), .Z(n1235) );
AND3_X1 U937 ( .A1(G214), .A2(n1104), .A3(n1238), .ZN(n1236) );
XOR2_X1 U938 ( .A(n1239), .B(n1240), .Z(n1234) );
NOR3_X1 U939 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1240) );
NOR2_X1 U940 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
INV_X1 U941 ( .A(KEYINPUT5), .ZN(n1245) );
NOR2_X1 U942 ( .A1(n1246), .A2(n1247), .ZN(n1244) );
AND3_X1 U943 ( .A1(KEYINPUT12), .A2(n1103), .A3(n1248), .ZN(n1247) );
NOR2_X1 U944 ( .A1(KEYINPUT12), .A2(n1248), .ZN(n1246) );
NOR2_X1 U945 ( .A1(KEYINPUT5), .A2(n1249), .ZN(n1242) );
NOR2_X1 U946 ( .A1(G125), .A2(n1250), .ZN(n1249) );
XOR2_X1 U947 ( .A(KEYINPUT12), .B(n1248), .Z(n1250) );
NOR2_X1 U948 ( .A1(n1248), .A2(n1103), .ZN(n1241) );
XOR2_X1 U949 ( .A(KEYINPUT0), .B(G140), .Z(n1248) );
NAND2_X1 U950 ( .A1(n1251), .A2(n1252), .ZN(n1239) );
NAND2_X1 U951 ( .A1(n1253), .A2(n1142), .ZN(n1252) );
XOR2_X1 U952 ( .A(KEYINPUT18), .B(n1254), .Z(n1251) );
NOR2_X1 U953 ( .A1(n1142), .A2(n1253), .ZN(n1254) );
XOR2_X1 U954 ( .A(G113), .B(n1255), .Z(n1253) );
NOR2_X1 U955 ( .A1(KEYINPUT9), .A2(n1256), .ZN(n1255) );
XOR2_X1 U956 ( .A(n1257), .B(KEYINPUT15), .Z(n1256) );
INV_X1 U957 ( .A(G122), .ZN(n1257) );
INV_X1 U958 ( .A(n1226), .ZN(n1232) );
XOR2_X1 U959 ( .A(n1258), .B(G478), .Z(n1226) );
NAND2_X1 U960 ( .A1(n1138), .A2(n1191), .ZN(n1258) );
XOR2_X1 U961 ( .A(n1259), .B(n1260), .Z(n1138) );
XOR2_X1 U962 ( .A(G116), .B(n1261), .Z(n1260) );
XOR2_X1 U963 ( .A(KEYINPUT48), .B(G122), .Z(n1261) );
XOR2_X1 U964 ( .A(n1262), .B(n1263), .Z(n1259) );
XNOR2_X1 U965 ( .A(n1264), .B(n1265), .ZN(n1263) );
NOR2_X1 U966 ( .A1(G107), .A2(KEYINPUT24), .ZN(n1265) );
NAND2_X1 U967 ( .A1(n1266), .A2(KEYINPUT61), .ZN(n1264) );
XOR2_X1 U968 ( .A(n1267), .B(n1268), .Z(n1266) );
NOR2_X1 U969 ( .A1(KEYINPUT23), .A2(n1269), .ZN(n1268) );
XNOR2_X1 U970 ( .A(G134), .B(G143), .ZN(n1267) );
NAND2_X1 U971 ( .A1(G217), .A2(n1270), .ZN(n1262) );
NOR2_X1 U972 ( .A1(n1035), .A2(n1189), .ZN(n1032) );
INV_X1 U973 ( .A(n1034), .ZN(n1189) );
NAND2_X1 U974 ( .A1(n1042), .A2(n1271), .ZN(n1034) );
NAND4_X1 U975 ( .A1(G953), .A2(G902), .A3(n1221), .A4(n1125), .ZN(n1271) );
INV_X1 U976 ( .A(G898), .ZN(n1125) );
NAND3_X1 U977 ( .A1(n1221), .A2(n1104), .A3(G952), .ZN(n1042) );
NAND2_X1 U978 ( .A1(G234), .A2(n1272), .ZN(n1221) );
XOR2_X1 U979 ( .A(KEYINPUT13), .B(G237), .Z(n1272) );
NAND2_X1 U980 ( .A1(n1063), .A2(n1064), .ZN(n1035) );
NAND2_X1 U981 ( .A1(n1273), .A2(n1274), .ZN(n1064) );
XOR2_X1 U982 ( .A(KEYINPUT49), .B(G214), .Z(n1273) );
XOR2_X1 U983 ( .A(n1080), .B(n1275), .Z(n1063) );
NOR2_X1 U984 ( .A1(n1086), .A2(KEYINPUT4), .ZN(n1275) );
INV_X1 U985 ( .A(n1079), .ZN(n1086) );
NAND2_X1 U986 ( .A1(G210), .A2(n1274), .ZN(n1079) );
NAND2_X1 U987 ( .A1(n1238), .A2(n1191), .ZN(n1274) );
NAND2_X1 U988 ( .A1(n1276), .A2(n1191), .ZN(n1080) );
XOR2_X1 U989 ( .A(n1277), .B(n1124), .Z(n1276) );
XNOR2_X1 U990 ( .A(n1278), .B(n1279), .ZN(n1124) );
XOR2_X1 U991 ( .A(n1280), .B(n1281), .Z(n1279) );
NAND2_X1 U992 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U993 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U994 ( .A(n1286), .B(KEYINPUT43), .Z(n1282) );
OR2_X1 U995 ( .A1(n1284), .A2(n1285), .ZN(n1286) );
INV_X1 U996 ( .A(G113), .ZN(n1285) );
XOR2_X1 U997 ( .A(G116), .B(n1287), .Z(n1284) );
NOR2_X1 U998 ( .A1(G119), .A2(KEYINPUT41), .ZN(n1287) );
NAND2_X1 U999 ( .A1(n1288), .A2(n1289), .ZN(n1280) );
NAND2_X1 U1000 ( .A1(G107), .A2(n1290), .ZN(n1289) );
XOR2_X1 U1001 ( .A(n1291), .B(KEYINPUT50), .Z(n1288) );
OR2_X1 U1002 ( .A1(n1290), .A2(G107), .ZN(n1291) );
XNOR2_X1 U1003 ( .A(n1142), .B(KEYINPUT31), .ZN(n1290) );
XOR2_X1 U1004 ( .A(n1213), .B(n1292), .Z(n1278) );
XOR2_X1 U1005 ( .A(G122), .B(G110), .Z(n1292) );
XNOR2_X1 U1006 ( .A(KEYINPUT33), .B(n1293), .ZN(n1277) );
NOR2_X1 U1007 ( .A1(KEYINPUT63), .A2(n1294), .ZN(n1293) );
XOR2_X1 U1008 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U1009 ( .A(n1196), .B(n1163), .ZN(n1296) );
NAND2_X1 U1010 ( .A1(G224), .A2(n1104), .ZN(n1163) );
XOR2_X1 U1011 ( .A(n1269), .B(n1297), .Z(n1196) );
XOR2_X1 U1012 ( .A(n1103), .B(KEYINPUT47), .Z(n1295) );
INV_X1 U1013 ( .A(G125), .ZN(n1103) );
INV_X1 U1014 ( .A(n1207), .ZN(n1026) );
NAND2_X1 U1015 ( .A1(n1052), .A2(n1053), .ZN(n1207) );
NAND2_X1 U1016 ( .A1(G221), .A2(n1298), .ZN(n1053) );
XNOR2_X1 U1017 ( .A(n1299), .B(G469), .ZN(n1052) );
NAND2_X1 U1018 ( .A1(n1300), .A2(n1191), .ZN(n1299) );
XOR2_X1 U1019 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1020 ( .A(n1303), .B(n1157), .Z(n1302) );
XOR2_X1 U1021 ( .A(n1304), .B(n1213), .Z(n1157) );
NAND3_X1 U1022 ( .A1(n1305), .A2(n1306), .A3(KEYINPUT51), .ZN(n1304) );
NAND2_X1 U1023 ( .A1(KEYINPUT14), .A2(n1307), .ZN(n1306) );
XOR2_X1 U1024 ( .A(n1142), .B(G107), .Z(n1307) );
NAND3_X1 U1025 ( .A1(G107), .A2(n1142), .A3(n1308), .ZN(n1305) );
INV_X1 U1026 ( .A(KEYINPUT14), .ZN(n1308) );
INV_X1 U1027 ( .A(G104), .ZN(n1142) );
XOR2_X1 U1028 ( .A(n1158), .B(n1309), .Z(n1303) );
NOR2_X1 U1029 ( .A1(KEYINPUT22), .A2(n1159), .ZN(n1309) );
XNOR2_X1 U1030 ( .A(n1310), .B(n1311), .ZN(n1159) );
XOR2_X1 U1031 ( .A(n1312), .B(n1313), .Z(n1158) );
XOR2_X1 U1032 ( .A(n1297), .B(n1314), .Z(n1313) );
XOR2_X1 U1033 ( .A(n1101), .B(n1315), .Z(n1312) );
AND2_X1 U1034 ( .A1(n1104), .A2(G227), .ZN(n1315) );
NAND2_X1 U1035 ( .A1(KEYINPUT25), .A2(G128), .ZN(n1101) );
XOR2_X1 U1036 ( .A(n1316), .B(KEYINPUT55), .Z(n1301) );
XNOR2_X1 U1037 ( .A(KEYINPUT60), .B(KEYINPUT56), .ZN(n1316) );
NOR2_X1 U1038 ( .A1(n1073), .A2(n1211), .ZN(n1068) );
XOR2_X1 U1039 ( .A(n1317), .B(n1135), .Z(n1211) );
AND2_X1 U1040 ( .A1(G217), .A2(n1298), .ZN(n1135) );
NAND2_X1 U1041 ( .A1(G234), .A2(n1191), .ZN(n1298) );
NAND2_X1 U1042 ( .A1(n1133), .A2(n1191), .ZN(n1317) );
XNOR2_X1 U1043 ( .A(n1318), .B(n1319), .ZN(n1133) );
XNOR2_X1 U1044 ( .A(n1314), .B(n1320), .ZN(n1319) );
XOR2_X1 U1045 ( .A(n1321), .B(n1322), .Z(n1320) );
NOR2_X1 U1046 ( .A1(KEYINPUT10), .A2(n1323), .ZN(n1322) );
INV_X1 U1047 ( .A(G146), .ZN(n1323) );
NAND2_X1 U1048 ( .A1(n1270), .A2(G221), .ZN(n1321) );
AND2_X1 U1049 ( .A1(G234), .A2(n1104), .ZN(n1270) );
XOR2_X1 U1050 ( .A(G110), .B(G140), .Z(n1314) );
XOR2_X1 U1051 ( .A(n1324), .B(n1325), .Z(n1318) );
XOR2_X1 U1052 ( .A(KEYINPUT0), .B(G125), .Z(n1325) );
XOR2_X1 U1053 ( .A(n1326), .B(n1327), .Z(n1324) );
NOR2_X1 U1054 ( .A1(KEYINPUT39), .A2(n1203), .ZN(n1327) );
NAND4_X1 U1055 ( .A1(n1328), .A2(n1329), .A3(n1330), .A4(n1331), .ZN(n1326) );
NAND3_X1 U1056 ( .A1(KEYINPUT38), .A2(n1332), .A3(n1269), .ZN(n1331) );
XOR2_X1 U1057 ( .A(KEYINPUT42), .B(n1227), .Z(n1332) );
OR2_X1 U1058 ( .A1(n1269), .A2(KEYINPUT38), .ZN(n1330) );
NAND3_X1 U1059 ( .A1(G119), .A2(n1333), .A3(n1334), .ZN(n1329) );
INV_X1 U1060 ( .A(KEYINPUT44), .ZN(n1334) );
OR2_X1 U1061 ( .A1(KEYINPUT42), .A2(G128), .ZN(n1333) );
NAND3_X1 U1062 ( .A1(n1335), .A2(n1227), .A3(KEYINPUT44), .ZN(n1328) );
INV_X1 U1063 ( .A(G119), .ZN(n1227) );
NAND2_X1 U1064 ( .A1(KEYINPUT42), .A2(n1269), .ZN(n1335) );
INV_X1 U1065 ( .A(G128), .ZN(n1269) );
INV_X1 U1066 ( .A(n1210), .ZN(n1073) );
XOR2_X1 U1067 ( .A(n1336), .B(G472), .Z(n1210) );
NAND2_X1 U1068 ( .A1(n1337), .A2(n1191), .ZN(n1336) );
INV_X1 U1069 ( .A(G902), .ZN(n1191) );
XOR2_X1 U1070 ( .A(n1338), .B(n1339), .Z(n1337) );
NOR2_X1 U1071 ( .A1(KEYINPUT45), .A2(n1146), .ZN(n1339) );
XNOR2_X1 U1072 ( .A(n1340), .B(n1341), .ZN(n1146) );
XOR2_X1 U1073 ( .A(G128), .B(G113), .Z(n1341) );
XOR2_X1 U1074 ( .A(n1342), .B(n1102), .Z(n1340) );
XNOR2_X1 U1075 ( .A(n1310), .B(n1237), .ZN(n1102) );
XOR2_X1 U1076 ( .A(n1311), .B(n1297), .Z(n1237) );
XOR2_X1 U1077 ( .A(G143), .B(G146), .Z(n1297) );
XOR2_X1 U1078 ( .A(G131), .B(KEYINPUT19), .Z(n1311) );
XOR2_X1 U1079 ( .A(G134), .B(n1203), .Z(n1310) );
INV_X1 U1080 ( .A(G137), .ZN(n1203) );
NAND2_X1 U1081 ( .A1(KEYINPUT1), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1082 ( .A(G119), .B(G116), .Z(n1343) );
NAND2_X1 U1083 ( .A1(n1344), .A2(n1151), .ZN(n1338) );
NAND4_X1 U1084 ( .A1(G210), .A2(G101), .A3(n1238), .A4(n1104), .ZN(n1151) );
XOR2_X1 U1085 ( .A(n1150), .B(KEYINPUT26), .Z(n1344) );
NAND2_X1 U1086 ( .A1(n1213), .A2(n1345), .ZN(n1150) );
NAND3_X1 U1087 ( .A1(n1238), .A2(n1104), .A3(G210), .ZN(n1345) );
INV_X1 U1088 ( .A(G953), .ZN(n1104) );
INV_X1 U1089 ( .A(G237), .ZN(n1238) );
INV_X1 U1090 ( .A(G101), .ZN(n1213) );
endmodule


