//Key = 1001101010011100100100010010011010101101111100100100010011100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389;

XNOR2_X1 U758 ( .A(G107), .B(n1047), .ZN(G9) );
NOR2_X1 U759 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR2_X1 U760 ( .A1(G952), .A2(n1050), .ZN(n1049) );
NOR3_X1 U761 ( .A1(n1051), .A2(n1052), .A3(n1050), .ZN(n1048) );
NAND2_X1 U762 ( .A1(n1053), .A2(n1054), .ZN(n1050) );
NAND4_X1 U763 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NOR3_X1 U764 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
XOR2_X1 U765 ( .A(n1062), .B(n1063), .Z(n1061) );
XNOR2_X1 U766 ( .A(n1064), .B(KEYINPUT4), .ZN(n1062) );
XOR2_X1 U767 ( .A(n1065), .B(n1066), .Z(n1059) );
XOR2_X1 U768 ( .A(KEYINPUT35), .B(G478), .Z(n1066) );
NAND2_X1 U769 ( .A1(KEYINPUT49), .A2(n1067), .ZN(n1065) );
NOR2_X1 U770 ( .A1(n1068), .A2(n1069), .ZN(n1052) );
NOR2_X1 U771 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U772 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U773 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR2_X1 U774 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR3_X1 U775 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1076) );
NOR3_X1 U776 ( .A1(n1081), .A2(KEYINPUT40), .A3(n1082), .ZN(n1080) );
NOR2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(n1079) );
NOR2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
AND2_X1 U779 ( .A1(n1087), .A2(KEYINPUT40), .ZN(n1085) );
NOR2_X1 U780 ( .A1(n1088), .A2(n1089), .ZN(n1078) );
NOR2_X1 U781 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
AND2_X1 U782 ( .A1(n1092), .A2(KEYINPUT62), .ZN(n1090) );
NOR2_X1 U783 ( .A1(n1093), .A2(n1089), .ZN(n1074) );
NOR2_X1 U784 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NOR2_X1 U785 ( .A1(n1096), .A2(n1084), .ZN(n1095) );
NOR3_X1 U786 ( .A1(n1097), .A2(KEYINPUT62), .A3(n1098), .ZN(n1094) );
INV_X1 U787 ( .A(n1092), .ZN(n1097) );
NOR3_X1 U788 ( .A1(n1084), .A2(n1099), .A3(n1089), .ZN(n1070) );
INV_X1 U789 ( .A(n1056), .ZN(n1089) );
NOR3_X1 U790 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
AND3_X1 U791 ( .A1(n1057), .A2(n1103), .A3(n1060), .ZN(n1102) );
NOR3_X1 U792 ( .A1(n1104), .A2(n1077), .A3(n1105), .ZN(n1101) );
INV_X1 U793 ( .A(n1098), .ZN(n1077) );
NOR2_X1 U794 ( .A1(n1106), .A2(n1107), .ZN(n1100) );
XOR2_X1 U795 ( .A(n1098), .B(KEYINPUT11), .Z(n1107) );
INV_X1 U796 ( .A(n1081), .ZN(n1084) );
NAND2_X1 U797 ( .A1(n1108), .A2(n1109), .ZN(G72) );
NAND2_X1 U798 ( .A1(n1110), .A2(n1053), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U800 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
OR2_X1 U801 ( .A1(n1113), .A2(n1115), .ZN(n1111) );
NAND4_X1 U802 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1113) );
NOR2_X1 U803 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U804 ( .A(n1122), .B(KEYINPUT3), .Z(n1121) );
XNOR2_X1 U805 ( .A(n1123), .B(KEYINPUT15), .ZN(n1120) );
NAND2_X1 U806 ( .A1(n1124), .A2(G953), .ZN(n1108) );
XOR2_X1 U807 ( .A(n1125), .B(n1115), .Z(n1124) );
XNOR2_X1 U808 ( .A(n1114), .B(KEYINPUT41), .ZN(n1115) );
NAND2_X1 U809 ( .A1(n1126), .A2(n1127), .ZN(n1114) );
NAND2_X1 U810 ( .A1(G953), .A2(n1128), .ZN(n1127) );
XOR2_X1 U811 ( .A(n1129), .B(n1130), .Z(n1126) );
NOR2_X1 U812 ( .A1(KEYINPUT31), .A2(n1131), .ZN(n1129) );
XNOR2_X1 U813 ( .A(n1132), .B(n1133), .ZN(n1131) );
NOR3_X1 U814 ( .A1(KEYINPUT17), .A2(n1134), .A3(n1135), .ZN(n1133) );
NOR3_X1 U815 ( .A1(G131), .A2(n1136), .A3(n1137), .ZN(n1135) );
NOR2_X1 U816 ( .A1(n1138), .A2(n1139), .ZN(n1134) );
NOR2_X1 U817 ( .A1(n1136), .A2(n1137), .ZN(n1138) );
INV_X1 U818 ( .A(n1140), .ZN(n1137) );
AND2_X1 U819 ( .A1(G227), .A2(G900), .ZN(n1125) );
NAND2_X1 U820 ( .A1(n1141), .A2(n1142), .ZN(G69) );
NAND2_X1 U821 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U822 ( .A1(n1145), .A2(n1146), .ZN(n1141) );
NAND2_X1 U823 ( .A1(n1147), .A2(n1144), .ZN(n1146) );
NAND2_X1 U824 ( .A1(G953), .A2(n1148), .ZN(n1144) );
INV_X1 U825 ( .A(G224), .ZN(n1148) );
INV_X1 U826 ( .A(n1143), .ZN(n1145) );
NAND2_X1 U827 ( .A1(n1149), .A2(n1150), .ZN(n1143) );
NAND3_X1 U828 ( .A1(n1151), .A2(n1147), .A3(n1152), .ZN(n1150) );
INV_X1 U829 ( .A(n1153), .ZN(n1147) );
XNOR2_X1 U830 ( .A(n1154), .B(KEYINPUT32), .ZN(n1151) );
OR3_X1 U831 ( .A1(n1154), .A2(G953), .A3(n1152), .ZN(n1149) );
XOR2_X1 U832 ( .A(n1155), .B(n1156), .Z(n1152) );
XOR2_X1 U833 ( .A(G122), .B(G110), .Z(n1156) );
NAND3_X1 U834 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1155) );
NAND2_X1 U835 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U836 ( .A1(KEYINPUT34), .A2(n1162), .ZN(n1161) );
XOR2_X1 U837 ( .A(KEYINPUT60), .B(n1163), .Z(n1162) );
NAND3_X1 U838 ( .A1(KEYINPUT34), .A2(n1164), .A3(n1163), .ZN(n1158) );
OR2_X1 U839 ( .A1(n1163), .A2(KEYINPUT34), .ZN(n1157) );
NOR2_X1 U840 ( .A1(n1165), .A2(n1166), .ZN(G66) );
XOR2_X1 U841 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U842 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
NOR2_X1 U843 ( .A1(n1165), .A2(n1171), .ZN(G63) );
XOR2_X1 U844 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U845 ( .A(KEYINPUT19), .B(n1174), .Z(n1173) );
NOR2_X1 U846 ( .A1(n1175), .A2(n1170), .ZN(n1174) );
NOR2_X1 U847 ( .A1(n1165), .A2(n1176), .ZN(G60) );
XOR2_X1 U848 ( .A(n1177), .B(n1178), .Z(n1176) );
AND2_X1 U849 ( .A1(G475), .A2(n1179), .ZN(n1177) );
XNOR2_X1 U850 ( .A(n1180), .B(n1181), .ZN(G6) );
XNOR2_X1 U851 ( .A(G104), .B(KEYINPUT63), .ZN(n1181) );
NOR2_X1 U852 ( .A1(n1165), .A2(n1182), .ZN(G57) );
XOR2_X1 U853 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND2_X1 U854 ( .A1(n1185), .A2(n1186), .ZN(n1183) );
NAND2_X1 U855 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U856 ( .A(KEYINPUT39), .B(n1189), .Z(n1185) );
NOR2_X1 U857 ( .A1(n1187), .A2(n1188), .ZN(n1189) );
NAND2_X1 U858 ( .A1(n1179), .A2(G472), .ZN(n1188) );
XOR2_X1 U859 ( .A(n1190), .B(n1191), .Z(n1187) );
XOR2_X1 U860 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U861 ( .A(n1194), .B(KEYINPUT1), .Z(n1190) );
NOR2_X1 U862 ( .A1(n1165), .A2(n1195), .ZN(G54) );
XOR2_X1 U863 ( .A(n1196), .B(n1197), .Z(n1195) );
XOR2_X1 U864 ( .A(n1198), .B(n1199), .Z(n1197) );
NOR2_X1 U865 ( .A1(KEYINPUT44), .A2(n1200), .ZN(n1199) );
XOR2_X1 U866 ( .A(KEYINPUT36), .B(n1201), .Z(n1200) );
NOR2_X1 U867 ( .A1(n1202), .A2(n1203), .ZN(n1198) );
NOR2_X1 U868 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
XOR2_X1 U869 ( .A(KEYINPUT0), .B(n1206), .Z(n1205) );
INV_X1 U870 ( .A(n1207), .ZN(n1204) );
XOR2_X1 U871 ( .A(n1192), .B(n1208), .Z(n1196) );
AND2_X1 U872 ( .A1(G469), .A2(n1179), .ZN(n1208) );
INV_X1 U873 ( .A(n1170), .ZN(n1179) );
NOR2_X1 U874 ( .A1(n1165), .A2(n1209), .ZN(G51) );
XOR2_X1 U875 ( .A(n1210), .B(n1211), .Z(n1209) );
NOR2_X1 U876 ( .A1(n1212), .A2(n1170), .ZN(n1211) );
NAND2_X1 U877 ( .A1(G902), .A2(n1051), .ZN(n1170) );
NAND4_X1 U878 ( .A1(n1123), .A2(n1118), .A3(n1154), .A4(n1213), .ZN(n1051) );
AND3_X1 U879 ( .A1(n1116), .A2(n1117), .A3(n1122), .ZN(n1213) );
AND4_X1 U880 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1154) );
AND4_X1 U881 ( .A1(n1047), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1217) );
NAND3_X1 U882 ( .A1(n1056), .A2(n1221), .A3(n1091), .ZN(n1047) );
NOR2_X1 U883 ( .A1(n1222), .A2(n1180), .ZN(n1216) );
AND3_X1 U884 ( .A1(n1056), .A2(n1221), .A3(n1092), .ZN(n1180) );
AND4_X1 U885 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1123) );
NAND2_X1 U886 ( .A1(n1227), .A2(n1228), .ZN(n1223) );
INV_X1 U887 ( .A(n1229), .ZN(n1228) );
XOR2_X1 U888 ( .A(n1230), .B(KEYINPUT59), .Z(n1227) );
NAND2_X1 U889 ( .A1(KEYINPUT6), .A2(n1231), .ZN(n1210) );
XOR2_X1 U890 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U891 ( .A(n1234), .B(n1235), .Z(n1233) );
NOR2_X1 U892 ( .A1(KEYINPUT51), .A2(n1236), .ZN(n1235) );
XOR2_X1 U893 ( .A(G125), .B(n1237), .Z(n1236) );
NOR2_X1 U894 ( .A1(n1053), .A2(G952), .ZN(n1165) );
NAND2_X1 U895 ( .A1(n1238), .A2(n1239), .ZN(G48) );
NAND2_X1 U896 ( .A1(G146), .A2(n1224), .ZN(n1239) );
XOR2_X1 U897 ( .A(KEYINPUT12), .B(n1240), .Z(n1238) );
NOR2_X1 U898 ( .A1(G146), .A2(n1224), .ZN(n1240) );
NAND3_X1 U899 ( .A1(n1092), .A2(n1241), .A3(n1242), .ZN(n1224) );
NAND3_X1 U900 ( .A1(n1243), .A2(n1244), .A3(n1245), .ZN(G45) );
NAND2_X1 U901 ( .A1(G143), .A2(n1225), .ZN(n1245) );
NAND2_X1 U902 ( .A1(KEYINPUT2), .A2(n1246), .ZN(n1244) );
NAND2_X1 U903 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
INV_X1 U904 ( .A(n1225), .ZN(n1248) );
XOR2_X1 U905 ( .A(KEYINPUT28), .B(n1249), .Z(n1247) );
NAND2_X1 U906 ( .A1(n1250), .A2(n1251), .ZN(n1243) );
INV_X1 U907 ( .A(KEYINPUT2), .ZN(n1251) );
NAND2_X1 U908 ( .A1(n1252), .A2(n1253), .ZN(n1250) );
OR3_X1 U909 ( .A1(n1225), .A2(G143), .A3(KEYINPUT28), .ZN(n1253) );
NAND4_X1 U910 ( .A1(n1254), .A2(n1241), .A3(n1255), .A4(n1256), .ZN(n1225) );
NAND2_X1 U911 ( .A1(KEYINPUT28), .A2(G143), .ZN(n1252) );
XOR2_X1 U912 ( .A(G140), .B(n1257), .Z(G42) );
NOR2_X1 U913 ( .A1(n1258), .A2(n1229), .ZN(n1257) );
NAND4_X1 U914 ( .A1(n1086), .A2(n1092), .A3(n1259), .A4(n1098), .ZN(n1229) );
XNOR2_X1 U915 ( .A(n1226), .B(n1260), .ZN(G39) );
NOR2_X1 U916 ( .A1(KEYINPUT5), .A2(n1261), .ZN(n1260) );
INV_X1 U917 ( .A(G137), .ZN(n1261) );
NAND3_X1 U918 ( .A1(n1081), .A2(n1098), .A3(n1242), .ZN(n1226) );
XOR2_X1 U919 ( .A(n1262), .B(n1118), .Z(G36) );
NAND3_X1 U920 ( .A1(n1091), .A2(n1098), .A3(n1254), .ZN(n1118) );
NAND2_X1 U921 ( .A1(n1263), .A2(n1264), .ZN(G33) );
NAND2_X1 U922 ( .A1(G131), .A2(n1265), .ZN(n1264) );
NAND2_X1 U923 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NAND2_X1 U924 ( .A1(KEYINPUT55), .A2(KEYINPUT43), .ZN(n1267) );
NAND3_X1 U925 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1263) );
INV_X1 U926 ( .A(KEYINPUT55), .ZN(n1270) );
OR2_X1 U927 ( .A1(n1116), .A2(KEYINPUT43), .ZN(n1269) );
NAND2_X1 U928 ( .A1(KEYINPUT43), .A2(n1271), .ZN(n1268) );
NAND2_X1 U929 ( .A1(n1266), .A2(n1139), .ZN(n1271) );
INV_X1 U930 ( .A(n1116), .ZN(n1266) );
NAND3_X1 U931 ( .A1(n1092), .A2(n1098), .A3(n1254), .ZN(n1116) );
NOR3_X1 U932 ( .A1(n1106), .A2(n1258), .A3(n1082), .ZN(n1254) );
NAND2_X1 U933 ( .A1(n1272), .A2(n1273), .ZN(n1098) );
OR2_X1 U934 ( .A1(n1096), .A2(KEYINPUT29), .ZN(n1273) );
NAND3_X1 U935 ( .A1(n1274), .A2(n1103), .A3(KEYINPUT29), .ZN(n1272) );
XOR2_X1 U936 ( .A(n1122), .B(n1275), .Z(G30) );
NAND2_X1 U937 ( .A1(KEYINPUT23), .A2(G128), .ZN(n1275) );
NAND3_X1 U938 ( .A1(n1091), .A2(n1241), .A3(n1242), .ZN(n1122) );
AND4_X1 U939 ( .A1(n1259), .A2(n1276), .A3(n1277), .A4(n1230), .ZN(n1242) );
XOR2_X1 U940 ( .A(n1222), .B(n1278), .Z(G3) );
NOR2_X1 U941 ( .A1(KEYINPUT38), .A2(n1279), .ZN(n1278) );
AND3_X1 U942 ( .A1(n1081), .A2(n1221), .A3(n1087), .ZN(n1222) );
XNOR2_X1 U943 ( .A(G125), .B(n1117), .ZN(G27) );
NAND4_X1 U944 ( .A1(n1086), .A2(n1092), .A3(n1280), .A4(n1057), .ZN(n1117) );
NOR2_X1 U945 ( .A1(n1258), .A2(n1096), .ZN(n1280) );
INV_X1 U946 ( .A(n1241), .ZN(n1096) );
INV_X1 U947 ( .A(n1230), .ZN(n1258) );
NAND2_X1 U948 ( .A1(n1069), .A2(n1281), .ZN(n1230) );
NAND4_X1 U949 ( .A1(G902), .A2(G953), .A3(n1282), .A4(n1128), .ZN(n1281) );
INV_X1 U950 ( .A(G900), .ZN(n1128) );
XNOR2_X1 U951 ( .A(G122), .B(n1214), .ZN(G24) );
NAND4_X1 U952 ( .A1(n1283), .A2(n1056), .A3(n1255), .A4(n1256), .ZN(n1214) );
NOR2_X1 U953 ( .A1(n1277), .A2(n1276), .ZN(n1056) );
XNOR2_X1 U954 ( .A(G119), .B(n1215), .ZN(G21) );
NAND4_X1 U955 ( .A1(n1283), .A2(n1081), .A3(n1276), .A4(n1277), .ZN(n1215) );
INV_X1 U956 ( .A(n1284), .ZN(n1276) );
XOR2_X1 U957 ( .A(n1220), .B(n1285), .Z(G18) );
NAND2_X1 U958 ( .A1(KEYINPUT56), .A2(G116), .ZN(n1285) );
NAND3_X1 U959 ( .A1(n1087), .A2(n1091), .A3(n1283), .ZN(n1220) );
AND2_X1 U960 ( .A1(n1055), .A2(n1255), .ZN(n1091) );
XNOR2_X1 U961 ( .A(G113), .B(n1219), .ZN(G15) );
NAND3_X1 U962 ( .A1(n1087), .A2(n1092), .A3(n1283), .ZN(n1219) );
AND2_X1 U963 ( .A1(n1057), .A2(n1286), .ZN(n1283) );
INV_X1 U964 ( .A(n1073), .ZN(n1057) );
NAND2_X1 U965 ( .A1(n1287), .A2(n1104), .ZN(n1073) );
NOR2_X1 U966 ( .A1(n1255), .A2(n1055), .ZN(n1092) );
INV_X1 U967 ( .A(n1082), .ZN(n1087) );
NAND2_X1 U968 ( .A1(n1284), .A2(n1277), .ZN(n1082) );
XOR2_X1 U969 ( .A(n1218), .B(n1288), .Z(G12) );
XOR2_X1 U970 ( .A(KEYINPUT13), .B(G110), .Z(n1288) );
NAND3_X1 U971 ( .A1(n1081), .A2(n1221), .A3(n1086), .ZN(n1218) );
NOR2_X1 U972 ( .A1(n1277), .A2(n1284), .ZN(n1086) );
XNOR2_X1 U973 ( .A(n1289), .B(n1169), .ZN(n1284) );
NAND2_X1 U974 ( .A1(G217), .A2(n1290), .ZN(n1169) );
OR2_X1 U975 ( .A1(n1168), .A2(G902), .ZN(n1289) );
XNOR2_X1 U976 ( .A(n1291), .B(n1292), .ZN(n1168) );
XOR2_X1 U977 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U978 ( .A(n1295), .B(n1296), .Z(n1294) );
AND3_X1 U979 ( .A1(G221), .A2(n1053), .A3(G234), .ZN(n1296) );
NOR2_X1 U980 ( .A1(KEYINPUT48), .A2(G140), .ZN(n1295) );
XOR2_X1 U981 ( .A(n1297), .B(n1298), .Z(n1291) );
XOR2_X1 U982 ( .A(G137), .B(G125), .Z(n1298) );
XNOR2_X1 U983 ( .A(G110), .B(G119), .ZN(n1297) );
XNOR2_X1 U984 ( .A(n1299), .B(G472), .ZN(n1277) );
NAND2_X1 U985 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
XOR2_X1 U986 ( .A(n1302), .B(n1303), .Z(n1300) );
XNOR2_X1 U987 ( .A(n1184), .B(n1193), .ZN(n1303) );
XOR2_X1 U988 ( .A(n1304), .B(n1305), .Z(n1193) );
NOR2_X1 U989 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NOR3_X1 U990 ( .A1(n1308), .A2(G119), .A3(n1309), .ZN(n1307) );
INV_X1 U991 ( .A(G116), .ZN(n1309) );
INV_X1 U992 ( .A(KEYINPUT50), .ZN(n1308) );
NOR2_X1 U993 ( .A1(KEYINPUT50), .A2(n1310), .ZN(n1306) );
XOR2_X1 U994 ( .A(n1311), .B(n1279), .Z(n1184) );
INV_X1 U995 ( .A(G101), .ZN(n1279) );
NAND2_X1 U996 ( .A1(G210), .A2(n1312), .ZN(n1311) );
XOR2_X1 U997 ( .A(n1237), .B(n1313), .Z(n1302) );
XNOR2_X1 U998 ( .A(n1314), .B(KEYINPUT54), .ZN(n1313) );
NAND2_X1 U999 ( .A1(KEYINPUT37), .A2(n1315), .ZN(n1314) );
AND2_X1 U1000 ( .A1(n1259), .A2(n1286), .ZN(n1221) );
AND2_X1 U1001 ( .A1(n1241), .A2(n1316), .ZN(n1286) );
NAND2_X1 U1002 ( .A1(n1069), .A2(n1317), .ZN(n1316) );
NAND3_X1 U1003 ( .A1(n1153), .A2(n1282), .A3(G902), .ZN(n1317) );
NOR2_X1 U1004 ( .A1(G898), .A2(n1053), .ZN(n1153) );
NAND3_X1 U1005 ( .A1(n1282), .A2(n1053), .A3(G952), .ZN(n1069) );
NAND2_X1 U1006 ( .A1(G237), .A2(G234), .ZN(n1282) );
NOR2_X1 U1007 ( .A1(n1103), .A2(n1060), .ZN(n1241) );
INV_X1 U1008 ( .A(n1274), .ZN(n1060) );
NAND2_X1 U1009 ( .A1(G214), .A2(n1318), .ZN(n1274) );
NAND3_X1 U1010 ( .A1(n1319), .A2(n1320), .A3(n1321), .ZN(n1103) );
NAND2_X1 U1011 ( .A1(n1064), .A2(n1322), .ZN(n1321) );
OR3_X1 U1012 ( .A1(n1322), .A2(n1064), .A3(KEYINPUT22), .ZN(n1320) );
AND2_X1 U1013 ( .A1(n1323), .A2(n1301), .ZN(n1064) );
XOR2_X1 U1014 ( .A(n1324), .B(n1325), .Z(n1323) );
INV_X1 U1015 ( .A(n1232), .ZN(n1325) );
XOR2_X1 U1016 ( .A(n1326), .B(n1327), .Z(n1232) );
XOR2_X1 U1017 ( .A(n1328), .B(n1329), .Z(n1327) );
XOR2_X1 U1018 ( .A(KEYINPUT16), .B(G110), .Z(n1329) );
XNOR2_X1 U1019 ( .A(n1330), .B(n1163), .ZN(n1326) );
XNOR2_X1 U1020 ( .A(n1304), .B(n1310), .ZN(n1163) );
XOR2_X1 U1021 ( .A(G116), .B(G119), .Z(n1310) );
XNOR2_X1 U1022 ( .A(G113), .B(KEYINPUT24), .ZN(n1304) );
NOR3_X1 U1023 ( .A1(KEYINPUT14), .A2(n1331), .A3(n1332), .ZN(n1324) );
NOR2_X1 U1024 ( .A1(n1237), .A2(n1333), .ZN(n1332) );
XOR2_X1 U1025 ( .A(KEYINPUT25), .B(n1334), .Z(n1333) );
AND2_X1 U1026 ( .A1(n1237), .A2(n1334), .ZN(n1331) );
XNOR2_X1 U1027 ( .A(n1234), .B(n1335), .ZN(n1334) );
XOR2_X1 U1028 ( .A(KEYINPUT8), .B(G125), .Z(n1335) );
NAND2_X1 U1029 ( .A1(n1336), .A2(n1053), .ZN(n1234) );
XOR2_X1 U1030 ( .A(KEYINPUT9), .B(G224), .Z(n1336) );
INV_X1 U1031 ( .A(n1194), .ZN(n1237) );
XOR2_X1 U1032 ( .A(n1249), .B(n1293), .Z(n1194) );
XOR2_X1 U1033 ( .A(G128), .B(G146), .Z(n1293) );
NAND2_X1 U1034 ( .A1(KEYINPUT53), .A2(n1212), .ZN(n1322) );
NAND2_X1 U1035 ( .A1(KEYINPUT22), .A2(n1063), .ZN(n1319) );
INV_X1 U1036 ( .A(n1212), .ZN(n1063) );
NAND2_X1 U1037 ( .A1(G210), .A2(n1318), .ZN(n1212) );
NAND2_X1 U1038 ( .A1(n1337), .A2(n1301), .ZN(n1318) );
INV_X1 U1039 ( .A(G237), .ZN(n1337) );
INV_X1 U1040 ( .A(n1106), .ZN(n1259) );
NAND2_X1 U1041 ( .A1(n1105), .A2(n1104), .ZN(n1106) );
NAND2_X1 U1042 ( .A1(G221), .A2(n1290), .ZN(n1104) );
NAND2_X1 U1043 ( .A1(G234), .A2(n1301), .ZN(n1290) );
INV_X1 U1044 ( .A(n1287), .ZN(n1105) );
XOR2_X1 U1045 ( .A(n1338), .B(G469), .Z(n1287) );
NAND2_X1 U1046 ( .A1(n1339), .A2(n1301), .ZN(n1338) );
XOR2_X1 U1047 ( .A(n1315), .B(n1340), .Z(n1339) );
XOR2_X1 U1048 ( .A(n1341), .B(n1201), .Z(n1340) );
XNOR2_X1 U1049 ( .A(n1342), .B(n1343), .ZN(n1201) );
NOR2_X1 U1050 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
NOR3_X1 U1051 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1345) );
XNOR2_X1 U1052 ( .A(G104), .B(G107), .ZN(n1348) );
INV_X1 U1053 ( .A(KEYINPUT61), .ZN(n1346) );
NOR2_X1 U1054 ( .A1(KEYINPUT61), .A2(n1160), .ZN(n1344) );
INV_X1 U1055 ( .A(n1164), .ZN(n1160) );
XOR2_X1 U1056 ( .A(n1328), .B(G104), .Z(n1164) );
XNOR2_X1 U1057 ( .A(G107), .B(n1347), .ZN(n1328) );
XNOR2_X1 U1058 ( .A(G101), .B(KEYINPUT27), .ZN(n1347) );
XOR2_X1 U1059 ( .A(n1132), .B(KEYINPUT18), .Z(n1342) );
NAND2_X1 U1060 ( .A1(n1349), .A2(n1350), .ZN(n1132) );
NAND4_X1 U1061 ( .A1(KEYINPUT30), .A2(G146), .A3(n1351), .A4(n1352), .ZN(n1350) );
NAND2_X1 U1062 ( .A1(n1353), .A2(n1249), .ZN(n1352) );
NAND2_X1 U1063 ( .A1(n1354), .A2(G143), .ZN(n1351) );
NAND3_X1 U1064 ( .A1(n1355), .A2(n1356), .A3(n1357), .ZN(n1349) );
NAND2_X1 U1065 ( .A1(KEYINPUT30), .A2(G146), .ZN(n1357) );
NAND2_X1 U1066 ( .A1(n1353), .A2(G143), .ZN(n1356) );
XOR2_X1 U1067 ( .A(G128), .B(KEYINPUT57), .Z(n1353) );
NAND2_X1 U1068 ( .A1(n1354), .A2(n1249), .ZN(n1355) );
XOR2_X1 U1069 ( .A(n1358), .B(KEYINPUT46), .Z(n1354) );
INV_X1 U1070 ( .A(G128), .ZN(n1358) );
NOR2_X1 U1071 ( .A1(n1202), .A2(n1359), .ZN(n1341) );
XOR2_X1 U1072 ( .A(n1360), .B(KEYINPUT58), .Z(n1359) );
NAND2_X1 U1073 ( .A1(n1206), .A2(n1207), .ZN(n1360) );
NOR2_X1 U1074 ( .A1(n1207), .A2(n1206), .ZN(n1202) );
XOR2_X1 U1075 ( .A(G110), .B(G140), .Z(n1206) );
NAND2_X1 U1076 ( .A1(G227), .A2(n1053), .ZN(n1207) );
INV_X1 U1077 ( .A(n1192), .ZN(n1315) );
XOR2_X1 U1078 ( .A(n1361), .B(n1362), .Z(n1192) );
NOR2_X1 U1079 ( .A1(G131), .A2(KEYINPUT21), .ZN(n1362) );
XOR2_X1 U1080 ( .A(n1363), .B(KEYINPUT20), .Z(n1361) );
NAND3_X1 U1081 ( .A1(n1364), .A2(n1365), .A3(n1140), .ZN(n1363) );
NAND2_X1 U1082 ( .A1(G137), .A2(n1262), .ZN(n1140) );
NAND2_X1 U1083 ( .A1(KEYINPUT47), .A2(n1262), .ZN(n1365) );
NAND2_X1 U1084 ( .A1(n1136), .A2(n1366), .ZN(n1364) );
INV_X1 U1085 ( .A(KEYINPUT47), .ZN(n1366) );
NOR2_X1 U1086 ( .A1(n1262), .A2(G137), .ZN(n1136) );
INV_X1 U1087 ( .A(G134), .ZN(n1262) );
NOR2_X1 U1088 ( .A1(n1255), .A2(n1256), .ZN(n1081) );
INV_X1 U1089 ( .A(n1055), .ZN(n1256) );
XOR2_X1 U1090 ( .A(n1367), .B(G475), .Z(n1055) );
OR2_X1 U1091 ( .A1(n1178), .A2(G902), .ZN(n1367) );
XNOR2_X1 U1092 ( .A(n1368), .B(n1369), .ZN(n1178) );
XOR2_X1 U1093 ( .A(n1370), .B(n1330), .Z(n1369) );
XOR2_X1 U1094 ( .A(G104), .B(G122), .Z(n1330) );
NOR2_X1 U1095 ( .A1(KEYINPUT45), .A2(n1371), .ZN(n1370) );
XOR2_X1 U1096 ( .A(n1249), .B(n1372), .Z(n1371) );
NAND2_X1 U1097 ( .A1(G214), .A2(n1312), .ZN(n1372) );
NOR2_X1 U1098 ( .A1(G953), .A2(G237), .ZN(n1312) );
XOR2_X1 U1099 ( .A(n1373), .B(n1374), .Z(n1368) );
NOR2_X1 U1100 ( .A1(KEYINPUT10), .A2(n1375), .ZN(n1374) );
XNOR2_X1 U1101 ( .A(G146), .B(n1130), .ZN(n1375) );
XOR2_X1 U1102 ( .A(G125), .B(G140), .Z(n1130) );
XOR2_X1 U1103 ( .A(G113), .B(n1139), .Z(n1373) );
INV_X1 U1104 ( .A(G131), .ZN(n1139) );
XOR2_X1 U1105 ( .A(n1175), .B(n1067), .Z(n1255) );
NAND2_X1 U1106 ( .A1(n1376), .A2(n1301), .ZN(n1067) );
INV_X1 U1107 ( .A(G902), .ZN(n1301) );
XNOR2_X1 U1108 ( .A(KEYINPUT42), .B(n1172), .ZN(n1376) );
NAND2_X1 U1109 ( .A1(n1377), .A2(n1378), .ZN(n1172) );
NAND4_X1 U1110 ( .A1(G234), .A2(G217), .A3(n1379), .A4(n1053), .ZN(n1378) );
XOR2_X1 U1111 ( .A(n1380), .B(KEYINPUT52), .Z(n1377) );
NAND2_X1 U1112 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
NAND3_X1 U1113 ( .A1(G217), .A2(n1053), .A3(G234), .ZN(n1382) );
INV_X1 U1114 ( .A(G953), .ZN(n1053) );
INV_X1 U1115 ( .A(n1379), .ZN(n1381) );
XOR2_X1 U1116 ( .A(n1383), .B(n1384), .Z(n1379) );
XOR2_X1 U1117 ( .A(G122), .B(n1385), .Z(n1384) );
XOR2_X1 U1118 ( .A(KEYINPUT33), .B(G134), .Z(n1385) );
XOR2_X1 U1119 ( .A(n1386), .B(n1387), .Z(n1383) );
XOR2_X1 U1120 ( .A(G116), .B(G107), .Z(n1387) );
NAND2_X1 U1121 ( .A1(n1388), .A2(KEYINPUT26), .ZN(n1386) );
XOR2_X1 U1122 ( .A(n1249), .B(n1389), .Z(n1388) );
NOR2_X1 U1123 ( .A1(G128), .A2(KEYINPUT7), .ZN(n1389) );
INV_X1 U1124 ( .A(G143), .ZN(n1249) );
INV_X1 U1125 ( .A(G478), .ZN(n1175) );
endmodule


