//Key = 1011010100111100010001111010000001010101000110010101101011111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341;

NAND2_X1 U743 ( .A1(n1030), .A2(n1031), .ZN(G9) );
NAND2_X1 U744 ( .A1(G107), .A2(n1032), .ZN(n1031) );
XOR2_X1 U745 ( .A(KEYINPUT13), .B(n1033), .Z(n1030) );
NOR2_X1 U746 ( .A1(G107), .A2(n1032), .ZN(n1033) );
NAND3_X1 U747 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1032) );
NOR2_X1 U748 ( .A1(n1037), .A2(n1038), .ZN(G75) );
NOR4_X1 U749 ( .A1(n1039), .A2(n1040), .A3(G953), .A4(n1041), .ZN(n1038) );
NOR3_X1 U750 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1040) );
NOR2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U752 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U753 ( .A1(n1049), .A2(n1050), .ZN(n1045) );
NOR2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U755 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR2_X1 U756 ( .A1(n1055), .A2(n1056), .ZN(n1051) );
XNOR2_X1 U757 ( .A(KEYINPUT62), .B(n1057), .ZN(n1056) );
NAND3_X1 U758 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1039) );
XOR2_X1 U759 ( .A(n1061), .B(KEYINPUT35), .Z(n1060) );
NAND2_X1 U760 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND3_X1 U761 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
INV_X1 U762 ( .A(n1042), .ZN(n1066) );
NAND3_X1 U763 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1065) );
NAND4_X1 U764 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
XNOR2_X1 U765 ( .A(n1074), .B(KEYINPUT56), .ZN(n1070) );
NAND4_X1 U766 ( .A1(n1075), .A2(n1074), .A3(n1035), .A4(n1076), .ZN(n1068) );
NAND3_X1 U767 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1067) );
NAND2_X1 U768 ( .A1(n1080), .A2(n1034), .ZN(n1062) );
NAND2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(n1059) );
NOR3_X1 U770 ( .A1(n1048), .A2(n1050), .A3(n1042), .ZN(n1080) );
INV_X1 U771 ( .A(n1078), .ZN(n1048) );
NOR2_X1 U772 ( .A1(n1053), .A2(n1057), .ZN(n1078) );
NOR3_X1 U773 ( .A1(n1041), .A2(G953), .A3(G952), .ZN(n1037) );
AND4_X1 U774 ( .A1(n1082), .A2(n1074), .A3(n1083), .A4(n1084), .ZN(n1041) );
NOR4_X1 U775 ( .A1(n1075), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1084) );
XNOR2_X1 U776 ( .A(G478), .B(n1088), .ZN(n1086) );
NOR2_X1 U777 ( .A1(KEYINPUT36), .A2(n1089), .ZN(n1088) );
XNOR2_X1 U778 ( .A(n1090), .B(KEYINPUT2), .ZN(n1089) );
XOR2_X1 U779 ( .A(n1091), .B(n1092), .Z(n1085) );
XOR2_X1 U780 ( .A(KEYINPUT12), .B(G469), .Z(n1092) );
XOR2_X1 U781 ( .A(n1093), .B(KEYINPUT55), .Z(n1083) );
INV_X1 U782 ( .A(n1050), .ZN(n1074) );
XNOR2_X1 U783 ( .A(n1094), .B(n1095), .ZN(n1082) );
XOR2_X1 U784 ( .A(n1096), .B(n1097), .Z(G72) );
NOR2_X1 U785 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U786 ( .A(n1100), .B(KEYINPUT26), .Z(n1098) );
NAND2_X1 U787 ( .A1(G900), .A2(G227), .ZN(n1100) );
NAND2_X1 U788 ( .A1(n1101), .A2(n1102), .ZN(n1096) );
NAND2_X1 U789 ( .A1(n1103), .A2(n1099), .ZN(n1102) );
XOR2_X1 U790 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND3_X1 U791 ( .A1(G900), .A2(n1105), .A3(G953), .ZN(n1101) );
XOR2_X1 U792 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U793 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U794 ( .A(KEYINPUT4), .B(G137), .Z(n1109) );
XOR2_X1 U795 ( .A(KEYINPUT52), .B(KEYINPUT51), .Z(n1108) );
XOR2_X1 U796 ( .A(n1110), .B(n1111), .Z(n1106) );
XOR2_X1 U797 ( .A(G131), .B(n1112), .Z(n1111) );
NOR2_X1 U798 ( .A1(G134), .A2(KEYINPUT1), .ZN(n1112) );
XOR2_X1 U799 ( .A(n1113), .B(n1114), .Z(n1110) );
NAND2_X1 U800 ( .A1(n1115), .A2(n1116), .ZN(G69) );
NAND2_X1 U801 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U802 ( .A1(G953), .A2(n1119), .ZN(n1118) );
NAND3_X1 U803 ( .A1(G953), .A2(n1120), .A3(n1121), .ZN(n1115) );
XNOR2_X1 U804 ( .A(n1117), .B(KEYINPUT14), .ZN(n1121) );
XNOR2_X1 U805 ( .A(n1122), .B(n1123), .ZN(n1117) );
AND2_X1 U806 ( .A1(n1124), .A2(n1099), .ZN(n1123) );
NAND2_X1 U807 ( .A1(n1125), .A2(n1126), .ZN(n1122) );
NAND2_X1 U808 ( .A1(G953), .A2(n1127), .ZN(n1126) );
XOR2_X1 U809 ( .A(n1128), .B(n1129), .Z(n1125) );
XOR2_X1 U810 ( .A(n1130), .B(n1131), .Z(n1128) );
NAND2_X1 U811 ( .A1(KEYINPUT49), .A2(n1132), .ZN(n1130) );
NAND2_X1 U812 ( .A1(G898), .A2(G224), .ZN(n1120) );
NOR2_X1 U813 ( .A1(n1133), .A2(n1134), .ZN(G66) );
NOR3_X1 U814 ( .A1(n1094), .A2(n1135), .A3(n1136), .ZN(n1134) );
AND4_X1 U815 ( .A1(n1137), .A2(KEYINPUT54), .A3(n1095), .A4(n1138), .ZN(n1136) );
NOR2_X1 U816 ( .A1(n1139), .A2(n1137), .ZN(n1135) );
NOR3_X1 U817 ( .A1(n1140), .A2(n1058), .A3(n1141), .ZN(n1139) );
INV_X1 U818 ( .A(KEYINPUT54), .ZN(n1140) );
NOR2_X1 U819 ( .A1(n1133), .A2(n1142), .ZN(G63) );
NOR3_X1 U820 ( .A1(n1090), .A2(n1143), .A3(n1144), .ZN(n1142) );
AND3_X1 U821 ( .A1(n1145), .A2(G478), .A3(n1138), .ZN(n1144) );
NOR2_X1 U822 ( .A1(n1146), .A2(n1145), .ZN(n1143) );
NOR2_X1 U823 ( .A1(n1058), .A2(n1147), .ZN(n1146) );
NOR2_X1 U824 ( .A1(n1133), .A2(n1148), .ZN(G60) );
XOR2_X1 U825 ( .A(n1149), .B(n1150), .Z(n1148) );
NAND2_X1 U826 ( .A1(n1138), .A2(G475), .ZN(n1149) );
XOR2_X1 U827 ( .A(G104), .B(n1151), .Z(G6) );
NOR2_X1 U828 ( .A1(n1133), .A2(n1152), .ZN(G57) );
XOR2_X1 U829 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U830 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U831 ( .A(n1157), .B(n1158), .Z(n1153) );
XOR2_X1 U832 ( .A(n1159), .B(KEYINPUT10), .Z(n1157) );
NAND2_X1 U833 ( .A1(n1138), .A2(G472), .ZN(n1159) );
NOR3_X1 U834 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(G54) );
AND2_X1 U835 ( .A1(KEYINPUT43), .A2(n1133), .ZN(n1162) );
NOR3_X1 U836 ( .A1(KEYINPUT43), .A2(G953), .A3(G952), .ZN(n1161) );
XOR2_X1 U837 ( .A(n1163), .B(n1164), .Z(n1160) );
XOR2_X1 U838 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND2_X1 U839 ( .A1(n1167), .A2(n1168), .ZN(n1165) );
NAND2_X1 U840 ( .A1(n1169), .A2(n1132), .ZN(n1168) );
NAND2_X1 U841 ( .A1(n1170), .A2(n1171), .ZN(n1167) );
XNOR2_X1 U842 ( .A(n1169), .B(KEYINPUT41), .ZN(n1171) );
XOR2_X1 U843 ( .A(n1172), .B(n1173), .Z(n1163) );
NAND3_X1 U844 ( .A1(n1138), .A2(G469), .A3(KEYINPUT33), .ZN(n1172) );
NOR2_X1 U845 ( .A1(n1133), .A2(n1174), .ZN(G51) );
XNOR2_X1 U846 ( .A(n1175), .B(n1176), .ZN(n1174) );
XOR2_X1 U847 ( .A(n1177), .B(n1178), .Z(n1176) );
NAND2_X1 U848 ( .A1(KEYINPUT0), .A2(n1179), .ZN(n1178) );
NAND2_X1 U849 ( .A1(n1138), .A2(G210), .ZN(n1177) );
NOR2_X1 U850 ( .A1(n1180), .A2(n1058), .ZN(n1138) );
NOR2_X1 U851 ( .A1(n1124), .A2(n1104), .ZN(n1058) );
NAND4_X1 U852 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1104) );
NOR4_X1 U853 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1184) );
NOR2_X1 U854 ( .A1(n1189), .A2(n1190), .ZN(n1183) );
NOR4_X1 U855 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1190) );
INV_X1 U856 ( .A(KEYINPUT42), .ZN(n1192) );
NOR2_X1 U857 ( .A1(n1195), .A2(n1047), .ZN(n1189) );
NOR3_X1 U858 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1195) );
NOR3_X1 U859 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1198) );
NOR3_X1 U860 ( .A1(n1194), .A2(KEYINPUT42), .A3(n1193), .ZN(n1196) );
NAND2_X1 U861 ( .A1(n1202), .A2(n1199), .ZN(n1181) );
INV_X1 U862 ( .A(KEYINPUT31), .ZN(n1199) );
NAND2_X1 U863 ( .A1(n1203), .A2(n1204), .ZN(n1124) );
AND4_X1 U864 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
NOR4_X1 U865 ( .A1(n1209), .A2(n1151), .A3(n1210), .A4(n1211), .ZN(n1203) );
NOR3_X1 U866 ( .A1(n1054), .A2(n1193), .A3(n1212), .ZN(n1211) );
NOR3_X1 U867 ( .A1(n1213), .A2(n1214), .A3(n1057), .ZN(n1210) );
XNOR2_X1 U868 ( .A(n1034), .B(KEYINPUT6), .ZN(n1214) );
AND3_X1 U869 ( .A1(n1036), .A2(n1035), .A3(n1081), .ZN(n1151) );
NOR2_X1 U870 ( .A1(n1099), .A2(G952), .ZN(n1133) );
XNOR2_X1 U871 ( .A(G146), .B(n1182), .ZN(G48) );
NAND2_X1 U872 ( .A1(n1215), .A2(n1081), .ZN(n1182) );
XNOR2_X1 U873 ( .A(n1216), .B(n1202), .ZN(G45) );
NOR3_X1 U874 ( .A1(n1047), .A2(n1217), .A3(n1200), .ZN(n1202) );
NAND4_X1 U875 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1200) );
XOR2_X1 U876 ( .A(G140), .B(n1188), .Z(G42) );
AND2_X1 U877 ( .A1(n1222), .A2(n1223), .ZN(n1188) );
XOR2_X1 U878 ( .A(G137), .B(n1187), .Z(G39) );
NOR3_X1 U879 ( .A1(n1050), .A2(n1044), .A3(n1194), .ZN(n1187) );
XNOR2_X1 U880 ( .A(n1224), .B(n1186), .ZN(G36) );
AND3_X1 U881 ( .A1(n1219), .A2(n1034), .A3(n1223), .ZN(n1186) );
XNOR2_X1 U882 ( .A(G131), .B(n1225), .ZN(G33) );
NAND2_X1 U883 ( .A1(KEYINPUT17), .A2(n1185), .ZN(n1225) );
AND3_X1 U884 ( .A1(n1219), .A2(n1081), .A3(n1223), .ZN(n1185) );
NOR3_X1 U885 ( .A1(n1055), .A2(n1217), .A3(n1050), .ZN(n1223) );
NAND2_X1 U886 ( .A1(n1077), .A2(n1226), .ZN(n1050) );
INV_X1 U887 ( .A(n1201), .ZN(n1217) );
INV_X1 U888 ( .A(n1220), .ZN(n1055) );
XNOR2_X1 U889 ( .A(G128), .B(n1227), .ZN(G30) );
NAND2_X1 U890 ( .A1(n1215), .A2(n1034), .ZN(n1227) );
INV_X1 U891 ( .A(n1193), .ZN(n1034) );
NOR2_X1 U892 ( .A1(n1194), .A2(n1047), .ZN(n1215) );
INV_X1 U893 ( .A(n1191), .ZN(n1047) );
NAND4_X1 U894 ( .A1(n1071), .A2(n1220), .A3(n1228), .A4(n1201), .ZN(n1194) );
XOR2_X1 U895 ( .A(G101), .B(n1209), .Z(G3) );
NOR3_X1 U896 ( .A1(n1213), .A2(n1044), .A3(n1054), .ZN(n1209) );
INV_X1 U897 ( .A(n1064), .ZN(n1044) );
NAND2_X1 U898 ( .A1(n1229), .A2(n1230), .ZN(G27) );
NAND2_X1 U899 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XOR2_X1 U900 ( .A(n1233), .B(KEYINPUT34), .Z(n1232) );
XNOR2_X1 U901 ( .A(KEYINPUT21), .B(G125), .ZN(n1231) );
NAND2_X1 U902 ( .A1(n1234), .A2(n1235), .ZN(n1229) );
XNOR2_X1 U903 ( .A(KEYINPUT28), .B(n1233), .ZN(n1235) );
NAND2_X1 U904 ( .A1(n1191), .A2(n1236), .ZN(n1233) );
XOR2_X1 U905 ( .A(KEYINPUT25), .B(n1197), .Z(n1236) );
AND3_X1 U906 ( .A1(n1073), .A2(n1201), .A3(n1222), .ZN(n1197) );
AND3_X1 U907 ( .A1(n1072), .A2(n1081), .A3(n1071), .ZN(n1222) );
NAND2_X1 U908 ( .A1(n1042), .A2(n1237), .ZN(n1201) );
NAND4_X1 U909 ( .A1(G902), .A2(G953), .A3(n1238), .A4(n1239), .ZN(n1237) );
INV_X1 U910 ( .A(G900), .ZN(n1239) );
XOR2_X1 U911 ( .A(KEYINPUT21), .B(G125), .Z(n1234) );
XNOR2_X1 U912 ( .A(G122), .B(n1208), .ZN(G24) );
NAND4_X1 U913 ( .A1(n1218), .A2(n1240), .A3(n1035), .A4(n1221), .ZN(n1208) );
INV_X1 U914 ( .A(n1057), .ZN(n1035) );
NAND2_X1 U915 ( .A1(n1072), .A2(n1241), .ZN(n1057) );
XNOR2_X1 U916 ( .A(G119), .B(n1205), .ZN(G21) );
NAND4_X1 U917 ( .A1(n1071), .A2(n1240), .A3(n1228), .A4(n1064), .ZN(n1205) );
XNOR2_X1 U918 ( .A(n1242), .B(KEYINPUT37), .ZN(n1228) );
XNOR2_X1 U919 ( .A(n1243), .B(n1244), .ZN(G18) );
NOR4_X1 U920 ( .A1(KEYINPUT30), .A2(n1193), .A3(n1212), .A4(n1054), .ZN(n1244) );
NAND2_X1 U921 ( .A1(n1245), .A2(n1221), .ZN(n1193) );
NAND3_X1 U922 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(G15) );
OR2_X1 U923 ( .A1(n1207), .A2(KEYINPUT7), .ZN(n1248) );
NAND3_X1 U924 ( .A1(KEYINPUT7), .A2(n1207), .A3(G113), .ZN(n1247) );
NAND2_X1 U925 ( .A1(n1249), .A2(n1250), .ZN(n1246) );
NAND2_X1 U926 ( .A1(KEYINPUT7), .A2(n1251), .ZN(n1249) );
XNOR2_X1 U927 ( .A(KEYINPUT39), .B(n1207), .ZN(n1251) );
NAND3_X1 U928 ( .A1(n1240), .A2(n1081), .A3(n1219), .ZN(n1207) );
INV_X1 U929 ( .A(n1054), .ZN(n1219) );
NAND2_X1 U930 ( .A1(n1242), .A2(n1241), .ZN(n1054) );
XOR2_X1 U931 ( .A(n1072), .B(KEYINPUT60), .Z(n1242) );
INV_X1 U932 ( .A(n1212), .ZN(n1240) );
NAND2_X1 U933 ( .A1(n1073), .A2(n1252), .ZN(n1212) );
INV_X1 U934 ( .A(n1053), .ZN(n1073) );
NAND2_X1 U935 ( .A1(n1076), .A2(n1253), .ZN(n1053) );
XNOR2_X1 U936 ( .A(G110), .B(n1206), .ZN(G12) );
NAND4_X1 U937 ( .A1(n1071), .A2(n1036), .A3(n1072), .A4(n1064), .ZN(n1206) );
NAND2_X1 U938 ( .A1(n1254), .A2(n1255), .ZN(n1064) );
OR3_X1 U939 ( .A1(n1218), .A2(n1221), .A3(KEYINPUT19), .ZN(n1255) );
INV_X1 U940 ( .A(n1245), .ZN(n1218) );
NAND2_X1 U941 ( .A1(KEYINPUT19), .A2(n1081), .ZN(n1254) );
NOR2_X1 U942 ( .A1(n1221), .A2(n1245), .ZN(n1081) );
XOR2_X1 U943 ( .A(n1087), .B(KEYINPUT23), .Z(n1245) );
XNOR2_X1 U944 ( .A(n1256), .B(G475), .ZN(n1087) );
NAND2_X1 U945 ( .A1(n1150), .A2(n1180), .ZN(n1256) );
XNOR2_X1 U946 ( .A(n1257), .B(n1258), .ZN(n1150) );
XNOR2_X1 U947 ( .A(n1259), .B(n1260), .ZN(n1258) );
NAND2_X1 U948 ( .A1(n1261), .A2(n1262), .ZN(n1259) );
NAND2_X1 U949 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
XOR2_X1 U950 ( .A(n1265), .B(KEYINPUT45), .Z(n1261) );
OR2_X1 U951 ( .A1(n1264), .A2(n1263), .ZN(n1265) );
XOR2_X1 U952 ( .A(n1266), .B(n1267), .Z(n1263) );
XNOR2_X1 U953 ( .A(n1216), .B(G131), .ZN(n1267) );
NAND2_X1 U954 ( .A1(n1268), .A2(G214), .ZN(n1266) );
XNOR2_X1 U955 ( .A(G113), .B(n1269), .ZN(n1257) );
XOR2_X1 U956 ( .A(KEYINPUT3), .B(G122), .Z(n1269) );
XNOR2_X1 U957 ( .A(n1090), .B(n1147), .ZN(n1221) );
INV_X1 U958 ( .A(G478), .ZN(n1147) );
NOR2_X1 U959 ( .A1(n1145), .A2(G902), .ZN(n1090) );
XNOR2_X1 U960 ( .A(n1270), .B(n1271), .ZN(n1145) );
XOR2_X1 U961 ( .A(G107), .B(n1272), .Z(n1271) );
XNOR2_X1 U962 ( .A(n1224), .B(G128), .ZN(n1272) );
INV_X1 U963 ( .A(G134), .ZN(n1224) );
XOR2_X1 U964 ( .A(n1273), .B(n1274), .Z(n1270) );
XOR2_X1 U965 ( .A(n1275), .B(n1276), .Z(n1274) );
AND2_X1 U966 ( .A1(n1277), .A2(G217), .ZN(n1276) );
NOR2_X1 U967 ( .A1(KEYINPUT48), .A2(n1278), .ZN(n1275) );
XNOR2_X1 U968 ( .A(n1243), .B(n1279), .ZN(n1278) );
NOR2_X1 U969 ( .A1(G122), .A2(KEYINPUT20), .ZN(n1279) );
NAND2_X1 U970 ( .A1(KEYINPUT57), .A2(n1216), .ZN(n1273) );
INV_X1 U971 ( .A(G143), .ZN(n1216) );
XOR2_X1 U972 ( .A(n1093), .B(KEYINPUT18), .Z(n1072) );
XOR2_X1 U973 ( .A(n1280), .B(G472), .Z(n1093) );
NAND2_X1 U974 ( .A1(n1281), .A2(n1180), .ZN(n1280) );
XNOR2_X1 U975 ( .A(n1158), .B(n1282), .ZN(n1281) );
NOR2_X1 U976 ( .A1(KEYINPUT40), .A2(n1283), .ZN(n1282) );
XOR2_X1 U977 ( .A(n1284), .B(n1155), .Z(n1283) );
NAND2_X1 U978 ( .A1(KEYINPUT47), .A2(n1156), .ZN(n1284) );
XNOR2_X1 U979 ( .A(n1285), .B(n1286), .ZN(n1158) );
XOR2_X1 U980 ( .A(n1287), .B(n1288), .Z(n1286) );
NAND2_X1 U981 ( .A1(n1268), .A2(G210), .ZN(n1288) );
NOR2_X1 U982 ( .A1(G953), .A2(G237), .ZN(n1268) );
NAND3_X1 U983 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1287) );
NAND2_X1 U984 ( .A1(n1292), .A2(n1243), .ZN(n1291) );
NAND2_X1 U985 ( .A1(KEYINPUT27), .A2(n1293), .ZN(n1290) );
NAND2_X1 U986 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
XNOR2_X1 U987 ( .A(KEYINPUT63), .B(n1243), .ZN(n1294) );
NAND2_X1 U988 ( .A1(n1296), .A2(n1297), .ZN(n1289) );
INV_X1 U989 ( .A(KEYINPUT27), .ZN(n1297) );
NAND2_X1 U990 ( .A1(n1298), .A2(n1299), .ZN(n1296) );
NAND2_X1 U991 ( .A1(KEYINPUT63), .A2(n1243), .ZN(n1299) );
OR3_X1 U992 ( .A1(n1292), .A2(KEYINPUT63), .A3(n1243), .ZN(n1298) );
XNOR2_X1 U993 ( .A(G101), .B(n1300), .ZN(n1285) );
NOR2_X1 U994 ( .A1(G113), .A2(KEYINPUT15), .ZN(n1300) );
INV_X1 U995 ( .A(n1213), .ZN(n1036) );
NAND2_X1 U996 ( .A1(n1220), .A2(n1252), .ZN(n1213) );
AND2_X1 U997 ( .A1(n1191), .A2(n1301), .ZN(n1252) );
NAND2_X1 U998 ( .A1(n1302), .A2(n1042), .ZN(n1301) );
NAND3_X1 U999 ( .A1(n1238), .A2(n1099), .A3(G952), .ZN(n1042) );
NAND4_X1 U1000 ( .A1(G902), .A2(n1303), .A3(n1238), .A4(n1127), .ZN(n1302) );
INV_X1 U1001 ( .A(G898), .ZN(n1127) );
NAND2_X1 U1002 ( .A1(G237), .A2(G234), .ZN(n1238) );
XNOR2_X1 U1003 ( .A(KEYINPUT8), .B(n1099), .ZN(n1303) );
NOR2_X1 U1004 ( .A1(n1077), .A2(n1079), .ZN(n1191) );
INV_X1 U1005 ( .A(n1226), .ZN(n1079) );
NAND2_X1 U1006 ( .A1(G214), .A2(n1304), .ZN(n1226) );
XOR2_X1 U1007 ( .A(n1305), .B(n1306), .Z(n1077) );
AND2_X1 U1008 ( .A1(n1304), .A2(G210), .ZN(n1306) );
NAND2_X1 U1009 ( .A1(n1307), .A2(n1180), .ZN(n1304) );
XNOR2_X1 U1010 ( .A(G237), .B(KEYINPUT29), .ZN(n1307) );
NAND2_X1 U1011 ( .A1(n1308), .A2(n1180), .ZN(n1305) );
XNOR2_X1 U1012 ( .A(n1309), .B(n1179), .ZN(n1308) );
XOR2_X1 U1013 ( .A(n1156), .B(n1310), .Z(n1179) );
XOR2_X1 U1014 ( .A(G125), .B(n1311), .Z(n1310) );
NOR2_X1 U1015 ( .A1(G953), .A2(n1119), .ZN(n1311) );
INV_X1 U1016 ( .A(G224), .ZN(n1119) );
XOR2_X1 U1017 ( .A(n1312), .B(n1313), .Z(n1156) );
INV_X1 U1018 ( .A(n1314), .ZN(n1313) );
NAND2_X1 U1019 ( .A1(KEYINPUT58), .A2(n1315), .ZN(n1312) );
INV_X1 U1020 ( .A(n1175), .ZN(n1309) );
XNOR2_X1 U1021 ( .A(n1316), .B(n1131), .ZN(n1175) );
XNOR2_X1 U1022 ( .A(n1317), .B(G122), .ZN(n1131) );
INV_X1 U1023 ( .A(G110), .ZN(n1317) );
NAND2_X1 U1024 ( .A1(KEYINPUT44), .A2(n1318), .ZN(n1316) );
XNOR2_X1 U1025 ( .A(n1129), .B(n1132), .ZN(n1318) );
INV_X1 U1026 ( .A(n1170), .ZN(n1132) );
XNOR2_X1 U1027 ( .A(n1250), .B(n1319), .ZN(n1129) );
NOR2_X1 U1028 ( .A1(KEYINPUT32), .A2(n1320), .ZN(n1319) );
XNOR2_X1 U1029 ( .A(n1243), .B(n1295), .ZN(n1320) );
INV_X1 U1030 ( .A(G116), .ZN(n1243) );
INV_X1 U1031 ( .A(G113), .ZN(n1250) );
NOR2_X1 U1032 ( .A1(n1076), .A2(n1075), .ZN(n1220) );
INV_X1 U1033 ( .A(n1253), .ZN(n1075) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1321), .ZN(n1253) );
XNOR2_X1 U1035 ( .A(n1091), .B(n1322), .ZN(n1076) );
NOR2_X1 U1036 ( .A1(G469), .A2(KEYINPUT38), .ZN(n1322) );
NAND2_X1 U1037 ( .A1(n1323), .A2(n1180), .ZN(n1091) );
XOR2_X1 U1038 ( .A(n1324), .B(n1325), .Z(n1323) );
XOR2_X1 U1039 ( .A(n1173), .B(n1326), .Z(n1325) );
NOR2_X1 U1040 ( .A1(KEYINPUT46), .A2(n1166), .ZN(n1326) );
XNOR2_X1 U1041 ( .A(n1327), .B(n1328), .ZN(n1166) );
XNOR2_X1 U1042 ( .A(G110), .B(KEYINPUT16), .ZN(n1327) );
AND2_X1 U1043 ( .A1(G227), .A2(n1099), .ZN(n1173) );
XNOR2_X1 U1044 ( .A(n1169), .B(n1170), .ZN(n1324) );
XNOR2_X1 U1045 ( .A(n1329), .B(n1260), .ZN(n1170) );
XOR2_X1 U1046 ( .A(G104), .B(KEYINPUT11), .Z(n1260) );
XNOR2_X1 U1047 ( .A(G101), .B(G107), .ZN(n1329) );
XNOR2_X1 U1048 ( .A(n1113), .B(n1155), .ZN(n1169) );
XOR2_X1 U1049 ( .A(G131), .B(n1330), .Z(n1155) );
NOR2_X1 U1050 ( .A1(KEYINPUT50), .A2(n1331), .ZN(n1330) );
XNOR2_X1 U1051 ( .A(G134), .B(G137), .ZN(n1331) );
XNOR2_X1 U1052 ( .A(n1314), .B(G128), .ZN(n1113) );
XOR2_X1 U1053 ( .A(G143), .B(n1332), .Z(n1314) );
INV_X1 U1054 ( .A(n1241), .ZN(n1071) );
XOR2_X1 U1055 ( .A(n1094), .B(n1333), .Z(n1241) );
NOR2_X1 U1056 ( .A1(n1095), .A2(KEYINPUT61), .ZN(n1333) );
INV_X1 U1057 ( .A(n1141), .ZN(n1095) );
NAND2_X1 U1058 ( .A1(G217), .A2(n1321), .ZN(n1141) );
NAND2_X1 U1059 ( .A1(G234), .A2(n1180), .ZN(n1321) );
INV_X1 U1060 ( .A(G902), .ZN(n1180) );
NOR2_X1 U1061 ( .A1(n1137), .A2(G902), .ZN(n1094) );
XOR2_X1 U1062 ( .A(n1334), .B(n1264), .Z(n1137) );
XOR2_X1 U1063 ( .A(n1114), .B(n1332), .Z(n1264) );
XOR2_X1 U1064 ( .A(G146), .B(KEYINPUT9), .Z(n1332) );
XOR2_X1 U1065 ( .A(G125), .B(n1328), .Z(n1114) );
XOR2_X1 U1066 ( .A(G140), .B(KEYINPUT24), .Z(n1328) );
XOR2_X1 U1067 ( .A(n1335), .B(n1336), .Z(n1334) );
XOR2_X1 U1068 ( .A(n1337), .B(n1338), .Z(n1336) );
XOR2_X1 U1069 ( .A(KEYINPUT22), .B(G137), .Z(n1338) );
XOR2_X1 U1070 ( .A(KEYINPUT59), .B(KEYINPUT53), .Z(n1337) );
XOR2_X1 U1071 ( .A(n1339), .B(n1340), .Z(n1335) );
XNOR2_X1 U1072 ( .A(n1315), .B(G110), .ZN(n1340) );
INV_X1 U1073 ( .A(G128), .ZN(n1315) );
XNOR2_X1 U1074 ( .A(n1341), .B(n1292), .ZN(n1339) );
INV_X1 U1075 ( .A(n1295), .ZN(n1292) );
XOR2_X1 U1076 ( .A(G119), .B(KEYINPUT5), .Z(n1295) );
NAND2_X1 U1077 ( .A1(n1277), .A2(G221), .ZN(n1341) );
AND2_X1 U1078 ( .A1(G234), .A2(n1099), .ZN(n1277) );
INV_X1 U1079 ( .A(G953), .ZN(n1099) );
endmodule


