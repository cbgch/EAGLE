//Key = 0000101111001000000101100010000010010100101110100001100111111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359;

XNOR2_X1 U749 ( .A(n1045), .B(n1046), .ZN(G9) );
NOR2_X1 U750 ( .A1(G107), .A2(KEYINPUT62), .ZN(n1046) );
NOR2_X1 U751 ( .A1(n1047), .A2(n1048), .ZN(G75) );
NOR4_X1 U752 ( .A1(n1049), .A2(n1050), .A3(G953), .A4(n1051), .ZN(n1048) );
NOR2_X1 U753 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U754 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U755 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U756 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U757 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U759 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
AND2_X1 U760 ( .A1(n1066), .A2(n1067), .ZN(n1062) );
NOR3_X1 U761 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1058) );
XNOR2_X1 U762 ( .A(n1071), .B(KEYINPUT50), .ZN(n1069) );
NOR4_X1 U763 ( .A1(n1065), .A2(n1061), .A3(n1072), .A4(n1068), .ZN(n1054) );
NAND3_X1 U764 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1049) );
XOR2_X1 U765 ( .A(n1076), .B(KEYINPUT37), .Z(n1075) );
NAND2_X1 U766 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND3_X1 U767 ( .A1(n1071), .A2(n1079), .A3(n1080), .ZN(n1078) );
NAND2_X1 U768 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
OR4_X1 U769 ( .A1(n1068), .A2(n1083), .A3(n1084), .A4(n1057), .ZN(n1082) );
INV_X1 U770 ( .A(n1085), .ZN(n1057) );
NAND2_X1 U771 ( .A1(n1086), .A2(n1087), .ZN(n1081) );
NAND2_X1 U772 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U773 ( .A1(n1090), .A2(n1091), .A3(n1085), .ZN(n1089) );
NAND2_X1 U774 ( .A1(KEYINPUT20), .A2(n1068), .ZN(n1091) );
INV_X1 U775 ( .A(n1067), .ZN(n1068) );
NAND2_X1 U776 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
INV_X1 U777 ( .A(KEYINPUT20), .ZN(n1093) );
OR2_X1 U778 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NAND2_X1 U779 ( .A1(n1067), .A2(n1096), .ZN(n1088) );
NAND4_X1 U780 ( .A1(n1080), .A2(n1067), .A3(n1097), .A4(n1086), .ZN(n1077) );
AND2_X1 U781 ( .A1(n1085), .A2(n1098), .ZN(n1097) );
INV_X1 U782 ( .A(n1053), .ZN(n1080) );
NOR3_X1 U783 ( .A1(n1051), .A2(G953), .A3(G952), .ZN(n1047) );
AND4_X1 U784 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1051) );
NOR4_X1 U785 ( .A1(n1103), .A2(n1104), .A3(n1065), .A4(n1105), .ZN(n1102) );
XOR2_X1 U786 ( .A(KEYINPUT23), .B(n1106), .Z(n1105) );
INV_X1 U787 ( .A(n1071), .ZN(n1065) );
XOR2_X1 U788 ( .A(n1107), .B(KEYINPUT57), .Z(n1103) );
AND2_X1 U789 ( .A1(n1094), .A2(n1108), .ZN(n1101) );
XNOR2_X1 U790 ( .A(n1109), .B(n1110), .ZN(n1100) );
XNOR2_X1 U791 ( .A(G469), .B(KEYINPUT58), .ZN(n1110) );
XNOR2_X1 U792 ( .A(KEYINPUT51), .B(n1084), .ZN(n1099) );
NAND3_X1 U793 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(G72) );
XOR2_X1 U794 ( .A(n1114), .B(KEYINPUT14), .Z(n1113) );
NAND3_X1 U795 ( .A1(n1115), .A2(n1116), .A3(G953), .ZN(n1114) );
NAND2_X1 U796 ( .A1(G900), .A2(G227), .ZN(n1115) );
NAND2_X1 U797 ( .A1(n1117), .A2(n1118), .ZN(n1112) );
XNOR2_X1 U798 ( .A(n1119), .B(n1120), .ZN(n1117) );
NAND2_X1 U799 ( .A1(KEYINPUT35), .A2(n1121), .ZN(n1120) );
NAND4_X1 U800 ( .A1(G900), .A2(G227), .A3(n1119), .A4(G953), .ZN(n1111) );
INV_X1 U801 ( .A(n1116), .ZN(n1119) );
NAND2_X1 U802 ( .A1(n1122), .A2(n1123), .ZN(n1116) );
NAND2_X1 U803 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XNOR2_X1 U804 ( .A(KEYINPUT47), .B(n1118), .ZN(n1124) );
XOR2_X1 U805 ( .A(n1126), .B(n1127), .Z(n1122) );
XNOR2_X1 U806 ( .A(n1128), .B(n1129), .ZN(n1127) );
XNOR2_X1 U807 ( .A(n1130), .B(n1131), .ZN(n1129) );
NOR2_X1 U808 ( .A1(G137), .A2(KEYINPUT53), .ZN(n1130) );
XNOR2_X1 U809 ( .A(G131), .B(n1132), .ZN(n1126) );
XNOR2_X1 U810 ( .A(KEYINPUT5), .B(n1133), .ZN(n1132) );
INV_X1 U811 ( .A(G134), .ZN(n1133) );
XOR2_X1 U812 ( .A(n1134), .B(n1135), .Z(G69) );
NOR2_X1 U813 ( .A1(n1136), .A2(n1118), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(n1134) );
NAND2_X1 U816 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NAND2_X1 U817 ( .A1(n1143), .A2(n1144), .ZN(n1139) );
XNOR2_X1 U818 ( .A(n1141), .B(KEYINPUT27), .ZN(n1144) );
NOR2_X1 U819 ( .A1(G953), .A2(n1073), .ZN(n1141) );
INV_X1 U820 ( .A(n1142), .ZN(n1143) );
NAND2_X1 U821 ( .A1(n1145), .A2(n1146), .ZN(n1142) );
NAND2_X1 U822 ( .A1(n1147), .A2(n1138), .ZN(n1146) );
XNOR2_X1 U823 ( .A(G953), .B(KEYINPUT12), .ZN(n1147) );
XOR2_X1 U824 ( .A(n1148), .B(n1149), .Z(n1145) );
NOR2_X1 U825 ( .A1(n1150), .A2(n1151), .ZN(G66) );
XNOR2_X1 U826 ( .A(n1152), .B(n1153), .ZN(n1151) );
NOR2_X1 U827 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NOR2_X1 U828 ( .A1(n1150), .A2(n1156), .ZN(G63) );
XOR2_X1 U829 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U830 ( .A(KEYINPUT28), .B(n1159), .Z(n1158) );
AND2_X1 U831 ( .A1(G478), .A2(n1160), .ZN(n1159) );
NOR2_X1 U832 ( .A1(n1150), .A2(n1161), .ZN(G60) );
XOR2_X1 U833 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U834 ( .A1(KEYINPUT18), .A2(n1164), .ZN(n1163) );
AND2_X1 U835 ( .A1(G475), .A2(n1160), .ZN(n1162) );
NAND3_X1 U836 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(G6) );
NAND2_X1 U837 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U838 ( .A1(n1170), .A2(n1171), .ZN(n1168) );
INV_X1 U839 ( .A(KEYINPUT31), .ZN(n1171) );
XNOR2_X1 U840 ( .A(G104), .B(KEYINPUT13), .ZN(n1170) );
OR3_X1 U841 ( .A1(n1169), .A2(G104), .A3(KEYINPUT31), .ZN(n1166) );
NAND2_X1 U842 ( .A1(G104), .A2(KEYINPUT31), .ZN(n1165) );
NOR2_X1 U843 ( .A1(n1150), .A2(n1172), .ZN(G57) );
XOR2_X1 U844 ( .A(n1173), .B(n1174), .Z(n1172) );
AND2_X1 U845 ( .A1(G472), .A2(n1160), .ZN(n1174) );
XOR2_X1 U846 ( .A(n1175), .B(n1176), .Z(n1173) );
NOR2_X1 U847 ( .A1(KEYINPUT30), .A2(n1177), .ZN(n1176) );
NAND3_X1 U848 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1175) );
NAND2_X1 U849 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
OR3_X1 U850 ( .A1(n1182), .A2(n1181), .A3(KEYINPUT33), .ZN(n1179) );
OR2_X1 U851 ( .A1(KEYINPUT16), .A2(n1183), .ZN(n1182) );
NAND2_X1 U852 ( .A1(KEYINPUT33), .A2(n1183), .ZN(n1178) );
NOR2_X1 U853 ( .A1(n1150), .A2(n1184), .ZN(G54) );
XOR2_X1 U854 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U855 ( .A1(n1187), .A2(n1155), .ZN(n1186) );
NOR2_X1 U856 ( .A1(n1188), .A2(n1189), .ZN(n1185) );
XOR2_X1 U857 ( .A(n1190), .B(KEYINPUT59), .Z(n1189) );
NAND2_X1 U858 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NOR2_X1 U859 ( .A1(n1191), .A2(n1192), .ZN(n1188) );
XOR2_X1 U860 ( .A(n1193), .B(n1194), .Z(n1192) );
XNOR2_X1 U861 ( .A(n1195), .B(n1196), .ZN(n1194) );
NOR2_X1 U862 ( .A1(KEYINPUT3), .A2(n1131), .ZN(n1196) );
XNOR2_X1 U863 ( .A(KEYINPUT52), .B(n1197), .ZN(n1191) );
NAND2_X1 U864 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NAND2_X1 U865 ( .A1(G110), .A2(n1200), .ZN(n1199) );
NAND2_X1 U866 ( .A1(n1201), .A2(n1202), .ZN(n1198) );
XNOR2_X1 U867 ( .A(KEYINPUT48), .B(n1200), .ZN(n1201) );
NOR2_X1 U868 ( .A1(n1150), .A2(n1203), .ZN(G51) );
XNOR2_X1 U869 ( .A(n1204), .B(n1205), .ZN(n1203) );
XNOR2_X1 U870 ( .A(n1206), .B(KEYINPUT25), .ZN(n1205) );
NAND3_X1 U871 ( .A1(n1160), .A2(G210), .A3(KEYINPUT7), .ZN(n1206) );
INV_X1 U872 ( .A(n1155), .ZN(n1160) );
NAND2_X1 U873 ( .A1(G902), .A2(n1207), .ZN(n1155) );
NAND2_X1 U874 ( .A1(n1073), .A2(n1074), .ZN(n1207) );
INV_X1 U875 ( .A(n1121), .ZN(n1074) );
NAND4_X1 U876 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1121) );
NOR4_X1 U877 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1211) );
INV_X1 U878 ( .A(n1216), .ZN(n1214) );
INV_X1 U879 ( .A(n1217), .ZN(n1212) );
NAND2_X1 U880 ( .A1(n1218), .A2(n1219), .ZN(n1210) );
NAND2_X1 U881 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NAND2_X1 U882 ( .A1(n1067), .A2(n1071), .ZN(n1221) );
NAND2_X1 U883 ( .A1(n1098), .A2(n1222), .ZN(n1220) );
AND4_X1 U884 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1073) );
NOR4_X1 U885 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1045), .ZN(n1226) );
AND3_X1 U886 ( .A1(n1098), .A2(n1085), .A3(n1230), .ZN(n1045) );
NOR3_X1 U887 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1225) );
NOR4_X1 U888 ( .A1(KEYINPUT32), .A2(n1234), .A3(n1061), .A4(n1072), .ZN(n1233) );
NAND3_X1 U889 ( .A1(n1064), .A2(n1235), .A3(n1098), .ZN(n1234) );
NOR2_X1 U890 ( .A1(n1236), .A2(n1237), .ZN(n1232) );
INV_X1 U891 ( .A(KEYINPUT32), .ZN(n1236) );
INV_X1 U892 ( .A(n1169), .ZN(n1231) );
NAND3_X1 U893 ( .A1(n1230), .A2(n1085), .A3(n1066), .ZN(n1169) );
NOR2_X1 U894 ( .A1(n1118), .A2(G952), .ZN(n1150) );
XNOR2_X1 U895 ( .A(G146), .B(n1208), .ZN(G48) );
NAND3_X1 U896 ( .A1(n1066), .A2(n1222), .A3(n1218), .ZN(n1208) );
XNOR2_X1 U897 ( .A(G143), .B(n1209), .ZN(G45) );
NAND3_X1 U898 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1209) );
NOR3_X1 U899 ( .A1(n1064), .A2(n1241), .A3(n1242), .ZN(n1240) );
XOR2_X1 U900 ( .A(G140), .B(n1215), .Z(G42) );
AND2_X1 U901 ( .A1(n1243), .A2(n1096), .ZN(n1215) );
XNOR2_X1 U902 ( .A(G137), .B(n1244), .ZN(G39) );
NAND3_X1 U903 ( .A1(n1218), .A2(n1071), .A3(n1245), .ZN(n1244) );
XNOR2_X1 U904 ( .A(n1067), .B(KEYINPUT22), .ZN(n1245) );
XNOR2_X1 U905 ( .A(G134), .B(n1216), .ZN(G36) );
NAND4_X1 U906 ( .A1(n1067), .A2(n1238), .A3(n1239), .A4(n1098), .ZN(n1216) );
XOR2_X1 U907 ( .A(G131), .B(n1213), .Z(G33) );
AND2_X1 U908 ( .A1(n1243), .A2(n1239), .ZN(n1213) );
AND3_X1 U909 ( .A1(n1238), .A2(n1066), .A3(n1067), .ZN(n1243) );
NOR2_X1 U910 ( .A1(n1095), .A2(n1246), .ZN(n1067) );
INV_X1 U911 ( .A(n1094), .ZN(n1246) );
XNOR2_X1 U912 ( .A(G128), .B(n1247), .ZN(G30) );
NAND3_X1 U913 ( .A1(n1218), .A2(n1098), .A3(n1248), .ZN(n1247) );
XNOR2_X1 U914 ( .A(n1222), .B(KEYINPUT61), .ZN(n1248) );
INV_X1 U915 ( .A(n1064), .ZN(n1222) );
AND3_X1 U916 ( .A1(n1104), .A2(n1106), .A3(n1238), .ZN(n1218) );
NOR2_X1 U917 ( .A1(n1070), .A2(n1249), .ZN(n1238) );
XNOR2_X1 U918 ( .A(G101), .B(n1250), .ZN(G3) );
NAND2_X1 U919 ( .A1(KEYINPUT40), .A2(n1229), .ZN(n1250) );
AND3_X1 U920 ( .A1(n1071), .A2(n1230), .A3(n1239), .ZN(n1229) );
XNOR2_X1 U921 ( .A(G125), .B(n1217), .ZN(G27) );
NAND4_X1 U922 ( .A1(n1096), .A2(n1066), .A3(n1251), .A4(n1086), .ZN(n1217) );
INV_X1 U923 ( .A(n1061), .ZN(n1086) );
NOR2_X1 U924 ( .A1(n1249), .A2(n1064), .ZN(n1251) );
AND2_X1 U925 ( .A1(n1053), .A2(n1252), .ZN(n1249) );
NAND2_X1 U926 ( .A1(n1253), .A2(n1125), .ZN(n1252) );
INV_X1 U927 ( .A(G900), .ZN(n1125) );
XNOR2_X1 U928 ( .A(G122), .B(n1254), .ZN(G24) );
NAND2_X1 U929 ( .A1(KEYINPUT44), .A2(n1228), .ZN(n1254) );
AND4_X1 U930 ( .A1(n1255), .A2(n1085), .A3(n1256), .A4(n1257), .ZN(n1228) );
NOR2_X1 U931 ( .A1(n1106), .A2(n1104), .ZN(n1085) );
XNOR2_X1 U932 ( .A(n1258), .B(n1259), .ZN(G21) );
NOR2_X1 U933 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NOR2_X1 U934 ( .A1(KEYINPUT11), .A2(n1262), .ZN(n1261) );
INV_X1 U935 ( .A(n1223), .ZN(n1262) );
NOR2_X1 U936 ( .A1(KEYINPUT21), .A2(n1223), .ZN(n1260) );
NAND4_X1 U937 ( .A1(n1255), .A2(n1071), .A3(n1104), .A4(n1106), .ZN(n1223) );
XOR2_X1 U938 ( .A(n1237), .B(n1263), .Z(G18) );
NAND2_X1 U939 ( .A1(KEYINPUT60), .A2(G116), .ZN(n1263) );
NAND3_X1 U940 ( .A1(n1239), .A2(n1098), .A3(n1255), .ZN(n1237) );
NOR2_X1 U941 ( .A1(n1257), .A2(n1242), .ZN(n1098) );
INV_X1 U942 ( .A(n1256), .ZN(n1242) );
XOR2_X1 U943 ( .A(G113), .B(n1227), .Z(G15) );
AND3_X1 U944 ( .A1(n1239), .A2(n1066), .A3(n1255), .ZN(n1227) );
NOR3_X1 U945 ( .A1(n1064), .A2(n1264), .A3(n1061), .ZN(n1255) );
NAND2_X1 U946 ( .A1(n1265), .A2(n1084), .ZN(n1061) );
INV_X1 U947 ( .A(n1083), .ZN(n1265) );
NOR2_X1 U948 ( .A1(n1256), .A2(n1241), .ZN(n1066) );
INV_X1 U949 ( .A(n1257), .ZN(n1241) );
INV_X1 U950 ( .A(n1072), .ZN(n1239) );
NAND2_X1 U951 ( .A1(n1266), .A2(n1106), .ZN(n1072) );
NAND2_X1 U952 ( .A1(n1267), .A2(n1268), .ZN(G12) );
NAND2_X1 U953 ( .A1(n1269), .A2(n1202), .ZN(n1268) );
XNOR2_X1 U954 ( .A(KEYINPUT49), .B(n1224), .ZN(n1269) );
NAND2_X1 U955 ( .A1(G110), .A2(n1270), .ZN(n1267) );
XOR2_X1 U956 ( .A(n1224), .B(KEYINPUT10), .Z(n1270) );
NAND3_X1 U957 ( .A1(n1071), .A2(n1230), .A3(n1096), .ZN(n1224) );
NOR2_X1 U958 ( .A1(n1106), .A2(n1266), .ZN(n1096) );
INV_X1 U959 ( .A(n1104), .ZN(n1266) );
XNOR2_X1 U960 ( .A(n1271), .B(n1272), .ZN(n1104) );
NOR2_X1 U961 ( .A1(n1273), .A2(n1154), .ZN(n1272) );
XOR2_X1 U962 ( .A(n1274), .B(KEYINPUT9), .Z(n1273) );
NAND2_X1 U963 ( .A1(n1152), .A2(n1275), .ZN(n1271) );
XNOR2_X1 U964 ( .A(n1276), .B(n1277), .ZN(n1152) );
XOR2_X1 U965 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U966 ( .A(n1280), .B(n1281), .Z(n1279) );
NOR2_X1 U967 ( .A1(G140), .A2(KEYINPUT54), .ZN(n1281) );
NOR2_X1 U968 ( .A1(n1282), .A2(n1283), .ZN(n1280) );
XOR2_X1 U969 ( .A(n1284), .B(KEYINPUT55), .Z(n1283) );
NAND2_X1 U970 ( .A1(n1285), .A2(n1258), .ZN(n1284) );
XOR2_X1 U971 ( .A(KEYINPUT36), .B(n1286), .Z(n1285) );
NOR2_X1 U972 ( .A1(n1258), .A2(n1286), .ZN(n1282) );
XOR2_X1 U973 ( .A(G128), .B(KEYINPUT0), .Z(n1286) );
NOR2_X1 U974 ( .A1(n1287), .A2(n1288), .ZN(n1278) );
INV_X1 U975 ( .A(G221), .ZN(n1287) );
XOR2_X1 U976 ( .A(n1289), .B(n1290), .Z(n1276) );
XNOR2_X1 U977 ( .A(n1291), .B(G137), .ZN(n1290) );
XNOR2_X1 U978 ( .A(G125), .B(G110), .ZN(n1289) );
XNOR2_X1 U979 ( .A(n1292), .B(G472), .ZN(n1106) );
NAND3_X1 U980 ( .A1(n1293), .A2(n1275), .A3(n1294), .ZN(n1292) );
NAND3_X1 U981 ( .A1(KEYINPUT56), .A2(n1181), .A3(n1295), .ZN(n1294) );
XNOR2_X1 U982 ( .A(n1177), .B(n1296), .ZN(n1295) );
AND2_X1 U983 ( .A1(n1183), .A2(KEYINPUT19), .ZN(n1296) );
NAND2_X1 U984 ( .A1(n1297), .A2(n1298), .ZN(n1293) );
NAND2_X1 U985 ( .A1(KEYINPUT56), .A2(n1181), .ZN(n1298) );
XOR2_X1 U986 ( .A(n1299), .B(n1131), .Z(n1181) );
XNOR2_X1 U987 ( .A(n1177), .B(n1300), .ZN(n1297) );
NOR2_X1 U988 ( .A1(n1183), .A2(n1301), .ZN(n1300) );
INV_X1 U989 ( .A(KEYINPUT19), .ZN(n1301) );
XOR2_X1 U990 ( .A(n1302), .B(n1303), .Z(n1183) );
XNOR2_X1 U991 ( .A(n1258), .B(n1304), .ZN(n1303) );
NOR2_X1 U992 ( .A1(G116), .A2(KEYINPUT38), .ZN(n1304) );
XNOR2_X1 U993 ( .A(n1305), .B(G101), .ZN(n1177) );
NAND2_X1 U994 ( .A1(n1306), .A2(G210), .ZN(n1305) );
NOR3_X1 U995 ( .A1(n1070), .A2(n1264), .A3(n1064), .ZN(n1230) );
NAND2_X1 U996 ( .A1(n1094), .A2(n1095), .ZN(n1064) );
NAND2_X1 U997 ( .A1(n1108), .A2(n1107), .ZN(n1095) );
NAND3_X1 U998 ( .A1(n1307), .A2(n1275), .A3(n1204), .ZN(n1107) );
NAND2_X1 U999 ( .A1(G210), .A2(G237), .ZN(n1307) );
NAND3_X1 U1000 ( .A1(n1308), .A2(n1309), .A3(G210), .ZN(n1108) );
NAND2_X1 U1001 ( .A1(n1204), .A2(n1275), .ZN(n1308) );
XOR2_X1 U1002 ( .A(n1310), .B(n1311), .Z(n1204) );
XOR2_X1 U1003 ( .A(n1312), .B(n1313), .Z(n1311) );
XNOR2_X1 U1004 ( .A(n1314), .B(n1315), .ZN(n1313) );
NOR2_X1 U1005 ( .A1(KEYINPUT24), .A2(n1148), .ZN(n1315) );
XOR2_X1 U1006 ( .A(n1316), .B(n1302), .Z(n1148) );
XOR2_X1 U1007 ( .A(G113), .B(KEYINPUT42), .Z(n1302) );
NAND2_X1 U1008 ( .A1(KEYINPUT43), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1009 ( .A(n1258), .B(G116), .ZN(n1317) );
INV_X1 U1010 ( .A(G119), .ZN(n1258) );
INV_X1 U1011 ( .A(G125), .ZN(n1314) );
NOR2_X1 U1012 ( .A1(G953), .A2(n1137), .ZN(n1312) );
INV_X1 U1013 ( .A(G224), .ZN(n1137) );
XNOR2_X1 U1014 ( .A(n1149), .B(n1131), .ZN(n1310) );
XOR2_X1 U1015 ( .A(n1318), .B(n1319), .Z(n1149) );
XOR2_X1 U1016 ( .A(KEYINPUT39), .B(G122), .Z(n1319) );
XNOR2_X1 U1017 ( .A(n1195), .B(n1202), .ZN(n1318) );
INV_X1 U1018 ( .A(G110), .ZN(n1202) );
NAND2_X1 U1019 ( .A1(G214), .A2(n1309), .ZN(n1094) );
OR2_X1 U1020 ( .A1(G237), .A2(G902), .ZN(n1309) );
INV_X1 U1021 ( .A(n1235), .ZN(n1264) );
NAND2_X1 U1022 ( .A1(n1320), .A2(n1053), .ZN(n1235) );
NAND3_X1 U1023 ( .A1(n1321), .A2(n1118), .A3(G952), .ZN(n1053) );
NAND2_X1 U1024 ( .A1(n1253), .A2(n1138), .ZN(n1320) );
INV_X1 U1025 ( .A(G898), .ZN(n1138) );
AND3_X1 U1026 ( .A1(G953), .A2(n1321), .A3(n1322), .ZN(n1253) );
XNOR2_X1 U1027 ( .A(G902), .B(KEYINPUT4), .ZN(n1322) );
NAND2_X1 U1028 ( .A1(G237), .A2(G234), .ZN(n1321) );
NAND2_X1 U1029 ( .A1(n1083), .A2(n1084), .ZN(n1070) );
NAND2_X1 U1030 ( .A1(G221), .A2(n1274), .ZN(n1084) );
NAND2_X1 U1031 ( .A1(G234), .A2(n1275), .ZN(n1274) );
NAND2_X1 U1032 ( .A1(n1323), .A2(n1324), .ZN(n1083) );
NAND2_X1 U1033 ( .A1(G469), .A2(n1325), .ZN(n1324) );
XOR2_X1 U1034 ( .A(n1326), .B(KEYINPUT15), .Z(n1323) );
NAND2_X1 U1035 ( .A1(n1109), .A2(n1327), .ZN(n1326) );
XNOR2_X1 U1036 ( .A(KEYINPUT26), .B(n1187), .ZN(n1327) );
INV_X1 U1037 ( .A(G469), .ZN(n1187) );
INV_X1 U1038 ( .A(n1325), .ZN(n1109) );
NAND2_X1 U1039 ( .A1(n1328), .A2(n1275), .ZN(n1325) );
XOR2_X1 U1040 ( .A(n1329), .B(n1330), .Z(n1328) );
XNOR2_X1 U1041 ( .A(n1195), .B(n1200), .ZN(n1330) );
XNOR2_X1 U1042 ( .A(G140), .B(n1331), .ZN(n1200) );
AND2_X1 U1043 ( .A1(n1118), .A2(G227), .ZN(n1331) );
XNOR2_X1 U1044 ( .A(G101), .B(n1332), .ZN(n1195) );
XOR2_X1 U1045 ( .A(G107), .B(G104), .Z(n1332) );
XNOR2_X1 U1046 ( .A(n1333), .B(n1131), .ZN(n1329) );
XOR2_X1 U1047 ( .A(n1334), .B(n1335), .Z(n1131) );
XNOR2_X1 U1048 ( .A(G146), .B(KEYINPUT63), .ZN(n1334) );
XNOR2_X1 U1049 ( .A(G110), .B(n1336), .ZN(n1333) );
NOR2_X1 U1050 ( .A1(KEYINPUT41), .A2(n1337), .ZN(n1336) );
XNOR2_X1 U1051 ( .A(n1193), .B(KEYINPUT46), .ZN(n1337) );
XNOR2_X1 U1052 ( .A(n1299), .B(KEYINPUT1), .ZN(n1193) );
XOR2_X1 U1053 ( .A(n1338), .B(n1339), .Z(n1299) );
NOR2_X1 U1054 ( .A1(KEYINPUT29), .A2(G131), .ZN(n1339) );
XNOR2_X1 U1055 ( .A(G134), .B(G137), .ZN(n1338) );
NOR2_X1 U1056 ( .A1(n1256), .A2(n1257), .ZN(n1071) );
XNOR2_X1 U1057 ( .A(n1340), .B(G475), .ZN(n1257) );
NAND2_X1 U1058 ( .A1(n1164), .A2(n1275), .ZN(n1340) );
INV_X1 U1059 ( .A(G902), .ZN(n1275) );
XNOR2_X1 U1060 ( .A(n1341), .B(n1342), .ZN(n1164) );
XOR2_X1 U1061 ( .A(G143), .B(G122), .Z(n1342) );
XOR2_X1 U1062 ( .A(n1343), .B(n1344), .Z(n1341) );
XOR2_X1 U1063 ( .A(n1345), .B(n1346), .Z(n1344) );
XNOR2_X1 U1064 ( .A(n1291), .B(G131), .ZN(n1346) );
INV_X1 U1065 ( .A(G146), .ZN(n1291) );
XOR2_X1 U1066 ( .A(KEYINPUT8), .B(KEYINPUT6), .Z(n1345) );
XOR2_X1 U1067 ( .A(n1347), .B(n1348), .Z(n1343) );
XOR2_X1 U1068 ( .A(G113), .B(G104), .Z(n1348) );
XOR2_X1 U1069 ( .A(n1349), .B(n1128), .Z(n1347) );
XOR2_X1 U1070 ( .A(G125), .B(G140), .Z(n1128) );
NAND2_X1 U1071 ( .A1(n1306), .A2(G214), .ZN(n1349) );
NOR2_X1 U1072 ( .A1(G953), .A2(G237), .ZN(n1306) );
XNOR2_X1 U1073 ( .A(n1350), .B(G478), .ZN(n1256) );
OR2_X1 U1074 ( .A1(n1157), .A2(G902), .ZN(n1350) );
XNOR2_X1 U1075 ( .A(n1351), .B(n1352), .ZN(n1157) );
XOR2_X1 U1076 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1077 ( .A(G107), .B(n1355), .Z(n1354) );
NOR2_X1 U1078 ( .A1(KEYINPUT45), .A2(n1356), .ZN(n1355) );
XOR2_X1 U1079 ( .A(n1357), .B(n1358), .Z(n1356) );
XOR2_X1 U1080 ( .A(KEYINPUT17), .B(G122), .Z(n1358) );
NOR2_X1 U1081 ( .A1(G116), .A2(KEYINPUT2), .ZN(n1357) );
NOR2_X1 U1082 ( .A1(G134), .A2(KEYINPUT34), .ZN(n1353) );
XOR2_X1 U1083 ( .A(n1359), .B(n1335), .Z(n1351) );
XOR2_X1 U1084 ( .A(G128), .B(G143), .Z(n1335) );
OR2_X1 U1085 ( .A1(n1154), .A2(n1288), .ZN(n1359) );
NAND2_X1 U1086 ( .A1(G234), .A2(n1118), .ZN(n1288) );
INV_X1 U1087 ( .A(G953), .ZN(n1118) );
INV_X1 U1088 ( .A(G217), .ZN(n1154) );
endmodule


