//Key = 0000101000000100111111000100110011110000001110100110111100001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351;

XOR2_X1 U739 ( .A(G107), .B(n1025), .Z(G9) );
NOR2_X1 U740 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR4_X1 U741 ( .A1(n1028), .A2(n1029), .A3(G953), .A4(n1030), .ZN(n1027) );
NOR2_X1 U742 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U743 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR3_X1 U744 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NOR2_X1 U745 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U747 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U748 ( .A1(n1044), .A2(n1045), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U750 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR3_X1 U751 ( .A1(n1041), .A2(n1050), .A3(n1045), .ZN(n1033) );
INV_X1 U752 ( .A(n1051), .ZN(n1045) );
NOR2_X1 U753 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U754 ( .A1(n1054), .A2(n1035), .ZN(n1053) );
INV_X1 U755 ( .A(n1055), .ZN(n1035) );
NOR2_X1 U756 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U757 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
XNOR2_X1 U758 ( .A(KEYINPUT9), .B(n1060), .ZN(n1059) );
NOR2_X1 U759 ( .A1(n1061), .A2(n1037), .ZN(n1052) );
INV_X1 U760 ( .A(n1062), .ZN(n1037) );
NOR2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U762 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
INV_X1 U763 ( .A(n1067), .ZN(n1041) );
INV_X1 U764 ( .A(n1068), .ZN(n1031) );
NAND3_X1 U765 ( .A1(n1069), .A2(G952), .A3(n1070), .ZN(n1028) );
XOR2_X1 U766 ( .A(n1071), .B(KEYINPUT34), .Z(n1070) );
NOR3_X1 U767 ( .A1(n1072), .A2(G953), .A3(n1030), .ZN(n1026) );
AND4_X1 U768 ( .A1(n1060), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1030) );
NOR4_X1 U769 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1066), .ZN(n1075) );
XNOR2_X1 U770 ( .A(n1079), .B(n1080), .ZN(n1078) );
XNOR2_X1 U771 ( .A(KEYINPUT42), .B(n1081), .ZN(n1079) );
NOR2_X1 U772 ( .A1(KEYINPUT7), .A2(n1082), .ZN(n1081) );
NOR2_X1 U773 ( .A1(n1049), .A2(n1083), .ZN(n1074) );
XNOR2_X1 U774 ( .A(n1084), .B(n1085), .ZN(n1083) );
XNOR2_X1 U775 ( .A(G478), .B(KEYINPUT8), .ZN(n1085) );
XNOR2_X1 U776 ( .A(G952), .B(KEYINPUT32), .ZN(n1072) );
XOR2_X1 U777 ( .A(n1086), .B(n1087), .Z(G72) );
NOR2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
AND2_X1 U779 ( .A1(G227), .A2(G900), .ZN(n1088) );
NOR2_X1 U780 ( .A1(KEYINPUT47), .A2(n1090), .ZN(n1086) );
NOR2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR3_X1 U782 ( .A1(G953), .A2(n1093), .A3(n1094), .ZN(n1092) );
NOR2_X1 U783 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
INV_X1 U784 ( .A(n1097), .ZN(n1096) );
AND2_X1 U785 ( .A1(n1095), .A2(n1069), .ZN(n1093) );
INV_X1 U786 ( .A(n1098), .ZN(n1069) );
NOR3_X1 U787 ( .A1(n1099), .A2(n1095), .A3(n1097), .ZN(n1091) );
XNOR2_X1 U788 ( .A(n1100), .B(KEYINPUT37), .ZN(n1097) );
NAND2_X1 U789 ( .A1(n1089), .A2(n1098), .ZN(n1100) );
NAND2_X1 U790 ( .A1(n1101), .A2(n1102), .ZN(n1095) );
NAND3_X1 U791 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
XOR2_X1 U792 ( .A(n1106), .B(n1107), .Z(n1105) );
NAND2_X1 U793 ( .A1(n1108), .A2(n1109), .ZN(n1101) );
NAND2_X1 U794 ( .A1(n1103), .A2(n1104), .ZN(n1109) );
NAND2_X1 U795 ( .A1(G125), .A2(n1110), .ZN(n1104) );
XNOR2_X1 U796 ( .A(KEYINPUT45), .B(n1111), .ZN(n1110) );
XNOR2_X1 U797 ( .A(KEYINPUT28), .B(n1112), .ZN(n1103) );
NAND2_X1 U798 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XNOR2_X1 U799 ( .A(KEYINPUT45), .B(n1115), .ZN(n1113) );
XNOR2_X1 U800 ( .A(n1107), .B(n1106), .ZN(n1108) );
XOR2_X1 U801 ( .A(n1116), .B(n1117), .Z(n1106) );
NOR2_X1 U802 ( .A1(G131), .A2(KEYINPUT12), .ZN(n1117) );
XOR2_X1 U803 ( .A(n1118), .B(n1119), .Z(G69) );
NOR4_X1 U804 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1119) );
INV_X1 U805 ( .A(n1124), .ZN(n1123) );
NOR2_X1 U806 ( .A1(n1125), .A2(n1126), .ZN(n1121) );
XOR2_X1 U807 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U808 ( .A(n1129), .B(G113), .Z(n1127) );
NOR3_X1 U809 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1120) );
NAND2_X1 U810 ( .A1(n1133), .A2(n1134), .ZN(n1118) );
NAND2_X1 U811 ( .A1(n1135), .A2(n1089), .ZN(n1134) );
NAND2_X1 U812 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XOR2_X1 U813 ( .A(n1138), .B(KEYINPUT0), .Z(n1136) );
NAND2_X1 U814 ( .A1(n1139), .A2(G953), .ZN(n1133) );
XOR2_X1 U815 ( .A(n1140), .B(KEYINPUT3), .Z(n1139) );
NAND2_X1 U816 ( .A1(G898), .A2(G224), .ZN(n1140) );
NOR3_X1 U817 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(G66) );
NOR2_X1 U818 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NOR2_X1 U819 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
AND2_X1 U820 ( .A1(n1148), .A2(KEYINPUT10), .ZN(n1147) );
NOR3_X1 U821 ( .A1(KEYINPUT10), .A2(n1148), .A3(n1149), .ZN(n1146) );
NOR2_X1 U822 ( .A1(n1150), .A2(n1151), .ZN(n1142) );
NOR2_X1 U823 ( .A1(n1148), .A2(n1149), .ZN(n1150) );
INV_X1 U824 ( .A(KEYINPUT54), .ZN(n1149) );
NAND3_X1 U825 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1148) );
XOR2_X1 U826 ( .A(KEYINPUT26), .B(G217), .Z(n1152) );
NOR2_X1 U827 ( .A1(n1141), .A2(n1155), .ZN(G63) );
NOR3_X1 U828 ( .A1(n1084), .A2(n1156), .A3(n1157), .ZN(n1155) );
AND3_X1 U829 ( .A1(n1158), .A2(G478), .A3(n1154), .ZN(n1157) );
NOR2_X1 U830 ( .A1(n1159), .A2(n1158), .ZN(n1156) );
NOR2_X1 U831 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR2_X1 U832 ( .A1(n1071), .A2(n1098), .ZN(n1160) );
NOR2_X1 U833 ( .A1(n1141), .A2(n1162), .ZN(G60) );
XOR2_X1 U834 ( .A(n1163), .B(n1164), .Z(n1162) );
AND2_X1 U835 ( .A1(G475), .A2(n1154), .ZN(n1163) );
XOR2_X1 U836 ( .A(n1165), .B(n1166), .Z(G6) );
NOR2_X1 U837 ( .A1(KEYINPUT39), .A2(n1167), .ZN(n1166) );
XOR2_X1 U838 ( .A(KEYINPUT33), .B(G104), .Z(n1167) );
NOR2_X1 U839 ( .A1(n1168), .A2(n1169), .ZN(n1165) );
XOR2_X1 U840 ( .A(n1170), .B(KEYINPUT30), .Z(n1168) );
NOR2_X1 U841 ( .A1(n1141), .A2(n1171), .ZN(G57) );
XOR2_X1 U842 ( .A(n1172), .B(n1173), .Z(n1171) );
AND2_X1 U843 ( .A1(G472), .A2(n1154), .ZN(n1172) );
NOR2_X1 U844 ( .A1(n1141), .A2(n1174), .ZN(G54) );
XOR2_X1 U845 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U846 ( .A(n1177), .B(n1178), .ZN(n1176) );
XNOR2_X1 U847 ( .A(n1179), .B(n1180), .ZN(n1178) );
NOR2_X1 U848 ( .A1(KEYINPUT63), .A2(n1181), .ZN(n1180) );
XOR2_X1 U849 ( .A(n1182), .B(n1183), .Z(n1175) );
XOR2_X1 U850 ( .A(KEYINPUT57), .B(n1184), .Z(n1183) );
NOR2_X1 U851 ( .A1(KEYINPUT36), .A2(n1185), .ZN(n1184) );
XOR2_X1 U852 ( .A(n1116), .B(n1186), .Z(n1185) );
NOR2_X1 U853 ( .A1(KEYINPUT31), .A2(n1187), .ZN(n1186) );
NAND2_X1 U854 ( .A1(n1154), .A2(G469), .ZN(n1182) );
NOR2_X1 U855 ( .A1(n1141), .A2(n1188), .ZN(G51) );
XOR2_X1 U856 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U857 ( .A(n1191), .B(n1192), .Z(n1190) );
NAND2_X1 U858 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NAND2_X1 U859 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XOR2_X1 U860 ( .A(n1197), .B(KEYINPUT38), .Z(n1193) );
OR2_X1 U861 ( .A1(n1196), .A2(n1195), .ZN(n1197) );
NAND2_X1 U862 ( .A1(n1154), .A2(n1198), .ZN(n1189) );
AND2_X1 U863 ( .A1(G902), .A2(n1199), .ZN(n1154) );
OR2_X1 U864 ( .A1(n1098), .A2(n1071), .ZN(n1199) );
NAND2_X1 U865 ( .A1(n1137), .A2(n1138), .ZN(n1071) );
AND4_X1 U866 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1137) );
NOR3_X1 U867 ( .A1(n1025), .A2(n1204), .A3(n1205), .ZN(n1203) );
AND2_X1 U868 ( .A1(n1206), .A2(n1207), .ZN(n1025) );
NAND2_X1 U869 ( .A1(n1047), .A2(n1208), .ZN(n1202) );
NAND2_X1 U870 ( .A1(n1209), .A2(n1170), .ZN(n1208) );
NAND3_X1 U871 ( .A1(n1210), .A2(n1064), .A3(n1207), .ZN(n1170) );
NAND4_X1 U872 ( .A1(n1211), .A2(n1051), .A3(n1066), .A4(n1212), .ZN(n1200) );
NAND4_X1 U873 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1098) );
NOR4_X1 U874 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1216) );
NOR2_X1 U875 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NOR2_X1 U876 ( .A1(n1042), .A2(n1223), .ZN(n1221) );
XNOR2_X1 U877 ( .A(n1043), .B(KEYINPUT53), .ZN(n1223) );
AND3_X1 U878 ( .A1(n1224), .A2(n1225), .A3(n1206), .ZN(n1219) );
NOR3_X1 U879 ( .A1(n1047), .A2(KEYINPUT43), .A3(n1226), .ZN(n1218) );
NOR2_X1 U880 ( .A1(n1227), .A2(n1169), .ZN(n1217) );
NOR2_X1 U881 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
INV_X1 U882 ( .A(n1230), .ZN(n1229) );
NOR2_X1 U883 ( .A1(n1226), .A2(n1231), .ZN(n1228) );
INV_X1 U884 ( .A(KEYINPUT43), .ZN(n1231) );
NOR2_X1 U885 ( .A1(n1089), .A2(G952), .ZN(n1141) );
XNOR2_X1 U886 ( .A(G146), .B(n1232), .ZN(G48) );
NAND2_X1 U887 ( .A1(n1233), .A2(n1047), .ZN(n1232) );
XOR2_X1 U888 ( .A(n1226), .B(KEYINPUT18), .Z(n1233) );
NAND3_X1 U889 ( .A1(n1234), .A2(n1064), .A3(n1224), .ZN(n1226) );
XNOR2_X1 U890 ( .A(G143), .B(n1215), .ZN(G45) );
NAND3_X1 U891 ( .A1(n1047), .A2(n1066), .A3(n1235), .ZN(n1215) );
XOR2_X1 U892 ( .A(G140), .B(n1236), .Z(G42) );
NOR2_X1 U893 ( .A1(n1237), .A2(n1222), .ZN(n1236) );
INV_X1 U894 ( .A(n1043), .ZN(n1237) );
XNOR2_X1 U895 ( .A(G137), .B(n1213), .ZN(G39) );
NAND4_X1 U896 ( .A1(n1055), .A2(n1224), .A3(n1067), .A4(n1234), .ZN(n1213) );
XNOR2_X1 U897 ( .A(G134), .B(n1214), .ZN(G36) );
NAND3_X1 U898 ( .A1(n1238), .A2(n1235), .A3(n1067), .ZN(n1214) );
AND3_X1 U899 ( .A1(n1042), .A2(n1212), .A3(n1234), .ZN(n1235) );
XOR2_X1 U900 ( .A(n1239), .B(n1240), .Z(G33) );
XNOR2_X1 U901 ( .A(KEYINPUT24), .B(n1241), .ZN(n1240) );
NOR2_X1 U902 ( .A1(n1242), .A2(n1222), .ZN(n1239) );
NAND3_X1 U903 ( .A1(n1234), .A2(n1064), .A3(n1067), .ZN(n1222) );
NOR2_X1 U904 ( .A1(n1243), .A2(n1049), .ZN(n1067) );
XNOR2_X1 U905 ( .A(n1048), .B(KEYINPUT22), .ZN(n1243) );
AND2_X1 U906 ( .A1(n1057), .A2(n1225), .ZN(n1234) );
XNOR2_X1 U907 ( .A(n1210), .B(KEYINPUT16), .ZN(n1057) );
INV_X1 U908 ( .A(n1042), .ZN(n1242) );
XNOR2_X1 U909 ( .A(G128), .B(n1244), .ZN(G30) );
NAND4_X1 U910 ( .A1(KEYINPUT49), .A2(n1206), .A3(n1245), .A4(n1225), .ZN(n1244) );
XOR2_X1 U911 ( .A(KEYINPUT27), .B(n1224), .Z(n1245) );
NOR4_X1 U912 ( .A1(n1246), .A2(n1169), .A3(n1066), .A4(n1065), .ZN(n1206) );
INV_X1 U913 ( .A(n1210), .ZN(n1246) );
XNOR2_X1 U914 ( .A(G101), .B(n1201), .ZN(G3) );
NAND3_X1 U915 ( .A1(n1042), .A2(n1047), .A3(n1247), .ZN(n1201) );
XOR2_X1 U916 ( .A(n1248), .B(n1249), .Z(G27) );
NOR2_X1 U917 ( .A1(n1250), .A2(n1230), .ZN(n1249) );
NAND4_X1 U918 ( .A1(n1043), .A2(n1062), .A3(n1064), .A4(n1225), .ZN(n1230) );
NAND2_X1 U919 ( .A1(n1251), .A2(n1252), .ZN(n1225) );
NAND4_X1 U920 ( .A1(G953), .A2(G902), .A3(n1068), .A4(n1099), .ZN(n1252) );
INV_X1 U921 ( .A(G900), .ZN(n1099) );
XNOR2_X1 U922 ( .A(n1047), .B(KEYINPUT11), .ZN(n1250) );
NAND2_X1 U923 ( .A1(KEYINPUT60), .A2(n1114), .ZN(n1248) );
XNOR2_X1 U924 ( .A(G122), .B(n1253), .ZN(G24) );
NAND4_X1 U925 ( .A1(n1207), .A2(n1254), .A3(n1255), .A4(n1062), .ZN(n1253) );
XOR2_X1 U926 ( .A(KEYINPUT1), .B(n1256), .Z(n1255) );
NOR2_X1 U927 ( .A1(n1065), .A2(n1238), .ZN(n1256) );
INV_X1 U928 ( .A(n1212), .ZN(n1065) );
XNOR2_X1 U929 ( .A(KEYINPUT40), .B(n1169), .ZN(n1254) );
AND2_X1 U930 ( .A1(n1051), .A2(n1257), .ZN(n1207) );
NOR2_X1 U931 ( .A1(n1258), .A2(n1259), .ZN(n1051) );
XOR2_X1 U932 ( .A(G119), .B(n1205), .Z(G21) );
AND3_X1 U933 ( .A1(n1055), .A2(n1224), .A3(n1211), .ZN(n1205) );
NOR2_X1 U934 ( .A1(n1260), .A2(n1073), .ZN(n1224) );
XOR2_X1 U935 ( .A(G116), .B(n1261), .Z(G18) );
NOR2_X1 U936 ( .A1(KEYINPUT59), .A2(n1138), .ZN(n1261) );
NAND4_X1 U937 ( .A1(n1211), .A2(n1042), .A3(n1238), .A4(n1212), .ZN(n1138) );
XOR2_X1 U938 ( .A(G113), .B(n1204), .Z(G15) );
AND3_X1 U939 ( .A1(n1042), .A2(n1064), .A3(n1211), .ZN(n1204) );
AND3_X1 U940 ( .A1(n1062), .A2(n1257), .A3(n1047), .ZN(n1211) );
INV_X1 U941 ( .A(n1169), .ZN(n1047) );
NAND2_X1 U942 ( .A1(n1262), .A2(n1263), .ZN(n1062) );
OR3_X1 U943 ( .A1(n1264), .A2(n1077), .A3(KEYINPUT9), .ZN(n1263) );
NAND2_X1 U944 ( .A1(KEYINPUT9), .A2(n1210), .ZN(n1262) );
NAND2_X1 U945 ( .A1(n1265), .A2(n1266), .ZN(n1064) );
OR3_X1 U946 ( .A1(n1238), .A2(n1212), .A3(KEYINPUT41), .ZN(n1266) );
INV_X1 U947 ( .A(n1066), .ZN(n1238) );
NAND2_X1 U948 ( .A1(KEYINPUT41), .A2(n1055), .ZN(n1265) );
NOR2_X1 U949 ( .A1(n1073), .A2(n1259), .ZN(n1042) );
INV_X1 U950 ( .A(n1260), .ZN(n1259) );
INV_X1 U951 ( .A(n1258), .ZN(n1073) );
XNOR2_X1 U952 ( .A(n1267), .B(n1268), .ZN(G12) );
NOR2_X1 U953 ( .A1(n1169), .A2(n1269), .ZN(n1268) );
XNOR2_X1 U954 ( .A(KEYINPUT17), .B(n1209), .ZN(n1269) );
NAND2_X1 U955 ( .A1(n1247), .A2(n1043), .ZN(n1209) );
NOR2_X1 U956 ( .A1(n1260), .A2(n1258), .ZN(n1043) );
XNOR2_X1 U957 ( .A(n1270), .B(G472), .ZN(n1258) );
OR2_X1 U958 ( .A1(n1173), .A2(G902), .ZN(n1270) );
XNOR2_X1 U959 ( .A(n1271), .B(n1272), .ZN(n1173) );
XOR2_X1 U960 ( .A(n1273), .B(n1274), .Z(n1272) );
XOR2_X1 U961 ( .A(n1275), .B(n1276), .Z(n1274) );
NOR2_X1 U962 ( .A1(G113), .A2(KEYINPUT23), .ZN(n1276) );
AND3_X1 U963 ( .A1(G210), .A2(n1089), .A3(n1277), .ZN(n1275) );
XNOR2_X1 U964 ( .A(n1129), .B(n1278), .ZN(n1271) );
XNOR2_X1 U965 ( .A(G101), .B(n1279), .ZN(n1129) );
XOR2_X1 U966 ( .A(n1280), .B(n1082), .Z(n1260) );
NAND2_X1 U967 ( .A1(n1281), .A2(n1282), .ZN(n1082) );
XNOR2_X1 U968 ( .A(KEYINPUT13), .B(n1151), .ZN(n1281) );
INV_X1 U969 ( .A(n1144), .ZN(n1151) );
XNOR2_X1 U970 ( .A(n1283), .B(n1284), .ZN(n1144) );
XOR2_X1 U971 ( .A(n1179), .B(n1285), .Z(n1284) );
XOR2_X1 U972 ( .A(n1286), .B(n1287), .Z(n1285) );
NOR2_X1 U973 ( .A1(G137), .A2(KEYINPUT58), .ZN(n1286) );
XOR2_X1 U974 ( .A(n1288), .B(n1289), .Z(n1283) );
XOR2_X1 U975 ( .A(KEYINPUT20), .B(G128), .Z(n1289) );
XOR2_X1 U976 ( .A(n1290), .B(G119), .Z(n1288) );
NAND3_X1 U977 ( .A1(G221), .A2(n1089), .A3(n1291), .ZN(n1290) );
NAND2_X1 U978 ( .A1(KEYINPUT55), .A2(n1080), .ZN(n1280) );
NAND2_X1 U979 ( .A1(G217), .A2(n1153), .ZN(n1080) );
AND3_X1 U980 ( .A1(n1210), .A2(n1257), .A3(n1055), .ZN(n1247) );
NOR2_X1 U981 ( .A1(n1212), .A2(n1066), .ZN(n1055) );
XNOR2_X1 U982 ( .A(n1292), .B(G475), .ZN(n1066) );
OR2_X1 U983 ( .A1(n1164), .A2(G902), .ZN(n1292) );
XNOR2_X1 U984 ( .A(n1293), .B(n1294), .ZN(n1164) );
XOR2_X1 U985 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U986 ( .A(n1297), .B(G104), .Z(n1296) );
NAND2_X1 U987 ( .A1(n1298), .A2(KEYINPUT46), .ZN(n1297) );
XNOR2_X1 U988 ( .A(G122), .B(n1299), .ZN(n1298) );
NOR2_X1 U989 ( .A1(G113), .A2(KEYINPUT2), .ZN(n1299) );
XNOR2_X1 U990 ( .A(G143), .B(G131), .ZN(n1295) );
XOR2_X1 U991 ( .A(n1300), .B(n1287), .Z(n1293) );
XNOR2_X1 U992 ( .A(n1114), .B(G146), .ZN(n1287) );
INV_X1 U993 ( .A(G125), .ZN(n1114) );
XOR2_X1 U994 ( .A(n1301), .B(n1302), .Z(n1300) );
NOR2_X1 U995 ( .A1(KEYINPUT56), .A2(n1111), .ZN(n1302) );
INV_X1 U996 ( .A(n1115), .ZN(n1111) );
NAND3_X1 U997 ( .A1(n1277), .A2(n1089), .A3(G214), .ZN(n1301) );
INV_X1 U998 ( .A(G237), .ZN(n1277) );
XOR2_X1 U999 ( .A(n1303), .B(n1161), .Z(n1212) );
INV_X1 U1000 ( .A(G478), .ZN(n1161) );
NAND2_X1 U1001 ( .A1(KEYINPUT29), .A2(n1084), .ZN(n1303) );
NOR2_X1 U1002 ( .A1(n1158), .A2(G902), .ZN(n1084) );
XOR2_X1 U1003 ( .A(n1304), .B(n1305), .Z(n1158) );
XOR2_X1 U1004 ( .A(G116), .B(n1306), .Z(n1305) );
XOR2_X1 U1005 ( .A(G134), .B(G122), .Z(n1306) );
XOR2_X1 U1006 ( .A(n1307), .B(n1308), .Z(n1304) );
XOR2_X1 U1007 ( .A(n1309), .B(G107), .Z(n1307) );
NAND3_X1 U1008 ( .A1(n1291), .A2(n1089), .A3(G217), .ZN(n1309) );
XNOR2_X1 U1009 ( .A(G234), .B(KEYINPUT19), .ZN(n1291) );
NAND2_X1 U1010 ( .A1(n1251), .A2(n1310), .ZN(n1257) );
NAND3_X1 U1011 ( .A1(G902), .A2(n1068), .A3(n1122), .ZN(n1310) );
AND2_X1 U1012 ( .A1(n1311), .A2(G953), .ZN(n1122) );
XNOR2_X1 U1013 ( .A(G898), .B(KEYINPUT5), .ZN(n1311) );
NAND3_X1 U1014 ( .A1(G952), .A2(n1068), .A3(n1312), .ZN(n1251) );
XNOR2_X1 U1015 ( .A(G953), .B(KEYINPUT14), .ZN(n1312) );
NAND2_X1 U1016 ( .A1(G237), .A2(G234), .ZN(n1068) );
NOR2_X1 U1017 ( .A1(n1060), .A2(n1077), .ZN(n1210) );
INV_X1 U1018 ( .A(n1058), .ZN(n1077) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1153), .ZN(n1058) );
NAND2_X1 U1020 ( .A1(G234), .A2(n1313), .ZN(n1153) );
INV_X1 U1021 ( .A(n1264), .ZN(n1060) );
XOR2_X1 U1022 ( .A(G469), .B(n1314), .Z(n1264) );
NOR2_X1 U1023 ( .A1(G902), .A2(n1315), .ZN(n1314) );
NOR2_X1 U1024 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XOR2_X1 U1025 ( .A(n1318), .B(KEYINPUT52), .Z(n1317) );
NAND2_X1 U1026 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
OR2_X1 U1027 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NOR3_X1 U1028 ( .A1(n1321), .A2(n1322), .A3(n1319), .ZN(n1316) );
XOR2_X1 U1029 ( .A(n1181), .B(n1179), .Z(n1319) );
XOR2_X1 U1030 ( .A(G110), .B(n1115), .Z(n1179) );
XOR2_X1 U1031 ( .A(G140), .B(KEYINPUT35), .Z(n1115) );
NAND2_X1 U1032 ( .A1(G227), .A2(n1089), .ZN(n1181) );
AND2_X1 U1033 ( .A1(n1278), .A2(n1323), .ZN(n1322) );
INV_X1 U1034 ( .A(n1177), .ZN(n1278) );
XNOR2_X1 U1035 ( .A(n1324), .B(KEYINPUT15), .ZN(n1321) );
NAND2_X1 U1036 ( .A1(n1325), .A2(n1177), .ZN(n1324) );
XOR2_X1 U1037 ( .A(n1107), .B(n1326), .Z(n1177) );
NOR2_X1 U1038 ( .A1(KEYINPUT51), .A2(n1241), .ZN(n1326) );
INV_X1 U1039 ( .A(G131), .ZN(n1241) );
XOR2_X1 U1040 ( .A(G134), .B(G137), .Z(n1107) );
XOR2_X1 U1041 ( .A(n1323), .B(KEYINPUT25), .Z(n1325) );
XOR2_X1 U1042 ( .A(n1116), .B(n1187), .Z(n1323) );
XNOR2_X1 U1043 ( .A(n1327), .B(G101), .ZN(n1187) );
NAND2_X1 U1044 ( .A1(KEYINPUT4), .A2(n1128), .ZN(n1327) );
NAND2_X1 U1045 ( .A1(n1328), .A2(n1329), .ZN(n1116) );
NAND2_X1 U1046 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
XOR2_X1 U1047 ( .A(KEYINPUT44), .B(n1308), .Z(n1330) );
NAND2_X1 U1048 ( .A1(n1308), .A2(G146), .ZN(n1328) );
NAND2_X1 U1049 ( .A1(n1332), .A2(n1049), .ZN(n1169) );
XNOR2_X1 U1050 ( .A(n1333), .B(n1198), .ZN(n1049) );
AND2_X1 U1051 ( .A1(G210), .A2(n1334), .ZN(n1198) );
NAND2_X1 U1052 ( .A1(n1335), .A2(n1282), .ZN(n1333) );
XOR2_X1 U1053 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1054 ( .A(n1191), .B(n1196), .Z(n1337) );
NAND2_X1 U1055 ( .A1(G224), .A2(n1089), .ZN(n1196) );
INV_X1 U1056 ( .A(G953), .ZN(n1089) );
NAND3_X1 U1057 ( .A1(n1338), .A2(n1339), .A3(n1124), .ZN(n1191) );
NAND3_X1 U1058 ( .A1(n1132), .A2(n1125), .A3(n1131), .ZN(n1124) );
NAND2_X1 U1059 ( .A1(n1340), .A2(n1132), .ZN(n1339) );
INV_X1 U1060 ( .A(n1341), .ZN(n1132) );
NAND2_X1 U1061 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
NAND2_X1 U1062 ( .A1(n1125), .A2(n1344), .ZN(n1343) );
NAND2_X1 U1063 ( .A1(n1345), .A2(n1130), .ZN(n1342) );
INV_X1 U1064 ( .A(n1125), .ZN(n1130) );
NAND2_X1 U1065 ( .A1(n1346), .A2(n1341), .ZN(n1338) );
XOR2_X1 U1066 ( .A(G113), .B(n1279), .Z(n1341) );
XOR2_X1 U1067 ( .A(G116), .B(G119), .Z(n1279) );
XNOR2_X1 U1068 ( .A(n1125), .B(n1345), .ZN(n1346) );
NOR2_X1 U1069 ( .A1(n1344), .A2(n1131), .ZN(n1345) );
XNOR2_X1 U1070 ( .A(G101), .B(n1128), .ZN(n1131) );
XOR2_X1 U1071 ( .A(G104), .B(G107), .Z(n1128) );
INV_X1 U1072 ( .A(KEYINPUT6), .ZN(n1344) );
NAND2_X1 U1073 ( .A1(n1347), .A2(n1348), .ZN(n1125) );
NAND2_X1 U1074 ( .A1(G122), .A2(n1267), .ZN(n1348) );
XOR2_X1 U1075 ( .A(KEYINPUT21), .B(n1349), .Z(n1347) );
NOR2_X1 U1076 ( .A1(G122), .A2(n1267), .ZN(n1349) );
NOR2_X1 U1077 ( .A1(KEYINPUT48), .A2(n1195), .ZN(n1336) );
XOR2_X1 U1078 ( .A(G125), .B(n1273), .Z(n1195) );
XNOR2_X1 U1079 ( .A(n1331), .B(n1308), .ZN(n1273) );
XOR2_X1 U1080 ( .A(G128), .B(G143), .Z(n1308) );
INV_X1 U1081 ( .A(G146), .ZN(n1331) );
XNOR2_X1 U1082 ( .A(n1076), .B(KEYINPUT22), .ZN(n1332) );
INV_X1 U1083 ( .A(n1048), .ZN(n1076) );
NAND2_X1 U1084 ( .A1(G214), .A2(n1334), .ZN(n1048) );
NAND2_X1 U1085 ( .A1(n1350), .A2(n1351), .ZN(n1334) );
XOR2_X1 U1086 ( .A(KEYINPUT61), .B(n1313), .Z(n1351) );
XNOR2_X1 U1087 ( .A(n1282), .B(KEYINPUT50), .ZN(n1313) );
INV_X1 U1088 ( .A(G902), .ZN(n1282) );
XNOR2_X1 U1089 ( .A(G237), .B(KEYINPUT62), .ZN(n1350) );
INV_X1 U1090 ( .A(G110), .ZN(n1267) );
endmodule


