//Key = 1011011111000000111101010000111111001011000101100110110100000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327;

XNOR2_X1 U726 ( .A(G107), .B(n998), .ZN(G9) );
NOR2_X1 U727 ( .A1(n999), .A2(n1000), .ZN(G75) );
NOR4_X1 U728 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n1000) );
NOR2_X1 U729 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NOR2_X1 U730 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
XOR2_X1 U731 ( .A(KEYINPUT1), .B(n1009), .Z(n1008) );
NOR2_X1 U732 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NOR3_X1 U733 ( .A1(n1012), .A2(n1013), .A3(n1011), .ZN(n1007) );
NOR2_X1 U734 ( .A1(n1014), .A2(n1015), .ZN(n1003) );
NOR2_X1 U735 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR2_X1 U736 ( .A1(n1018), .A2(n1011), .ZN(n1017) );
INV_X1 U737 ( .A(n1019), .ZN(n1011) );
NOR2_X1 U738 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR2_X1 U739 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR4_X1 U740 ( .A1(n1024), .A2(n1025), .A3(n1006), .A4(n1026), .ZN(n1016) );
NOR3_X1 U741 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1025) );
NOR2_X1 U742 ( .A1(n1030), .A2(n1031), .ZN(n1024) );
NOR2_X1 U743 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U744 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
INV_X1 U745 ( .A(n1036), .ZN(n1002) );
NAND3_X1 U746 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1001) );
NAND2_X1 U747 ( .A1(n1040), .A2(n1012), .ZN(n1039) );
INV_X1 U748 ( .A(KEYINPUT49), .ZN(n1012) );
NAND2_X1 U749 ( .A1(n1019), .A2(n1041), .ZN(n1040) );
NOR3_X1 U750 ( .A1(n1027), .A2(n1033), .A3(n1026), .ZN(n1019) );
INV_X1 U751 ( .A(n1042), .ZN(n1033) );
NOR3_X1 U752 ( .A1(n1043), .A2(G953), .A3(G952), .ZN(n999) );
INV_X1 U753 ( .A(n1037), .ZN(n1043) );
NAND4_X1 U754 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1037) );
NOR4_X1 U755 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
XNOR2_X1 U756 ( .A(n1052), .B(n1053), .ZN(n1050) );
XNOR2_X1 U757 ( .A(G478), .B(KEYINPUT43), .ZN(n1052) );
NOR2_X1 U758 ( .A1(n1015), .A2(n1054), .ZN(n1046) );
XNOR2_X1 U759 ( .A(G469), .B(n1055), .ZN(n1054) );
NAND2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(n1045) );
INV_X1 U761 ( .A(KEYINPUT9), .ZN(n1057) );
NAND2_X1 U762 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NAND2_X1 U763 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(n1058) );
NAND2_X1 U765 ( .A1(KEYINPUT9), .A2(n1064), .ZN(n1044) );
NAND2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U767 ( .A1(n1062), .A2(n1061), .ZN(n1066) );
XNOR2_X1 U768 ( .A(n1067), .B(KEYINPUT22), .ZN(n1062) );
NAND2_X1 U769 ( .A1(n1063), .A2(n1060), .ZN(n1065) );
XNOR2_X1 U770 ( .A(n1067), .B(KEYINPUT30), .ZN(n1060) );
XOR2_X1 U771 ( .A(n1068), .B(KEYINPUT13), .Z(n1067) );
XOR2_X1 U772 ( .A(n1069), .B(n1070), .Z(G72) );
XOR2_X1 U773 ( .A(n1071), .B(n1072), .Z(n1070) );
NOR2_X1 U774 ( .A1(n1073), .A2(G953), .ZN(n1072) );
NOR2_X1 U775 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U776 ( .A1(n1076), .A2(n1077), .ZN(n1071) );
XOR2_X1 U777 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U778 ( .A1(G900), .A2(n1038), .ZN(n1076) );
NOR2_X1 U779 ( .A1(n1080), .A2(n1038), .ZN(n1069) );
AND2_X1 U780 ( .A1(G227), .A2(G900), .ZN(n1080) );
XOR2_X1 U781 ( .A(n1081), .B(n1082), .Z(G69) );
XOR2_X1 U782 ( .A(n1083), .B(n1084), .Z(n1082) );
NAND2_X1 U783 ( .A1(G953), .A2(n1085), .ZN(n1084) );
NAND2_X1 U784 ( .A1(G898), .A2(G224), .ZN(n1085) );
NAND4_X1 U785 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1083) );
NAND2_X1 U786 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
INV_X1 U787 ( .A(KEYINPUT39), .ZN(n1091) );
NAND2_X1 U788 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
XNOR2_X1 U789 ( .A(n1094), .B(KEYINPUT27), .ZN(n1092) );
NAND2_X1 U790 ( .A1(KEYINPUT39), .A2(n1095), .ZN(n1088) );
NAND2_X1 U791 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
OR3_X1 U792 ( .A1(n1094), .A2(n1098), .A3(KEYINPUT27), .ZN(n1097) );
NAND2_X1 U793 ( .A1(KEYINPUT27), .A2(n1094), .ZN(n1096) );
NAND2_X1 U794 ( .A1(n1094), .A2(n1098), .ZN(n1087) );
NAND2_X1 U795 ( .A1(G953), .A2(n1099), .ZN(n1086) );
NOR2_X1 U796 ( .A1(n1100), .A2(G953), .ZN(n1081) );
NOR3_X1 U797 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1100) );
XOR2_X1 U798 ( .A(KEYINPUT34), .B(n1104), .Z(n1103) );
NAND3_X1 U799 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1101) );
NOR2_X1 U800 ( .A1(n1108), .A2(n1109), .ZN(G66) );
XOR2_X1 U801 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U802 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U803 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
XNOR2_X1 U804 ( .A(KEYINPUT5), .B(KEYINPUT45), .ZN(n1110) );
NOR2_X1 U805 ( .A1(G952), .A2(n1116), .ZN(n1108) );
XNOR2_X1 U806 ( .A(KEYINPUT52), .B(n1038), .ZN(n1116) );
NOR2_X1 U807 ( .A1(n1117), .A2(n1118), .ZN(G63) );
NOR3_X1 U808 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1118) );
AND3_X1 U809 ( .A1(n1122), .A2(G478), .A3(n1123), .ZN(n1121) );
NOR2_X1 U810 ( .A1(n1124), .A2(n1122), .ZN(n1120) );
NOR2_X1 U811 ( .A1(n1036), .A2(n1125), .ZN(n1124) );
NOR2_X1 U812 ( .A1(n1117), .A2(n1126), .ZN(G60) );
XOR2_X1 U813 ( .A(n1127), .B(n1128), .Z(n1126) );
AND2_X1 U814 ( .A1(G475), .A2(n1123), .ZN(n1127) );
XNOR2_X1 U815 ( .A(G104), .B(n1129), .ZN(G6) );
NOR2_X1 U816 ( .A1(n1117), .A2(n1130), .ZN(G57) );
XOR2_X1 U817 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U818 ( .A(n1133), .B(n1134), .ZN(n1132) );
NOR2_X1 U819 ( .A1(KEYINPUT47), .A2(n1135), .ZN(n1134) );
XOR2_X1 U820 ( .A(n1136), .B(n1137), .Z(n1131) );
AND2_X1 U821 ( .A1(G472), .A2(n1123), .ZN(n1137) );
NOR2_X1 U822 ( .A1(n1117), .A2(n1138), .ZN(G54) );
XOR2_X1 U823 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U824 ( .A(n1141), .B(n1142), .Z(n1140) );
XNOR2_X1 U825 ( .A(G134), .B(n1143), .ZN(n1142) );
AND2_X1 U826 ( .A1(G469), .A2(n1123), .ZN(n1141) );
XOR2_X1 U827 ( .A(n1144), .B(n1145), .Z(n1139) );
XOR2_X1 U828 ( .A(n1146), .B(n1147), .Z(n1144) );
NAND3_X1 U829 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1146) );
NAND2_X1 U830 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
OR3_X1 U831 ( .A1(n1152), .A2(n1151), .A3(n1153), .ZN(n1149) );
INV_X1 U832 ( .A(KEYINPUT31), .ZN(n1152) );
NAND2_X1 U833 ( .A1(n1153), .A2(n1154), .ZN(n1148) );
NAND2_X1 U834 ( .A1(n1155), .A2(KEYINPUT31), .ZN(n1154) );
XNOR2_X1 U835 ( .A(n1156), .B(KEYINPUT53), .ZN(n1155) );
XOR2_X1 U836 ( .A(G128), .B(n1157), .Z(n1153) );
NOR2_X1 U837 ( .A1(n1117), .A2(n1158), .ZN(G51) );
NOR2_X1 U838 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U839 ( .A(n1161), .B(KEYINPUT3), .Z(n1160) );
NAND2_X1 U840 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U841 ( .A(n1164), .B(KEYINPUT37), .Z(n1162) );
OR2_X1 U842 ( .A1(n1115), .A2(n1068), .ZN(n1164) );
NOR3_X1 U843 ( .A1(n1115), .A2(n1165), .A3(n1068), .ZN(n1159) );
XOR2_X1 U844 ( .A(n1163), .B(KEYINPUT40), .Z(n1165) );
XOR2_X1 U845 ( .A(n1166), .B(n1167), .Z(n1163) );
XOR2_X1 U846 ( .A(KEYINPUT41), .B(G125), .Z(n1167) );
XOR2_X1 U847 ( .A(n1168), .B(n1169), .Z(n1166) );
NAND2_X1 U848 ( .A1(KEYINPUT55), .A2(n1170), .ZN(n1168) );
INV_X1 U849 ( .A(n1171), .ZN(n1170) );
INV_X1 U850 ( .A(n1123), .ZN(n1115) );
NOR2_X1 U851 ( .A1(n1172), .A2(n1036), .ZN(n1123) );
NOR4_X1 U852 ( .A1(n1075), .A2(n1102), .A3(n1173), .A4(n1174), .ZN(n1036) );
XNOR2_X1 U853 ( .A(KEYINPUT10), .B(n1175), .ZN(n1174) );
NOR4_X1 U854 ( .A1(n1104), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1175) );
XOR2_X1 U855 ( .A(n1107), .B(KEYINPUT38), .Z(n1178) );
INV_X1 U856 ( .A(n1105), .ZN(n1177) );
INV_X1 U857 ( .A(n1106), .ZN(n1176) );
AND2_X1 U858 ( .A1(n1021), .A2(n1179), .ZN(n1104) );
XNOR2_X1 U859 ( .A(KEYINPUT14), .B(n1180), .ZN(n1179) );
XOR2_X1 U860 ( .A(KEYINPUT25), .B(n1074), .Z(n1173) );
NAND4_X1 U861 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1074) );
NAND4_X1 U862 ( .A1(n1129), .A2(n1185), .A3(n1186), .A4(n998), .ZN(n1102) );
NAND3_X1 U863 ( .A1(n1187), .A2(n1028), .A3(n1188), .ZN(n998) );
NAND3_X1 U864 ( .A1(n1188), .A2(n1187), .A3(n1029), .ZN(n1129) );
NAND3_X1 U865 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1075) );
NAND2_X1 U866 ( .A1(n1021), .A2(n1192), .ZN(n1191) );
NAND2_X1 U867 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NAND3_X1 U868 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1194) );
XNOR2_X1 U869 ( .A(KEYINPUT58), .B(n1013), .ZN(n1196) );
NAND2_X1 U870 ( .A1(n1029), .A2(n1198), .ZN(n1193) );
NAND2_X1 U871 ( .A1(n1199), .A2(n1200), .ZN(n1189) );
XOR2_X1 U872 ( .A(KEYINPUT61), .B(n1201), .Z(n1200) );
NOR2_X1 U873 ( .A1(n1038), .A2(G952), .ZN(n1117) );
XOR2_X1 U874 ( .A(G146), .B(n1202), .Z(G48) );
NOR3_X1 U875 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1202) );
XNOR2_X1 U876 ( .A(n1021), .B(KEYINPUT51), .ZN(n1204) );
XNOR2_X1 U877 ( .A(G143), .B(n1206), .ZN(G45) );
NAND4_X1 U878 ( .A1(n1207), .A2(KEYINPUT36), .A3(n1208), .A4(n1209), .ZN(n1206) );
NOR2_X1 U879 ( .A1(n1210), .A2(n1211), .ZN(n1208) );
XNOR2_X1 U880 ( .A(n1197), .B(KEYINPUT18), .ZN(n1207) );
XNOR2_X1 U881 ( .A(G140), .B(n1212), .ZN(G42) );
NAND3_X1 U882 ( .A1(n1201), .A2(n1199), .A3(KEYINPUT0), .ZN(n1212) );
NOR3_X1 U883 ( .A1(n1211), .A2(n1010), .A3(n1203), .ZN(n1201) );
INV_X1 U884 ( .A(n1195), .ZN(n1211) );
XNOR2_X1 U885 ( .A(G137), .B(n1190), .ZN(G39) );
NAND3_X1 U886 ( .A1(n1199), .A2(n1198), .A3(n1042), .ZN(n1190) );
XNOR2_X1 U887 ( .A(G134), .B(n1181), .ZN(G36) );
NAND3_X1 U888 ( .A1(n1195), .A2(n1028), .A3(n1041), .ZN(n1181) );
XNOR2_X1 U889 ( .A(G131), .B(n1182), .ZN(G33) );
NAND3_X1 U890 ( .A1(n1029), .A2(n1195), .A3(n1041), .ZN(n1182) );
NOR2_X1 U891 ( .A1(n1013), .A2(n1006), .ZN(n1041) );
INV_X1 U892 ( .A(n1199), .ZN(n1006) );
NOR2_X1 U893 ( .A1(n1022), .A2(n1048), .ZN(n1199) );
INV_X1 U894 ( .A(n1023), .ZN(n1048) );
INV_X1 U895 ( .A(n1209), .ZN(n1013) );
XNOR2_X1 U896 ( .A(G128), .B(n1183), .ZN(G30) );
NAND3_X1 U897 ( .A1(n1028), .A2(n1021), .A3(n1198), .ZN(n1183) );
INV_X1 U898 ( .A(n1205), .ZN(n1198) );
NAND3_X1 U899 ( .A1(n1213), .A2(n1214), .A3(n1195), .ZN(n1205) );
NOR3_X1 U900 ( .A1(n1215), .A2(n1049), .A3(n1034), .ZN(n1195) );
INV_X1 U901 ( .A(n1210), .ZN(n1021) );
XNOR2_X1 U902 ( .A(G101), .B(n1185), .ZN(G3) );
NAND3_X1 U903 ( .A1(n1042), .A2(n1188), .A3(n1209), .ZN(n1185) );
XNOR2_X1 U904 ( .A(G125), .B(n1184), .ZN(G27) );
NAND3_X1 U905 ( .A1(n1030), .A2(n1029), .A3(n1216), .ZN(n1184) );
NOR3_X1 U906 ( .A1(n1210), .A2(n1215), .A3(n1010), .ZN(n1216) );
INV_X1 U907 ( .A(n1217), .ZN(n1010) );
AND2_X1 U908 ( .A1(n1026), .A2(n1218), .ZN(n1215) );
NAND3_X1 U909 ( .A1(G953), .A2(n1219), .A3(n1220), .ZN(n1218) );
INV_X1 U910 ( .A(G900), .ZN(n1219) );
XNOR2_X1 U911 ( .A(n1221), .B(n1222), .ZN(G24) );
NOR2_X1 U912 ( .A1(n1210), .A2(n1180), .ZN(n1222) );
NAND4_X1 U913 ( .A1(n1030), .A2(n1197), .A3(n1187), .A4(n1223), .ZN(n1180) );
AND2_X1 U914 ( .A1(n1224), .A2(n1051), .ZN(n1197) );
INV_X1 U915 ( .A(n1027), .ZN(n1030) );
XNOR2_X1 U916 ( .A(G119), .B(n1105), .ZN(G21) );
NAND4_X1 U917 ( .A1(n1225), .A2(n1042), .A3(n1213), .A4(n1214), .ZN(n1105) );
XNOR2_X1 U918 ( .A(G116), .B(n1106), .ZN(G18) );
NAND3_X1 U919 ( .A1(n1209), .A2(n1028), .A3(n1225), .ZN(n1106) );
NOR2_X1 U920 ( .A1(n1051), .A2(n1226), .ZN(n1028) );
XNOR2_X1 U921 ( .A(n1107), .B(n1227), .ZN(G15) );
NOR2_X1 U922 ( .A1(KEYINPUT56), .A2(n1228), .ZN(n1227) );
NAND3_X1 U923 ( .A1(n1209), .A2(n1029), .A3(n1225), .ZN(n1107) );
NOR3_X1 U924 ( .A1(n1210), .A2(n1229), .A3(n1027), .ZN(n1225) );
NAND2_X1 U925 ( .A1(n1034), .A2(n1035), .ZN(n1027) );
INV_X1 U926 ( .A(n1203), .ZN(n1029) );
NAND2_X1 U927 ( .A1(n1226), .A2(n1051), .ZN(n1203) );
NOR2_X1 U928 ( .A1(n1214), .A2(n1230), .ZN(n1209) );
XNOR2_X1 U929 ( .A(G110), .B(n1186), .ZN(G12) );
NAND3_X1 U930 ( .A1(n1188), .A2(n1217), .A3(n1042), .ZN(n1186) );
NOR2_X1 U931 ( .A1(n1051), .A2(n1224), .ZN(n1042) );
INV_X1 U932 ( .A(n1226), .ZN(n1224) );
XOR2_X1 U933 ( .A(n1231), .B(n1125), .Z(n1226) );
INV_X1 U934 ( .A(G478), .ZN(n1125) );
NAND2_X1 U935 ( .A1(KEYINPUT29), .A2(n1053), .ZN(n1231) );
INV_X1 U936 ( .A(n1119), .ZN(n1053) );
NOR2_X1 U937 ( .A1(n1122), .A2(G902), .ZN(n1119) );
NAND2_X1 U938 ( .A1(n1232), .A2(n1233), .ZN(n1122) );
NAND2_X1 U939 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U940 ( .A1(KEYINPUT6), .A2(n1236), .ZN(n1235) );
NAND4_X1 U941 ( .A1(n1237), .A2(G217), .A3(n1238), .A4(n1239), .ZN(n1236) );
INV_X1 U942 ( .A(n1240), .ZN(n1234) );
NAND2_X1 U943 ( .A1(n1241), .A2(n1242), .ZN(n1232) );
NAND3_X1 U944 ( .A1(n1237), .A2(n1238), .A3(G217), .ZN(n1242) );
XNOR2_X1 U945 ( .A(n1038), .B(KEYINPUT23), .ZN(n1238) );
NAND2_X1 U946 ( .A1(n1243), .A2(n1239), .ZN(n1241) );
INV_X1 U947 ( .A(KEYINPUT57), .ZN(n1239) );
NAND2_X1 U948 ( .A1(KEYINPUT6), .A2(n1240), .ZN(n1243) );
XNOR2_X1 U949 ( .A(n1244), .B(n1245), .ZN(n1240) );
XOR2_X1 U950 ( .A(G107), .B(n1246), .Z(n1245) );
XNOR2_X1 U951 ( .A(KEYINPUT2), .B(n1247), .ZN(n1246) );
INV_X1 U952 ( .A(G116), .ZN(n1247) );
XOR2_X1 U953 ( .A(n1248), .B(n1249), .Z(n1244) );
XOR2_X1 U954 ( .A(n1250), .B(n1251), .Z(n1248) );
NAND2_X1 U955 ( .A1(KEYINPUT28), .A2(n1221), .ZN(n1250) );
XNOR2_X1 U956 ( .A(n1252), .B(G475), .ZN(n1051) );
OR2_X1 U957 ( .A1(n1128), .A2(G902), .ZN(n1252) );
XNOR2_X1 U958 ( .A(n1253), .B(n1254), .ZN(n1128) );
XNOR2_X1 U959 ( .A(n1255), .B(n1256), .ZN(n1254) );
NAND2_X1 U960 ( .A1(n1257), .A2(KEYINPUT21), .ZN(n1255) );
XOR2_X1 U961 ( .A(n1258), .B(n1259), .Z(n1257) );
NOR2_X1 U962 ( .A1(KEYINPUT11), .A2(n1249), .ZN(n1259) );
XNOR2_X1 U963 ( .A(n1260), .B(n1261), .ZN(n1258) );
INV_X1 U964 ( .A(G131), .ZN(n1261) );
NAND2_X1 U965 ( .A1(n1262), .A2(G214), .ZN(n1260) );
XNOR2_X1 U966 ( .A(G104), .B(n1263), .ZN(n1253) );
XNOR2_X1 U967 ( .A(n1221), .B(G113), .ZN(n1263) );
NAND2_X1 U968 ( .A1(n1264), .A2(n1265), .ZN(n1217) );
OR2_X1 U969 ( .A1(n1015), .A2(KEYINPUT32), .ZN(n1265) );
INV_X1 U970 ( .A(n1187), .ZN(n1015) );
NOR2_X1 U971 ( .A1(n1214), .A2(n1213), .ZN(n1187) );
NAND3_X1 U972 ( .A1(n1214), .A2(n1230), .A3(KEYINPUT32), .ZN(n1264) );
INV_X1 U973 ( .A(n1213), .ZN(n1230) );
XNOR2_X1 U974 ( .A(n1266), .B(G472), .ZN(n1213) );
NAND2_X1 U975 ( .A1(n1267), .A2(n1172), .ZN(n1266) );
XOR2_X1 U976 ( .A(n1268), .B(n1269), .Z(n1267) );
XNOR2_X1 U977 ( .A(n1135), .B(n1270), .ZN(n1269) );
NOR2_X1 U978 ( .A1(KEYINPUT60), .A2(n1136), .ZN(n1270) );
NAND2_X1 U979 ( .A1(n1262), .A2(G210), .ZN(n1136) );
NOR2_X1 U980 ( .A1(G953), .A2(G237), .ZN(n1262) );
INV_X1 U981 ( .A(G101), .ZN(n1135) );
NOR2_X1 U982 ( .A1(KEYINPUT44), .A2(n1133), .ZN(n1268) );
XNOR2_X1 U983 ( .A(n1271), .B(n1272), .ZN(n1133) );
XNOR2_X1 U984 ( .A(G113), .B(n1273), .ZN(n1272) );
XNOR2_X1 U985 ( .A(n1274), .B(n1275), .ZN(n1271) );
XOR2_X1 U986 ( .A(n1276), .B(n1114), .Z(n1214) );
NAND2_X1 U987 ( .A1(G217), .A2(n1277), .ZN(n1114) );
NAND2_X1 U988 ( .A1(n1278), .A2(n1172), .ZN(n1276) );
XOR2_X1 U989 ( .A(KEYINPUT12), .B(n1113), .Z(n1278) );
XNOR2_X1 U990 ( .A(n1279), .B(n1280), .ZN(n1113) );
XNOR2_X1 U991 ( .A(n1281), .B(n1282), .ZN(n1280) );
INV_X1 U992 ( .A(n1256), .ZN(n1282) );
XOR2_X1 U993 ( .A(G146), .B(n1078), .Z(n1256) );
XOR2_X1 U994 ( .A(G140), .B(G125), .Z(n1078) );
NOR2_X1 U995 ( .A1(n1283), .A2(n1284), .ZN(n1281) );
XOR2_X1 U996 ( .A(n1285), .B(KEYINPUT33), .Z(n1284) );
NAND2_X1 U997 ( .A1(G128), .A2(n1286), .ZN(n1285) );
NOR2_X1 U998 ( .A1(G128), .A2(n1286), .ZN(n1283) );
XOR2_X1 U999 ( .A(n1287), .B(G110), .Z(n1279) );
NAND3_X1 U1000 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n1287) );
NAND2_X1 U1001 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
INV_X1 U1002 ( .A(KEYINPUT19), .ZN(n1292) );
NAND3_X1 U1003 ( .A1(KEYINPUT19), .A2(n1293), .A3(n1294), .ZN(n1289) );
OR2_X1 U1004 ( .A1(n1294), .A2(n1293), .ZN(n1288) );
NOR2_X1 U1005 ( .A1(KEYINPUT4), .A2(n1291), .ZN(n1293) );
NAND3_X1 U1006 ( .A1(G221), .A2(n1038), .A3(n1237), .ZN(n1291) );
XNOR2_X1 U1007 ( .A(G234), .B(KEYINPUT8), .ZN(n1237) );
NOR4_X1 U1008 ( .A1(n1034), .A2(n1210), .A3(n1229), .A4(n1049), .ZN(n1188) );
INV_X1 U1009 ( .A(n1035), .ZN(n1049) );
NAND2_X1 U1010 ( .A1(G221), .A2(n1277), .ZN(n1035) );
NAND2_X1 U1011 ( .A1(G234), .A2(n1172), .ZN(n1277) );
INV_X1 U1012 ( .A(n1223), .ZN(n1229) );
NAND2_X1 U1013 ( .A1(n1026), .A2(n1295), .ZN(n1223) );
NAND3_X1 U1014 ( .A1(n1296), .A2(n1099), .A3(n1220), .ZN(n1295) );
AND2_X1 U1015 ( .A1(n1297), .A2(n1298), .ZN(n1220) );
XNOR2_X1 U1016 ( .A(KEYINPUT59), .B(n1172), .ZN(n1297) );
INV_X1 U1017 ( .A(G898), .ZN(n1099) );
XNOR2_X1 U1018 ( .A(KEYINPUT15), .B(n1038), .ZN(n1296) );
NAND3_X1 U1019 ( .A1(n1298), .A2(n1038), .A3(G952), .ZN(n1026) );
NAND2_X1 U1020 ( .A1(G237), .A2(G234), .ZN(n1298) );
NAND2_X1 U1021 ( .A1(n1022), .A2(n1023), .ZN(n1210) );
NAND2_X1 U1022 ( .A1(G214), .A2(n1299), .ZN(n1023) );
XOR2_X1 U1023 ( .A(n1068), .B(n1300), .Z(n1022) );
NOR2_X1 U1024 ( .A1(n1063), .A2(KEYINPUT20), .ZN(n1300) );
INV_X1 U1025 ( .A(n1061), .ZN(n1063) );
NAND2_X1 U1026 ( .A1(n1301), .A2(n1172), .ZN(n1061) );
XOR2_X1 U1027 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U1028 ( .A(n1304), .B(n1169), .Z(n1303) );
XNOR2_X1 U1029 ( .A(n1305), .B(n1306), .ZN(n1169) );
XNOR2_X1 U1030 ( .A(n1098), .B(n1307), .ZN(n1306) );
INV_X1 U1031 ( .A(n1094), .ZN(n1307) );
XNOR2_X1 U1032 ( .A(n1308), .B(n1309), .ZN(n1094) );
XOR2_X1 U1033 ( .A(n1310), .B(n1311), .Z(n1309) );
NAND2_X1 U1034 ( .A1(KEYINPUT7), .A2(n1312), .ZN(n1310) );
INV_X1 U1035 ( .A(G104), .ZN(n1312) );
XNOR2_X1 U1036 ( .A(n1313), .B(n1228), .ZN(n1308) );
INV_X1 U1037 ( .A(G113), .ZN(n1228) );
NAND2_X1 U1038 ( .A1(KEYINPUT16), .A2(n1274), .ZN(n1313) );
XNOR2_X1 U1039 ( .A(G116), .B(n1286), .ZN(n1274) );
INV_X1 U1040 ( .A(G119), .ZN(n1286) );
INV_X1 U1041 ( .A(n1093), .ZN(n1098) );
XOR2_X1 U1042 ( .A(G110), .B(n1221), .Z(n1093) );
INV_X1 U1043 ( .A(G122), .ZN(n1221) );
XOR2_X1 U1044 ( .A(n1273), .B(n1314), .Z(n1305) );
XOR2_X1 U1045 ( .A(KEYINPUT17), .B(G128), .Z(n1314) );
NAND2_X1 U1046 ( .A1(n1315), .A2(n1316), .ZN(n1273) );
OR2_X1 U1047 ( .A1(n1249), .A2(G146), .ZN(n1316) );
XOR2_X1 U1048 ( .A(n1317), .B(KEYINPUT42), .Z(n1315) );
NAND2_X1 U1049 ( .A1(G146), .A2(n1249), .ZN(n1317) );
NOR2_X1 U1050 ( .A1(G125), .A2(KEYINPUT24), .ZN(n1304) );
XOR2_X1 U1051 ( .A(n1318), .B(n1319), .Z(n1302) );
XOR2_X1 U1052 ( .A(KEYINPUT63), .B(KEYINPUT46), .Z(n1319) );
NOR2_X1 U1053 ( .A1(KEYINPUT26), .A2(n1171), .ZN(n1318) );
NAND2_X1 U1054 ( .A1(G224), .A2(n1038), .ZN(n1171) );
NAND2_X1 U1055 ( .A1(G210), .A2(n1299), .ZN(n1068) );
NAND2_X1 U1056 ( .A1(n1320), .A2(n1172), .ZN(n1299) );
INV_X1 U1057 ( .A(G237), .ZN(n1320) );
XNOR2_X1 U1058 ( .A(n1055), .B(n1321), .ZN(n1034) );
NOR2_X1 U1059 ( .A1(G469), .A2(KEYINPUT54), .ZN(n1321) );
NAND2_X1 U1060 ( .A1(n1322), .A2(n1172), .ZN(n1055) );
INV_X1 U1061 ( .A(G902), .ZN(n1172) );
XOR2_X1 U1062 ( .A(n1323), .B(n1324), .Z(n1322) );
XNOR2_X1 U1063 ( .A(n1325), .B(n1151), .ZN(n1324) );
INV_X1 U1064 ( .A(n1156), .ZN(n1151) );
XNOR2_X1 U1065 ( .A(n1311), .B(n1326), .ZN(n1156) );
NOR2_X1 U1066 ( .A1(G104), .A2(KEYINPUT48), .ZN(n1326) );
XNOR2_X1 U1067 ( .A(G107), .B(G101), .ZN(n1311) );
NOR2_X1 U1068 ( .A1(KEYINPUT35), .A2(n1143), .ZN(n1325) );
NAND2_X1 U1069 ( .A1(G227), .A2(n1038), .ZN(n1143) );
INV_X1 U1070 ( .A(G953), .ZN(n1038) );
XNOR2_X1 U1071 ( .A(n1145), .B(n1079), .ZN(n1323) );
XOR2_X1 U1072 ( .A(n1275), .B(n1157), .Z(n1079) );
XOR2_X1 U1073 ( .A(n1249), .B(n1327), .Z(n1157) );
NOR2_X1 U1074 ( .A1(G146), .A2(KEYINPUT62), .ZN(n1327) );
XOR2_X1 U1075 ( .A(G143), .B(KEYINPUT50), .Z(n1249) );
XOR2_X1 U1076 ( .A(n1147), .B(n1251), .Z(n1275) );
XOR2_X1 U1077 ( .A(G134), .B(G128), .Z(n1251) );
XNOR2_X1 U1078 ( .A(G131), .B(n1294), .ZN(n1147) );
INV_X1 U1079 ( .A(G137), .ZN(n1294) );
XOR2_X1 U1080 ( .A(G140), .B(G110), .Z(n1145) );
endmodule


