//Key = 0100100000101101010000110011100000010110101101111010101001011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338;

XOR2_X1 U731 ( .A(G107), .B(n1022), .Z(G9) );
NOR2_X1 U732 ( .A1(n1023), .A2(n1024), .ZN(G75) );
XOR2_X1 U733 ( .A(KEYINPUT56), .B(n1025), .Z(n1024) );
NOR3_X1 U734 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NAND3_X1 U735 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1026) );
NAND2_X1 U736 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NAND2_X1 U737 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND3_X1 U738 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NAND2_X1 U739 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NAND3_X1 U740 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NAND2_X1 U741 ( .A1(n1044), .A2(n1045), .ZN(n1039) );
NAND2_X1 U742 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U743 ( .A1(n1042), .A2(n1048), .ZN(n1034) );
NAND2_X1 U744 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND3_X1 U745 ( .A1(n1038), .A2(n1051), .A3(n1044), .ZN(n1050) );
OR2_X1 U746 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U747 ( .A1(n1036), .A2(n1054), .ZN(n1049) );
NAND2_X1 U748 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U749 ( .A1(n1044), .A2(n1057), .ZN(n1056) );
NAND2_X1 U750 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U751 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U752 ( .A1(n1038), .A2(n1062), .ZN(n1055) );
XNOR2_X1 U753 ( .A(KEYINPUT49), .B(n1063), .ZN(n1062) );
INV_X1 U754 ( .A(n1064), .ZN(n1032) );
INV_X1 U755 ( .A(n1065), .ZN(n1029) );
NOR2_X1 U756 ( .A1(G952), .A2(n1065), .ZN(n1023) );
NAND2_X1 U757 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND4_X1 U758 ( .A1(n1068), .A2(n1036), .A3(n1069), .A4(n1070), .ZN(n1067) );
NOR4_X1 U759 ( .A1(n1061), .A2(n1043), .A3(n1071), .A4(n1072), .ZN(n1070) );
XOR2_X1 U760 ( .A(n1073), .B(n1074), .Z(n1071) );
NOR2_X1 U761 ( .A1(n1075), .A2(KEYINPUT2), .ZN(n1074) );
INV_X1 U762 ( .A(n1076), .ZN(n1075) );
XOR2_X1 U763 ( .A(n1077), .B(n1078), .Z(n1069) );
XNOR2_X1 U764 ( .A(n1079), .B(n1080), .ZN(n1068) );
XOR2_X1 U765 ( .A(n1081), .B(n1082), .Z(G72) );
XOR2_X1 U766 ( .A(n1083), .B(n1084), .Z(n1082) );
NOR3_X1 U767 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
NOR2_X1 U768 ( .A1(KEYINPUT8), .A2(n1027), .ZN(n1087) );
NOR2_X1 U769 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
INV_X1 U770 ( .A(KEYINPUT8), .ZN(n1089) );
XNOR2_X1 U771 ( .A(G953), .B(KEYINPUT48), .ZN(n1085) );
NAND2_X1 U772 ( .A1(n1090), .A2(n1091), .ZN(n1083) );
NAND2_X1 U773 ( .A1(G953), .A2(n1092), .ZN(n1091) );
XOR2_X1 U774 ( .A(n1093), .B(n1094), .Z(n1090) );
XNOR2_X1 U775 ( .A(n1095), .B(n1096), .ZN(n1094) );
NOR2_X1 U776 ( .A1(KEYINPUT19), .A2(n1097), .ZN(n1096) );
XNOR2_X1 U777 ( .A(G134), .B(n1098), .ZN(n1093) );
NAND2_X1 U778 ( .A1(G953), .A2(n1099), .ZN(n1081) );
NAND2_X1 U779 ( .A1(G900), .A2(G227), .ZN(n1099) );
XOR2_X1 U780 ( .A(n1100), .B(n1101), .Z(G69) );
NOR2_X1 U781 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR3_X1 U782 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1103) );
NOR2_X1 U783 ( .A1(G953), .A2(n1107), .ZN(n1106) );
AND2_X1 U784 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U785 ( .A1(G224), .A2(n1066), .ZN(n1105) );
NOR2_X1 U786 ( .A1(KEYINPUT54), .A2(G953), .ZN(n1102) );
NOR2_X1 U787 ( .A1(n1104), .A2(n1110), .ZN(n1100) );
XOR2_X1 U788 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U789 ( .A1(KEYINPUT53), .A2(n1113), .ZN(n1111) );
NOR2_X1 U790 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U791 ( .A(KEYINPUT3), .B(n1116), .Z(n1115) );
NOR2_X1 U792 ( .A1(n1117), .A2(n1118), .ZN(G66) );
XOR2_X1 U793 ( .A(n1119), .B(n1120), .Z(n1118) );
NOR2_X1 U794 ( .A1(n1076), .A2(n1121), .ZN(n1120) );
NOR2_X1 U795 ( .A1(n1117), .A2(n1122), .ZN(G63) );
XOR2_X1 U796 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND3_X1 U797 ( .A1(n1125), .A2(G478), .A3(KEYINPUT59), .ZN(n1123) );
NOR2_X1 U798 ( .A1(n1117), .A2(n1126), .ZN(G60) );
XOR2_X1 U799 ( .A(n1127), .B(n1128), .Z(n1126) );
AND2_X1 U800 ( .A1(G475), .A2(n1125), .ZN(n1127) );
XOR2_X1 U801 ( .A(G104), .B(n1129), .Z(G6) );
NOR2_X1 U802 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U803 ( .A1(n1117), .A2(n1132), .ZN(G57) );
XOR2_X1 U804 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U805 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U806 ( .A1(n1080), .A2(n1121), .ZN(n1136) );
INV_X1 U807 ( .A(G472), .ZN(n1080) );
NAND2_X1 U808 ( .A1(KEYINPUT1), .A2(n1137), .ZN(n1135) );
XOR2_X1 U809 ( .A(n1138), .B(KEYINPUT41), .Z(n1137) );
XNOR2_X1 U810 ( .A(n1139), .B(n1140), .ZN(n1133) );
NOR2_X1 U811 ( .A1(n1117), .A2(n1141), .ZN(G54) );
XOR2_X1 U812 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U813 ( .A(n1144), .B(n1145), .Z(n1143) );
NAND2_X1 U814 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
INV_X1 U815 ( .A(n1148), .ZN(n1147) );
NAND2_X1 U816 ( .A1(n1149), .A2(n1150), .ZN(n1146) );
XNOR2_X1 U817 ( .A(KEYINPUT4), .B(n1151), .ZN(n1150) );
XNOR2_X1 U818 ( .A(G140), .B(KEYINPUT46), .ZN(n1149) );
NAND2_X1 U819 ( .A1(n1152), .A2(n1153), .ZN(n1144) );
NAND2_X1 U820 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XOR2_X1 U821 ( .A(KEYINPUT26), .B(n1156), .Z(n1152) );
NOR2_X1 U822 ( .A1(n1154), .A2(n1155), .ZN(n1156) );
NAND2_X1 U823 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
OR2_X1 U824 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U825 ( .A(n1161), .B(KEYINPUT55), .Z(n1157) );
NAND2_X1 U826 ( .A1(n1159), .A2(n1160), .ZN(n1161) );
INV_X1 U827 ( .A(n1162), .ZN(n1154) );
XOR2_X1 U828 ( .A(n1163), .B(n1164), .Z(n1142) );
AND2_X1 U829 ( .A1(G469), .A2(n1125), .ZN(n1163) );
INV_X1 U830 ( .A(n1121), .ZN(n1125) );
NOR2_X1 U831 ( .A1(n1117), .A2(n1165), .ZN(G51) );
XOR2_X1 U832 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U833 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U834 ( .A(n1170), .B(n1171), .Z(n1166) );
XOR2_X1 U835 ( .A(KEYINPUT25), .B(G125), .Z(n1171) );
NOR2_X1 U836 ( .A1(n1078), .A2(n1121), .ZN(n1170) );
NAND2_X1 U837 ( .A1(G902), .A2(n1172), .ZN(n1121) );
NAND3_X1 U838 ( .A1(n1031), .A2(n1109), .A3(n1173), .ZN(n1172) );
XOR2_X1 U839 ( .A(n1027), .B(KEYINPUT17), .Z(n1173) );
NAND3_X1 U840 ( .A1(n1088), .A2(n1174), .A3(n1175), .ZN(n1027) );
NOR3_X1 U841 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1175) );
AND4_X1 U842 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1088) );
NAND3_X1 U843 ( .A1(n1053), .A2(n1183), .A3(n1184), .ZN(n1179) );
INV_X1 U844 ( .A(n1028), .ZN(n1109) );
NAND4_X1 U845 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1028) );
NOR4_X1 U846 ( .A1(n1189), .A2(n1190), .A3(n1022), .A4(n1191), .ZN(n1188) );
AND3_X1 U847 ( .A1(n1053), .A2(n1042), .A3(n1192), .ZN(n1022) );
NAND2_X1 U848 ( .A1(KEYINPUT13), .A2(n1193), .ZN(n1187) );
NAND3_X1 U849 ( .A1(n1194), .A2(n1195), .A3(n1192), .ZN(n1186) );
NAND2_X1 U850 ( .A1(n1036), .A2(n1046), .ZN(n1195) );
INV_X1 U851 ( .A(n1196), .ZN(n1046) );
NAND2_X1 U852 ( .A1(n1197), .A2(n1198), .ZN(n1194) );
INV_X1 U853 ( .A(n1036), .ZN(n1198) );
OR2_X1 U854 ( .A1(n1047), .A2(KEYINPUT13), .ZN(n1197) );
NAND2_X1 U855 ( .A1(n1199), .A2(n1200), .ZN(n1185) );
XOR2_X1 U856 ( .A(n1131), .B(KEYINPUT50), .Z(n1199) );
NAND4_X1 U857 ( .A1(n1052), .A2(n1042), .A3(n1201), .A4(n1202), .ZN(n1131) );
XOR2_X1 U858 ( .A(n1108), .B(KEYINPUT20), .Z(n1031) );
NOR2_X1 U859 ( .A1(n1066), .A2(G952), .ZN(n1117) );
XOR2_X1 U860 ( .A(n1203), .B(n1176), .Z(G48) );
AND3_X1 U861 ( .A1(n1052), .A2(n1183), .A3(n1184), .ZN(n1176) );
XNOR2_X1 U862 ( .A(G146), .B(KEYINPUT57), .ZN(n1203) );
XOR2_X1 U863 ( .A(n1174), .B(n1204), .Z(G45) );
XOR2_X1 U864 ( .A(KEYINPUT42), .B(G143), .Z(n1204) );
NAND4_X1 U865 ( .A1(n1205), .A2(n1183), .A3(n1206), .A4(n1207), .ZN(n1174) );
XOR2_X1 U866 ( .A(G140), .B(n1178), .Z(G42) );
AND3_X1 U867 ( .A1(n1196), .A2(n1044), .A3(n1208), .ZN(n1178) );
NOR3_X1 U868 ( .A1(n1209), .A2(n1210), .A3(n1058), .ZN(n1208) );
XOR2_X1 U869 ( .A(G137), .B(n1177), .Z(G39) );
AND3_X1 U870 ( .A1(n1044), .A2(n1036), .A3(n1184), .ZN(n1177) );
XOR2_X1 U871 ( .A(n1180), .B(n1211), .Z(G36) );
NAND2_X1 U872 ( .A1(KEYINPUT10), .A2(G134), .ZN(n1211) );
NAND3_X1 U873 ( .A1(n1044), .A2(n1053), .A3(n1205), .ZN(n1180) );
XNOR2_X1 U874 ( .A(G131), .B(n1181), .ZN(G33) );
NAND3_X1 U875 ( .A1(n1044), .A2(n1052), .A3(n1205), .ZN(n1181) );
NOR3_X1 U876 ( .A1(n1058), .A2(n1210), .A3(n1047), .ZN(n1205) );
NOR2_X1 U877 ( .A1(n1212), .A2(n1043), .ZN(n1044) );
XNOR2_X1 U878 ( .A(G128), .B(n1213), .ZN(G30) );
NAND4_X1 U879 ( .A1(KEYINPUT38), .A2(n1184), .A3(n1053), .A4(n1183), .ZN(n1213) );
AND4_X1 U880 ( .A1(n1214), .A2(n1201), .A3(n1215), .A4(n1216), .ZN(n1184) );
XOR2_X1 U881 ( .A(n1217), .B(n1193), .Z(G3) );
AND3_X1 U882 ( .A1(n1036), .A2(n1192), .A3(n1218), .ZN(n1193) );
NAND2_X1 U883 ( .A1(KEYINPUT27), .A2(n1140), .ZN(n1217) );
XNOR2_X1 U884 ( .A(G125), .B(n1182), .ZN(G27) );
NAND3_X1 U885 ( .A1(n1196), .A2(n1052), .A3(n1219), .ZN(n1182) );
NOR3_X1 U886 ( .A1(n1220), .A2(n1210), .A3(n1063), .ZN(n1219) );
INV_X1 U887 ( .A(n1216), .ZN(n1210) );
NAND2_X1 U888 ( .A1(n1064), .A2(n1221), .ZN(n1216) );
NAND4_X1 U889 ( .A1(G902), .A2(G953), .A3(n1222), .A4(n1092), .ZN(n1221) );
INV_X1 U890 ( .A(G900), .ZN(n1092) );
INV_X1 U891 ( .A(n1209), .ZN(n1052) );
XOR2_X1 U892 ( .A(n1190), .B(n1223), .Z(G24) );
NOR2_X1 U893 ( .A1(KEYINPUT11), .A2(n1224), .ZN(n1223) );
AND4_X1 U894 ( .A1(n1225), .A2(n1042), .A3(n1206), .A4(n1207), .ZN(n1190) );
NOR2_X1 U895 ( .A1(n1215), .A2(n1226), .ZN(n1042) );
XOR2_X1 U896 ( .A(G119), .B(n1191), .Z(G21) );
AND4_X1 U897 ( .A1(n1214), .A2(n1225), .A3(n1036), .A4(n1215), .ZN(n1191) );
XNOR2_X1 U898 ( .A(n1227), .B(n1189), .ZN(G18) );
AND3_X1 U899 ( .A1(n1225), .A2(n1053), .A3(n1218), .ZN(n1189) );
INV_X1 U900 ( .A(n1047), .ZN(n1218) );
NOR2_X1 U901 ( .A1(n1207), .A2(n1228), .ZN(n1053) );
NOR3_X1 U902 ( .A1(n1063), .A2(n1229), .A3(n1220), .ZN(n1225) );
INV_X1 U903 ( .A(n1183), .ZN(n1063) );
XNOR2_X1 U904 ( .A(G113), .B(n1108), .ZN(G15) );
NAND4_X1 U905 ( .A1(n1200), .A2(n1202), .A3(n1038), .A4(n1230), .ZN(n1108) );
NOR2_X1 U906 ( .A1(n1047), .A2(n1209), .ZN(n1230) );
NAND2_X1 U907 ( .A1(n1228), .A2(n1207), .ZN(n1209) );
INV_X1 U908 ( .A(n1206), .ZN(n1228) );
NAND2_X1 U909 ( .A1(n1214), .A2(n1231), .ZN(n1047) );
XNOR2_X1 U910 ( .A(n1232), .B(KEYINPUT16), .ZN(n1214) );
INV_X1 U911 ( .A(n1220), .ZN(n1038) );
NAND2_X1 U912 ( .A1(n1233), .A2(n1060), .ZN(n1220) );
INV_X1 U913 ( .A(n1072), .ZN(n1060) );
XNOR2_X1 U914 ( .A(G110), .B(n1234), .ZN(G12) );
NAND4_X1 U915 ( .A1(n1196), .A2(n1036), .A3(n1235), .A4(n1236), .ZN(n1234) );
OR2_X1 U916 ( .A1(n1192), .A2(KEYINPUT34), .ZN(n1236) );
NOR3_X1 U917 ( .A1(n1130), .A2(n1229), .A3(n1058), .ZN(n1192) );
NAND2_X1 U918 ( .A1(KEYINPUT34), .A2(n1237), .ZN(n1235) );
NAND3_X1 U919 ( .A1(n1200), .A2(n1201), .A3(n1229), .ZN(n1237) );
INV_X1 U920 ( .A(n1202), .ZN(n1229) );
NAND2_X1 U921 ( .A1(n1064), .A2(n1238), .ZN(n1202) );
NAND3_X1 U922 ( .A1(n1104), .A2(n1222), .A3(G902), .ZN(n1238) );
NOR2_X1 U923 ( .A1(G898), .A2(n1066), .ZN(n1104) );
NAND3_X1 U924 ( .A1(n1222), .A2(n1066), .A3(G952), .ZN(n1064) );
NAND2_X1 U925 ( .A1(G237), .A2(G234), .ZN(n1222) );
INV_X1 U926 ( .A(n1058), .ZN(n1201) );
NAND2_X1 U927 ( .A1(n1233), .A2(n1072), .ZN(n1058) );
XNOR2_X1 U928 ( .A(n1239), .B(G469), .ZN(n1072) );
NAND2_X1 U929 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
XOR2_X1 U930 ( .A(n1242), .B(n1243), .Z(n1240) );
NOR2_X1 U931 ( .A1(n1244), .A2(n1148), .ZN(n1243) );
NOR2_X1 U932 ( .A1(n1151), .A2(G140), .ZN(n1148) );
NOR2_X1 U933 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
XNOR2_X1 U934 ( .A(KEYINPUT33), .B(n1151), .ZN(n1246) );
XOR2_X1 U935 ( .A(KEYINPUT62), .B(G140), .Z(n1245) );
XOR2_X1 U936 ( .A(n1247), .B(n1164), .Z(n1242) );
AND2_X1 U937 ( .A1(G227), .A2(n1066), .ZN(n1164) );
NAND2_X1 U938 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND2_X1 U939 ( .A1(n1162), .A2(n1250), .ZN(n1249) );
XOR2_X1 U940 ( .A(KEYINPUT45), .B(n1251), .Z(n1248) );
NOR2_X1 U941 ( .A1(n1162), .A2(n1250), .ZN(n1251) );
XNOR2_X1 U942 ( .A(n1252), .B(n1159), .ZN(n1250) );
XOR2_X1 U943 ( .A(n1098), .B(n1253), .Z(n1159) );
NOR2_X1 U944 ( .A1(KEYINPUT39), .A2(n1254), .ZN(n1098) );
INV_X1 U945 ( .A(G128), .ZN(n1254) );
XOR2_X1 U946 ( .A(n1160), .B(KEYINPUT15), .Z(n1252) );
NAND2_X1 U947 ( .A1(n1255), .A2(n1256), .ZN(n1160) );
NAND2_X1 U948 ( .A1(n1257), .A2(n1140), .ZN(n1256) );
XNOR2_X1 U949 ( .A(n1258), .B(n1259), .ZN(n1162) );
XNOR2_X1 U950 ( .A(KEYINPUT32), .B(G134), .ZN(n1258) );
XNOR2_X1 U951 ( .A(KEYINPUT63), .B(n1061), .ZN(n1233) );
AND2_X1 U952 ( .A1(G221), .A2(n1260), .ZN(n1061) );
INV_X1 U953 ( .A(n1130), .ZN(n1200) );
XOR2_X1 U954 ( .A(n1183), .B(KEYINPUT60), .Z(n1130) );
NOR2_X1 U955 ( .A1(n1041), .A2(n1043), .ZN(n1183) );
AND2_X1 U956 ( .A1(G214), .A2(n1261), .ZN(n1043) );
INV_X1 U957 ( .A(n1212), .ZN(n1041) );
XOR2_X1 U958 ( .A(n1262), .B(n1078), .Z(n1212) );
NAND2_X1 U959 ( .A1(G210), .A2(n1261), .ZN(n1078) );
NAND2_X1 U960 ( .A1(n1241), .A2(n1263), .ZN(n1261) );
NAND2_X1 U961 ( .A1(KEYINPUT52), .A2(n1077), .ZN(n1262) );
AND2_X1 U962 ( .A1(n1264), .A2(n1241), .ZN(n1077) );
XOR2_X1 U963 ( .A(n1265), .B(n1168), .Z(n1264) );
XNOR2_X1 U964 ( .A(n1266), .B(n1112), .ZN(n1168) );
XNOR2_X1 U965 ( .A(n1267), .B(n1268), .ZN(n1112) );
XNOR2_X1 U966 ( .A(n1224), .B(G110), .ZN(n1268) );
XNOR2_X1 U967 ( .A(KEYINPUT40), .B(KEYINPUT36), .ZN(n1267) );
XOR2_X1 U968 ( .A(n1269), .B(n1270), .Z(n1266) );
NOR2_X1 U969 ( .A1(n1114), .A2(n1271), .ZN(n1270) );
XNOR2_X1 U970 ( .A(n1116), .B(KEYINPUT12), .ZN(n1271) );
NOR2_X1 U971 ( .A1(n1272), .A2(n1273), .ZN(n1116) );
XNOR2_X1 U972 ( .A(n1140), .B(n1274), .ZN(n1272) );
NAND2_X1 U973 ( .A1(KEYINPUT28), .A2(n1257), .ZN(n1274) );
AND3_X1 U974 ( .A1(n1275), .A2(n1255), .A3(n1273), .ZN(n1114) );
XOR2_X1 U975 ( .A(n1276), .B(n1277), .Z(n1273) );
NAND2_X1 U976 ( .A1(KEYINPUT23), .A2(n1278), .ZN(n1276) );
OR2_X1 U977 ( .A1(n1140), .A2(n1257), .ZN(n1255) );
NAND2_X1 U978 ( .A1(n1279), .A2(n1257), .ZN(n1275) );
XOR2_X1 U979 ( .A(G104), .B(G107), .Z(n1257) );
XNOR2_X1 U980 ( .A(KEYINPUT28), .B(n1140), .ZN(n1279) );
NAND2_X1 U981 ( .A1(G224), .A2(n1066), .ZN(n1269) );
NAND3_X1 U982 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1265) );
NAND2_X1 U983 ( .A1(G125), .A2(n1283), .ZN(n1282) );
OR3_X1 U984 ( .A1(n1283), .A2(G125), .A3(KEYINPUT44), .ZN(n1281) );
NAND2_X1 U985 ( .A1(KEYINPUT47), .A2(n1284), .ZN(n1283) );
INV_X1 U986 ( .A(n1169), .ZN(n1284) );
NAND2_X1 U987 ( .A1(n1169), .A2(KEYINPUT44), .ZN(n1280) );
XOR2_X1 U988 ( .A(G128), .B(n1253), .Z(n1169) );
NOR2_X1 U989 ( .A1(n1206), .A2(n1207), .ZN(n1036) );
XNOR2_X1 U990 ( .A(n1285), .B(G475), .ZN(n1207) );
OR2_X1 U991 ( .A1(n1128), .A2(G902), .ZN(n1285) );
XNOR2_X1 U992 ( .A(n1286), .B(n1287), .ZN(n1128) );
XNOR2_X1 U993 ( .A(n1288), .B(n1289), .ZN(n1287) );
NOR2_X1 U994 ( .A1(KEYINPUT14), .A2(n1290), .ZN(n1289) );
XOR2_X1 U995 ( .A(n1291), .B(n1292), .Z(n1290) );
NOR2_X1 U996 ( .A1(KEYINPUT5), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U997 ( .A(G131), .B(n1294), .ZN(n1291) );
NOR2_X1 U998 ( .A1(KEYINPUT6), .A2(n1295), .ZN(n1294) );
XNOR2_X1 U999 ( .A(G143), .B(n1296), .ZN(n1295) );
AND3_X1 U1000 ( .A1(G214), .A2(n1066), .A3(n1263), .ZN(n1296) );
NAND2_X1 U1001 ( .A1(KEYINPUT37), .A2(n1297), .ZN(n1288) );
XNOR2_X1 U1002 ( .A(n1224), .B(G113), .ZN(n1297) );
XNOR2_X1 U1003 ( .A(G104), .B(KEYINPUT51), .ZN(n1286) );
XNOR2_X1 U1004 ( .A(n1298), .B(G478), .ZN(n1206) );
NAND2_X1 U1005 ( .A1(n1124), .A2(n1241), .ZN(n1298) );
XOR2_X1 U1006 ( .A(n1299), .B(n1300), .Z(n1124) );
XOR2_X1 U1007 ( .A(n1301), .B(n1302), .Z(n1300) );
NAND2_X1 U1008 ( .A1(n1303), .A2(KEYINPUT35), .ZN(n1301) );
XNOR2_X1 U1009 ( .A(G107), .B(n1304), .ZN(n1303) );
XNOR2_X1 U1010 ( .A(n1224), .B(G116), .ZN(n1304) );
INV_X1 U1011 ( .A(G122), .ZN(n1224) );
XOR2_X1 U1012 ( .A(n1305), .B(G143), .Z(n1299) );
NAND2_X1 U1013 ( .A1(G217), .A2(n1306), .ZN(n1305) );
NOR2_X1 U1014 ( .A1(n1226), .A2(n1231), .ZN(n1196) );
INV_X1 U1015 ( .A(n1215), .ZN(n1231) );
XOR2_X1 U1016 ( .A(n1073), .B(n1076), .Z(n1215) );
NAND2_X1 U1017 ( .A1(G217), .A2(n1260), .ZN(n1076) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1241), .ZN(n1260) );
NAND2_X1 U1019 ( .A1(n1307), .A2(n1241), .ZN(n1073) );
XOR2_X1 U1020 ( .A(KEYINPUT22), .B(n1119), .Z(n1307) );
AND2_X1 U1021 ( .A1(n1308), .A2(n1309), .ZN(n1119) );
NAND2_X1 U1022 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
XOR2_X1 U1023 ( .A(n1312), .B(KEYINPUT7), .Z(n1308) );
OR2_X1 U1024 ( .A1(n1311), .A2(n1310), .ZN(n1312) );
XOR2_X1 U1025 ( .A(n1313), .B(n1314), .Z(n1310) );
XNOR2_X1 U1026 ( .A(KEYINPUT58), .B(n1151), .ZN(n1314) );
INV_X1 U1027 ( .A(G110), .ZN(n1151) );
XNOR2_X1 U1028 ( .A(n1293), .B(n1315), .ZN(n1313) );
NOR2_X1 U1029 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
NOR2_X1 U1030 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NOR2_X1 U1031 ( .A1(KEYINPUT0), .A2(G119), .ZN(n1319) );
NOR2_X1 U1032 ( .A1(G128), .A2(n1320), .ZN(n1318) );
AND2_X1 U1033 ( .A1(G119), .A2(KEYINPUT24), .ZN(n1320) );
NOR4_X1 U1034 ( .A1(KEYINPUT24), .A2(KEYINPUT0), .A3(G128), .A4(G119), .ZN(n1316) );
XOR2_X1 U1035 ( .A(G146), .B(n1097), .Z(n1293) );
XOR2_X1 U1036 ( .A(G125), .B(G140), .Z(n1097) );
XNOR2_X1 U1037 ( .A(n1321), .B(G137), .ZN(n1311) );
NAND2_X1 U1038 ( .A1(n1306), .A2(G221), .ZN(n1321) );
AND2_X1 U1039 ( .A1(G234), .A2(n1066), .ZN(n1306) );
INV_X1 U1040 ( .A(n1232), .ZN(n1226) );
XOR2_X1 U1041 ( .A(G472), .B(n1322), .Z(n1232) );
NOR2_X1 U1042 ( .A1(KEYINPUT31), .A2(n1323), .ZN(n1322) );
XNOR2_X1 U1043 ( .A(KEYINPUT21), .B(n1079), .ZN(n1323) );
NAND2_X1 U1044 ( .A1(n1324), .A2(n1241), .ZN(n1079) );
INV_X1 U1045 ( .A(G902), .ZN(n1241) );
XOR2_X1 U1046 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1047 ( .A(n1138), .B(n1327), .Z(n1326) );
NOR2_X1 U1048 ( .A1(KEYINPUT9), .A2(n1139), .ZN(n1327) );
NAND3_X1 U1049 ( .A1(n1263), .A2(n1066), .A3(G210), .ZN(n1139) );
INV_X1 U1050 ( .A(G953), .ZN(n1066) );
INV_X1 U1051 ( .A(G237), .ZN(n1263) );
XOR2_X1 U1052 ( .A(n1328), .B(n1329), .Z(n1138) );
XOR2_X1 U1053 ( .A(n1278), .B(n1330), .Z(n1329) );
XOR2_X1 U1054 ( .A(KEYINPUT32), .B(KEYINPUT29), .Z(n1330) );
XOR2_X1 U1055 ( .A(G113), .B(KEYINPUT18), .Z(n1278) );
XOR2_X1 U1056 ( .A(n1331), .B(n1332), .Z(n1328) );
NOR2_X1 U1057 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
NOR3_X1 U1058 ( .A1(n1335), .A2(G119), .A3(n1227), .ZN(n1334) );
INV_X1 U1059 ( .A(KEYINPUT30), .ZN(n1335) );
NOR2_X1 U1060 ( .A1(KEYINPUT30), .A2(n1277), .ZN(n1333) );
XNOR2_X1 U1061 ( .A(n1227), .B(G119), .ZN(n1277) );
INV_X1 U1062 ( .A(G116), .ZN(n1227) );
XNOR2_X1 U1063 ( .A(n1302), .B(n1336), .ZN(n1331) );
INV_X1 U1064 ( .A(n1095), .ZN(n1336) );
XOR2_X1 U1065 ( .A(n1253), .B(n1259), .Z(n1095) );
XNOR2_X1 U1066 ( .A(n1337), .B(G137), .ZN(n1259) );
INV_X1 U1067 ( .A(G131), .ZN(n1337) );
XOR2_X1 U1068 ( .A(G146), .B(G143), .Z(n1253) );
XNOR2_X1 U1069 ( .A(G134), .B(G128), .ZN(n1302) );
XNOR2_X1 U1070 ( .A(n1338), .B(n1140), .ZN(n1325) );
INV_X1 U1071 ( .A(G101), .ZN(n1140) );
XNOR2_X1 U1072 ( .A(KEYINPUT61), .B(KEYINPUT43), .ZN(n1338) );
endmodule


