//Key = 0001011011101100101010110011000011010110101000101011111011100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288;

XNOR2_X1 U713 ( .A(G107), .B(n987), .ZN(G9) );
NOR2_X1 U714 ( .A1(n988), .A2(n989), .ZN(G75) );
NOR4_X1 U715 ( .A1(n990), .A2(n991), .A3(n992), .A4(n993), .ZN(n989) );
INV_X1 U716 ( .A(G952), .ZN(n992) );
NAND3_X1 U717 ( .A1(n994), .A2(n995), .A3(n996), .ZN(n990) );
NAND2_X1 U718 ( .A1(n997), .A2(n998), .ZN(n996) );
NAND2_X1 U719 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND3_X1 U720 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n1000) );
NAND2_X1 U721 ( .A1(n1004), .A2(n1005), .ZN(n1002) );
NAND2_X1 U722 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
OR2_X1 U723 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND2_X1 U724 ( .A1(n1010), .A2(n1011), .ZN(n1004) );
NAND2_X1 U725 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND2_X1 U726 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND3_X1 U727 ( .A1(n1010), .A2(n1016), .A3(n1006), .ZN(n999) );
NAND3_X1 U728 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1016) );
NAND2_X1 U729 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
XNOR2_X1 U730 ( .A(n1001), .B(KEYINPUT8), .ZN(n1020) );
NAND3_X1 U731 ( .A1(n1022), .A2(n1001), .A3(n1023), .ZN(n1018) );
NAND2_X1 U732 ( .A1(n1003), .A2(n1024), .ZN(n1017) );
OR2_X1 U733 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
INV_X1 U734 ( .A(n1027), .ZN(n997) );
NOR3_X1 U735 ( .A1(n1028), .A2(G953), .A3(n1029), .ZN(n988) );
XOR2_X1 U736 ( .A(KEYINPUT36), .B(G952), .Z(n1029) );
XNOR2_X1 U737 ( .A(KEYINPUT25), .B(n994), .ZN(n1028) );
NAND4_X1 U738 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n994) );
NOR4_X1 U739 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1033) );
XOR2_X1 U740 ( .A(n1038), .B(n1039), .Z(n1037) );
XNOR2_X1 U741 ( .A(KEYINPUT53), .B(n1040), .ZN(n1036) );
XOR2_X1 U742 ( .A(n1041), .B(n1042), .Z(n1035) );
NAND2_X1 U743 ( .A1(KEYINPUT22), .A2(n1043), .ZN(n1041) );
NOR3_X1 U744 ( .A1(n1044), .A2(n1023), .A3(n1045), .ZN(n1032) );
INV_X1 U745 ( .A(n1046), .ZN(n1044) );
XOR2_X1 U746 ( .A(n1047), .B(n1048), .Z(n1030) );
NOR2_X1 U747 ( .A1(G475), .A2(KEYINPUT45), .ZN(n1048) );
XOR2_X1 U748 ( .A(n1049), .B(n1050), .Z(G72) );
NOR2_X1 U749 ( .A1(n1051), .A2(n995), .ZN(n1050) );
NOR2_X1 U750 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U751 ( .A1(n1054), .A2(n1055), .ZN(n1049) );
NAND2_X1 U752 ( .A1(n1056), .A2(n995), .ZN(n1055) );
XOR2_X1 U753 ( .A(n993), .B(n1057), .Z(n1056) );
NAND3_X1 U754 ( .A1(G900), .A2(n1057), .A3(G953), .ZN(n1054) );
XNOR2_X1 U755 ( .A(n1058), .B(n1059), .ZN(n1057) );
XOR2_X1 U756 ( .A(n1060), .B(n1061), .Z(n1059) );
XOR2_X1 U757 ( .A(n1062), .B(G131), .Z(n1061) );
NAND2_X1 U758 ( .A1(KEYINPUT52), .A2(n1063), .ZN(n1062) );
NAND2_X1 U759 ( .A1(KEYINPUT5), .A2(n1064), .ZN(n1060) );
XNOR2_X1 U760 ( .A(n1065), .B(n1066), .ZN(n1058) );
XOR2_X1 U761 ( .A(n1067), .B(n1068), .Z(G69) );
NOR2_X1 U762 ( .A1(KEYINPUT41), .A2(n1069), .ZN(n1068) );
XOR2_X1 U763 ( .A(n1070), .B(n1071), .Z(n1069) );
AND2_X1 U764 ( .A1(n991), .A2(n995), .ZN(n1071) );
NOR2_X1 U765 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
XOR2_X1 U766 ( .A(n1074), .B(n1075), .Z(n1073) );
XOR2_X1 U767 ( .A(n1076), .B(n1077), .Z(n1075) );
NAND2_X1 U768 ( .A1(KEYINPUT26), .A2(n1078), .ZN(n1076) );
XOR2_X1 U769 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U770 ( .A1(G898), .A2(n995), .ZN(n1072) );
NAND2_X1 U771 ( .A1(G953), .A2(n1081), .ZN(n1067) );
NAND2_X1 U772 ( .A1(G898), .A2(G224), .ZN(n1081) );
NOR2_X1 U773 ( .A1(n1082), .A2(n1083), .ZN(G66) );
XNOR2_X1 U774 ( .A(n1084), .B(n1085), .ZN(n1083) );
XNOR2_X1 U775 ( .A(KEYINPUT16), .B(n1086), .ZN(n1085) );
NOR3_X1 U776 ( .A1(n1087), .A2(KEYINPUT24), .A3(n1088), .ZN(n1086) );
NOR2_X1 U777 ( .A1(n1082), .A2(n1089), .ZN(G63) );
XOR2_X1 U778 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR3_X1 U779 ( .A1(n1087), .A2(KEYINPUT11), .A3(n1092), .ZN(n1091) );
NOR2_X1 U780 ( .A1(n1082), .A2(n1093), .ZN(G60) );
XOR2_X1 U781 ( .A(n1094), .B(n1095), .Z(n1093) );
XNOR2_X1 U782 ( .A(n1096), .B(KEYINPUT19), .ZN(n1095) );
NAND3_X1 U783 ( .A1(G475), .A2(n1097), .A3(KEYINPUT18), .ZN(n1096) );
XOR2_X1 U784 ( .A(G104), .B(n1098), .Z(G6) );
NOR3_X1 U785 ( .A1(n1099), .A2(KEYINPUT44), .A3(n1100), .ZN(n1098) );
NOR2_X1 U786 ( .A1(n1082), .A2(n1101), .ZN(G57) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U788 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U789 ( .A1(n1038), .A2(n1087), .ZN(n1104) );
XOR2_X1 U790 ( .A(n1106), .B(n1107), .Z(n1102) );
NOR2_X1 U791 ( .A1(n1082), .A2(n1108), .ZN(G54) );
XOR2_X1 U792 ( .A(n1109), .B(n1110), .Z(n1108) );
XOR2_X1 U793 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U794 ( .A(n1113), .B(n1114), .Z(n1112) );
AND2_X1 U795 ( .A1(G469), .A2(n1097), .ZN(n1113) );
XOR2_X1 U796 ( .A(n1115), .B(n1116), .Z(n1109) );
NOR2_X1 U797 ( .A1(n1117), .A2(KEYINPUT31), .ZN(n1116) );
XOR2_X1 U798 ( .A(n1118), .B(KEYINPUT63), .Z(n1115) );
NOR2_X1 U799 ( .A1(n1082), .A2(n1119), .ZN(G51) );
XOR2_X1 U800 ( .A(n1120), .B(n1121), .Z(n1119) );
AND2_X1 U801 ( .A1(G210), .A2(n1097), .ZN(n1121) );
INV_X1 U802 ( .A(n1087), .ZN(n1097) );
NAND2_X1 U803 ( .A1(G902), .A2(n1122), .ZN(n1087) );
OR2_X1 U804 ( .A1(n991), .A2(n993), .ZN(n1122) );
NAND4_X1 U805 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n993) );
NOR4_X1 U806 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1126) );
INV_X1 U807 ( .A(n1131), .ZN(n1130) );
NAND2_X1 U808 ( .A1(n1021), .A2(n1132), .ZN(n1125) );
NAND2_X1 U809 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U810 ( .A1(n1008), .A2(n1135), .ZN(n1134) );
NAND2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND3_X1 U812 ( .A1(n1025), .A2(n1138), .A3(n1006), .ZN(n1137) );
NAND2_X1 U813 ( .A1(KEYINPUT13), .A2(n1139), .ZN(n1136) );
OR2_X1 U814 ( .A1(n1140), .A2(KEYINPUT13), .ZN(n1133) );
NAND4_X1 U815 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n991) );
AND4_X1 U816 ( .A1(n987), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1144) );
NAND4_X1 U817 ( .A1(n1148), .A2(n1001), .A3(n1149), .A4(n1009), .ZN(n987) );
NOR2_X1 U818 ( .A1(n1150), .A2(n1151), .ZN(n1143) );
NOR2_X1 U819 ( .A1(n1100), .A2(n1099), .ZN(n1151) );
NAND3_X1 U820 ( .A1(n1001), .A2(n1149), .A3(n1008), .ZN(n1099) );
NOR2_X1 U821 ( .A1(n995), .A2(G952), .ZN(n1082) );
XNOR2_X1 U822 ( .A(G146), .B(n1152), .ZN(G48) );
NAND3_X1 U823 ( .A1(n1140), .A2(n1021), .A3(KEYINPUT9), .ZN(n1152) );
AND2_X1 U824 ( .A1(n1139), .A2(n1008), .ZN(n1140) );
XOR2_X1 U825 ( .A(n1123), .B(n1153), .Z(G45) );
NAND2_X1 U826 ( .A1(KEYINPUT3), .A2(G143), .ZN(n1153) );
NAND4_X1 U827 ( .A1(n1040), .A2(n1021), .A3(n1154), .A4(n1155), .ZN(n1123) );
AND2_X1 U828 ( .A1(n1026), .A2(n1156), .ZN(n1155) );
XOR2_X1 U829 ( .A(n1157), .B(n1124), .Z(G42) );
NAND4_X1 U830 ( .A1(n1003), .A2(n1156), .A3(n1008), .A4(n1025), .ZN(n1124) );
XOR2_X1 U831 ( .A(n1158), .B(n1131), .Z(G39) );
NAND3_X1 U832 ( .A1(n1003), .A2(n1010), .A3(n1139), .ZN(n1131) );
XOR2_X1 U833 ( .A(G134), .B(n1128), .Z(G36) );
AND2_X1 U834 ( .A1(n1159), .A2(n1009), .ZN(n1128) );
XOR2_X1 U835 ( .A(G131), .B(n1127), .Z(G33) );
AND2_X1 U836 ( .A1(n1159), .A2(n1008), .ZN(n1127) );
AND3_X1 U837 ( .A1(n1156), .A2(n1026), .A3(n1003), .ZN(n1159) );
NOR2_X1 U838 ( .A1(n1160), .A2(n1023), .ZN(n1003) );
NAND2_X1 U839 ( .A1(n1161), .A2(n1162), .ZN(G30) );
NAND2_X1 U840 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NAND2_X1 U841 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
OR2_X1 U842 ( .A1(KEYINPUT14), .A2(KEYINPUT27), .ZN(n1166) );
NAND3_X1 U843 ( .A1(n1167), .A2(n1168), .A3(KEYINPUT27), .ZN(n1161) );
NAND2_X1 U844 ( .A1(n1129), .A2(n1169), .ZN(n1168) );
INV_X1 U845 ( .A(n1165), .ZN(n1129) );
NAND2_X1 U846 ( .A1(n1170), .A2(n1165), .ZN(n1167) );
NAND3_X1 U847 ( .A1(n1009), .A2(n1021), .A3(n1139), .ZN(n1165) );
AND3_X1 U848 ( .A1(n1171), .A2(n1172), .A3(n1156), .ZN(n1139) );
NOR2_X1 U849 ( .A1(n1012), .A2(n1173), .ZN(n1156) );
INV_X1 U850 ( .A(n1149), .ZN(n1012) );
NAND2_X1 U851 ( .A1(G128), .A2(n1169), .ZN(n1170) );
INV_X1 U852 ( .A(KEYINPUT14), .ZN(n1169) );
XOR2_X1 U853 ( .A(G101), .B(n1150), .Z(G3) );
AND2_X1 U854 ( .A1(n1026), .A2(n1174), .ZN(n1150) );
XOR2_X1 U855 ( .A(n1064), .B(n1175), .Z(G27) );
NAND4_X1 U856 ( .A1(n1008), .A2(n1006), .A3(n1176), .A4(n1021), .ZN(n1175) );
NOR2_X1 U857 ( .A1(n1173), .A2(n1177), .ZN(n1176) );
XNOR2_X1 U858 ( .A(n1025), .B(KEYINPUT29), .ZN(n1177) );
INV_X1 U859 ( .A(n1138), .ZN(n1173) );
NAND2_X1 U860 ( .A1(n1027), .A2(n1178), .ZN(n1138) );
NAND4_X1 U861 ( .A1(G953), .A2(G902), .A3(n1179), .A4(n1053), .ZN(n1178) );
INV_X1 U862 ( .A(G900), .ZN(n1053) );
NAND2_X1 U863 ( .A1(n1180), .A2(n1181), .ZN(G24) );
OR2_X1 U864 ( .A1(n1141), .A2(G122), .ZN(n1181) );
XOR2_X1 U865 ( .A(n1182), .B(KEYINPUT21), .Z(n1180) );
NAND2_X1 U866 ( .A1(G122), .A2(n1141), .ZN(n1182) );
NAND4_X1 U867 ( .A1(n1154), .A2(n1183), .A3(n1040), .A4(n1001), .ZN(n1141) );
NOR2_X1 U868 ( .A1(n1171), .A2(n1172), .ZN(n1001) );
XOR2_X1 U869 ( .A(n1184), .B(n1142), .Z(G21) );
NAND4_X1 U870 ( .A1(n1171), .A2(n1183), .A3(n1172), .A4(n1010), .ZN(n1142) );
INV_X1 U871 ( .A(n1185), .ZN(n1171) );
XOR2_X1 U872 ( .A(n1147), .B(n1186), .Z(G18) );
NAND2_X1 U873 ( .A1(KEYINPUT35), .A2(G116), .ZN(n1186) );
NAND3_X1 U874 ( .A1(n1183), .A2(n1009), .A3(n1026), .ZN(n1147) );
AND2_X1 U875 ( .A1(n1040), .A2(n1187), .ZN(n1009) );
XOR2_X1 U876 ( .A(n1188), .B(n1146), .Z(G15) );
NAND3_X1 U877 ( .A1(n1026), .A2(n1183), .A3(n1008), .ZN(n1146) );
NOR2_X1 U878 ( .A1(n1187), .A2(n1040), .ZN(n1008) );
INV_X1 U879 ( .A(n1154), .ZN(n1187) );
AND2_X1 U880 ( .A1(n1006), .A2(n1148), .ZN(n1183) );
AND2_X1 U881 ( .A1(n1189), .A2(n1015), .ZN(n1006) );
XOR2_X1 U882 ( .A(KEYINPUT0), .B(n1031), .Z(n1189) );
NOR2_X1 U883 ( .A1(n1185), .A2(n1172), .ZN(n1026) );
XOR2_X1 U884 ( .A(n1190), .B(G110), .Z(G12) );
NAND2_X1 U885 ( .A1(KEYINPUT20), .A2(n1145), .ZN(n1190) );
NAND2_X1 U886 ( .A1(n1025), .A2(n1174), .ZN(n1145) );
AND3_X1 U887 ( .A1(n1148), .A2(n1149), .A3(n1010), .ZN(n1174) );
NOR2_X1 U888 ( .A1(n1154), .A2(n1040), .ZN(n1010) );
XOR2_X1 U889 ( .A(n1191), .B(n1192), .Z(n1040) );
NOR2_X1 U890 ( .A1(n1090), .A2(G902), .ZN(n1192) );
AND2_X1 U891 ( .A1(n1193), .A2(n1194), .ZN(n1090) );
NAND2_X1 U892 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XOR2_X1 U893 ( .A(KEYINPUT10), .B(n1197), .Z(n1193) );
NOR2_X1 U894 ( .A1(n1195), .A2(n1196), .ZN(n1197) );
XNOR2_X1 U895 ( .A(n1198), .B(n1199), .ZN(n1196) );
XOR2_X1 U896 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U897 ( .A(G116), .B(G107), .Z(n1201) );
XOR2_X1 U898 ( .A(KEYINPUT32), .B(G128), .Z(n1200) );
XOR2_X1 U899 ( .A(n1063), .B(n1202), .Z(n1198) );
XNOR2_X1 U900 ( .A(n1203), .B(n1204), .ZN(n1202) );
NOR2_X1 U901 ( .A1(G143), .A2(KEYINPUT47), .ZN(n1204) );
NAND2_X1 U902 ( .A1(KEYINPUT51), .A2(n1205), .ZN(n1203) );
AND3_X1 U903 ( .A1(G234), .A2(n995), .A3(G217), .ZN(n1195) );
XOR2_X1 U904 ( .A(n1092), .B(KEYINPUT56), .Z(n1191) );
INV_X1 U905 ( .A(G478), .ZN(n1092) );
XOR2_X1 U906 ( .A(n1206), .B(n1047), .Z(n1154) );
NOR2_X1 U907 ( .A1(n1094), .A2(G902), .ZN(n1047) );
XOR2_X1 U908 ( .A(n1207), .B(n1208), .Z(n1094) );
XOR2_X1 U909 ( .A(n1209), .B(n1210), .Z(n1208) );
XOR2_X1 U910 ( .A(G104), .B(n1211), .Z(n1210) );
NOR2_X1 U911 ( .A1(KEYINPUT55), .A2(n1212), .ZN(n1211) );
XOR2_X1 U912 ( .A(G140), .B(n1213), .Z(n1212) );
XOR2_X1 U913 ( .A(G131), .B(G113), .Z(n1209) );
XOR2_X1 U914 ( .A(n1205), .B(n1214), .Z(n1207) );
XOR2_X1 U915 ( .A(n1215), .B(n1216), .Z(n1214) );
NAND2_X1 U916 ( .A1(KEYINPUT40), .A2(n1217), .ZN(n1216) );
NAND2_X1 U917 ( .A1(n1218), .A2(G214), .ZN(n1215) );
NAND2_X1 U918 ( .A1(KEYINPUT42), .A2(n1219), .ZN(n1206) );
INV_X1 U919 ( .A(G475), .ZN(n1219) );
NOR2_X1 U920 ( .A1(n1220), .A2(n1015), .ZN(n1149) );
XNOR2_X1 U921 ( .A(n1043), .B(n1221), .ZN(n1015) );
INV_X1 U922 ( .A(n1042), .ZN(n1221) );
XNOR2_X1 U923 ( .A(G469), .B(KEYINPUT6), .ZN(n1042) );
NAND2_X1 U924 ( .A1(n1222), .A2(n1223), .ZN(n1043) );
XOR2_X1 U925 ( .A(n1224), .B(n1225), .Z(n1222) );
XNOR2_X1 U926 ( .A(n1117), .B(n1226), .ZN(n1225) );
NOR2_X1 U927 ( .A1(KEYINPUT60), .A2(n1111), .ZN(n1226) );
XOR2_X1 U928 ( .A(n1227), .B(G140), .Z(n1111) );
INV_X1 U929 ( .A(G110), .ZN(n1227) );
NOR2_X1 U930 ( .A1(n1052), .A2(G953), .ZN(n1117) );
INV_X1 U931 ( .A(G227), .ZN(n1052) );
XOR2_X1 U932 ( .A(n1228), .B(KEYINPUT43), .Z(n1224) );
NAND2_X1 U933 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NAND3_X1 U934 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1230) );
NAND2_X1 U935 ( .A1(n1234), .A2(n1235), .ZN(n1232) );
OR2_X1 U936 ( .A1(n1118), .A2(n1235), .ZN(n1231) );
NAND2_X1 U937 ( .A1(n1236), .A2(n1237), .ZN(n1118) );
XOR2_X1 U938 ( .A(n1238), .B(KEYINPUT62), .Z(n1229) );
NAND3_X1 U939 ( .A1(n1114), .A2(n1237), .A3(n1239), .ZN(n1238) );
XOR2_X1 U940 ( .A(n1235), .B(n1236), .Z(n1239) );
INV_X1 U941 ( .A(n1234), .ZN(n1236) );
NOR2_X1 U942 ( .A1(n1065), .A2(n1077), .ZN(n1234) );
INV_X1 U943 ( .A(KEYINPUT12), .ZN(n1235) );
NAND2_X1 U944 ( .A1(n1077), .A2(n1065), .ZN(n1237) );
XNOR2_X1 U945 ( .A(n1240), .B(n1241), .ZN(n1065) );
NAND2_X1 U946 ( .A1(KEYINPUT58), .A2(n1217), .ZN(n1240) );
INV_X1 U947 ( .A(G143), .ZN(n1217) );
XOR2_X1 U948 ( .A(KEYINPUT0), .B(n1014), .Z(n1220) );
INV_X1 U949 ( .A(n1031), .ZN(n1014) );
NAND2_X1 U950 ( .A1(G221), .A2(n1242), .ZN(n1031) );
INV_X1 U951 ( .A(n1100), .ZN(n1148) );
NAND2_X1 U952 ( .A1(n1021), .A2(n1243), .ZN(n1100) );
NAND2_X1 U953 ( .A1(n1027), .A2(n1244), .ZN(n1243) );
NAND4_X1 U954 ( .A1(G953), .A2(G902), .A3(n1179), .A4(n1245), .ZN(n1244) );
INV_X1 U955 ( .A(G898), .ZN(n1245) );
NAND3_X1 U956 ( .A1(n1179), .A2(n995), .A3(G952), .ZN(n1027) );
NAND2_X1 U957 ( .A1(G237), .A2(G234), .ZN(n1179) );
NOR2_X1 U958 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
AND2_X1 U959 ( .A1(G214), .A2(n1246), .ZN(n1023) );
INV_X1 U960 ( .A(n1160), .ZN(n1022) );
NAND2_X1 U961 ( .A1(n1247), .A2(n1046), .ZN(n1160) );
NAND2_X1 U962 ( .A1(n1248), .A2(n1249), .ZN(n1046) );
XNOR2_X1 U963 ( .A(n1045), .B(KEYINPUT7), .ZN(n1247) );
NOR2_X1 U964 ( .A1(n1249), .A2(n1248), .ZN(n1045) );
AND2_X1 U965 ( .A1(n1250), .A2(n1223), .ZN(n1248) );
XOR2_X1 U966 ( .A(KEYINPUT30), .B(n1251), .Z(n1250) );
INV_X1 U967 ( .A(n1120), .ZN(n1251) );
XOR2_X1 U968 ( .A(n1252), .B(n1253), .Z(n1120) );
XOR2_X1 U969 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U970 ( .A(n1256), .B(n1079), .Z(n1255) );
NOR2_X1 U971 ( .A1(KEYINPUT59), .A2(n1184), .ZN(n1079) );
INV_X1 U972 ( .A(G119), .ZN(n1184) );
NAND2_X1 U973 ( .A1(KEYINPUT38), .A2(n1257), .ZN(n1256) );
INV_X1 U974 ( .A(n1077), .ZN(n1257) );
XOR2_X1 U975 ( .A(n1106), .B(n1258), .Z(n1077) );
XOR2_X1 U976 ( .A(G107), .B(G104), .Z(n1258) );
INV_X1 U977 ( .A(G101), .ZN(n1106) );
XOR2_X1 U978 ( .A(n1064), .B(KEYINPUT17), .Z(n1254) );
INV_X1 U979 ( .A(G125), .ZN(n1064) );
XOR2_X1 U980 ( .A(n1259), .B(n1074), .Z(n1252) );
XNOR2_X1 U981 ( .A(n1205), .B(n1260), .ZN(n1074) );
NOR2_X1 U982 ( .A1(G110), .A2(KEYINPUT49), .ZN(n1260) );
XNOR2_X1 U983 ( .A(G122), .B(KEYINPUT39), .ZN(n1205) );
XOR2_X1 U984 ( .A(n1261), .B(n1262), .Z(n1259) );
AND2_X1 U985 ( .A1(n995), .A2(G224), .ZN(n1262) );
NAND2_X1 U986 ( .A1(G210), .A2(n1263), .ZN(n1249) );
XNOR2_X1 U987 ( .A(KEYINPUT57), .B(n1246), .ZN(n1263) );
OR2_X1 U988 ( .A1(G902), .A2(G237), .ZN(n1246) );
AND2_X1 U989 ( .A1(n1172), .A2(n1185), .ZN(n1025) );
NAND2_X1 U990 ( .A1(n1264), .A2(n1265), .ZN(n1185) );
NAND2_X1 U991 ( .A1(n1266), .A2(n1038), .ZN(n1265) );
INV_X1 U992 ( .A(G472), .ZN(n1038) );
XOR2_X1 U993 ( .A(n1039), .B(KEYINPUT1), .Z(n1266) );
NAND2_X1 U994 ( .A1(n1267), .A2(G472), .ZN(n1264) );
XOR2_X1 U995 ( .A(n1039), .B(KEYINPUT48), .Z(n1267) );
NAND2_X1 U996 ( .A1(n1268), .A2(n1223), .ZN(n1039) );
XOR2_X1 U997 ( .A(n1269), .B(n1105), .Z(n1268) );
XNOR2_X1 U998 ( .A(n1261), .B(n1270), .ZN(n1105) );
XOR2_X1 U999 ( .A(G119), .B(n1114), .Z(n1270) );
INV_X1 U1000 ( .A(n1233), .ZN(n1114) );
XOR2_X1 U1001 ( .A(n1063), .B(n1271), .Z(n1233) );
XNOR2_X1 U1002 ( .A(n1272), .B(n1273), .ZN(n1271) );
NOR2_X1 U1003 ( .A1(KEYINPUT4), .A2(n1158), .ZN(n1273) );
NAND2_X1 U1004 ( .A1(KEYINPUT33), .A2(G131), .ZN(n1272) );
XNOR2_X1 U1005 ( .A(G134), .B(KEYINPUT2), .ZN(n1063) );
XOR2_X1 U1006 ( .A(n1274), .B(n1275), .Z(n1261) );
XOR2_X1 U1007 ( .A(KEYINPUT28), .B(G143), .Z(n1275) );
XNOR2_X1 U1008 ( .A(n1080), .B(n1241), .ZN(n1274) );
XOR2_X1 U1009 ( .A(G146), .B(G128), .Z(n1241) );
XNOR2_X1 U1010 ( .A(n1188), .B(n1276), .ZN(n1080) );
XOR2_X1 U1011 ( .A(KEYINPUT54), .B(G116), .Z(n1276) );
INV_X1 U1012 ( .A(G113), .ZN(n1188) );
NAND2_X1 U1013 ( .A1(n1277), .A2(KEYINPUT50), .ZN(n1269) );
XNOR2_X1 U1014 ( .A(n1278), .B(n1107), .ZN(n1277) );
NAND2_X1 U1015 ( .A1(n1218), .A2(G210), .ZN(n1107) );
NOR2_X1 U1016 ( .A1(G953), .A2(G237), .ZN(n1218) );
XNOR2_X1 U1017 ( .A(KEYINPUT23), .B(n1279), .ZN(n1278) );
NOR2_X1 U1018 ( .A1(KEYINPUT34), .A2(n1280), .ZN(n1279) );
XOR2_X1 U1019 ( .A(KEYINPUT46), .B(G101), .Z(n1280) );
XNOR2_X1 U1020 ( .A(n1034), .B(KEYINPUT37), .ZN(n1172) );
XOR2_X1 U1021 ( .A(n1281), .B(n1088), .Z(n1034) );
NAND2_X1 U1022 ( .A1(G217), .A2(n1242), .ZN(n1088) );
NAND2_X1 U1023 ( .A1(G234), .A2(n1223), .ZN(n1242) );
NAND2_X1 U1024 ( .A1(n1084), .A2(n1223), .ZN(n1281) );
INV_X1 U1025 ( .A(G902), .ZN(n1223) );
XNOR2_X1 U1026 ( .A(n1282), .B(n1283), .ZN(n1084) );
XOR2_X1 U1027 ( .A(n1284), .B(n1285), .Z(n1283) );
XOR2_X1 U1028 ( .A(G110), .B(n1286), .Z(n1285) );
AND3_X1 U1029 ( .A1(G221), .A2(n995), .A3(G234), .ZN(n1286) );
INV_X1 U1030 ( .A(G953), .ZN(n995) );
XOR2_X1 U1031 ( .A(KEYINPUT15), .B(G119), .Z(n1284) );
XNOR2_X1 U1032 ( .A(n1066), .B(n1287), .ZN(n1282) );
XOR2_X1 U1033 ( .A(n1288), .B(n1213), .Z(n1287) );
XOR2_X1 U1034 ( .A(G146), .B(G125), .Z(n1213) );
NOR2_X1 U1035 ( .A1(KEYINPUT61), .A2(n1164), .ZN(n1288) );
INV_X1 U1036 ( .A(G128), .ZN(n1164) );
XOR2_X1 U1037 ( .A(n1158), .B(n1157), .Z(n1066) );
INV_X1 U1038 ( .A(G140), .ZN(n1157) );
INV_X1 U1039 ( .A(G137), .ZN(n1158) );
endmodule


