//Key = 1100001110001111010011100000001001001001011110011110000010010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321;

XNOR2_X1 U723 ( .A(G107), .B(n1017), .ZN(G9) );
NAND2_X1 U724 ( .A1(KEYINPUT20), .A2(n1018), .ZN(n1017) );
NOR2_X1 U725 ( .A1(n1019), .A2(n1020), .ZN(G75) );
NOR3_X1 U726 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NAND3_X1 U727 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1021) );
NAND2_X1 U728 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U729 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND3_X1 U730 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
NAND2_X1 U731 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NAND3_X1 U732 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NAND2_X1 U733 ( .A1(n1039), .A2(n1040), .ZN(n1034) );
XNOR2_X1 U734 ( .A(KEYINPUT46), .B(n1041), .ZN(n1040) );
NAND3_X1 U735 ( .A1(n1036), .A2(n1042), .A3(n1043), .ZN(n1029) );
NAND3_X1 U736 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1042) );
NAND2_X1 U737 ( .A1(n1033), .A2(n1047), .ZN(n1046) );
NAND2_X1 U738 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U739 ( .A1(n1038), .A2(n1050), .ZN(n1049) );
NAND2_X1 U740 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U741 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U742 ( .A1(n1031), .A2(n1055), .ZN(n1048) );
NAND2_X1 U743 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U744 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND3_X1 U745 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1045) );
XNOR2_X1 U746 ( .A(n1038), .B(KEYINPUT47), .ZN(n1062) );
XNOR2_X1 U747 ( .A(n1031), .B(KEYINPUT13), .ZN(n1060) );
NAND3_X1 U748 ( .A1(n1031), .A2(n1063), .A3(n1038), .ZN(n1044) );
INV_X1 U749 ( .A(n1064), .ZN(n1027) );
NOR3_X1 U750 ( .A1(n1065), .A2(G953), .A3(G952), .ZN(n1019) );
INV_X1 U751 ( .A(n1024), .ZN(n1065) );
NAND4_X1 U752 ( .A1(n1033), .A2(n1031), .A3(n1066), .A4(n1067), .ZN(n1024) );
NOR4_X1 U753 ( .A1(n1068), .A2(n1058), .A3(n1069), .A4(n1070), .ZN(n1067) );
XNOR2_X1 U754 ( .A(n1071), .B(n1072), .ZN(n1070) );
XNOR2_X1 U755 ( .A(n1073), .B(KEYINPUT14), .ZN(n1071) );
XNOR2_X1 U756 ( .A(n1037), .B(KEYINPUT63), .ZN(n1066) );
XOR2_X1 U757 ( .A(n1074), .B(n1075), .Z(G72) );
NOR2_X1 U758 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR3_X1 U759 ( .A1(n1022), .A2(n1078), .A3(n1079), .ZN(n1077) );
NOR2_X1 U760 ( .A1(G900), .A2(n1025), .ZN(n1078) );
NOR2_X1 U761 ( .A1(n1080), .A2(n1081), .ZN(n1076) );
XOR2_X1 U762 ( .A(n1082), .B(KEYINPUT45), .Z(n1081) );
NAND2_X1 U763 ( .A1(n1079), .A2(n1025), .ZN(n1082) );
XNOR2_X1 U764 ( .A(n1083), .B(n1084), .ZN(n1079) );
XOR2_X1 U765 ( .A(n1085), .B(n1086), .Z(n1084) );
XNOR2_X1 U766 ( .A(KEYINPUT32), .B(KEYINPUT17), .ZN(n1086) );
XNOR2_X1 U767 ( .A(KEYINPUT34), .B(KEYINPUT33), .ZN(n1085) );
XOR2_X1 U768 ( .A(n1087), .B(n1088), .Z(n1083) );
XNOR2_X1 U769 ( .A(G131), .B(n1089), .ZN(n1088) );
XNOR2_X1 U770 ( .A(n1090), .B(n1091), .ZN(n1087) );
NAND3_X1 U771 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1090) );
NAND2_X1 U772 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
INV_X1 U773 ( .A(KEYINPUT43), .ZN(n1096) );
NAND3_X1 U774 ( .A1(KEYINPUT43), .A2(n1097), .A3(n1098), .ZN(n1093) );
OR2_X1 U775 ( .A1(n1098), .A2(n1097), .ZN(n1092) );
NOR2_X1 U776 ( .A1(KEYINPUT23), .A2(n1095), .ZN(n1097) );
INV_X1 U777 ( .A(n1022), .ZN(n1080) );
NAND2_X1 U778 ( .A1(G953), .A2(n1099), .ZN(n1074) );
NAND2_X1 U779 ( .A1(G227), .A2(n1100), .ZN(n1099) );
XNOR2_X1 U780 ( .A(KEYINPUT28), .B(n1101), .ZN(n1100) );
NAND2_X1 U781 ( .A1(n1102), .A2(n1103), .ZN(G69) );
NAND2_X1 U782 ( .A1(n1104), .A2(n1025), .ZN(n1103) );
XNOR2_X1 U783 ( .A(n1023), .B(n1105), .ZN(n1104) );
NAND2_X1 U784 ( .A1(n1106), .A2(G953), .ZN(n1102) );
NAND2_X1 U785 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U786 ( .A1(n1105), .A2(n1109), .ZN(n1108) );
NAND2_X1 U787 ( .A1(G224), .A2(n1110), .ZN(n1107) );
NAND2_X1 U788 ( .A1(G898), .A2(n1105), .ZN(n1110) );
NAND2_X1 U789 ( .A1(n1111), .A2(n1112), .ZN(n1105) );
NAND2_X1 U790 ( .A1(G953), .A2(n1113), .ZN(n1112) );
XOR2_X1 U791 ( .A(n1114), .B(n1115), .Z(n1111) );
NOR2_X1 U792 ( .A1(n1116), .A2(n1117), .ZN(G66) );
XOR2_X1 U793 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND2_X1 U794 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
NOR2_X1 U795 ( .A1(n1116), .A2(n1122), .ZN(G63) );
XOR2_X1 U796 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U797 ( .A1(KEYINPUT10), .A2(n1125), .ZN(n1124) );
AND2_X1 U798 ( .A1(G478), .A2(n1120), .ZN(n1123) );
NOR2_X1 U799 ( .A1(n1116), .A2(n1126), .ZN(G60) );
XOR2_X1 U800 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U801 ( .A(n1129), .B(KEYINPUT29), .Z(n1127) );
NAND2_X1 U802 ( .A1(n1120), .A2(G475), .ZN(n1129) );
XNOR2_X1 U803 ( .A(G104), .B(n1130), .ZN(G6) );
NOR2_X1 U804 ( .A1(n1116), .A2(n1131), .ZN(G57) );
XOR2_X1 U805 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U806 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U807 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U808 ( .A1(KEYINPUT41), .A2(n1138), .ZN(n1137) );
NOR2_X1 U809 ( .A1(KEYINPUT2), .A2(n1139), .ZN(n1134) );
XOR2_X1 U810 ( .A(n1140), .B(n1141), .Z(n1132) );
NOR2_X1 U811 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
AND2_X1 U812 ( .A1(KEYINPUT24), .A2(n1144), .ZN(n1143) );
NOR2_X1 U813 ( .A1(KEYINPUT37), .A2(n1144), .ZN(n1142) );
NAND2_X1 U814 ( .A1(n1120), .A2(G472), .ZN(n1144) );
XOR2_X1 U815 ( .A(n1145), .B(n1146), .Z(n1140) );
NAND2_X1 U816 ( .A1(KEYINPUT1), .A2(n1147), .ZN(n1145) );
INV_X1 U817 ( .A(G101), .ZN(n1147) );
NOR2_X1 U818 ( .A1(n1116), .A2(n1148), .ZN(G54) );
XOR2_X1 U819 ( .A(n1149), .B(n1150), .Z(n1148) );
XNOR2_X1 U820 ( .A(n1146), .B(n1151), .ZN(n1150) );
XOR2_X1 U821 ( .A(n1152), .B(n1153), .Z(n1149) );
XOR2_X1 U822 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND2_X1 U823 ( .A1(KEYINPUT12), .A2(n1156), .ZN(n1154) );
NAND2_X1 U824 ( .A1(n1120), .A2(G469), .ZN(n1152) );
INV_X1 U825 ( .A(n1157), .ZN(n1120) );
NOR2_X1 U826 ( .A1(n1116), .A2(n1158), .ZN(G51) );
NOR2_X1 U827 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U828 ( .A(KEYINPUT9), .B(n1161), .Z(n1160) );
NOR2_X1 U829 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U830 ( .A(KEYINPUT35), .B(n1164), .Z(n1163) );
NOR2_X1 U831 ( .A1(n1072), .A2(n1157), .ZN(n1164) );
INV_X1 U832 ( .A(n1165), .ZN(n1162) );
NOR3_X1 U833 ( .A1(n1165), .A2(n1072), .A3(n1157), .ZN(n1159) );
NAND2_X1 U834 ( .A1(G902), .A2(n1166), .ZN(n1157) );
OR2_X1 U835 ( .A1(n1023), .A2(n1022), .ZN(n1166) );
NAND4_X1 U836 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1022) );
AND3_X1 U837 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1170) );
NAND2_X1 U838 ( .A1(n1038), .A2(n1174), .ZN(n1169) );
NAND3_X1 U839 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1174) );
NAND2_X1 U840 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND3_X1 U841 ( .A1(n1180), .A2(n1033), .A3(n1181), .ZN(n1175) );
NAND4_X1 U842 ( .A1(n1182), .A2(n1130), .A3(n1183), .A4(n1184), .ZN(n1023) );
NOR3_X1 U843 ( .A1(n1018), .A2(n1185), .A3(n1186), .ZN(n1184) );
AND3_X1 U844 ( .A1(n1043), .A2(n1063), .A3(n1187), .ZN(n1018) );
NAND2_X1 U845 ( .A1(n1188), .A2(n1189), .ZN(n1183) );
NAND2_X1 U846 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND4_X1 U847 ( .A1(n1039), .A2(n1033), .A3(n1179), .A4(n1192), .ZN(n1191) );
XNOR2_X1 U848 ( .A(KEYINPUT59), .B(n1193), .ZN(n1190) );
NAND3_X1 U849 ( .A1(n1043), .A2(n1187), .A3(n1061), .ZN(n1130) );
NAND2_X1 U850 ( .A1(n1194), .A2(n1195), .ZN(n1182) );
OR2_X1 U851 ( .A1(n1061), .A2(n1063), .ZN(n1195) );
XNOR2_X1 U852 ( .A(n1196), .B(n1197), .ZN(n1165) );
NAND2_X1 U853 ( .A1(KEYINPUT50), .A2(n1198), .ZN(n1196) );
XOR2_X1 U854 ( .A(KEYINPUT21), .B(n1199), .Z(n1198) );
AND2_X1 U855 ( .A1(G953), .A2(n1200), .ZN(n1116) );
XOR2_X1 U856 ( .A(KEYINPUT36), .B(G952), .Z(n1200) );
XNOR2_X1 U857 ( .A(G146), .B(n1167), .ZN(G48) );
NAND2_X1 U858 ( .A1(n1201), .A2(n1061), .ZN(n1167) );
XNOR2_X1 U859 ( .A(G143), .B(n1168), .ZN(G45) );
NAND4_X1 U860 ( .A1(n1181), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1168) );
XOR2_X1 U861 ( .A(G140), .B(n1205), .Z(G42) );
NOR3_X1 U862 ( .A1(n1206), .A2(n1207), .A3(n1051), .ZN(n1205) );
INV_X1 U863 ( .A(n1179), .ZN(n1051) );
XNOR2_X1 U864 ( .A(n1038), .B(KEYINPUT40), .ZN(n1207) );
XNOR2_X1 U865 ( .A(G137), .B(n1208), .ZN(G39) );
NAND2_X1 U866 ( .A1(n1209), .A2(n1038), .ZN(n1208) );
XOR2_X1 U867 ( .A(n1210), .B(KEYINPUT15), .Z(n1209) );
NAND3_X1 U868 ( .A1(n1033), .A2(n1211), .A3(n1181), .ZN(n1210) );
XOR2_X1 U869 ( .A(KEYINPUT54), .B(n1180), .Z(n1211) );
XNOR2_X1 U870 ( .A(n1098), .B(n1212), .ZN(G36) );
NOR2_X1 U871 ( .A1(n1213), .A2(n1041), .ZN(n1212) );
XOR2_X1 U872 ( .A(n1176), .B(KEYINPUT4), .Z(n1213) );
NAND3_X1 U873 ( .A1(n1039), .A2(n1063), .A3(n1181), .ZN(n1176) );
XNOR2_X1 U874 ( .A(G131), .B(n1171), .ZN(G33) );
NAND4_X1 U875 ( .A1(n1038), .A2(n1181), .A3(n1039), .A4(n1061), .ZN(n1171) );
INV_X1 U876 ( .A(n1041), .ZN(n1038) );
NAND2_X1 U877 ( .A1(n1059), .A2(n1214), .ZN(n1041) );
XNOR2_X1 U878 ( .A(G128), .B(n1173), .ZN(G30) );
NAND2_X1 U879 ( .A1(n1201), .A2(n1063), .ZN(n1173) );
AND3_X1 U880 ( .A1(n1180), .A2(n1188), .A3(n1181), .ZN(n1201) );
AND2_X1 U881 ( .A1(n1179), .A2(n1215), .ZN(n1181) );
XNOR2_X1 U882 ( .A(G101), .B(n1216), .ZN(G3) );
NAND4_X1 U883 ( .A1(n1217), .A2(n1202), .A3(n1033), .A4(n1179), .ZN(n1216) );
XNOR2_X1 U884 ( .A(n1218), .B(KEYINPUT31), .ZN(n1217) );
XNOR2_X1 U885 ( .A(G125), .B(n1172), .ZN(G27) );
NAND3_X1 U886 ( .A1(n1031), .A2(n1188), .A3(n1178), .ZN(n1172) );
INV_X1 U887 ( .A(n1206), .ZN(n1178) );
NAND4_X1 U888 ( .A1(n1061), .A2(n1036), .A3(n1037), .A4(n1215), .ZN(n1206) );
NAND2_X1 U889 ( .A1(n1064), .A2(n1219), .ZN(n1215) );
NAND4_X1 U890 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1101), .ZN(n1219) );
INV_X1 U891 ( .A(G900), .ZN(n1101) );
XOR2_X1 U892 ( .A(G122), .B(n1221), .Z(G24) );
NOR2_X1 U893 ( .A1(n1056), .A2(n1193), .ZN(n1221) );
NAND4_X1 U894 ( .A1(n1043), .A2(n1036), .A3(n1031), .A4(n1222), .ZN(n1193) );
NOR3_X1 U895 ( .A1(n1223), .A2(n1218), .A3(n1224), .ZN(n1222) );
XOR2_X1 U896 ( .A(n1186), .B(n1225), .Z(G21) );
NOR2_X1 U897 ( .A1(KEYINPUT26), .A2(n1226), .ZN(n1225) );
AND4_X1 U898 ( .A1(n1180), .A2(n1033), .A3(n1227), .A4(n1031), .ZN(n1186) );
NOR2_X1 U899 ( .A1(n1218), .A2(n1056), .ZN(n1227) );
INV_X1 U900 ( .A(n1188), .ZN(n1056) );
INV_X1 U901 ( .A(n1192), .ZN(n1218) );
NOR2_X1 U902 ( .A1(n1043), .A2(n1036), .ZN(n1180) );
INV_X1 U903 ( .A(n1037), .ZN(n1043) );
XNOR2_X1 U904 ( .A(G116), .B(n1228), .ZN(G18) );
NAND3_X1 U905 ( .A1(n1194), .A2(n1063), .A3(KEYINPUT7), .ZN(n1228) );
NOR2_X1 U906 ( .A1(n1204), .A2(n1223), .ZN(n1063) );
INV_X1 U907 ( .A(n1203), .ZN(n1223) );
INV_X1 U908 ( .A(n1229), .ZN(n1194) );
XNOR2_X1 U909 ( .A(n1230), .B(n1231), .ZN(G15) );
NOR2_X1 U910 ( .A1(n1232), .A2(n1229), .ZN(n1231) );
NAND3_X1 U911 ( .A1(n1031), .A2(n1192), .A3(n1202), .ZN(n1229) );
AND2_X1 U912 ( .A1(n1039), .A2(n1188), .ZN(n1202) );
NOR2_X1 U913 ( .A1(n1037), .A2(n1036), .ZN(n1039) );
NOR2_X1 U914 ( .A1(n1233), .A2(n1053), .ZN(n1031) );
XNOR2_X1 U915 ( .A(n1061), .B(KEYINPUT18), .ZN(n1232) );
NOR2_X1 U916 ( .A1(n1203), .A2(n1224), .ZN(n1061) );
INV_X1 U917 ( .A(n1204), .ZN(n1224) );
XOR2_X1 U918 ( .A(G110), .B(n1185), .Z(G12) );
AND3_X1 U919 ( .A1(n1187), .A2(n1037), .A3(n1033), .ZN(n1185) );
NOR2_X1 U920 ( .A1(n1203), .A2(n1204), .ZN(n1033) );
XNOR2_X1 U921 ( .A(n1234), .B(G475), .ZN(n1204) );
NAND2_X1 U922 ( .A1(n1128), .A2(n1235), .ZN(n1234) );
XNOR2_X1 U923 ( .A(n1236), .B(n1237), .ZN(n1128) );
XOR2_X1 U924 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U925 ( .A(G131), .B(G104), .Z(n1239) );
NOR2_X1 U926 ( .A1(KEYINPUT38), .A2(n1240), .ZN(n1238) );
XOR2_X1 U927 ( .A(G143), .B(n1241), .Z(n1240) );
AND3_X1 U928 ( .A1(G214), .A2(n1025), .A3(n1242), .ZN(n1241) );
XOR2_X1 U929 ( .A(n1243), .B(n1244), .Z(n1236) );
NOR3_X1 U930 ( .A1(n1245), .A2(KEYINPUT58), .A3(n1246), .ZN(n1244) );
AND2_X1 U931 ( .A1(n1230), .A2(G122), .ZN(n1246) );
XOR2_X1 U932 ( .A(KEYINPUT3), .B(n1247), .Z(n1245) );
NOR2_X1 U933 ( .A1(G122), .A2(n1230), .ZN(n1247) );
NAND2_X1 U934 ( .A1(n1248), .A2(n1249), .ZN(n1243) );
NAND2_X1 U935 ( .A1(G146), .A2(n1250), .ZN(n1249) );
XOR2_X1 U936 ( .A(n1251), .B(KEYINPUT27), .Z(n1248) );
NAND2_X1 U937 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
XNOR2_X1 U938 ( .A(n1250), .B(KEYINPUT55), .ZN(n1252) );
XNOR2_X1 U939 ( .A(n1254), .B(G478), .ZN(n1203) );
NAND2_X1 U940 ( .A1(n1125), .A2(n1235), .ZN(n1254) );
XOR2_X1 U941 ( .A(n1255), .B(n1256), .Z(n1125) );
XOR2_X1 U942 ( .A(n1257), .B(n1258), .Z(n1256) );
XOR2_X1 U943 ( .A(G107), .B(n1259), .Z(n1258) );
NOR2_X1 U944 ( .A1(KEYINPUT61), .A2(n1260), .ZN(n1259) );
XNOR2_X1 U945 ( .A(G116), .B(n1261), .ZN(n1260) );
XOR2_X1 U946 ( .A(KEYINPUT5), .B(G122), .Z(n1261) );
XOR2_X1 U947 ( .A(KEYINPUT62), .B(KEYINPUT19), .Z(n1257) );
XOR2_X1 U948 ( .A(n1262), .B(n1263), .Z(n1255) );
XNOR2_X1 U949 ( .A(n1264), .B(n1265), .ZN(n1262) );
NAND2_X1 U950 ( .A1(KEYINPUT39), .A2(n1098), .ZN(n1265) );
INV_X1 U951 ( .A(G134), .ZN(n1098) );
NAND3_X1 U952 ( .A1(G217), .A2(n1266), .A3(KEYINPUT48), .ZN(n1264) );
XNOR2_X1 U953 ( .A(n1267), .B(n1121), .ZN(n1037) );
AND2_X1 U954 ( .A1(G217), .A2(n1268), .ZN(n1121) );
NAND2_X1 U955 ( .A1(n1119), .A2(n1235), .ZN(n1267) );
XNOR2_X1 U956 ( .A(n1269), .B(n1270), .ZN(n1119) );
XOR2_X1 U957 ( .A(n1271), .B(n1272), .Z(n1270) );
XNOR2_X1 U958 ( .A(n1226), .B(G110), .ZN(n1272) );
INV_X1 U959 ( .A(G119), .ZN(n1226) );
XNOR2_X1 U960 ( .A(n1253), .B(G128), .ZN(n1271) );
XOR2_X1 U961 ( .A(n1273), .B(n1095), .Z(n1269) );
XNOR2_X1 U962 ( .A(n1274), .B(n1091), .ZN(n1273) );
INV_X1 U963 ( .A(n1250), .ZN(n1091) );
XOR2_X1 U964 ( .A(G140), .B(n1275), .Z(n1250) );
NAND3_X1 U965 ( .A1(n1266), .A2(G221), .A3(KEYINPUT49), .ZN(n1274) );
AND2_X1 U966 ( .A1(G234), .A2(n1025), .ZN(n1266) );
AND4_X1 U967 ( .A1(n1188), .A2(n1179), .A3(n1036), .A4(n1192), .ZN(n1187) );
NAND2_X1 U968 ( .A1(n1064), .A2(n1276), .ZN(n1192) );
NAND4_X1 U969 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1113), .ZN(n1276) );
INV_X1 U970 ( .A(G898), .ZN(n1113) );
NAND3_X1 U971 ( .A1(n1220), .A2(n1025), .A3(G952), .ZN(n1064) );
NAND2_X1 U972 ( .A1(G237), .A2(G234), .ZN(n1220) );
NOR2_X1 U973 ( .A1(n1277), .A2(n1069), .ZN(n1036) );
NOR2_X1 U974 ( .A1(n1278), .A2(G472), .ZN(n1069) );
XOR2_X1 U975 ( .A(n1068), .B(KEYINPUT11), .Z(n1277) );
AND2_X1 U976 ( .A1(G472), .A2(n1278), .ZN(n1068) );
NAND2_X1 U977 ( .A1(n1279), .A2(n1235), .ZN(n1278) );
XOR2_X1 U978 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U979 ( .A(n1139), .B(n1282), .Z(n1281) );
XNOR2_X1 U980 ( .A(n1283), .B(n1146), .ZN(n1282) );
NAND2_X1 U981 ( .A1(KEYINPUT30), .A2(n1138), .ZN(n1283) );
XOR2_X1 U982 ( .A(n1284), .B(n1285), .Z(n1138) );
NAND2_X1 U983 ( .A1(KEYINPUT56), .A2(n1230), .ZN(n1284) );
XOR2_X1 U984 ( .A(n1136), .B(n1286), .Z(n1280) );
XNOR2_X1 U985 ( .A(G101), .B(KEYINPUT44), .ZN(n1286) );
NAND3_X1 U986 ( .A1(n1242), .A2(n1025), .A3(G210), .ZN(n1136) );
NOR2_X1 U987 ( .A1(n1054), .A2(n1053), .ZN(n1179) );
AND2_X1 U988 ( .A1(G221), .A2(n1268), .ZN(n1053) );
NAND2_X1 U989 ( .A1(G234), .A2(n1235), .ZN(n1268) );
INV_X1 U990 ( .A(n1233), .ZN(n1054) );
XNOR2_X1 U991 ( .A(n1287), .B(G469), .ZN(n1233) );
NAND2_X1 U992 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
XNOR2_X1 U993 ( .A(n1156), .B(n1290), .ZN(n1289) );
XOR2_X1 U994 ( .A(n1291), .B(n1155), .Z(n1290) );
AND2_X1 U995 ( .A1(G227), .A2(n1025), .ZN(n1155) );
INV_X1 U996 ( .A(G953), .ZN(n1025) );
NAND2_X1 U997 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND2_X1 U998 ( .A1(n1151), .A2(n1146), .ZN(n1293) );
XOR2_X1 U999 ( .A(KEYINPUT42), .B(n1294), .Z(n1292) );
NOR2_X1 U1000 ( .A1(n1151), .A2(n1146), .ZN(n1294) );
XNOR2_X1 U1001 ( .A(n1295), .B(n1296), .ZN(n1146) );
NOR2_X1 U1002 ( .A1(n1095), .A2(n1297), .ZN(n1296) );
XOR2_X1 U1003 ( .A(KEYINPUT60), .B(KEYINPUT16), .Z(n1297) );
XOR2_X1 U1004 ( .A(G137), .B(KEYINPUT52), .Z(n1095) );
XNOR2_X1 U1005 ( .A(G131), .B(G134), .ZN(n1295) );
XNOR2_X1 U1006 ( .A(n1298), .B(n1299), .ZN(n1151) );
XNOR2_X1 U1007 ( .A(G101), .B(n1089), .ZN(n1299) );
NAND2_X1 U1008 ( .A1(n1300), .A2(n1301), .ZN(n1089) );
NAND2_X1 U1009 ( .A1(G128), .A2(n1302), .ZN(n1301) );
XOR2_X1 U1010 ( .A(n1303), .B(KEYINPUT53), .Z(n1300) );
OR2_X1 U1011 ( .A1(n1302), .A2(G128), .ZN(n1303) );
NAND2_X1 U1012 ( .A1(n1304), .A2(n1305), .ZN(n1302) );
NAND2_X1 U1013 ( .A1(G143), .A2(n1253), .ZN(n1305) );
XOR2_X1 U1014 ( .A(KEYINPUT0), .B(n1306), .Z(n1304) );
NOR2_X1 U1015 ( .A1(G143), .A2(n1253), .ZN(n1306) );
INV_X1 U1016 ( .A(G146), .ZN(n1253) );
XOR2_X1 U1017 ( .A(G140), .B(G110), .Z(n1156) );
XNOR2_X1 U1018 ( .A(KEYINPUT6), .B(n1235), .ZN(n1288) );
NOR2_X1 U1019 ( .A1(n1059), .A2(n1058), .ZN(n1188) );
INV_X1 U1020 ( .A(n1214), .ZN(n1058) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1307), .ZN(n1214) );
XNOR2_X1 U1022 ( .A(n1072), .B(n1308), .ZN(n1059) );
NOR2_X1 U1023 ( .A1(n1073), .A2(KEYINPUT57), .ZN(n1308) );
AND2_X1 U1024 ( .A1(n1309), .A2(n1235), .ZN(n1073) );
XOR2_X1 U1025 ( .A(n1310), .B(n1199), .Z(n1309) );
XOR2_X1 U1026 ( .A(n1139), .B(n1275), .Z(n1199) );
XOR2_X1 U1027 ( .A(G125), .B(KEYINPUT51), .Z(n1275) );
XOR2_X1 U1028 ( .A(G146), .B(n1263), .Z(n1139) );
XOR2_X1 U1029 ( .A(G128), .B(G143), .Z(n1263) );
XNOR2_X1 U1030 ( .A(n1197), .B(KEYINPUT25), .ZN(n1310) );
XNOR2_X1 U1031 ( .A(n1311), .B(n1312), .ZN(n1197) );
NOR2_X1 U1032 ( .A1(G953), .A2(n1109), .ZN(n1312) );
INV_X1 U1033 ( .A(G224), .ZN(n1109) );
NAND2_X1 U1034 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
NAND2_X1 U1035 ( .A1(n1114), .A2(n1115), .ZN(n1314) );
XOR2_X1 U1036 ( .A(KEYINPUT22), .B(n1315), .Z(n1313) );
NOR2_X1 U1037 ( .A1(n1114), .A2(n1115), .ZN(n1315) );
XOR2_X1 U1038 ( .A(G110), .B(G122), .Z(n1115) );
XOR2_X1 U1039 ( .A(n1316), .B(n1285), .Z(n1114) );
XNOR2_X1 U1040 ( .A(n1317), .B(G119), .ZN(n1285) );
INV_X1 U1041 ( .A(G116), .ZN(n1317) );
XNOR2_X1 U1042 ( .A(n1318), .B(n1230), .ZN(n1316) );
INV_X1 U1043 ( .A(G113), .ZN(n1230) );
NAND2_X1 U1044 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
NAND2_X1 U1045 ( .A1(G101), .A2(n1298), .ZN(n1320) );
XOR2_X1 U1046 ( .A(KEYINPUT8), .B(n1321), .Z(n1319) );
NOR2_X1 U1047 ( .A1(G101), .A2(n1298), .ZN(n1321) );
XOR2_X1 U1048 ( .A(G104), .B(G107), .Z(n1298) );
NAND2_X1 U1049 ( .A1(G210), .A2(n1307), .ZN(n1072) );
NAND2_X1 U1050 ( .A1(n1242), .A2(n1235), .ZN(n1307) );
INV_X1 U1051 ( .A(G902), .ZN(n1235) );
INV_X1 U1052 ( .A(G237), .ZN(n1242) );
endmodule


