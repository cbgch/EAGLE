//Key = 0001010010110001010110100101001101001000101011100001111101000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342;

XOR2_X1 U733 ( .A(G107), .B(n1011), .Z(G9) );
NOR2_X1 U734 ( .A1(n1012), .A2(n1013), .ZN(G75) );
NOR3_X1 U735 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NOR2_X1 U736 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NOR2_X1 U737 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR2_X1 U738 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
INV_X1 U739 ( .A(n1023), .ZN(n1022) );
NOR2_X1 U740 ( .A1(n1024), .A2(n1025), .ZN(n1021) );
NOR2_X1 U741 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR3_X1 U742 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1026) );
NOR3_X1 U743 ( .A1(n1031), .A2(KEYINPUT46), .A3(n1032), .ZN(n1030) );
NOR2_X1 U744 ( .A1(n1033), .A2(n1034), .ZN(n1029) );
NOR3_X1 U745 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1033) );
AND2_X1 U746 ( .A1(n1038), .A2(KEYINPUT46), .ZN(n1037) );
AND2_X1 U747 ( .A1(n1039), .A2(KEYINPUT26), .ZN(n1036) );
NOR2_X1 U748 ( .A1(KEYINPUT49), .A2(n1040), .ZN(n1035) );
NOR2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1028) );
NOR2_X1 U750 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
INV_X1 U751 ( .A(n1045), .ZN(n1044) );
NOR3_X1 U752 ( .A1(n1046), .A2(KEYINPUT26), .A3(n1047), .ZN(n1043) );
NOR3_X1 U753 ( .A1(n1034), .A2(n1048), .A3(n1042), .ZN(n1024) );
NOR2_X1 U754 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR4_X1 U755 ( .A1(n1051), .A2(n1027), .A3(n1042), .A4(n1034), .ZN(n1019) );
INV_X1 U756 ( .A(n1052), .ZN(n1027) );
NOR2_X1 U757 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
XNOR2_X1 U758 ( .A(n1055), .B(KEYINPUT52), .ZN(n1054) );
NOR2_X1 U759 ( .A1(n1056), .A2(n1057), .ZN(n1053) );
NAND3_X1 U760 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1014) );
NAND3_X1 U761 ( .A1(n1023), .A2(n1061), .A3(KEYINPUT49), .ZN(n1060) );
NAND4_X1 U762 ( .A1(n1062), .A2(n1031), .A3(n1063), .A4(n1052), .ZN(n1061) );
AND3_X1 U763 ( .A1(n1058), .A2(n1059), .A3(n1064), .ZN(n1012) );
NAND4_X1 U764 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1058) );
NOR3_X1 U765 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1068) );
XNOR2_X1 U766 ( .A(n1072), .B(n1073), .ZN(n1071) );
XOR2_X1 U767 ( .A(KEYINPUT37), .B(KEYINPUT12), .Z(n1073) );
NAND3_X1 U768 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1069) );
XNOR2_X1 U769 ( .A(n1077), .B(KEYINPUT7), .ZN(n1076) );
OR2_X1 U770 ( .A1(n1031), .A2(KEYINPUT23), .ZN(n1075) );
NAND2_X1 U771 ( .A1(KEYINPUT23), .A2(n1078), .ZN(n1074) );
NAND3_X1 U772 ( .A1(n1079), .A2(n1046), .A3(G469), .ZN(n1078) );
NOR3_X1 U773 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1067) );
NAND2_X1 U774 ( .A1(G478), .A2(n1083), .ZN(n1066) );
XOR2_X1 U775 ( .A(n1084), .B(n1085), .Z(n1065) );
NAND2_X1 U776 ( .A1(KEYINPUT25), .A2(n1086), .ZN(n1085) );
NAND2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(G72) );
NAND2_X1 U778 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U779 ( .A1(G953), .A2(n1091), .ZN(n1089) );
NAND2_X1 U780 ( .A1(G900), .A2(G227), .ZN(n1091) );
NAND2_X1 U781 ( .A1(n1092), .A2(n1093), .ZN(n1087) );
NAND2_X1 U782 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U783 ( .A1(G953), .A2(n1096), .ZN(n1095) );
INV_X1 U784 ( .A(n1090), .ZN(n1092) );
NAND2_X1 U785 ( .A1(n1097), .A2(KEYINPUT15), .ZN(n1090) );
XOR2_X1 U786 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U787 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XOR2_X1 U788 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND2_X1 U789 ( .A1(n1104), .A2(KEYINPUT30), .ZN(n1102) );
XNOR2_X1 U790 ( .A(n1105), .B(n1106), .ZN(n1104) );
XNOR2_X1 U791 ( .A(n1107), .B(KEYINPUT0), .ZN(n1105) );
NAND2_X1 U792 ( .A1(n1059), .A2(n1108), .ZN(n1098) );
NAND2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U794 ( .A(n1111), .B(n1112), .Z(G69) );
XOR2_X1 U795 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U796 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U797 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U798 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U799 ( .A(n1121), .B(n1122), .Z(n1117) );
NOR2_X1 U800 ( .A1(KEYINPUT4), .A2(n1123), .ZN(n1122) );
XNOR2_X1 U801 ( .A(G122), .B(n1124), .ZN(n1123) );
NOR2_X1 U802 ( .A1(G898), .A2(n1059), .ZN(n1115) );
NOR2_X1 U803 ( .A1(n1125), .A2(n1126), .ZN(n1113) );
XNOR2_X1 U804 ( .A(KEYINPUT32), .B(n1059), .ZN(n1126) );
NOR2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
XNOR2_X1 U806 ( .A(KEYINPUT56), .B(n1129), .ZN(n1128) );
NOR2_X1 U807 ( .A1(n1130), .A2(n1059), .ZN(n1111) );
AND2_X1 U808 ( .A1(G224), .A2(G898), .ZN(n1130) );
NOR2_X1 U809 ( .A1(n1131), .A2(n1132), .ZN(G66) );
XNOR2_X1 U810 ( .A(n1133), .B(n1134), .ZN(n1132) );
NOR2_X1 U811 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NOR2_X1 U812 ( .A1(n1131), .A2(n1137), .ZN(G63) );
XNOR2_X1 U813 ( .A(n1138), .B(n1139), .ZN(n1137) );
AND2_X1 U814 ( .A1(G478), .A2(n1140), .ZN(n1139) );
NOR2_X1 U815 ( .A1(n1131), .A2(n1141), .ZN(G60) );
XNOR2_X1 U816 ( .A(n1142), .B(n1143), .ZN(n1141) );
AND2_X1 U817 ( .A1(G475), .A2(n1140), .ZN(n1142) );
XNOR2_X1 U818 ( .A(G104), .B(n1129), .ZN(G6) );
NOR3_X1 U819 ( .A1(n1131), .A2(n1144), .A3(n1145), .ZN(G57) );
NOR2_X1 U820 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XNOR2_X1 U821 ( .A(n1148), .B(KEYINPUT42), .ZN(n1147) );
INV_X1 U822 ( .A(G101), .ZN(n1146) );
NOR2_X1 U823 ( .A1(G101), .A2(n1149), .ZN(n1144) );
XNOR2_X1 U824 ( .A(KEYINPUT17), .B(n1150), .ZN(n1149) );
INV_X1 U825 ( .A(n1148), .ZN(n1150) );
XNOR2_X1 U826 ( .A(n1151), .B(n1152), .ZN(n1148) );
XOR2_X1 U827 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND2_X1 U829 ( .A1(n1140), .A2(G472), .ZN(n1156) );
NOR2_X1 U830 ( .A1(KEYINPUT35), .A2(n1107), .ZN(n1153) );
XNOR2_X1 U831 ( .A(n1157), .B(n1106), .ZN(n1151) );
NAND2_X1 U832 ( .A1(KEYINPUT44), .A2(n1158), .ZN(n1157) );
NOR2_X1 U833 ( .A1(n1131), .A2(n1159), .ZN(G54) );
XOR2_X1 U834 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U835 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U836 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U837 ( .A1(KEYINPUT61), .A2(n1166), .ZN(n1165) );
AND2_X1 U838 ( .A1(G469), .A2(n1140), .ZN(n1162) );
XOR2_X1 U839 ( .A(n1167), .B(n1168), .Z(n1160) );
XNOR2_X1 U840 ( .A(n1169), .B(n1170), .ZN(n1167) );
NOR2_X1 U841 ( .A1(KEYINPUT59), .A2(n1171), .ZN(n1170) );
NOR2_X1 U842 ( .A1(n1131), .A2(n1172), .ZN(G51) );
XOR2_X1 U843 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U844 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U845 ( .A1(n1140), .A2(G210), .ZN(n1176) );
INV_X1 U846 ( .A(n1136), .ZN(n1140) );
NAND2_X1 U847 ( .A1(G902), .A2(n1016), .ZN(n1136) );
NAND4_X1 U848 ( .A1(n1177), .A2(n1178), .A3(n1109), .A4(n1129), .ZN(n1016) );
NAND3_X1 U849 ( .A1(n1179), .A2(n1039), .A3(n1050), .ZN(n1129) );
AND4_X1 U850 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1109) );
NOR4_X1 U851 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1183) );
NAND2_X1 U852 ( .A1(n1188), .A2(n1189), .ZN(n1182) );
INV_X1 U853 ( .A(n1190), .ZN(n1189) );
XNOR2_X1 U854 ( .A(n1038), .B(KEYINPUT11), .ZN(n1188) );
INV_X1 U855 ( .A(n1127), .ZN(n1178) );
NAND4_X1 U856 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1127) );
NOR3_X1 U857 ( .A1(n1195), .A2(n1011), .A3(n1196), .ZN(n1194) );
AND3_X1 U858 ( .A1(n1049), .A2(n1039), .A3(n1179), .ZN(n1011) );
NAND2_X1 U859 ( .A1(n1055), .A2(n1197), .ZN(n1193) );
NAND2_X1 U860 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U861 ( .A(n1200), .B(KEYINPUT24), .Z(n1198) );
NAND2_X1 U862 ( .A1(n1201), .A2(n1050), .ZN(n1200) );
XOR2_X1 U863 ( .A(n1110), .B(KEYINPUT41), .Z(n1177) );
NAND2_X1 U864 ( .A1(n1202), .A2(n1203), .ZN(n1175) );
NAND2_X1 U865 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NOR2_X1 U866 ( .A1(n1059), .A2(G952), .ZN(n1131) );
XNOR2_X1 U867 ( .A(G146), .B(n1180), .ZN(G48) );
NAND4_X1 U868 ( .A1(n1206), .A2(n1207), .A3(n1050), .A4(n1055), .ZN(n1180) );
XOR2_X1 U869 ( .A(n1208), .B(G143), .Z(G45) );
NAND2_X1 U870 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
OR2_X1 U871 ( .A1(n1110), .A2(KEYINPUT6), .ZN(n1210) );
OR2_X1 U872 ( .A1(n1211), .A2(n1212), .ZN(n1110) );
NAND3_X1 U873 ( .A1(n1055), .A2(n1211), .A3(KEYINPUT6), .ZN(n1209) );
NAND4_X1 U874 ( .A1(n1206), .A2(n1038), .A3(n1070), .A4(n1213), .ZN(n1211) );
XOR2_X1 U875 ( .A(n1214), .B(n1187), .Z(G42) );
NOR2_X1 U876 ( .A1(n1190), .A2(n1040), .ZN(n1187) );
NAND2_X1 U877 ( .A1(KEYINPUT45), .A2(n1215), .ZN(n1214) );
XOR2_X1 U878 ( .A(n1216), .B(n1186), .Z(G39) );
AND4_X1 U879 ( .A1(n1206), .A2(n1023), .A3(n1207), .A4(n1052), .ZN(n1186) );
NAND2_X1 U880 ( .A1(KEYINPUT19), .A2(n1217), .ZN(n1216) );
XNOR2_X1 U881 ( .A(G134), .B(n1181), .ZN(G36) );
NAND4_X1 U882 ( .A1(n1206), .A2(n1023), .A3(n1038), .A4(n1049), .ZN(n1181) );
XOR2_X1 U883 ( .A(n1218), .B(n1219), .Z(G33) );
XOR2_X1 U884 ( .A(KEYINPUT21), .B(G131), .Z(n1219) );
NOR2_X1 U885 ( .A1(n1032), .A2(n1190), .ZN(n1218) );
NAND3_X1 U886 ( .A1(n1023), .A2(n1050), .A3(n1206), .ZN(n1190) );
NOR2_X1 U887 ( .A1(n1045), .A2(n1220), .ZN(n1206) );
NOR2_X1 U888 ( .A1(n1056), .A2(n1080), .ZN(n1023) );
INV_X1 U889 ( .A(n1221), .ZN(n1056) );
XOR2_X1 U890 ( .A(n1222), .B(n1185), .Z(G30) );
AND4_X1 U891 ( .A1(n1223), .A2(n1224), .A3(n1055), .A4(n1225), .ZN(n1185) );
NOR2_X1 U892 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
NAND2_X1 U893 ( .A1(KEYINPUT63), .A2(n1228), .ZN(n1222) );
INV_X1 U894 ( .A(G128), .ZN(n1228) );
XOR2_X1 U895 ( .A(n1191), .B(n1229), .Z(G3) );
NOR2_X1 U896 ( .A1(G101), .A2(KEYINPUT38), .ZN(n1229) );
NAND3_X1 U897 ( .A1(n1179), .A2(n1052), .A3(n1038), .ZN(n1191) );
XOR2_X1 U898 ( .A(G125), .B(n1184), .Z(G27) );
AND3_X1 U899 ( .A1(n1031), .A2(n1063), .A3(n1230), .ZN(n1184) );
NOR3_X1 U900 ( .A1(n1231), .A2(n1220), .A3(n1212), .ZN(n1230) );
INV_X1 U901 ( .A(n1224), .ZN(n1220) );
NAND2_X1 U902 ( .A1(n1018), .A2(n1232), .ZN(n1224) );
OR3_X1 U903 ( .A1(n1233), .A2(n1234), .A3(n1094), .ZN(n1232) );
INV_X1 U904 ( .A(n1100), .ZN(n1094) );
NOR2_X1 U905 ( .A1(n1059), .A2(G900), .ZN(n1100) );
XNOR2_X1 U906 ( .A(G122), .B(n1192), .ZN(G24) );
NAND3_X1 U907 ( .A1(n1235), .A2(n1039), .A3(n1236), .ZN(n1192) );
NOR3_X1 U908 ( .A1(n1212), .A2(n1237), .A3(n1238), .ZN(n1236) );
INV_X1 U909 ( .A(n1055), .ZN(n1212) );
INV_X1 U910 ( .A(n1042), .ZN(n1039) );
NAND2_X1 U911 ( .A1(n1072), .A2(n1239), .ZN(n1042) );
NAND2_X1 U912 ( .A1(n1240), .A2(n1241), .ZN(G21) );
NAND2_X1 U913 ( .A1(G119), .A2(n1242), .ZN(n1241) );
XOR2_X1 U914 ( .A(n1243), .B(KEYINPUT48), .Z(n1240) );
OR2_X1 U915 ( .A1(n1242), .A2(G119), .ZN(n1243) );
NAND2_X1 U916 ( .A1(n1244), .A2(n1055), .ZN(n1242) );
XOR2_X1 U917 ( .A(n1199), .B(KEYINPUT33), .Z(n1244) );
NAND3_X1 U918 ( .A1(n1235), .A2(n1052), .A3(n1207), .ZN(n1199) );
INV_X1 U919 ( .A(n1227), .ZN(n1207) );
NAND2_X1 U920 ( .A1(n1245), .A2(n1246), .ZN(n1227) );
XOR2_X1 U921 ( .A(G116), .B(n1195), .Z(G18) );
AND3_X1 U922 ( .A1(n1049), .A2(n1055), .A3(n1201), .ZN(n1195) );
INV_X1 U923 ( .A(n1226), .ZN(n1049) );
NAND2_X1 U924 ( .A1(n1247), .A2(n1213), .ZN(n1226) );
XNOR2_X1 U925 ( .A(KEYINPUT51), .B(n1238), .ZN(n1247) );
XNOR2_X1 U926 ( .A(G113), .B(n1248), .ZN(G15) );
NAND3_X1 U927 ( .A1(n1055), .A2(n1249), .A3(n1201), .ZN(n1248) );
AND2_X1 U928 ( .A1(n1038), .A2(n1235), .ZN(n1201) );
AND2_X1 U929 ( .A1(n1031), .A2(n1250), .ZN(n1235) );
INV_X1 U930 ( .A(n1034), .ZN(n1031) );
NAND2_X1 U931 ( .A1(n1251), .A2(n1046), .ZN(n1034) );
INV_X1 U932 ( .A(n1047), .ZN(n1251) );
INV_X1 U933 ( .A(n1032), .ZN(n1038) );
NAND2_X1 U934 ( .A1(n1072), .A2(n1246), .ZN(n1032) );
XNOR2_X1 U935 ( .A(KEYINPUT47), .B(n1231), .ZN(n1249) );
XOR2_X1 U936 ( .A(G110), .B(n1196), .Z(G12) );
AND3_X1 U937 ( .A1(n1179), .A2(n1052), .A3(n1063), .ZN(n1196) );
INV_X1 U938 ( .A(n1040), .ZN(n1063) );
NAND2_X1 U939 ( .A1(n1245), .A2(n1239), .ZN(n1040) );
XOR2_X1 U940 ( .A(n1246), .B(KEYINPUT10), .Z(n1239) );
XOR2_X1 U941 ( .A(n1084), .B(n1086), .Z(n1246) );
INV_X1 U942 ( .A(G472), .ZN(n1086) );
NAND2_X1 U943 ( .A1(n1252), .A2(n1253), .ZN(n1084) );
NAND2_X1 U944 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U945 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XOR2_X1 U946 ( .A(KEYINPUT20), .B(n1258), .Z(n1254) );
NOR2_X1 U947 ( .A1(n1256), .A2(n1257), .ZN(n1258) );
XNOR2_X1 U948 ( .A(n1259), .B(G101), .ZN(n1257) );
NAND2_X1 U949 ( .A1(KEYINPUT22), .A2(n1155), .ZN(n1259) );
NAND3_X1 U950 ( .A1(n1260), .A2(n1059), .A3(G210), .ZN(n1155) );
XNOR2_X1 U951 ( .A(n1261), .B(n1158), .ZN(n1256) );
XOR2_X1 U952 ( .A(n1262), .B(n1263), .Z(n1158) );
NAND2_X1 U953 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
NAND2_X1 U954 ( .A1(n1120), .A2(n1266), .ZN(n1265) );
INV_X1 U955 ( .A(KEYINPUT50), .ZN(n1266) );
XNOR2_X1 U956 ( .A(G119), .B(n1267), .ZN(n1120) );
NAND3_X1 U957 ( .A1(n1267), .A2(n1268), .A3(KEYINPUT50), .ZN(n1264) );
NAND2_X1 U958 ( .A1(n1269), .A2(n1270), .ZN(n1261) );
NAND2_X1 U959 ( .A1(n1169), .A2(n1107), .ZN(n1270) );
XOR2_X1 U960 ( .A(n1271), .B(KEYINPUT1), .Z(n1269) );
NAND2_X1 U961 ( .A1(n1106), .A2(n1272), .ZN(n1271) );
INV_X1 U962 ( .A(n1107), .ZN(n1272) );
XNOR2_X1 U963 ( .A(n1072), .B(KEYINPUT28), .ZN(n1245) );
XNOR2_X1 U964 ( .A(n1273), .B(n1135), .ZN(n1072) );
NAND2_X1 U965 ( .A1(G217), .A2(n1274), .ZN(n1135) );
NAND2_X1 U966 ( .A1(n1134), .A2(n1252), .ZN(n1273) );
XOR2_X1 U967 ( .A(n1275), .B(n1276), .Z(n1134) );
NOR2_X1 U968 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
XOR2_X1 U969 ( .A(KEYINPUT58), .B(n1279), .Z(n1278) );
NOR4_X1 U970 ( .A1(G953), .A2(n1280), .A3(n1281), .A4(n1217), .ZN(n1279) );
NOR2_X1 U971 ( .A1(n1282), .A2(G137), .ZN(n1277) );
NOR3_X1 U972 ( .A1(n1281), .A2(G953), .A3(n1280), .ZN(n1282) );
INV_X1 U973 ( .A(G221), .ZN(n1281) );
NAND2_X1 U974 ( .A1(n1283), .A2(n1284), .ZN(n1275) );
NAND2_X1 U975 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
XOR2_X1 U976 ( .A(KEYINPUT53), .B(n1287), .Z(n1283) );
NOR2_X1 U977 ( .A1(n1286), .A2(n1285), .ZN(n1287) );
XNOR2_X1 U978 ( .A(G146), .B(n1103), .ZN(n1285) );
XNOR2_X1 U979 ( .A(G125), .B(n1215), .ZN(n1103) );
XOR2_X1 U980 ( .A(n1288), .B(n1289), .Z(n1286) );
XNOR2_X1 U981 ( .A(G128), .B(KEYINPUT13), .ZN(n1288) );
NAND2_X1 U982 ( .A1(n1290), .A2(n1291), .ZN(n1052) );
OR2_X1 U983 ( .A1(n1231), .A2(KEYINPUT51), .ZN(n1291) );
INV_X1 U984 ( .A(n1050), .ZN(n1231) );
NOR2_X1 U985 ( .A1(n1213), .A2(n1238), .ZN(n1050) );
INV_X1 U986 ( .A(n1237), .ZN(n1213) );
NAND3_X1 U987 ( .A1(n1237), .A2(n1238), .A3(KEYINPUT51), .ZN(n1290) );
INV_X1 U988 ( .A(n1070), .ZN(n1238) );
XNOR2_X1 U989 ( .A(n1292), .B(G475), .ZN(n1070) );
NAND2_X1 U990 ( .A1(n1143), .A2(n1252), .ZN(n1292) );
XOR2_X1 U991 ( .A(n1293), .B(n1294), .Z(n1143) );
XOR2_X1 U992 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U993 ( .A(n1297), .B(n1298), .Z(n1296) );
NOR2_X1 U994 ( .A1(G125), .A2(KEYINPUT2), .ZN(n1298) );
AND3_X1 U995 ( .A1(G214), .A2(n1059), .A3(n1260), .ZN(n1297) );
XOR2_X1 U996 ( .A(n1299), .B(n1300), .Z(n1293) );
XNOR2_X1 U997 ( .A(n1215), .B(G131), .ZN(n1300) );
XNOR2_X1 U998 ( .A(G104), .B(n1301), .ZN(n1299) );
NOR2_X1 U999 ( .A1(KEYINPUT9), .A2(n1302), .ZN(n1301) );
XNOR2_X1 U1000 ( .A(G113), .B(G122), .ZN(n1302) );
NOR2_X1 U1001 ( .A1(n1303), .A2(n1082), .ZN(n1237) );
NOR2_X1 U1002 ( .A1(n1083), .A2(G478), .ZN(n1082) );
AND2_X1 U1003 ( .A1(n1304), .A2(G478), .ZN(n1303) );
XOR2_X1 U1004 ( .A(n1083), .B(KEYINPUT18), .Z(n1304) );
NAND2_X1 U1005 ( .A1(n1252), .A2(n1305), .ZN(n1083) );
XNOR2_X1 U1006 ( .A(KEYINPUT34), .B(n1306), .ZN(n1305) );
INV_X1 U1007 ( .A(n1138), .ZN(n1306) );
XNOR2_X1 U1008 ( .A(n1307), .B(n1308), .ZN(n1138) );
XOR2_X1 U1009 ( .A(n1309), .B(n1310), .Z(n1308) );
XNOR2_X1 U1010 ( .A(n1311), .B(n1312), .ZN(n1310) );
NOR4_X1 U1011 ( .A1(KEYINPUT39), .A2(G953), .A3(n1280), .A4(n1313), .ZN(n1312) );
INV_X1 U1012 ( .A(G217), .ZN(n1313) );
NAND2_X1 U1013 ( .A1(KEYINPUT54), .A2(G128), .ZN(n1311) );
XNOR2_X1 U1014 ( .A(G107), .B(n1314), .ZN(n1307) );
XOR2_X1 U1015 ( .A(G143), .B(G134), .Z(n1314) );
AND3_X1 U1016 ( .A1(n1223), .A2(n1250), .A3(n1055), .ZN(n1179) );
NOR2_X1 U1017 ( .A1(n1221), .A2(n1080), .ZN(n1055) );
INV_X1 U1018 ( .A(n1057), .ZN(n1080) );
NAND2_X1 U1019 ( .A1(G214), .A2(n1315), .ZN(n1057) );
NOR2_X1 U1020 ( .A1(n1077), .A2(n1081), .ZN(n1221) );
NOR2_X1 U1021 ( .A1(n1316), .A2(n1317), .ZN(n1081) );
AND2_X1 U1022 ( .A1(G210), .A2(n1315), .ZN(n1317) );
AND3_X1 U1023 ( .A1(n1315), .A2(n1316), .A3(G210), .ZN(n1077) );
NAND2_X1 U1024 ( .A1(n1252), .A2(n1318), .ZN(n1316) );
XOR2_X1 U1025 ( .A(n1319), .B(n1173), .Z(n1318) );
XOR2_X1 U1026 ( .A(n1320), .B(n1321), .Z(n1173) );
XOR2_X1 U1027 ( .A(n1289), .B(n1309), .Z(n1321) );
XOR2_X1 U1028 ( .A(G122), .B(n1267), .Z(n1309) );
XOR2_X1 U1029 ( .A(G116), .B(KEYINPUT62), .Z(n1267) );
XNOR2_X1 U1030 ( .A(n1268), .B(n1124), .ZN(n1289) );
INV_X1 U1031 ( .A(G119), .ZN(n1268) );
XOR2_X1 U1032 ( .A(n1322), .B(n1121), .Z(n1320) );
AND2_X1 U1033 ( .A1(KEYINPUT31), .A2(n1263), .ZN(n1121) );
INV_X1 U1034 ( .A(G113), .ZN(n1263) );
NAND2_X1 U1035 ( .A1(KEYINPUT36), .A2(n1119), .ZN(n1322) );
NAND2_X1 U1036 ( .A1(n1323), .A2(n1324), .ZN(n1119) );
OR2_X1 U1037 ( .A1(n1325), .A2(G101), .ZN(n1324) );
XOR2_X1 U1038 ( .A(n1326), .B(KEYINPUT43), .Z(n1323) );
NAND2_X1 U1039 ( .A1(G101), .A2(n1325), .ZN(n1326) );
XOR2_X1 U1040 ( .A(G104), .B(G107), .Z(n1325) );
NAND3_X1 U1041 ( .A1(n1327), .A2(n1328), .A3(KEYINPUT27), .ZN(n1319) );
NAND2_X1 U1042 ( .A1(n1204), .A2(n1329), .ZN(n1328) );
XNOR2_X1 U1043 ( .A(KEYINPUT57), .B(n1205), .ZN(n1329) );
XNOR2_X1 U1044 ( .A(KEYINPUT8), .B(n1202), .ZN(n1327) );
OR2_X1 U1045 ( .A1(n1205), .A2(n1204), .ZN(n1202) );
AND2_X1 U1046 ( .A1(G224), .A2(n1059), .ZN(n1204) );
XNOR2_X1 U1047 ( .A(G125), .B(n1107), .ZN(n1205) );
NAND2_X1 U1048 ( .A1(n1233), .A2(n1260), .ZN(n1315) );
NAND2_X1 U1049 ( .A1(n1330), .A2(n1018), .ZN(n1250) );
INV_X1 U1050 ( .A(n1062), .ZN(n1018) );
NOR3_X1 U1051 ( .A1(n1234), .A2(G953), .A3(n1064), .ZN(n1062) );
INV_X1 U1052 ( .A(G952), .ZN(n1064) );
XOR2_X1 U1053 ( .A(KEYINPUT5), .B(n1331), .Z(n1330) );
NOR4_X1 U1054 ( .A1(G898), .A2(n1234), .A3(n1233), .A4(n1059), .ZN(n1331) );
INV_X1 U1055 ( .A(G953), .ZN(n1059) );
INV_X1 U1056 ( .A(G902), .ZN(n1233) );
NOR2_X1 U1057 ( .A1(n1260), .A2(n1280), .ZN(n1234) );
INV_X1 U1058 ( .A(G234), .ZN(n1280) );
INV_X1 U1059 ( .A(G237), .ZN(n1260) );
XNOR2_X1 U1060 ( .A(n1045), .B(KEYINPUT60), .ZN(n1223) );
NAND2_X1 U1061 ( .A1(n1047), .A2(n1046), .ZN(n1045) );
NAND2_X1 U1062 ( .A1(G221), .A2(n1274), .ZN(n1046) );
NAND2_X1 U1063 ( .A1(n1332), .A2(G234), .ZN(n1274) );
XNOR2_X1 U1064 ( .A(G902), .B(KEYINPUT29), .ZN(n1332) );
XNOR2_X1 U1065 ( .A(n1079), .B(G469), .ZN(n1047) );
NAND2_X1 U1066 ( .A1(n1252), .A2(n1333), .ZN(n1079) );
XOR2_X1 U1067 ( .A(n1334), .B(n1335), .Z(n1333) );
XNOR2_X1 U1068 ( .A(n1166), .B(n1106), .ZN(n1335) );
INV_X1 U1069 ( .A(n1169), .ZN(n1106) );
XOR2_X1 U1070 ( .A(G131), .B(n1336), .Z(n1169) );
XNOR2_X1 U1071 ( .A(n1217), .B(G134), .ZN(n1336) );
INV_X1 U1072 ( .A(G137), .ZN(n1217) );
XOR2_X1 U1073 ( .A(n1337), .B(n1338), .Z(n1166) );
XNOR2_X1 U1074 ( .A(n1339), .B(n1107), .ZN(n1338) );
XOR2_X1 U1075 ( .A(G128), .B(n1295), .Z(n1107) );
XOR2_X1 U1076 ( .A(G143), .B(G146), .Z(n1295) );
NAND2_X1 U1077 ( .A1(KEYINPUT3), .A2(n1340), .ZN(n1339) );
INV_X1 U1078 ( .A(G104), .ZN(n1340) );
XNOR2_X1 U1079 ( .A(G107), .B(G101), .ZN(n1337) );
XOR2_X1 U1080 ( .A(n1341), .B(n1164), .Z(n1334) );
NOR2_X1 U1081 ( .A1(n1096), .A2(G953), .ZN(n1164) );
INV_X1 U1082 ( .A(G227), .ZN(n1096) );
NAND2_X1 U1083 ( .A1(KEYINPUT55), .A2(n1342), .ZN(n1341) );
XNOR2_X1 U1084 ( .A(n1171), .B(n1168), .ZN(n1342) );
XNOR2_X1 U1085 ( .A(n1215), .B(KEYINPUT16), .ZN(n1168) );
INV_X1 U1086 ( .A(G140), .ZN(n1215) );
INV_X1 U1087 ( .A(n1124), .ZN(n1171) );
XOR2_X1 U1088 ( .A(G110), .B(KEYINPUT40), .Z(n1124) );
XNOR2_X1 U1089 ( .A(G902), .B(KEYINPUT14), .ZN(n1252) );
endmodule


