//Key = 1010011000101000010011000010000000111010011111011001000111110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311;

XNOR2_X1 U729 ( .A(n993), .B(n994), .ZN(G9) );
NAND2_X1 U730 ( .A1(KEYINPUT42), .A2(n995), .ZN(n993) );
OR2_X1 U731 ( .A1(n996), .A2(n997), .ZN(n995) );
NOR2_X1 U732 ( .A1(n998), .A2(n999), .ZN(G75) );
NOR4_X1 U733 ( .A1(n1000), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(n999) );
NOR2_X1 U734 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NOR2_X1 U735 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NOR2_X1 U736 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NOR2_X1 U737 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NOR2_X1 U738 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR2_X1 U739 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR2_X1 U740 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR2_X1 U741 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
AND3_X1 U742 ( .A1(n1020), .A2(n1021), .A3(G214), .ZN(n1018) );
INV_X1 U743 ( .A(n1022), .ZN(n1020) );
NOR2_X1 U744 ( .A1(n1023), .A2(n1024), .ZN(n1014) );
NOR2_X1 U745 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR4_X1 U746 ( .A1(KEYINPUT47), .A2(n1027), .A3(n1028), .A4(n1024), .ZN(n1010) );
NOR3_X1 U747 ( .A1(n1024), .A2(n1029), .A3(n1017), .ZN(n1006) );
NOR2_X1 U748 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR2_X1 U749 ( .A1(n1032), .A2(n1013), .ZN(n1031) );
NOR3_X1 U750 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1032) );
AND3_X1 U751 ( .A1(KEYINPUT17), .A2(n1036), .A3(n1037), .ZN(n1035) );
NOR2_X1 U752 ( .A1(KEYINPUT17), .A2(n1009), .ZN(n1034) );
NOR2_X1 U753 ( .A1(n1038), .A2(n1009), .ZN(n1030) );
NOR2_X1 U754 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
AND2_X1 U755 ( .A1(n1041), .A2(KEYINPUT47), .ZN(n1039) );
INV_X1 U756 ( .A(n1042), .ZN(n1004) );
NOR3_X1 U757 ( .A1(n1001), .A2(G952), .A3(n1002), .ZN(n998) );
AND4_X1 U758 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1002) );
NOR4_X1 U759 ( .A1(n1047), .A2(n1048), .A3(n1024), .A4(n1049), .ZN(n1046) );
XNOR2_X1 U760 ( .A(KEYINPUT9), .B(n1050), .ZN(n1049) );
XOR2_X1 U761 ( .A(n1051), .B(KEYINPUT0), .Z(n1047) );
NOR2_X1 U762 ( .A1(n1052), .A2(n1037), .ZN(n1045) );
NAND2_X1 U763 ( .A1(G478), .A2(n1053), .ZN(n1044) );
XOR2_X1 U764 ( .A(G469), .B(n1054), .Z(n1043) );
NOR2_X1 U765 ( .A1(n1055), .A2(KEYINPUT31), .ZN(n1054) );
NAND2_X1 U766 ( .A1(n1056), .A2(n1057), .ZN(G72) );
NAND2_X1 U767 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
OR2_X1 U768 ( .A1(n1060), .A2(G227), .ZN(n1059) );
NAND3_X1 U769 ( .A1(G953), .A2(n1061), .A3(n1062), .ZN(n1056) );
INV_X1 U770 ( .A(n1058), .ZN(n1062) );
XNOR2_X1 U771 ( .A(n1063), .B(n1064), .ZN(n1058) );
NOR2_X1 U772 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U773 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR2_X1 U774 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
INV_X1 U775 ( .A(n1071), .ZN(n1070) );
NOR2_X1 U776 ( .A1(KEYINPUT22), .A2(n1072), .ZN(n1069) );
NOR2_X1 U777 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U778 ( .A1(n1075), .A2(n1076), .ZN(n1067) );
INV_X1 U779 ( .A(n1073), .ZN(n1076) );
NOR2_X1 U780 ( .A1(n1077), .A2(n1074), .ZN(n1075) );
INV_X1 U781 ( .A(KEYINPUT55), .ZN(n1074) );
NOR2_X1 U782 ( .A1(KEYINPUT22), .A2(n1071), .ZN(n1077) );
XNOR2_X1 U783 ( .A(n1078), .B(n1079), .ZN(n1071) );
NOR2_X1 U784 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U785 ( .A(KEYINPUT49), .B(KEYINPUT1), .Z(n1081) );
NOR2_X1 U786 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
XOR2_X1 U787 ( .A(n1084), .B(KEYINPUT38), .Z(n1083) );
NAND2_X1 U788 ( .A1(G131), .A2(n1085), .ZN(n1084) );
OR2_X1 U789 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR3_X1 U790 ( .A1(n1086), .A2(G131), .A3(n1087), .ZN(n1082) );
XNOR2_X1 U791 ( .A(n1088), .B(KEYINPUT3), .ZN(n1086) );
NAND2_X1 U792 ( .A1(G137), .A2(n1089), .ZN(n1088) );
NAND3_X1 U793 ( .A1(n1090), .A2(n1060), .A3(KEYINPUT57), .ZN(n1063) );
NAND2_X1 U794 ( .A1(G900), .A2(G227), .ZN(n1061) );
NAND2_X1 U795 ( .A1(n1091), .A2(n1092), .ZN(G69) );
NAND2_X1 U796 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U797 ( .A1(n1095), .A2(n1096), .ZN(n1091) );
NAND2_X1 U798 ( .A1(n1097), .A2(n1094), .ZN(n1096) );
NAND2_X1 U799 ( .A1(G953), .A2(n1098), .ZN(n1094) );
INV_X1 U800 ( .A(n1093), .ZN(n1095) );
XNOR2_X1 U801 ( .A(n1099), .B(n1100), .ZN(n1093) );
NOR2_X1 U802 ( .A1(G953), .A2(n1101), .ZN(n1100) );
NOR2_X1 U803 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XNOR2_X1 U804 ( .A(n1104), .B(KEYINPUT32), .ZN(n1102) );
NAND2_X1 U805 ( .A1(n1105), .A2(n1097), .ZN(n1099) );
INV_X1 U806 ( .A(n1106), .ZN(n1097) );
XNOR2_X1 U807 ( .A(n1107), .B(n1108), .ZN(n1105) );
NOR2_X1 U808 ( .A1(n1109), .A2(n1110), .ZN(G66) );
XNOR2_X1 U809 ( .A(n1111), .B(n1112), .ZN(n1110) );
NOR2_X1 U810 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U811 ( .A1(n1109), .A2(n1115), .ZN(G63) );
XNOR2_X1 U812 ( .A(n1116), .B(n1117), .ZN(n1115) );
AND2_X1 U813 ( .A1(G478), .A2(n1118), .ZN(n1116) );
NOR2_X1 U814 ( .A1(n1109), .A2(n1119), .ZN(G60) );
XNOR2_X1 U815 ( .A(n1120), .B(n1121), .ZN(n1119) );
AND2_X1 U816 ( .A1(G475), .A2(n1118), .ZN(n1121) );
XNOR2_X1 U817 ( .A(G104), .B(n1122), .ZN(G6) );
NAND4_X1 U818 ( .A1(KEYINPUT12), .A2(n1123), .A3(n1124), .A4(n1040), .ZN(n1122) );
NOR2_X1 U819 ( .A1(n1125), .A2(n1017), .ZN(n1124) );
XNOR2_X1 U820 ( .A(n1033), .B(KEYINPUT60), .ZN(n1125) );
NOR2_X1 U821 ( .A1(n1109), .A2(n1126), .ZN(G57) );
XOR2_X1 U822 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U823 ( .A(n1129), .B(n1130), .Z(n1128) );
XNOR2_X1 U824 ( .A(n1131), .B(n1132), .ZN(n1127) );
NOR3_X1 U825 ( .A1(n1114), .A2(KEYINPUT13), .A3(n1133), .ZN(n1132) );
NOR2_X1 U826 ( .A1(KEYINPUT54), .A2(n1134), .ZN(n1131) );
NOR2_X1 U827 ( .A1(n1109), .A2(n1135), .ZN(G54) );
XOR2_X1 U828 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U829 ( .A(n1078), .B(n1138), .Z(n1137) );
XOR2_X1 U830 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U831 ( .A1(KEYINPUT26), .A2(n1141), .ZN(n1139) );
XOR2_X1 U832 ( .A(n1142), .B(n1143), .Z(n1136) );
XNOR2_X1 U833 ( .A(G140), .B(n1144), .ZN(n1143) );
XNOR2_X1 U834 ( .A(n1145), .B(n1146), .ZN(n1142) );
NAND2_X1 U835 ( .A1(KEYINPUT62), .A2(G110), .ZN(n1146) );
NAND3_X1 U836 ( .A1(n1118), .A2(G469), .A3(KEYINPUT58), .ZN(n1145) );
INV_X1 U837 ( .A(n1114), .ZN(n1118) );
NOR2_X1 U838 ( .A1(n1109), .A2(n1147), .ZN(G51) );
XOR2_X1 U839 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U840 ( .A(n1150), .B(n1151), .ZN(n1149) );
XOR2_X1 U841 ( .A(n1152), .B(n1153), .Z(n1148) );
NOR2_X1 U842 ( .A1(n1154), .A2(n1114), .ZN(n1152) );
NAND2_X1 U843 ( .A1(G902), .A2(n1000), .ZN(n1114) );
NAND3_X1 U844 ( .A1(n1155), .A2(n1104), .A3(n1156), .ZN(n1000) );
INV_X1 U845 ( .A(n1090), .ZN(n1156) );
NAND2_X1 U846 ( .A1(n1157), .A2(n1158), .ZN(n1090) );
NOR4_X1 U847 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1158) );
INV_X1 U848 ( .A(n1163), .ZN(n1161) );
INV_X1 U849 ( .A(n1164), .ZN(n1160) );
NOR4_X1 U850 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1157) );
NOR2_X1 U851 ( .A1(KEYINPUT29), .A2(n1169), .ZN(n1168) );
NOR3_X1 U852 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1167) );
NOR2_X1 U853 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NOR3_X1 U854 ( .A1(n1009), .A2(n996), .A3(n1175), .ZN(n1174) );
AND4_X1 U855 ( .A1(n1024), .A2(n1033), .A3(n1026), .A4(KEYINPUT29), .ZN(n1173) );
INV_X1 U856 ( .A(n1040), .ZN(n1170) );
INV_X1 U857 ( .A(n1176), .ZN(n1166) );
AND3_X1 U858 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1104) );
NAND2_X1 U859 ( .A1(n1019), .A2(n1180), .ZN(n1179) );
NAND2_X1 U860 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND2_X1 U861 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XNOR2_X1 U862 ( .A(KEYINPUT51), .B(n1185), .ZN(n1181) );
NAND3_X1 U863 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1177) );
XNOR2_X1 U864 ( .A(KEYINPUT24), .B(n1009), .ZN(n1187) );
XOR2_X1 U865 ( .A(n1103), .B(KEYINPUT6), .Z(n1155) );
OR3_X1 U866 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1103) );
AND2_X1 U867 ( .A1(n1019), .A2(n1192), .ZN(n1191) );
NAND2_X1 U868 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NAND2_X1 U869 ( .A1(n1040), .A2(n1195), .ZN(n1194) );
XOR2_X1 U870 ( .A(n997), .B(KEYINPUT15), .Z(n1193) );
NAND2_X1 U871 ( .A1(n1041), .A2(n1195), .ZN(n997) );
AND3_X1 U872 ( .A1(n1027), .A2(n1184), .A3(n1033), .ZN(n1195) );
NOR2_X1 U873 ( .A1(n1060), .A2(G952), .ZN(n1109) );
XOR2_X1 U874 ( .A(n1162), .B(n1196), .Z(G48) );
NOR2_X1 U875 ( .A1(KEYINPUT4), .A2(n1197), .ZN(n1196) );
INV_X1 U876 ( .A(G146), .ZN(n1197) );
AND2_X1 U877 ( .A1(n1040), .A2(n1198), .ZN(n1162) );
XNOR2_X1 U878 ( .A(G143), .B(n1176), .ZN(G45) );
NAND4_X1 U879 ( .A1(n1019), .A2(n1033), .A3(n1026), .A4(n1199), .ZN(n1176) );
NOR3_X1 U880 ( .A1(n1051), .A2(n1200), .A3(n1171), .ZN(n1199) );
XOR2_X1 U881 ( .A(G140), .B(n1165), .Z(G42) );
AND3_X1 U882 ( .A1(n1040), .A2(n1201), .A3(n1025), .ZN(n1165) );
XNOR2_X1 U883 ( .A(G137), .B(n1163), .ZN(G39) );
NAND3_X1 U884 ( .A1(n1201), .A2(n1186), .A3(n1202), .ZN(n1163) );
XNOR2_X1 U885 ( .A(G134), .B(n1164), .ZN(G36) );
NAND3_X1 U886 ( .A1(n1201), .A2(n1041), .A3(n1026), .ZN(n1164) );
XOR2_X1 U887 ( .A(n1169), .B(n1203), .Z(G33) );
XNOR2_X1 U888 ( .A(KEYINPUT45), .B(n1204), .ZN(n1203) );
NAND3_X1 U889 ( .A1(n1026), .A2(n1201), .A3(n1040), .ZN(n1169) );
NOR3_X1 U890 ( .A1(n1205), .A2(n1171), .A3(n1024), .ZN(n1201) );
OR2_X1 U891 ( .A1(n1022), .A2(n1206), .ZN(n1024) );
AND2_X1 U892 ( .A1(G214), .A2(n1021), .ZN(n1206) );
INV_X1 U893 ( .A(n1207), .ZN(n1171) );
XNOR2_X1 U894 ( .A(n1208), .B(n1159), .ZN(G30) );
AND2_X1 U895 ( .A1(n1198), .A2(n1041), .ZN(n1159) );
AND4_X1 U896 ( .A1(n1186), .A2(n1019), .A3(n1033), .A4(n1207), .ZN(n1198) );
XOR2_X1 U897 ( .A(G101), .B(n1189), .Z(G3) );
AND3_X1 U898 ( .A1(n1026), .A2(n1033), .A3(n1188), .ZN(n1189) );
INV_X1 U899 ( .A(n1209), .ZN(n1188) );
XNOR2_X1 U900 ( .A(n1210), .B(n1211), .ZN(G27) );
NOR3_X1 U901 ( .A1(n1212), .A2(n1009), .A3(n1213), .ZN(n1211) );
XNOR2_X1 U902 ( .A(KEYINPUT8), .B(n1207), .ZN(n1213) );
NAND2_X1 U903 ( .A1(n1214), .A2(n1215), .ZN(n1207) );
NAND3_X1 U904 ( .A1(G902), .A2(n1042), .A3(n1066), .ZN(n1214) );
NOR2_X1 U905 ( .A1(n1060), .A2(G900), .ZN(n1066) );
NAND3_X1 U906 ( .A1(n1040), .A2(n1019), .A3(n1025), .ZN(n1212) );
INV_X1 U907 ( .A(n1175), .ZN(n1025) );
XNOR2_X1 U908 ( .A(G122), .B(n1216), .ZN(G24) );
NAND3_X1 U909 ( .A1(n1183), .A2(n1019), .A3(n1217), .ZN(n1216) );
XOR2_X1 U910 ( .A(n1184), .B(KEYINPUT40), .Z(n1217) );
NOR4_X1 U911 ( .A1(n1009), .A2(n1017), .A3(n1051), .A4(n1200), .ZN(n1183) );
INV_X1 U912 ( .A(n1027), .ZN(n1017) );
NOR2_X1 U913 ( .A1(n1048), .A2(n1218), .ZN(n1027) );
XOR2_X1 U914 ( .A(G119), .B(n1219), .Z(G21) );
NOR3_X1 U915 ( .A1(n1220), .A2(n1009), .A3(n1209), .ZN(n1219) );
XOR2_X1 U916 ( .A(KEYINPUT35), .B(n1186), .Z(n1220) );
AND2_X1 U917 ( .A1(n1218), .A2(n1048), .ZN(n1186) );
XNOR2_X1 U918 ( .A(n1221), .B(n1222), .ZN(G18) );
NOR2_X1 U919 ( .A1(n996), .A2(n1185), .ZN(n1222) );
NAND4_X1 U920 ( .A1(n1223), .A2(n1026), .A3(n1041), .A4(n1184), .ZN(n1185) );
INV_X1 U921 ( .A(n1028), .ZN(n1041) );
NAND2_X1 U922 ( .A1(n1224), .A2(n1225), .ZN(n1028) );
XOR2_X1 U923 ( .A(n1051), .B(KEYINPUT14), .Z(n1224) );
XOR2_X1 U924 ( .A(n1178), .B(n1226), .Z(G15) );
XNOR2_X1 U925 ( .A(G113), .B(KEYINPUT33), .ZN(n1226) );
NAND4_X1 U926 ( .A1(n1123), .A2(n1223), .A3(n1040), .A4(n1026), .ZN(n1178) );
NOR2_X1 U927 ( .A1(n1048), .A2(n1050), .ZN(n1026) );
NOR2_X1 U928 ( .A1(n1225), .A2(n1051), .ZN(n1040) );
INV_X1 U929 ( .A(n1200), .ZN(n1225) );
INV_X1 U930 ( .A(n1009), .ZN(n1223) );
NAND2_X1 U931 ( .A1(n1036), .A2(n1227), .ZN(n1009) );
XOR2_X1 U932 ( .A(G110), .B(n1190), .Z(G12) );
NOR3_X1 U933 ( .A1(n1175), .A2(n1205), .A3(n1209), .ZN(n1190) );
NAND2_X1 U934 ( .A1(n1123), .A2(n1202), .ZN(n1209) );
INV_X1 U935 ( .A(n1013), .ZN(n1202) );
NAND2_X1 U936 ( .A1(n1200), .A2(n1051), .ZN(n1013) );
XOR2_X1 U937 ( .A(n1228), .B(G475), .Z(n1051) );
NAND2_X1 U938 ( .A1(n1120), .A2(n1229), .ZN(n1228) );
XNOR2_X1 U939 ( .A(n1230), .B(n1231), .ZN(n1120) );
XNOR2_X1 U940 ( .A(n1232), .B(n1233), .ZN(n1231) );
XOR2_X1 U941 ( .A(n1234), .B(n1235), .Z(n1233) );
NOR2_X1 U942 ( .A1(KEYINPUT39), .A2(n1236), .ZN(n1235) );
XNOR2_X1 U943 ( .A(G146), .B(n1073), .ZN(n1236) );
XOR2_X1 U944 ( .A(G125), .B(G140), .Z(n1073) );
NAND3_X1 U945 ( .A1(n1237), .A2(n1060), .A3(G214), .ZN(n1234) );
XOR2_X1 U946 ( .A(n1238), .B(n1239), .Z(n1230) );
XNOR2_X1 U947 ( .A(KEYINPUT50), .B(n1204), .ZN(n1239) );
XNOR2_X1 U948 ( .A(G113), .B(G104), .ZN(n1238) );
NOR2_X1 U949 ( .A1(n1240), .A2(n1052), .ZN(n1200) );
NOR3_X1 U950 ( .A1(G478), .A2(G902), .A3(n1241), .ZN(n1052) );
AND2_X1 U951 ( .A1(n1242), .A2(n1053), .ZN(n1240) );
NAND2_X1 U952 ( .A1(n1117), .A2(n1229), .ZN(n1053) );
INV_X1 U953 ( .A(n1241), .ZN(n1117) );
XNOR2_X1 U954 ( .A(n1243), .B(n1244), .ZN(n1241) );
AND3_X1 U955 ( .A1(G234), .A2(n1060), .A3(G217), .ZN(n1244) );
NAND2_X1 U956 ( .A1(n1245), .A2(KEYINPUT41), .ZN(n1243) );
XOR2_X1 U957 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U958 ( .A(n1248), .B(n1232), .Z(n1247) );
XNOR2_X1 U959 ( .A(G122), .B(n1249), .ZN(n1232) );
XNOR2_X1 U960 ( .A(G128), .B(n1250), .ZN(n1246) );
XNOR2_X1 U961 ( .A(KEYINPUT18), .B(n1089), .ZN(n1250) );
XNOR2_X1 U962 ( .A(G478), .B(KEYINPUT43), .ZN(n1242) );
AND2_X1 U963 ( .A1(n1019), .A2(n1184), .ZN(n1123) );
NAND2_X1 U964 ( .A1(n1215), .A2(n1251), .ZN(n1184) );
NAND3_X1 U965 ( .A1(G902), .A2(n1042), .A3(n1106), .ZN(n1251) );
NOR2_X1 U966 ( .A1(G898), .A2(n1060), .ZN(n1106) );
NAND3_X1 U967 ( .A1(n1252), .A2(n1042), .A3(G952), .ZN(n1215) );
NAND2_X1 U968 ( .A1(G237), .A2(G234), .ZN(n1042) );
XOR2_X1 U969 ( .A(KEYINPUT48), .B(n1001), .Z(n1252) );
XNOR2_X1 U970 ( .A(n1060), .B(KEYINPUT25), .ZN(n1001) );
INV_X1 U971 ( .A(n996), .ZN(n1019) );
NAND2_X1 U972 ( .A1(n1022), .A2(n1253), .ZN(n996) );
NAND2_X1 U973 ( .A1(G214), .A2(n1021), .ZN(n1253) );
XOR2_X1 U974 ( .A(n1254), .B(n1154), .Z(n1022) );
NAND2_X1 U975 ( .A1(G210), .A2(n1021), .ZN(n1154) );
NAND2_X1 U976 ( .A1(n1255), .A2(n1237), .ZN(n1021) );
NAND3_X1 U977 ( .A1(n1256), .A2(n1229), .A3(n1257), .ZN(n1254) );
XOR2_X1 U978 ( .A(n1258), .B(KEYINPUT46), .Z(n1257) );
NAND2_X1 U979 ( .A1(n1151), .A2(n1259), .ZN(n1258) );
OR2_X1 U980 ( .A1(n1259), .A2(n1151), .ZN(n1256) );
XNOR2_X1 U981 ( .A(n1107), .B(n1260), .ZN(n1151) );
XOR2_X1 U982 ( .A(KEYINPUT59), .B(n1261), .Z(n1260) );
NOR2_X1 U983 ( .A1(KEYINPUT11), .A2(n1108), .ZN(n1261) );
XOR2_X1 U984 ( .A(n1262), .B(G110), .Z(n1108) );
NAND2_X1 U985 ( .A1(KEYINPUT2), .A2(n1263), .ZN(n1262) );
INV_X1 U986 ( .A(G122), .ZN(n1263) );
XOR2_X1 U987 ( .A(n1130), .B(n1264), .Z(n1107) );
XOR2_X1 U988 ( .A(G104), .B(n1248), .Z(n1264) );
XNOR2_X1 U989 ( .A(n994), .B(G116), .ZN(n1248) );
XNOR2_X1 U990 ( .A(G101), .B(n1265), .ZN(n1130) );
XNOR2_X1 U991 ( .A(n1266), .B(n1153), .ZN(n1259) );
XNOR2_X1 U992 ( .A(n1210), .B(n1267), .ZN(n1153) );
NOR2_X1 U993 ( .A1(n1098), .A2(G953), .ZN(n1267) );
INV_X1 U994 ( .A(G224), .ZN(n1098) );
INV_X1 U995 ( .A(G125), .ZN(n1210) );
NAND2_X1 U996 ( .A1(KEYINPUT34), .A2(n1150), .ZN(n1266) );
INV_X1 U997 ( .A(n1033), .ZN(n1205) );
NOR2_X1 U998 ( .A1(n1036), .A2(n1037), .ZN(n1033) );
INV_X1 U999 ( .A(n1227), .ZN(n1037) );
NAND2_X1 U1000 ( .A1(G221), .A2(n1268), .ZN(n1227) );
XNOR2_X1 U1001 ( .A(n1055), .B(G469), .ZN(n1036) );
AND2_X1 U1002 ( .A1(n1269), .A2(n1229), .ZN(n1055) );
XOR2_X1 U1003 ( .A(n1270), .B(n1271), .Z(n1269) );
XNOR2_X1 U1004 ( .A(n1272), .B(n1144), .ZN(n1271) );
NAND2_X1 U1005 ( .A1(n1273), .A2(n1060), .ZN(n1144) );
XOR2_X1 U1006 ( .A(KEYINPUT7), .B(G227), .Z(n1273) );
NAND2_X1 U1007 ( .A1(KEYINPUT10), .A2(n1274), .ZN(n1272) );
XOR2_X1 U1008 ( .A(G140), .B(G110), .Z(n1274) );
XNOR2_X1 U1009 ( .A(KEYINPUT27), .B(n1275), .ZN(n1270) );
NOR2_X1 U1010 ( .A1(KEYINPUT23), .A2(n1276), .ZN(n1275) );
XOR2_X1 U1011 ( .A(n1277), .B(n1140), .Z(n1276) );
XOR2_X1 U1012 ( .A(G101), .B(n1278), .Z(n1140) );
NOR2_X1 U1013 ( .A1(KEYINPUT52), .A2(n1279), .ZN(n1278) );
XNOR2_X1 U1014 ( .A(G104), .B(n1280), .ZN(n1279) );
NOR2_X1 U1015 ( .A1(KEYINPUT16), .A2(n994), .ZN(n1280) );
INV_X1 U1016 ( .A(G107), .ZN(n994) );
XNOR2_X1 U1017 ( .A(n1141), .B(n1281), .ZN(n1277) );
NOR2_X1 U1018 ( .A1(KEYINPUT30), .A2(n1078), .ZN(n1281) );
XNOR2_X1 U1019 ( .A(G128), .B(n1282), .ZN(n1078) );
NOR2_X1 U1020 ( .A1(KEYINPUT61), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U1021 ( .A(G146), .B(n1284), .ZN(n1283) );
NAND2_X1 U1022 ( .A1(KEYINPUT20), .A2(n1249), .ZN(n1284) );
INV_X1 U1023 ( .A(G143), .ZN(n1249) );
NAND2_X1 U1024 ( .A1(n1050), .A2(n1048), .ZN(n1175) );
XOR2_X1 U1025 ( .A(n1285), .B(n1113), .Z(n1048) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1268), .ZN(n1113) );
NAND2_X1 U1027 ( .A1(G234), .A2(n1255), .ZN(n1268) );
XNOR2_X1 U1028 ( .A(G902), .B(KEYINPUT19), .ZN(n1255) );
NAND2_X1 U1029 ( .A1(n1111), .A2(n1229), .ZN(n1285) );
XNOR2_X1 U1030 ( .A(n1286), .B(n1287), .ZN(n1111) );
XOR2_X1 U1031 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U1032 ( .A(G110), .B(n1290), .Z(n1289) );
AND3_X1 U1033 ( .A1(G221), .A2(n1060), .A3(G234), .ZN(n1290) );
INV_X1 U1034 ( .A(G953), .ZN(n1060) );
XOR2_X1 U1035 ( .A(KEYINPUT28), .B(G119), .Z(n1288) );
XOR2_X1 U1036 ( .A(n1291), .B(n1292), .Z(n1286) );
XNOR2_X1 U1037 ( .A(n1293), .B(n1294), .ZN(n1291) );
NAND2_X1 U1038 ( .A1(KEYINPUT5), .A2(n1295), .ZN(n1294) );
NAND2_X1 U1039 ( .A1(n1296), .A2(KEYINPUT44), .ZN(n1293) );
XOR2_X1 U1040 ( .A(n1297), .B(G140), .Z(n1296) );
NAND2_X1 U1041 ( .A1(KEYINPUT56), .A2(G125), .ZN(n1297) );
INV_X1 U1042 ( .A(n1218), .ZN(n1050) );
XNOR2_X1 U1043 ( .A(n1298), .B(n1299), .ZN(n1218) );
XNOR2_X1 U1044 ( .A(KEYINPUT37), .B(n1133), .ZN(n1299) );
INV_X1 U1045 ( .A(G472), .ZN(n1133) );
NAND2_X1 U1046 ( .A1(n1300), .A2(n1229), .ZN(n1298) );
INV_X1 U1047 ( .A(G902), .ZN(n1229) );
XOR2_X1 U1048 ( .A(n1265), .B(n1301), .Z(n1300) );
XNOR2_X1 U1049 ( .A(n1129), .B(n1302), .ZN(n1301) );
NOR2_X1 U1050 ( .A1(KEYINPUT63), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1051 ( .A(G101), .B(n1134), .Z(n1303) );
NAND3_X1 U1052 ( .A1(G210), .A2(n1237), .A3(n1304), .ZN(n1134) );
XNOR2_X1 U1053 ( .A(G953), .B(KEYINPUT53), .ZN(n1304) );
INV_X1 U1054 ( .A(G237), .ZN(n1237) );
XOR2_X1 U1055 ( .A(n1150), .B(n1305), .Z(n1129) );
XNOR2_X1 U1056 ( .A(n1141), .B(n1306), .ZN(n1305) );
NAND2_X1 U1057 ( .A1(KEYINPUT36), .A2(n1221), .ZN(n1306) );
INV_X1 U1058 ( .A(G116), .ZN(n1221) );
AND3_X1 U1059 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1141) );
NAND2_X1 U1060 ( .A1(G137), .A2(n1310), .ZN(n1309) );
XNOR2_X1 U1061 ( .A(n1089), .B(G131), .ZN(n1310) );
NAND3_X1 U1062 ( .A1(n1089), .A2(n1295), .A3(n1204), .ZN(n1308) );
INV_X1 U1063 ( .A(G131), .ZN(n1204) );
INV_X1 U1064 ( .A(G137), .ZN(n1295) );
NAND2_X1 U1065 ( .A1(n1087), .A2(G131), .ZN(n1307) );
NOR2_X1 U1066 ( .A1(n1089), .A2(G137), .ZN(n1087) );
INV_X1 U1067 ( .A(G134), .ZN(n1089) );
XNOR2_X1 U1068 ( .A(n1311), .B(n1292), .ZN(n1150) );
XNOR2_X1 U1069 ( .A(n1208), .B(G146), .ZN(n1292) );
INV_X1 U1070 ( .A(G128), .ZN(n1208) );
XNOR2_X1 U1071 ( .A(G143), .B(KEYINPUT21), .ZN(n1311) );
XNOR2_X1 U1072 ( .A(G113), .B(G119), .ZN(n1265) );
endmodule


