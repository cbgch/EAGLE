//Key = 0110010101000101011001000111000001000110111111000011111100100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351;

XNOR2_X1 U749 ( .A(G107), .B(n1036), .ZN(G9) );
NAND2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
XOR2_X1 U751 ( .A(n1039), .B(KEYINPUT38), .Z(n1037) );
NOR2_X1 U752 ( .A1(n1040), .A2(n1041), .ZN(G75) );
NOR4_X1 U753 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1041) );
NOR2_X1 U754 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR3_X1 U755 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1044) );
NOR2_X1 U756 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U757 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR3_X1 U758 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1053) );
NOR3_X1 U759 ( .A1(n1058), .A2(KEYINPUT41), .A3(n1059), .ZN(n1057) );
INV_X1 U760 ( .A(n1060), .ZN(n1059) );
NOR2_X1 U761 ( .A1(n1061), .A2(n1062), .ZN(n1056) );
NOR2_X1 U762 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
AND2_X1 U763 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
AND2_X1 U764 ( .A1(n1060), .A2(KEYINPUT41), .ZN(n1063) );
NOR2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1055) );
NOR2_X1 U766 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR3_X1 U767 ( .A1(n1062), .A2(n1071), .A3(n1068), .ZN(n1051) );
NOR2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NAND3_X1 U770 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1042) );
NAND3_X1 U771 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
XOR2_X1 U772 ( .A(n1047), .B(KEYINPUT58), .Z(n1081) );
OR4_X1 U773 ( .A1(n1048), .A2(n1054), .A3(n1062), .A4(n1068), .ZN(n1047) );
NOR3_X1 U774 ( .A1(n1082), .A2(G953), .A3(G952), .ZN(n1040) );
INV_X1 U775 ( .A(n1076), .ZN(n1082) );
NAND4_X1 U776 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1076) );
NOR3_X1 U777 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
XOR2_X1 U778 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U779 ( .A1(n1092), .A2(KEYINPUT10), .ZN(n1091) );
INV_X1 U780 ( .A(n1093), .ZN(n1092) );
NAND3_X1 U781 ( .A1(n1075), .A2(n1094), .A3(n1095), .ZN(n1087) );
NOR3_X1 U782 ( .A1(n1065), .A2(n1096), .A3(n1097), .ZN(n1085) );
AND2_X1 U783 ( .A1(G469), .A2(n1098), .ZN(n1097) );
NOR2_X1 U784 ( .A1(G469), .A2(n1099), .ZN(n1096) );
NOR2_X1 U785 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U786 ( .A1(KEYINPUT59), .A2(n1098), .ZN(n1101) );
NOR2_X1 U787 ( .A1(n1102), .A2(KEYINPUT63), .ZN(n1098) );
INV_X1 U788 ( .A(n1103), .ZN(n1102) );
AND2_X1 U789 ( .A1(n1103), .A2(KEYINPUT59), .ZN(n1100) );
XNOR2_X1 U790 ( .A(n1104), .B(n1105), .ZN(n1084) );
XNOR2_X1 U791 ( .A(G475), .B(KEYINPUT18), .ZN(n1105) );
XNOR2_X1 U792 ( .A(n1106), .B(n1107), .ZN(n1083) );
XNOR2_X1 U793 ( .A(G472), .B(KEYINPUT44), .ZN(n1107) );
XOR2_X1 U794 ( .A(n1108), .B(n1109), .Z(G72) );
NOR2_X1 U795 ( .A1(n1110), .A2(n1077), .ZN(n1109) );
NOR2_X1 U796 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1108) );
NAND3_X1 U798 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
NAND2_X1 U799 ( .A1(G953), .A2(n1112), .ZN(n1116) );
OR2_X1 U800 ( .A1(n1115), .A2(n1117), .ZN(n1113) );
NAND2_X1 U801 ( .A1(n1077), .A2(n1118), .ZN(n1117) );
NAND3_X1 U802 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1118) );
XOR2_X1 U803 ( .A(n1122), .B(KEYINPUT25), .Z(n1121) );
INV_X1 U804 ( .A(n1123), .ZN(n1119) );
XNOR2_X1 U805 ( .A(n1124), .B(n1125), .ZN(n1115) );
NOR2_X1 U806 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U807 ( .A(n1128), .B(KEYINPUT1), .Z(n1127) );
NAND2_X1 U808 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(n1126) );
XOR2_X1 U810 ( .A(n1131), .B(G134), .Z(n1129) );
XOR2_X1 U811 ( .A(n1132), .B(n1133), .Z(G69) );
XOR2_X1 U812 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U813 ( .A1(n1136), .A2(n1077), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XNOR2_X1 U815 ( .A(G224), .B(KEYINPUT32), .ZN(n1137) );
NAND2_X1 U816 ( .A1(n1139), .A2(n1140), .ZN(n1134) );
XNOR2_X1 U817 ( .A(n1141), .B(n1142), .ZN(n1140) );
XNOR2_X1 U818 ( .A(n1143), .B(n1144), .ZN(n1141) );
XOR2_X1 U819 ( .A(n1145), .B(KEYINPUT56), .Z(n1139) );
NAND2_X1 U820 ( .A1(G953), .A2(n1138), .ZN(n1145) );
NAND2_X1 U821 ( .A1(n1077), .A2(n1146), .ZN(n1132) );
NOR2_X1 U822 ( .A1(n1147), .A2(n1148), .ZN(G66) );
XOR2_X1 U823 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U824 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
NOR2_X1 U825 ( .A1(n1153), .A2(n1154), .ZN(G63) );
XNOR2_X1 U826 ( .A(n1155), .B(n1156), .ZN(n1154) );
NOR2_X1 U827 ( .A1(n1157), .A2(n1152), .ZN(n1155) );
XNOR2_X1 U828 ( .A(n1147), .B(KEYINPUT33), .ZN(n1153) );
NOR2_X1 U829 ( .A1(n1147), .A2(n1158), .ZN(G60) );
NOR3_X1 U830 ( .A1(n1104), .A2(n1159), .A3(n1160), .ZN(n1158) );
AND3_X1 U831 ( .A1(n1161), .A2(G475), .A3(n1162), .ZN(n1160) );
NOR2_X1 U832 ( .A1(n1163), .A2(n1161), .ZN(n1159) );
AND2_X1 U833 ( .A1(n1043), .A2(G475), .ZN(n1163) );
XNOR2_X1 U834 ( .A(G104), .B(n1164), .ZN(G6) );
NOR2_X1 U835 ( .A1(n1147), .A2(n1165), .ZN(G57) );
XOR2_X1 U836 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U837 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U838 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U839 ( .A1(n1172), .A2(n1173), .ZN(n1168) );
AND2_X1 U840 ( .A1(KEYINPUT31), .A2(n1174), .ZN(n1173) );
NOR2_X1 U841 ( .A1(KEYINPUT19), .A2(n1174), .ZN(n1172) );
XOR2_X1 U842 ( .A(n1175), .B(n1176), .Z(n1166) );
XOR2_X1 U843 ( .A(n1177), .B(KEYINPUT39), .Z(n1176) );
NAND2_X1 U844 ( .A1(n1162), .A2(G472), .ZN(n1177) );
NOR2_X1 U845 ( .A1(n1178), .A2(n1179), .ZN(G54) );
XOR2_X1 U846 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U847 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U848 ( .A(n1184), .B(n1185), .Z(n1180) );
AND2_X1 U849 ( .A1(G469), .A2(n1162), .ZN(n1185) );
INV_X1 U850 ( .A(n1152), .ZN(n1162) );
NAND2_X1 U851 ( .A1(KEYINPUT9), .A2(n1130), .ZN(n1184) );
INV_X1 U852 ( .A(n1186), .ZN(n1130) );
XNOR2_X1 U853 ( .A(n1147), .B(KEYINPUT13), .ZN(n1178) );
NOR2_X1 U854 ( .A1(n1147), .A2(n1187), .ZN(G51) );
XOR2_X1 U855 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U856 ( .A(n1190), .B(n1191), .Z(n1189) );
XOR2_X1 U857 ( .A(n1192), .B(n1193), .Z(n1188) );
NOR2_X1 U858 ( .A1(n1093), .A2(n1152), .ZN(n1193) );
NAND2_X1 U859 ( .A1(G902), .A2(n1043), .ZN(n1152) );
OR4_X1 U860 ( .A1(n1123), .A2(n1122), .A3(n1146), .A4(n1194), .ZN(n1043) );
INV_X1 U861 ( .A(n1120), .ZN(n1194) );
NAND4_X1 U862 ( .A1(n1195), .A2(n1164), .A3(n1196), .A4(n1197), .ZN(n1146) );
AND4_X1 U863 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
NAND2_X1 U864 ( .A1(n1202), .A2(n1203), .ZN(n1196) );
INV_X1 U865 ( .A(KEYINPUT0), .ZN(n1203) );
NAND4_X1 U866 ( .A1(n1204), .A2(n1070), .A3(n1073), .A4(n1205), .ZN(n1164) );
NAND2_X1 U867 ( .A1(n1038), .A2(n1206), .ZN(n1195) );
NAND3_X1 U868 ( .A1(n1207), .A2(n1039), .A3(n1208), .ZN(n1206) );
XNOR2_X1 U869 ( .A(KEYINPUT54), .B(n1209), .ZN(n1208) );
NAND4_X1 U870 ( .A1(n1073), .A2(n1069), .A3(n1205), .A4(n1210), .ZN(n1039) );
NAND3_X1 U871 ( .A1(n1211), .A2(n1212), .A3(KEYINPUT0), .ZN(n1207) );
NAND4_X1 U872 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1122) );
NAND4_X1 U873 ( .A1(n1217), .A2(n1218), .A3(n1069), .A4(n1219), .ZN(n1213) );
NAND3_X1 U874 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1123) );
NOR2_X1 U875 ( .A1(n1077), .A2(G952), .ZN(n1147) );
XOR2_X1 U876 ( .A(n1223), .B(n1222), .Z(G48) );
NAND3_X1 U877 ( .A1(n1224), .A2(n1038), .A3(n1070), .ZN(n1222) );
XNOR2_X1 U878 ( .A(G143), .B(n1220), .ZN(G45) );
NAND3_X1 U879 ( .A1(n1225), .A2(n1217), .A3(n1226), .ZN(n1220) );
AND3_X1 U880 ( .A1(n1038), .A2(n1227), .A3(n1219), .ZN(n1226) );
XOR2_X1 U881 ( .A(n1228), .B(G140), .Z(G42) );
NAND2_X1 U882 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
OR2_X1 U883 ( .A1(n1120), .A2(KEYINPUT36), .ZN(n1230) );
NAND3_X1 U884 ( .A1(n1218), .A2(n1073), .A3(n1231), .ZN(n1120) );
NAND4_X1 U885 ( .A1(n1073), .A2(n1050), .A3(n1231), .A4(KEYINPUT36), .ZN(n1229) );
XNOR2_X1 U886 ( .A(G137), .B(n1221), .ZN(G39) );
NAND3_X1 U887 ( .A1(n1224), .A2(n1218), .A3(n1058), .ZN(n1221) );
XOR2_X1 U888 ( .A(n1232), .B(n1233), .Z(G36) );
XOR2_X1 U889 ( .A(KEYINPUT52), .B(G134), .Z(n1233) );
NAND4_X1 U890 ( .A1(n1217), .A2(n1218), .A3(n1069), .A4(n1234), .ZN(n1232) );
XNOR2_X1 U891 ( .A(KEYINPUT7), .B(n1219), .ZN(n1234) );
XNOR2_X1 U892 ( .A(n1215), .B(n1235), .ZN(G33) );
NOR2_X1 U893 ( .A1(KEYINPUT34), .A2(n1236), .ZN(n1235) );
INV_X1 U894 ( .A(G131), .ZN(n1236) );
NAND4_X1 U895 ( .A1(n1070), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1215) );
INV_X1 U896 ( .A(n1050), .ZN(n1218) );
NAND2_X1 U897 ( .A1(n1237), .A2(n1095), .ZN(n1050) );
XNOR2_X1 U898 ( .A(KEYINPUT45), .B(n1079), .ZN(n1237) );
XNOR2_X1 U899 ( .A(G128), .B(n1216), .ZN(G30) );
NAND3_X1 U900 ( .A1(n1038), .A2(n1069), .A3(n1224), .ZN(n1216) );
AND4_X1 U901 ( .A1(n1238), .A2(n1073), .A3(n1065), .A4(n1219), .ZN(n1224) );
XNOR2_X1 U902 ( .A(G101), .B(n1201), .ZN(G3) );
NAND2_X1 U903 ( .A1(n1239), .A2(n1217), .ZN(n1201) );
AND2_X1 U904 ( .A1(n1060), .A2(n1073), .ZN(n1217) );
NAND2_X1 U905 ( .A1(n1240), .A2(n1241), .ZN(G27) );
NAND2_X1 U906 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND2_X1 U907 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
OR2_X1 U908 ( .A1(n1246), .A2(KEYINPUT42), .ZN(n1245) );
INV_X1 U909 ( .A(n1214), .ZN(n1242) );
NAND3_X1 U910 ( .A1(n1247), .A2(n1248), .A3(KEYINPUT42), .ZN(n1240) );
NAND2_X1 U911 ( .A1(KEYINPUT27), .A2(n1249), .ZN(n1248) );
NAND2_X1 U912 ( .A1(n1244), .A2(n1214), .ZN(n1249) );
NAND3_X1 U913 ( .A1(n1231), .A2(n1038), .A3(n1250), .ZN(n1214) );
AND4_X1 U914 ( .A1(n1070), .A2(n1066), .A3(n1065), .A4(n1219), .ZN(n1231) );
NAND2_X1 U915 ( .A1(n1048), .A2(n1251), .ZN(n1219) );
NAND4_X1 U916 ( .A1(G953), .A2(G902), .A3(n1252), .A4(n1112), .ZN(n1251) );
INV_X1 U917 ( .A(G900), .ZN(n1112) );
NAND2_X1 U918 ( .A1(n1244), .A2(n1246), .ZN(n1247) );
INV_X1 U919 ( .A(KEYINPUT27), .ZN(n1246) );
XOR2_X1 U920 ( .A(G125), .B(KEYINPUT22), .Z(n1244) );
XOR2_X1 U921 ( .A(G122), .B(n1202), .Z(G24) );
AND2_X1 U922 ( .A1(n1211), .A2(n1204), .ZN(n1202) );
NOR4_X1 U923 ( .A1(n1253), .A2(n1054), .A3(n1068), .A4(n1254), .ZN(n1211) );
INV_X1 U924 ( .A(n1205), .ZN(n1068) );
NOR2_X1 U925 ( .A1(n1065), .A2(n1238), .ZN(n1205) );
XOR2_X1 U926 ( .A(n1255), .B(n1200), .Z(G21) );
NAND4_X1 U927 ( .A1(n1239), .A2(n1250), .A3(n1238), .A4(n1065), .ZN(n1200) );
XOR2_X1 U928 ( .A(G116), .B(n1256), .Z(G18) );
NOR2_X1 U929 ( .A1(n1046), .A2(n1209), .ZN(n1256) );
NAND4_X1 U930 ( .A1(n1250), .A2(n1060), .A3(n1069), .A4(n1210), .ZN(n1209) );
NOR2_X1 U931 ( .A1(n1225), .A2(n1254), .ZN(n1069) );
XOR2_X1 U932 ( .A(n1257), .B(n1199), .Z(G15) );
NAND4_X1 U933 ( .A1(n1204), .A2(n1250), .A3(n1070), .A4(n1060), .ZN(n1199) );
NOR2_X1 U934 ( .A1(n1066), .A2(n1065), .ZN(n1060) );
NOR2_X1 U935 ( .A1(n1253), .A2(n1227), .ZN(n1070) );
INV_X1 U936 ( .A(n1054), .ZN(n1250) );
NAND2_X1 U937 ( .A1(n1258), .A2(n1075), .ZN(n1054) );
INV_X1 U938 ( .A(n1074), .ZN(n1258) );
XNOR2_X1 U939 ( .A(G110), .B(n1198), .ZN(G12) );
NAND4_X1 U940 ( .A1(n1239), .A2(n1073), .A3(n1066), .A4(n1065), .ZN(n1198) );
XNOR2_X1 U941 ( .A(n1259), .B(n1260), .ZN(n1065) );
NOR2_X1 U942 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U943 ( .A(KEYINPUT50), .B(G217), .Z(n1262) );
INV_X1 U944 ( .A(n1263), .ZN(n1261) );
OR2_X1 U945 ( .A1(n1150), .A2(G902), .ZN(n1259) );
XNOR2_X1 U946 ( .A(n1264), .B(n1265), .ZN(n1150) );
XOR2_X1 U947 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U948 ( .A(n1268), .B(n1269), .Z(n1267) );
NOR2_X1 U949 ( .A1(KEYINPUT16), .A2(n1270), .ZN(n1269) );
XOR2_X1 U950 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U951 ( .A(n1255), .B(G128), .Z(n1271) );
NAND3_X1 U952 ( .A1(G234), .A2(n1077), .A3(G221), .ZN(n1268) );
XNOR2_X1 U953 ( .A(G137), .B(n1273), .ZN(n1264) );
XOR2_X1 U954 ( .A(KEYINPUT60), .B(G146), .Z(n1273) );
INV_X1 U955 ( .A(n1238), .ZN(n1066) );
XNOR2_X1 U956 ( .A(G472), .B(n1274), .ZN(n1238) );
NOR2_X1 U957 ( .A1(n1106), .A2(KEYINPUT57), .ZN(n1274) );
AND2_X1 U958 ( .A1(n1275), .A2(n1276), .ZN(n1106) );
XOR2_X1 U959 ( .A(KEYINPUT12), .B(n1277), .Z(n1275) );
NOR2_X1 U960 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
AND2_X1 U961 ( .A1(n1280), .A2(n1170), .ZN(n1279) );
NOR2_X1 U962 ( .A1(n1280), .A2(n1281), .ZN(n1278) );
XOR2_X1 U963 ( .A(n1170), .B(KEYINPUT23), .Z(n1281) );
XNOR2_X1 U964 ( .A(G101), .B(n1282), .ZN(n1170) );
AND3_X1 U965 ( .A1(G210), .A2(n1077), .A3(n1283), .ZN(n1282) );
XOR2_X1 U966 ( .A(n1284), .B(n1171), .Z(n1280) );
NAND2_X1 U967 ( .A1(n1285), .A2(n1286), .ZN(n1171) );
NAND2_X1 U968 ( .A1(n1287), .A2(G119), .ZN(n1286) );
NAND2_X1 U969 ( .A1(n1288), .A2(n1255), .ZN(n1285) );
INV_X1 U970 ( .A(G119), .ZN(n1255) );
XNOR2_X1 U971 ( .A(n1287), .B(KEYINPUT46), .ZN(n1288) );
XNOR2_X1 U972 ( .A(n1289), .B(G116), .ZN(n1287) );
NAND2_X1 U973 ( .A1(KEYINPUT5), .A2(n1257), .ZN(n1289) );
NAND2_X1 U974 ( .A1(n1290), .A2(n1291), .ZN(n1284) );
NAND2_X1 U975 ( .A1(n1174), .A2(n1292), .ZN(n1291) );
XOR2_X1 U976 ( .A(n1293), .B(KEYINPUT6), .Z(n1290) );
NAND2_X1 U977 ( .A1(n1175), .A2(n1294), .ZN(n1293) );
AND2_X1 U978 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U979 ( .A1(G221), .A2(n1263), .ZN(n1075) );
NAND2_X1 U980 ( .A1(G234), .A2(n1276), .ZN(n1263) );
XNOR2_X1 U981 ( .A(n1103), .B(G469), .ZN(n1074) );
NAND2_X1 U982 ( .A1(n1295), .A2(n1276), .ZN(n1103) );
XOR2_X1 U983 ( .A(n1296), .B(n1297), .Z(n1295) );
INV_X1 U984 ( .A(n1182), .ZN(n1297) );
XOR2_X1 U985 ( .A(n1298), .B(n1299), .Z(n1182) );
XOR2_X1 U986 ( .A(n1294), .B(n1272), .Z(n1299) );
INV_X1 U987 ( .A(n1174), .ZN(n1294) );
XOR2_X1 U988 ( .A(n1131), .B(n1300), .Z(n1174) );
NOR2_X1 U989 ( .A1(G134), .A2(KEYINPUT35), .ZN(n1300) );
XNOR2_X1 U990 ( .A(G137), .B(n1301), .ZN(n1131) );
XNOR2_X1 U991 ( .A(G140), .B(n1302), .ZN(n1298) );
NOR2_X1 U992 ( .A1(G953), .A2(n1111), .ZN(n1302) );
INV_X1 U993 ( .A(G227), .ZN(n1111) );
XNOR2_X1 U994 ( .A(KEYINPUT11), .B(n1303), .ZN(n1296) );
NOR2_X1 U995 ( .A1(KEYINPUT61), .A2(n1304), .ZN(n1303) );
XNOR2_X1 U996 ( .A(n1305), .B(n1183), .ZN(n1304) );
NAND2_X1 U997 ( .A1(KEYINPUT21), .A2(n1186), .ZN(n1305) );
XNOR2_X1 U998 ( .A(n1306), .B(n1307), .ZN(n1186) );
NOR2_X1 U999 ( .A1(G143), .A2(KEYINPUT62), .ZN(n1307) );
AND2_X1 U1000 ( .A1(n1204), .A2(n1058), .ZN(n1239) );
INV_X1 U1001 ( .A(n1062), .ZN(n1058) );
NAND2_X1 U1002 ( .A1(n1254), .A2(n1253), .ZN(n1062) );
INV_X1 U1003 ( .A(n1225), .ZN(n1253) );
XNOR2_X1 U1004 ( .A(n1104), .B(n1308), .ZN(n1225) );
NOR2_X1 U1005 ( .A1(G475), .A2(KEYINPUT48), .ZN(n1308) );
NOR2_X1 U1006 ( .A1(n1161), .A2(G902), .ZN(n1104) );
XNOR2_X1 U1007 ( .A(n1309), .B(KEYINPUT8), .ZN(n1161) );
XOR2_X1 U1008 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1009 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U1010 ( .A(n1301), .B(n1124), .Z(n1313) );
INV_X1 U1011 ( .A(n1266), .ZN(n1124) );
XNOR2_X1 U1012 ( .A(G125), .B(G140), .ZN(n1266) );
XOR2_X1 U1013 ( .A(G131), .B(KEYINPUT29), .Z(n1301) );
XOR2_X1 U1014 ( .A(n1314), .B(n1315), .Z(n1312) );
NAND2_X1 U1015 ( .A1(KEYINPUT2), .A2(n1223), .ZN(n1315) );
INV_X1 U1016 ( .A(G146), .ZN(n1223) );
NAND3_X1 U1017 ( .A1(G214), .A2(n1077), .A3(n1316), .ZN(n1314) );
XOR2_X1 U1018 ( .A(n1283), .B(KEYINPUT3), .Z(n1316) );
XOR2_X1 U1019 ( .A(n1317), .B(n1318), .Z(n1310) );
XOR2_X1 U1020 ( .A(G143), .B(G122), .Z(n1318) );
XOR2_X1 U1021 ( .A(G104), .B(n1257), .Z(n1317) );
INV_X1 U1022 ( .A(n1227), .ZN(n1254) );
NAND2_X1 U1023 ( .A1(n1319), .A2(n1094), .ZN(n1227) );
NAND3_X1 U1024 ( .A1(n1157), .A2(n1276), .A3(n1156), .ZN(n1094) );
INV_X1 U1025 ( .A(G478), .ZN(n1157) );
XNOR2_X1 U1026 ( .A(n1088), .B(KEYINPUT4), .ZN(n1319) );
AND2_X1 U1027 ( .A1(G478), .A2(n1320), .ZN(n1088) );
NAND2_X1 U1028 ( .A1(n1156), .A2(n1276), .ZN(n1320) );
XOR2_X1 U1029 ( .A(n1321), .B(n1322), .Z(n1156) );
XOR2_X1 U1030 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1031 ( .A(G122), .B(G116), .Z(n1324) );
XOR2_X1 U1032 ( .A(KEYINPUT15), .B(G134), .Z(n1323) );
XOR2_X1 U1033 ( .A(n1325), .B(n1326), .Z(n1321) );
NOR4_X1 U1034 ( .A1(KEYINPUT14), .A2(G953), .A3(n1327), .A4(n1151), .ZN(n1326) );
INV_X1 U1035 ( .A(G217), .ZN(n1151) );
INV_X1 U1036 ( .A(G234), .ZN(n1327) );
XNOR2_X1 U1037 ( .A(G107), .B(n1328), .ZN(n1325) );
NOR2_X1 U1038 ( .A1(KEYINPUT30), .A2(n1329), .ZN(n1328) );
XNOR2_X1 U1039 ( .A(G128), .B(G143), .ZN(n1329) );
NOR2_X1 U1040 ( .A1(n1046), .A2(n1212), .ZN(n1204) );
INV_X1 U1041 ( .A(n1210), .ZN(n1212) );
NAND2_X1 U1042 ( .A1(n1048), .A2(n1330), .ZN(n1210) );
NAND4_X1 U1043 ( .A1(G953), .A2(G902), .A3(n1252), .A4(n1138), .ZN(n1330) );
INV_X1 U1044 ( .A(G898), .ZN(n1138) );
NAND3_X1 U1045 ( .A1(n1252), .A2(n1077), .A3(n1331), .ZN(n1048) );
XOR2_X1 U1046 ( .A(KEYINPUT47), .B(G952), .Z(n1331) );
NAND2_X1 U1047 ( .A1(G237), .A2(G234), .ZN(n1252) );
INV_X1 U1048 ( .A(n1038), .ZN(n1046) );
NOR2_X1 U1049 ( .A1(n1079), .A2(n1080), .ZN(n1038) );
INV_X1 U1050 ( .A(n1095), .ZN(n1080) );
NAND2_X1 U1051 ( .A1(G214), .A2(n1332), .ZN(n1095) );
XNOR2_X1 U1052 ( .A(n1090), .B(n1093), .ZN(n1079) );
NAND2_X1 U1053 ( .A1(G210), .A2(n1332), .ZN(n1093) );
NAND2_X1 U1054 ( .A1(n1283), .A2(n1276), .ZN(n1332) );
INV_X1 U1055 ( .A(G902), .ZN(n1276) );
INV_X1 U1056 ( .A(G237), .ZN(n1283) );
NAND2_X1 U1057 ( .A1(n1333), .A2(n1334), .ZN(n1090) );
XOR2_X1 U1058 ( .A(KEYINPUT43), .B(G902), .Z(n1334) );
XOR2_X1 U1059 ( .A(n1335), .B(n1336), .Z(n1333) );
NOR2_X1 U1060 ( .A1(KEYINPUT28), .A2(n1190), .ZN(n1336) );
XNOR2_X1 U1061 ( .A(n1337), .B(n1143), .ZN(n1190) );
XNOR2_X1 U1062 ( .A(n1338), .B(G122), .ZN(n1143) );
NAND2_X1 U1063 ( .A1(KEYINPUT51), .A2(n1272), .ZN(n1338) );
XOR2_X1 U1064 ( .A(G110), .B(KEYINPUT55), .Z(n1272) );
NAND2_X1 U1065 ( .A1(n1339), .A2(KEYINPUT17), .ZN(n1337) );
XOR2_X1 U1066 ( .A(n1340), .B(n1144), .Z(n1339) );
XNOR2_X1 U1067 ( .A(n1341), .B(n1342), .ZN(n1144) );
XOR2_X1 U1068 ( .A(KEYINPUT20), .B(G119), .Z(n1342) );
XOR2_X1 U1069 ( .A(n1257), .B(G116), .Z(n1341) );
INV_X1 U1070 ( .A(G113), .ZN(n1257) );
NAND2_X1 U1071 ( .A1(KEYINPUT26), .A2(n1142), .ZN(n1340) );
XNOR2_X1 U1072 ( .A(n1183), .B(n1343), .ZN(n1142) );
XOR2_X1 U1073 ( .A(KEYINPUT49), .B(KEYINPUT40), .Z(n1343) );
XOR2_X1 U1074 ( .A(G101), .B(n1344), .Z(n1183) );
XOR2_X1 U1075 ( .A(G107), .B(G104), .Z(n1344) );
NAND3_X1 U1076 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1335) );
NAND2_X1 U1077 ( .A1(n1191), .A2(n1348), .ZN(n1347) );
INV_X1 U1078 ( .A(KEYINPUT37), .ZN(n1348) );
NAND3_X1 U1079 ( .A1(KEYINPUT37), .A2(n1349), .A3(n1192), .ZN(n1346) );
OR2_X1 U1080 ( .A1(n1192), .A2(n1349), .ZN(n1345) );
NOR2_X1 U1081 ( .A1(n1350), .A2(n1191), .ZN(n1349) );
XOR2_X1 U1082 ( .A(G125), .B(n1292), .Z(n1191) );
INV_X1 U1083 ( .A(n1175), .ZN(n1292) );
XOR2_X1 U1084 ( .A(n1351), .B(n1306), .Z(n1175) );
XOR2_X1 U1085 ( .A(G128), .B(G146), .Z(n1306) );
XNOR2_X1 U1086 ( .A(G143), .B(KEYINPUT24), .ZN(n1351) );
INV_X1 U1087 ( .A(KEYINPUT53), .ZN(n1350) );
NAND2_X1 U1088 ( .A1(G224), .A2(n1077), .ZN(n1192) );
INV_X1 U1089 ( .A(G953), .ZN(n1077) );
endmodule


