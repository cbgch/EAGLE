//Key = 1101000111110000000100000001011001111010101001110111000000111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421;

XNOR2_X1 U773 ( .A(G107), .B(n1082), .ZN(G9) );
NAND2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U775 ( .A(KEYINPUT17), .B(n1085), .Z(n1084) );
NOR2_X1 U776 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U777 ( .A1(n1088), .A2(n1089), .ZN(G75) );
NOR4_X1 U778 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1089) );
NOR2_X1 U779 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NOR2_X1 U780 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NOR2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
INV_X1 U782 ( .A(n1100), .ZN(n1099) );
NOR2_X1 U783 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
NOR2_X1 U784 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U785 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NOR2_X1 U786 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U787 ( .A1(n1109), .A2(n1083), .ZN(n1107) );
NOR2_X1 U788 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR2_X1 U789 ( .A1(n1112), .A2(n1113), .ZN(n1105) );
NOR2_X1 U790 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NOR2_X1 U791 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NOR3_X1 U792 ( .A1(n1113), .A2(n1118), .A3(n1108), .ZN(n1101) );
NOR2_X1 U793 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XOR2_X1 U794 ( .A(KEYINPUT12), .B(n1121), .Z(n1120) );
AND2_X1 U795 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
NOR4_X1 U796 ( .A1(n1124), .A2(n1108), .A3(n1113), .A4(n1104), .ZN(n1096) );
INV_X1 U797 ( .A(n1125), .ZN(n1108) );
NOR2_X1 U798 ( .A1(n1126), .A2(n1127), .ZN(n1124) );
NAND2_X1 U799 ( .A1(n1128), .A2(n1129), .ZN(n1090) );
NOR3_X1 U800 ( .A1(n1091), .A2(G952), .A3(n1092), .ZN(n1088) );
AND4_X1 U801 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1092) );
NOR3_X1 U802 ( .A1(n1134), .A2(n1116), .A3(n1135), .ZN(n1133) );
NAND3_X1 U803 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1134) );
XOR2_X1 U804 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U805 ( .A1(KEYINPUT4), .A2(n1141), .ZN(n1140) );
XOR2_X1 U806 ( .A(n1142), .B(KEYINPUT53), .Z(n1139) );
NAND2_X1 U807 ( .A1(n1143), .A2(n1144), .ZN(n1137) );
OR2_X1 U808 ( .A1(n1144), .A2(G469), .ZN(n1136) );
INV_X1 U809 ( .A(KEYINPUT22), .ZN(n1144) );
NOR3_X1 U810 ( .A1(n1123), .A2(n1145), .A3(n1146), .ZN(n1132) );
XNOR2_X1 U811 ( .A(n1147), .B(n1148), .ZN(n1131) );
NAND2_X1 U812 ( .A1(KEYINPUT3), .A2(n1149), .ZN(n1148) );
XOR2_X1 U813 ( .A(n1150), .B(n1151), .Z(n1130) );
NAND2_X1 U814 ( .A1(KEYINPUT35), .A2(n1152), .ZN(n1151) );
INV_X1 U815 ( .A(n1153), .ZN(n1091) );
XOR2_X1 U816 ( .A(n1154), .B(n1155), .Z(G72) );
NOR2_X1 U817 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U818 ( .A(n1158), .B(n1159), .Z(n1157) );
XNOR2_X1 U819 ( .A(n1160), .B(n1161), .ZN(n1159) );
XNOR2_X1 U820 ( .A(n1162), .B(n1163), .ZN(n1158) );
XNOR2_X1 U821 ( .A(n1164), .B(n1165), .ZN(n1163) );
NOR2_X1 U822 ( .A1(G140), .A2(KEYINPUT55), .ZN(n1165) );
NAND2_X1 U823 ( .A1(n1166), .A2(n1167), .ZN(n1154) );
NAND2_X1 U824 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND3_X1 U825 ( .A1(KEYINPUT59), .A2(n1170), .A3(G953), .ZN(n1166) );
NAND2_X1 U826 ( .A1(G900), .A2(G227), .ZN(n1170) );
NAND2_X1 U827 ( .A1(n1171), .A2(n1172), .ZN(G69) );
NAND2_X1 U828 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NAND2_X1 U829 ( .A1(G953), .A2(n1175), .ZN(n1174) );
NAND3_X1 U830 ( .A1(G953), .A2(n1176), .A3(n1177), .ZN(n1171) );
INV_X1 U831 ( .A(n1173), .ZN(n1177) );
XNOR2_X1 U832 ( .A(n1178), .B(n1179), .ZN(n1173) );
NOR2_X1 U833 ( .A1(n1180), .A2(G953), .ZN(n1179) );
NOR2_X1 U834 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND2_X1 U835 ( .A1(n1183), .A2(n1184), .ZN(n1178) );
NAND2_X1 U836 ( .A1(G953), .A2(n1185), .ZN(n1184) );
XNOR2_X1 U837 ( .A(n1186), .B(n1187), .ZN(n1183) );
NAND2_X1 U838 ( .A1(n1188), .A2(n1189), .ZN(n1186) );
XOR2_X1 U839 ( .A(KEYINPUT61), .B(KEYINPUT45), .Z(n1189) );
NAND2_X1 U840 ( .A1(G898), .A2(G224), .ZN(n1176) );
NOR2_X1 U841 ( .A1(n1190), .A2(n1191), .ZN(G66) );
NOR3_X1 U842 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1191) );
NOR3_X1 U843 ( .A1(n1195), .A2(n1142), .A3(n1196), .ZN(n1194) );
NOR2_X1 U844 ( .A1(n1197), .A2(n1198), .ZN(n1193) );
NOR2_X1 U845 ( .A1(n1199), .A2(n1142), .ZN(n1198) );
NOR2_X1 U846 ( .A1(n1190), .A2(n1200), .ZN(G63) );
XOR2_X1 U847 ( .A(n1201), .B(n1202), .Z(n1200) );
XOR2_X1 U848 ( .A(KEYINPUT29), .B(n1203), .Z(n1202) );
NOR2_X1 U849 ( .A1(n1204), .A2(n1196), .ZN(n1203) );
NOR2_X1 U850 ( .A1(n1190), .A2(n1205), .ZN(G60) );
NOR3_X1 U851 ( .A1(n1147), .A2(n1206), .A3(n1207), .ZN(n1205) );
NOR3_X1 U852 ( .A1(n1208), .A2(n1196), .A3(n1149), .ZN(n1207) );
NOR2_X1 U853 ( .A1(n1209), .A2(n1210), .ZN(n1206) );
NOR2_X1 U854 ( .A1(n1199), .A2(n1149), .ZN(n1209) );
INV_X1 U855 ( .A(G475), .ZN(n1149) );
XNOR2_X1 U856 ( .A(G104), .B(n1211), .ZN(G6) );
NOR2_X1 U857 ( .A1(n1190), .A2(n1212), .ZN(G57) );
XOR2_X1 U858 ( .A(n1213), .B(n1214), .Z(n1212) );
XNOR2_X1 U859 ( .A(n1215), .B(n1216), .ZN(n1214) );
NOR2_X1 U860 ( .A1(KEYINPUT39), .A2(n1217), .ZN(n1216) );
XOR2_X1 U861 ( .A(n1218), .B(n1219), .Z(n1213) );
NOR2_X1 U862 ( .A1(n1220), .A2(n1196), .ZN(n1219) );
XNOR2_X1 U863 ( .A(n1221), .B(n1222), .ZN(n1218) );
NOR2_X1 U864 ( .A1(KEYINPUT57), .A2(n1223), .ZN(n1222) );
NOR2_X1 U865 ( .A1(KEYINPUT16), .A2(n1160), .ZN(n1221) );
NOR2_X1 U866 ( .A1(n1190), .A2(n1224), .ZN(G54) );
XOR2_X1 U867 ( .A(n1225), .B(n1226), .Z(n1224) );
NOR2_X1 U868 ( .A1(KEYINPUT56), .A2(n1227), .ZN(n1226) );
XOR2_X1 U869 ( .A(n1228), .B(n1229), .Z(n1227) );
XOR2_X1 U870 ( .A(n1230), .B(n1231), .Z(n1229) );
NOR2_X1 U871 ( .A1(G110), .A2(KEYINPUT54), .ZN(n1231) );
NOR3_X1 U872 ( .A1(n1232), .A2(KEYINPUT13), .A3(G953), .ZN(n1230) );
INV_X1 U873 ( .A(G227), .ZN(n1232) );
XOR2_X1 U874 ( .A(G140), .B(n1233), .Z(n1228) );
NOR2_X1 U875 ( .A1(KEYINPUT37), .A2(n1234), .ZN(n1233) );
XNOR2_X1 U876 ( .A(n1235), .B(n1236), .ZN(n1234) );
XOR2_X1 U877 ( .A(n1237), .B(KEYINPUT21), .Z(n1235) );
NAND3_X1 U878 ( .A1(G469), .A2(n1238), .A3(n1239), .ZN(n1225) );
XNOR2_X1 U879 ( .A(G902), .B(KEYINPUT10), .ZN(n1239) );
NOR2_X1 U880 ( .A1(n1190), .A2(n1240), .ZN(G51) );
NOR3_X1 U881 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1240) );
NOR3_X1 U882 ( .A1(n1244), .A2(n1150), .A3(n1196), .ZN(n1243) );
NAND2_X1 U883 ( .A1(G902), .A2(n1238), .ZN(n1196) );
NOR2_X1 U884 ( .A1(n1245), .A2(n1246), .ZN(n1242) );
NOR2_X1 U885 ( .A1(n1199), .A2(n1150), .ZN(n1245) );
INV_X1 U886 ( .A(n1238), .ZN(n1199) );
NAND2_X1 U887 ( .A1(n1128), .A2(n1247), .ZN(n1238) );
XOR2_X1 U888 ( .A(KEYINPUT31), .B(n1129), .Z(n1247) );
NOR2_X1 U889 ( .A1(n1182), .A2(n1248), .ZN(n1129) );
XOR2_X1 U890 ( .A(KEYINPUT52), .B(n1181), .Z(n1248) );
NAND4_X1 U891 ( .A1(n1249), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1181) );
NAND3_X1 U892 ( .A1(n1115), .A2(n1126), .A3(n1253), .ZN(n1249) );
NAND3_X1 U893 ( .A1(n1254), .A2(n1211), .A3(n1255), .ZN(n1182) );
NAND2_X1 U894 ( .A1(KEYINPUT30), .A2(n1256), .ZN(n1255) );
NAND3_X1 U895 ( .A1(n1083), .A2(n1257), .A3(n1127), .ZN(n1211) );
NAND2_X1 U896 ( .A1(n1083), .A2(n1258), .ZN(n1254) );
NAND3_X1 U897 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1258) );
NAND2_X1 U898 ( .A1(n1126), .A2(n1257), .ZN(n1261) );
INV_X1 U899 ( .A(n1086), .ZN(n1257) );
NAND3_X1 U900 ( .A1(n1125), .A2(n1262), .A3(n1121), .ZN(n1086) );
OR3_X1 U901 ( .A1(n1121), .A2(KEYINPUT30), .A3(n1263), .ZN(n1259) );
INV_X1 U902 ( .A(n1168), .ZN(n1128) );
NAND4_X1 U903 ( .A1(n1264), .A2(n1265), .A3(n1266), .A4(n1267), .ZN(n1168) );
AND4_X1 U904 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1267) );
AND2_X1 U905 ( .A1(n1272), .A2(n1273), .ZN(n1266) );
NAND3_X1 U906 ( .A1(n1274), .A2(n1126), .A3(n1275), .ZN(n1264) );
NOR2_X1 U907 ( .A1(n1169), .A2(G952), .ZN(n1190) );
XNOR2_X1 U908 ( .A(G146), .B(n1270), .ZN(G48) );
NAND3_X1 U909 ( .A1(n1127), .A2(n1083), .A3(n1276), .ZN(n1270) );
XNOR2_X1 U910 ( .A(G143), .B(n1265), .ZN(G45) );
NAND4_X1 U911 ( .A1(n1277), .A2(n1274), .A3(n1278), .A4(n1083), .ZN(n1265) );
XOR2_X1 U912 ( .A(G140), .B(n1279), .Z(G42) );
NOR2_X1 U913 ( .A1(KEYINPUT41), .A2(n1273), .ZN(n1279) );
NAND3_X1 U914 ( .A1(n1275), .A2(n1121), .A3(n1280), .ZN(n1273) );
XNOR2_X1 U915 ( .A(G137), .B(n1269), .ZN(G39) );
NAND3_X1 U916 ( .A1(n1276), .A2(n1275), .A3(n1100), .ZN(n1269) );
XOR2_X1 U917 ( .A(n1281), .B(n1282), .Z(G36) );
NOR2_X1 U918 ( .A1(KEYINPUT5), .A2(n1283), .ZN(n1282) );
NOR3_X1 U919 ( .A1(n1284), .A2(n1087), .A3(n1285), .ZN(n1281) );
INV_X1 U920 ( .A(n1126), .ZN(n1087) );
XNOR2_X1 U921 ( .A(KEYINPUT49), .B(n1113), .ZN(n1284) );
INV_X1 U922 ( .A(n1275), .ZN(n1113) );
XNOR2_X1 U923 ( .A(G131), .B(n1268), .ZN(G33) );
NAND3_X1 U924 ( .A1(n1274), .A2(n1127), .A3(n1275), .ZN(n1268) );
NOR2_X1 U925 ( .A1(n1110), .A2(n1145), .ZN(n1275) );
INV_X1 U926 ( .A(n1111), .ZN(n1145) );
INV_X1 U927 ( .A(n1285), .ZN(n1274) );
NAND3_X1 U928 ( .A1(n1121), .A2(n1286), .A3(n1115), .ZN(n1285) );
NAND3_X1 U929 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(G30) );
NAND2_X1 U930 ( .A1(G128), .A2(n1272), .ZN(n1289) );
NAND2_X1 U931 ( .A1(KEYINPUT20), .A2(n1290), .ZN(n1288) );
NAND2_X1 U932 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XNOR2_X1 U933 ( .A(KEYINPUT19), .B(n1293), .ZN(n1292) );
NAND2_X1 U934 ( .A1(n1294), .A2(n1295), .ZN(n1287) );
INV_X1 U935 ( .A(KEYINPUT20), .ZN(n1295) );
NAND2_X1 U936 ( .A1(n1296), .A2(n1297), .ZN(n1294) );
NAND3_X1 U937 ( .A1(KEYINPUT19), .A2(n1291), .A3(n1293), .ZN(n1297) );
INV_X1 U938 ( .A(n1272), .ZN(n1291) );
NAND3_X1 U939 ( .A1(n1083), .A2(n1126), .A3(n1276), .ZN(n1272) );
AND4_X1 U940 ( .A1(n1298), .A2(n1121), .A3(n1116), .A4(n1286), .ZN(n1276) );
OR2_X1 U941 ( .A1(n1293), .A2(KEYINPUT19), .ZN(n1296) );
XNOR2_X1 U942 ( .A(G101), .B(n1299), .ZN(G3) );
NAND2_X1 U943 ( .A1(n1300), .A2(n1083), .ZN(n1299) );
XOR2_X1 U944 ( .A(n1260), .B(KEYINPUT8), .Z(n1300) );
NAND4_X1 U945 ( .A1(n1100), .A2(n1115), .A3(n1121), .A4(n1262), .ZN(n1260) );
XNOR2_X1 U946 ( .A(G125), .B(n1271), .ZN(G27) );
NAND3_X1 U947 ( .A1(n1280), .A2(n1083), .A3(n1301), .ZN(n1271) );
AND4_X1 U948 ( .A1(n1298), .A2(n1127), .A3(n1302), .A4(n1286), .ZN(n1280) );
NAND2_X1 U949 ( .A1(n1095), .A2(n1303), .ZN(n1286) );
NAND3_X1 U950 ( .A1(G902), .A2(n1304), .A3(n1156), .ZN(n1303) );
AND2_X1 U951 ( .A1(G953), .A2(n1305), .ZN(n1156) );
XOR2_X1 U952 ( .A(KEYINPUT47), .B(G900), .Z(n1305) );
XNOR2_X1 U953 ( .A(G122), .B(n1250), .ZN(G24) );
NAND4_X1 U954 ( .A1(n1277), .A2(n1253), .A3(n1278), .A4(n1125), .ZN(n1250) );
NOR2_X1 U955 ( .A1(n1116), .A2(n1298), .ZN(n1125) );
NAND2_X1 U956 ( .A1(n1306), .A2(n1307), .ZN(G21) );
OR2_X1 U957 ( .A1(n1251), .A2(G119), .ZN(n1307) );
XOR2_X1 U958 ( .A(n1308), .B(KEYINPUT26), .Z(n1306) );
NAND2_X1 U959 ( .A1(G119), .A2(n1251), .ZN(n1308) );
NAND4_X1 U960 ( .A1(n1253), .A2(n1100), .A3(n1298), .A4(n1116), .ZN(n1251) );
NAND2_X1 U961 ( .A1(n1309), .A2(n1310), .ZN(G18) );
NAND2_X1 U962 ( .A1(G116), .A2(n1311), .ZN(n1310) );
XOR2_X1 U963 ( .A(KEYINPUT36), .B(n1312), .Z(n1309) );
NOR2_X1 U964 ( .A1(G116), .A2(n1311), .ZN(n1312) );
NAND4_X1 U965 ( .A1(n1313), .A2(n1262), .A3(n1126), .A4(n1314), .ZN(n1311) );
NOR2_X1 U966 ( .A1(n1315), .A2(n1104), .ZN(n1314) );
NOR2_X1 U967 ( .A1(n1316), .A2(n1277), .ZN(n1126) );
XOR2_X1 U968 ( .A(KEYINPUT14), .B(n1083), .Z(n1313) );
XNOR2_X1 U969 ( .A(G113), .B(n1252), .ZN(G15) );
NAND3_X1 U970 ( .A1(n1127), .A2(n1115), .A3(n1253), .ZN(n1252) );
AND3_X1 U971 ( .A1(n1083), .A2(n1262), .A3(n1301), .ZN(n1253) );
INV_X1 U972 ( .A(n1104), .ZN(n1301) );
NAND2_X1 U973 ( .A1(n1122), .A2(n1317), .ZN(n1104) );
INV_X1 U974 ( .A(n1315), .ZN(n1115) );
NAND2_X1 U975 ( .A1(n1318), .A2(n1116), .ZN(n1315) );
XNOR2_X1 U976 ( .A(KEYINPUT44), .B(n1298), .ZN(n1318) );
AND2_X1 U977 ( .A1(n1277), .A2(n1319), .ZN(n1127) );
XNOR2_X1 U978 ( .A(KEYINPUT15), .B(n1278), .ZN(n1319) );
XOR2_X1 U979 ( .A(G110), .B(n1256), .Z(G12) );
AND3_X1 U980 ( .A1(n1083), .A2(n1121), .A3(n1320), .ZN(n1256) );
INV_X1 U981 ( .A(n1263), .ZN(n1320) );
NAND4_X1 U982 ( .A1(n1298), .A2(n1100), .A3(n1302), .A4(n1262), .ZN(n1263) );
NAND2_X1 U983 ( .A1(n1095), .A2(n1321), .ZN(n1262) );
NAND4_X1 U984 ( .A1(G953), .A2(G902), .A3(n1304), .A4(n1185), .ZN(n1321) );
INV_X1 U985 ( .A(G898), .ZN(n1185) );
NAND3_X1 U986 ( .A1(n1153), .A2(n1304), .A3(G952), .ZN(n1095) );
NAND2_X1 U987 ( .A1(G237), .A2(G234), .ZN(n1304) );
XOR2_X1 U988 ( .A(G953), .B(KEYINPUT7), .Z(n1153) );
INV_X1 U989 ( .A(n1116), .ZN(n1302) );
XOR2_X1 U990 ( .A(n1322), .B(n1220), .Z(n1116) );
INV_X1 U991 ( .A(G472), .ZN(n1220) );
NAND2_X1 U992 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U993 ( .A(n1325), .B(n1217), .Z(n1323) );
XNOR2_X1 U994 ( .A(n1326), .B(G101), .ZN(n1217) );
NAND3_X1 U995 ( .A1(n1327), .A2(n1169), .A3(G210), .ZN(n1326) );
NAND3_X1 U996 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1325) );
NAND2_X1 U997 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NAND2_X1 U998 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
XNOR2_X1 U999 ( .A(KEYINPUT42), .B(n1223), .ZN(n1331) );
NAND4_X1 U1000 ( .A1(n1335), .A2(n1334), .A3(n1336), .A4(n1333), .ZN(n1329) );
INV_X1 U1001 ( .A(n1337), .ZN(n1333) );
XOR2_X1 U1002 ( .A(KEYINPUT42), .B(n1223), .Z(n1336) );
XNOR2_X1 U1003 ( .A(n1338), .B(n1339), .ZN(n1223) );
NOR2_X1 U1004 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
NOR2_X1 U1005 ( .A1(G119), .A2(n1342), .ZN(n1341) );
XNOR2_X1 U1006 ( .A(KEYINPUT60), .B(n1343), .ZN(n1342) );
INV_X1 U1007 ( .A(KEYINPUT62), .ZN(n1334) );
INV_X1 U1008 ( .A(KEYINPUT25), .ZN(n1335) );
NAND2_X1 U1009 ( .A1(KEYINPUT25), .A2(n1337), .ZN(n1328) );
XNOR2_X1 U1010 ( .A(n1215), .B(n1160), .ZN(n1337) );
NOR2_X1 U1011 ( .A1(n1278), .A2(n1277), .ZN(n1100) );
XNOR2_X1 U1012 ( .A(n1147), .B(n1344), .ZN(n1277) );
NOR2_X1 U1013 ( .A1(G475), .A2(KEYINPUT43), .ZN(n1344) );
NOR2_X1 U1014 ( .A1(n1210), .A2(G902), .ZN(n1147) );
INV_X1 U1015 ( .A(n1208), .ZN(n1210) );
XNOR2_X1 U1016 ( .A(n1345), .B(n1346), .ZN(n1208) );
XNOR2_X1 U1017 ( .A(G104), .B(n1347), .ZN(n1346) );
NAND2_X1 U1018 ( .A1(n1348), .A2(KEYINPUT58), .ZN(n1347) );
XOR2_X1 U1019 ( .A(n1349), .B(n1350), .Z(n1348) );
XNOR2_X1 U1020 ( .A(KEYINPUT27), .B(n1351), .ZN(n1350) );
INV_X1 U1021 ( .A(G131), .ZN(n1351) );
XOR2_X1 U1022 ( .A(n1352), .B(n1353), .Z(n1349) );
NAND2_X1 U1023 ( .A1(n1354), .A2(n1355), .ZN(n1352) );
NAND4_X1 U1024 ( .A1(G143), .A2(G214), .A3(n1327), .A4(n1169), .ZN(n1355) );
XOR2_X1 U1025 ( .A(n1356), .B(KEYINPUT24), .Z(n1354) );
NAND2_X1 U1026 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
NAND3_X1 U1027 ( .A1(n1327), .A2(n1169), .A3(G214), .ZN(n1358) );
XNOR2_X1 U1028 ( .A(G113), .B(G122), .ZN(n1345) );
INV_X1 U1029 ( .A(n1316), .ZN(n1278) );
XOR2_X1 U1030 ( .A(n1135), .B(KEYINPUT1), .Z(n1316) );
XOR2_X1 U1031 ( .A(n1359), .B(n1204), .Z(n1135) );
INV_X1 U1032 ( .A(G478), .ZN(n1204) );
NAND2_X1 U1033 ( .A1(n1201), .A2(n1324), .ZN(n1359) );
XNOR2_X1 U1034 ( .A(n1360), .B(n1361), .ZN(n1201) );
XNOR2_X1 U1035 ( .A(n1343), .B(n1362), .ZN(n1361) );
XNOR2_X1 U1036 ( .A(n1283), .B(G122), .ZN(n1362) );
INV_X1 U1037 ( .A(G134), .ZN(n1283) );
XOR2_X1 U1038 ( .A(n1363), .B(n1364), .Z(n1360) );
XOR2_X1 U1039 ( .A(n1365), .B(G107), .Z(n1363) );
NAND2_X1 U1040 ( .A1(G217), .A2(n1366), .ZN(n1365) );
INV_X1 U1041 ( .A(n1117), .ZN(n1298) );
XNOR2_X1 U1042 ( .A(n1142), .B(n1367), .ZN(n1117) );
XNOR2_X1 U1043 ( .A(KEYINPUT46), .B(n1141), .ZN(n1367) );
INV_X1 U1044 ( .A(n1192), .ZN(n1141) );
NOR2_X1 U1045 ( .A1(n1197), .A2(G902), .ZN(n1192) );
INV_X1 U1046 ( .A(n1195), .ZN(n1197) );
NAND2_X1 U1047 ( .A1(n1368), .A2(n1369), .ZN(n1195) );
NAND2_X1 U1048 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
XOR2_X1 U1049 ( .A(KEYINPUT0), .B(n1372), .Z(n1368) );
NOR2_X1 U1050 ( .A1(n1370), .A2(n1371), .ZN(n1372) );
XNOR2_X1 U1051 ( .A(n1373), .B(G137), .ZN(n1371) );
NAND2_X1 U1052 ( .A1(G221), .A2(n1366), .ZN(n1373) );
AND2_X1 U1053 ( .A1(G234), .A2(n1169), .ZN(n1366) );
XNOR2_X1 U1054 ( .A(n1374), .B(n1375), .ZN(n1370) );
XNOR2_X1 U1055 ( .A(n1293), .B(G119), .ZN(n1375) );
INV_X1 U1056 ( .A(G128), .ZN(n1293) );
XNOR2_X1 U1057 ( .A(n1353), .B(n1376), .ZN(n1374) );
NOR2_X1 U1058 ( .A1(G110), .A2(KEYINPUT6), .ZN(n1376) );
XOR2_X1 U1059 ( .A(G125), .B(n1377), .Z(n1353) );
XNOR2_X1 U1060 ( .A(n1378), .B(G140), .ZN(n1377) );
INV_X1 U1061 ( .A(G146), .ZN(n1378) );
NAND2_X1 U1062 ( .A1(G217), .A2(n1379), .ZN(n1142) );
NOR2_X1 U1063 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
INV_X1 U1064 ( .A(n1317), .ZN(n1123) );
NAND2_X1 U1065 ( .A1(G221), .A2(n1379), .ZN(n1317) );
NAND2_X1 U1066 ( .A1(G234), .A2(n1324), .ZN(n1379) );
NOR2_X1 U1067 ( .A1(n1146), .A2(n1143), .ZN(n1122) );
AND2_X1 U1068 ( .A1(G469), .A2(n1380), .ZN(n1143) );
NOR2_X1 U1069 ( .A1(n1380), .A2(G469), .ZN(n1146) );
NAND2_X1 U1070 ( .A1(n1381), .A2(n1324), .ZN(n1380) );
XOR2_X1 U1071 ( .A(n1382), .B(n1383), .Z(n1381) );
XOR2_X1 U1072 ( .A(n1384), .B(n1237), .Z(n1383) );
XOR2_X1 U1073 ( .A(n1385), .B(n1386), .Z(n1237) );
XOR2_X1 U1074 ( .A(G107), .B(G104), .Z(n1386) );
XNOR2_X1 U1075 ( .A(n1387), .B(G101), .ZN(n1385) );
NAND2_X1 U1076 ( .A1(KEYINPUT38), .A2(n1215), .ZN(n1384) );
INV_X1 U1077 ( .A(n1236), .ZN(n1215) );
NAND2_X1 U1078 ( .A1(n1388), .A2(n1389), .ZN(n1236) );
OR2_X1 U1079 ( .A1(n1161), .A2(n1162), .ZN(n1389) );
NAND2_X1 U1080 ( .A1(n1390), .A2(n1161), .ZN(n1388) );
XNOR2_X1 U1081 ( .A(G134), .B(KEYINPUT33), .ZN(n1161) );
XOR2_X1 U1082 ( .A(KEYINPUT2), .B(n1162), .Z(n1390) );
XOR2_X1 U1083 ( .A(G131), .B(G137), .Z(n1162) );
XOR2_X1 U1084 ( .A(n1391), .B(n1392), .Z(n1382) );
XOR2_X1 U1085 ( .A(n1393), .B(KEYINPUT11), .Z(n1392) );
NAND2_X1 U1086 ( .A1(n1394), .A2(n1395), .ZN(n1393) );
NAND2_X1 U1087 ( .A1(G110), .A2(n1396), .ZN(n1395) );
XOR2_X1 U1088 ( .A(n1397), .B(KEYINPUT48), .Z(n1394) );
OR2_X1 U1089 ( .A1(n1396), .A2(G110), .ZN(n1397) );
XOR2_X1 U1090 ( .A(G140), .B(KEYINPUT50), .Z(n1396) );
NAND3_X1 U1091 ( .A1(G227), .A2(n1169), .A3(KEYINPUT40), .ZN(n1391) );
INV_X1 U1092 ( .A(G953), .ZN(n1169) );
AND2_X1 U1093 ( .A1(n1110), .A2(n1111), .ZN(n1083) );
NAND2_X1 U1094 ( .A1(n1398), .A2(G214), .ZN(n1111) );
XOR2_X1 U1095 ( .A(n1399), .B(KEYINPUT23), .Z(n1398) );
XOR2_X1 U1096 ( .A(n1150), .B(n1400), .Z(n1110) );
NOR2_X1 U1097 ( .A1(n1401), .A2(n1402), .ZN(n1400) );
NOR2_X1 U1098 ( .A1(KEYINPUT51), .A2(n1241), .ZN(n1402) );
NOR2_X1 U1099 ( .A1(KEYINPUT63), .A2(n1152), .ZN(n1401) );
INV_X1 U1100 ( .A(n1241), .ZN(n1152) );
NOR2_X1 U1101 ( .A1(n1246), .A2(G902), .ZN(n1241) );
INV_X1 U1102 ( .A(n1244), .ZN(n1246) );
XNOR2_X1 U1103 ( .A(n1403), .B(n1404), .ZN(n1244) );
XOR2_X1 U1104 ( .A(n1405), .B(n1406), .Z(n1404) );
XNOR2_X1 U1105 ( .A(KEYINPUT32), .B(n1164), .ZN(n1406) );
INV_X1 U1106 ( .A(G125), .ZN(n1164) );
NOR2_X1 U1107 ( .A1(G953), .A2(n1175), .ZN(n1405) );
INV_X1 U1108 ( .A(G224), .ZN(n1175) );
XOR2_X1 U1109 ( .A(n1407), .B(n1187), .Z(n1403) );
XOR2_X1 U1110 ( .A(G122), .B(G110), .Z(n1187) );
XNOR2_X1 U1111 ( .A(n1188), .B(n1160), .ZN(n1407) );
INV_X1 U1112 ( .A(n1387), .ZN(n1160) );
XOR2_X1 U1113 ( .A(G146), .B(n1364), .Z(n1387) );
XNOR2_X1 U1114 ( .A(n1357), .B(G128), .ZN(n1364) );
INV_X1 U1115 ( .A(G143), .ZN(n1357) );
XOR2_X1 U1116 ( .A(n1408), .B(n1409), .Z(n1188) );
NOR2_X1 U1117 ( .A1(G101), .A2(KEYINPUT18), .ZN(n1409) );
XOR2_X1 U1118 ( .A(n1410), .B(n1411), .Z(n1408) );
NOR2_X1 U1119 ( .A1(n1412), .A2(n1413), .ZN(n1411) );
XOR2_X1 U1120 ( .A(KEYINPUT28), .B(n1414), .Z(n1413) );
NOR2_X1 U1121 ( .A1(G107), .A2(n1415), .ZN(n1414) );
AND2_X1 U1122 ( .A1(n1415), .A2(G107), .ZN(n1412) );
XOR2_X1 U1123 ( .A(G104), .B(KEYINPUT9), .Z(n1415) );
NAND2_X1 U1124 ( .A1(n1416), .A2(n1417), .ZN(n1410) );
NAND2_X1 U1125 ( .A1(n1418), .A2(n1338), .ZN(n1417) );
XNOR2_X1 U1126 ( .A(G116), .B(G119), .ZN(n1418) );
XOR2_X1 U1127 ( .A(KEYINPUT34), .B(n1419), .Z(n1416) );
NOR2_X1 U1128 ( .A1(n1420), .A2(n1338), .ZN(n1419) );
INV_X1 U1129 ( .A(G113), .ZN(n1338) );
NOR2_X1 U1130 ( .A1(n1421), .A2(n1340), .ZN(n1420) );
AND2_X1 U1131 ( .A1(G119), .A2(n1343), .ZN(n1340) );
NOR2_X1 U1132 ( .A1(G119), .A2(n1343), .ZN(n1421) );
INV_X1 U1133 ( .A(G116), .ZN(n1343) );
NAND2_X1 U1134 ( .A1(G210), .A2(n1399), .ZN(n1150) );
NAND2_X1 U1135 ( .A1(n1324), .A2(n1327), .ZN(n1399) );
INV_X1 U1136 ( .A(G237), .ZN(n1327) );
INV_X1 U1137 ( .A(G902), .ZN(n1324) );
endmodule


