//Key = 1101001011101100010010011011110000101110001111001000010110111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336;

XNOR2_X1 U736 ( .A(G107), .B(n1021), .ZN(G9) );
NOR2_X1 U737 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR3_X1 U738 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
NOR2_X1 U739 ( .A1(KEYINPUT12), .A2(n1027), .ZN(n1025) );
NOR4_X1 U740 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1027) );
INV_X1 U741 ( .A(n1032), .ZN(n1029) );
NAND2_X1 U742 ( .A1(n1033), .A2(n1034), .ZN(n1028) );
NAND3_X1 U743 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1024) );
NAND2_X1 U744 ( .A1(n1033), .A2(n1038), .ZN(n1037) );
NAND2_X1 U745 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND3_X1 U746 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NAND2_X1 U747 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NAND2_X1 U748 ( .A1(n1034), .A2(n1046), .ZN(n1045) );
NAND2_X1 U749 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U750 ( .A1(KEYINPUT12), .A2(n1032), .ZN(n1048) );
NAND2_X1 U751 ( .A1(n1049), .A2(n1050), .ZN(n1044) );
NAND2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND3_X1 U754 ( .A1(n1049), .A2(n1055), .A3(n1034), .ZN(n1039) );
NAND2_X1 U755 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U756 ( .A1(n1041), .A2(n1058), .ZN(n1057) );
OR2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U758 ( .A1(n1043), .A2(n1061), .ZN(n1056) );
NAND2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
INV_X1 U761 ( .A(n1066), .ZN(n1062) );
INV_X1 U762 ( .A(n1067), .ZN(n1033) );
NOR3_X1 U763 ( .A1(n1068), .A2(G953), .A3(G952), .ZN(n1022) );
INV_X1 U764 ( .A(n1035), .ZN(n1068) );
NAND4_X1 U765 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1035) );
NOR4_X1 U766 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1072) );
XNOR2_X1 U767 ( .A(G469), .B(n1077), .ZN(n1076) );
XNOR2_X1 U768 ( .A(n1078), .B(n1079), .ZN(n1073) );
XNOR2_X1 U769 ( .A(n1080), .B(KEYINPUT42), .ZN(n1078) );
NOR3_X1 U770 ( .A1(n1053), .A2(n1081), .A3(n1064), .ZN(n1071) );
NAND2_X1 U771 ( .A1(G475), .A2(n1082), .ZN(n1070) );
XNOR2_X1 U772 ( .A(n1083), .B(n1084), .ZN(n1069) );
XNOR2_X1 U773 ( .A(n1085), .B(KEYINPUT34), .ZN(n1084) );
NAND2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(G72) );
NAND2_X1 U775 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NAND2_X1 U776 ( .A1(G900), .A2(n1089), .ZN(n1088) );
XOR2_X1 U777 ( .A(n1090), .B(n1091), .Z(n1089) );
XOR2_X1 U778 ( .A(KEYINPUT31), .B(G227), .Z(n1091) );
NAND2_X1 U779 ( .A1(n1092), .A2(n1036), .ZN(n1086) );
XOR2_X1 U780 ( .A(n1093), .B(n1090), .Z(n1092) );
XNOR2_X1 U781 ( .A(n1094), .B(n1095), .ZN(n1090) );
XOR2_X1 U782 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U783 ( .A1(KEYINPUT48), .A2(n1098), .ZN(n1097) );
NAND2_X1 U784 ( .A1(n1099), .A2(n1100), .ZN(n1096) );
XOR2_X1 U785 ( .A(n1101), .B(KEYINPUT23), .Z(n1099) );
NAND2_X1 U786 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
OR3_X1 U787 ( .A1(n1104), .A2(G131), .A3(KEYINPUT15), .ZN(n1103) );
NAND2_X1 U788 ( .A1(KEYINPUT15), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U789 ( .A(G125), .B(n1105), .ZN(n1094) );
XOR2_X1 U790 ( .A(KEYINPUT36), .B(G140), .Z(n1105) );
NOR2_X1 U791 ( .A1(n1106), .A2(KEYINPUT19), .ZN(n1093) );
XOR2_X1 U792 ( .A(n1107), .B(n1108), .Z(G69) );
XOR2_X1 U793 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND2_X1 U794 ( .A1(G953), .A2(n1111), .ZN(n1110) );
NAND2_X1 U795 ( .A1(G224), .A2(n1112), .ZN(n1111) );
XNOR2_X1 U796 ( .A(KEYINPUT4), .B(n1113), .ZN(n1112) );
NAND2_X1 U797 ( .A1(n1114), .A2(n1115), .ZN(n1109) );
NAND2_X1 U798 ( .A1(G953), .A2(n1113), .ZN(n1115) );
XOR2_X1 U799 ( .A(n1116), .B(n1117), .Z(n1114) );
NOR2_X1 U800 ( .A1(KEYINPUT30), .A2(n1118), .ZN(n1117) );
NOR2_X1 U801 ( .A1(n1119), .A2(G953), .ZN(n1107) );
NOR2_X1 U802 ( .A1(n1120), .A2(n1121), .ZN(G66) );
XOR2_X1 U803 ( .A(KEYINPUT32), .B(n1122), .Z(n1121) );
NOR3_X1 U804 ( .A1(n1085), .A2(n1123), .A3(n1124), .ZN(n1120) );
AND3_X1 U805 ( .A1(n1125), .A2(n1083), .A3(n1126), .ZN(n1124) );
NOR2_X1 U806 ( .A1(n1127), .A2(n1125), .ZN(n1123) );
AND2_X1 U807 ( .A1(n1026), .A2(n1083), .ZN(n1127) );
NOR3_X1 U808 ( .A1(n1122), .A2(n1128), .A3(n1129), .ZN(G63) );
NOR3_X1 U809 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1129) );
NOR2_X1 U810 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
INV_X1 U811 ( .A(KEYINPUT5), .ZN(n1134) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1128) );
NOR2_X1 U813 ( .A1(KEYINPUT5), .A2(n1133), .ZN(n1135) );
XOR2_X1 U814 ( .A(n1131), .B(KEYINPUT57), .Z(n1133) );
AND2_X1 U815 ( .A1(n1126), .A2(G478), .ZN(n1131) );
NOR2_X1 U816 ( .A1(n1122), .A2(n1137), .ZN(G60) );
XNOR2_X1 U817 ( .A(n1138), .B(n1139), .ZN(n1137) );
NAND2_X1 U818 ( .A1(KEYINPUT24), .A2(n1140), .ZN(n1138) );
NAND2_X1 U819 ( .A1(n1126), .A2(G475), .ZN(n1140) );
XNOR2_X1 U820 ( .A(G104), .B(n1141), .ZN(G6) );
NOR2_X1 U821 ( .A1(n1122), .A2(n1142), .ZN(G57) );
XOR2_X1 U822 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U823 ( .A(n1145), .B(n1146), .Z(n1144) );
XNOR2_X1 U824 ( .A(n1147), .B(n1148), .ZN(n1146) );
NOR2_X1 U825 ( .A1(KEYINPUT35), .A2(n1149), .ZN(n1148) );
AND2_X1 U826 ( .A1(G472), .A2(n1126), .ZN(n1145) );
INV_X1 U827 ( .A(n1150), .ZN(n1126) );
XNOR2_X1 U828 ( .A(n1151), .B(n1152), .ZN(n1143) );
NOR2_X1 U829 ( .A1(n1122), .A2(n1153), .ZN(G54) );
XOR2_X1 U830 ( .A(n1154), .B(n1155), .Z(n1153) );
XNOR2_X1 U831 ( .A(n1156), .B(n1157), .ZN(n1155) );
XNOR2_X1 U832 ( .A(G110), .B(KEYINPUT28), .ZN(n1157) );
XOR2_X1 U833 ( .A(n1158), .B(n1159), .Z(n1154) );
XOR2_X1 U834 ( .A(n1160), .B(n1161), .Z(n1158) );
NOR2_X1 U835 ( .A1(n1162), .A2(n1150), .ZN(n1161) );
NAND2_X1 U836 ( .A1(KEYINPUT26), .A2(G140), .ZN(n1160) );
NOR2_X1 U837 ( .A1(n1122), .A2(n1163), .ZN(G51) );
XOR2_X1 U838 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U839 ( .A(n1166), .B(n1167), .Z(n1165) );
XNOR2_X1 U840 ( .A(n1168), .B(n1169), .ZN(n1167) );
NOR2_X1 U841 ( .A1(n1079), .A2(n1150), .ZN(n1166) );
NAND2_X1 U842 ( .A1(G902), .A2(n1026), .ZN(n1150) );
NAND2_X1 U843 ( .A1(n1119), .A2(n1106), .ZN(n1026) );
AND4_X1 U844 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1106) );
NOR4_X1 U845 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1173) );
NOR2_X1 U846 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NOR2_X1 U847 ( .A1(n1180), .A2(n1181), .ZN(n1172) );
NAND2_X1 U848 ( .A1(n1034), .A2(n1182), .ZN(n1170) );
NAND2_X1 U849 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NAND4_X1 U850 ( .A1(n1066), .A2(n1179), .A3(n1059), .A4(n1185), .ZN(n1184) );
NOR2_X1 U851 ( .A1(n1047), .A2(n1186), .ZN(n1185) );
INV_X1 U852 ( .A(n1187), .ZN(n1047) );
INV_X1 U853 ( .A(KEYINPUT55), .ZN(n1179) );
XOR2_X1 U854 ( .A(KEYINPUT3), .B(n1188), .Z(n1183) );
AND4_X1 U855 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1119) );
AND4_X1 U856 ( .A1(n1141), .A2(n1021), .A3(n1193), .A4(n1194), .ZN(n1192) );
NAND3_X1 U857 ( .A1(n1049), .A2(n1195), .A3(n1060), .ZN(n1021) );
NAND3_X1 U858 ( .A1(n1049), .A2(n1195), .A3(n1059), .ZN(n1141) );
NOR2_X1 U859 ( .A1(n1196), .A2(n1197), .ZN(n1191) );
NOR4_X1 U860 ( .A1(n1198), .A2(n1199), .A3(KEYINPUT58), .A4(n1051), .ZN(n1197) );
NAND3_X1 U861 ( .A1(n1032), .A2(n1043), .A3(n1200), .ZN(n1198) );
NOR2_X1 U862 ( .A1(n1201), .A2(n1202), .ZN(n1196) );
XNOR2_X1 U863 ( .A(KEYINPUT38), .B(n1031), .ZN(n1202) );
NAND2_X1 U864 ( .A1(n1203), .A2(n1204), .ZN(n1189) );
NAND2_X1 U865 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NAND2_X1 U866 ( .A1(KEYINPUT58), .A2(n1032), .ZN(n1206) );
XNOR2_X1 U867 ( .A(n1187), .B(KEYINPUT16), .ZN(n1205) );
XOR2_X1 U868 ( .A(n1207), .B(n1149), .Z(n1164) );
NAND2_X1 U869 ( .A1(KEYINPUT27), .A2(n1208), .ZN(n1207) );
NOR2_X1 U870 ( .A1(n1036), .A2(G952), .ZN(n1122) );
XOR2_X1 U871 ( .A(G146), .B(n1176), .Z(G48) );
AND4_X1 U872 ( .A1(n1209), .A2(n1059), .A3(n1210), .A4(n1066), .ZN(n1176) );
XOR2_X1 U873 ( .A(G143), .B(n1175), .Z(G45) );
AND4_X1 U874 ( .A1(n1211), .A2(n1210), .A3(n1075), .A4(n1212), .ZN(n1175) );
XOR2_X1 U875 ( .A(n1213), .B(n1214), .Z(G42) );
NAND2_X1 U876 ( .A1(KEYINPUT29), .A2(G140), .ZN(n1214) );
NAND2_X1 U877 ( .A1(n1188), .A2(n1034), .ZN(n1213) );
AND2_X1 U878 ( .A1(n1215), .A2(n1066), .ZN(n1188) );
XNOR2_X1 U879 ( .A(G137), .B(n1171), .ZN(G39) );
NAND4_X1 U880 ( .A1(n1034), .A2(n1209), .A3(n1043), .A4(n1066), .ZN(n1171) );
XOR2_X1 U881 ( .A(G134), .B(n1174), .Z(G36) );
AND3_X1 U882 ( .A1(n1034), .A2(n1060), .A3(n1211), .ZN(n1174) );
XNOR2_X1 U883 ( .A(G131), .B(n1178), .ZN(G33) );
NAND3_X1 U884 ( .A1(n1034), .A2(n1059), .A3(n1211), .ZN(n1178) );
AND3_X1 U885 ( .A1(n1066), .A2(n1186), .A3(n1187), .ZN(n1211) );
XOR2_X1 U886 ( .A(n1216), .B(KEYINPUT54), .Z(n1066) );
AND2_X1 U887 ( .A1(n1054), .A2(n1217), .ZN(n1034) );
XNOR2_X1 U888 ( .A(n1181), .B(n1218), .ZN(G30) );
XOR2_X1 U889 ( .A(KEYINPUT61), .B(G128), .Z(n1218) );
AND4_X1 U890 ( .A1(n1209), .A2(n1060), .A3(n1216), .A4(n1210), .ZN(n1181) );
AND3_X1 U891 ( .A1(n1074), .A2(n1186), .A3(n1219), .ZN(n1209) );
XNOR2_X1 U892 ( .A(G101), .B(n1220), .ZN(G3) );
NAND2_X1 U893 ( .A1(n1203), .A2(n1187), .ZN(n1220) );
XNOR2_X1 U894 ( .A(n1168), .B(n1180), .ZN(G27) );
AND3_X1 U895 ( .A1(n1041), .A2(n1210), .A3(n1215), .ZN(n1180) );
AND3_X1 U896 ( .A1(n1059), .A2(n1186), .A3(n1032), .ZN(n1215) );
NAND2_X1 U897 ( .A1(n1067), .A2(n1221), .ZN(n1186) );
NAND4_X1 U898 ( .A1(G902), .A2(G953), .A3(n1222), .A4(n1223), .ZN(n1221) );
INV_X1 U899 ( .A(G900), .ZN(n1223) );
INV_X1 U900 ( .A(n1030), .ZN(n1041) );
XNOR2_X1 U901 ( .A(G122), .B(n1190), .ZN(G24) );
NAND4_X1 U902 ( .A1(n1224), .A2(n1049), .A3(n1075), .A4(n1212), .ZN(n1190) );
NOR2_X1 U903 ( .A1(n1074), .A2(n1219), .ZN(n1049) );
XOR2_X1 U904 ( .A(G119), .B(n1225), .Z(G21) );
NOR2_X1 U905 ( .A1(n1031), .A2(n1201), .ZN(n1225) );
NAND3_X1 U906 ( .A1(n1224), .A2(n1074), .A3(n1219), .ZN(n1201) );
INV_X1 U907 ( .A(n1043), .ZN(n1031) );
NAND2_X1 U908 ( .A1(n1226), .A2(n1227), .ZN(G18) );
NAND2_X1 U909 ( .A1(G116), .A2(n1194), .ZN(n1227) );
XOR2_X1 U910 ( .A(KEYINPUT56), .B(n1228), .Z(n1226) );
NOR2_X1 U911 ( .A1(G116), .A2(n1194), .ZN(n1228) );
NAND3_X1 U912 ( .A1(n1187), .A2(n1060), .A3(n1224), .ZN(n1194) );
NOR2_X1 U913 ( .A1(n1212), .A2(n1229), .ZN(n1060) );
INV_X1 U914 ( .A(n1075), .ZN(n1229) );
XNOR2_X1 U915 ( .A(G113), .B(n1193), .ZN(G15) );
NAND3_X1 U916 ( .A1(n1187), .A2(n1059), .A3(n1224), .ZN(n1193) );
NOR3_X1 U917 ( .A1(n1051), .A2(n1200), .A3(n1030), .ZN(n1224) );
NAND2_X1 U918 ( .A1(n1065), .A2(n1230), .ZN(n1030) );
XOR2_X1 U919 ( .A(n1231), .B(KEYINPUT41), .Z(n1065) );
NOR2_X1 U920 ( .A1(n1075), .A2(n1232), .ZN(n1059) );
NOR2_X1 U921 ( .A1(n1219), .A2(n1233), .ZN(n1187) );
INV_X1 U922 ( .A(n1074), .ZN(n1233) );
INV_X1 U923 ( .A(n1234), .ZN(n1219) );
XNOR2_X1 U924 ( .A(G110), .B(n1235), .ZN(G12) );
NAND2_X1 U925 ( .A1(n1203), .A2(n1032), .ZN(n1235) );
NOR2_X1 U926 ( .A1(n1234), .A2(n1074), .ZN(n1032) );
XNOR2_X1 U927 ( .A(n1236), .B(G472), .ZN(n1074) );
NAND2_X1 U928 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XOR2_X1 U929 ( .A(n1239), .B(n1240), .Z(n1237) );
XOR2_X1 U930 ( .A(n1147), .B(G101), .Z(n1240) );
NAND2_X1 U931 ( .A1(G210), .A2(n1241), .ZN(n1147) );
NAND2_X1 U932 ( .A1(KEYINPUT17), .A2(n1242), .ZN(n1239) );
XNOR2_X1 U933 ( .A(n1243), .B(n1152), .ZN(n1242) );
INV_X1 U934 ( .A(n1244), .ZN(n1152) );
NOR2_X1 U935 ( .A1(n1245), .A2(n1246), .ZN(n1243) );
XOR2_X1 U936 ( .A(n1247), .B(KEYINPUT63), .Z(n1246) );
NAND2_X1 U937 ( .A1(n1248), .A2(n1149), .ZN(n1247) );
NOR2_X1 U938 ( .A1(n1248), .A2(n1149), .ZN(n1245) );
XOR2_X1 U939 ( .A(n1249), .B(KEYINPUT11), .Z(n1248) );
XOR2_X1 U940 ( .A(n1085), .B(n1250), .Z(n1234) );
NOR2_X1 U941 ( .A1(n1083), .A2(KEYINPUT22), .ZN(n1250) );
AND2_X1 U942 ( .A1(G217), .A2(n1251), .ZN(n1083) );
NOR2_X1 U943 ( .A1(n1125), .A2(G902), .ZN(n1085) );
XNOR2_X1 U944 ( .A(n1252), .B(n1253), .ZN(n1125) );
XOR2_X1 U945 ( .A(G119), .B(G110), .Z(n1253) );
XOR2_X1 U946 ( .A(n1254), .B(n1255), .Z(n1252) );
NOR3_X1 U947 ( .A1(n1256), .A2(G953), .A3(n1257), .ZN(n1255) );
INV_X1 U948 ( .A(G221), .ZN(n1257) );
XOR2_X1 U949 ( .A(KEYINPUT43), .B(G234), .Z(n1256) );
XOR2_X1 U950 ( .A(n1258), .B(n1259), .Z(n1254) );
XNOR2_X1 U951 ( .A(G137), .B(n1260), .ZN(n1259) );
XNOR2_X1 U952 ( .A(KEYINPUT40), .B(KEYINPUT39), .ZN(n1260) );
XNOR2_X1 U953 ( .A(n1261), .B(n1262), .ZN(n1258) );
INV_X1 U954 ( .A(n1263), .ZN(n1262) );
XNOR2_X1 U955 ( .A(n1264), .B(n1168), .ZN(n1261) );
AND2_X1 U956 ( .A1(n1043), .A2(n1195), .ZN(n1203) );
NOR3_X1 U957 ( .A1(n1051), .A2(n1200), .A3(n1199), .ZN(n1195) );
INV_X1 U958 ( .A(n1216), .ZN(n1199) );
NOR2_X1 U959 ( .A1(n1231), .A2(n1064), .ZN(n1216) );
INV_X1 U960 ( .A(n1230), .ZN(n1064) );
NAND2_X1 U961 ( .A1(G221), .A2(n1251), .ZN(n1230) );
NAND2_X1 U962 ( .A1(G234), .A2(n1238), .ZN(n1251) );
NAND3_X1 U963 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1231) );
OR2_X1 U964 ( .A1(n1162), .A2(n1268), .ZN(n1267) );
NAND3_X1 U965 ( .A1(n1268), .A2(n1162), .A3(KEYINPUT9), .ZN(n1266) );
INV_X1 U966 ( .A(G469), .ZN(n1162) );
NOR2_X1 U967 ( .A1(n1269), .A2(KEYINPUT47), .ZN(n1268) );
INV_X1 U968 ( .A(n1077), .ZN(n1269) );
OR2_X1 U969 ( .A1(n1077), .A2(KEYINPUT9), .ZN(n1265) );
NAND2_X1 U970 ( .A1(n1270), .A2(n1238), .ZN(n1077) );
XNOR2_X1 U971 ( .A(n1159), .B(n1271), .ZN(n1270) );
NOR3_X1 U972 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n1271) );
NOR2_X1 U973 ( .A1(KEYINPUT13), .A2(n1156), .ZN(n1274) );
NOR3_X1 U974 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1273) );
INV_X1 U975 ( .A(KEYINPUT13), .ZN(n1275) );
AND2_X1 U976 ( .A1(n1277), .A2(n1276), .ZN(n1272) );
XNOR2_X1 U977 ( .A(G110), .B(G140), .ZN(n1276) );
NAND2_X1 U978 ( .A1(KEYINPUT45), .A2(n1156), .ZN(n1277) );
AND2_X1 U979 ( .A1(G227), .A2(n1278), .ZN(n1156) );
XNOR2_X1 U980 ( .A(KEYINPUT53), .B(n1036), .ZN(n1278) );
XOR2_X1 U981 ( .A(n1279), .B(n1098), .Z(n1159) );
XOR2_X1 U982 ( .A(n1264), .B(n1280), .Z(n1098) );
XOR2_X1 U983 ( .A(KEYINPUT62), .B(G143), .Z(n1280) );
XOR2_X1 U984 ( .A(n1151), .B(n1281), .Z(n1279) );
XOR2_X1 U985 ( .A(n1249), .B(G101), .Z(n1151) );
NAND2_X1 U986 ( .A1(n1282), .A2(n1283), .ZN(n1249) );
OR2_X1 U987 ( .A1(n1104), .A2(G131), .ZN(n1283) );
XOR2_X1 U988 ( .A(n1100), .B(KEYINPUT46), .Z(n1282) );
NAND2_X1 U989 ( .A1(n1104), .A2(G131), .ZN(n1100) );
XNOR2_X1 U990 ( .A(G134), .B(n1284), .ZN(n1104) );
XOR2_X1 U991 ( .A(KEYINPUT8), .B(G137), .Z(n1284) );
AND2_X1 U992 ( .A1(n1067), .A2(n1285), .ZN(n1200) );
NAND4_X1 U993 ( .A1(G902), .A2(G953), .A3(n1222), .A4(n1113), .ZN(n1285) );
INV_X1 U994 ( .A(G898), .ZN(n1113) );
NAND3_X1 U995 ( .A1(n1222), .A2(n1036), .A3(G952), .ZN(n1067) );
NAND2_X1 U996 ( .A1(G237), .A2(G234), .ZN(n1222) );
INV_X1 U997 ( .A(n1210), .ZN(n1051) );
NOR2_X1 U998 ( .A1(n1054), .A2(n1053), .ZN(n1210) );
INV_X1 U999 ( .A(n1217), .ZN(n1053) );
NAND2_X1 U1000 ( .A1(G214), .A2(n1286), .ZN(n1217) );
XOR2_X1 U1001 ( .A(n1287), .B(n1079), .Z(n1054) );
NAND2_X1 U1002 ( .A1(G210), .A2(n1286), .ZN(n1079) );
NAND2_X1 U1003 ( .A1(n1288), .A2(n1238), .ZN(n1286) );
INV_X1 U1004 ( .A(G237), .ZN(n1288) );
XNOR2_X1 U1005 ( .A(KEYINPUT21), .B(n1289), .ZN(n1287) );
NOR2_X1 U1006 ( .A1(KEYINPUT33), .A2(n1080), .ZN(n1289) );
AND2_X1 U1007 ( .A1(n1290), .A2(n1238), .ZN(n1080) );
XNOR2_X1 U1008 ( .A(n1291), .B(n1208), .ZN(n1290) );
XOR2_X1 U1009 ( .A(n1116), .B(n1292), .Z(n1208) );
XOR2_X1 U1010 ( .A(KEYINPUT0), .B(n1118), .Z(n1292) );
XNOR2_X1 U1011 ( .A(G110), .B(n1293), .ZN(n1118) );
XNOR2_X1 U1012 ( .A(n1244), .B(n1294), .ZN(n1116) );
XOR2_X1 U1013 ( .A(n1295), .B(n1281), .Z(n1294) );
XNOR2_X1 U1014 ( .A(n1296), .B(n1297), .ZN(n1281) );
XNOR2_X1 U1015 ( .A(G107), .B(KEYINPUT59), .ZN(n1296) );
NOR2_X1 U1016 ( .A1(G101), .A2(KEYINPUT50), .ZN(n1295) );
XOR2_X1 U1017 ( .A(G113), .B(n1298), .Z(n1244) );
XOR2_X1 U1018 ( .A(G119), .B(G116), .Z(n1298) );
NOR2_X1 U1019 ( .A1(KEYINPUT51), .A2(n1299), .ZN(n1291) );
XNOR2_X1 U1020 ( .A(n1169), .B(n1300), .ZN(n1299) );
NAND2_X1 U1021 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U1022 ( .A1(G125), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1023 ( .A(n1304), .B(KEYINPUT25), .Z(n1301) );
OR2_X1 U1024 ( .A1(n1303), .A2(G125), .ZN(n1304) );
XOR2_X1 U1025 ( .A(n1149), .B(KEYINPUT52), .Z(n1303) );
XNOR2_X1 U1026 ( .A(n1264), .B(n1305), .ZN(n1149) );
NOR2_X1 U1027 ( .A1(KEYINPUT2), .A2(n1306), .ZN(n1305) );
XOR2_X1 U1028 ( .A(KEYINPUT10), .B(G143), .Z(n1306) );
XNOR2_X1 U1029 ( .A(G128), .B(n1307), .ZN(n1264) );
AND2_X1 U1030 ( .A1(G224), .A2(n1036), .ZN(n1169) );
NOR2_X1 U1031 ( .A1(n1075), .A2(n1212), .ZN(n1043) );
INV_X1 U1032 ( .A(n1232), .ZN(n1212) );
NOR2_X1 U1033 ( .A1(n1308), .A2(n1081), .ZN(n1232) );
NOR2_X1 U1034 ( .A1(n1082), .A2(G475), .ZN(n1081) );
AND2_X1 U1035 ( .A1(n1309), .A2(G475), .ZN(n1308) );
XOR2_X1 U1036 ( .A(n1082), .B(KEYINPUT18), .Z(n1309) );
NAND2_X1 U1037 ( .A1(n1139), .A2(n1238), .ZN(n1082) );
INV_X1 U1038 ( .A(G902), .ZN(n1238) );
XNOR2_X1 U1039 ( .A(n1310), .B(n1311), .ZN(n1139) );
XNOR2_X1 U1040 ( .A(n1263), .B(n1312), .ZN(n1311) );
XNOR2_X1 U1041 ( .A(n1307), .B(n1297), .ZN(n1312) );
XOR2_X1 U1042 ( .A(G104), .B(KEYINPUT37), .Z(n1297) );
XOR2_X1 U1043 ( .A(G146), .B(KEYINPUT6), .Z(n1307) );
XOR2_X1 U1044 ( .A(G140), .B(KEYINPUT14), .Z(n1263) );
XOR2_X1 U1045 ( .A(n1313), .B(n1314), .Z(n1310) );
XOR2_X1 U1046 ( .A(n1315), .B(n1316), .Z(n1314) );
NAND2_X1 U1047 ( .A1(KEYINPUT44), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1048 ( .A(KEYINPUT1), .B(n1168), .ZN(n1317) );
INV_X1 U1049 ( .A(G125), .ZN(n1168) );
NAND3_X1 U1050 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1315) );
NAND2_X1 U1051 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NAND2_X1 U1052 ( .A1(n1323), .A2(KEYINPUT20), .ZN(n1322) );
XNOR2_X1 U1053 ( .A(G131), .B(KEYINPUT7), .ZN(n1323) );
INV_X1 U1054 ( .A(n1324), .ZN(n1321) );
NAND3_X1 U1055 ( .A1(KEYINPUT20), .A2(n1324), .A3(n1325), .ZN(n1319) );
XNOR2_X1 U1056 ( .A(n1326), .B(G143), .ZN(n1324) );
NAND2_X1 U1057 ( .A1(G214), .A2(n1241), .ZN(n1326) );
NOR2_X1 U1058 ( .A1(G953), .A2(G237), .ZN(n1241) );
OR2_X1 U1059 ( .A1(n1325), .A2(KEYINPUT20), .ZN(n1318) );
INV_X1 U1060 ( .A(G131), .ZN(n1325) );
XNOR2_X1 U1061 ( .A(G113), .B(G122), .ZN(n1313) );
XOR2_X1 U1062 ( .A(G478), .B(n1327), .Z(n1075) );
NOR2_X1 U1063 ( .A1(G902), .A2(n1136), .ZN(n1327) );
INV_X1 U1064 ( .A(n1130), .ZN(n1136) );
XNOR2_X1 U1065 ( .A(n1328), .B(n1329), .ZN(n1130) );
NOR2_X1 U1066 ( .A1(KEYINPUT49), .A2(n1330), .ZN(n1329) );
XOR2_X1 U1067 ( .A(n1331), .B(n1332), .Z(n1330) );
XNOR2_X1 U1068 ( .A(n1333), .B(n1334), .ZN(n1332) );
XNOR2_X1 U1069 ( .A(n1293), .B(G116), .ZN(n1334) );
INV_X1 U1070 ( .A(G122), .ZN(n1293) );
INV_X1 U1071 ( .A(G107), .ZN(n1333) );
XOR2_X1 U1072 ( .A(n1335), .B(n1336), .Z(n1331) );
XOR2_X1 U1073 ( .A(G134), .B(G128), .Z(n1336) );
XOR2_X1 U1074 ( .A(KEYINPUT60), .B(G143), .Z(n1335) );
NAND3_X1 U1075 ( .A1(G217), .A2(n1036), .A3(G234), .ZN(n1328) );
INV_X1 U1076 ( .A(G953), .ZN(n1036) );
endmodule


