//Key = 0010001110111111001011010111011101010100011011101010001011110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;

XOR2_X1 U734 ( .A(n1008), .B(n1009), .Z(G9) );
XNOR2_X1 U735 ( .A(KEYINPUT10), .B(n1010), .ZN(n1009) );
NOR2_X1 U736 ( .A1(n1011), .A2(n1012), .ZN(G75) );
NOR4_X1 U737 ( .A1(G953), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1012) );
XOR2_X1 U738 ( .A(KEYINPUT15), .B(n1016), .Z(n1015) );
NOR4_X1 U739 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
NOR3_X1 U740 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
INV_X1 U741 ( .A(n1024), .ZN(n1023) );
NOR2_X1 U742 ( .A1(n1025), .A2(n1026), .ZN(n1022) );
NOR2_X1 U743 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
AND2_X1 U744 ( .A1(n1029), .A2(n1030), .ZN(n1025) );
NOR4_X1 U745 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1028), .ZN(n1019) );
XNOR2_X1 U746 ( .A(n1034), .B(KEYINPUT24), .ZN(n1033) );
INV_X1 U747 ( .A(n1035), .ZN(n1032) );
NAND2_X1 U748 ( .A1(n1036), .A2(n1029), .ZN(n1031) );
NOR4_X1 U749 ( .A1(n1028), .A2(n1037), .A3(n1038), .A4(n1021), .ZN(n1018) );
INV_X1 U750 ( .A(n1039), .ZN(n1021) );
INV_X1 U751 ( .A(n1040), .ZN(n1028) );
NAND3_X1 U752 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1017) );
NAND2_X1 U753 ( .A1(n1024), .A2(n1044), .ZN(n1042) );
NAND2_X1 U754 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND3_X1 U755 ( .A1(n1047), .A2(n1029), .A3(n1039), .ZN(n1046) );
NOR2_X1 U756 ( .A1(n1048), .A2(n1049), .ZN(n1039) );
NAND3_X1 U757 ( .A1(n1040), .A2(n1050), .A3(n1036), .ZN(n1045) );
INV_X1 U758 ( .A(n1048), .ZN(n1036) );
NAND2_X1 U759 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND4_X1 U760 ( .A1(n1053), .A2(n1034), .A3(G214), .A4(n1054), .ZN(n1052) );
NAND2_X1 U761 ( .A1(n1029), .A2(n1055), .ZN(n1051) );
NAND2_X1 U762 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U763 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
INV_X1 U764 ( .A(G952), .ZN(n1014) );
NOR3_X1 U765 ( .A1(n1060), .A2(G953), .A3(n1013), .ZN(n1011) );
AND4_X1 U766 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1013) );
NOR4_X1 U767 ( .A1(n1065), .A2(n1066), .A3(n1037), .A4(n1067), .ZN(n1064) );
XOR2_X1 U768 ( .A(n1068), .B(n1069), .Z(n1066) );
XNOR2_X1 U769 ( .A(KEYINPUT58), .B(n1070), .ZN(n1069) );
XNOR2_X1 U770 ( .A(n1071), .B(n1072), .ZN(n1065) );
NAND2_X1 U771 ( .A1(KEYINPUT50), .A2(n1073), .ZN(n1071) );
NOR3_X1 U772 ( .A1(n1074), .A2(n1075), .A3(n1059), .ZN(n1063) );
NAND2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1061) );
XNOR2_X1 U774 ( .A(KEYINPUT0), .B(n1078), .ZN(n1076) );
XNOR2_X1 U775 ( .A(G952), .B(KEYINPUT23), .ZN(n1060) );
NAND2_X1 U776 ( .A1(n1079), .A2(n1080), .ZN(G72) );
NAND2_X1 U777 ( .A1(n1081), .A2(G953), .ZN(n1080) );
XNOR2_X1 U778 ( .A(n1082), .B(n1083), .ZN(n1081) );
NOR2_X1 U779 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U780 ( .A1(n1086), .A2(n1087), .ZN(n1079) );
NAND2_X1 U781 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NAND2_X1 U782 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U783 ( .A1(n1082), .A2(n1041), .ZN(n1088) );
XNOR2_X1 U784 ( .A(n1090), .B(KEYINPUT49), .ZN(n1082) );
NAND2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NAND2_X1 U786 ( .A1(G953), .A2(n1085), .ZN(n1093) );
XOR2_X1 U787 ( .A(n1094), .B(n1095), .Z(n1092) );
XOR2_X1 U788 ( .A(n1096), .B(n1097), .Z(n1095) );
XNOR2_X1 U789 ( .A(n1098), .B(n1099), .ZN(n1094) );
XNOR2_X1 U790 ( .A(n1100), .B(G134), .ZN(n1099) );
XOR2_X1 U791 ( .A(n1101), .B(n1102), .Z(G69) );
XOR2_X1 U792 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR3_X1 U793 ( .A1(n1043), .A2(KEYINPUT32), .A3(G953), .ZN(n1104) );
NOR2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
XOR2_X1 U795 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U796 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U797 ( .A1(KEYINPUT4), .A2(n1111), .ZN(n1109) );
XNOR2_X1 U798 ( .A(G113), .B(n1112), .ZN(n1111) );
NOR2_X1 U799 ( .A1(G898), .A2(n1113), .ZN(n1105) );
XNOR2_X1 U800 ( .A(G953), .B(KEYINPUT60), .ZN(n1113) );
NOR2_X1 U801 ( .A1(n1114), .A2(n1087), .ZN(n1101) );
NOR2_X1 U802 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U803 ( .A1(n1117), .A2(n1118), .ZN(G66) );
NOR2_X1 U804 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XOR2_X1 U805 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U806 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U807 ( .A1(KEYINPUT36), .A2(n1125), .ZN(n1121) );
AND2_X1 U808 ( .A1(n1125), .A2(KEYINPUT36), .ZN(n1119) );
NOR2_X1 U809 ( .A1(n1117), .A2(n1126), .ZN(G63) );
XNOR2_X1 U810 ( .A(n1127), .B(n1128), .ZN(n1126) );
NOR2_X1 U811 ( .A1(n1078), .A2(n1124), .ZN(n1128) );
INV_X1 U812 ( .A(G478), .ZN(n1078) );
NOR2_X1 U813 ( .A1(n1117), .A2(n1129), .ZN(G60) );
XOR2_X1 U814 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U815 ( .A1(n1132), .A2(n1124), .ZN(n1131) );
NAND2_X1 U816 ( .A1(KEYINPUT41), .A2(n1133), .ZN(n1130) );
XNOR2_X1 U817 ( .A(G104), .B(n1134), .ZN(G6) );
NOR2_X1 U818 ( .A1(n1117), .A2(n1135), .ZN(G57) );
XOR2_X1 U819 ( .A(n1136), .B(n1137), .Z(n1135) );
XNOR2_X1 U820 ( .A(n1138), .B(n1139), .ZN(n1137) );
XOR2_X1 U821 ( .A(n1140), .B(n1141), .Z(n1136) );
NOR2_X1 U822 ( .A1(n1142), .A2(KEYINPUT1), .ZN(n1141) );
XOR2_X1 U823 ( .A(n1143), .B(n1144), .Z(n1140) );
NOR2_X1 U824 ( .A1(n1072), .A2(n1124), .ZN(n1144) );
INV_X1 U825 ( .A(G472), .ZN(n1072) );
NOR2_X1 U826 ( .A1(n1117), .A2(n1145), .ZN(G54) );
XOR2_X1 U827 ( .A(n1146), .B(n1147), .Z(n1145) );
XNOR2_X1 U828 ( .A(n1148), .B(n1149), .ZN(n1147) );
XOR2_X1 U829 ( .A(n1150), .B(n1151), .Z(n1146) );
NOR2_X1 U830 ( .A1(n1070), .A2(n1124), .ZN(n1151) );
INV_X1 U831 ( .A(G469), .ZN(n1070) );
NOR3_X1 U832 ( .A1(n1084), .A2(KEYINPUT5), .A3(G953), .ZN(n1150) );
NOR2_X1 U833 ( .A1(n1087), .A2(G952), .ZN(n1117) );
NOR2_X1 U834 ( .A1(n1152), .A2(n1153), .ZN(G51) );
XOR2_X1 U835 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U836 ( .A1(n1156), .A2(n1124), .ZN(n1155) );
NAND2_X1 U837 ( .A1(G902), .A2(n1157), .ZN(n1124) );
NAND2_X1 U838 ( .A1(n1043), .A2(n1041), .ZN(n1157) );
INV_X1 U839 ( .A(n1091), .ZN(n1041) );
NAND4_X1 U840 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1091) );
NOR4_X1 U841 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1161) );
AND2_X1 U842 ( .A1(n1166), .A2(n1167), .ZN(n1160) );
NAND2_X1 U843 ( .A1(n1168), .A2(n1169), .ZN(n1158) );
XOR2_X1 U844 ( .A(n1170), .B(KEYINPUT12), .Z(n1168) );
AND4_X1 U845 ( .A1(n1134), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1043) );
AND4_X1 U846 ( .A1(n1008), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1173) );
NAND3_X1 U847 ( .A1(n1040), .A2(n1177), .A3(n1035), .ZN(n1008) );
AND2_X1 U848 ( .A1(n1178), .A2(n1179), .ZN(n1172) );
NAND4_X1 U849 ( .A1(n1180), .A2(n1030), .A3(n1035), .A4(n1181), .ZN(n1171) );
XNOR2_X1 U850 ( .A(n1034), .B(KEYINPUT59), .ZN(n1180) );
NAND3_X1 U851 ( .A1(n1040), .A2(n1177), .A3(n1182), .ZN(n1134) );
NOR2_X1 U852 ( .A1(G952), .A2(n1183), .ZN(n1152) );
XNOR2_X1 U853 ( .A(G953), .B(KEYINPUT3), .ZN(n1183) );
XOR2_X1 U854 ( .A(n1159), .B(n1184), .Z(G48) );
NOR2_X1 U855 ( .A1(KEYINPUT51), .A2(n1185), .ZN(n1184) );
XNOR2_X1 U856 ( .A(G146), .B(KEYINPUT14), .ZN(n1185) );
NAND3_X1 U857 ( .A1(n1182), .A2(n1169), .A3(n1186), .ZN(n1159) );
XNOR2_X1 U858 ( .A(n1187), .B(n1188), .ZN(G45) );
NOR2_X1 U859 ( .A1(n1027), .A2(n1170), .ZN(n1188) );
NAND3_X1 U860 ( .A1(n1030), .A2(n1189), .A3(n1190), .ZN(n1170) );
AND3_X1 U861 ( .A1(n1067), .A2(n1191), .A3(n1192), .ZN(n1190) );
INV_X1 U862 ( .A(n1169), .ZN(n1027) );
XOR2_X1 U863 ( .A(n1166), .B(n1193), .Z(G42) );
NOR2_X1 U864 ( .A1(KEYINPUT9), .A2(n1194), .ZN(n1193) );
XNOR2_X1 U865 ( .A(G140), .B(KEYINPUT11), .ZN(n1194) );
NAND3_X1 U866 ( .A1(n1182), .A2(n1047), .A3(n1195), .ZN(n1166) );
XOR2_X1 U867 ( .A(G137), .B(n1165), .Z(G39) );
AND3_X1 U868 ( .A1(n1024), .A2(n1029), .A3(n1186), .ZN(n1165) );
XOR2_X1 U869 ( .A(n1164), .B(n1196), .Z(G36) );
NOR2_X1 U870 ( .A1(KEYINPUT40), .A2(n1197), .ZN(n1196) );
AND3_X1 U871 ( .A1(n1030), .A2(n1035), .A3(n1195), .ZN(n1164) );
XOR2_X1 U872 ( .A(n1163), .B(n1198), .Z(G33) );
NOR2_X1 U873 ( .A1(KEYINPUT62), .A2(n1199), .ZN(n1198) );
AND3_X1 U874 ( .A1(n1182), .A2(n1030), .A3(n1195), .ZN(n1163) );
AND3_X1 U875 ( .A1(n1189), .A2(n1192), .A3(n1029), .ZN(n1195) );
INV_X1 U876 ( .A(n1037), .ZN(n1029) );
NAND2_X1 U877 ( .A1(n1053), .A2(n1200), .ZN(n1037) );
NAND2_X1 U878 ( .A1(G214), .A2(n1054), .ZN(n1200) );
XNOR2_X1 U879 ( .A(n1201), .B(n1162), .ZN(G30) );
AND3_X1 U880 ( .A1(n1035), .A2(n1169), .A3(n1186), .ZN(n1162) );
AND4_X1 U881 ( .A1(n1189), .A2(n1202), .A3(n1203), .A4(n1192), .ZN(n1186) );
XNOR2_X1 U882 ( .A(G101), .B(n1179), .ZN(G3) );
NAND3_X1 U883 ( .A1(n1024), .A2(n1177), .A3(n1030), .ZN(n1179) );
XNOR2_X1 U884 ( .A(G125), .B(n1167), .ZN(G27) );
NAND4_X1 U885 ( .A1(n1169), .A2(n1192), .A3(n1047), .A4(n1204), .ZN(n1167) );
NOR2_X1 U886 ( .A1(n1049), .A2(n1038), .ZN(n1204) );
INV_X1 U887 ( .A(n1182), .ZN(n1038) );
NAND2_X1 U888 ( .A1(n1205), .A2(n1048), .ZN(n1192) );
NAND4_X1 U889 ( .A1(G902), .A2(G953), .A3(n1206), .A4(n1085), .ZN(n1205) );
INV_X1 U890 ( .A(G900), .ZN(n1085) );
XNOR2_X1 U891 ( .A(G122), .B(n1178), .ZN(G24) );
NAND4_X1 U892 ( .A1(n1207), .A2(n1040), .A3(n1067), .A4(n1191), .ZN(n1178) );
NOR2_X1 U893 ( .A1(n1203), .A2(n1202), .ZN(n1040) );
XOR2_X1 U894 ( .A(n1176), .B(n1208), .Z(G21) );
NOR2_X1 U895 ( .A1(G119), .A2(KEYINPUT38), .ZN(n1208) );
NAND4_X1 U896 ( .A1(n1207), .A2(n1024), .A3(n1202), .A4(n1203), .ZN(n1176) );
INV_X1 U897 ( .A(n1209), .ZN(n1202) );
XNOR2_X1 U898 ( .A(G116), .B(n1210), .ZN(G18) );
NAND4_X1 U899 ( .A1(KEYINPUT46), .A2(n1030), .A3(n1207), .A4(n1035), .ZN(n1210) );
NOR2_X1 U900 ( .A1(n1067), .A2(n1211), .ZN(n1035) );
XOR2_X1 U901 ( .A(n1175), .B(n1212), .Z(G15) );
XNOR2_X1 U902 ( .A(KEYINPUT54), .B(n1213), .ZN(n1212) );
NAND3_X1 U903 ( .A1(n1030), .A2(n1207), .A3(n1182), .ZN(n1175) );
NOR2_X1 U904 ( .A1(n1191), .A2(n1214), .ZN(n1182) );
INV_X1 U905 ( .A(n1067), .ZN(n1214) );
AND2_X1 U906 ( .A1(n1034), .A2(n1181), .ZN(n1207) );
INV_X1 U907 ( .A(n1049), .ZN(n1034) );
NAND2_X1 U908 ( .A1(n1058), .A2(n1215), .ZN(n1049) );
XOR2_X1 U909 ( .A(n1216), .B(KEYINPUT44), .Z(n1058) );
NOR2_X1 U910 ( .A1(n1203), .A2(n1209), .ZN(n1030) );
XNOR2_X1 U911 ( .A(G110), .B(n1174), .ZN(G12) );
NAND3_X1 U912 ( .A1(n1047), .A2(n1177), .A3(n1024), .ZN(n1174) );
NOR2_X1 U913 ( .A1(n1191), .A2(n1067), .ZN(n1024) );
XOR2_X1 U914 ( .A(n1217), .B(n1132), .Z(n1067) );
INV_X1 U915 ( .A(G475), .ZN(n1132) );
NAND2_X1 U916 ( .A1(n1133), .A2(n1218), .ZN(n1217) );
XOR2_X1 U917 ( .A(n1219), .B(n1220), .Z(n1133) );
XOR2_X1 U918 ( .A(n1221), .B(n1222), .Z(n1220) );
XNOR2_X1 U919 ( .A(n1223), .B(n1098), .ZN(n1222) );
INV_X1 U920 ( .A(G125), .ZN(n1098) );
NAND2_X1 U921 ( .A1(KEYINPUT7), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U922 ( .A(KEYINPUT25), .B(n1187), .ZN(n1224) );
XNOR2_X1 U923 ( .A(G131), .B(G146), .ZN(n1221) );
XOR2_X1 U924 ( .A(n1225), .B(n1226), .Z(n1219) );
XOR2_X1 U925 ( .A(n1227), .B(n1228), .Z(n1225) );
AND2_X1 U926 ( .A1(n1229), .A2(G214), .ZN(n1228) );
NAND2_X1 U927 ( .A1(n1230), .A2(KEYINPUT45), .ZN(n1227) );
XOR2_X1 U928 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U929 ( .A(KEYINPUT30), .B(G122), .Z(n1232) );
XNOR2_X1 U930 ( .A(G104), .B(G113), .ZN(n1231) );
INV_X1 U931 ( .A(n1211), .ZN(n1191) );
NOR2_X1 U932 ( .A1(n1233), .A2(n1075), .ZN(n1211) );
NOR2_X1 U933 ( .A1(n1077), .A2(G478), .ZN(n1075) );
AND2_X1 U934 ( .A1(G478), .A2(n1077), .ZN(n1233) );
NAND2_X1 U935 ( .A1(n1127), .A2(n1218), .ZN(n1077) );
XNOR2_X1 U936 ( .A(n1234), .B(n1235), .ZN(n1127) );
XOR2_X1 U937 ( .A(n1236), .B(n1237), .Z(n1235) );
XNOR2_X1 U938 ( .A(n1010), .B(n1238), .ZN(n1237) );
NOR2_X1 U939 ( .A1(KEYINPUT17), .A2(n1239), .ZN(n1238) );
XNOR2_X1 U940 ( .A(n1240), .B(n1197), .ZN(n1239) );
NAND3_X1 U941 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1240) );
NAND2_X1 U942 ( .A1(G143), .A2(n1201), .ZN(n1243) );
NAND2_X1 U943 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
INV_X1 U944 ( .A(KEYINPUT6), .ZN(n1245) );
NAND2_X1 U945 ( .A1(n1246), .A2(n1187), .ZN(n1244) );
XNOR2_X1 U946 ( .A(KEYINPUT27), .B(G128), .ZN(n1246) );
NAND2_X1 U947 ( .A1(KEYINPUT6), .A2(n1247), .ZN(n1241) );
NAND2_X1 U948 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
OR2_X1 U949 ( .A1(G128), .A2(KEYINPUT27), .ZN(n1249) );
NAND3_X1 U950 ( .A1(G128), .A2(n1187), .A3(KEYINPUT27), .ZN(n1248) );
AND3_X1 U951 ( .A1(G234), .A2(n1087), .A3(G217), .ZN(n1236) );
XNOR2_X1 U952 ( .A(G116), .B(n1250), .ZN(n1234) );
XOR2_X1 U953 ( .A(KEYINPUT56), .B(G122), .Z(n1250) );
AND2_X1 U954 ( .A1(n1181), .A2(n1189), .ZN(n1177) );
INV_X1 U955 ( .A(n1056), .ZN(n1189) );
NAND2_X1 U956 ( .A1(n1215), .A2(n1216), .ZN(n1056) );
NAND2_X1 U957 ( .A1(n1251), .A2(n1252), .ZN(n1216) );
NAND2_X1 U958 ( .A1(G469), .A2(n1068), .ZN(n1252) );
XOR2_X1 U959 ( .A(KEYINPUT20), .B(n1253), .Z(n1251) );
NOR2_X1 U960 ( .A1(G469), .A2(n1068), .ZN(n1253) );
NAND2_X1 U961 ( .A1(n1254), .A2(n1218), .ZN(n1068) );
XOR2_X1 U962 ( .A(n1149), .B(n1255), .Z(n1254) );
XNOR2_X1 U963 ( .A(n1084), .B(n1148), .ZN(n1255) );
XNOR2_X1 U964 ( .A(G110), .B(n1100), .ZN(n1148) );
INV_X1 U965 ( .A(G140), .ZN(n1100) );
INV_X1 U966 ( .A(G227), .ZN(n1084) );
XOR2_X1 U967 ( .A(n1256), .B(n1257), .Z(n1149) );
XOR2_X1 U968 ( .A(n1139), .B(n1258), .Z(n1257) );
XNOR2_X1 U969 ( .A(n1010), .B(G104), .ZN(n1258) );
XOR2_X1 U970 ( .A(n1259), .B(n1096), .Z(n1256) );
XNOR2_X1 U971 ( .A(n1187), .B(n1260), .ZN(n1096) );
XOR2_X1 U972 ( .A(n1059), .B(KEYINPUT33), .Z(n1215) );
AND2_X1 U973 ( .A1(G221), .A2(n1261), .ZN(n1059) );
AND2_X1 U974 ( .A1(n1169), .A2(n1262), .ZN(n1181) );
NAND2_X1 U975 ( .A1(n1048), .A2(n1263), .ZN(n1262) );
NAND4_X1 U976 ( .A1(G902), .A2(G953), .A3(n1206), .A4(n1116), .ZN(n1263) );
INV_X1 U977 ( .A(G898), .ZN(n1116) );
NAND3_X1 U978 ( .A1(n1206), .A2(n1087), .A3(G952), .ZN(n1048) );
NAND2_X1 U979 ( .A1(G237), .A2(G234), .ZN(n1206) );
NOR2_X1 U980 ( .A1(n1053), .A2(n1264), .ZN(n1169) );
AND2_X1 U981 ( .A1(G214), .A2(n1054), .ZN(n1264) );
XNOR2_X1 U982 ( .A(n1265), .B(n1156), .ZN(n1053) );
NAND2_X1 U983 ( .A1(G210), .A2(n1054), .ZN(n1156) );
NAND2_X1 U984 ( .A1(n1266), .A2(n1267), .ZN(n1054) );
INV_X1 U985 ( .A(G237), .ZN(n1267) );
XNOR2_X1 U986 ( .A(G902), .B(KEYINPUT43), .ZN(n1266) );
NAND2_X1 U987 ( .A1(n1268), .A2(n1218), .ZN(n1265) );
XOR2_X1 U988 ( .A(n1154), .B(KEYINPUT18), .Z(n1268) );
XOR2_X1 U989 ( .A(n1269), .B(n1270), .Z(n1154) );
XNOR2_X1 U990 ( .A(n1271), .B(n1272), .ZN(n1270) );
XOR2_X1 U991 ( .A(n1107), .B(n1273), .Z(n1272) );
NOR2_X1 U992 ( .A1(G953), .A2(n1115), .ZN(n1273) );
INV_X1 U993 ( .A(G224), .ZN(n1115) );
XOR2_X1 U994 ( .A(n1274), .B(n1275), .Z(n1107) );
XOR2_X1 U995 ( .A(KEYINPUT8), .B(KEYINPUT35), .Z(n1275) );
XOR2_X1 U996 ( .A(n1276), .B(n1139), .Z(n1274) );
NAND2_X1 U997 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND2_X1 U998 ( .A1(G104), .A2(n1010), .ZN(n1278) );
XOR2_X1 U999 ( .A(KEYINPUT2), .B(n1279), .Z(n1277) );
NOR2_X1 U1000 ( .A1(G104), .A2(n1010), .ZN(n1279) );
INV_X1 U1001 ( .A(G107), .ZN(n1010) );
XOR2_X1 U1002 ( .A(n1280), .B(n1281), .Z(n1269) );
NOR2_X1 U1003 ( .A1(KEYINPUT19), .A2(n1110), .ZN(n1281) );
XOR2_X1 U1004 ( .A(G110), .B(G122), .Z(n1110) );
XNOR2_X1 U1005 ( .A(G125), .B(n1282), .ZN(n1280) );
NOR2_X1 U1006 ( .A1(KEYINPUT28), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U1007 ( .A(n1213), .B(n1112), .ZN(n1283) );
AND2_X1 U1008 ( .A1(n1284), .A2(n1285), .ZN(n1112) );
NAND2_X1 U1009 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XNOR2_X1 U1010 ( .A(G119), .B(KEYINPUT31), .ZN(n1286) );
XOR2_X1 U1011 ( .A(KEYINPUT42), .B(n1288), .Z(n1284) );
NOR2_X1 U1012 ( .A1(G119), .A2(n1289), .ZN(n1288) );
XNOR2_X1 U1013 ( .A(G116), .B(KEYINPUT22), .ZN(n1289) );
AND2_X1 U1014 ( .A1(n1209), .A2(n1203), .ZN(n1047) );
NAND3_X1 U1015 ( .A1(n1290), .A2(n1291), .A3(n1062), .ZN(n1203) );
NAND3_X1 U1016 ( .A1(n1123), .A2(n1218), .A3(n1292), .ZN(n1062) );
INV_X1 U1017 ( .A(n1125), .ZN(n1292) );
NAND2_X1 U1018 ( .A1(n1123), .A2(n1293), .ZN(n1291) );
INV_X1 U1019 ( .A(KEYINPUT63), .ZN(n1293) );
NAND2_X1 U1020 ( .A1(n1074), .A2(KEYINPUT63), .ZN(n1290) );
NOR2_X1 U1021 ( .A1(n1123), .A2(n1294), .ZN(n1074) );
NOR2_X1 U1022 ( .A1(n1125), .A2(G902), .ZN(n1294) );
XNOR2_X1 U1023 ( .A(n1295), .B(n1296), .ZN(n1125) );
XNOR2_X1 U1024 ( .A(n1226), .B(n1297), .ZN(n1296) );
XOR2_X1 U1025 ( .A(n1298), .B(n1260), .Z(n1297) );
NAND2_X1 U1026 ( .A1(KEYINPUT48), .A2(G110), .ZN(n1298) );
XOR2_X1 U1027 ( .A(G140), .B(KEYINPUT53), .Z(n1226) );
XOR2_X1 U1028 ( .A(n1299), .B(n1300), .Z(n1295) );
NOR2_X1 U1029 ( .A1(G125), .A2(KEYINPUT55), .ZN(n1300) );
XOR2_X1 U1030 ( .A(n1301), .B(G119), .Z(n1299) );
NAND2_X1 U1031 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
XNOR2_X1 U1032 ( .A(G137), .B(n1304), .ZN(n1303) );
NAND3_X1 U1033 ( .A1(G234), .A2(n1305), .A3(G221), .ZN(n1304) );
XNOR2_X1 U1034 ( .A(KEYINPUT29), .B(n1087), .ZN(n1305) );
INV_X1 U1035 ( .A(G953), .ZN(n1087) );
XOR2_X1 U1036 ( .A(KEYINPUT57), .B(KEYINPUT47), .Z(n1302) );
NAND2_X1 U1037 ( .A1(G217), .A2(n1261), .ZN(n1123) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1218), .ZN(n1261) );
INV_X1 U1039 ( .A(G902), .ZN(n1218) );
XOR2_X1 U1040 ( .A(G472), .B(n1073), .Z(n1209) );
NAND2_X1 U1041 ( .A1(n1306), .A2(n1307), .ZN(n1073) );
XOR2_X1 U1042 ( .A(n1308), .B(n1309), .Z(n1307) );
NOR2_X1 U1043 ( .A1(KEYINPUT34), .A2(n1310), .ZN(n1309) );
XNOR2_X1 U1044 ( .A(n1142), .B(n1311), .ZN(n1310) );
INV_X1 U1045 ( .A(n1138), .ZN(n1311) );
XOR2_X1 U1046 ( .A(n1259), .B(n1312), .Z(n1138) );
INV_X1 U1047 ( .A(n1271), .ZN(n1312) );
XNOR2_X1 U1048 ( .A(n1313), .B(n1260), .ZN(n1271) );
XNOR2_X1 U1049 ( .A(G146), .B(n1201), .ZN(n1260) );
INV_X1 U1050 ( .A(G128), .ZN(n1201) );
NAND2_X1 U1051 ( .A1(KEYINPUT13), .A2(n1187), .ZN(n1313) );
INV_X1 U1052 ( .A(G143), .ZN(n1187) );
NAND2_X1 U1053 ( .A1(n1314), .A2(n1315), .ZN(n1259) );
NAND2_X1 U1054 ( .A1(n1097), .A2(n1197), .ZN(n1315) );
INV_X1 U1055 ( .A(G134), .ZN(n1197) );
NAND2_X1 U1056 ( .A1(n1316), .A2(G134), .ZN(n1314) );
XOR2_X1 U1057 ( .A(KEYINPUT21), .B(n1097), .Z(n1316) );
XNOR2_X1 U1058 ( .A(n1199), .B(n1317), .ZN(n1097) );
XOR2_X1 U1059 ( .A(KEYINPUT61), .B(G137), .Z(n1317) );
INV_X1 U1060 ( .A(G131), .ZN(n1199) );
AND3_X1 U1061 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1142) );
NAND2_X1 U1062 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NAND2_X1 U1063 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XNOR2_X1 U1064 ( .A(KEYINPUT16), .B(n1213), .ZN(n1323) );
XNOR2_X1 U1065 ( .A(G116), .B(G119), .ZN(n1321) );
NAND3_X1 U1066 ( .A1(G113), .A2(n1325), .A3(n1324), .ZN(n1319) );
INV_X1 U1067 ( .A(KEYINPUT52), .ZN(n1324) );
XNOR2_X1 U1068 ( .A(G119), .B(n1287), .ZN(n1325) );
INV_X1 U1069 ( .A(G116), .ZN(n1287) );
NAND2_X1 U1070 ( .A1(KEYINPUT52), .A2(n1213), .ZN(n1318) );
INV_X1 U1071 ( .A(G113), .ZN(n1213) );
XNOR2_X1 U1072 ( .A(n1326), .B(n1143), .ZN(n1308) );
NAND2_X1 U1073 ( .A1(G210), .A2(n1229), .ZN(n1143) );
NOR2_X1 U1074 ( .A1(G953), .A2(G237), .ZN(n1229) );
NAND2_X1 U1075 ( .A1(KEYINPUT26), .A2(n1139), .ZN(n1326) );
XOR2_X1 U1076 ( .A(G101), .B(KEYINPUT37), .Z(n1139) );
XNOR2_X1 U1077 ( .A(G902), .B(KEYINPUT39), .ZN(n1306) );
endmodule


