//Key = 1100010011111110011000001010110101110011101011111111001110011111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338;

NAND2_X1 U739 ( .A1(n1019), .A2(n1020), .ZN(G9) );
NAND2_X1 U740 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
XOR2_X1 U741 ( .A(KEYINPUT50), .B(n1023), .Z(n1019) );
NOR2_X1 U742 ( .A1(n1021), .A2(n1022), .ZN(n1023) );
XNOR2_X1 U743 ( .A(KEYINPUT33), .B(G107), .ZN(n1021) );
NOR2_X1 U744 ( .A1(n1024), .A2(n1025), .ZN(G75) );
XOR2_X1 U745 ( .A(KEYINPUT4), .B(n1026), .Z(n1025) );
NOR4_X1 U746 ( .A1(n1027), .A2(n1028), .A3(G953), .A4(n1029), .ZN(n1026) );
NOR2_X1 U747 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR2_X1 U748 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR3_X1 U749 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NOR2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U751 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U752 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U753 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U754 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(n1041) );
NOR2_X1 U756 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR3_X1 U757 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1049) );
INV_X1 U758 ( .A(KEYINPUT14), .ZN(n1051) );
NOR3_X1 U759 ( .A1(n1044), .A2(n1054), .A3(n1048), .ZN(n1037) );
NOR3_X1 U760 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NOR2_X1 U761 ( .A1(KEYINPUT14), .A2(n1040), .ZN(n1057) );
XOR2_X1 U762 ( .A(KEYINPUT52), .B(n1058), .Z(n1055) );
NOR4_X1 U763 ( .A1(n1059), .A2(n1048), .A3(n1044), .A4(n1040), .ZN(n1032) );
INV_X1 U764 ( .A(n1060), .ZN(n1048) );
NOR2_X1 U765 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR2_X1 U766 ( .A1(n1063), .A2(n1034), .ZN(n1061) );
NOR3_X1 U767 ( .A1(n1028), .A2(G953), .A3(G952), .ZN(n1024) );
AND4_X1 U768 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1028) );
NOR4_X1 U769 ( .A1(n1068), .A2(n1036), .A3(n1069), .A4(n1070), .ZN(n1067) );
XNOR2_X1 U770 ( .A(n1071), .B(KEYINPUT56), .ZN(n1069) );
INV_X1 U771 ( .A(n1072), .ZN(n1068) );
NOR3_X1 U772 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1066) );
NOR3_X1 U773 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
AND2_X1 U774 ( .A1(n1076), .A2(n1078), .ZN(n1074) );
INV_X1 U775 ( .A(KEYINPUT44), .ZN(n1076) );
XNOR2_X1 U776 ( .A(n1079), .B(n1080), .ZN(n1073) );
XNOR2_X1 U777 ( .A(G478), .B(KEYINPUT32), .ZN(n1080) );
XOR2_X1 U778 ( .A(n1081), .B(n1082), .Z(G72) );
XOR2_X1 U779 ( .A(n1083), .B(n1084), .Z(n1082) );
NOR2_X1 U780 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U781 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NAND2_X1 U782 ( .A1(n1089), .A2(n1090), .ZN(n1083) );
NAND2_X1 U783 ( .A1(G953), .A2(n1088), .ZN(n1090) );
XNOR2_X1 U784 ( .A(n1091), .B(n1092), .ZN(n1089) );
XNOR2_X1 U785 ( .A(KEYINPUT57), .B(n1093), .ZN(n1092) );
NOR2_X1 U786 ( .A1(KEYINPUT27), .A2(n1094), .ZN(n1093) );
XOR2_X1 U787 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U788 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U789 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U790 ( .A(KEYINPUT15), .B(G131), .Z(n1099) );
AND2_X1 U791 ( .A1(n1100), .A2(G131), .ZN(n1097) );
XNOR2_X1 U792 ( .A(n1101), .B(n1102), .ZN(n1100) );
NAND2_X1 U793 ( .A1(KEYINPUT11), .A2(G137), .ZN(n1101) );
NAND2_X1 U794 ( .A1(n1086), .A2(n1103), .ZN(n1081) );
XOR2_X1 U795 ( .A(n1104), .B(n1105), .Z(G69) );
XOR2_X1 U796 ( .A(n1106), .B(n1107), .Z(n1105) );
NAND2_X1 U797 ( .A1(G953), .A2(n1108), .ZN(n1107) );
NAND2_X1 U798 ( .A1(G898), .A2(G224), .ZN(n1108) );
NAND2_X1 U799 ( .A1(n1109), .A2(n1110), .ZN(n1106) );
XOR2_X1 U800 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U801 ( .A(n1113), .B(KEYINPUT36), .Z(n1109) );
NAND2_X1 U802 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XNOR2_X1 U803 ( .A(G953), .B(KEYINPUT26), .ZN(n1114) );
NOR2_X1 U804 ( .A1(n1116), .A2(G953), .ZN(n1104) );
NOR2_X1 U805 ( .A1(n1117), .A2(n1118), .ZN(G66) );
XNOR2_X1 U806 ( .A(n1119), .B(n1120), .ZN(n1118) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NOR2_X1 U808 ( .A1(n1117), .A2(n1123), .ZN(G63) );
XOR2_X1 U809 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND2_X1 U810 ( .A1(KEYINPUT34), .A2(n1126), .ZN(n1125) );
OR2_X1 U811 ( .A1(n1122), .A2(n1127), .ZN(n1124) );
NOR2_X1 U812 ( .A1(n1117), .A2(n1128), .ZN(G60) );
XOR2_X1 U813 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U814 ( .A1(n1131), .A2(n1122), .ZN(n1129) );
XOR2_X1 U815 ( .A(n1132), .B(n1133), .Z(G6) );
NAND2_X1 U816 ( .A1(KEYINPUT28), .A2(G104), .ZN(n1133) );
NOR2_X1 U817 ( .A1(n1117), .A2(n1134), .ZN(G57) );
XOR2_X1 U818 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U819 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U820 ( .A1(n1139), .A2(n1122), .ZN(n1138) );
XOR2_X1 U821 ( .A(n1140), .B(KEYINPUT10), .Z(n1135) );
NAND2_X1 U822 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NAND2_X1 U823 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U824 ( .A(KEYINPUT42), .B(n1145), .Z(n1141) );
NOR2_X1 U825 ( .A1(n1144), .A2(n1143), .ZN(n1145) );
XOR2_X1 U826 ( .A(n1146), .B(n1147), .Z(n1143) );
NAND2_X1 U827 ( .A1(KEYINPUT31), .A2(n1148), .ZN(n1146) );
XNOR2_X1 U828 ( .A(KEYINPUT62), .B(n1149), .ZN(n1148) );
NOR2_X1 U829 ( .A1(n1117), .A2(n1150), .ZN(G54) );
XOR2_X1 U830 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U831 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U832 ( .A1(n1155), .A2(n1122), .ZN(n1154) );
NAND2_X1 U833 ( .A1(KEYINPUT55), .A2(n1156), .ZN(n1153) );
XOR2_X1 U834 ( .A(n1157), .B(n1158), .Z(n1151) );
NAND2_X1 U835 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NAND2_X1 U836 ( .A1(G140), .A2(n1161), .ZN(n1160) );
XOR2_X1 U837 ( .A(KEYINPUT61), .B(n1162), .Z(n1159) );
NOR2_X1 U838 ( .A1(G140), .A2(n1161), .ZN(n1162) );
NOR2_X1 U839 ( .A1(n1117), .A2(n1163), .ZN(G51) );
XOR2_X1 U840 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U841 ( .A1(n1078), .A2(n1122), .ZN(n1165) );
NAND2_X1 U842 ( .A1(G902), .A2(n1027), .ZN(n1122) );
NAND2_X1 U843 ( .A1(n1116), .A2(n1166), .ZN(n1027) );
INV_X1 U844 ( .A(n1103), .ZN(n1166) );
NAND4_X1 U845 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1103) );
NOR4_X1 U846 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1170) );
INV_X1 U847 ( .A(n1175), .ZN(n1171) );
AND2_X1 U848 ( .A1(n1176), .A2(n1177), .ZN(n1169) );
NAND2_X1 U849 ( .A1(n1178), .A2(n1179), .ZN(n1167) );
INV_X1 U850 ( .A(n1180), .ZN(n1179) );
AND4_X1 U851 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1116) );
AND4_X1 U852 ( .A1(n1185), .A2(n1186), .A3(n1132), .A4(n1022), .ZN(n1184) );
NAND3_X1 U853 ( .A1(n1060), .A2(n1187), .A3(n1058), .ZN(n1022) );
NAND3_X1 U854 ( .A1(n1060), .A2(n1187), .A3(n1056), .ZN(n1132) );
NOR2_X1 U855 ( .A1(n1188), .A2(n1189), .ZN(n1183) );
NOR2_X1 U856 ( .A1(n1190), .A2(n1180), .ZN(n1189) );
NOR3_X1 U857 ( .A1(n1191), .A2(n1192), .A3(n1040), .ZN(n1188) );
INV_X1 U858 ( .A(n1193), .ZN(n1040) );
NAND3_X1 U859 ( .A1(n1194), .A2(n1195), .A3(n1046), .ZN(n1191) );
NAND2_X1 U860 ( .A1(KEYINPUT0), .A2(n1196), .ZN(n1195) );
NAND2_X1 U861 ( .A1(n1197), .A2(n1198), .ZN(n1194) );
INV_X1 U862 ( .A(KEYINPUT0), .ZN(n1198) );
NAND2_X1 U863 ( .A1(n1050), .A2(n1199), .ZN(n1197) );
NOR2_X1 U864 ( .A1(n1086), .A2(G952), .ZN(n1117) );
XNOR2_X1 U865 ( .A(G146), .B(n1168), .ZN(G48) );
NAND3_X1 U866 ( .A1(n1056), .A2(n1200), .A3(n1201), .ZN(n1168) );
XOR2_X1 U867 ( .A(n1177), .B(n1202), .Z(G45) );
XOR2_X1 U868 ( .A(KEYINPUT13), .B(G143), .Z(n1202) );
NAND3_X1 U869 ( .A1(n1046), .A2(n1200), .A3(n1203), .ZN(n1177) );
NOR3_X1 U870 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1203) );
XOR2_X1 U871 ( .A(n1174), .B(n1207), .Z(G42) );
XOR2_X1 U872 ( .A(KEYINPUT3), .B(G140), .Z(n1207) );
AND3_X1 U873 ( .A1(n1056), .A2(n1045), .A3(n1178), .ZN(n1174) );
XNOR2_X1 U874 ( .A(G137), .B(n1208), .ZN(G39) );
NAND4_X1 U875 ( .A1(n1209), .A2(n1201), .A3(n1210), .A4(n1193), .ZN(n1208) );
NOR2_X1 U876 ( .A1(n1036), .A2(n1034), .ZN(n1210) );
XNOR2_X1 U877 ( .A(n1050), .B(KEYINPUT54), .ZN(n1209) );
INV_X1 U878 ( .A(n1211), .ZN(n1050) );
XNOR2_X1 U879 ( .A(n1102), .B(n1173), .ZN(G36) );
AND3_X1 U880 ( .A1(n1046), .A2(n1058), .A3(n1178), .ZN(n1173) );
XOR2_X1 U881 ( .A(G131), .B(n1172), .Z(G33) );
AND3_X1 U882 ( .A1(n1056), .A2(n1046), .A3(n1178), .ZN(n1172) );
NOR4_X1 U883 ( .A1(n1034), .A2(n1211), .A3(n1036), .A4(n1205), .ZN(n1178) );
INV_X1 U884 ( .A(n1212), .ZN(n1205) );
XNOR2_X1 U885 ( .A(n1213), .B(n1214), .ZN(G30) );
NAND2_X1 U886 ( .A1(KEYINPUT47), .A2(n1176), .ZN(n1213) );
NAND3_X1 U887 ( .A1(n1058), .A2(n1200), .A3(n1201), .ZN(n1176) );
AND3_X1 U888 ( .A1(n1215), .A2(n1212), .A3(n1216), .ZN(n1201) );
XNOR2_X1 U889 ( .A(G101), .B(n1217), .ZN(G3) );
NAND3_X1 U890 ( .A1(n1193), .A2(n1187), .A3(n1046), .ZN(n1217) );
XNOR2_X1 U891 ( .A(G125), .B(n1175), .ZN(G27) );
NAND4_X1 U892 ( .A1(n1062), .A2(n1212), .A3(n1065), .A4(n1218), .ZN(n1175) );
AND2_X1 U893 ( .A1(n1045), .A2(n1056), .ZN(n1218) );
NAND2_X1 U894 ( .A1(n1219), .A2(n1031), .ZN(n1212) );
NAND4_X1 U895 ( .A1(G902), .A2(G953), .A3(n1220), .A4(n1088), .ZN(n1219) );
INV_X1 U896 ( .A(G900), .ZN(n1088) );
INV_X1 U897 ( .A(n1199), .ZN(n1062) );
XNOR2_X1 U898 ( .A(G122), .B(n1181), .ZN(G24) );
NAND4_X1 U899 ( .A1(n1221), .A2(n1060), .A3(n1071), .A4(n1222), .ZN(n1181) );
NOR2_X1 U900 ( .A1(n1215), .A2(n1216), .ZN(n1060) );
XNOR2_X1 U901 ( .A(n1223), .B(n1224), .ZN(G21) );
NOR3_X1 U902 ( .A1(n1180), .A2(KEYINPUT19), .A3(n1190), .ZN(n1224) );
INV_X1 U903 ( .A(n1221), .ZN(n1190) );
NAND3_X1 U904 ( .A1(n1216), .A2(n1215), .A3(n1193), .ZN(n1180) );
NAND2_X1 U905 ( .A1(n1225), .A2(n1226), .ZN(G18) );
NAND2_X1 U906 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NAND2_X1 U907 ( .A1(G116), .A2(n1229), .ZN(n1225) );
NAND2_X1 U908 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND2_X1 U909 ( .A1(KEYINPUT30), .A2(n1232), .ZN(n1231) );
INV_X1 U910 ( .A(n1182), .ZN(n1232) );
OR2_X1 U911 ( .A1(n1227), .A2(KEYINPUT30), .ZN(n1230) );
NOR2_X1 U912 ( .A1(KEYINPUT37), .A2(n1182), .ZN(n1227) );
NAND3_X1 U913 ( .A1(n1046), .A2(n1058), .A3(n1221), .ZN(n1182) );
NOR2_X1 U914 ( .A1(n1071), .A2(n1206), .ZN(n1058) );
INV_X1 U915 ( .A(n1222), .ZN(n1206) );
XNOR2_X1 U916 ( .A(n1186), .B(n1233), .ZN(G15) );
XNOR2_X1 U917 ( .A(KEYINPUT53), .B(n1234), .ZN(n1233) );
NAND3_X1 U918 ( .A1(n1221), .A2(n1046), .A3(n1056), .ZN(n1186) );
NOR2_X1 U919 ( .A1(n1222), .A2(n1204), .ZN(n1056) );
INV_X1 U920 ( .A(n1071), .ZN(n1204) );
NOR2_X1 U921 ( .A1(n1215), .A2(n1064), .ZN(n1046) );
NOR3_X1 U922 ( .A1(n1199), .A2(n1192), .A3(n1044), .ZN(n1221) );
INV_X1 U923 ( .A(n1065), .ZN(n1044) );
NOR2_X1 U924 ( .A1(n1053), .A2(n1235), .ZN(n1065) );
INV_X1 U925 ( .A(n1052), .ZN(n1235) );
NAND2_X1 U926 ( .A1(n1236), .A2(n1237), .ZN(G12) );
NAND2_X1 U927 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND2_X1 U928 ( .A1(G110), .A2(n1240), .ZN(n1239) );
OR2_X1 U929 ( .A1(KEYINPUT23), .A2(KEYINPUT29), .ZN(n1240) );
NAND3_X1 U930 ( .A1(n1241), .A2(n1242), .A3(KEYINPUT29), .ZN(n1236) );
OR2_X1 U931 ( .A1(G110), .A2(KEYINPUT23), .ZN(n1242) );
NAND2_X1 U932 ( .A1(G110), .A2(n1243), .ZN(n1241) );
OR2_X1 U933 ( .A1(n1238), .A2(KEYINPUT23), .ZN(n1243) );
INV_X1 U934 ( .A(n1185), .ZN(n1238) );
NAND3_X1 U935 ( .A1(n1193), .A2(n1187), .A3(n1045), .ZN(n1185) );
AND2_X1 U936 ( .A1(n1064), .A2(n1215), .ZN(n1045) );
XOR2_X1 U937 ( .A(n1070), .B(KEYINPUT25), .Z(n1215) );
XOR2_X1 U938 ( .A(n1244), .B(n1121), .Z(n1070) );
NAND2_X1 U939 ( .A1(G217), .A2(n1245), .ZN(n1121) );
NAND2_X1 U940 ( .A1(G234), .A2(n1246), .ZN(n1245) );
NAND2_X1 U941 ( .A1(n1119), .A2(n1246), .ZN(n1244) );
XNOR2_X1 U942 ( .A(n1247), .B(n1248), .ZN(n1119) );
XOR2_X1 U943 ( .A(n1249), .B(n1250), .Z(n1248) );
XNOR2_X1 U944 ( .A(G137), .B(n1223), .ZN(n1250) );
XOR2_X1 U945 ( .A(KEYINPUT6), .B(G146), .Z(n1249) );
XOR2_X1 U946 ( .A(n1251), .B(n1252), .Z(n1247) );
XNOR2_X1 U947 ( .A(n1161), .B(n1253), .ZN(n1252) );
XOR2_X1 U948 ( .A(n1254), .B(n1255), .Z(n1251) );
NOR2_X1 U949 ( .A1(G128), .A2(KEYINPUT2), .ZN(n1255) );
NAND3_X1 U950 ( .A1(G234), .A2(n1256), .A3(G221), .ZN(n1254) );
XNOR2_X1 U951 ( .A(KEYINPUT59), .B(n1257), .ZN(n1256) );
INV_X1 U952 ( .A(n1216), .ZN(n1064) );
XOR2_X1 U953 ( .A(n1258), .B(n1139), .Z(n1216) );
INV_X1 U954 ( .A(G472), .ZN(n1139) );
NAND2_X1 U955 ( .A1(n1259), .A2(n1246), .ZN(n1258) );
XOR2_X1 U956 ( .A(n1260), .B(n1261), .Z(n1259) );
XOR2_X1 U957 ( .A(n1144), .B(n1137), .Z(n1261) );
XOR2_X1 U958 ( .A(n1262), .B(G101), .Z(n1137) );
NAND2_X1 U959 ( .A1(G210), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U960 ( .A(G113), .B(n1264), .ZN(n1144) );
XNOR2_X1 U961 ( .A(n1223), .B(G116), .ZN(n1264) );
INV_X1 U962 ( .A(G119), .ZN(n1223) );
XNOR2_X1 U963 ( .A(n1147), .B(n1265), .ZN(n1260) );
NOR2_X1 U964 ( .A1(KEYINPUT43), .A2(n1149), .ZN(n1265) );
NOR2_X1 U965 ( .A1(n1196), .A2(n1192), .ZN(n1187) );
AND2_X1 U966 ( .A1(n1031), .A2(n1266), .ZN(n1192) );
NAND4_X1 U967 ( .A1(G902), .A2(G953), .A3(n1220), .A4(n1115), .ZN(n1266) );
INV_X1 U968 ( .A(G898), .ZN(n1115) );
NAND3_X1 U969 ( .A1(n1220), .A2(n1086), .A3(G952), .ZN(n1031) );
INV_X1 U970 ( .A(G953), .ZN(n1086) );
NAND2_X1 U971 ( .A1(G237), .A2(G234), .ZN(n1220) );
INV_X1 U972 ( .A(n1200), .ZN(n1196) );
NOR2_X1 U973 ( .A1(n1199), .A2(n1211), .ZN(n1200) );
NAND2_X1 U974 ( .A1(n1053), .A2(n1052), .ZN(n1211) );
NAND2_X1 U975 ( .A1(G221), .A2(n1267), .ZN(n1052) );
XOR2_X1 U976 ( .A(KEYINPUT38), .B(n1268), .Z(n1267) );
AND2_X1 U977 ( .A1(n1246), .A2(G234), .ZN(n1268) );
XOR2_X1 U978 ( .A(n1269), .B(n1155), .Z(n1053) );
INV_X1 U979 ( .A(G469), .ZN(n1155) );
NAND2_X1 U980 ( .A1(n1270), .A2(n1246), .ZN(n1269) );
XOR2_X1 U981 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U982 ( .A(n1158), .B(n1273), .Z(n1272) );
XOR2_X1 U983 ( .A(KEYINPUT49), .B(KEYINPUT16), .Z(n1273) );
NOR2_X1 U984 ( .A1(n1087), .A2(n1274), .ZN(n1158) );
INV_X1 U985 ( .A(G227), .ZN(n1087) );
XNOR2_X1 U986 ( .A(n1275), .B(n1156), .ZN(n1271) );
XOR2_X1 U987 ( .A(n1276), .B(n1277), .Z(n1156) );
XOR2_X1 U988 ( .A(n1147), .B(n1278), .Z(n1277) );
XNOR2_X1 U989 ( .A(n1279), .B(G104), .ZN(n1278) );
XOR2_X1 U990 ( .A(G131), .B(n1280), .Z(n1147) );
XNOR2_X1 U991 ( .A(G137), .B(n1102), .ZN(n1280) );
XNOR2_X1 U992 ( .A(n1095), .B(n1281), .ZN(n1276) );
XOR2_X1 U993 ( .A(n1282), .B(n1283), .Z(n1095) );
NAND2_X1 U994 ( .A1(KEYINPUT45), .A2(n1214), .ZN(n1282) );
NAND2_X1 U995 ( .A1(KEYINPUT51), .A2(n1284), .ZN(n1275) );
XOR2_X1 U996 ( .A(n1161), .B(n1285), .Z(n1284) );
XOR2_X1 U997 ( .A(KEYINPUT58), .B(G140), .Z(n1285) );
NAND2_X1 U998 ( .A1(n1286), .A2(n1034), .ZN(n1199) );
NAND2_X1 U999 ( .A1(n1287), .A2(n1072), .ZN(n1034) );
NAND2_X1 U1000 ( .A1(n1077), .A2(n1078), .ZN(n1072) );
OR2_X1 U1001 ( .A1(n1078), .A2(n1077), .ZN(n1287) );
NOR2_X1 U1002 ( .A1(n1164), .A2(G902), .ZN(n1077) );
XOR2_X1 U1003 ( .A(n1288), .B(n1289), .Z(n1164) );
XNOR2_X1 U1004 ( .A(n1290), .B(n1291), .ZN(n1289) );
INV_X1 U1005 ( .A(n1149), .ZN(n1291) );
XOR2_X1 U1006 ( .A(n1283), .B(n1214), .Z(n1149) );
XNOR2_X1 U1007 ( .A(G146), .B(n1292), .ZN(n1283) );
NAND2_X1 U1008 ( .A1(G224), .A2(n1257), .ZN(n1290) );
XNOR2_X1 U1009 ( .A(n1293), .B(n1294), .ZN(n1288) );
INV_X1 U1010 ( .A(G125), .ZN(n1294) );
NAND2_X1 U1011 ( .A1(n1295), .A2(n1296), .ZN(n1293) );
NAND2_X1 U1012 ( .A1(n1297), .A2(n1111), .ZN(n1296) );
XOR2_X1 U1013 ( .A(KEYINPUT18), .B(n1298), .Z(n1295) );
NOR2_X1 U1014 ( .A1(n1297), .A2(n1111), .ZN(n1298) );
NAND2_X1 U1015 ( .A1(n1299), .A2(n1300), .ZN(n1111) );
NAND2_X1 U1016 ( .A1(n1301), .A2(n1234), .ZN(n1300) );
XOR2_X1 U1017 ( .A(KEYINPUT40), .B(n1302), .Z(n1301) );
NAND2_X1 U1018 ( .A1(n1302), .A2(G113), .ZN(n1299) );
XNOR2_X1 U1019 ( .A(n1303), .B(n1304), .ZN(n1302) );
NOR2_X1 U1020 ( .A1(G116), .A2(KEYINPUT7), .ZN(n1304) );
XNOR2_X1 U1021 ( .A(G119), .B(n1305), .ZN(n1303) );
NOR2_X1 U1022 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XOR2_X1 U1023 ( .A(n1308), .B(KEYINPUT9), .Z(n1307) );
NAND2_X1 U1024 ( .A1(n1309), .A2(n1281), .ZN(n1308) );
NOR2_X1 U1025 ( .A1(n1281), .A2(n1309), .ZN(n1306) );
XOR2_X1 U1026 ( .A(n1310), .B(G104), .Z(n1309) );
NAND2_X1 U1027 ( .A1(KEYINPUT46), .A2(n1279), .ZN(n1310) );
XNOR2_X1 U1028 ( .A(G101), .B(KEYINPUT17), .ZN(n1281) );
XNOR2_X1 U1029 ( .A(KEYINPUT8), .B(n1112), .ZN(n1297) );
XNOR2_X1 U1030 ( .A(n1311), .B(n1161), .ZN(n1112) );
XOR2_X1 U1031 ( .A(G110), .B(KEYINPUT1), .Z(n1161) );
XNOR2_X1 U1032 ( .A(G122), .B(KEYINPUT22), .ZN(n1311) );
NAND2_X1 U1033 ( .A1(G210), .A2(n1312), .ZN(n1078) );
XNOR2_X1 U1034 ( .A(n1036), .B(KEYINPUT21), .ZN(n1286) );
INV_X1 U1035 ( .A(n1063), .ZN(n1036) );
NAND2_X1 U1036 ( .A1(G214), .A2(n1312), .ZN(n1063) );
NAND2_X1 U1037 ( .A1(n1313), .A2(n1246), .ZN(n1312) );
INV_X1 U1038 ( .A(G902), .ZN(n1246) );
INV_X1 U1039 ( .A(G237), .ZN(n1313) );
NOR2_X1 U1040 ( .A1(n1222), .A2(n1071), .ZN(n1193) );
XOR2_X1 U1041 ( .A(n1314), .B(n1131), .Z(n1071) );
INV_X1 U1042 ( .A(G475), .ZN(n1131) );
OR2_X1 U1043 ( .A1(n1130), .A2(G902), .ZN(n1314) );
XNOR2_X1 U1044 ( .A(n1315), .B(n1316), .ZN(n1130) );
XOR2_X1 U1045 ( .A(n1317), .B(n1318), .Z(n1316) );
XNOR2_X1 U1046 ( .A(n1234), .B(n1319), .ZN(n1318) );
NOR2_X1 U1047 ( .A1(KEYINPUT41), .A2(n1320), .ZN(n1319) );
XNOR2_X1 U1048 ( .A(n1321), .B(n1322), .ZN(n1320) );
XOR2_X1 U1049 ( .A(n1323), .B(KEYINPUT5), .Z(n1322) );
NAND2_X1 U1050 ( .A1(G214), .A2(n1263), .ZN(n1323) );
NOR2_X1 U1051 ( .A1(n1274), .A2(G237), .ZN(n1263) );
INV_X1 U1052 ( .A(G113), .ZN(n1234) );
XOR2_X1 U1053 ( .A(G131), .B(G122), .Z(n1317) );
XNOR2_X1 U1054 ( .A(n1324), .B(n1253), .ZN(n1315) );
INV_X1 U1055 ( .A(n1091), .ZN(n1253) );
XOR2_X1 U1056 ( .A(G125), .B(G140), .Z(n1091) );
XNOR2_X1 U1057 ( .A(n1325), .B(n1326), .ZN(n1324) );
NAND2_X1 U1058 ( .A1(KEYINPUT60), .A2(G146), .ZN(n1326) );
NAND2_X1 U1059 ( .A1(n1327), .A2(KEYINPUT35), .ZN(n1325) );
XNOR2_X1 U1060 ( .A(G104), .B(KEYINPUT12), .ZN(n1327) );
XOR2_X1 U1061 ( .A(n1328), .B(n1127), .Z(n1222) );
INV_X1 U1062 ( .A(G478), .ZN(n1127) );
NAND2_X1 U1063 ( .A1(KEYINPUT24), .A2(n1079), .ZN(n1328) );
NOR2_X1 U1064 ( .A1(G902), .A2(n1126), .ZN(n1079) );
AND2_X1 U1065 ( .A1(n1329), .A2(n1330), .ZN(n1126) );
NAND4_X1 U1066 ( .A1(G234), .A2(G217), .A3(n1257), .A4(n1331), .ZN(n1330) );
XOR2_X1 U1067 ( .A(KEYINPUT63), .B(n1332), .Z(n1331) );
NAND2_X1 U1068 ( .A1(n1332), .A2(n1333), .ZN(n1329) );
NAND3_X1 U1069 ( .A1(n1257), .A2(G217), .A3(G234), .ZN(n1333) );
INV_X1 U1070 ( .A(n1274), .ZN(n1257) );
XOR2_X1 U1071 ( .A(G953), .B(KEYINPUT20), .Z(n1274) );
XNOR2_X1 U1072 ( .A(n1334), .B(n1335), .ZN(n1332) );
XNOR2_X1 U1073 ( .A(n1228), .B(n1336), .ZN(n1335) );
XNOR2_X1 U1074 ( .A(n1214), .B(G122), .ZN(n1336) );
INV_X1 U1075 ( .A(G128), .ZN(n1214) );
INV_X1 U1076 ( .A(G116), .ZN(n1228) );
XNOR2_X1 U1077 ( .A(n1337), .B(n1292), .ZN(n1334) );
INV_X1 U1078 ( .A(n1321), .ZN(n1292) );
XOR2_X1 U1079 ( .A(G143), .B(KEYINPUT48), .Z(n1321) );
XNOR2_X1 U1080 ( .A(n1338), .B(n1279), .ZN(n1337) );
INV_X1 U1081 ( .A(G107), .ZN(n1279) );
NAND2_X1 U1082 ( .A1(KEYINPUT39), .A2(n1102), .ZN(n1338) );
INV_X1 U1083 ( .A(G134), .ZN(n1102) );
endmodule


