//Key = 0111101001101110001110011111110110100010111101011001100010100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290;

XOR2_X1 U720 ( .A(G107), .B(n986), .Z(G9) );
NOR2_X1 U721 ( .A1(n987), .A2(n988), .ZN(G75) );
NOR2_X1 U722 ( .A1(n989), .A2(n990), .ZN(n988) );
NAND4_X1 U723 ( .A1(n991), .A2(n992), .A3(n993), .A4(n994), .ZN(n990) );
NAND2_X1 U724 ( .A1(n995), .A2(n996), .ZN(n994) );
NAND2_X1 U725 ( .A1(n997), .A2(n998), .ZN(n996) );
NAND3_X1 U726 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n998) );
NAND2_X1 U727 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NAND2_X1 U728 ( .A1(n1004), .A2(n1005), .ZN(n1002) );
INV_X1 U729 ( .A(KEYINPUT1), .ZN(n1005) );
NAND4_X1 U730 ( .A1(n1006), .A2(n1007), .A3(n1008), .A4(n1009), .ZN(n999) );
NAND2_X1 U731 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NAND3_X1 U732 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1007) );
NAND2_X1 U733 ( .A1(n1015), .A2(n1016), .ZN(n1012) );
NAND2_X1 U734 ( .A1(KEYINPUT1), .A2(n1004), .ZN(n1006) );
AND3_X1 U735 ( .A1(n1010), .A2(n1014), .A3(n1017), .ZN(n1004) );
NAND2_X1 U736 ( .A1(n1018), .A2(n1019), .ZN(n997) );
NAND2_X1 U737 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U738 ( .A1(KEYINPUT51), .A2(n1022), .ZN(n1021) );
NAND4_X1 U739 ( .A1(n1022), .A2(n1023), .A3(n1018), .A4(n1024), .ZN(n993) );
INV_X1 U740 ( .A(KEYINPUT51), .ZN(n1023) );
NAND4_X1 U741 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n989) );
NAND3_X1 U742 ( .A1(n1001), .A2(n1029), .A3(n1018), .ZN(n1026) );
AND4_X1 U743 ( .A1(n1009), .A2(n1010), .A3(n1014), .A4(n1013), .ZN(n1018) );
INV_X1 U744 ( .A(n1003), .ZN(n1009) );
NAND2_X1 U745 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U746 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
XNOR2_X1 U747 ( .A(KEYINPUT63), .B(n1034), .ZN(n1033) );
NOR3_X1 U748 ( .A1(n1035), .A2(G953), .A3(G952), .ZN(n987) );
INV_X1 U749 ( .A(n1027), .ZN(n1035) );
NAND4_X1 U750 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1027) );
NOR4_X1 U751 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
XNOR2_X1 U752 ( .A(KEYINPUT0), .B(n1044), .ZN(n1043) );
XNOR2_X1 U753 ( .A(G475), .B(n1045), .ZN(n1042) );
NAND2_X1 U754 ( .A1(KEYINPUT27), .A2(n1046), .ZN(n1045) );
NOR2_X1 U755 ( .A1(n1032), .A2(n1017), .ZN(n1038) );
XNOR2_X1 U756 ( .A(G469), .B(n1047), .ZN(n1037) );
NAND2_X1 U757 ( .A1(KEYINPUT24), .A2(n1048), .ZN(n1047) );
XOR2_X1 U758 ( .A(n1049), .B(n1050), .Z(G72) );
XOR2_X1 U759 ( .A(n1051), .B(n1052), .Z(n1050) );
NOR3_X1 U760 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NOR2_X1 U761 ( .A1(G900), .A2(n1028), .ZN(n1055) );
NOR2_X1 U762 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
XOR2_X1 U763 ( .A(n1058), .B(KEYINPUT61), .Z(n1053) );
NAND2_X1 U764 ( .A1(n1057), .A2(n1056), .ZN(n1058) );
XNOR2_X1 U765 ( .A(n1059), .B(n1060), .ZN(n1057) );
NAND2_X1 U766 ( .A1(n1061), .A2(n1062), .ZN(n1051) );
NAND2_X1 U767 ( .A1(G900), .A2(G227), .ZN(n1062) );
XNOR2_X1 U768 ( .A(G953), .B(KEYINPUT45), .ZN(n1061) );
NAND2_X1 U769 ( .A1(n1028), .A2(n1063), .ZN(n1049) );
XOR2_X1 U770 ( .A(n1064), .B(n1065), .Z(G69) );
XOR2_X1 U771 ( .A(n1066), .B(n1067), .Z(n1065) );
NOR2_X1 U772 ( .A1(n1068), .A2(n1028), .ZN(n1067) );
AND2_X1 U773 ( .A1(G224), .A2(G898), .ZN(n1068) );
NAND2_X1 U774 ( .A1(n1069), .A2(n1070), .ZN(n1066) );
NAND2_X1 U775 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XNOR2_X1 U776 ( .A(G953), .B(KEYINPUT34), .ZN(n1071) );
XOR2_X1 U777 ( .A(n1073), .B(n1074), .Z(n1069) );
XOR2_X1 U778 ( .A(n1075), .B(KEYINPUT13), .Z(n1074) );
NAND2_X1 U779 ( .A1(n1028), .A2(n1076), .ZN(n1064) );
NAND2_X1 U780 ( .A1(n992), .A2(n1077), .ZN(n1076) );
NOR2_X1 U781 ( .A1(n1078), .A2(n1079), .ZN(G66) );
XOR2_X1 U782 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U783 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NOR2_X1 U784 ( .A1(n1078), .A2(n1084), .ZN(G63) );
XOR2_X1 U785 ( .A(n1085), .B(n1086), .Z(n1084) );
XNOR2_X1 U786 ( .A(KEYINPUT60), .B(n1087), .ZN(n1086) );
AND2_X1 U787 ( .A1(G478), .A2(n1088), .ZN(n1085) );
NOR2_X1 U788 ( .A1(n1078), .A2(n1089), .ZN(G60) );
XOR2_X1 U789 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U790 ( .A1(n1092), .A2(KEYINPUT50), .ZN(n1091) );
AND2_X1 U791 ( .A1(G475), .A2(n1088), .ZN(n1092) );
XNOR2_X1 U792 ( .A(G104), .B(n1093), .ZN(G6) );
NOR2_X1 U793 ( .A1(n1078), .A2(n1094), .ZN(G57) );
XOR2_X1 U794 ( .A(n1095), .B(n1096), .Z(n1094) );
XOR2_X1 U795 ( .A(n1097), .B(n1098), .Z(n1095) );
NOR2_X1 U796 ( .A1(n1099), .A2(n1083), .ZN(n1098) );
XNOR2_X1 U797 ( .A(G472), .B(KEYINPUT46), .ZN(n1099) );
NAND2_X1 U798 ( .A1(KEYINPUT43), .A2(n1100), .ZN(n1097) );
NOR2_X1 U799 ( .A1(n1078), .A2(n1101), .ZN(G54) );
XOR2_X1 U800 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U801 ( .A(n1104), .B(n1105), .Z(n1103) );
XNOR2_X1 U802 ( .A(n1106), .B(n1107), .ZN(n1105) );
NAND2_X1 U803 ( .A1(KEYINPUT38), .A2(n1108), .ZN(n1107) );
NAND2_X1 U804 ( .A1(KEYINPUT23), .A2(n1060), .ZN(n1106) );
XOR2_X1 U805 ( .A(n1059), .B(n1109), .Z(n1104) );
AND2_X1 U806 ( .A1(G469), .A2(n1088), .ZN(n1109) );
XOR2_X1 U807 ( .A(n1110), .B(n1111), .Z(n1102) );
XOR2_X1 U808 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U809 ( .A1(KEYINPUT15), .A2(n1114), .ZN(n1113) );
XNOR2_X1 U810 ( .A(n1115), .B(KEYINPUT47), .ZN(n1114) );
XNOR2_X1 U811 ( .A(KEYINPUT35), .B(n1116), .ZN(n1110) );
NOR2_X1 U812 ( .A1(n1078), .A2(n1117), .ZN(G51) );
XOR2_X1 U813 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND3_X1 U814 ( .A1(n1088), .A2(n1120), .A3(KEYINPUT52), .ZN(n1118) );
INV_X1 U815 ( .A(n1083), .ZN(n1088) );
NAND2_X1 U816 ( .A1(G902), .A2(n1121), .ZN(n1083) );
NAND3_X1 U817 ( .A1(n992), .A2(n1025), .A3(n991), .ZN(n1121) );
INV_X1 U818 ( .A(n1063), .ZN(n991) );
NAND4_X1 U819 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1063) );
NOR4_X1 U820 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n1125) );
NAND2_X1 U821 ( .A1(n1130), .A2(n1131), .ZN(n1124) );
NAND2_X1 U822 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NAND2_X1 U823 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XNOR2_X1 U824 ( .A(KEYINPUT14), .B(n1136), .ZN(n1135) );
INV_X1 U825 ( .A(n1137), .ZN(n1134) );
NAND2_X1 U826 ( .A1(n1138), .A2(n1139), .ZN(n1132) );
XNOR2_X1 U827 ( .A(n1077), .B(KEYINPUT56), .ZN(n1025) );
AND4_X1 U828 ( .A1(n1093), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n992) );
NOR4_X1 U829 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n986), .ZN(n1142) );
AND3_X1 U830 ( .A1(n1146), .A2(n1001), .A3(n1147), .ZN(n986) );
NAND3_X1 U831 ( .A1(n1148), .A2(n1001), .A3(n1149), .ZN(n1141) );
NAND3_X1 U832 ( .A1(n1147), .A2(n1001), .A3(n1130), .ZN(n1093) );
NOR2_X1 U833 ( .A1(n1028), .A2(G952), .ZN(n1078) );
XNOR2_X1 U834 ( .A(n1150), .B(n1151), .ZN(G48) );
NOR3_X1 U835 ( .A1(n1137), .A2(n1152), .A3(n1015), .ZN(n1151) );
XNOR2_X1 U836 ( .A(G143), .B(n1122), .ZN(G45) );
NAND4_X1 U837 ( .A1(n1148), .A2(n1022), .A3(n1153), .A4(n1011), .ZN(n1122) );
NOR2_X1 U838 ( .A1(n1152), .A2(n1031), .ZN(n1153) );
XOR2_X1 U839 ( .A(n1154), .B(n1155), .Z(G42) );
XNOR2_X1 U840 ( .A(KEYINPUT49), .B(n1116), .ZN(n1155) );
NOR3_X1 U841 ( .A1(n1156), .A2(n1015), .A3(n1157), .ZN(n1154) );
XNOR2_X1 U842 ( .A(KEYINPUT2), .B(n1020), .ZN(n1156) );
XNOR2_X1 U843 ( .A(G137), .B(n1123), .ZN(G39) );
NAND4_X1 U844 ( .A1(n1010), .A2(n1138), .A3(n1158), .A4(n1041), .ZN(n1123) );
XOR2_X1 U845 ( .A(G134), .B(n1129), .Z(G36) );
AND3_X1 U846 ( .A1(n1138), .A2(n1146), .A3(n1022), .ZN(n1129) );
NAND2_X1 U847 ( .A1(n1159), .A2(n1160), .ZN(G33) );
NAND2_X1 U848 ( .A1(n1128), .A2(n1161), .ZN(n1160) );
XOR2_X1 U849 ( .A(KEYINPUT6), .B(n1162), .Z(n1159) );
NOR2_X1 U850 ( .A1(n1128), .A2(n1161), .ZN(n1162) );
INV_X1 U851 ( .A(G131), .ZN(n1161) );
AND3_X1 U852 ( .A1(n1138), .A2(n1130), .A3(n1022), .ZN(n1128) );
INV_X1 U853 ( .A(n1157), .ZN(n1138) );
NAND4_X1 U854 ( .A1(n1163), .A2(n1014), .A3(n1136), .A4(n1013), .ZN(n1157) );
XNOR2_X1 U855 ( .A(n1164), .B(KEYINPUT4), .ZN(n1014) );
XOR2_X1 U856 ( .A(G128), .B(n1127), .Z(G30) );
NOR3_X1 U857 ( .A1(n1016), .A2(n1152), .A3(n1137), .ZN(n1127) );
NAND4_X1 U858 ( .A1(n1011), .A2(n1158), .A3(n1163), .A4(n1041), .ZN(n1137) );
INV_X1 U859 ( .A(n1146), .ZN(n1016) );
XNOR2_X1 U860 ( .A(G101), .B(n1140), .ZN(G3) );
NAND3_X1 U861 ( .A1(n1022), .A2(n1147), .A3(n1010), .ZN(n1140) );
XOR2_X1 U862 ( .A(G125), .B(n1126), .Z(G27) );
AND4_X1 U863 ( .A1(n1139), .A2(n1130), .A3(n1165), .A4(n1011), .ZN(n1126) );
NOR2_X1 U864 ( .A1(n1152), .A2(n1024), .ZN(n1165) );
INV_X1 U865 ( .A(n995), .ZN(n1024) );
INV_X1 U866 ( .A(n1136), .ZN(n1152) );
NAND2_X1 U867 ( .A1(n1003), .A2(n1166), .ZN(n1136) );
NAND4_X1 U868 ( .A1(G953), .A2(G902), .A3(n1167), .A4(n1168), .ZN(n1166) );
INV_X1 U869 ( .A(G900), .ZN(n1168) );
XOR2_X1 U870 ( .A(n1169), .B(n1170), .Z(G24) );
NOR2_X1 U871 ( .A1(KEYINPUT11), .A2(n1171), .ZN(n1170) );
NOR3_X1 U872 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1169) );
INV_X1 U873 ( .A(n1001), .ZN(n1174) );
NOR2_X1 U874 ( .A1(n1041), .A2(n1158), .ZN(n1001) );
XNOR2_X1 U875 ( .A(n1148), .B(KEYINPUT44), .ZN(n1173) );
AND2_X1 U876 ( .A1(n1175), .A2(n1176), .ZN(n1148) );
XOR2_X1 U877 ( .A(n1145), .B(n1177), .Z(G21) );
NOR2_X1 U878 ( .A1(KEYINPUT8), .A2(n1178), .ZN(n1177) );
AND4_X1 U879 ( .A1(n1149), .A2(n1010), .A3(n1158), .A4(n1041), .ZN(n1145) );
INV_X1 U880 ( .A(n1179), .ZN(n1158) );
XOR2_X1 U881 ( .A(G116), .B(n1144), .Z(G18) );
AND3_X1 U882 ( .A1(n1022), .A2(n1146), .A3(n1149), .ZN(n1144) );
INV_X1 U883 ( .A(n1172), .ZN(n1149) );
NAND3_X1 U884 ( .A1(n995), .A2(n1180), .A3(n1011), .ZN(n1172) );
XNOR2_X1 U885 ( .A(n1181), .B(KEYINPUT58), .ZN(n1011) );
NOR2_X1 U886 ( .A1(n1176), .A2(n1044), .ZN(n1146) );
XOR2_X1 U887 ( .A(G113), .B(n1143), .Z(G15) );
AND4_X1 U888 ( .A1(n1022), .A2(n1130), .A3(n1182), .A4(n1181), .ZN(n1143) );
AND2_X1 U889 ( .A1(n1180), .A2(n995), .ZN(n1182) );
NAND2_X1 U890 ( .A1(n1183), .A2(n1184), .ZN(n995) );
OR2_X1 U891 ( .A1(n1031), .A2(KEYINPUT63), .ZN(n1184) );
INV_X1 U892 ( .A(n1163), .ZN(n1031) );
NAND3_X1 U893 ( .A1(n1034), .A2(n1185), .A3(KEYINPUT63), .ZN(n1183) );
INV_X1 U894 ( .A(n1015), .ZN(n1130) );
NAND2_X1 U895 ( .A1(n1044), .A2(n1176), .ZN(n1015) );
INV_X1 U896 ( .A(n1175), .ZN(n1044) );
NOR2_X1 U897 ( .A1(n1179), .A2(n1041), .ZN(n1022) );
XNOR2_X1 U898 ( .A(G110), .B(n1077), .ZN(G12) );
NAND3_X1 U899 ( .A1(n1139), .A2(n1147), .A3(n1010), .ZN(n1077) );
NOR2_X1 U900 ( .A1(n1175), .A2(n1176), .ZN(n1010) );
XOR2_X1 U901 ( .A(G475), .B(n1046), .Z(n1176) );
AND2_X1 U902 ( .A1(n1090), .A2(n1186), .ZN(n1046) );
XOR2_X1 U903 ( .A(n1187), .B(n1188), .Z(n1090) );
XNOR2_X1 U904 ( .A(n1189), .B(n1190), .ZN(n1188) );
INV_X1 U905 ( .A(n1191), .ZN(n1190) );
NOR2_X1 U906 ( .A1(n1192), .A2(n1193), .ZN(n1189) );
INV_X1 U907 ( .A(G214), .ZN(n1192) );
XOR2_X1 U908 ( .A(n1194), .B(n1195), .Z(n1187) );
NOR2_X1 U909 ( .A1(KEYINPUT59), .A2(n1196), .ZN(n1195) );
XOR2_X1 U910 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U911 ( .A(n1199), .B(G104), .Z(n1198) );
NAND2_X1 U912 ( .A1(KEYINPUT12), .A2(n1171), .ZN(n1199) );
XNOR2_X1 U913 ( .A(G113), .B(KEYINPUT41), .ZN(n1197) );
XNOR2_X1 U914 ( .A(G131), .B(G143), .ZN(n1194) );
XNOR2_X1 U915 ( .A(n1200), .B(G478), .ZN(n1175) );
NAND2_X1 U916 ( .A1(n1186), .A2(n1087), .ZN(n1200) );
NAND2_X1 U917 ( .A1(n1201), .A2(n1202), .ZN(n1087) );
NAND2_X1 U918 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NAND3_X1 U919 ( .A1(n1205), .A2(n1028), .A3(G217), .ZN(n1204) );
XNOR2_X1 U920 ( .A(n1206), .B(n1207), .ZN(n1203) );
XOR2_X1 U921 ( .A(n1208), .B(KEYINPUT39), .Z(n1201) );
NAND4_X1 U922 ( .A1(n1209), .A2(G217), .A3(n1205), .A4(n1028), .ZN(n1208) );
XNOR2_X1 U923 ( .A(G234), .B(KEYINPUT3), .ZN(n1205) );
XNOR2_X1 U924 ( .A(n1206), .B(n1210), .ZN(n1209) );
INV_X1 U925 ( .A(n1207), .ZN(n1210) );
XNOR2_X1 U926 ( .A(n1211), .B(n1212), .ZN(n1207) );
XNOR2_X1 U927 ( .A(G134), .B(G143), .ZN(n1211) );
NAND2_X1 U928 ( .A1(n1213), .A2(KEYINPUT42), .ZN(n1206) );
XNOR2_X1 U929 ( .A(G107), .B(n1214), .ZN(n1213) );
XNOR2_X1 U930 ( .A(n1171), .B(G116), .ZN(n1214) );
AND3_X1 U931 ( .A1(n1163), .A2(n1180), .A3(n1181), .ZN(n1147) );
NOR2_X1 U932 ( .A1(n1164), .A2(n1017), .ZN(n1181) );
INV_X1 U933 ( .A(n1013), .ZN(n1017) );
NAND2_X1 U934 ( .A1(G214), .A2(n1215), .ZN(n1013) );
XOR2_X1 U935 ( .A(n1036), .B(n1216), .Z(n1164) );
XOR2_X1 U936 ( .A(KEYINPUT36), .B(KEYINPUT17), .Z(n1216) );
XOR2_X1 U937 ( .A(n1217), .B(n1120), .Z(n1036) );
AND2_X1 U938 ( .A1(G210), .A2(n1215), .ZN(n1120) );
NAND2_X1 U939 ( .A1(n1218), .A2(n1186), .ZN(n1215) );
NAND2_X1 U940 ( .A1(n1219), .A2(n1186), .ZN(n1217) );
XOR2_X1 U941 ( .A(n1119), .B(KEYINPUT53), .Z(n1219) );
XOR2_X1 U942 ( .A(n1220), .B(n1221), .Z(n1119) );
XOR2_X1 U943 ( .A(n1222), .B(n1223), .Z(n1221) );
XOR2_X1 U944 ( .A(n1224), .B(G125), .Z(n1223) );
NAND2_X1 U945 ( .A1(n1225), .A2(n1028), .ZN(n1224) );
XOR2_X1 U946 ( .A(KEYINPUT54), .B(G224), .Z(n1225) );
NAND2_X1 U947 ( .A1(KEYINPUT31), .A2(n1075), .ZN(n1222) );
XOR2_X1 U948 ( .A(n1226), .B(n1227), .Z(n1075) );
XOR2_X1 U949 ( .A(n1228), .B(n1229), .Z(n1227) );
NOR2_X1 U950 ( .A1(G113), .A2(KEYINPUT57), .ZN(n1228) );
XOR2_X1 U951 ( .A(n1230), .B(n1231), .Z(n1226) );
XNOR2_X1 U952 ( .A(n1178), .B(G116), .ZN(n1231) );
NAND2_X1 U953 ( .A1(n1232), .A2(KEYINPUT29), .ZN(n1230) );
XNOR2_X1 U954 ( .A(KEYINPUT21), .B(G101), .ZN(n1232) );
XNOR2_X1 U955 ( .A(n1073), .B(n1100), .ZN(n1220) );
XOR2_X1 U956 ( .A(n1233), .B(n1234), .Z(n1073) );
XNOR2_X1 U957 ( .A(n1171), .B(G110), .ZN(n1234) );
INV_X1 U958 ( .A(G122), .ZN(n1171) );
XNOR2_X1 U959 ( .A(KEYINPUT26), .B(KEYINPUT10), .ZN(n1233) );
NAND2_X1 U960 ( .A1(n1003), .A2(n1235), .ZN(n1180) );
NAND4_X1 U961 ( .A1(G953), .A2(G902), .A3(n1167), .A4(n1072), .ZN(n1235) );
INV_X1 U962 ( .A(G898), .ZN(n1072) );
NAND3_X1 U963 ( .A1(n1167), .A2(n1028), .A3(G952), .ZN(n1003) );
NAND2_X1 U964 ( .A1(G237), .A2(G234), .ZN(n1167) );
NOR2_X1 U965 ( .A1(n1034), .A2(n1032), .ZN(n1163) );
INV_X1 U966 ( .A(n1185), .ZN(n1032) );
NAND2_X1 U967 ( .A1(G221), .A2(n1236), .ZN(n1185) );
XOR2_X1 U968 ( .A(n1048), .B(G469), .Z(n1034) );
NAND2_X1 U969 ( .A1(n1237), .A2(n1186), .ZN(n1048) );
XOR2_X1 U970 ( .A(n1238), .B(n1239), .Z(n1237) );
XNOR2_X1 U971 ( .A(n1240), .B(n1115), .ZN(n1239) );
XNOR2_X1 U972 ( .A(n1241), .B(n1229), .ZN(n1115) );
XOR2_X1 U973 ( .A(G104), .B(G107), .Z(n1229) );
XNOR2_X1 U974 ( .A(KEYINPUT20), .B(n1242), .ZN(n1241) );
NOR2_X1 U975 ( .A1(KEYINPUT55), .A2(n1243), .ZN(n1242) );
XOR2_X1 U976 ( .A(KEYINPUT21), .B(G101), .Z(n1243) );
XOR2_X1 U977 ( .A(n1244), .B(n1245), .Z(n1238) );
NOR2_X1 U978 ( .A1(KEYINPUT37), .A2(n1059), .ZN(n1245) );
NAND3_X1 U979 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1059) );
NAND2_X1 U980 ( .A1(KEYINPUT7), .A2(n1249), .ZN(n1248) );
NAND3_X1 U981 ( .A1(n1250), .A2(n1251), .A3(n1212), .ZN(n1247) );
INV_X1 U982 ( .A(KEYINPUT7), .ZN(n1251) );
OR2_X1 U983 ( .A1(n1212), .A2(n1250), .ZN(n1246) );
NOR2_X1 U984 ( .A1(KEYINPUT30), .A2(n1249), .ZN(n1250) );
XNOR2_X1 U985 ( .A(G146), .B(G143), .ZN(n1249) );
NAND2_X1 U986 ( .A1(n1252), .A2(n1253), .ZN(n1244) );
XOR2_X1 U987 ( .A(n1254), .B(n1112), .Z(n1253) );
AND2_X1 U988 ( .A1(G227), .A2(n1028), .ZN(n1112) );
NAND3_X1 U989 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1254) );
NAND2_X1 U990 ( .A1(G140), .A2(n1108), .ZN(n1257) );
INV_X1 U991 ( .A(G110), .ZN(n1108) );
NAND2_X1 U992 ( .A1(n1258), .A2(n1259), .ZN(n1256) );
INV_X1 U993 ( .A(KEYINPUT32), .ZN(n1259) );
NAND2_X1 U994 ( .A1(n1260), .A2(n1116), .ZN(n1258) );
XNOR2_X1 U995 ( .A(KEYINPUT40), .B(G110), .ZN(n1260) );
NAND2_X1 U996 ( .A1(KEYINPUT32), .A2(n1261), .ZN(n1255) );
NAND2_X1 U997 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
OR2_X1 U998 ( .A1(G110), .A2(KEYINPUT40), .ZN(n1263) );
NAND3_X1 U999 ( .A1(G110), .A2(n1116), .A3(KEYINPUT40), .ZN(n1262) );
XNOR2_X1 U1000 ( .A(KEYINPUT62), .B(KEYINPUT18), .ZN(n1252) );
INV_X1 U1001 ( .A(n1020), .ZN(n1139) );
NAND2_X1 U1002 ( .A1(n1179), .A2(n1041), .ZN(n1020) );
XOR2_X1 U1003 ( .A(n1264), .B(n1082), .Z(n1041) );
NAND2_X1 U1004 ( .A1(G217), .A2(n1236), .ZN(n1082) );
NAND2_X1 U1005 ( .A1(G234), .A2(n1186), .ZN(n1236) );
OR2_X1 U1006 ( .A1(n1081), .A2(G902), .ZN(n1264) );
XNOR2_X1 U1007 ( .A(n1265), .B(n1266), .ZN(n1081) );
XNOR2_X1 U1008 ( .A(n1191), .B(n1267), .ZN(n1266) );
XOR2_X1 U1009 ( .A(n1268), .B(n1269), .Z(n1267) );
NOR2_X1 U1010 ( .A1(KEYINPUT16), .A2(n1270), .ZN(n1269) );
XOR2_X1 U1011 ( .A(n1271), .B(n1212), .Z(n1270) );
XNOR2_X1 U1012 ( .A(G119), .B(G110), .ZN(n1271) );
NAND3_X1 U1013 ( .A1(G234), .A2(n1028), .A3(G221), .ZN(n1268) );
XOR2_X1 U1014 ( .A(G146), .B(n1056), .Z(n1191) );
XNOR2_X1 U1015 ( .A(G125), .B(n1116), .ZN(n1056) );
INV_X1 U1016 ( .A(G140), .ZN(n1116) );
XOR2_X1 U1017 ( .A(n1272), .B(G137), .Z(n1265) );
XNOR2_X1 U1018 ( .A(KEYINPUT5), .B(KEYINPUT22), .ZN(n1272) );
XOR2_X1 U1019 ( .A(n1040), .B(KEYINPUT19), .Z(n1179) );
XNOR2_X1 U1020 ( .A(n1273), .B(G472), .ZN(n1040) );
NAND2_X1 U1021 ( .A1(n1274), .A2(n1186), .ZN(n1273) );
INV_X1 U1022 ( .A(G902), .ZN(n1186) );
XOR2_X1 U1023 ( .A(n1096), .B(n1100), .Z(n1274) );
XOR2_X1 U1024 ( .A(n1275), .B(n1212), .Z(n1100) );
XOR2_X1 U1025 ( .A(G128), .B(KEYINPUT9), .Z(n1212) );
NAND3_X1 U1026 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1275) );
OR2_X1 U1027 ( .A1(n1279), .A2(KEYINPUT28), .ZN(n1278) );
NAND3_X1 U1028 ( .A1(KEYINPUT28), .A2(n1279), .A3(G146), .ZN(n1277) );
NAND2_X1 U1029 ( .A1(n1280), .A2(n1150), .ZN(n1276) );
INV_X1 U1030 ( .A(G146), .ZN(n1150) );
NAND2_X1 U1031 ( .A1(KEYINPUT28), .A2(n1281), .ZN(n1280) );
XNOR2_X1 U1032 ( .A(KEYINPUT48), .B(n1279), .ZN(n1281) );
INV_X1 U1033 ( .A(G143), .ZN(n1279) );
XNOR2_X1 U1034 ( .A(n1282), .B(n1283), .ZN(n1096) );
XNOR2_X1 U1035 ( .A(n1240), .B(n1284), .ZN(n1283) );
XOR2_X1 U1036 ( .A(n1285), .B(n1286), .Z(n1284) );
NOR2_X1 U1037 ( .A1(n1287), .A2(n1193), .ZN(n1286) );
NAND2_X1 U1038 ( .A1(n1028), .A2(n1218), .ZN(n1193) );
INV_X1 U1039 ( .A(G237), .ZN(n1218) );
INV_X1 U1040 ( .A(G953), .ZN(n1028) );
INV_X1 U1041 ( .A(G210), .ZN(n1287) );
NOR2_X1 U1042 ( .A1(KEYINPUT33), .A2(n1288), .ZN(n1285) );
XNOR2_X1 U1043 ( .A(G116), .B(KEYINPUT25), .ZN(n1288) );
INV_X1 U1044 ( .A(n1060), .ZN(n1240) );
XOR2_X1 U1045 ( .A(G131), .B(n1289), .Z(n1060) );
XOR2_X1 U1046 ( .A(G137), .B(G134), .Z(n1289) );
XNOR2_X1 U1047 ( .A(G101), .B(n1290), .ZN(n1282) );
XNOR2_X1 U1048 ( .A(n1178), .B(G113), .ZN(n1290) );
INV_X1 U1049 ( .A(G119), .ZN(n1178) );
endmodule


