//Key = 0011010000011000111100010010000000001000011100011000100001110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365;

XOR2_X1 U757 ( .A(G107), .B(n1045), .Z(G9) );
NOR2_X1 U758 ( .A1(n1046), .A2(n1047), .ZN(G75) );
NOR4_X1 U759 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
INV_X1 U760 ( .A(G952), .ZN(n1050) );
NAND4_X1 U761 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1048) );
NAND3_X1 U762 ( .A1(n1056), .A2(n1057), .A3(KEYINPUT55), .ZN(n1053) );
NAND4_X1 U763 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1057) );
NAND2_X1 U764 ( .A1(n1058), .A2(n1062), .ZN(n1052) );
NAND2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U766 ( .A1(n1065), .A2(n1066), .A3(n1056), .ZN(n1064) );
NAND3_X1 U767 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
NAND2_X1 U768 ( .A1(n1059), .A2(n1070), .ZN(n1069) );
OR2_X1 U769 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U770 ( .A1(n1060), .A2(n1073), .A3(n1074), .ZN(n1068) );
NAND3_X1 U771 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1067) );
XOR2_X1 U772 ( .A(KEYINPUT50), .B(n1060), .Z(n1075) );
NAND3_X1 U773 ( .A1(n1060), .A2(n1078), .A3(n1059), .ZN(n1063) );
NAND2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U775 ( .A1(n1056), .A2(n1081), .ZN(n1080) );
NAND2_X1 U776 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
OR2_X1 U777 ( .A1(n1084), .A2(KEYINPUT55), .ZN(n1083) );
NAND2_X1 U778 ( .A1(n1065), .A2(n1085), .ZN(n1079) );
NAND2_X1 U779 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U780 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
INV_X1 U781 ( .A(n1090), .ZN(n1058) );
NOR3_X1 U782 ( .A1(n1091), .A2(G953), .A3(n1092), .ZN(n1046) );
INV_X1 U783 ( .A(n1054), .ZN(n1092) );
NAND4_X1 U784 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1054) );
NOR4_X1 U785 ( .A1(n1077), .A2(n1088), .A3(n1097), .A4(n1098), .ZN(n1096) );
NOR2_X1 U786 ( .A1(n1099), .A2(n1100), .ZN(n1095) );
XNOR2_X1 U787 ( .A(n1101), .B(n1102), .ZN(n1094) );
XOR2_X1 U788 ( .A(n1103), .B(KEYINPUT33), .Z(n1101) );
XNOR2_X1 U789 ( .A(n1104), .B(n1105), .ZN(n1093) );
XNOR2_X1 U790 ( .A(G952), .B(KEYINPUT12), .ZN(n1091) );
XOR2_X1 U791 ( .A(n1106), .B(n1107), .Z(G72) );
XOR2_X1 U792 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U793 ( .A1(G953), .A2(n1110), .ZN(n1109) );
NAND2_X1 U794 ( .A1(G900), .A2(G227), .ZN(n1110) );
NAND2_X1 U795 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
NAND2_X1 U796 ( .A1(n1113), .A2(G953), .ZN(n1112) );
XOR2_X1 U797 ( .A(n1114), .B(n1115), .Z(n1111) );
XOR2_X1 U798 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U799 ( .A(n1118), .B(n1119), .Z(n1114) );
XNOR2_X1 U800 ( .A(KEYINPUT44), .B(n1120), .ZN(n1119) );
NAND2_X1 U801 ( .A1(KEYINPUT47), .A2(n1121), .ZN(n1118) );
AND2_X1 U802 ( .A1(n1049), .A2(n1055), .ZN(n1106) );
XOR2_X1 U803 ( .A(n1122), .B(n1123), .Z(G69) );
NOR2_X1 U804 ( .A1(n1124), .A2(n1055), .ZN(n1123) );
NOR2_X1 U805 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XNOR2_X1 U806 ( .A(KEYINPUT11), .B(n1127), .ZN(n1126) );
NAND2_X1 U807 ( .A1(n1128), .A2(n1129), .ZN(n1122) );
NAND2_X1 U808 ( .A1(n1130), .A2(n1055), .ZN(n1129) );
XNOR2_X1 U809 ( .A(n1051), .B(n1131), .ZN(n1130) );
OR3_X1 U810 ( .A1(n1127), .A2(n1131), .A3(n1055), .ZN(n1128) );
XNOR2_X1 U811 ( .A(n1132), .B(n1133), .ZN(n1131) );
XNOR2_X1 U812 ( .A(n1134), .B(n1135), .ZN(n1133) );
XNOR2_X1 U813 ( .A(KEYINPUT38), .B(n1136), .ZN(n1132) );
NOR2_X1 U814 ( .A1(KEYINPUT49), .A2(n1137), .ZN(n1136) );
XNOR2_X1 U815 ( .A(n1138), .B(KEYINPUT18), .ZN(n1137) );
NOR2_X1 U816 ( .A1(n1139), .A2(n1140), .ZN(G66) );
XOR2_X1 U817 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U818 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NOR2_X1 U819 ( .A1(n1139), .A2(n1145), .ZN(G63) );
XOR2_X1 U820 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U821 ( .A1(n1148), .A2(n1144), .ZN(n1146) );
NOR2_X1 U822 ( .A1(n1139), .A2(n1149), .ZN(G60) );
XOR2_X1 U823 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR3_X1 U824 ( .A1(n1144), .A2(KEYINPUT30), .A3(n1152), .ZN(n1150) );
XNOR2_X1 U825 ( .A(n1153), .B(n1154), .ZN(G6) );
NOR2_X1 U826 ( .A1(G104), .A2(KEYINPUT25), .ZN(n1154) );
NOR2_X1 U827 ( .A1(n1139), .A2(n1155), .ZN(G57) );
XOR2_X1 U828 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U829 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U830 ( .A1(n1160), .A2(n1144), .ZN(n1159) );
NAND2_X1 U831 ( .A1(KEYINPUT63), .A2(n1161), .ZN(n1158) );
NOR2_X1 U832 ( .A1(n1139), .A2(n1162), .ZN(G54) );
XOR2_X1 U833 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U834 ( .A1(n1105), .A2(n1144), .ZN(n1164) );
INV_X1 U835 ( .A(G469), .ZN(n1105) );
NOR2_X1 U836 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
XOR2_X1 U837 ( .A(KEYINPUT24), .B(n1167), .Z(n1166) );
NOR3_X1 U838 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1167) );
INV_X1 U839 ( .A(n1171), .ZN(n1168) );
NOR2_X1 U840 ( .A1(n1172), .A2(n1171), .ZN(n1165) );
XNOR2_X1 U841 ( .A(n1173), .B(n1174), .ZN(n1171) );
XNOR2_X1 U842 ( .A(n1175), .B(n1176), .ZN(n1174) );
NOR2_X1 U843 ( .A1(G140), .A2(KEYINPUT40), .ZN(n1176) );
XNOR2_X1 U844 ( .A(G110), .B(KEYINPUT46), .ZN(n1173) );
NOR2_X1 U845 ( .A1(n1169), .A2(n1170), .ZN(n1172) );
NOR2_X1 U846 ( .A1(n1139), .A2(n1177), .ZN(G51) );
XOR2_X1 U847 ( .A(n1178), .B(n1179), .Z(n1177) );
XNOR2_X1 U848 ( .A(n1180), .B(n1181), .ZN(n1179) );
NOR2_X1 U849 ( .A1(n1102), .A2(n1144), .ZN(n1181) );
NAND2_X1 U850 ( .A1(G902), .A2(n1182), .ZN(n1144) );
OR2_X1 U851 ( .A1(n1049), .A2(n1051), .ZN(n1182) );
NAND4_X1 U852 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1051) );
NOR4_X1 U853 ( .A1(n1187), .A2(n1188), .A3(n1153), .A4(n1045), .ZN(n1186) );
AND3_X1 U854 ( .A1(n1072), .A2(n1065), .A3(n1189), .ZN(n1045) );
AND3_X1 U855 ( .A1(n1189), .A2(n1065), .A3(n1071), .ZN(n1153) );
NOR3_X1 U856 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1185) );
NOR2_X1 U857 ( .A1(n1086), .A2(n1193), .ZN(n1192) );
NOR4_X1 U858 ( .A1(n1194), .A2(n1195), .A3(KEYINPUT17), .A4(n1196), .ZN(n1191) );
NOR2_X1 U859 ( .A1(n1197), .A2(n1198), .ZN(n1190) );
INV_X1 U860 ( .A(KEYINPUT17), .ZN(n1198) );
NAND4_X1 U861 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1049) );
NOR4_X1 U862 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
INV_X1 U863 ( .A(n1207), .ZN(n1206) );
AND4_X1 U864 ( .A1(n1072), .A2(n1061), .A3(n1208), .A4(n1056), .ZN(n1204) );
INV_X1 U865 ( .A(n1209), .ZN(n1203) );
NOR2_X1 U866 ( .A1(n1210), .A2(n1211), .ZN(n1201) );
AND2_X1 U867 ( .A1(n1212), .A2(n1059), .ZN(n1211) );
XNOR2_X1 U868 ( .A(G125), .B(n1213), .ZN(n1178) );
NOR2_X1 U869 ( .A1(KEYINPUT56), .A2(n1214), .ZN(n1213) );
NOR2_X1 U870 ( .A1(n1055), .A2(G952), .ZN(n1139) );
XNOR2_X1 U871 ( .A(n1215), .B(n1210), .ZN(G48) );
AND2_X1 U872 ( .A1(n1216), .A2(n1217), .ZN(n1210) );
XNOR2_X1 U873 ( .A(G143), .B(n1209), .ZN(G45) );
NAND3_X1 U874 ( .A1(n1208), .A2(n1061), .A3(n1218), .ZN(n1209) );
XNOR2_X1 U875 ( .A(G140), .B(n1199), .ZN(G42) );
NAND2_X1 U876 ( .A1(n1219), .A2(n1220), .ZN(n1199) );
XNOR2_X1 U877 ( .A(G137), .B(n1200), .ZN(G39) );
NAND3_X1 U878 ( .A1(n1217), .A2(n1056), .A3(n1060), .ZN(n1200) );
XNOR2_X1 U879 ( .A(G134), .B(n1221), .ZN(G36) );
NAND4_X1 U880 ( .A1(n1222), .A2(n1208), .A3(n1061), .A4(n1072), .ZN(n1221) );
XNOR2_X1 U881 ( .A(n1056), .B(KEYINPUT41), .ZN(n1222) );
XNOR2_X1 U882 ( .A(G131), .B(n1207), .ZN(G33) );
NAND2_X1 U883 ( .A1(n1220), .A2(n1061), .ZN(n1207) );
AND3_X1 U884 ( .A1(n1056), .A2(n1208), .A3(n1071), .ZN(n1220) );
AND2_X1 U885 ( .A1(n1089), .A2(n1223), .ZN(n1056) );
NAND2_X1 U886 ( .A1(n1224), .A2(n1225), .ZN(G30) );
NAND2_X1 U887 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
XOR2_X1 U888 ( .A(KEYINPUT45), .B(n1205), .Z(n1226) );
NAND2_X1 U889 ( .A1(n1228), .A2(G128), .ZN(n1224) );
XOR2_X1 U890 ( .A(KEYINPUT19), .B(n1205), .Z(n1228) );
AND3_X1 U891 ( .A1(n1072), .A2(n1194), .A3(n1217), .ZN(n1205) );
AND3_X1 U892 ( .A1(n1208), .A2(n1099), .A3(n1229), .ZN(n1217) );
AND3_X1 U893 ( .A1(n1230), .A2(n1074), .A3(n1073), .ZN(n1208) );
XOR2_X1 U894 ( .A(n1188), .B(n1231), .Z(G3) );
NOR2_X1 U895 ( .A1(KEYINPUT13), .A2(n1232), .ZN(n1231) );
AND3_X1 U896 ( .A1(n1061), .A2(n1189), .A3(n1060), .ZN(n1188) );
XOR2_X1 U897 ( .A(n1233), .B(n1234), .Z(G27) );
NOR2_X1 U898 ( .A1(G125), .A2(KEYINPUT53), .ZN(n1234) );
NAND2_X1 U899 ( .A1(n1212), .A2(n1235), .ZN(n1233) );
XOR2_X1 U900 ( .A(KEYINPUT28), .B(n1059), .Z(n1235) );
AND3_X1 U901 ( .A1(n1219), .A2(n1230), .A3(n1216), .ZN(n1212) );
NAND2_X1 U902 ( .A1(n1236), .A2(n1090), .ZN(n1230) );
NAND2_X1 U903 ( .A1(n1113), .A2(n1237), .ZN(n1236) );
XNOR2_X1 U904 ( .A(G900), .B(KEYINPUT10), .ZN(n1113) );
XNOR2_X1 U905 ( .A(G122), .B(n1183), .ZN(G24) );
NAND3_X1 U906 ( .A1(n1238), .A2(n1065), .A3(n1218), .ZN(n1183) );
NOR3_X1 U907 ( .A1(n1086), .A2(n1239), .A3(n1240), .ZN(n1218) );
AND2_X1 U908 ( .A1(n1241), .A2(n1242), .ZN(n1065) );
XNOR2_X1 U909 ( .A(G119), .B(n1197), .ZN(G21) );
OR3_X1 U910 ( .A1(n1196), .A2(n1086), .A3(n1195), .ZN(n1197) );
NAND3_X1 U911 ( .A1(n1229), .A2(n1099), .A3(n1060), .ZN(n1195) );
INV_X1 U912 ( .A(n1194), .ZN(n1086) );
XNOR2_X1 U913 ( .A(G116), .B(n1243), .ZN(G18) );
NAND2_X1 U914 ( .A1(n1244), .A2(n1194), .ZN(n1243) );
XOR2_X1 U915 ( .A(n1193), .B(KEYINPUT5), .Z(n1244) );
NAND3_X1 U916 ( .A1(n1061), .A2(n1072), .A3(n1238), .ZN(n1193) );
NOR2_X1 U917 ( .A1(n1098), .A2(n1240), .ZN(n1072) );
INV_X1 U918 ( .A(n1245), .ZN(n1240) );
XNOR2_X1 U919 ( .A(n1246), .B(n1184), .ZN(G15) );
NAND3_X1 U920 ( .A1(n1216), .A2(n1061), .A3(n1238), .ZN(n1184) );
INV_X1 U921 ( .A(n1196), .ZN(n1238) );
NAND2_X1 U922 ( .A1(n1059), .A2(n1247), .ZN(n1196) );
NOR2_X1 U923 ( .A1(n1073), .A2(n1077), .ZN(n1059) );
INV_X1 U924 ( .A(n1074), .ZN(n1077) );
INV_X1 U925 ( .A(n1084), .ZN(n1061) );
NAND2_X1 U926 ( .A1(n1241), .A2(n1099), .ZN(n1084) );
XNOR2_X1 U927 ( .A(n1100), .B(KEYINPUT1), .ZN(n1241) );
AND2_X1 U928 ( .A1(n1071), .A2(n1194), .ZN(n1216) );
NOR2_X1 U929 ( .A1(n1245), .A2(n1239), .ZN(n1071) );
INV_X1 U930 ( .A(n1098), .ZN(n1239) );
NAND2_X1 U931 ( .A1(KEYINPUT48), .A2(n1248), .ZN(n1246) );
XNOR2_X1 U932 ( .A(n1249), .B(n1187), .ZN(G12) );
AND3_X1 U933 ( .A1(n1060), .A2(n1189), .A3(n1219), .ZN(n1187) );
INV_X1 U934 ( .A(n1082), .ZN(n1219) );
NAND2_X1 U935 ( .A1(n1229), .A2(n1242), .ZN(n1082) );
INV_X1 U936 ( .A(n1099), .ZN(n1242) );
XOR2_X1 U937 ( .A(n1250), .B(n1160), .Z(n1099) );
INV_X1 U938 ( .A(G472), .ZN(n1160) );
NAND2_X1 U939 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XOR2_X1 U940 ( .A(n1156), .B(n1161), .Z(n1251) );
AND2_X1 U941 ( .A1(n1253), .A2(n1254), .ZN(n1161) );
NAND2_X1 U942 ( .A1(n1255), .A2(n1248), .ZN(n1254) );
XNOR2_X1 U943 ( .A(n1256), .B(n1257), .ZN(n1255) );
INV_X1 U944 ( .A(G116), .ZN(n1256) );
NAND2_X1 U945 ( .A1(G113), .A2(n1258), .ZN(n1253) );
XNOR2_X1 U946 ( .A(G116), .B(n1257), .ZN(n1258) );
NOR2_X1 U947 ( .A1(G119), .A2(KEYINPUT7), .ZN(n1257) );
XOR2_X1 U948 ( .A(n1259), .B(n1260), .Z(n1156) );
XNOR2_X1 U949 ( .A(n1214), .B(n1261), .ZN(n1260) );
INV_X1 U950 ( .A(n1262), .ZN(n1214) );
XNOR2_X1 U951 ( .A(n1263), .B(n1232), .ZN(n1259) );
NAND2_X1 U952 ( .A1(n1264), .A2(G210), .ZN(n1263) );
XNOR2_X1 U953 ( .A(n1100), .B(KEYINPUT36), .ZN(n1229) );
XNOR2_X1 U954 ( .A(n1143), .B(n1265), .ZN(n1100) );
NOR2_X1 U955 ( .A1(G902), .A2(n1141), .ZN(n1265) );
NAND2_X1 U956 ( .A1(n1266), .A2(n1267), .ZN(n1141) );
NAND2_X1 U957 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND2_X1 U958 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
OR2_X1 U959 ( .A1(n1272), .A2(KEYINPUT8), .ZN(n1271) );
INV_X1 U960 ( .A(KEYINPUT32), .ZN(n1270) );
NAND2_X1 U961 ( .A1(n1272), .A2(n1273), .ZN(n1266) );
NAND2_X1 U962 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
OR2_X1 U963 ( .A1(n1268), .A2(KEYINPUT32), .ZN(n1275) );
XNOR2_X1 U964 ( .A(G137), .B(n1276), .ZN(n1268) );
NOR2_X1 U965 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
INV_X1 U966 ( .A(KEYINPUT8), .ZN(n1274) );
XOR2_X1 U967 ( .A(n1117), .B(n1279), .Z(n1272) );
XNOR2_X1 U968 ( .A(n1215), .B(n1280), .ZN(n1279) );
NOR2_X1 U969 ( .A1(KEYINPUT54), .A2(n1281), .ZN(n1280) );
XOR2_X1 U970 ( .A(n1282), .B(n1283), .Z(n1281) );
XNOR2_X1 U971 ( .A(KEYINPUT61), .B(n1249), .ZN(n1283) );
NAND2_X1 U972 ( .A1(n1284), .A2(n1285), .ZN(n1282) );
NAND2_X1 U973 ( .A1(G119), .A2(n1227), .ZN(n1285) );
XOR2_X1 U974 ( .A(KEYINPUT26), .B(n1286), .Z(n1284) );
NOR2_X1 U975 ( .A1(G119), .A2(n1227), .ZN(n1286) );
NAND2_X1 U976 ( .A1(G217), .A2(n1287), .ZN(n1143) );
AND4_X1 U977 ( .A1(n1073), .A2(n1194), .A3(n1247), .A4(n1074), .ZN(n1189) );
NAND2_X1 U978 ( .A1(n1288), .A2(n1287), .ZN(n1074) );
NAND2_X1 U979 ( .A1(G234), .A2(n1252), .ZN(n1287) );
XNOR2_X1 U980 ( .A(KEYINPUT15), .B(n1277), .ZN(n1288) );
INV_X1 U981 ( .A(G221), .ZN(n1277) );
NAND2_X1 U982 ( .A1(n1090), .A2(n1289), .ZN(n1247) );
NAND2_X1 U983 ( .A1(n1237), .A2(n1127), .ZN(n1289) );
INV_X1 U984 ( .A(G898), .ZN(n1127) );
AND3_X1 U985 ( .A1(n1290), .A2(n1291), .A3(G953), .ZN(n1237) );
XNOR2_X1 U986 ( .A(KEYINPUT22), .B(n1252), .ZN(n1290) );
NAND3_X1 U987 ( .A1(n1291), .A2(n1055), .A3(G952), .ZN(n1090) );
NAND2_X1 U988 ( .A1(G237), .A2(G234), .ZN(n1291) );
NOR2_X1 U989 ( .A1(n1089), .A2(n1088), .ZN(n1194) );
INV_X1 U990 ( .A(n1223), .ZN(n1088) );
NAND2_X1 U991 ( .A1(G214), .A2(n1292), .ZN(n1223) );
XNOR2_X1 U992 ( .A(n1103), .B(n1293), .ZN(n1089) );
NOR2_X1 U993 ( .A1(n1294), .A2(KEYINPUT4), .ZN(n1293) );
INV_X1 U994 ( .A(n1102), .ZN(n1294) );
NAND2_X1 U995 ( .A1(G210), .A2(n1292), .ZN(n1102) );
NAND2_X1 U996 ( .A1(n1295), .A2(n1252), .ZN(n1292) );
INV_X1 U997 ( .A(G237), .ZN(n1295) );
NAND2_X1 U998 ( .A1(n1296), .A2(n1252), .ZN(n1103) );
XNOR2_X1 U999 ( .A(n1297), .B(n1298), .ZN(n1296) );
XNOR2_X1 U1000 ( .A(n1299), .B(n1262), .ZN(n1298) );
XOR2_X1 U1001 ( .A(n1300), .B(n1227), .Z(n1262) );
NAND2_X1 U1002 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U1003 ( .A1(n1303), .A2(n1215), .ZN(n1302) );
XOR2_X1 U1004 ( .A(KEYINPUT9), .B(n1304), .Z(n1303) );
XNOR2_X1 U1005 ( .A(n1305), .B(KEYINPUT14), .ZN(n1301) );
NAND2_X1 U1006 ( .A1(KEYINPUT62), .A2(n1306), .ZN(n1299) );
INV_X1 U1007 ( .A(G125), .ZN(n1306) );
INV_X1 U1008 ( .A(n1180), .ZN(n1297) );
XNOR2_X1 U1009 ( .A(n1307), .B(n1308), .ZN(n1180) );
NOR2_X1 U1010 ( .A1(G953), .A2(n1125), .ZN(n1308) );
INV_X1 U1011 ( .A(G224), .ZN(n1125) );
NAND2_X1 U1012 ( .A1(n1309), .A2(n1310), .ZN(n1307) );
NAND2_X1 U1013 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U1014 ( .A(KEYINPUT21), .B(n1134), .Z(n1312) );
XNOR2_X1 U1015 ( .A(n1313), .B(n1138), .ZN(n1311) );
NAND2_X1 U1016 ( .A1(n1314), .A2(n1315), .ZN(n1309) );
XNOR2_X1 U1017 ( .A(n1135), .B(n1138), .ZN(n1315) );
XOR2_X1 U1018 ( .A(G113), .B(n1316), .Z(n1138) );
NOR2_X1 U1019 ( .A1(KEYINPUT60), .A2(n1317), .ZN(n1316) );
XOR2_X1 U1020 ( .A(n1318), .B(G119), .Z(n1317) );
NAND2_X1 U1021 ( .A1(KEYINPUT57), .A2(G116), .ZN(n1318) );
INV_X1 U1022 ( .A(n1313), .ZN(n1135) );
XNOR2_X1 U1023 ( .A(n1319), .B(n1320), .ZN(n1313) );
XNOR2_X1 U1024 ( .A(KEYINPUT2), .B(n1232), .ZN(n1320) );
NAND2_X1 U1025 ( .A1(KEYINPUT58), .A2(n1321), .ZN(n1319) );
XNOR2_X1 U1026 ( .A(n1134), .B(KEYINPUT31), .ZN(n1314) );
XNOR2_X1 U1027 ( .A(n1249), .B(G122), .ZN(n1134) );
INV_X1 U1028 ( .A(n1076), .ZN(n1073) );
XNOR2_X1 U1029 ( .A(n1104), .B(n1322), .ZN(n1076) );
XOR2_X1 U1030 ( .A(KEYINPUT34), .B(n1323), .Z(n1322) );
NOR2_X1 U1031 ( .A1(KEYINPUT20), .A2(G469), .ZN(n1323) );
NAND2_X1 U1032 ( .A1(n1324), .A2(n1252), .ZN(n1104) );
INV_X1 U1033 ( .A(G902), .ZN(n1252) );
XOR2_X1 U1034 ( .A(n1175), .B(n1325), .Z(n1324) );
XOR2_X1 U1035 ( .A(n1326), .B(n1327), .Z(n1325) );
NOR2_X1 U1036 ( .A1(n1169), .A2(n1328), .ZN(n1327) );
XNOR2_X1 U1037 ( .A(n1170), .B(KEYINPUT43), .ZN(n1328) );
AND2_X1 U1038 ( .A1(n1329), .A2(n1261), .ZN(n1170) );
NOR2_X1 U1039 ( .A1(n1261), .A2(n1329), .ZN(n1169) );
XOR2_X1 U1040 ( .A(n1330), .B(n1331), .Z(n1329) );
XNOR2_X1 U1041 ( .A(KEYINPUT59), .B(n1232), .ZN(n1331) );
INV_X1 U1042 ( .A(G101), .ZN(n1232) );
XOR2_X1 U1043 ( .A(n1116), .B(n1332), .Z(n1330) );
NOR2_X1 U1044 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
NOR3_X1 U1045 ( .A1(KEYINPUT23), .A2(G107), .A3(n1335), .ZN(n1334) );
NOR2_X1 U1046 ( .A1(n1321), .A2(n1336), .ZN(n1333) );
INV_X1 U1047 ( .A(KEYINPUT23), .ZN(n1336) );
XNOR2_X1 U1048 ( .A(n1335), .B(G107), .ZN(n1321) );
XOR2_X1 U1049 ( .A(n1337), .B(n1338), .Z(n1116) );
NOR2_X1 U1050 ( .A1(G128), .A2(KEYINPUT29), .ZN(n1338) );
NAND2_X1 U1051 ( .A1(n1339), .A2(n1340), .ZN(n1337) );
NAND2_X1 U1052 ( .A1(n1341), .A2(n1215), .ZN(n1340) );
XOR2_X1 U1053 ( .A(KEYINPUT39), .B(n1304), .Z(n1341) );
XOR2_X1 U1054 ( .A(KEYINPUT42), .B(n1305), .Z(n1339) );
NOR2_X1 U1055 ( .A1(n1215), .A2(n1304), .ZN(n1305) );
XOR2_X1 U1056 ( .A(G143), .B(KEYINPUT51), .Z(n1304) );
INV_X1 U1057 ( .A(G146), .ZN(n1215) );
XNOR2_X1 U1058 ( .A(G131), .B(n1121), .ZN(n1261) );
XNOR2_X1 U1059 ( .A(G134), .B(G137), .ZN(n1121) );
NAND2_X1 U1060 ( .A1(KEYINPUT3), .A2(n1342), .ZN(n1326) );
XNOR2_X1 U1061 ( .A(G140), .B(n1249), .ZN(n1342) );
NAND2_X1 U1062 ( .A1(G227), .A2(n1055), .ZN(n1175) );
NOR2_X1 U1063 ( .A1(n1245), .A2(n1098), .ZN(n1060) );
XOR2_X1 U1064 ( .A(n1343), .B(n1152), .Z(n1098) );
INV_X1 U1065 ( .A(G475), .ZN(n1152) );
OR2_X1 U1066 ( .A1(n1151), .A2(G902), .ZN(n1343) );
XNOR2_X1 U1067 ( .A(n1344), .B(n1345), .ZN(n1151) );
XNOR2_X1 U1068 ( .A(n1248), .B(n1346), .ZN(n1345) );
XNOR2_X1 U1069 ( .A(n1120), .B(G122), .ZN(n1346) );
INV_X1 U1070 ( .A(G131), .ZN(n1120) );
INV_X1 U1071 ( .A(G113), .ZN(n1248) );
XOR2_X1 U1072 ( .A(n1347), .B(n1348), .Z(n1344) );
XNOR2_X1 U1073 ( .A(n1335), .B(n1349), .ZN(n1348) );
NOR2_X1 U1074 ( .A1(KEYINPUT35), .A2(n1350), .ZN(n1349) );
XNOR2_X1 U1075 ( .A(n1351), .B(n1117), .ZN(n1350) );
XOR2_X1 U1076 ( .A(G125), .B(G140), .Z(n1117) );
NAND2_X1 U1077 ( .A1(KEYINPUT52), .A2(G146), .ZN(n1351) );
INV_X1 U1078 ( .A(G104), .ZN(n1335) );
NAND2_X1 U1079 ( .A1(KEYINPUT16), .A2(n1352), .ZN(n1347) );
XNOR2_X1 U1080 ( .A(G143), .B(n1353), .ZN(n1352) );
NAND2_X1 U1081 ( .A1(n1264), .A2(G214), .ZN(n1353) );
NOR2_X1 U1082 ( .A1(G953), .A2(G237), .ZN(n1264) );
XOR2_X1 U1083 ( .A(n1097), .B(KEYINPUT37), .Z(n1245) );
XOR2_X1 U1084 ( .A(n1354), .B(n1148), .Z(n1097) );
INV_X1 U1085 ( .A(G478), .ZN(n1148) );
OR2_X1 U1086 ( .A1(n1147), .A2(G902), .ZN(n1354) );
XNOR2_X1 U1087 ( .A(n1355), .B(n1356), .ZN(n1147) );
XOR2_X1 U1088 ( .A(n1357), .B(n1358), .Z(n1356) );
XNOR2_X1 U1089 ( .A(G134), .B(n1227), .ZN(n1358) );
INV_X1 U1090 ( .A(G128), .ZN(n1227) );
XNOR2_X1 U1091 ( .A(KEYINPUT6), .B(n1359), .ZN(n1357) );
INV_X1 U1092 ( .A(G143), .ZN(n1359) );
XOR2_X1 U1093 ( .A(n1360), .B(n1361), .Z(n1355) );
XOR2_X1 U1094 ( .A(n1362), .B(n1363), .Z(n1361) );
NOR2_X1 U1095 ( .A1(n1278), .A2(n1364), .ZN(n1363) );
INV_X1 U1096 ( .A(G217), .ZN(n1364) );
NAND2_X1 U1097 ( .A1(n1365), .A2(n1055), .ZN(n1278) );
INV_X1 U1098 ( .A(G953), .ZN(n1055) );
XOR2_X1 U1099 ( .A(KEYINPUT0), .B(G234), .Z(n1365) );
NOR2_X1 U1100 ( .A1(G122), .A2(KEYINPUT27), .ZN(n1362) );
XNOR2_X1 U1101 ( .A(G107), .B(G116), .ZN(n1360) );
INV_X1 U1102 ( .A(G110), .ZN(n1249) );
endmodule


