//Key = 0000001101111000100100111000001001110111001010110000100111001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369;

XOR2_X1 U750 ( .A(G107), .B(n1038), .Z(G9) );
NOR2_X1 U751 ( .A1(n1039), .A2(n1040), .ZN(G75) );
NOR4_X1 U752 ( .A1(G953), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1040) );
NOR2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U754 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR4_X1 U755 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
NOR3_X1 U756 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1049) );
NOR2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U758 ( .A1(n1057), .A2(n1058), .ZN(n1053) );
NOR2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U760 ( .A1(n1061), .A2(n1062), .ZN(n1048) );
NOR2_X1 U761 ( .A1(n1063), .A2(n1056), .ZN(n1061) );
NOR4_X1 U762 ( .A1(n1064), .A2(n1058), .A3(n1056), .A4(n1052), .ZN(n1046) );
NOR3_X1 U763 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NOR2_X1 U764 ( .A1(n1068), .A2(n1050), .ZN(n1067) );
NOR2_X1 U765 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NOR2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
AND3_X1 U767 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1066) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1065) );
XNOR2_X1 U769 ( .A(n1073), .B(KEYINPUT49), .ZN(n1076) );
NOR3_X1 U770 ( .A1(n1041), .A2(G953), .A3(G952), .ZN(n1039) );
AND4_X1 U771 ( .A1(n1078), .A2(n1073), .A3(n1079), .A4(n1080), .ZN(n1041) );
NOR4_X1 U772 ( .A1(n1081), .A2(n1063), .A3(n1082), .A4(n1083), .ZN(n1080) );
XNOR2_X1 U773 ( .A(n1084), .B(n1085), .ZN(n1083) );
NOR2_X1 U774 ( .A1(G478), .A2(KEYINPUT40), .ZN(n1085) );
AND2_X1 U775 ( .A1(n1086), .A2(G475), .ZN(n1082) );
NOR2_X1 U776 ( .A1(n1087), .A2(n1052), .ZN(n1079) );
XNOR2_X1 U777 ( .A(n1074), .B(KEYINPUT63), .ZN(n1087) );
XNOR2_X1 U778 ( .A(n1088), .B(G472), .ZN(n1078) );
XOR2_X1 U779 ( .A(n1089), .B(n1090), .Z(G72) );
XOR2_X1 U780 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U781 ( .A1(G953), .A2(n1093), .ZN(n1092) );
NAND2_X1 U782 ( .A1(G900), .A2(G227), .ZN(n1093) );
NAND2_X1 U783 ( .A1(n1094), .A2(n1095), .ZN(n1091) );
NAND2_X1 U784 ( .A1(G953), .A2(n1096), .ZN(n1095) );
XNOR2_X1 U785 ( .A(n1097), .B(n1098), .ZN(n1094) );
NAND3_X1 U786 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1097) );
NAND2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
OR3_X1 U788 ( .A1(n1103), .A2(n1102), .A3(KEYINPUT25), .ZN(n1100) );
NAND2_X1 U789 ( .A1(KEYINPUT9), .A2(n1104), .ZN(n1103) );
NAND2_X1 U790 ( .A1(n1105), .A2(KEYINPUT25), .ZN(n1099) );
INV_X1 U791 ( .A(n1104), .ZN(n1105) );
XOR2_X1 U792 ( .A(n1106), .B(n1107), .Z(n1104) );
XNOR2_X1 U793 ( .A(n1108), .B(G134), .ZN(n1107) );
NAND2_X1 U794 ( .A1(KEYINPUT34), .A2(G131), .ZN(n1106) );
NOR2_X1 U795 ( .A1(n1109), .A2(G953), .ZN(n1089) );
NAND2_X1 U796 ( .A1(n1110), .A2(n1111), .ZN(G69) );
NAND2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U798 ( .A1(G953), .A2(n1114), .ZN(n1113) );
NAND3_X1 U799 ( .A1(n1115), .A2(n1116), .A3(G953), .ZN(n1110) );
NAND2_X1 U800 ( .A1(G898), .A2(G224), .ZN(n1116) );
XOR2_X1 U801 ( .A(KEYINPUT38), .B(n1112), .Z(n1115) );
XNOR2_X1 U802 ( .A(n1117), .B(n1118), .ZN(n1112) );
NOR2_X1 U803 ( .A1(n1119), .A2(G953), .ZN(n1118) );
NAND2_X1 U804 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
INV_X1 U805 ( .A(n1122), .ZN(n1121) );
XNOR2_X1 U806 ( .A(n1123), .B(n1124), .ZN(n1120) );
XNOR2_X1 U807 ( .A(n1125), .B(n1126), .ZN(n1124) );
NOR2_X1 U808 ( .A1(KEYINPUT29), .A2(n1127), .ZN(n1126) );
NOR3_X1 U809 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(G66) );
AND3_X1 U810 ( .A1(KEYINPUT14), .A2(G953), .A3(G952), .ZN(n1130) );
NOR2_X1 U811 ( .A1(KEYINPUT14), .A2(n1131), .ZN(n1129) );
INV_X1 U812 ( .A(n1132), .ZN(n1131) );
NOR2_X1 U813 ( .A1(n1133), .A2(n1134), .ZN(n1128) );
XOR2_X1 U814 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U815 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U816 ( .A1(KEYINPUT17), .A2(n1139), .ZN(n1135) );
AND2_X1 U817 ( .A1(n1139), .A2(KEYINPUT17), .ZN(n1133) );
NOR2_X1 U818 ( .A1(n1132), .A2(n1140), .ZN(G63) );
NOR3_X1 U819 ( .A1(n1084), .A2(n1141), .A3(n1142), .ZN(n1140) );
NOR2_X1 U820 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
AND2_X1 U821 ( .A1(n1043), .A2(G478), .ZN(n1143) );
AND3_X1 U822 ( .A1(n1144), .A2(G478), .A3(n1145), .ZN(n1141) );
NOR2_X1 U823 ( .A1(n1132), .A2(n1146), .ZN(G60) );
XOR2_X1 U824 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U825 ( .A1(n1149), .A2(KEYINPUT4), .ZN(n1148) );
AND2_X1 U826 ( .A1(G475), .A2(n1145), .ZN(n1149) );
NAND2_X1 U827 ( .A1(n1150), .A2(n1151), .ZN(G6) );
NAND2_X1 U828 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XNOR2_X1 U829 ( .A(KEYINPUT8), .B(n1154), .ZN(n1152) );
NAND2_X1 U830 ( .A1(G104), .A2(n1155), .ZN(n1150) );
XOR2_X1 U831 ( .A(n1154), .B(KEYINPUT48), .Z(n1155) );
NOR2_X1 U832 ( .A1(n1132), .A2(n1156), .ZN(G57) );
XOR2_X1 U833 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U834 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U835 ( .A1(KEYINPUT59), .A2(n1161), .ZN(n1160) );
XOR2_X1 U836 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U837 ( .A1(n1145), .A2(G472), .ZN(n1163) );
NAND2_X1 U838 ( .A1(n1164), .A2(KEYINPUT52), .ZN(n1162) );
XNOR2_X1 U839 ( .A(n1165), .B(n1166), .ZN(n1164) );
NOR2_X1 U840 ( .A1(G101), .A2(KEYINPUT31), .ZN(n1157) );
NOR2_X1 U841 ( .A1(n1132), .A2(n1167), .ZN(G54) );
XOR2_X1 U842 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U844 ( .A1(KEYINPUT20), .A2(n1172), .ZN(n1171) );
NAND2_X1 U845 ( .A1(KEYINPUT7), .A2(n1173), .ZN(n1170) );
XOR2_X1 U846 ( .A(n1174), .B(n1175), .Z(n1168) );
AND2_X1 U847 ( .A1(G469), .A2(n1145), .ZN(n1175) );
INV_X1 U848 ( .A(n1138), .ZN(n1145) );
NAND3_X1 U849 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1174) );
NAND2_X1 U850 ( .A1(KEYINPUT15), .A2(n1127), .ZN(n1178) );
OR3_X1 U851 ( .A1(n1179), .A2(KEYINPUT15), .A3(n1102), .ZN(n1177) );
NAND2_X1 U852 ( .A1(n1102), .A2(n1179), .ZN(n1176) );
NAND2_X1 U853 ( .A1(KEYINPUT46), .A2(n1180), .ZN(n1179) );
NOR2_X1 U854 ( .A1(n1132), .A2(n1181), .ZN(G51) );
XOR2_X1 U855 ( .A(n1182), .B(n1183), .Z(n1181) );
NOR2_X1 U856 ( .A1(n1184), .A2(n1138), .ZN(n1183) );
NAND2_X1 U857 ( .A1(G902), .A2(n1043), .ZN(n1138) );
NAND2_X1 U858 ( .A1(n1109), .A2(n1119), .ZN(n1043) );
AND4_X1 U859 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1119) );
NOR4_X1 U860 ( .A1(n1189), .A2(n1190), .A3(n1038), .A4(n1191), .ZN(n1188) );
NOR2_X1 U861 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NOR3_X1 U862 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1192) );
NOR3_X1 U863 ( .A1(n1197), .A2(n1198), .A3(n1077), .ZN(n1196) );
XOR2_X1 U864 ( .A(KEYINPUT50), .B(n1199), .Z(n1194) );
NOR3_X1 U865 ( .A1(n1198), .A2(n1050), .A3(n1200), .ZN(n1038) );
INV_X1 U866 ( .A(n1201), .ZN(n1050) );
AND4_X1 U867 ( .A1(KEYINPUT1), .A2(n1202), .A3(n1203), .A4(n1201), .ZN(n1190) );
NOR2_X1 U868 ( .A1(KEYINPUT1), .A2(n1154), .ZN(n1189) );
NAND3_X1 U869 ( .A1(n1202), .A2(n1201), .A3(n1060), .ZN(n1154) );
AND4_X1 U870 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1109) );
AND4_X1 U871 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1207) );
NAND2_X1 U872 ( .A1(n1060), .A2(n1212), .ZN(n1206) );
NAND2_X1 U873 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
OR2_X1 U874 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND3_X1 U875 ( .A1(n1217), .A2(n1218), .A3(n1059), .ZN(n1204) );
OR2_X1 U876 ( .A1(n1219), .A2(KEYINPUT0), .ZN(n1218) );
NAND2_X1 U877 ( .A1(KEYINPUT0), .A2(n1220), .ZN(n1217) );
NAND2_X1 U878 ( .A1(n1221), .A2(n1077), .ZN(n1220) );
NOR2_X1 U879 ( .A1(n1222), .A2(G952), .ZN(n1132) );
XOR2_X1 U880 ( .A(G146), .B(n1223), .Z(G48) );
NOR3_X1 U881 ( .A1(n1224), .A2(n1203), .A3(n1215), .ZN(n1223) );
XOR2_X1 U882 ( .A(KEYINPUT41), .B(n1216), .Z(n1224) );
NAND2_X1 U883 ( .A1(n1225), .A2(n1226), .ZN(G45) );
OR2_X1 U884 ( .A1(n1205), .A2(G143), .ZN(n1226) );
XOR2_X1 U885 ( .A(n1227), .B(KEYINPUT26), .Z(n1225) );
NAND2_X1 U886 ( .A1(G143), .A2(n1205), .ZN(n1227) );
NAND3_X1 U887 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1205) );
NOR3_X1 U888 ( .A1(n1231), .A2(n1232), .A3(n1216), .ZN(n1230) );
XNOR2_X1 U889 ( .A(G140), .B(n1211), .ZN(G42) );
NAND2_X1 U890 ( .A1(n1221), .A2(n1233), .ZN(n1211) );
XNOR2_X1 U891 ( .A(n1108), .B(n1234), .ZN(G39) );
NOR2_X1 U892 ( .A1(KEYINPUT54), .A2(n1210), .ZN(n1234) );
NAND2_X1 U893 ( .A1(n1221), .A2(n1235), .ZN(n1210) );
XNOR2_X1 U894 ( .A(G134), .B(n1236), .ZN(G36) );
NAND2_X1 U895 ( .A1(n1219), .A2(n1059), .ZN(n1236) );
XNOR2_X1 U896 ( .A(G131), .B(n1237), .ZN(G33) );
NAND2_X1 U897 ( .A1(n1219), .A2(n1238), .ZN(n1237) );
XNOR2_X1 U898 ( .A(KEYINPUT2), .B(n1203), .ZN(n1238) );
INV_X1 U899 ( .A(n1213), .ZN(n1219) );
NAND2_X1 U900 ( .A1(n1228), .A2(n1221), .ZN(n1213) );
NOR4_X1 U901 ( .A1(n1051), .A2(n1062), .A3(n1216), .A4(n1063), .ZN(n1221) );
INV_X1 U902 ( .A(n1073), .ZN(n1051) );
NOR2_X1 U903 ( .A1(n1071), .A2(n1239), .ZN(n1073) );
INV_X1 U904 ( .A(n1072), .ZN(n1239) );
XOR2_X1 U905 ( .A(n1209), .B(n1240), .Z(G30) );
NAND2_X1 U906 ( .A1(KEYINPUT23), .A2(G128), .ZN(n1240) );
OR3_X1 U907 ( .A1(n1198), .A2(n1216), .A3(n1215), .ZN(n1209) );
NAND3_X1 U908 ( .A1(n1074), .A2(n1241), .A3(n1229), .ZN(n1215) );
XNOR2_X1 U909 ( .A(G101), .B(n1187), .ZN(G3) );
NAND3_X1 U910 ( .A1(n1242), .A2(n1202), .A3(n1228), .ZN(n1187) );
XNOR2_X1 U911 ( .A(G125), .B(n1208), .ZN(G27) );
NAND3_X1 U912 ( .A1(n1062), .A2(n1233), .A3(n1243), .ZN(n1208) );
NOR3_X1 U913 ( .A1(n1193), .A2(n1216), .A3(n1058), .ZN(n1243) );
AND2_X1 U914 ( .A1(n1244), .A2(n1045), .ZN(n1216) );
XOR2_X1 U915 ( .A(KEYINPUT24), .B(n1245), .Z(n1244) );
AND4_X1 U916 ( .A1(n1096), .A2(n1246), .A3(G953), .A4(G902), .ZN(n1245) );
INV_X1 U917 ( .A(G900), .ZN(n1096) );
AND3_X1 U918 ( .A1(n1075), .A2(n1074), .A3(n1060), .ZN(n1233) );
XNOR2_X1 U919 ( .A(G122), .B(n1185), .ZN(G24) );
NAND3_X1 U920 ( .A1(n1247), .A2(n1201), .A3(n1248), .ZN(n1185) );
NOR3_X1 U921 ( .A1(n1193), .A2(n1232), .A3(n1231), .ZN(n1248) );
NOR2_X1 U922 ( .A1(n1241), .A2(n1074), .ZN(n1201) );
XNOR2_X1 U923 ( .A(G119), .B(n1249), .ZN(G21) );
NAND2_X1 U924 ( .A1(n1199), .A2(n1070), .ZN(n1249) );
AND2_X1 U925 ( .A1(n1247), .A2(n1235), .ZN(n1199) );
AND3_X1 U926 ( .A1(n1074), .A2(n1241), .A3(n1242), .ZN(n1235) );
XOR2_X1 U927 ( .A(n1250), .B(n1251), .Z(G18) );
NOR2_X1 U928 ( .A1(G116), .A2(KEYINPUT43), .ZN(n1251) );
NAND4_X1 U929 ( .A1(n1252), .A2(n1247), .A3(n1059), .A4(n1070), .ZN(n1250) );
INV_X1 U930 ( .A(n1193), .ZN(n1070) );
INV_X1 U931 ( .A(n1198), .ZN(n1059) );
NAND2_X1 U932 ( .A1(n1232), .A2(n1253), .ZN(n1198) );
INV_X1 U933 ( .A(n1197), .ZN(n1247) );
XNOR2_X1 U934 ( .A(n1228), .B(KEYINPUT16), .ZN(n1252) );
XNOR2_X1 U935 ( .A(n1254), .B(n1255), .ZN(G15) );
NOR2_X1 U936 ( .A1(n1256), .A2(n1193), .ZN(n1255) );
XNOR2_X1 U937 ( .A(n1195), .B(KEYINPUT5), .ZN(n1256) );
NOR3_X1 U938 ( .A1(n1077), .A2(n1203), .A3(n1197), .ZN(n1195) );
NAND3_X1 U939 ( .A1(n1257), .A2(n1258), .A3(n1062), .ZN(n1197) );
INV_X1 U940 ( .A(n1058), .ZN(n1257) );
XNOR2_X1 U941 ( .A(n1063), .B(KEYINPUT6), .ZN(n1058) );
INV_X1 U942 ( .A(n1060), .ZN(n1203) );
NOR2_X1 U943 ( .A1(n1253), .A2(n1232), .ZN(n1060) );
INV_X1 U944 ( .A(n1231), .ZN(n1253) );
INV_X1 U945 ( .A(n1228), .ZN(n1077) );
NOR2_X1 U946 ( .A1(n1074), .A2(n1075), .ZN(n1228) );
XOR2_X1 U947 ( .A(n1186), .B(n1259), .Z(G12) );
NAND2_X1 U948 ( .A1(KEYINPUT55), .A2(G110), .ZN(n1259) );
NAND4_X1 U949 ( .A1(n1242), .A2(n1202), .A3(n1075), .A4(n1074), .ZN(n1186) );
XOR2_X1 U950 ( .A(n1260), .B(n1137), .Z(n1074) );
NAND2_X1 U951 ( .A1(G217), .A2(n1261), .ZN(n1137) );
OR2_X1 U952 ( .A1(n1139), .A2(G902), .ZN(n1260) );
XNOR2_X1 U953 ( .A(n1262), .B(n1263), .ZN(n1139) );
XOR2_X1 U954 ( .A(n1264), .B(n1265), .Z(n1263) );
NAND2_X1 U955 ( .A1(KEYINPUT12), .A2(n1266), .ZN(n1265) );
XNOR2_X1 U956 ( .A(KEYINPUT57), .B(n1267), .ZN(n1266) );
NAND2_X1 U957 ( .A1(n1268), .A2(n1269), .ZN(n1264) );
NAND2_X1 U958 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U959 ( .A1(n1272), .A2(G221), .ZN(n1271) );
XNOR2_X1 U960 ( .A(KEYINPUT51), .B(G137), .ZN(n1270) );
XOR2_X1 U961 ( .A(n1273), .B(KEYINPUT18), .Z(n1268) );
NAND3_X1 U962 ( .A1(G221), .A2(n1274), .A3(n1272), .ZN(n1273) );
XNOR2_X1 U963 ( .A(KEYINPUT51), .B(n1108), .ZN(n1274) );
XOR2_X1 U964 ( .A(n1275), .B(n1276), .Z(n1262) );
XOR2_X1 U965 ( .A(G146), .B(G110), .Z(n1276) );
NAND2_X1 U966 ( .A1(n1277), .A2(KEYINPUT60), .ZN(n1275) );
XNOR2_X1 U967 ( .A(n1278), .B(n1279), .ZN(n1277) );
NAND2_X1 U968 ( .A1(KEYINPUT11), .A2(n1280), .ZN(n1278) );
INV_X1 U969 ( .A(n1241), .ZN(n1075) );
XNOR2_X1 U970 ( .A(n1281), .B(G472), .ZN(n1241) );
NAND2_X1 U971 ( .A1(KEYINPUT47), .A2(n1088), .ZN(n1281) );
AND2_X1 U972 ( .A1(n1282), .A2(n1283), .ZN(n1088) );
XOR2_X1 U973 ( .A(n1165), .B(n1284), .Z(n1282) );
XOR2_X1 U974 ( .A(n1285), .B(n1286), .Z(n1284) );
NOR2_X1 U975 ( .A1(KEYINPUT28), .A2(n1166), .ZN(n1286) );
NAND2_X1 U976 ( .A1(n1287), .A2(n1288), .ZN(n1285) );
OR2_X1 U977 ( .A1(n1159), .A2(G101), .ZN(n1288) );
XOR2_X1 U978 ( .A(n1289), .B(KEYINPUT53), .Z(n1287) );
NAND2_X1 U979 ( .A1(n1159), .A2(G101), .ZN(n1289) );
NOR3_X1 U980 ( .A1(G237), .A2(G953), .A3(n1184), .ZN(n1159) );
INV_X1 U981 ( .A(G210), .ZN(n1184) );
XOR2_X1 U982 ( .A(n1290), .B(n1291), .Z(n1165) );
XOR2_X1 U983 ( .A(n1292), .B(n1293), .Z(n1290) );
NAND2_X1 U984 ( .A1(KEYINPUT19), .A2(n1254), .ZN(n1292) );
INV_X1 U985 ( .A(n1200), .ZN(n1202) );
NAND2_X1 U986 ( .A1(n1229), .A2(n1258), .ZN(n1200) );
NAND2_X1 U987 ( .A1(n1045), .A2(n1294), .ZN(n1258) );
NAND3_X1 U988 ( .A1(n1122), .A2(n1246), .A3(G902), .ZN(n1294) );
NOR2_X1 U989 ( .A1(n1222), .A2(G898), .ZN(n1122) );
NAND3_X1 U990 ( .A1(n1246), .A2(n1222), .A3(G952), .ZN(n1045) );
NAND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1246) );
NOR3_X1 U992 ( .A1(n1062), .A2(n1063), .A3(n1193), .ZN(n1229) );
NAND2_X1 U993 ( .A1(n1071), .A2(n1072), .ZN(n1193) );
NAND2_X1 U994 ( .A1(G214), .A2(n1295), .ZN(n1072) );
NAND2_X1 U995 ( .A1(n1296), .A2(n1283), .ZN(n1295) );
NAND2_X1 U996 ( .A1(n1297), .A2(n1298), .ZN(n1071) );
NAND2_X1 U997 ( .A1(G210), .A2(n1299), .ZN(n1298) );
NAND2_X1 U998 ( .A1(n1283), .A2(n1300), .ZN(n1299) );
OR2_X1 U999 ( .A1(n1296), .A2(n1301), .ZN(n1300) );
NAND3_X1 U1000 ( .A1(n1302), .A2(n1283), .A3(n1301), .ZN(n1297) );
XOR2_X1 U1001 ( .A(n1182), .B(KEYINPUT30), .Z(n1301) );
XOR2_X1 U1002 ( .A(n1303), .B(n1304), .Z(n1182) );
XNOR2_X1 U1003 ( .A(n1293), .B(n1305), .ZN(n1304) );
INV_X1 U1004 ( .A(n1123), .ZN(n1305) );
XOR2_X1 U1005 ( .A(G110), .B(n1306), .Z(n1123) );
XNOR2_X1 U1006 ( .A(KEYINPUT61), .B(n1307), .ZN(n1306) );
INV_X1 U1007 ( .A(G122), .ZN(n1307) );
XNOR2_X1 U1008 ( .A(n1308), .B(n1309), .ZN(n1293) );
NAND2_X1 U1009 ( .A1(KEYINPUT10), .A2(G143), .ZN(n1308) );
XOR2_X1 U1010 ( .A(n1310), .B(n1311), .Z(n1303) );
XNOR2_X1 U1011 ( .A(n1312), .B(n1313), .ZN(n1311) );
NOR2_X1 U1012 ( .A1(n1114), .A2(n1314), .ZN(n1313) );
XNOR2_X1 U1013 ( .A(KEYINPUT62), .B(n1222), .ZN(n1314) );
INV_X1 U1014 ( .A(G224), .ZN(n1114) );
INV_X1 U1015 ( .A(G125), .ZN(n1312) );
NAND3_X1 U1016 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n1310) );
NAND2_X1 U1017 ( .A1(KEYINPUT27), .A2(n1125), .ZN(n1317) );
NAND3_X1 U1018 ( .A1(n1318), .A2(n1319), .A3(n1180), .ZN(n1316) );
INV_X1 U1019 ( .A(n1125), .ZN(n1318) );
NAND2_X1 U1020 ( .A1(n1127), .A2(n1320), .ZN(n1315) );
NAND2_X1 U1021 ( .A1(n1321), .A2(n1319), .ZN(n1320) );
INV_X1 U1022 ( .A(KEYINPUT27), .ZN(n1319) );
XNOR2_X1 U1023 ( .A(n1125), .B(KEYINPUT36), .ZN(n1321) );
XNOR2_X1 U1024 ( .A(n1322), .B(n1291), .ZN(n1125) );
XNOR2_X1 U1025 ( .A(G116), .B(n1280), .ZN(n1291) );
INV_X1 U1026 ( .A(G119), .ZN(n1280) );
XNOR2_X1 U1027 ( .A(G113), .B(KEYINPUT3), .ZN(n1322) );
NAND2_X1 U1028 ( .A1(G210), .A2(G237), .ZN(n1302) );
INV_X1 U1029 ( .A(n1055), .ZN(n1063) );
NAND2_X1 U1030 ( .A1(G221), .A2(n1261), .ZN(n1055) );
NAND2_X1 U1031 ( .A1(G234), .A2(n1283), .ZN(n1261) );
INV_X1 U1032 ( .A(n1052), .ZN(n1062) );
XNOR2_X1 U1033 ( .A(n1323), .B(G469), .ZN(n1052) );
NAND2_X1 U1034 ( .A1(n1324), .A2(n1283), .ZN(n1323) );
XNOR2_X1 U1035 ( .A(n1325), .B(n1172), .ZN(n1324) );
XNOR2_X1 U1036 ( .A(n1326), .B(n1327), .ZN(n1172) );
XOR2_X1 U1037 ( .A(G140), .B(G110), .Z(n1327) );
NAND2_X1 U1038 ( .A1(G227), .A2(n1222), .ZN(n1326) );
NAND2_X1 U1039 ( .A1(KEYINPUT42), .A2(n1328), .ZN(n1325) );
XNOR2_X1 U1040 ( .A(n1180), .B(n1329), .ZN(n1328) );
XOR2_X1 U1041 ( .A(n1330), .B(n1102), .Z(n1329) );
XNOR2_X1 U1042 ( .A(n1309), .B(n1331), .ZN(n1102) );
XNOR2_X1 U1043 ( .A(KEYINPUT21), .B(n1332), .ZN(n1331) );
XOR2_X1 U1044 ( .A(G128), .B(n1333), .Z(n1309) );
XOR2_X1 U1045 ( .A(KEYINPUT58), .B(G146), .Z(n1333) );
NAND2_X1 U1046 ( .A1(KEYINPUT22), .A2(n1166), .ZN(n1330) );
INV_X1 U1047 ( .A(n1173), .ZN(n1166) );
XNOR2_X1 U1048 ( .A(n1334), .B(G131), .ZN(n1173) );
NAND3_X1 U1049 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1334) );
NAND2_X1 U1050 ( .A1(G134), .A2(n1108), .ZN(n1337) );
INV_X1 U1051 ( .A(G137), .ZN(n1108) );
NAND2_X1 U1052 ( .A1(n1338), .A2(n1339), .ZN(n1336) );
INV_X1 U1053 ( .A(KEYINPUT33), .ZN(n1339) );
NAND2_X1 U1054 ( .A1(n1340), .A2(n1341), .ZN(n1338) );
XNOR2_X1 U1055 ( .A(KEYINPUT37), .B(G137), .ZN(n1340) );
NAND2_X1 U1056 ( .A1(KEYINPUT33), .A2(n1342), .ZN(n1335) );
NAND2_X1 U1057 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
OR2_X1 U1058 ( .A1(G137), .A2(KEYINPUT37), .ZN(n1344) );
NAND3_X1 U1059 ( .A1(G137), .A2(n1341), .A3(KEYINPUT37), .ZN(n1343) );
INV_X1 U1060 ( .A(n1127), .ZN(n1180) );
XOR2_X1 U1061 ( .A(G101), .B(n1345), .Z(n1127) );
XNOR2_X1 U1062 ( .A(G107), .B(n1153), .ZN(n1345) );
INV_X1 U1063 ( .A(n1056), .ZN(n1242) );
NAND2_X1 U1064 ( .A1(n1231), .A2(n1232), .ZN(n1056) );
NOR2_X1 U1065 ( .A1(n1346), .A2(n1081), .ZN(n1232) );
NOR2_X1 U1066 ( .A1(n1086), .A2(G475), .ZN(n1081) );
AND2_X1 U1067 ( .A1(n1347), .A2(n1086), .ZN(n1346) );
NAND2_X1 U1068 ( .A1(n1147), .A2(n1283), .ZN(n1086) );
INV_X1 U1069 ( .A(G902), .ZN(n1283) );
XOR2_X1 U1070 ( .A(n1348), .B(n1349), .Z(n1147) );
XOR2_X1 U1071 ( .A(n1350), .B(n1351), .Z(n1349) );
XNOR2_X1 U1072 ( .A(n1352), .B(n1353), .ZN(n1351) );
NOR2_X1 U1073 ( .A1(KEYINPUT13), .A2(n1354), .ZN(n1353) );
XOR2_X1 U1074 ( .A(n1355), .B(G146), .Z(n1354) );
NAND2_X1 U1075 ( .A1(KEYINPUT39), .A2(n1267), .ZN(n1355) );
INV_X1 U1076 ( .A(n1098), .ZN(n1267) );
XOR2_X1 U1077 ( .A(G125), .B(G140), .Z(n1098) );
NAND2_X1 U1078 ( .A1(KEYINPUT56), .A2(n1153), .ZN(n1352) );
INV_X1 U1079 ( .A(G104), .ZN(n1153) );
XNOR2_X1 U1080 ( .A(n1254), .B(n1356), .ZN(n1350) );
AND3_X1 U1081 ( .A1(G214), .A2(n1222), .A3(n1296), .ZN(n1356) );
INV_X1 U1082 ( .A(G237), .ZN(n1296) );
INV_X1 U1083 ( .A(G113), .ZN(n1254) );
XOR2_X1 U1084 ( .A(n1357), .B(n1358), .Z(n1348) );
XNOR2_X1 U1085 ( .A(KEYINPUT35), .B(n1332), .ZN(n1358) );
XNOR2_X1 U1086 ( .A(G122), .B(G131), .ZN(n1357) );
XNOR2_X1 U1087 ( .A(G475), .B(KEYINPUT44), .ZN(n1347) );
XNOR2_X1 U1088 ( .A(n1084), .B(G478), .ZN(n1231) );
NOR2_X1 U1089 ( .A1(n1144), .A2(G902), .ZN(n1084) );
XOR2_X1 U1090 ( .A(n1359), .B(n1360), .Z(n1144) );
XNOR2_X1 U1091 ( .A(n1341), .B(G122), .ZN(n1360) );
INV_X1 U1092 ( .A(G134), .ZN(n1341) );
XOR2_X1 U1093 ( .A(n1361), .B(G116), .Z(n1359) );
NAND2_X1 U1094 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
NAND2_X1 U1095 ( .A1(n1364), .A2(n1332), .ZN(n1363) );
INV_X1 U1096 ( .A(G143), .ZN(n1332) );
XNOR2_X1 U1097 ( .A(n1365), .B(KEYINPUT32), .ZN(n1364) );
NAND2_X1 U1098 ( .A1(n1366), .A2(G143), .ZN(n1362) );
XNOR2_X1 U1099 ( .A(KEYINPUT45), .B(n1367), .ZN(n1366) );
INV_X1 U1100 ( .A(n1365), .ZN(n1367) );
XNOR2_X1 U1101 ( .A(n1368), .B(n1369), .ZN(n1365) );
XNOR2_X1 U1102 ( .A(n1279), .B(G107), .ZN(n1369) );
INV_X1 U1103 ( .A(G128), .ZN(n1279) );
NAND2_X1 U1104 ( .A1(G217), .A2(n1272), .ZN(n1368) );
AND2_X1 U1105 ( .A1(G234), .A2(n1222), .ZN(n1272) );
INV_X1 U1106 ( .A(G953), .ZN(n1222) );
endmodule


