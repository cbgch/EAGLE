//Key = 0101010010011101011001001101010100010010101001010000011110001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323;

XOR2_X1 U739 ( .A(G107), .B(n1011), .Z(G9) );
NOR2_X1 U740 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR2_X1 U741 ( .A1(n1014), .A2(n1015), .ZN(G75) );
NOR4_X1 U742 ( .A1(G953), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(n1015) );
NOR2_X1 U743 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR2_X1 U744 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR3_X1 U745 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NOR2_X1 U746 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U747 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR2_X1 U748 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR2_X1 U749 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR3_X1 U750 ( .A1(n1034), .A2(n1035), .A3(n1029), .ZN(n1021) );
INV_X1 U751 ( .A(n1036), .ZN(n1029) );
NOR3_X1 U752 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1035) );
AND3_X1 U753 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
NOR2_X1 U754 ( .A1(n1043), .A2(n1025), .ZN(n1037) );
NOR2_X1 U755 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR3_X1 U756 ( .A1(n1016), .A2(G953), .A3(G952), .ZN(n1014) );
AND4_X1 U757 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1016) );
NOR4_X1 U758 ( .A1(n1050), .A2(n1042), .A3(n1051), .A4(n1052), .ZN(n1049) );
XOR2_X1 U759 ( .A(n1053), .B(n1054), .Z(n1052) );
XNOR2_X1 U760 ( .A(KEYINPUT58), .B(n1055), .ZN(n1053) );
NOR2_X1 U761 ( .A1(KEYINPUT49), .A2(n1056), .ZN(n1055) );
NOR2_X1 U762 ( .A1(n1057), .A2(n1058), .ZN(n1051) );
XNOR2_X1 U763 ( .A(KEYINPUT46), .B(n1059), .ZN(n1058) );
NOR2_X1 U764 ( .A1(n1034), .A2(n1060), .ZN(n1048) );
XOR2_X1 U765 ( .A(n1061), .B(n1062), .Z(n1047) );
XOR2_X1 U766 ( .A(KEYINPUT42), .B(G469), .Z(n1062) );
NAND2_X1 U767 ( .A1(KEYINPUT29), .A2(n1063), .ZN(n1061) );
XNOR2_X1 U768 ( .A(n1064), .B(KEYINPUT7), .ZN(n1046) );
XOR2_X1 U769 ( .A(n1065), .B(n1066), .Z(G72) );
NOR2_X1 U770 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
AND2_X1 U771 ( .A1(G227), .A2(G900), .ZN(n1067) );
NAND2_X1 U772 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
NAND2_X1 U773 ( .A1(n1071), .A2(n1068), .ZN(n1070) );
XNOR2_X1 U774 ( .A(n1072), .B(n1073), .ZN(n1071) );
NAND3_X1 U775 ( .A1(G900), .A2(n1073), .A3(G953), .ZN(n1069) );
XNOR2_X1 U776 ( .A(n1074), .B(n1075), .ZN(n1073) );
XOR2_X1 U777 ( .A(n1076), .B(n1077), .Z(n1075) );
XNOR2_X1 U778 ( .A(KEYINPUT36), .B(n1078), .ZN(n1077) );
NOR2_X1 U779 ( .A1(KEYINPUT28), .A2(n1079), .ZN(n1078) );
NAND2_X1 U780 ( .A1(KEYINPUT3), .A2(n1080), .ZN(n1076) );
XNOR2_X1 U781 ( .A(n1081), .B(n1082), .ZN(n1074) );
XOR2_X1 U782 ( .A(n1083), .B(n1084), .Z(G69) );
NAND2_X1 U783 ( .A1(G953), .A2(n1085), .ZN(n1084) );
NAND2_X1 U784 ( .A1(G898), .A2(G224), .ZN(n1085) );
NAND3_X1 U785 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1083) );
OR2_X1 U786 ( .A1(n1089), .A2(KEYINPUT47), .ZN(n1088) );
NAND3_X1 U787 ( .A1(KEYINPUT47), .A2(n1090), .A3(n1091), .ZN(n1087) );
OR2_X1 U788 ( .A1(n1091), .A2(n1090), .ZN(n1086) );
AND2_X1 U789 ( .A1(KEYINPUT18), .A2(n1089), .ZN(n1090) );
NAND2_X1 U790 ( .A1(n1092), .A2(n1093), .ZN(n1089) );
NAND2_X1 U791 ( .A1(G953), .A2(n1094), .ZN(n1093) );
XOR2_X1 U792 ( .A(n1095), .B(n1096), .Z(n1092) );
XOR2_X1 U793 ( .A(n1097), .B(KEYINPUT33), .Z(n1095) );
NAND2_X1 U794 ( .A1(n1068), .A2(n1098), .ZN(n1091) );
NAND2_X1 U795 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U796 ( .A(KEYINPUT55), .B(n1101), .ZN(n1100) );
NOR2_X1 U797 ( .A1(n1102), .A2(n1103), .ZN(G66) );
XOR2_X1 U798 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U799 ( .A1(KEYINPUT26), .A2(n1106), .ZN(n1105) );
NAND2_X1 U800 ( .A1(n1107), .A2(n1054), .ZN(n1104) );
NOR2_X1 U801 ( .A1(n1102), .A2(n1108), .ZN(G63) );
XNOR2_X1 U802 ( .A(n1109), .B(n1110), .ZN(n1108) );
AND2_X1 U803 ( .A1(G478), .A2(n1107), .ZN(n1110) );
NOR2_X1 U804 ( .A1(n1102), .A2(n1111), .ZN(G60) );
XNOR2_X1 U805 ( .A(n1112), .B(n1113), .ZN(n1111) );
NOR2_X1 U806 ( .A1(n1057), .A2(n1114), .ZN(n1113) );
INV_X1 U807 ( .A(G475), .ZN(n1057) );
XOR2_X1 U808 ( .A(n1115), .B(n1116), .Z(G6) );
XNOR2_X1 U809 ( .A(G104), .B(KEYINPUT0), .ZN(n1116) );
NOR2_X1 U810 ( .A1(n1102), .A2(n1117), .ZN(G57) );
XOR2_X1 U811 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U812 ( .A(G101), .B(n1120), .Z(n1119) );
NOR2_X1 U813 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XNOR2_X1 U814 ( .A(KEYINPUT56), .B(KEYINPUT20), .ZN(n1121) );
XOR2_X1 U815 ( .A(n1123), .B(n1124), .Z(n1118) );
AND2_X1 U816 ( .A1(G472), .A2(n1107), .ZN(n1124) );
INV_X1 U817 ( .A(n1114), .ZN(n1107) );
NOR2_X1 U818 ( .A1(n1102), .A2(n1125), .ZN(G54) );
XOR2_X1 U819 ( .A(n1126), .B(n1127), .Z(n1125) );
XNOR2_X1 U820 ( .A(n1079), .B(n1128), .ZN(n1127) );
XNOR2_X1 U821 ( .A(n1129), .B(n1130), .ZN(n1128) );
NAND2_X1 U822 ( .A1(KEYINPUT15), .A2(n1131), .ZN(n1130) );
NAND2_X1 U823 ( .A1(KEYINPUT12), .A2(n1132), .ZN(n1129) );
XOR2_X1 U824 ( .A(n1133), .B(n1134), .Z(n1126) );
XOR2_X1 U825 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U826 ( .A1(KEYINPUT22), .A2(n1137), .ZN(n1136) );
NOR3_X1 U827 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1135) );
INV_X1 U828 ( .A(G469), .ZN(n1140) );
XOR2_X1 U829 ( .A(n1018), .B(KEYINPUT38), .Z(n1139) );
XOR2_X1 U830 ( .A(n1141), .B(G110), .Z(n1133) );
NOR2_X1 U831 ( .A1(n1102), .A2(n1142), .ZN(G51) );
XOR2_X1 U832 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U833 ( .A1(n1145), .A2(n1114), .ZN(n1143) );
NAND2_X1 U834 ( .A1(G902), .A2(n1018), .ZN(n1114) );
NAND3_X1 U835 ( .A1(n1099), .A2(n1101), .A3(n1072), .ZN(n1018) );
AND4_X1 U836 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1072) );
NOR4_X1 U837 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1149) );
INV_X1 U838 ( .A(n1154), .ZN(n1153) );
INV_X1 U839 ( .A(n1155), .ZN(n1150) );
NAND3_X1 U840 ( .A1(n1156), .A2(n1044), .A3(n1026), .ZN(n1148) );
AND2_X1 U841 ( .A1(n1157), .A2(n1158), .ZN(n1026) );
OR2_X1 U842 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
AND4_X1 U843 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1099) );
AND3_X1 U844 ( .A1(n1115), .A2(n1165), .A3(n1166), .ZN(n1164) );
OR2_X1 U845 ( .A1(n1167), .A2(n1013), .ZN(n1166) );
NOR2_X1 U846 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XNOR2_X1 U847 ( .A(KEYINPUT6), .B(n1012), .ZN(n1169) );
NAND4_X1 U848 ( .A1(n1045), .A2(n1170), .A3(n1036), .A4(n1171), .ZN(n1012) );
NOR3_X1 U849 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1168) );
NAND4_X1 U850 ( .A1(n1036), .A2(n1171), .A3(n1170), .A4(n1175), .ZN(n1115) );
NOR2_X1 U851 ( .A1(n1013), .A2(n1176), .ZN(n1175) );
NOR2_X1 U852 ( .A1(n1177), .A2(G952), .ZN(n1102) );
XOR2_X1 U853 ( .A(KEYINPUT2), .B(n1068), .Z(n1177) );
XOR2_X1 U854 ( .A(n1178), .B(n1146), .Z(G48) );
NAND3_X1 U855 ( .A1(n1044), .A2(n1030), .A3(n1179), .ZN(n1146) );
XOR2_X1 U856 ( .A(n1180), .B(n1147), .Z(G45) );
NAND4_X1 U857 ( .A1(n1181), .A2(n1030), .A3(n1060), .A4(n1182), .ZN(n1147) );
XOR2_X1 U858 ( .A(n1132), .B(n1183), .Z(G42) );
NAND4_X1 U859 ( .A1(n1156), .A2(n1044), .A3(n1157), .A4(n1184), .ZN(n1183) );
XOR2_X1 U860 ( .A(KEYINPUT10), .B(n1159), .Z(n1184) );
XOR2_X1 U861 ( .A(n1080), .B(n1154), .Z(G39) );
NAND3_X1 U862 ( .A1(n1179), .A2(n1157), .A3(n1040), .ZN(n1154) );
XOR2_X1 U863 ( .A(G134), .B(n1152), .Z(G36) );
AND3_X1 U864 ( .A1(n1157), .A2(n1045), .A3(n1181), .ZN(n1152) );
INV_X1 U865 ( .A(n1185), .ZN(n1181) );
XNOR2_X1 U866 ( .A(G131), .B(n1186), .ZN(G33) );
NAND2_X1 U867 ( .A1(n1157), .A2(n1187), .ZN(n1186) );
XOR2_X1 U868 ( .A(KEYINPUT34), .B(n1188), .Z(n1187) );
NOR2_X1 U869 ( .A1(n1176), .A2(n1185), .ZN(n1188) );
NAND2_X1 U870 ( .A1(n1160), .A2(n1156), .ZN(n1185) );
INV_X1 U871 ( .A(n1034), .ZN(n1157) );
NAND2_X1 U872 ( .A1(n1189), .A2(n1033), .ZN(n1034) );
XOR2_X1 U873 ( .A(G128), .B(n1151), .Z(G30) );
AND3_X1 U874 ( .A1(n1030), .A2(n1045), .A3(n1179), .ZN(n1151) );
AND3_X1 U875 ( .A1(n1064), .A2(n1190), .A3(n1156), .ZN(n1179) );
AND2_X1 U876 ( .A1(n1170), .A2(n1191), .ZN(n1156) );
XOR2_X1 U877 ( .A(n1192), .B(n1193), .Z(G3) );
NAND4_X1 U878 ( .A1(n1194), .A2(KEYINPUT63), .A3(n1195), .A4(n1038), .ZN(n1193) );
NOR2_X1 U879 ( .A1(n1013), .A2(n1174), .ZN(n1195) );
XOR2_X1 U880 ( .A(n1171), .B(KEYINPUT4), .Z(n1194) );
XOR2_X1 U881 ( .A(G125), .B(n1196), .Z(G27) );
NOR2_X1 U882 ( .A1(KEYINPUT57), .A2(n1155), .ZN(n1196) );
NAND4_X1 U883 ( .A1(n1044), .A2(n1159), .A3(n1197), .A4(n1198), .ZN(n1155) );
INV_X1 U884 ( .A(n1025), .ZN(n1198) );
AND2_X1 U885 ( .A1(n1191), .A2(n1030), .ZN(n1197) );
NAND2_X1 U886 ( .A1(n1199), .A2(n1200), .ZN(n1191) );
NAND2_X1 U887 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
INV_X1 U888 ( .A(G900), .ZN(n1202) );
XNOR2_X1 U889 ( .A(G122), .B(n1163), .ZN(G24) );
NAND4_X1 U890 ( .A1(n1203), .A2(n1036), .A3(n1060), .A4(n1182), .ZN(n1163) );
INV_X1 U891 ( .A(n1204), .ZN(n1060) );
NOR2_X1 U892 ( .A1(n1190), .A2(n1064), .ZN(n1036) );
NAND2_X1 U893 ( .A1(n1205), .A2(n1206), .ZN(G21) );
NAND2_X1 U894 ( .A1(G119), .A2(n1101), .ZN(n1206) );
XOR2_X1 U895 ( .A(KEYINPUT13), .B(n1207), .Z(n1205) );
NOR2_X1 U896 ( .A1(G119), .A2(n1101), .ZN(n1207) );
NAND4_X1 U897 ( .A1(n1203), .A2(n1040), .A3(n1064), .A4(n1190), .ZN(n1101) );
INV_X1 U898 ( .A(n1208), .ZN(n1190) );
XOR2_X1 U899 ( .A(n1209), .B(n1161), .Z(G18) );
NAND3_X1 U900 ( .A1(n1160), .A2(n1045), .A3(n1203), .ZN(n1161) );
NOR2_X1 U901 ( .A1(n1182), .A2(n1204), .ZN(n1045) );
XOR2_X1 U902 ( .A(n1165), .B(n1210), .Z(G15) );
NAND2_X1 U903 ( .A1(KEYINPUT45), .A2(G113), .ZN(n1210) );
NAND3_X1 U904 ( .A1(n1160), .A2(n1044), .A3(n1203), .ZN(n1165) );
NOR3_X1 U905 ( .A1(n1013), .A2(n1173), .A3(n1025), .ZN(n1203) );
NAND2_X1 U906 ( .A1(n1211), .A2(n1041), .ZN(n1025) );
XOR2_X1 U907 ( .A(KEYINPUT53), .B(n1042), .Z(n1211) );
INV_X1 U908 ( .A(n1171), .ZN(n1173) );
INV_X1 U909 ( .A(n1176), .ZN(n1044) );
NAND2_X1 U910 ( .A1(n1204), .A2(n1182), .ZN(n1176) );
INV_X1 U911 ( .A(n1212), .ZN(n1182) );
INV_X1 U912 ( .A(n1174), .ZN(n1160) );
NAND2_X1 U913 ( .A1(n1208), .A2(n1064), .ZN(n1174) );
NAND2_X1 U914 ( .A1(n1213), .A2(n1214), .ZN(G12) );
OR2_X1 U915 ( .A1(n1162), .A2(G110), .ZN(n1214) );
XOR2_X1 U916 ( .A(n1215), .B(KEYINPUT32), .Z(n1213) );
NAND2_X1 U917 ( .A1(G110), .A2(n1162), .ZN(n1215) );
NAND4_X1 U918 ( .A1(n1038), .A2(n1159), .A3(n1030), .A4(n1171), .ZN(n1162) );
NAND2_X1 U919 ( .A1(n1199), .A2(n1216), .ZN(n1171) );
NAND2_X1 U920 ( .A1(n1201), .A2(n1094), .ZN(n1216) );
INV_X1 U921 ( .A(G898), .ZN(n1094) );
NOR3_X1 U922 ( .A1(n1068), .A2(n1020), .A3(n1138), .ZN(n1201) );
INV_X1 U923 ( .A(n1217), .ZN(n1020) );
NAND3_X1 U924 ( .A1(n1217), .A2(n1068), .A3(G952), .ZN(n1199) );
NAND2_X1 U925 ( .A1(G237), .A2(n1218), .ZN(n1217) );
INV_X1 U926 ( .A(n1013), .ZN(n1030) );
NAND2_X1 U927 ( .A1(n1032), .A2(n1033), .ZN(n1013) );
NAND2_X1 U928 ( .A1(G214), .A2(n1219), .ZN(n1033) );
INV_X1 U929 ( .A(n1189), .ZN(n1032) );
XOR2_X1 U930 ( .A(n1220), .B(n1221), .Z(n1189) );
NOR2_X1 U931 ( .A1(n1222), .A2(n1145), .ZN(n1221) );
INV_X1 U932 ( .A(G210), .ZN(n1145) );
XOR2_X1 U933 ( .A(n1219), .B(KEYINPUT31), .Z(n1222) );
OR2_X1 U934 ( .A1(G902), .A2(G237), .ZN(n1219) );
OR2_X1 U935 ( .A1(n1144), .A2(G902), .ZN(n1220) );
XNOR2_X1 U936 ( .A(n1223), .B(n1224), .ZN(n1144) );
XOR2_X1 U937 ( .A(n1097), .B(n1225), .Z(n1224) );
NAND2_X1 U938 ( .A1(n1226), .A2(n1227), .ZN(n1097) );
NAND2_X1 U939 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
XOR2_X1 U940 ( .A(n1230), .B(G104), .Z(n1228) );
NAND2_X1 U941 ( .A1(n1231), .A2(n1232), .ZN(n1226) );
XOR2_X1 U942 ( .A(G107), .B(G104), .Z(n1232) );
XNOR2_X1 U943 ( .A(n1229), .B(KEYINPUT9), .ZN(n1231) );
XNOR2_X1 U944 ( .A(n1233), .B(G101), .ZN(n1229) );
NAND2_X1 U945 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U946 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U947 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND2_X1 U948 ( .A1(G113), .A2(n1240), .ZN(n1239) );
INV_X1 U949 ( .A(KEYINPUT51), .ZN(n1238) );
NAND2_X1 U950 ( .A1(n1241), .A2(n1242), .ZN(n1234) );
NAND2_X1 U951 ( .A1(n1240), .A2(n1243), .ZN(n1241) );
OR2_X1 U952 ( .A1(n1236), .A2(KEYINPUT51), .ZN(n1243) );
NAND2_X1 U953 ( .A1(n1244), .A2(n1245), .ZN(n1236) );
NAND2_X1 U954 ( .A1(KEYINPUT21), .A2(n1246), .ZN(n1245) );
OR3_X1 U955 ( .A1(n1209), .A2(G119), .A3(KEYINPUT21), .ZN(n1244) );
INV_X1 U956 ( .A(KEYINPUT50), .ZN(n1240) );
XOR2_X1 U957 ( .A(n1247), .B(n1248), .Z(n1223) );
XOR2_X1 U958 ( .A(G125), .B(n1249), .Z(n1248) );
NOR2_X1 U959 ( .A1(KEYINPUT48), .A2(n1096), .ZN(n1249) );
XOR2_X1 U960 ( .A(G122), .B(G110), .Z(n1096) );
NAND2_X1 U961 ( .A1(G224), .A2(n1068), .ZN(n1247) );
NOR2_X1 U962 ( .A1(n1064), .A2(n1208), .ZN(n1159) );
XNOR2_X1 U963 ( .A(n1056), .B(n1054), .ZN(n1208) );
AND2_X1 U964 ( .A1(G217), .A2(n1250), .ZN(n1054) );
NOR2_X1 U965 ( .A1(n1106), .A2(G902), .ZN(n1056) );
XNOR2_X1 U966 ( .A(n1251), .B(n1252), .ZN(n1106) );
XOR2_X1 U967 ( .A(n1253), .B(n1254), .Z(n1252) );
XNOR2_X1 U968 ( .A(n1255), .B(n1256), .ZN(n1254) );
NOR2_X1 U969 ( .A1(KEYINPUT19), .A2(n1257), .ZN(n1256) );
NAND2_X1 U970 ( .A1(KEYINPUT54), .A2(G110), .ZN(n1255) );
AND2_X1 U971 ( .A1(n1258), .A2(G221), .ZN(n1253) );
XOR2_X1 U972 ( .A(n1259), .B(n1260), .Z(n1251) );
NOR2_X1 U973 ( .A1(KEYINPUT14), .A2(G119), .ZN(n1260) );
XOR2_X1 U974 ( .A(n1261), .B(G137), .Z(n1259) );
XNOR2_X1 U975 ( .A(n1262), .B(G472), .ZN(n1064) );
NAND2_X1 U976 ( .A1(n1263), .A2(n1138), .ZN(n1262) );
XOR2_X1 U977 ( .A(n1123), .B(n1264), .Z(n1263) );
NOR2_X1 U978 ( .A1(KEYINPUT30), .A2(n1265), .ZN(n1264) );
XOR2_X1 U979 ( .A(n1122), .B(n1266), .Z(n1265) );
NOR2_X1 U980 ( .A1(G101), .A2(KEYINPUT43), .ZN(n1266) );
NAND2_X1 U981 ( .A1(n1267), .A2(G210), .ZN(n1122) );
XOR2_X1 U982 ( .A(n1268), .B(n1269), .Z(n1123) );
XOR2_X1 U983 ( .A(n1225), .B(n1246), .Z(n1269) );
XOR2_X1 U984 ( .A(n1209), .B(G119), .Z(n1246) );
INV_X1 U985 ( .A(G116), .ZN(n1209) );
XOR2_X1 U986 ( .A(n1270), .B(G128), .Z(n1225) );
NAND2_X1 U987 ( .A1(n1271), .A2(KEYINPUT11), .ZN(n1270) );
XOR2_X1 U988 ( .A(n1272), .B(G143), .Z(n1271) );
NAND2_X1 U989 ( .A1(KEYINPUT17), .A2(n1178), .ZN(n1272) );
XOR2_X1 U990 ( .A(n1137), .B(n1273), .Z(n1268) );
XOR2_X1 U991 ( .A(KEYINPUT37), .B(G113), .Z(n1273) );
INV_X1 U992 ( .A(n1172), .ZN(n1038) );
NAND2_X1 U993 ( .A1(n1040), .A2(n1170), .ZN(n1172) );
NOR2_X1 U994 ( .A1(n1041), .A2(n1042), .ZN(n1170) );
AND2_X1 U995 ( .A1(G221), .A2(n1250), .ZN(n1042) );
NAND2_X1 U996 ( .A1(n1218), .A2(n1138), .ZN(n1250) );
XNOR2_X1 U997 ( .A(G234), .B(KEYINPUT25), .ZN(n1218) );
XNOR2_X1 U998 ( .A(n1063), .B(n1274), .ZN(n1041) );
XOR2_X1 U999 ( .A(KEYINPUT8), .B(G469), .Z(n1274) );
NAND2_X1 U1000 ( .A1(n1275), .A2(n1138), .ZN(n1063) );
XOR2_X1 U1001 ( .A(n1137), .B(n1276), .Z(n1275) );
XOR2_X1 U1002 ( .A(n1277), .B(n1278), .Z(n1276) );
NOR2_X1 U1003 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
XOR2_X1 U1004 ( .A(n1281), .B(KEYINPUT5), .Z(n1280) );
NAND4_X1 U1005 ( .A1(n1282), .A2(n1131), .A3(n1283), .A4(n1284), .ZN(n1281) );
NOR2_X1 U1006 ( .A1(n1285), .A2(n1131), .ZN(n1279) );
NAND2_X1 U1007 ( .A1(n1286), .A2(G227), .ZN(n1131) );
XOR2_X1 U1008 ( .A(n1068), .B(KEYINPUT16), .Z(n1286) );
AND3_X1 U1009 ( .A1(n1282), .A2(n1284), .A3(n1283), .ZN(n1285) );
NAND2_X1 U1010 ( .A1(G140), .A2(n1287), .ZN(n1283) );
NAND2_X1 U1011 ( .A1(KEYINPUT40), .A2(n1288), .ZN(n1287) );
NAND4_X1 U1012 ( .A1(KEYINPUT60), .A2(KEYINPUT40), .A3(n1288), .A4(n1132), .ZN(n1284) );
INV_X1 U1013 ( .A(G140), .ZN(n1132) );
OR2_X1 U1014 ( .A1(n1288), .A2(KEYINPUT60), .ZN(n1282) );
INV_X1 U1015 ( .A(G110), .ZN(n1288) );
NAND2_X1 U1016 ( .A1(n1289), .A2(KEYINPUT27), .ZN(n1277) );
XNOR2_X1 U1017 ( .A(n1290), .B(n1141), .ZN(n1289) );
NAND2_X1 U1018 ( .A1(n1291), .A2(n1292), .ZN(n1141) );
NAND2_X1 U1019 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
NAND2_X1 U1020 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
NAND2_X1 U1021 ( .A1(G101), .A2(n1297), .ZN(n1295) );
XNOR2_X1 U1022 ( .A(G104), .B(n1298), .ZN(n1293) );
NAND2_X1 U1023 ( .A1(n1192), .A2(n1299), .ZN(n1291) );
NAND2_X1 U1024 ( .A1(n1300), .A2(n1297), .ZN(n1299) );
INV_X1 U1025 ( .A(KEYINPUT23), .ZN(n1297) );
NAND2_X1 U1026 ( .A1(n1301), .A2(n1296), .ZN(n1300) );
INV_X1 U1027 ( .A(KEYINPUT39), .ZN(n1296) );
XOR2_X1 U1028 ( .A(n1298), .B(G104), .Z(n1301) );
NAND2_X1 U1029 ( .A1(KEYINPUT61), .A2(n1230), .ZN(n1298) );
INV_X1 U1030 ( .A(G101), .ZN(n1192) );
NAND2_X1 U1031 ( .A1(KEYINPUT1), .A2(n1079), .ZN(n1290) );
XNOR2_X1 U1032 ( .A(n1302), .B(n1303), .ZN(n1079) );
XOR2_X1 U1033 ( .A(G146), .B(G128), .Z(n1303) );
NAND2_X1 U1034 ( .A1(KEYINPUT35), .A2(n1180), .ZN(n1302) );
INV_X1 U1035 ( .A(G143), .ZN(n1180) );
XOR2_X1 U1036 ( .A(n1080), .B(n1082), .Z(n1137) );
XOR2_X1 U1037 ( .A(G131), .B(G134), .Z(n1082) );
INV_X1 U1038 ( .A(G137), .ZN(n1080) );
INV_X1 U1039 ( .A(n1023), .ZN(n1040) );
NAND2_X1 U1040 ( .A1(n1204), .A2(n1212), .ZN(n1023) );
NOR2_X1 U1041 ( .A1(n1050), .A2(n1304), .ZN(n1212) );
AND2_X1 U1042 ( .A1(G475), .A2(n1059), .ZN(n1304) );
NOR2_X1 U1043 ( .A1(n1059), .A2(G475), .ZN(n1050) );
NAND2_X1 U1044 ( .A1(n1112), .A2(n1138), .ZN(n1059) );
XNOR2_X1 U1045 ( .A(n1305), .B(n1306), .ZN(n1112) );
XNOR2_X1 U1046 ( .A(n1307), .B(n1308), .ZN(n1306) );
NOR2_X1 U1047 ( .A1(G104), .A2(KEYINPUT59), .ZN(n1308) );
NAND2_X1 U1048 ( .A1(n1309), .A2(KEYINPUT24), .ZN(n1307) );
XOR2_X1 U1049 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1050 ( .A(G143), .B(G131), .Z(n1311) );
XOR2_X1 U1051 ( .A(n1257), .B(n1312), .Z(n1310) );
AND2_X1 U1052 ( .A1(G214), .A2(n1267), .ZN(n1312) );
NOR2_X1 U1053 ( .A1(G953), .A2(G237), .ZN(n1267) );
XOR2_X1 U1054 ( .A(n1178), .B(n1081), .Z(n1257) );
XOR2_X1 U1055 ( .A(G125), .B(G140), .Z(n1081) );
INV_X1 U1056 ( .A(G146), .ZN(n1178) );
XOR2_X1 U1057 ( .A(n1242), .B(n1313), .Z(n1305) );
XOR2_X1 U1058 ( .A(KEYINPUT52), .B(G122), .Z(n1313) );
INV_X1 U1059 ( .A(G113), .ZN(n1242) );
XOR2_X1 U1060 ( .A(n1314), .B(G478), .Z(n1204) );
NAND2_X1 U1061 ( .A1(n1109), .A2(n1138), .ZN(n1314) );
INV_X1 U1062 ( .A(G902), .ZN(n1138) );
XNOR2_X1 U1063 ( .A(n1315), .B(n1316), .ZN(n1109) );
XOR2_X1 U1064 ( .A(n1317), .B(n1318), .Z(n1316) );
XOR2_X1 U1065 ( .A(G134), .B(G116), .Z(n1318) );
XOR2_X1 U1066 ( .A(KEYINPUT44), .B(G143), .Z(n1317) );
XOR2_X1 U1067 ( .A(n1319), .B(n1320), .Z(n1315) );
XOR2_X1 U1068 ( .A(n1321), .B(n1322), .Z(n1320) );
NAND2_X1 U1069 ( .A1(KEYINPUT62), .A2(n1261), .ZN(n1322) );
INV_X1 U1070 ( .A(G128), .ZN(n1261) );
NAND2_X1 U1071 ( .A1(G217), .A2(n1258), .ZN(n1321) );
AND2_X1 U1072 ( .A1(G234), .A2(n1068), .ZN(n1258) );
INV_X1 U1073 ( .A(G953), .ZN(n1068) );
XOR2_X1 U1074 ( .A(n1230), .B(n1323), .Z(n1319) );
NOR2_X1 U1075 ( .A1(G122), .A2(KEYINPUT41), .ZN(n1323) );
INV_X1 U1076 ( .A(G107), .ZN(n1230) );
endmodule


