//Key = 0000010110111001010011011110011000110001000011001010001100110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
n1513, n1514;

XOR2_X1 U815 ( .A(n1143), .B(n1144), .Z(G9) );
NAND2_X1 U816 ( .A1(KEYINPUT35), .A2(n1145), .ZN(n1143) );
NOR2_X1 U817 ( .A1(n1146), .A2(n1147), .ZN(G75) );
NOR4_X1 U818 ( .A1(G953), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1147) );
NOR2_X1 U819 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
NOR2_X1 U820 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U821 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U822 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
NOR2_X1 U823 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U824 ( .A1(n1161), .A2(n1162), .ZN(n1159) );
NOR2_X1 U825 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U826 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
AND3_X1 U827 ( .A1(KEYINPUT33), .A2(n1167), .A3(n1168), .ZN(n1161) );
NOR3_X1 U828 ( .A1(n1169), .A2(n1170), .A3(n1167), .ZN(n1157) );
NOR2_X1 U829 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U830 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NOR2_X1 U831 ( .A1(n1175), .A2(n1176), .ZN(n1173) );
NOR2_X1 U832 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
XOR2_X1 U833 ( .A(n1179), .B(KEYINPUT60), .Z(n1177) );
NOR3_X1 U834 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1171) );
NOR3_X1 U835 ( .A1(n1160), .A2(n1181), .A3(n1167), .ZN(n1153) );
INV_X1 U836 ( .A(n1183), .ZN(n1167) );
AND3_X1 U837 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1181) );
NAND2_X1 U838 ( .A1(n1187), .A2(n1188), .ZN(n1185) );
NAND2_X1 U839 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U840 ( .A1(n1191), .A2(n1192), .ZN(n1184) );
NAND2_X1 U841 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NAND3_X1 U842 ( .A1(n1195), .A2(n1180), .A3(n1196), .ZN(n1194) );
INV_X1 U843 ( .A(KEYINPUT47), .ZN(n1180) );
NAND2_X1 U844 ( .A1(n1168), .A2(n1197), .ZN(n1193) );
INV_X1 U845 ( .A(KEYINPUT33), .ZN(n1197) );
INV_X1 U846 ( .A(n1186), .ZN(n1160) );
INV_X1 U847 ( .A(n1198), .ZN(n1151) );
NOR3_X1 U848 ( .A1(n1148), .A2(G953), .A3(G952), .ZN(n1146) );
AND4_X1 U849 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1148) );
NOR3_X1 U850 ( .A1(n1203), .A2(n1195), .A3(n1204), .ZN(n1202) );
NAND3_X1 U851 ( .A1(n1179), .A2(n1205), .A3(n1206), .ZN(n1203) );
NOR3_X1 U852 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1201) );
XOR2_X1 U853 ( .A(n1196), .B(KEYINPUT29), .Z(n1209) );
NOR2_X1 U854 ( .A1(n1210), .A2(n1211), .ZN(n1208) );
AND2_X1 U855 ( .A1(n1212), .A2(n1213), .ZN(n1210) );
XOR2_X1 U856 ( .A(n1214), .B(n1215), .Z(n1199) );
NAND2_X1 U857 ( .A1(KEYINPUT17), .A2(n1216), .ZN(n1214) );
INV_X1 U858 ( .A(n1217), .ZN(n1216) );
XOR2_X1 U859 ( .A(n1218), .B(n1219), .Z(G72) );
XOR2_X1 U860 ( .A(n1220), .B(n1221), .Z(n1219) );
NOR3_X1 U861 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1221) );
NOR2_X1 U862 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XNOR2_X1 U863 ( .A(KEYINPUT16), .B(n1227), .ZN(n1226) );
INV_X1 U864 ( .A(n1228), .ZN(n1225) );
NOR2_X1 U865 ( .A1(n1228), .A2(n1227), .ZN(n1223) );
NAND2_X1 U866 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
XOR2_X1 U867 ( .A(KEYINPUT10), .B(n1231), .Z(n1229) );
NAND2_X1 U868 ( .A1(n1232), .A2(n1233), .ZN(n1228) );
NAND2_X1 U869 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U870 ( .A(KEYINPUT54), .B(n1236), .Z(n1232) );
NOR2_X1 U871 ( .A1(n1234), .A2(n1235), .ZN(n1236) );
INV_X1 U872 ( .A(n1237), .ZN(n1235) );
AND3_X1 U873 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1234) );
OR2_X1 U874 ( .A1(n1241), .A2(G131), .ZN(n1240) );
NAND2_X1 U875 ( .A1(n1242), .A2(n1243), .ZN(n1239) );
INV_X1 U876 ( .A(KEYINPUT59), .ZN(n1243) );
NAND2_X1 U877 ( .A1(n1244), .A2(n1241), .ZN(n1242) );
XNOR2_X1 U878 ( .A(KEYINPUT61), .B(G131), .ZN(n1244) );
NAND2_X1 U879 ( .A1(KEYINPUT59), .A2(n1245), .ZN(n1238) );
NAND2_X1 U880 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
OR2_X1 U881 ( .A1(G131), .A2(KEYINPUT61), .ZN(n1247) );
NAND3_X1 U882 ( .A1(G131), .A2(n1241), .A3(KEYINPUT61), .ZN(n1246) );
XOR2_X1 U883 ( .A(G134), .B(G137), .Z(n1241) );
NAND3_X1 U884 ( .A1(G953), .A2(n1248), .A3(KEYINPUT48), .ZN(n1220) );
NAND2_X1 U885 ( .A1(G900), .A2(G227), .ZN(n1248) );
NAND2_X1 U886 ( .A1(n1249), .A2(n1250), .ZN(n1218) );
NAND2_X1 U887 ( .A1(n1251), .A2(n1252), .ZN(G69) );
NAND2_X1 U888 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
OR2_X1 U889 ( .A1(n1249), .A2(G224), .ZN(n1254) );
NAND3_X1 U890 ( .A1(G953), .A2(n1255), .A3(n1256), .ZN(n1251) );
INV_X1 U891 ( .A(n1253), .ZN(n1256) );
NOR2_X1 U892 ( .A1(KEYINPUT4), .A2(n1257), .ZN(n1253) );
XOR2_X1 U893 ( .A(n1258), .B(n1259), .Z(n1257) );
NOR3_X1 U894 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1259) );
INV_X1 U895 ( .A(n1263), .ZN(n1261) );
XOR2_X1 U896 ( .A(n1264), .B(KEYINPUT20), .Z(n1260) );
NAND2_X1 U897 ( .A1(n1249), .A2(n1265), .ZN(n1258) );
NAND2_X1 U898 ( .A1(G898), .A2(G224), .ZN(n1255) );
NOR2_X1 U899 ( .A1(n1266), .A2(n1267), .ZN(G66) );
NOR3_X1 U900 ( .A1(n1268), .A2(n1215), .A3(n1269), .ZN(n1267) );
NOR2_X1 U901 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XOR2_X1 U902 ( .A(KEYINPUT49), .B(n1272), .Z(n1268) );
AND3_X1 U903 ( .A1(n1270), .A2(n1271), .A3(G902), .ZN(n1272) );
AND3_X1 U904 ( .A1(n1150), .A2(n1273), .A3(G217), .ZN(n1270) );
NOR2_X1 U905 ( .A1(n1266), .A2(n1274), .ZN(G63) );
XOR2_X1 U906 ( .A(n1275), .B(n1213), .Z(n1274) );
NAND2_X1 U907 ( .A1(n1276), .A2(G478), .ZN(n1275) );
NOR2_X1 U908 ( .A1(n1266), .A2(n1277), .ZN(G60) );
XOR2_X1 U909 ( .A(n1278), .B(n1279), .Z(n1277) );
NOR2_X1 U910 ( .A1(KEYINPUT28), .A2(n1280), .ZN(n1279) );
XOR2_X1 U911 ( .A(n1281), .B(n1282), .Z(n1280) );
NAND2_X1 U912 ( .A1(n1276), .A2(G475), .ZN(n1278) );
XNOR2_X1 U913 ( .A(G104), .B(n1283), .ZN(G6) );
NOR2_X1 U914 ( .A1(n1266), .A2(n1284), .ZN(G57) );
XOR2_X1 U915 ( .A(n1285), .B(n1286), .Z(n1284) );
NAND2_X1 U916 ( .A1(KEYINPUT58), .A2(n1287), .ZN(n1285) );
XNOR2_X1 U917 ( .A(n1288), .B(n1289), .ZN(n1287) );
XOR2_X1 U918 ( .A(n1290), .B(n1291), .Z(n1289) );
NOR2_X1 U919 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XOR2_X1 U920 ( .A(KEYINPUT3), .B(n1294), .Z(n1293) );
NOR2_X1 U921 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
NOR2_X1 U922 ( .A1(n1297), .A2(n1298), .ZN(n1292) );
NAND2_X1 U923 ( .A1(n1276), .A2(G472), .ZN(n1290) );
NOR2_X1 U924 ( .A1(n1266), .A2(n1299), .ZN(G54) );
XOR2_X1 U925 ( .A(n1300), .B(n1301), .Z(n1299) );
XOR2_X1 U926 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U927 ( .A(n1237), .B(n1304), .Z(n1303) );
XOR2_X1 U928 ( .A(n1305), .B(n1296), .Z(n1300) );
XOR2_X1 U929 ( .A(n1306), .B(n1307), .Z(n1305) );
NOR2_X1 U930 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
XOR2_X1 U931 ( .A(KEYINPUT19), .B(n1310), .Z(n1309) );
NAND3_X1 U932 ( .A1(n1276), .A2(G469), .A3(KEYINPUT15), .ZN(n1306) );
NOR2_X1 U933 ( .A1(n1266), .A2(n1311), .ZN(G51) );
NOR2_X1 U934 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
XOR2_X1 U935 ( .A(n1314), .B(KEYINPUT8), .Z(n1313) );
NAND2_X1 U936 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NOR2_X1 U937 ( .A1(n1315), .A2(n1316), .ZN(n1312) );
XOR2_X1 U938 ( .A(n1317), .B(n1318), .Z(n1316) );
NOR2_X1 U939 ( .A1(KEYINPUT0), .A2(n1319), .ZN(n1318) );
NOR3_X1 U940 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1319) );
AND3_X1 U941 ( .A1(KEYINPUT30), .A2(n1323), .A3(n1324), .ZN(n1322) );
NOR2_X1 U942 ( .A1(KEYINPUT30), .A2(n1324), .ZN(n1321) );
AND3_X1 U943 ( .A1(G210), .A2(n1325), .A3(n1276), .ZN(n1315) );
AND2_X1 U944 ( .A1(G902), .A2(n1150), .ZN(n1276) );
OR2_X1 U945 ( .A1(n1250), .A2(n1265), .ZN(n1150) );
NAND4_X1 U946 ( .A1(n1283), .A2(n1326), .A3(n1327), .A4(n1328), .ZN(n1265) );
NOR4_X1 U947 ( .A1(n1144), .A2(n1329), .A3(n1330), .A4(n1331), .ZN(n1328) );
AND3_X1 U948 ( .A1(n1183), .A2(n1332), .A3(n1333), .ZN(n1144) );
NAND2_X1 U949 ( .A1(n1176), .A2(n1334), .ZN(n1327) );
NAND2_X1 U950 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
NAND3_X1 U951 ( .A1(n1166), .A2(n1337), .A3(n1338), .ZN(n1336) );
XOR2_X1 U952 ( .A(n1339), .B(KEYINPUT40), .Z(n1335) );
NAND3_X1 U953 ( .A1(n1333), .A2(n1183), .A3(n1337), .ZN(n1283) );
NAND4_X1 U954 ( .A1(n1340), .A2(n1341), .A3(n1342), .A4(n1343), .ZN(n1250) );
NOR4_X1 U955 ( .A1(n1344), .A2(n1345), .A3(n1346), .A4(n1347), .ZN(n1343) );
NOR3_X1 U956 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1342) );
NOR4_X1 U957 ( .A1(n1351), .A2(n1352), .A3(n1353), .A4(n1354), .ZN(n1350) );
NAND3_X1 U958 ( .A1(n1168), .A2(n1176), .A3(n1332), .ZN(n1352) );
INV_X1 U959 ( .A(KEYINPUT6), .ZN(n1351) );
NOR2_X1 U960 ( .A1(KEYINPUT6), .A2(n1355), .ZN(n1349) );
NOR3_X1 U961 ( .A1(n1356), .A2(n1357), .A3(n1156), .ZN(n1348) );
XOR2_X1 U962 ( .A(KEYINPUT39), .B(n1358), .Z(n1356) );
NOR2_X1 U963 ( .A1(n1249), .A2(G952), .ZN(n1266) );
XOR2_X1 U964 ( .A(n1359), .B(n1340), .Z(G48) );
NAND3_X1 U965 ( .A1(n1360), .A2(n1337), .A3(n1358), .ZN(n1340) );
XNOR2_X1 U966 ( .A(n1361), .B(n1341), .ZN(G45) );
NAND4_X1 U967 ( .A1(n1360), .A2(n1166), .A3(n1362), .A4(n1363), .ZN(n1341) );
NAND2_X1 U968 ( .A1(KEYINPUT55), .A2(n1364), .ZN(n1361) );
XOR2_X1 U969 ( .A(G140), .B(n1347), .Z(G42) );
AND3_X1 U970 ( .A1(n1337), .A2(n1165), .A3(n1365), .ZN(n1347) );
XOR2_X1 U971 ( .A(G137), .B(n1366), .Z(G39) );
AND2_X1 U972 ( .A1(n1365), .A2(n1367), .ZN(n1366) );
XOR2_X1 U973 ( .A(G134), .B(n1346), .Z(G36) );
AND3_X1 U974 ( .A1(n1365), .A2(n1332), .A3(n1166), .ZN(n1346) );
XOR2_X1 U975 ( .A(G131), .B(n1345), .Z(G33) );
AND3_X1 U976 ( .A1(n1365), .A2(n1337), .A3(n1166), .ZN(n1345) );
INV_X1 U977 ( .A(n1357), .ZN(n1365) );
NAND3_X1 U978 ( .A1(n1168), .A2(n1354), .A3(n1186), .ZN(n1357) );
NOR2_X1 U979 ( .A1(n1368), .A2(n1178), .ZN(n1186) );
XNOR2_X1 U980 ( .A(n1179), .B(KEYINPUT14), .ZN(n1368) );
XOR2_X1 U981 ( .A(n1369), .B(n1355), .Z(G30) );
NAND3_X1 U982 ( .A1(n1360), .A2(n1332), .A3(n1358), .ZN(n1355) );
INV_X1 U983 ( .A(n1353), .ZN(n1358) );
AND3_X1 U984 ( .A1(n1176), .A2(n1354), .A3(n1168), .ZN(n1360) );
XOR2_X1 U985 ( .A(n1370), .B(n1326), .Z(G3) );
NAND3_X1 U986 ( .A1(n1166), .A2(n1333), .A3(n1191), .ZN(n1326) );
NAND2_X1 U987 ( .A1(n1371), .A2(n1372), .ZN(G27) );
NAND2_X1 U988 ( .A1(n1344), .A2(n1373), .ZN(n1372) );
XOR2_X1 U989 ( .A(KEYINPUT12), .B(n1374), .Z(n1371) );
NOR2_X1 U990 ( .A1(n1344), .A2(n1373), .ZN(n1374) );
AND4_X1 U991 ( .A1(n1176), .A2(n1354), .A3(n1165), .A4(n1375), .ZN(n1344) );
NOR2_X1 U992 ( .A1(n1164), .A2(n1190), .ZN(n1375) );
INV_X1 U993 ( .A(n1187), .ZN(n1164) );
NAND2_X1 U994 ( .A1(n1376), .A2(n1377), .ZN(n1354) );
NAND3_X1 U995 ( .A1(G902), .A2(n1198), .A3(n1222), .ZN(n1377) );
NOR2_X1 U996 ( .A1(n1249), .A2(G900), .ZN(n1222) );
XOR2_X1 U997 ( .A(G122), .B(n1331), .Z(G24) );
AND4_X1 U998 ( .A1(n1338), .A2(n1183), .A3(n1378), .A4(n1176), .ZN(n1331) );
NOR2_X1 U999 ( .A1(n1379), .A2(n1200), .ZN(n1378) );
NOR2_X1 U1000 ( .A1(n1380), .A2(n1207), .ZN(n1183) );
XOR2_X1 U1001 ( .A(G119), .B(n1381), .Z(G21) );
NOR2_X1 U1002 ( .A1(n1382), .A2(n1339), .ZN(n1381) );
NAND2_X1 U1003 ( .A1(n1367), .A2(n1338), .ZN(n1339) );
NOR2_X1 U1004 ( .A1(n1156), .A2(n1353), .ZN(n1367) );
NAND2_X1 U1005 ( .A1(n1207), .A2(n1380), .ZN(n1353) );
NAND2_X1 U1006 ( .A1(n1383), .A2(n1384), .ZN(G18) );
NAND2_X1 U1007 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
XOR2_X1 U1008 ( .A(KEYINPUT36), .B(n1330), .Z(n1385) );
INV_X1 U1009 ( .A(n1387), .ZN(n1330) );
NAND2_X1 U1010 ( .A1(G116), .A2(n1388), .ZN(n1383) );
XOR2_X1 U1011 ( .A(n1387), .B(KEYINPUT9), .Z(n1388) );
NAND4_X1 U1012 ( .A1(n1338), .A2(n1166), .A3(n1332), .A4(n1176), .ZN(n1387) );
INV_X1 U1013 ( .A(n1189), .ZN(n1332) );
NAND2_X1 U1014 ( .A1(n1389), .A2(n1363), .ZN(n1189) );
XNOR2_X1 U1015 ( .A(G113), .B(n1390), .ZN(G15) );
NAND4_X1 U1016 ( .A1(n1338), .A2(n1166), .A3(n1337), .A4(n1391), .ZN(n1390) );
XOR2_X1 U1017 ( .A(KEYINPUT41), .B(n1176), .Z(n1391) );
INV_X1 U1018 ( .A(n1190), .ZN(n1337) );
NAND2_X1 U1019 ( .A1(n1379), .A2(n1362), .ZN(n1190) );
INV_X1 U1020 ( .A(n1200), .ZN(n1362) );
AND2_X1 U1021 ( .A1(n1392), .A2(n1207), .ZN(n1166) );
AND2_X1 U1022 ( .A1(n1187), .A2(n1393), .ZN(n1338) );
NOR2_X1 U1023 ( .A1(n1169), .A2(n1174), .ZN(n1187) );
INV_X1 U1024 ( .A(n1196), .ZN(n1169) );
XOR2_X1 U1025 ( .A(G110), .B(n1329), .Z(G12) );
AND3_X1 U1026 ( .A1(n1165), .A2(n1333), .A3(n1191), .ZN(n1329) );
INV_X1 U1027 ( .A(n1156), .ZN(n1191) );
NAND2_X1 U1028 ( .A1(n1379), .A2(n1389), .ZN(n1156) );
XOR2_X1 U1029 ( .A(n1200), .B(KEYINPUT32), .Z(n1389) );
XOR2_X1 U1030 ( .A(n1394), .B(G475), .Z(n1200) );
NAND2_X1 U1031 ( .A1(n1395), .A2(n1212), .ZN(n1394) );
XNOR2_X1 U1032 ( .A(n1282), .B(n1281), .ZN(n1395) );
XOR2_X1 U1033 ( .A(n1396), .B(n1397), .Z(n1281) );
XOR2_X1 U1034 ( .A(n1398), .B(n1399), .Z(n1397) );
NAND3_X1 U1035 ( .A1(n1400), .A2(n1401), .A3(n1402), .ZN(n1399) );
NAND2_X1 U1036 ( .A1(n1403), .A2(G146), .ZN(n1402) );
NAND2_X1 U1037 ( .A1(n1404), .A2(n1405), .ZN(n1401) );
INV_X1 U1038 ( .A(KEYINPUT51), .ZN(n1405) );
NAND2_X1 U1039 ( .A1(n1406), .A2(KEYINPUT51), .ZN(n1400) );
XOR2_X1 U1040 ( .A(G146), .B(n1231), .Z(n1406) );
NAND3_X1 U1041 ( .A1(G214), .A2(n1407), .A3(n1408), .ZN(n1398) );
XOR2_X1 U1042 ( .A(n1249), .B(KEYINPUT37), .Z(n1408) );
XNOR2_X1 U1043 ( .A(n1409), .B(n1410), .ZN(n1282) );
XOR2_X1 U1044 ( .A(KEYINPUT44), .B(G143), .Z(n1410) );
XNOR2_X1 U1045 ( .A(G122), .B(G131), .ZN(n1409) );
INV_X1 U1046 ( .A(n1363), .ZN(n1379) );
NAND2_X1 U1047 ( .A1(n1411), .A2(n1205), .ZN(n1363) );
NAND3_X1 U1048 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1205) );
INV_X1 U1049 ( .A(G478), .ZN(n1211) );
NAND2_X1 U1050 ( .A1(n1412), .A2(n1413), .ZN(n1411) );
NAND2_X1 U1051 ( .A1(n1213), .A2(n1212), .ZN(n1413) );
XNOR2_X1 U1052 ( .A(n1414), .B(n1415), .ZN(n1213) );
XOR2_X1 U1053 ( .A(n1416), .B(n1417), .Z(n1415) );
XOR2_X1 U1054 ( .A(n1386), .B(G134), .Z(n1417) );
NAND3_X1 U1055 ( .A1(n1418), .A2(n1419), .A3(n1420), .ZN(n1416) );
OR3_X1 U1056 ( .A1(G128), .A2(G143), .A3(KEYINPUT18), .ZN(n1419) );
NAND2_X1 U1057 ( .A1(KEYINPUT18), .A2(G128), .ZN(n1418) );
XOR2_X1 U1058 ( .A(n1421), .B(n1422), .Z(n1414) );
NAND3_X1 U1059 ( .A1(G234), .A2(n1249), .A3(G217), .ZN(n1421) );
XOR2_X1 U1060 ( .A(KEYINPUT31), .B(G478), .Z(n1412) );
AND3_X1 U1061 ( .A1(n1176), .A2(n1393), .A3(n1168), .ZN(n1333) );
NOR2_X1 U1062 ( .A1(n1196), .A2(n1174), .ZN(n1168) );
XNOR2_X1 U1063 ( .A(n1195), .B(KEYINPUT45), .ZN(n1174) );
INV_X1 U1064 ( .A(n1182), .ZN(n1195) );
NAND2_X1 U1065 ( .A1(G221), .A2(n1273), .ZN(n1182) );
XNOR2_X1 U1066 ( .A(G469), .B(n1423), .ZN(n1196) );
NOR2_X1 U1067 ( .A1(G902), .A2(n1424), .ZN(n1423) );
NOR2_X1 U1068 ( .A1(n1425), .A2(n1426), .ZN(n1424) );
XOR2_X1 U1069 ( .A(n1427), .B(KEYINPUT7), .Z(n1426) );
NAND2_X1 U1070 ( .A1(n1428), .A2(n1429), .ZN(n1427) );
OR2_X1 U1071 ( .A1(n1430), .A2(n1431), .ZN(n1429) );
NOR3_X1 U1072 ( .A1(n1430), .A2(n1431), .A3(n1428), .ZN(n1425) );
XOR2_X1 U1073 ( .A(n1432), .B(n1296), .Z(n1428) );
INV_X1 U1074 ( .A(n1297), .ZN(n1296) );
NAND3_X1 U1075 ( .A1(n1433), .A2(n1434), .A3(n1435), .ZN(n1432) );
NAND2_X1 U1076 ( .A1(n1302), .A2(n1436), .ZN(n1435) );
INV_X1 U1077 ( .A(KEYINPUT50), .ZN(n1436) );
NAND3_X1 U1078 ( .A1(KEYINPUT50), .A2(n1437), .A3(n1237), .ZN(n1434) );
OR2_X1 U1079 ( .A1(n1237), .A2(n1437), .ZN(n1433) );
NOR2_X1 U1080 ( .A1(KEYINPUT22), .A2(n1302), .ZN(n1437) );
NAND2_X1 U1081 ( .A1(n1438), .A2(n1439), .ZN(n1302) );
NAND2_X1 U1082 ( .A1(n1440), .A2(n1370), .ZN(n1439) );
XOR2_X1 U1083 ( .A(KEYINPUT11), .B(n1441), .Z(n1438) );
NOR2_X1 U1084 ( .A1(n1370), .A2(n1440), .ZN(n1441) );
XNOR2_X1 U1085 ( .A(G104), .B(n1442), .ZN(n1440) );
NOR2_X1 U1086 ( .A1(n1443), .A2(n1444), .ZN(n1442) );
NOR2_X1 U1087 ( .A1(KEYINPUT38), .A2(G107), .ZN(n1444) );
NOR2_X1 U1088 ( .A1(KEYINPUT63), .A2(n1145), .ZN(n1443) );
INV_X1 U1089 ( .A(G107), .ZN(n1145) );
INV_X1 U1090 ( .A(G101), .ZN(n1370) );
NAND4_X1 U1091 ( .A1(n1445), .A2(n1446), .A3(n1447), .A4(n1448), .ZN(n1237) );
NAND3_X1 U1092 ( .A1(G146), .A2(n1449), .A3(KEYINPUT34), .ZN(n1448) );
NAND2_X1 U1093 ( .A1(n1450), .A2(n1451), .ZN(n1447) );
INV_X1 U1094 ( .A(KEYINPUT34), .ZN(n1451) );
NAND2_X1 U1095 ( .A1(n1420), .A2(n1452), .ZN(n1450) );
NAND2_X1 U1096 ( .A1(G128), .A2(n1359), .ZN(n1452) );
NAND3_X1 U1097 ( .A1(n1369), .A2(n1364), .A3(n1453), .ZN(n1446) );
XOR2_X1 U1098 ( .A(KEYINPUT34), .B(G146), .Z(n1453) );
INV_X1 U1099 ( .A(G143), .ZN(n1364) );
INV_X1 U1100 ( .A(G128), .ZN(n1369) );
OR2_X1 U1101 ( .A1(n1420), .A2(G146), .ZN(n1445) );
NAND2_X1 U1102 ( .A1(G143), .A2(G128), .ZN(n1420) );
NOR2_X1 U1103 ( .A1(n1454), .A2(n1304), .ZN(n1431) );
XNOR2_X1 U1104 ( .A(n1455), .B(KEYINPUT53), .ZN(n1430) );
NAND2_X1 U1105 ( .A1(n1304), .A2(n1454), .ZN(n1455) );
NOR2_X1 U1106 ( .A1(n1308), .A2(n1310), .ZN(n1454) );
NOR2_X1 U1107 ( .A1(n1456), .A2(n1457), .ZN(n1310) );
INV_X1 U1108 ( .A(G110), .ZN(n1457) );
NOR2_X1 U1109 ( .A1(n1458), .A2(G110), .ZN(n1308) );
AND2_X1 U1110 ( .A1(G227), .A2(n1249), .ZN(n1304) );
NAND2_X1 U1111 ( .A1(n1376), .A2(n1459), .ZN(n1393) );
NAND3_X1 U1112 ( .A1(G902), .A2(n1198), .A3(n1262), .ZN(n1459) );
NOR2_X1 U1113 ( .A1(n1249), .A2(G898), .ZN(n1262) );
NAND3_X1 U1114 ( .A1(n1198), .A2(n1249), .A3(n1460), .ZN(n1376) );
XOR2_X1 U1115 ( .A(KEYINPUT46), .B(G952), .Z(n1460) );
NAND2_X1 U1116 ( .A1(G237), .A2(G234), .ZN(n1198) );
INV_X1 U1117 ( .A(n1382), .ZN(n1176) );
NAND2_X1 U1118 ( .A1(n1178), .A2(n1179), .ZN(n1382) );
NAND2_X1 U1119 ( .A1(G214), .A2(n1325), .ZN(n1179) );
NAND2_X1 U1120 ( .A1(n1461), .A2(n1206), .ZN(n1178) );
NAND3_X1 U1121 ( .A1(n1462), .A2(n1325), .A3(G210), .ZN(n1206) );
XNOR2_X1 U1122 ( .A(n1204), .B(KEYINPUT27), .ZN(n1461) );
NOR2_X1 U1123 ( .A1(n1462), .A2(n1463), .ZN(n1204) );
AND2_X1 U1124 ( .A1(G210), .A2(n1325), .ZN(n1463) );
NAND2_X1 U1125 ( .A1(n1464), .A2(n1407), .ZN(n1325) );
NAND3_X1 U1126 ( .A1(n1465), .A2(n1212), .A3(n1466), .ZN(n1462) );
XOR2_X1 U1127 ( .A(n1467), .B(KEYINPUT43), .Z(n1466) );
NAND2_X1 U1128 ( .A1(n1468), .A2(n1317), .ZN(n1467) );
OR2_X1 U1129 ( .A1(n1317), .A2(n1468), .ZN(n1465) );
NOR2_X1 U1130 ( .A1(n1320), .A2(n1469), .ZN(n1468) );
AND2_X1 U1131 ( .A1(n1324), .A2(n1323), .ZN(n1469) );
NOR2_X1 U1132 ( .A1(n1323), .A2(n1324), .ZN(n1320) );
XOR2_X1 U1133 ( .A(n1373), .B(n1295), .Z(n1324) );
INV_X1 U1134 ( .A(G125), .ZN(n1373) );
NAND2_X1 U1135 ( .A1(G224), .A2(n1249), .ZN(n1323) );
NAND2_X1 U1136 ( .A1(n1470), .A2(n1471), .ZN(n1317) );
NAND2_X1 U1137 ( .A1(KEYINPUT13), .A2(n1472), .ZN(n1471) );
XOR2_X1 U1138 ( .A(n1473), .B(n1474), .Z(n1472) );
XOR2_X1 U1139 ( .A(G110), .B(n1422), .Z(n1474) );
XOR2_X1 U1140 ( .A(G107), .B(G122), .Z(n1422) );
NAND3_X1 U1141 ( .A1(n1264), .A2(n1263), .A3(n1475), .ZN(n1470) );
INV_X1 U1142 ( .A(KEYINPUT13), .ZN(n1475) );
NAND2_X1 U1143 ( .A1(n1476), .A2(n1477), .ZN(n1263) );
OR2_X1 U1144 ( .A1(n1477), .A2(n1476), .ZN(n1264) );
XNOR2_X1 U1145 ( .A(n1473), .B(G107), .ZN(n1476) );
XOR2_X1 U1146 ( .A(n1478), .B(n1479), .Z(n1473) );
XOR2_X1 U1147 ( .A(G116), .B(G101), .Z(n1479) );
XOR2_X1 U1148 ( .A(n1480), .B(n1396), .Z(n1478) );
XOR2_X1 U1149 ( .A(G113), .B(G104), .Z(n1396) );
NAND2_X1 U1150 ( .A1(KEYINPUT26), .A2(n1481), .ZN(n1480) );
XOR2_X1 U1151 ( .A(G122), .B(G110), .Z(n1477) );
NOR2_X1 U1152 ( .A1(n1207), .A2(n1392), .ZN(n1165) );
INV_X1 U1153 ( .A(n1380), .ZN(n1392) );
NAND2_X1 U1154 ( .A1(n1482), .A2(n1483), .ZN(n1380) );
OR2_X1 U1155 ( .A1(n1217), .A2(n1215), .ZN(n1483) );
XOR2_X1 U1156 ( .A(n1484), .B(KEYINPUT52), .Z(n1482) );
NAND2_X1 U1157 ( .A1(n1215), .A2(n1217), .ZN(n1484) );
NAND2_X1 U1158 ( .A1(n1485), .A2(n1273), .ZN(n1217) );
NAND2_X1 U1159 ( .A1(G234), .A2(n1464), .ZN(n1273) );
XOR2_X1 U1160 ( .A(n1212), .B(KEYINPUT57), .Z(n1464) );
XOR2_X1 U1161 ( .A(KEYINPUT42), .B(G217), .Z(n1485) );
NOR2_X1 U1162 ( .A1(n1271), .A2(G902), .ZN(n1215) );
XNOR2_X1 U1163 ( .A(n1486), .B(n1487), .ZN(n1271) );
XOR2_X1 U1164 ( .A(n1488), .B(n1489), .Z(n1487) );
XOR2_X1 U1165 ( .A(G110), .B(n1490), .Z(n1489) );
NOR2_X1 U1166 ( .A1(n1491), .A2(n1404), .ZN(n1490) );
NAND2_X1 U1167 ( .A1(n1492), .A2(n1493), .ZN(n1404) );
OR3_X1 U1168 ( .A1(n1403), .A2(n1231), .A3(G146), .ZN(n1493) );
INV_X1 U1169 ( .A(n1230), .ZN(n1403) );
NAND2_X1 U1170 ( .A1(n1231), .A2(G146), .ZN(n1492) );
NOR2_X1 U1171 ( .A1(n1458), .A2(G125), .ZN(n1231) );
NOR2_X1 U1172 ( .A1(n1359), .A2(n1230), .ZN(n1491) );
NAND2_X1 U1173 ( .A1(G125), .A2(n1458), .ZN(n1230) );
INV_X1 U1174 ( .A(n1456), .ZN(n1458) );
XNOR2_X1 U1175 ( .A(G140), .B(KEYINPUT5), .ZN(n1456) );
NOR2_X1 U1176 ( .A1(n1494), .A2(n1495), .ZN(n1488) );
XOR2_X1 U1177 ( .A(n1496), .B(KEYINPUT25), .Z(n1495) );
NAND2_X1 U1178 ( .A1(n1497), .A2(G137), .ZN(n1496) );
NOR2_X1 U1179 ( .A1(G137), .A2(n1497), .ZN(n1494) );
AND3_X1 U1180 ( .A1(G234), .A2(n1249), .A3(G221), .ZN(n1497) );
XOR2_X1 U1181 ( .A(n1481), .B(n1498), .Z(n1486) );
XOR2_X1 U1182 ( .A(KEYINPUT23), .B(G128), .Z(n1498) );
INV_X1 U1183 ( .A(G119), .ZN(n1481) );
XNOR2_X1 U1184 ( .A(n1499), .B(G472), .ZN(n1207) );
NAND2_X1 U1185 ( .A1(n1500), .A2(n1212), .ZN(n1499) );
INV_X1 U1186 ( .A(G902), .ZN(n1212) );
XOR2_X1 U1187 ( .A(n1501), .B(n1502), .Z(n1500) );
XOR2_X1 U1188 ( .A(n1503), .B(n1298), .Z(n1502) );
INV_X1 U1189 ( .A(n1295), .ZN(n1298) );
XOR2_X1 U1190 ( .A(n1359), .B(n1449), .Z(n1295) );
XOR2_X1 U1191 ( .A(G143), .B(G128), .Z(n1449) );
INV_X1 U1192 ( .A(G146), .ZN(n1359) );
INV_X1 U1193 ( .A(n1286), .ZN(n1503) );
XOR2_X1 U1194 ( .A(n1504), .B(G101), .Z(n1286) );
NAND3_X1 U1195 ( .A1(n1407), .A2(n1249), .A3(G210), .ZN(n1504) );
INV_X1 U1196 ( .A(G953), .ZN(n1249) );
INV_X1 U1197 ( .A(G237), .ZN(n1407) );
XNOR2_X1 U1198 ( .A(n1505), .B(n1506), .ZN(n1501) );
NOR2_X1 U1199 ( .A1(KEYINPUT56), .A2(n1288), .ZN(n1506) );
XNOR2_X1 U1200 ( .A(n1507), .B(G113), .ZN(n1288) );
NAND2_X1 U1201 ( .A1(n1508), .A2(KEYINPUT21), .ZN(n1507) );
XOR2_X1 U1202 ( .A(n1386), .B(G119), .Z(n1508) );
INV_X1 U1203 ( .A(G116), .ZN(n1386) );
NAND2_X1 U1204 ( .A1(KEYINPUT24), .A2(n1297), .ZN(n1505) );
XNOR2_X1 U1205 ( .A(G131), .B(n1509), .ZN(n1297) );
NOR2_X1 U1206 ( .A1(n1510), .A2(n1511), .ZN(n1509) );
XOR2_X1 U1207 ( .A(KEYINPUT2), .B(n1512), .Z(n1511) );
NOR2_X1 U1208 ( .A1(G134), .A2(n1513), .ZN(n1512) );
XOR2_X1 U1209 ( .A(KEYINPUT1), .B(n1514), .Z(n1513) );
AND2_X1 U1210 ( .A1(n1514), .A2(G134), .ZN(n1510) );
XOR2_X1 U1211 ( .A(G137), .B(KEYINPUT62), .Z(n1514) );
endmodule


