//Key = 110000000000010000000000000000000000000000000000010000101000000001010000000000000000000100100100000000000000000000000000100000000000000000110110001100000001100000001000000000000000000000
module c7552 ( G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, 
        G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, 
        G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, 
        G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, 
        G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, 
        G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, 
        G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, 
        G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, 
        G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, 
        G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, 
        G239, G240, G1197, G1455, G1459, G1462, G1469, G1480, G1486, 
        G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, 
        G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, 
        G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, 
        G4427, G4432, G4437, G4526, G4528, KEYINPUT0, KEYINPUT1, KEYINPUT2, 
        KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, 
        KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, 
        KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, 
        KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, 
        KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, 
        KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, 
        KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, 
        KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, 
        KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, 
        KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, 
        KEYINPUT63, KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, 
        KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, 
        KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, 
        KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, 
        KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, 
        KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, 
        KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, 
        KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, 
        KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, 
        KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, 
        KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, 
        KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT128, 
        KEYINPUT129, KEYINPUT130, KEYINPUT131, KEYINPUT132, KEYINPUT133, 
        KEYINPUT134, KEYINPUT135, KEYINPUT136, KEYINPUT137, KEYINPUT138, 
        KEYINPUT139, KEYINPUT140, KEYINPUT141, KEYINPUT142, KEYINPUT143, 
        KEYINPUT144, KEYINPUT145, KEYINPUT146, KEYINPUT147, KEYINPUT148, 
        KEYINPUT149, KEYINPUT150, KEYINPUT151, KEYINPUT152, KEYINPUT153, 
        KEYINPUT154, KEYINPUT155, KEYINPUT156, KEYINPUT157, KEYINPUT158, 
        KEYINPUT159, KEYINPUT160, KEYINPUT161, KEYINPUT162, KEYINPUT163, 
        KEYINPUT164, KEYINPUT165, KEYINPUT166, KEYINPUT167, KEYINPUT168, 
        KEYINPUT169, KEYINPUT170, KEYINPUT171, KEYINPUT172, KEYINPUT173, 
        KEYINPUT174, KEYINPUT175, KEYINPUT176, KEYINPUT177, KEYINPUT178, 
        KEYINPUT179, KEYINPUT180, KEYINPUT181, KEYINPUT182, KEYINPUT183, 
        KEYINPUT184, KEYINPUT185, G2, G3, G450, G448, G444, G442, G440, G438, 
        G496, G494, G492, G490, G488, G486, G484, G482, G480, G560, G542, G558, 
        G556, G554, G552, G550, G548, G546, G544, G540, G538, G536, G534, G532, 
        G530, G528, G526, G524, G279, G436, G478, G522, G402, G404, G406, G408, 
        G410, G432, G446, G284, G286, G289, G292, G341, G281, G453, G278, G373, 
        G246, G258, G264, G270, G388, G391, G394, G397, G376, G379, G382, G385, 
        G412_enc, G414_enc, G416_enc, G249, G295, G324, G252, G276, G310, G313,         
        G316, G319, G327, G330, G333, G336, G418_enc, G273, G298, G301, G304,  G307, 
        G344, G422, G469, G419, G471, G359, G362, G365, G368, G347, G350,  G353, G356, G321, G338, G370, G399 );
  input G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47,
         G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65,
         G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83,
         G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110,
         G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133,
         G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
         G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165,
         G166, G167, G168, G169, G170, G171, G172, G173, G174, G175, G176,
         G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G187,
         G188, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198,
         G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209,
         G210, G211, G212, G213, G214, G215, G216, G217, G218, G219, G220,
         G221, G222, G223, G224, G225, G226, G227, G228, G229, G230, G231,
         G232, G233, G234, G235, G236, G237, G238, G239, G240, G1197,
         G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208,
         G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698,
         G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393,
         G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526,
         G4528, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
         KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
         KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15,
         KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
         KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
         KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
         KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
         KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
         KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45,
         KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
         KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
         KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
         KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
         KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
         KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
         KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
         KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85,
         KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90,
         KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
         KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
         KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
         KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
         KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
         KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
         KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
         KEYINPUT126, KEYINPUT127, KEYINPUT128, KEYINPUT129, KEYINPUT130,
         KEYINPUT131, KEYINPUT132, KEYINPUT133, KEYINPUT134, KEYINPUT135,
         KEYINPUT136, KEYINPUT137, KEYINPUT138, KEYINPUT139, KEYINPUT140,
         KEYINPUT141, KEYINPUT142, KEYINPUT143, KEYINPUT144, KEYINPUT145,
         KEYINPUT146, KEYINPUT147, KEYINPUT148, KEYINPUT149, KEYINPUT150,
         KEYINPUT151, KEYINPUT152, KEYINPUT153, KEYINPUT154, KEYINPUT155,
         KEYINPUT156, KEYINPUT157, KEYINPUT158, KEYINPUT159, KEYINPUT160,
         KEYINPUT161, KEYINPUT162, KEYINPUT163, KEYINPUT164, KEYINPUT165,
         KEYINPUT166, KEYINPUT167, KEYINPUT168, KEYINPUT169, KEYINPUT170,
         KEYINPUT171, KEYINPUT172, KEYINPUT173, KEYINPUT174, KEYINPUT175,
         KEYINPUT176, KEYINPUT177, KEYINPUT178, KEYINPUT179, KEYINPUT180,
         KEYINPUT181, KEYINPUT182, KEYINPUT183, KEYINPUT184, KEYINPUT185;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
         G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552,
         G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528,
         G526, G524, G279, G436, G478, G522, G402, G404, G406, G408, G410,
         G432, G446, G284, G286, G289, G292, G341, G281, G453, G278, G373,
         G246, G258, G264, G270, G388, G391, G394, G397, G376, G379, G382,
         G385, G412_enc, G414_enc, G416_enc, G249, G295, G324, G252, G276,         
         G310, G313, G316, G319, G327, G330, G333, G336, G418_enc, G273, G298, 
         G301, G304, G307, G344, G422, G469, G419, G471, G359, G362, G365, G368, 
         G347, G350, G353, G356, G321, G338, G370, G399;

  wire   n3797, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018;

  INV_X4 U2579 ( .A(G18), .ZN(n3844) );
  BUF_X1 U2580 ( .A(G1459), .Z(G450) );
  BUF_X1 U2581 ( .A(G1469), .Z(G448) );
  BUF_X1 U2582 ( .A(G1480), .Z(G444) );
  BUF_X1 U2583 ( .A(G1486), .Z(G442) );
  BUF_X1 U2584 ( .A(G1492), .Z(G440) );
  BUF_X1 U2585 ( .A(G1496), .Z(G438) );
  BUF_X1 U2586 ( .A(G2208), .Z(G496) );
  BUF_X1 U2587 ( .A(G2218), .Z(G494) );
  BUF_X1 U2588 ( .A(G2224), .Z(G492) );
  BUF_X1 U2589 ( .A(G2230), .Z(G490) );
  BUF_X1 U2590 ( .A(G2236), .Z(G488) );
  BUF_X1 U2591 ( .A(G2239), .Z(G486) );
  BUF_X1 U2592 ( .A(G2247), .Z(G484) );
  BUF_X1 U2593 ( .A(G2253), .Z(G482) );
  BUF_X1 U2594 ( .A(G2256), .Z(G480) );
  BUF_X1 U2595 ( .A(G3698), .Z(G560) );
  BUF_X1 U2596 ( .A(G3701), .Z(G542) );
  BUF_X1 U2597 ( .A(G3705), .Z(G558) );
  BUF_X1 U2598 ( .A(G3711), .Z(G556) );
  BUF_X1 U2599 ( .A(G3717), .Z(G554) );
  BUF_X1 U2600 ( .A(G3723), .Z(G552) );
  BUF_X1 U2601 ( .A(G3729), .Z(G550) );
  BUF_X1 U2602 ( .A(G3737), .Z(G548) );
  BUF_X1 U2603 ( .A(G3743), .Z(G546) );
  BUF_X1 U2604 ( .A(G3749), .Z(G544) );
  BUF_X1 U2605 ( .A(G4393), .Z(G540) );
  BUF_X1 U2606 ( .A(G4400), .Z(G538) );
  BUF_X1 U2607 ( .A(G4405), .Z(G536) );
  BUF_X1 U2608 ( .A(G4410), .Z(G534) );
  BUF_X1 U2609 ( .A(G4415), .Z(G532) );
  BUF_X1 U2610 ( .A(G4420), .Z(G530) );
  BUF_X1 U2611 ( .A(G4427), .Z(G528) );
  BUF_X1 U2612 ( .A(G4432), .Z(G526) );
  BUF_X1 U2613 ( .A(G4437), .Z(G524) );
  BUF_X1 U2614 ( .A(G1462), .Z(G436) );
  BUF_X1 U2615 ( .A(G2211), .Z(G478) );
  BUF_X1 U2616 ( .A(G4394), .Z(G522) );
  BUF_X1 U2617 ( .A(G106), .Z(G446) );
  BUF_X1 U2618 ( .A(G279), .Z(G341) );
  BUF_X1 U2619 ( .A(G279), .Z(G286) );
  INV_X1 U2620 ( .A(G1), .ZN(n3797) );
  INV_X1 U2621 ( .A(n3797), .ZN(G2) );
  INV_X1 U2622 ( .A(n3797), .ZN(G3) );
  INV_X1 U2623 ( .A(n3797), .ZN(G453) );
  INV_X1 U2624 ( .A(n3797), .ZN(G432) );
  BUF_X1 U2625 ( .A(G471), .Z(G419) );
  BUF_X1 U2626 ( .A(G469), .Z(G422) );
  BUF_X1 U2627 ( .A(G292), .Z(G281) );
  BUF_X1 U2628 ( .A(G289), .Z(G284) );
  XNOR2_X1 U2629 ( .A(n3806), .B(n3807), .ZN(G471) );
  NAND2_X1 U2630 ( .A1(n3808), .A2(n3809), .ZN(G469) );
  NAND3_X1 U2631 ( .A1(n3810), .A2(n3811), .A3(KEYINPUT142), .ZN(n3809) );
  NAND2_X1 U2632 ( .A1(n3812), .A2(n3813), .ZN(n3811) );
  NAND2_X1 U2633 ( .A1(n3806), .A2(n3814), .ZN(n3813) );
  OR2_X1 U2634 ( .A1(n3815), .A2(n3806), .ZN(n3808) );
  NOR3_X1 U2635 ( .A1(n3816), .A2(KEYINPUT14), .A3(n3817), .ZN(G418_enc) );
  NOR3_X1 U2636 ( .A1(n3818), .A2(n3819), .A3(n3820), .ZN(n3817) );
  NOR2_X1 U2637 ( .A1(KEYINPUT44), .A2(n3821), .ZN(n3820) );
  NOR2_X1 U2638 ( .A1(G410), .A2(G408), .ZN(n3821) );
  NOR2_X1 U2639 ( .A1(KEYINPUT43), .A2(n3822), .ZN(n3819) );
  NOR2_X1 U2640 ( .A1(G406), .A2(G404), .ZN(n3822) );
  NOR2_X1 U2641 ( .A1(KEYINPUT24), .A2(n3823), .ZN(n3818) );
  NOR3_X1 U2642 ( .A1(n3824), .A2(n3825), .A3(n3826), .ZN(n3823) );
  INV_X1 U2643 ( .A(KEYINPUT13), .ZN(n3816) );
  AND2_X1 U2644 ( .A1(KEYINPUT139), .A2(n3824), .ZN(G416_enc) );
  NOR2_X1 U2645 ( .A1(KEYINPUT136), .A2(n3827), .ZN(n3824) );
  NOR4_X1 U2646 ( .A1(n3828), .A2(n3829), .A3(n3830), .A4(n3831), .ZN(n3827) );
  XNOR2_X1 U2647 ( .A(n3832), .B(n3833), .ZN(n3831) );
  XNOR2_X1 U2648 ( .A(n3834), .B(n3835), .ZN(n3833) );
  XOR2_X1 U2649 ( .A(n3836), .B(n3837), .Z(n3834) );
  XOR2_X1 U2650 ( .A(n3838), .B(n3839), .Z(n3837) );
  XOR2_X1 U2651 ( .A(n3840), .B(n3841), .Z(n3839) );
  NAND2_X1 U2652 ( .A1(n3842), .A2(n3843), .ZN(n3841) );
  NAND2_X1 U2653 ( .A1(G44), .A2(n3844), .ZN(n3843) );
  NAND2_X1 U2654 ( .A1(G208), .A2(G18), .ZN(n3842) );
  XOR2_X1 U2655 ( .A(n3845), .B(n3846), .Z(n3838) );
  XOR2_X1 U2656 ( .A(n3847), .B(n3848), .Z(n3836) );
  XNOR2_X1 U2657 ( .A(n3849), .B(n3850), .ZN(n3848) );
  XOR2_X1 U2658 ( .A(n3851), .B(n3852), .Z(n3847) );
  XOR2_X1 U2659 ( .A(n3853), .B(n3854), .Z(n3830) );
  XOR2_X1 U2660 ( .A(n3855), .B(n3856), .Z(n3854) );
  XOR2_X1 U2661 ( .A(n3857), .B(n3858), .Z(n3856) );
  NAND3_X1 U2662 ( .A1(n3859), .A2(n3860), .A3(G18), .ZN(n3855) );
  XOR2_X1 U2663 ( .A(G165), .B(G164), .Z(n3859) );
  XOR2_X1 U2664 ( .A(n3861), .B(n3862), .Z(n3853) );
  NOR2_X1 U2665 ( .A1(n3863), .A2(n3864), .ZN(n3862) );
  NOR3_X1 U2666 ( .A1(n3865), .A2(n3866), .A3(n3867), .ZN(n3864) );
  AND2_X1 U2667 ( .A1(n3860), .A2(G170), .ZN(n3867) );
  NOR2_X1 U2668 ( .A1(n3868), .A2(n3869), .ZN(n3863) );
  NOR2_X1 U2669 ( .A1(G170), .A2(n3866), .ZN(n3868) );
  XNOR2_X1 U2670 ( .A(n3870), .B(n3871), .ZN(n3861) );
  XOR2_X1 U2671 ( .A(n3872), .B(n3873), .Z(n3829) );
  XOR2_X1 U2672 ( .A(n3874), .B(n3875), .Z(n3873) );
  XOR2_X1 U2673 ( .A(n3876), .B(n3877), .Z(n3872) );
  XOR2_X1 U2674 ( .A(n3878), .B(n3879), .Z(n3877) );
  XOR2_X1 U2675 ( .A(n3880), .B(n3881), .Z(n3879) );
  XNOR2_X1 U2676 ( .A(n3882), .B(n3883), .ZN(n3878) );
  NOR2_X1 U2677 ( .A1(n3884), .A2(n3885), .ZN(n3883) );
  NOR2_X1 U2678 ( .A1(G18), .A2(G141), .ZN(n3885) );
  NOR2_X1 U2679 ( .A1(G181), .A2(n3844), .ZN(n3884) );
  XOR2_X1 U2680 ( .A(n3886), .B(n3887), .Z(n3876) );
  XOR2_X1 U2681 ( .A(n3888), .B(n3889), .Z(n3887) );
  XOR2_X1 U2682 ( .A(n3890), .B(n3891), .Z(n3886) );
  XNOR2_X1 U2683 ( .A(n3892), .B(n3893), .ZN(n3828) );
  XNOR2_X1 U2684 ( .A(n3894), .B(n3895), .ZN(n3892) );
  XOR2_X1 U2685 ( .A(n3896), .B(n3897), .Z(n3894) );
  XOR2_X1 U2686 ( .A(n3898), .B(n3899), .Z(n3897) );
  XOR2_X1 U2687 ( .A(n3900), .B(n3901), .Z(n3899) );
  NOR2_X1 U2688 ( .A1(n3902), .A2(n3903), .ZN(n3901) );
  NOR2_X1 U2689 ( .A1(G18), .A2(G115), .ZN(n3903) );
  NOR2_X1 U2690 ( .A1(G197), .A2(n3844), .ZN(n3902) );
  XNOR2_X1 U2691 ( .A(n3904), .B(n3905), .ZN(n3898) );
  XOR2_X1 U2692 ( .A(n3906), .B(n3907), .Z(n3896) );
  XNOR2_X1 U2693 ( .A(n3908), .B(n3909), .ZN(n3907) );
  XNOR2_X1 U2694 ( .A(n3910), .B(n3911), .ZN(n3906) );
  AND2_X1 U2695 ( .A1(KEYINPUT141), .A2(n3826), .ZN(G414_enc) );
  NOR2_X1 U2696 ( .A1(KEYINPUT140), .A2(n3912), .ZN(n3826) );
  NOR4_X1 U2697 ( .A1(n3913), .A2(n3914), .A3(n3915), .A4(n3916), .ZN(n3912) );
  XOR2_X1 U2698 ( .A(n3917), .B(n3918), .Z(n3916) );
  XOR2_X1 U2699 ( .A(n3919), .B(n3920), .Z(n3918) );
  XNOR2_X1 U2700 ( .A(n3921), .B(n3922), .ZN(n3920) );
  XNOR2_X1 U2701 ( .A(n3923), .B(n3924), .ZN(n3919) );
  NAND2_X1 U2702 ( .A1(n3925), .A2(n3926), .ZN(n3923) );
  NAND2_X1 U2703 ( .A1(n3927), .A2(n3844), .ZN(n3926) );
  XNOR2_X1 U2704 ( .A(n3928), .B(G82), .ZN(n3927) );
  NAND2_X1 U2705 ( .A1(n3929), .A2(G18), .ZN(n3925) );
  XOR2_X1 U2706 ( .A(G2208), .B(n3928), .Z(n3929) );
  XOR2_X1 U2707 ( .A(n3930), .B(n3931), .Z(n3928) );
  XOR2_X1 U2708 ( .A(n3932), .B(n3933), .Z(n3917) );
  XOR2_X1 U2709 ( .A(n3934), .B(n3935), .Z(n3933) );
  XOR2_X1 U2710 ( .A(n3936), .B(n3937), .Z(n3932) );
  XOR2_X1 U2711 ( .A(n3938), .B(n3939), .Z(n3915) );
  XOR2_X1 U2712 ( .A(n3940), .B(n3941), .Z(n3939) );
  XOR2_X1 U2713 ( .A(n3942), .B(n3943), .Z(n3941) );
  XNOR2_X1 U2714 ( .A(n3944), .B(n3945), .ZN(n3940) );
  XOR2_X1 U2715 ( .A(n3946), .B(n3947), .Z(n3938) );
  XOR2_X1 U2716 ( .A(n3948), .B(n3949), .Z(n3947) );
  NAND2_X1 U2717 ( .A1(n3950), .A2(n3951), .ZN(n3949) );
  NAND2_X1 U2718 ( .A1(n3952), .A2(n3844), .ZN(n3951) );
  XOR2_X1 U2719 ( .A(n3953), .B(n3954), .Z(n3952) );
  XNOR2_X1 U2720 ( .A(G70), .B(G69), .ZN(n3954) );
  NAND2_X1 U2721 ( .A1(n3955), .A2(G18), .ZN(n3950) );
  XOR2_X1 U2722 ( .A(n3953), .B(n3956), .Z(n3955) );
  XNOR2_X1 U2723 ( .A(G3701), .B(G3698), .ZN(n3956) );
  XNOR2_X1 U2724 ( .A(n3957), .B(n3958), .ZN(n3946) );
  XOR2_X1 U2725 ( .A(n3959), .B(n3960), .Z(n3914) );
  XOR2_X1 U2726 ( .A(n3961), .B(n3962), .Z(n3960) );
  XOR2_X1 U2727 ( .A(n3963), .B(n3964), .Z(n3962) );
  XNOR2_X1 U2728 ( .A(n3965), .B(n3966), .ZN(n3961) );
  XOR2_X1 U2729 ( .A(n3967), .B(n3968), .Z(n3959) );
  XNOR2_X1 U2730 ( .A(n3969), .B(n3970), .ZN(n3968) );
  XNOR2_X1 U2731 ( .A(n3971), .B(n3972), .ZN(n3967) );
  NAND2_X1 U2732 ( .A1(n3973), .A2(n3974), .ZN(n3971) );
  NAND2_X1 U2733 ( .A1(n3975), .A2(n3844), .ZN(n3974) );
  XNOR2_X1 U2734 ( .A(n3976), .B(G58), .ZN(n3975) );
  NAND2_X1 U2735 ( .A1(n3977), .A2(G18), .ZN(n3973) );
  XOR2_X1 U2736 ( .A(G4393), .B(n3976), .Z(n3977) );
  XOR2_X1 U2737 ( .A(n3978), .B(n3979), .Z(n3976) );
  XOR2_X1 U2738 ( .A(n3980), .B(n3981), .Z(n3913) );
  XOR2_X1 U2739 ( .A(n3982), .B(n3983), .Z(n3981) );
  NAND2_X1 U2740 ( .A1(n3984), .A2(n3985), .ZN(n3983) );
  NAND2_X1 U2741 ( .A1(n3986), .A2(n3844), .ZN(n3985) );
  XOR2_X1 U2742 ( .A(n3987), .B(n3988), .Z(n3986) );
  XNOR2_X1 U2743 ( .A(G1455), .B(G2204), .ZN(n3988) );
  NAND2_X1 U2744 ( .A1(n3989), .A2(G18), .ZN(n3984) );
  XOR2_X1 U2745 ( .A(n3987), .B(n3990), .Z(n3989) );
  XNOR2_X1 U2746 ( .A(G1496), .B(G1492), .ZN(n3990) );
  XNOR2_X1 U2747 ( .A(n3991), .B(n3992), .ZN(n3980) );
  NAND2_X1 U2748 ( .A1(n3993), .A2(n3994), .ZN(n3991) );
  NAND2_X1 U2749 ( .A1(n3995), .A2(n3844), .ZN(n3994) );
  XNOR2_X1 U2750 ( .A(n3996), .B(G114), .ZN(n3995) );
  NAND2_X1 U2751 ( .A1(n3997), .A2(G18), .ZN(n3993) );
  XNOR2_X1 U2752 ( .A(G1459), .B(n3998), .ZN(n3997) );
  INV_X1 U2753 ( .A(n3996), .ZN(n3998) );
  XNOR2_X1 U2754 ( .A(n3999), .B(n4000), .ZN(n3996) );
  AND2_X1 U2755 ( .A1(KEYINPUT138), .A2(n3825), .ZN(G412_enc) );
  NOR2_X1 U2756 ( .A1(KEYINPUT137), .A2(n4001), .ZN(n3825) );
  NOR4_X1 U2757 ( .A1(n4002), .A2(n4003), .A3(n4004), .A4(n4005), .ZN(n4001) );
  XOR2_X1 U2758 ( .A(n4006), .B(n4007), .Z(n4005) );
  XOR2_X1 U2759 ( .A(n4008), .B(n4009), .Z(n4007) );
  XNOR2_X1 U2760 ( .A(n4010), .B(n4011), .ZN(n4009) );
  XOR2_X1 U2761 ( .A(n4012), .B(n4013), .Z(n4008) );
  XOR2_X1 U2762 ( .A(n4014), .B(n4015), .Z(n4006) );
  XNOR2_X1 U2763 ( .A(n4016), .B(n4017), .ZN(n4015) );
  NAND2_X1 U2764 ( .A1(n4018), .A2(n4019), .ZN(n4017) );
  NAND2_X1 U2765 ( .A1(n4020), .A2(n3844), .ZN(n4019) );
  XNOR2_X1 U2766 ( .A(G141), .B(n4021), .ZN(n4020) );
  NAND2_X1 U2767 ( .A1(n4022), .A2(G18), .ZN(n4018) );
  XNOR2_X1 U2768 ( .A(n4021), .B(G161), .ZN(n4022) );
  XNOR2_X1 U2769 ( .A(n4023), .B(n4024), .ZN(n4021) );
  XNOR2_X1 U2770 ( .A(n4025), .B(n4026), .ZN(n4014) );
  XOR2_X1 U2771 ( .A(n4027), .B(n4028), .Z(n4004) );
  XOR2_X1 U2772 ( .A(n4029), .B(n4030), .Z(n4028) );
  XNOR2_X1 U2773 ( .A(n4031), .B(n4032), .ZN(n4030) );
  NAND2_X1 U2774 ( .A1(KEYINPUT1), .A2(n3860), .ZN(n4029) );
  XOR2_X1 U2775 ( .A(n4033), .B(n4034), .Z(n4027) );
  XOR2_X1 U2776 ( .A(n4035), .B(n4036), .Z(n4034) );
  NAND3_X1 U2777 ( .A1(n4037), .A2(n3860), .A3(G18), .ZN(n4035) );
  XOR2_X1 U2778 ( .A(G212), .B(G211), .Z(n4037) );
  XNOR2_X1 U2779 ( .A(n4038), .B(n4039), .ZN(n4033) );
  XOR2_X1 U2780 ( .A(n4040), .B(n4041), .Z(n4003) );
  XOR2_X1 U2781 ( .A(n4042), .B(n4043), .Z(n4041) );
  XOR2_X1 U2782 ( .A(n4044), .B(n4045), .Z(n4043) );
  XOR2_X1 U2783 ( .A(n4046), .B(n4047), .Z(n4045) );
  NAND2_X1 U2784 ( .A1(n4048), .A2(n4049), .ZN(n4047) );
  NAND2_X1 U2785 ( .A1(n4050), .A2(n3844), .ZN(n4049) );
  XOR2_X1 U2786 ( .A(G44), .B(n4051), .Z(n4050) );
  NAND2_X1 U2787 ( .A1(n4052), .A2(G18), .ZN(n4048) );
  XOR2_X1 U2788 ( .A(G239), .B(n4051), .Z(n4052) );
  XNOR2_X1 U2789 ( .A(n4053), .B(n4054), .ZN(n4044) );
  XOR2_X1 U2790 ( .A(n4055), .B(n4056), .Z(n4042) );
  XNOR2_X1 U2791 ( .A(n4057), .B(n4058), .ZN(n4056) );
  XNOR2_X1 U2792 ( .A(n4059), .B(n4060), .ZN(n4055) );
  XOR2_X1 U2793 ( .A(n4061), .B(n4062), .Z(n4002) );
  XOR2_X1 U2794 ( .A(n4063), .B(n4064), .Z(n4062) );
  XOR2_X1 U2795 ( .A(n4065), .B(n4066), .Z(n4064) );
  NAND2_X1 U2796 ( .A1(n4067), .A2(n4068), .ZN(n4066) );
  NAND2_X1 U2797 ( .A1(n4069), .A2(n3844), .ZN(n4068) );
  XNOR2_X1 U2798 ( .A(G115), .B(n4070), .ZN(n4069) );
  NAND2_X1 U2799 ( .A1(n4071), .A2(G18), .ZN(n4067) );
  XNOR2_X1 U2800 ( .A(n4070), .B(G227), .ZN(n4071) );
  XNOR2_X1 U2801 ( .A(n4072), .B(n4073), .ZN(n4070) );
  XNOR2_X1 U2802 ( .A(n4074), .B(n4075), .ZN(n4063) );
  XOR2_X1 U2803 ( .A(n4076), .B(n4077), .Z(n4061) );
  XNOR2_X1 U2804 ( .A(n4078), .B(n4079), .ZN(n4077) );
  XNOR2_X1 U2805 ( .A(n4080), .B(n4081), .ZN(n4076) );
  NAND4_X1 U2806 ( .A1(G199), .A2(G188), .A3(G172), .A4(G162), .ZN(G410) );
  NAND4_X1 U2807 ( .A1(G186), .A2(G185), .A3(G183), .A4(G182), .ZN(G408) );
  NAND4_X1 U2808 ( .A1(G230), .A2(G218), .A3(G210), .A4(G152), .ZN(G406) );
  NAND4_X1 U2809 ( .A1(G240), .A2(G228), .A3(G184), .A4(G150), .ZN(G404) );
  OR2_X1 U2810 ( .A1(G5), .A2(G57), .ZN(G402) );
  NAND2_X1 U2811 ( .A1(n4082), .A2(n4083), .ZN(G399) );
  NAND2_X1 U2812 ( .A1(n4084), .A2(n4085), .ZN(n4083) );
  XOR2_X1 U2813 ( .A(n4086), .B(n4087), .Z(n4084) );
  XOR2_X1 U2814 ( .A(n4088), .B(n4089), .Z(n4087) );
  NAND2_X1 U2815 ( .A1(n4090), .A2(KEYINPUT164), .ZN(n4088) );
  XNOR2_X1 U2816 ( .A(n4091), .B(n4092), .ZN(n4090) );
  NOR4_X1 U2817 ( .A1(KEYINPUT133), .A2(n4093), .A3(n4094), .A4(n4095), .ZN(n4092) );
  AND2_X1 U2818 ( .A1(n4096), .A2(n4097), .ZN(n4095) );
  XNOR2_X1 U2819 ( .A(n4098), .B(n4099), .ZN(n4086) );
  NAND4_X1 U2820 ( .A1(n4100), .A2(n4101), .A3(n4102), .A4(n4103), .ZN(n4099) );
  NAND2_X1 U2821 ( .A1(n4094), .A2(n4104), .ZN(n4103) );
  NOR2_X1 U2822 ( .A1(n4105), .A2(n4106), .ZN(n4094) );
  NOR2_X1 U2823 ( .A1(KEYINPUT72), .A2(KEYINPUT182), .ZN(n4102) );
  NAND2_X1 U2824 ( .A1(n4097), .A2(n4107), .ZN(n4101) );
  NAND2_X1 U2825 ( .A1(n4108), .A2(G4526), .ZN(n4082) );
  XOR2_X1 U2826 ( .A(n4109), .B(n4110), .Z(n4108) );
  XOR2_X1 U2827 ( .A(n4111), .B(n4112), .Z(n4110) );
  NOR4_X1 U2828 ( .A1(KEYINPUT71), .A2(KEYINPUT181), .A3(n4113), .A4(n4114),  .ZN(n4112) );
  INV_X1 U2829 ( .A(n4115), .ZN(n4113) );
  XOR2_X1 U2830 ( .A(n4089), .B(n4116), .Z(n4109) );
  NOR2_X1 U2831 ( .A1(n4117), .A2(n4118), .ZN(n4116) );
  NOR3_X1 U2832 ( .A1(n4119), .A2(KEYINPUT132), .A3(n4093), .ZN(n4118) );
  NOR2_X1 U2833 ( .A1(n4120), .A2(n4121), .ZN(n4117) );
  NOR3_X1 U2834 ( .A1(n4096), .A2(KEYINPUT132), .A3(n4093), .ZN(n4121) );
  INV_X1 U2835 ( .A(n4119), .ZN(n4120) );
  XNOR2_X1 U2836 ( .A(n4122), .B(n4123), .ZN(n4089) );
  XOR2_X1 U2837 ( .A(n4124), .B(n4125), .Z(n4122) );
  NOR2_X1 U2838 ( .A1(n4126), .A2(n4127), .ZN(n4125) );
  NOR2_X1 U2839 ( .A1(n4128), .A2(n4129), .ZN(n4127) );
  XOR2_X1 U2840 ( .A(n4130), .B(n4131), .Z(n4129) );
  XNOR2_X1 U2841 ( .A(n4132), .B(n4133), .ZN(n4131) );
  NAND3_X1 U2842 ( .A1(n4134), .A2(n4135), .A3(n4136), .ZN(n4132) );
  NAND3_X1 U2843 ( .A1(n4137), .A2(n4138), .A3(n4139), .ZN(n4136) );
  INV_X1 U2844 ( .A(n4140), .ZN(n4135) );
  XOR2_X1 U2845 ( .A(n4141), .B(n4142), .Z(n4130) );
  NOR3_X1 U2846 ( .A1(n4143), .A2(KEYINPUT178), .A3(n4140), .ZN(n4142) );
  NOR2_X1 U2847 ( .A1(n4144), .A2(n4145), .ZN(n4128) );
  NOR3_X1 U2848 ( .A1(n4146), .A2(n4144), .A3(n4145), .ZN(n4126) );
  NOR2_X1 U2849 ( .A1(KEYINPUT120), .A2(n4085), .ZN(n4144) );
  XOR2_X1 U2850 ( .A(n4147), .B(n4148), .Z(n4146) );
  NOR2_X1 U2851 ( .A1(KEYINPUT179), .A2(n4143), .ZN(n4148) );
  NAND2_X1 U2852 ( .A1(n4149), .A2(n4150), .ZN(n4147) );
  NAND2_X1 U2853 ( .A1(n4151), .A2(n4152), .ZN(n4150) );
  NAND2_X1 U2854 ( .A1(n4153), .A2(n4154), .ZN(n4151) );
  NAND2_X1 U2855 ( .A1(n4155), .A2(n4133), .ZN(n4154) );
  NAND2_X1 U2856 ( .A1(n4156), .A2(n4157), .ZN(n4153) );
  NAND2_X1 U2857 ( .A1(n4158), .A2(n4159), .ZN(n4149) );
  NAND2_X1 U2858 ( .A1(n4160), .A2(n4161), .ZN(n4158) );
  NAND2_X1 U2859 ( .A1(n4156), .A2(n4155), .ZN(n4161) );
  XNOR2_X1 U2860 ( .A(n4162), .B(n4137), .ZN(n4155) );
  INV_X1 U2861 ( .A(n4133), .ZN(n4156) );
  NAND2_X1 U2862 ( .A1(n4133), .A2(n4157), .ZN(n4160) );
  NAND2_X1 U2863 ( .A1(n4134), .A2(n4163), .ZN(n4157) );
  NAND2_X1 U2864 ( .A1(n4139), .A2(n4137), .ZN(n4163) );
  XOR2_X1 U2865 ( .A(n4164), .B(n4165), .Z(n4133) );
  NAND2_X1 U2866 ( .A1(n4138), .A2(n4166), .ZN(n4164) );
  NAND2_X1 U2867 ( .A1(n4167), .A2(n4168), .ZN(n4166) );
  NAND3_X1 U2868 ( .A1(n4169), .A2(n4170), .A3(n4171), .ZN(n4124) );
  NAND2_X1 U2869 ( .A1(n4172), .A2(n4173), .ZN(n4171) );
  XNOR2_X1 U2870 ( .A(n4174), .B(n4096), .ZN(n4172) );
  NAND3_X1 U2871 ( .A1(n4104), .A2(n4106), .A3(n4174), .ZN(n4170) );
  NAND2_X1 U2872 ( .A1(n4175), .A2(n4107), .ZN(n4169) );
  INV_X1 U2873 ( .A(n4174), .ZN(n4175) );
  XOR2_X1 U2874 ( .A(n4176), .B(n4177), .Z(n4174) );
  XNOR2_X1 U2875 ( .A(n4178), .B(n4179), .ZN(G397) );
  NAND2_X1 U2876 ( .A1(n4180), .A2(n4181), .ZN(n4178) );
  NAND2_X1 U2877 ( .A1(G4526), .A2(n4177), .ZN(n4181) );
  XNOR2_X1 U2878 ( .A(n4106), .B(n4182), .ZN(G394) );
  XNOR2_X1 U2879 ( .A(n4104), .B(n4183), .ZN(G391) );
  NOR3_X1 U2880 ( .A1(n4184), .A2(KEYINPUT131), .A3(n4093), .ZN(n4183) );
  NOR2_X1 U2881 ( .A1(n4106), .A2(n4185), .ZN(n4184) );
  XNOR2_X1 U2882 ( .A(n4186), .B(n4123), .ZN(G388) );
  NAND3_X1 U2883 ( .A1(n4100), .A2(n4187), .A3(n4188), .ZN(n4186) );
  NOR3_X1 U2884 ( .A1(KEYINPUT130), .A2(KEYINPUT70), .A3(KEYINPUT176), .ZN(n4188) );
  NAND2_X1 U2885 ( .A1(n4182), .A2(n4107), .ZN(n4187) );
  INV_X1 U2886 ( .A(n4185), .ZN(n4182) );
  NAND2_X1 U2887 ( .A1(n4119), .A2(n4189), .ZN(n4185) );
  NAND2_X1 U2888 ( .A1(n4098), .A2(n4085), .ZN(n4189) );
  NAND2_X1 U2889 ( .A1(n4098), .A2(n4190), .ZN(n4119) );
  NAND2_X1 U2890 ( .A1(n4177), .A2(n4176), .ZN(n4190) );
  XOR2_X1 U2891 ( .A(n4168), .B(n4191), .Z(G385) );
  XOR2_X1 U2892 ( .A(n4192), .B(n4167), .Z(G382) );
  NAND2_X1 U2893 ( .A1(n4141), .A2(n4193), .ZN(n4192) );
  NAND2_X1 U2894 ( .A1(n4191), .A2(n4152), .ZN(n4193) );
  XOR2_X1 U2895 ( .A(n4194), .B(n4137), .Z(G379) );
  NOR2_X1 U2896 ( .A1(n4195), .A2(n4162), .ZN(n4194) );
  NOR2_X1 U2897 ( .A1(n4191), .A2(n4138), .ZN(n4195) );
  XOR2_X1 U2898 ( .A(n4196), .B(n4165), .Z(G376) );
  NAND3_X1 U2899 ( .A1(n4197), .A2(n4198), .A3(n4199), .ZN(n4196) );
  INV_X1 U2900 ( .A(n4143), .ZN(n4199) );
  NAND2_X1 U2901 ( .A1(KEYINPUT169), .A2(n4191), .ZN(n4198) );
  OR2_X1 U2902 ( .A1(n4191), .A2(n4200), .ZN(n4197) );
  NOR2_X1 U2903 ( .A1(KEYINPUT168), .A2(n4140), .ZN(n4200) );
  XNOR2_X1 U2904 ( .A(n4085), .B(n4177), .ZN(G373) );
  INV_X1 U2905 ( .A(G4526), .ZN(n4085) );
  NAND2_X1 U2906 ( .A1(n4201), .A2(n4202), .ZN(G370) );
  NAND2_X1 U2907 ( .A1(n4203), .A2(n4204), .ZN(n4202) );
  XOR2_X1 U2908 ( .A(n4205), .B(n4206), .Z(n4203) );
  XNOR2_X1 U2909 ( .A(n4207), .B(n4208), .ZN(n4206) );
  XOR2_X1 U2910 ( .A(n4209), .B(n4210), .Z(n4208) );
  NOR4_X1 U2911 ( .A1(KEYINPUT154), .A2(KEYINPUT113), .A3(n4211), .A4(n4212),  .ZN(n4210) );
  NOR2_X1 U2912 ( .A1(n4209), .A2(n4213), .ZN(n4211) );
  AND2_X1 U2913 ( .A1(n4214), .A2(n4215), .ZN(n4209) );
  XOR2_X1 U2914 ( .A(n4216), .B(n4217), .Z(n4205) );
  NAND2_X1 U2915 ( .A1(n4218), .A2(n4219), .ZN(n4201) );
  XOR2_X1 U2916 ( .A(n4220), .B(n4221), .Z(n4218) );
  XNOR2_X1 U2917 ( .A(n4214), .B(n4222), .ZN(n4221) );
  XNOR2_X1 U2918 ( .A(n4223), .B(n4224), .ZN(n4222) );
  XNOR2_X1 U2919 ( .A(n4217), .B(n4225), .ZN(n4220) );
  NOR2_X1 U2920 ( .A1(KEYINPUT114), .A2(n4226), .ZN(n4225) );
  XNOR2_X1 U2921 ( .A(n4227), .B(n4228), .ZN(n4217) );
  XOR2_X1 U2922 ( .A(n4229), .B(n4230), .Z(n4228) );
  XNOR2_X1 U2923 ( .A(n4231), .B(n4232), .ZN(n4230) );
  NAND2_X1 U2924 ( .A1(n4233), .A2(n4234), .ZN(n4229) );
  NAND2_X1 U2925 ( .A1(n4235), .A2(n4236), .ZN(n4234) );
  INV_X1 U2926 ( .A(n4237), .ZN(n4236) );
  XOR2_X1 U2927 ( .A(n4238), .B(n4239), .Z(n4235) );
  XOR2_X1 U2928 ( .A(n4240), .B(n4241), .Z(n4239) );
  NOR3_X1 U2929 ( .A1(n4242), .A2(n4243), .A3(n4244), .ZN(n4240) );
  NOR3_X1 U2930 ( .A1(n4245), .A2(n4246), .A3(n4247), .ZN(n4242) );
  INV_X1 U2931 ( .A(n4248), .ZN(n4247) );
  XOR2_X1 U2932 ( .A(n4249), .B(n4250), .Z(n4238) );
  NAND2_X1 U2933 ( .A1(n4251), .A2(n4237), .ZN(n4233) );
  NOR4_X1 U2934 ( .A1(n4252), .A2(n4253), .A3(KEYINPUT112), .A4(KEYINPUT60),  .ZN(n4237) );
  AND2_X1 U2935 ( .A1(n4254), .A2(n4204), .ZN(n4253) );
  INV_X1 U2936 ( .A(n4219), .ZN(n4204) );
  NOR4_X1 U2937 ( .A1(n4255), .A2(n4256), .A3(KEYINPUT106), .A4(KEYINPUT177),  .ZN(n4219) );
  AND2_X1 U2938 ( .A1(n4257), .A2(n4258), .ZN(n4256) );
  NAND3_X1 U2939 ( .A1(n4259), .A2(n4260), .A3(KEYINPUT156), .ZN(n4258) );
  NAND2_X1 U2940 ( .A1(KEYINPUT67), .A2(n4261), .ZN(n4257) );
  INV_X1 U2941 ( .A(n4145), .ZN(n4261) );
  OR3_X1 U2942 ( .A1(n4262), .A2(KEYINPUT92), .A3(n4263), .ZN(n4254) );
  INV_X1 U2943 ( .A(KEYINPUT90), .ZN(n4263) );
  XNOR2_X1 U2944 ( .A(n4264), .B(n4265), .ZN(n4251) );
  NAND3_X1 U2945 ( .A1(n4266), .A2(n4267), .A3(n4268), .ZN(n4265) );
  NAND2_X1 U2946 ( .A1(n4269), .A2(n4248), .ZN(n4268) );
  XNOR2_X1 U2947 ( .A(n4270), .B(n4271), .ZN(n4269) );
  NAND2_X1 U2948 ( .A1(n4243), .A2(n4271), .ZN(n4267) );
  OR3_X1 U2949 ( .A1(n4245), .A2(n4248), .A3(n4271), .ZN(n4266) );
  XNOR2_X1 U2950 ( .A(n4272), .B(n4241), .ZN(n4271) );
  XNOR2_X1 U2951 ( .A(n4273), .B(n4274), .ZN(n4241) );
  NAND2_X1 U2952 ( .A1(n4275), .A2(n4276), .ZN(n4273) );
  OR2_X1 U2953 ( .A1(n4277), .A2(n4278), .ZN(n4276) );
  XNOR2_X1 U2954 ( .A(n4279), .B(n4280), .ZN(n4227) );
  XNOR2_X1 U2955 ( .A(n4213), .B(n4281), .ZN(n4280) );
  XOR2_X1 U2956 ( .A(n4282), .B(n4232), .Z(G368) );
  NAND2_X1 U2957 ( .A1(n4283), .A2(n4284), .ZN(n4282) );
  NAND2_X1 U2958 ( .A1(n4279), .A2(n4285), .ZN(n4284) );
  XNOR2_X1 U2959 ( .A(n4281), .B(n4286), .ZN(G365) );
  XOR2_X1 U2960 ( .A(n4213), .B(n4287), .Z(G362) );
  NOR2_X1 U2961 ( .A1(KEYINPUT134), .A2(n4288), .ZN(n4287) );
  XNOR2_X1 U2962 ( .A(n4231), .B(n4289), .ZN(G359) );
  NOR4_X1 U2963 ( .A1(KEYINPUT73), .A2(KEYINPUT110), .A3(n4212), .A4(n4290),  .ZN(n4289) );
  NOR2_X1 U2964 ( .A1(n4291), .A2(n4213), .ZN(n4290) );
  INV_X1 U2965 ( .A(n4288), .ZN(n4291) );
  NAND2_X1 U2966 ( .A1(n4292), .A2(n4293), .ZN(n4288) );
  OR2_X1 U2967 ( .A1(n4286), .A2(n4294), .ZN(n4293) );
  NAND2_X1 U2968 ( .A1(n4207), .A2(n4295), .ZN(n4286) );
  NAND2_X1 U2969 ( .A1(n4296), .A2(n4223), .ZN(n4295) );
  NAND2_X1 U2970 ( .A1(n4223), .A2(n4297), .ZN(n4207) );
  NAND2_X1 U2971 ( .A1(n4279), .A2(n4232), .ZN(n4297) );
  INV_X1 U2972 ( .A(n4298), .ZN(n4223) );
  XNOR2_X1 U2973 ( .A(n4299), .B(n4278), .ZN(G356) );
  XOR2_X1 U2974 ( .A(n4300), .B(n4277), .Z(G353) );
  NOR2_X1 U2975 ( .A1(n4301), .A2(n4249), .ZN(n4300) );
  NOR2_X1 U2976 ( .A1(n4264), .A2(n4302), .ZN(n4301) );
  XNOR2_X1 U2977 ( .A(n4303), .B(n4248), .ZN(G350) );
  NAND2_X1 U2978 ( .A1(n4270), .A2(n4304), .ZN(n4303) );
  NAND2_X1 U2979 ( .A1(n4246), .A2(n4302), .ZN(n4304) );
  INV_X1 U2980 ( .A(n4275), .ZN(n4246) );
  XOR2_X1 U2981 ( .A(n4305), .B(n4274), .Z(G347) );
  NOR2_X1 U2982 ( .A1(n4306), .A2(n4307), .ZN(n4305) );
  NOR3_X1 U2983 ( .A1(n4302), .A2(KEYINPUT185), .A3(n4272), .ZN(n4307) );
  NOR3_X1 U2984 ( .A1(n4299), .A2(KEYINPUT184), .A3(n4250), .ZN(n4306) );
  OR2_X1 U2985 ( .A1(n4272), .A2(n4244), .ZN(n4250) );
  INV_X1 U2986 ( .A(n4302), .ZN(n4299) );
  NAND3_X1 U2987 ( .A1(n4308), .A2(n4309), .A3(n4310), .ZN(n4302) );
  NOR3_X1 U2988 ( .A1(KEYINPUT109), .A2(KEYINPUT59), .A3(KEYINPUT52), .ZN(n4310) );
  NAND2_X1 U2989 ( .A1(n4311), .A2(n4285), .ZN(n4309) );
  INV_X1 U2990 ( .A(n4296), .ZN(n4285) );
  OR2_X1 U2991 ( .A1(KEYINPUT91), .A2(n4262), .ZN(n4311) );
  INV_X1 U2992 ( .A(n4252), .ZN(n4308) );
  XNOR2_X1 U2993 ( .A(n4296), .B(n4279), .ZN(G344) );
  NOR4_X1 U2994 ( .A1(n4255), .A2(n4312), .A3(KEYINPUT101), .A4(KEYINPUT167),  .ZN(n4296) );
  NOR2_X1 U2995 ( .A1(n4191), .A2(n4313), .ZN(n4312) );
  AND3_X1 U2996 ( .A1(n4259), .A2(n4314), .A3(KEYINPUT155), .ZN(n4313) );
  NOR3_X1 U2997 ( .A1(KEYINPUT66), .A2(n4315), .A3(n4316), .ZN(n4191) );
  INV_X1 U2998 ( .A(n4317), .ZN(n4316) );
  INV_X1 U2999 ( .A(G15), .ZN(G279) );
  NAND2_X1 U3000 ( .A1(n4318), .A2(n4319), .ZN(G338) );
  NAND2_X1 U3001 ( .A1(n4320), .A2(n4321), .ZN(n4319) );
  XOR2_X1 U3002 ( .A(n4322), .B(n4323), .Z(n4320) );
  XNOR2_X1 U3003 ( .A(n4324), .B(n4325), .ZN(n4323) );
  XOR2_X1 U3004 ( .A(n4326), .B(n4327), .Z(n4322) );
  XOR2_X1 U3005 ( .A(n4328), .B(n4329), .Z(n4327) );
  NOR4_X1 U3006 ( .A1(KEYINPUT157), .A2(KEYINPUT124), .A3(n4330), .A4(n4331),  .ZN(n4329) );
  NOR2_X1 U3007 ( .A1(n4328), .A2(n4332), .ZN(n4330) );
  NOR2_X1 U3008 ( .A1(n4333), .A2(n4334), .ZN(n4328) );
  NAND2_X1 U3009 ( .A1(n4335), .A2(n4336), .ZN(n4318) );
  XOR2_X1 U3010 ( .A(n4337), .B(n4338), .Z(n4335) );
  XOR2_X1 U3011 ( .A(n4324), .B(n4339), .Z(n4338) );
  NOR2_X1 U3012 ( .A1(KEYINPUT125), .A2(n4340), .ZN(n4339) );
  XOR2_X1 U3013 ( .A(n4341), .B(n4342), .Z(n4324) );
  XNOR2_X1 U3014 ( .A(n4343), .B(n4344), .ZN(n4342) );
  XNOR2_X1 U3015 ( .A(n4345), .B(n4332), .ZN(n4344) );
  XNOR2_X1 U3016 ( .A(n4346), .B(n4347), .ZN(n4341) );
  XOR2_X1 U3017 ( .A(n4348), .B(n4349), .Z(n4346) );
  NAND2_X1 U3018 ( .A1(n4350), .A2(n4351), .ZN(n4348) );
  NAND3_X1 U3019 ( .A1(n4352), .A2(n4353), .A3(n3807), .ZN(n4351) );
  NAND2_X1 U3020 ( .A1(n3810), .A2(n4354), .ZN(n4353) );
  NAND2_X1 U3021 ( .A1(n4355), .A2(n3814), .ZN(n3810) );
  INV_X1 U3022 ( .A(n3812), .ZN(n4355) );
  NAND2_X1 U3023 ( .A1(n3815), .A2(n4356), .ZN(n4352) );
  XOR2_X1 U3024 ( .A(n3812), .B(n4357), .Z(n3815) );
  NOR2_X1 U3025 ( .A1(n4358), .A2(n4359), .ZN(n4357) );
  NAND2_X1 U3026 ( .A1(n3812), .A2(n4360), .ZN(n4350) );
  NAND2_X1 U3027 ( .A1(n3807), .A2(n4361), .ZN(n4360) );
  OR2_X1 U3028 ( .A1(n3814), .A2(n4356), .ZN(n4361) );
  INV_X1 U3029 ( .A(n4354), .ZN(n4356) );
  NAND2_X1 U3030 ( .A1(n4362), .A2(n4363), .ZN(n4354) );
  OR2_X1 U3031 ( .A1(KEYINPUT93), .A2(n4336), .ZN(n4363) );
  XOR2_X1 U3032 ( .A(n4333), .B(n4364), .Z(n4337) );
  XNOR2_X1 U3033 ( .A(n4365), .B(n4366), .ZN(n4364) );
  XNOR2_X1 U3034 ( .A(n4367), .B(n4368), .ZN(G336) );
  NAND2_X1 U3035 ( .A1(n4369), .A2(n4370), .ZN(n4367) );
  NAND2_X1 U3036 ( .A1(n4345), .A2(n4371), .ZN(n4370) );
  XNOR2_X1 U3037 ( .A(n4372), .B(n4373), .ZN(G333) );
  XNOR2_X1 U3038 ( .A(n4374), .B(n4375), .ZN(G330) );
  NOR2_X1 U3039 ( .A1(KEYINPUT143), .A2(n4376), .ZN(n4375) );
  XNOR2_X1 U3040 ( .A(n4349), .B(n4377), .ZN(G327) );
  NOR4_X1 U3041 ( .A1(KEYINPUT85), .A2(KEYINPUT127), .A3(n4331), .A4(n4378),  .ZN(n4377) );
  AND2_X1 U3042 ( .A1(n4376), .A2(n4374), .ZN(n4378) );
  NAND2_X1 U3043 ( .A1(n4379), .A2(n4380), .ZN(n4376) );
  OR2_X1 U3044 ( .A1(n4373), .A2(n4343), .ZN(n4380) );
  NAND2_X1 U3045 ( .A1(n4325), .A2(n4381), .ZN(n4373) );
  NAND2_X1 U3046 ( .A1(n4382), .A2(n4383), .ZN(n4381) );
  NAND2_X1 U3047 ( .A1(n4383), .A2(n4384), .ZN(n4325) );
  NAND2_X1 U3048 ( .A1(n4345), .A2(n4347), .ZN(n4384) );
  INV_X1 U3049 ( .A(n4366), .ZN(n4383) );
  XNOR2_X1 U3050 ( .A(n4382), .B(n4345), .ZN(G324) );
  INV_X1 U3051 ( .A(n4385), .ZN(n4345) );
  NAND2_X1 U3052 ( .A1(n4386), .A2(n4387), .ZN(G321) );
  NAND2_X1 U3053 ( .A1(n4388), .A2(n4389), .ZN(n4387) );
  XOR2_X1 U3054 ( .A(n4390), .B(n4391), .Z(n4388) );
  XOR2_X1 U3055 ( .A(n4392), .B(n4393), .Z(n4391) );
  NOR2_X1 U3056 ( .A1(n4394), .A2(n4395), .ZN(n4393) );
  NOR3_X1 U3057 ( .A1(n4396), .A2(KEYINPUT173), .A3(n4397), .ZN(n4395) );
  NOR2_X1 U3058 ( .A1(n4398), .A2(n4399), .ZN(n4394) );
  NOR3_X1 U3059 ( .A1(n4400), .A2(KEYINPUT173), .A3(n4397), .ZN(n4399) );
  XOR2_X1 U3060 ( .A(n4401), .B(n4402), .Z(n4390) );
  XOR2_X1 U3061 ( .A(n4403), .B(n4404), .Z(n4402) );
  NAND3_X1 U3062 ( .A1(n4405), .A2(n4406), .A3(n4407), .ZN(n4404) );
  NAND2_X1 U3063 ( .A1(n4408), .A2(n4409), .ZN(n4407) );
  NAND3_X1 U3064 ( .A1(n4410), .A2(n4411), .A3(n4412), .ZN(n4406) );
  NAND2_X1 U3065 ( .A1(n4413), .A2(n4414), .ZN(n4405) );
  INV_X1 U3066 ( .A(n4412), .ZN(n4414) );
  NAND3_X1 U3067 ( .A1(n4415), .A2(n4416), .A3(n4417), .ZN(n4403) );
  NOR3_X1 U3068 ( .A1(KEYINPUT103), .A2(KEYINPUT171), .A3(KEYINPUT150), .ZN(n4417) );
  INV_X1 U3069 ( .A(n4418), .ZN(n4415) );
  NAND2_X1 U3070 ( .A1(n4419), .A2(n4420), .ZN(n4386) );
  XOR2_X1 U3071 ( .A(n4421), .B(n4422), .Z(n4420) );
  XOR2_X1 U3072 ( .A(n4423), .B(n4424), .Z(n4422) );
  XNOR2_X1 U3073 ( .A(n4425), .B(n4426), .ZN(n4424) );
  NAND4_X1 U3074 ( .A1(n4427), .A2(n4428), .A3(n4429), .A4(n4430), .ZN(n4426) );
  NAND3_X1 U3075 ( .A1(n4413), .A2(n4431), .A3(n4432), .ZN(n4430) );
  NOR2_X1 U3076 ( .A1(KEYINPUT172), .A2(KEYINPUT104), .ZN(n4429) );
  NAND2_X1 U3077 ( .A1(n4433), .A2(n4410), .ZN(n4428) );
  XNOR2_X1 U3078 ( .A(n4434), .B(n4435), .ZN(n4423) );
  NOR4_X1 U3079 ( .A1(KEYINPUT174), .A2(n4397), .A3(n4433), .A4(n4436), .ZN(n4435) );
  NOR3_X1 U3080 ( .A1(n4434), .A2(n4411), .A3(n4437), .ZN(n4436) );
  NOR2_X1 U3081 ( .A1(n4438), .A2(n4411), .ZN(n4433) );
  XOR2_X1 U3082 ( .A(n4408), .B(n4439), .Z(n4421) );
  XNOR2_X1 U3083 ( .A(n4409), .B(n4392), .ZN(n4439) );
  XNOR2_X1 U3084 ( .A(n4440), .B(n4441), .ZN(n4392) );
  NAND2_X1 U3085 ( .A1(n4442), .A2(n4443), .ZN(n4440) );
  NAND2_X1 U3086 ( .A1(n4444), .A2(n4445), .ZN(n4443) );
  INV_X1 U3087 ( .A(n4446), .ZN(n4445) );
  XOR2_X1 U3088 ( .A(n4447), .B(n4448), .Z(n4444) );
  XOR2_X1 U3089 ( .A(n4449), .B(n4450), .Z(n4448) );
  XOR2_X1 U3090 ( .A(n4451), .B(n4452), .Z(n4447) );
  NOR2_X1 U3091 ( .A1(n4453), .A2(n4454), .ZN(n4452) );
  NAND2_X1 U3092 ( .A1(n4455), .A2(n4446), .ZN(n4442) );
  NOR4_X1 U3093 ( .A1(n4456), .A2(n4457), .A3(KEYINPUT115), .A4(KEYINPUT61),  .ZN(n4446) );
  AND2_X1 U3094 ( .A1(n4458), .A2(n4389), .ZN(n4457) );
  INV_X1 U3095 ( .A(n4419), .ZN(n4389) );
  OR3_X1 U3096 ( .A1(n4459), .A2(KEYINPUT88), .A3(n4460), .ZN(n4458) );
  INV_X1 U3097 ( .A(KEYINPUT87), .ZN(n4460) );
  XOR2_X1 U3098 ( .A(n4461), .B(n4462), .Z(n4455) );
  XNOR2_X1 U3099 ( .A(n4463), .B(n4451), .ZN(n4462) );
  XNOR2_X1 U3100 ( .A(n4464), .B(n4465), .ZN(n4451) );
  NAND2_X1 U3101 ( .A1(n4466), .A2(n4467), .ZN(n4464) );
  NAND2_X1 U3102 ( .A1(n4468), .A2(n4469), .ZN(n4467) );
  NAND2_X1 U3103 ( .A1(n4470), .A2(n4471), .ZN(n4469) );
  OR2_X1 U3104 ( .A1(n4472), .A2(n4473), .ZN(n4471) );
  NAND2_X1 U3105 ( .A1(n4474), .A2(n4475), .ZN(n4466) );
  XOR2_X1 U3106 ( .A(n4473), .B(n4472), .Z(n4474) );
  XNOR2_X1 U3107 ( .A(n4454), .B(n4476), .ZN(n4461) );
  XNOR2_X1 U3108 ( .A(n4412), .B(n4400), .ZN(n4408) );
  NOR2_X1 U3109 ( .A1(n4477), .A2(n4478), .ZN(n4412) );
  AND2_X1 U3110 ( .A1(n4479), .A2(n4437), .ZN(n4477) );
  NOR3_X1 U3111 ( .A1(KEYINPUT26), .A2(KEYINPUT18), .A3(n4480), .ZN(n4419) );
  XNOR2_X1 U3112 ( .A(n4431), .B(n4481), .ZN(G319) );
  NOR2_X1 U3113 ( .A1(n4482), .A2(n4432), .ZN(n4481) );
  NOR2_X1 U3114 ( .A1(n4483), .A2(n4479), .ZN(n4482) );
  XNOR2_X1 U3115 ( .A(n4484), .B(n4411), .ZN(G316) );
  XNOR2_X1 U3116 ( .A(n4410), .B(n4485), .ZN(G313) );
  NOR4_X1 U3117 ( .A1(KEYINPUT166), .A2(KEYINPUT135), .A3(n4397), .A4(n4486),  .ZN(n4485) );
  NOR2_X1 U3118 ( .A1(n4411), .A2(n4487), .ZN(n4486) );
  XNOR2_X1 U3119 ( .A(n4488), .B(n4489), .ZN(G310) );
  NAND3_X1 U3120 ( .A1(n4427), .A2(n4490), .A3(n4491), .ZN(n4488) );
  NOR3_X1 U3121 ( .A1(KEYINPUT105), .A2(KEYINPUT79), .A3(KEYINPUT175), .ZN(n4491) );
  NAND2_X1 U3122 ( .A1(n4484), .A2(n4413), .ZN(n4490) );
  INV_X1 U3123 ( .A(n4487), .ZN(n4484) );
  NAND2_X1 U3124 ( .A1(n4492), .A2(n4396), .ZN(n4487) );
  INV_X1 U3125 ( .A(n4398), .ZN(n4396) );
  NOR2_X1 U3126 ( .A1(n4493), .A2(n4478), .ZN(n4398) );
  NAND2_X1 U3127 ( .A1(n4483), .A2(n4425), .ZN(n4492) );
  INV_X1 U3128 ( .A(n4493), .ZN(n4425) );
  XNOR2_X1 U3129 ( .A(n4472), .B(n4494), .ZN(G307) );
  XNOR2_X1 U3130 ( .A(n4495), .B(n4473), .ZN(G304) );
  NAND2_X1 U3131 ( .A1(n4496), .A2(n4450), .ZN(n4495) );
  NAND2_X1 U3132 ( .A1(n4011), .A2(G2239), .ZN(n4450) );
  NAND2_X1 U3133 ( .A1(n4494), .A2(n4476), .ZN(n4496) );
  INV_X1 U3134 ( .A(n4497), .ZN(n4476) );
  XNOR2_X1 U3135 ( .A(n4498), .B(n4499), .ZN(G301) );
  NOR2_X1 U3136 ( .A1(n4500), .A2(n4454), .ZN(n4499) );
  NOR2_X1 U3137 ( .A1(n4494), .A2(n4470), .ZN(n4500) );
  XNOR2_X1 U3138 ( .A(n4501), .B(n4468), .ZN(G298) );
  NAND2_X1 U3139 ( .A1(n4449), .A2(n4502), .ZN(n4501) );
  NAND2_X1 U3140 ( .A1(n4494), .A2(n4463), .ZN(n4502) );
  NOR3_X1 U3141 ( .A1(KEYINPUT53), .A2(n4503), .A3(n4504), .ZN(n4494) );
  NOR2_X1 U3142 ( .A1(n4483), .A2(n4505), .ZN(n4503) );
  NAND2_X1 U3143 ( .A1(n4463), .A2(n4506), .ZN(n4449) );
  NAND2_X1 U3144 ( .A1(n4453), .A2(n4498), .ZN(n4506) );
  INV_X1 U3145 ( .A(n4470), .ZN(n4453) );
  INV_X1 U3146 ( .A(n4507), .ZN(n4463) );
  XOR2_X1 U3147 ( .A(n4479), .B(n4483), .Z(G295) );
  NOR3_X1 U3148 ( .A1(KEYINPUT27), .A2(KEYINPUT19), .A3(n4508), .ZN(n4483) );
  NAND3_X1 U3149 ( .A1(G133), .A2(n4509), .A3(G134), .ZN(G292) );
  NAND2_X1 U3150 ( .A1(G1197), .A2(n4509), .ZN(G289) );
  INV_X1 U3151 ( .A(G5), .ZN(n4509) );
  AND2_X1 U3152 ( .A1(G1), .A2(G163), .ZN(G278) );
  NAND2_X1 U3153 ( .A1(n4510), .A2(n4511), .ZN(G276) );
  NAND2_X1 U3154 ( .A1(n4512), .A2(n4513), .ZN(n4511) );
  NAND2_X1 U3155 ( .A1(KEYINPUT56), .A2(n4362), .ZN(n4513) );
  AND2_X1 U3156 ( .A1(n4514), .A2(n4515), .ZN(n4362) );
  NAND2_X1 U3157 ( .A1(n4516), .A2(n4321), .ZN(n4515) );
  INV_X1 U3158 ( .A(n4336), .ZN(n4321) );
  NOR4_X1 U3159 ( .A1(KEYINPUT16), .A2(n4517), .A3(KEYINPUT7), .A4(KEYINPUT28),  .ZN(n4336) );
  NAND2_X1 U3160 ( .A1(n4510), .A2(n4518), .ZN(G273) );
  NAND2_X1 U3161 ( .A1(n4512), .A2(n3806), .ZN(n4518) );
  NAND3_X1 U3162 ( .A1(n4519), .A2(n4520), .A3(n4521), .ZN(n3806) );
  NOR3_X1 U3163 ( .A1(KEYINPUT126), .A2(KEYINPUT64), .A3(KEYINPUT55), .ZN(n4521) );
  NAND2_X1 U3164 ( .A1(n4371), .A2(n4522), .ZN(n4520) );
  INV_X1 U3165 ( .A(n4382), .ZN(n4371) );
  NOR4_X1 U3166 ( .A1(KEYINPUT17), .A2(n4523), .A3(KEYINPUT8), .A4(KEYINPUT29),  .ZN(n4382) );
  INV_X1 U3167 ( .A(n4524), .ZN(n4519) );
  NAND4_X1 U3168 ( .A1(n4525), .A2(n4510), .A3(n4526), .A4(n4527), .ZN(G270) );
  NOR4_X1 U3169 ( .A1(KEYINPUT5), .A2(KEYINPUT42), .A3(KEYINPUT23), .A4(KEYINPUT12), .ZN(n4527) );
  NAND2_X1 U3170 ( .A1(KEYINPUT45), .A2(n4517), .ZN(n4526) );
  NAND2_X1 U3171 ( .A1(n4512), .A2(n4528), .ZN(n4525) );
  NAND2_X1 U3172 ( .A1(n4514), .A2(n4529), .ZN(n4528) );
  NAND2_X1 U3173 ( .A1(n4516), .A2(n4517), .ZN(n4529) );
  NAND3_X1 U3174 ( .A1(n4530), .A2(n4531), .A3(n4532), .ZN(n4517) );
  NOR3_X1 U3175 ( .A1(n4533), .A2(KEYINPUT81), .A3(KEYINPUT128), .ZN(n4532) );
  NOR2_X1 U3176 ( .A1(n4534), .A2(n4535), .ZN(n4533) );
  NOR3_X1 U3177 ( .A1(n4456), .A2(KEYINPUT61), .A3(KEYINPUT115), .ZN(n4534) );
  NAND2_X1 U3178 ( .A1(n4480), .A2(n4536), .ZN(n4531) );
  OR2_X1 U3179 ( .A1(KEYINPUT32), .A2(n4537), .ZN(n4536) );
  NOR2_X1 U3180 ( .A1(n4535), .A2(n4538), .ZN(n4537) );
  NOR2_X1 U3181 ( .A1(KEYINPUT88), .A2(n4459), .ZN(n4538) );
  NOR2_X1 U3182 ( .A1(KEYINPUT158), .A2(n4539), .ZN(n4535) );
  NAND3_X1 U3183 ( .A1(n4540), .A2(n4541), .A3(n4542), .ZN(n4480) );
  NOR3_X1 U3184 ( .A1(n4543), .A2(KEYINPUT78), .A3(KEYINPUT111), .ZN(n4542) );
  NOR2_X1 U3185 ( .A1(n4544), .A2(n4545), .ZN(n4543) );
  NOR3_X1 U3186 ( .A1(n4252), .A2(KEYINPUT60), .A3(KEYINPUT112), .ZN(n4544) );
  NAND2_X1 U3187 ( .A1(n4546), .A2(n4547), .ZN(n4541) );
  OR2_X1 U3188 ( .A1(KEYINPUT35), .A2(n4548), .ZN(n4547) );
  NOR2_X1 U3189 ( .A1(n4549), .A2(n4545), .ZN(n4548) );
  NOR2_X1 U3190 ( .A1(KEYINPUT153), .A2(n4550), .ZN(n4545) );
  NOR2_X1 U3191 ( .A1(KEYINPUT92), .A2(n4262), .ZN(n4549) );
  NAND4_X1 U3192 ( .A1(n4551), .A2(n4552), .A3(n4553), .A4(n4554), .ZN(n4546) );
  NOR3_X1 U3193 ( .A1(KEYINPUT106), .A2(KEYINPUT76), .A3(KEYINPUT177), .ZN(n4554) );
  NAND2_X1 U3194 ( .A1(n4555), .A2(n4145), .ZN(n4552) );
  NAND3_X1 U3195 ( .A1(n4556), .A2(n4557), .A3(n4558), .ZN(n4145) );
  NOR3_X1 U3196 ( .A1(KEYINPUT107), .A2(KEYINPUT51), .A3(KEYINPUT180), .ZN(n4558) );
  NAND2_X1 U3197 ( .A1(G4526), .A2(n4559), .ZN(n4557) );
  OR2_X1 U3198 ( .A1(n4560), .A2(KEYINPUT122), .ZN(n4559) );
  INV_X1 U3199 ( .A(n4561), .ZN(n4556) );
  NAND2_X1 U3200 ( .A1(n4260), .A2(n4259), .ZN(n4555) );
  INV_X1 U3201 ( .A(KEYINPUT151), .ZN(n4260) );
  NAND2_X1 U3202 ( .A1(KEYINPUT38), .A2(G4526), .ZN(n4551) );
  NAND2_X1 U3203 ( .A1(n4562), .A2(n4563), .ZN(n4516) );
  INV_X1 U3204 ( .A(KEYINPUT94), .ZN(n4563) );
  NOR3_X1 U3205 ( .A1(KEYINPUT63), .A2(KEYINPUT123), .A3(n4524), .ZN(n4514) );
  OR3_X1 U3206 ( .A1(KEYINPUT10), .A2(n4564), .A3(n4565), .ZN(G264) );
  OR3_X1 U3207 ( .A1(KEYINPUT40), .A2(KEYINPUT3), .A3(KEYINPUT21), .ZN(n4565) );
  OR3_X1 U3208 ( .A1(KEYINPUT2), .A2(n4564), .A3(n4566), .ZN(G258) );
  OR3_X1 U3209 ( .A1(KEYINPUT9), .A2(KEYINPUT39), .A3(KEYINPUT20), .ZN(n4566) );
  NAND2_X1 U3210 ( .A1(n4567), .A2(n4568), .ZN(n4564) );
  NAND2_X1 U3211 ( .A1(KEYINPUT47), .A2(n4569), .ZN(n4568) );
  NAND2_X1 U3212 ( .A1(n4570), .A2(n4571), .ZN(G252) );
  NAND2_X1 U3213 ( .A1(n4572), .A2(n4573), .ZN(n4571) );
  NAND3_X1 U3214 ( .A1(n4574), .A2(n4575), .A3(KEYINPUT49), .ZN(n4573) );
  NAND2_X1 U3215 ( .A1(n4576), .A2(n4577), .ZN(n4575) );
  NAND2_X1 U3216 ( .A1(n4578), .A2(n4579), .ZN(n4577) );
  NAND2_X1 U3217 ( .A1(n4580), .A2(n4581), .ZN(n4579) );
  NAND2_X1 U3218 ( .A1(KEYINPUT65), .A2(n4582), .ZN(n4581) );
  NAND2_X1 U3219 ( .A1(KEYINPUT147), .A2(n4583), .ZN(n4580) );
  INV_X1 U3220 ( .A(n4584), .ZN(n4576) );
  NAND2_X1 U3221 ( .A1(KEYINPUT146), .A2(n4585), .ZN(n4572) );
  NAND2_X1 U3222 ( .A1(n4567), .A2(n4586), .ZN(G249) );
  NAND2_X1 U3223 ( .A1(n4587), .A2(n4588), .ZN(n4586) );
  NAND2_X1 U3224 ( .A1(KEYINPUT54), .A2(n4589), .ZN(n4587) );
  NAND2_X1 U3225 ( .A1(n4590), .A2(n4591), .ZN(n4589) );
  OR3_X1 U3226 ( .A1(KEYINPUT6), .A2(KEYINPUT25), .A3(KEYINPUT15), .ZN(n4591) );
  AND2_X1 U3227 ( .A1(n4592), .A2(n4593), .ZN(n4567) );
  NAND2_X1 U3228 ( .A1(G38), .A2(n4594), .ZN(n4593) );
  OR3_X1 U3229 ( .A1(G1455), .A2(G2204), .A3(n4595), .ZN(n4594) );
  INV_X1 U3230 ( .A(G4528), .ZN(n4595) );
  NAND2_X1 U3231 ( .A1(n4588), .A2(n4596), .ZN(n4592) );
  NAND4_X1 U3232 ( .A1(n4597), .A2(n4598), .A3(n4599), .A4(n4600), .ZN(n4596) );
  NAND2_X1 U3233 ( .A1(n4590), .A2(n4569), .ZN(n4600) );
  NAND4_X1 U3234 ( .A1(n4601), .A2(n4602), .A3(n4603), .A4(n4604), .ZN(n4569) );
  NOR3_X1 U3235 ( .A1(n4605), .A2(KEYINPUT80), .A3(KEYINPUT117), .ZN(n4604) );
  NOR2_X1 U3236 ( .A1(n4606), .A2(n4607), .ZN(n4605) );
  NOR2_X1 U3237 ( .A1(n4608), .A2(KEYINPUT148), .ZN(n4607) );
  NOR4_X1 U3238 ( .A1(n4609), .A2(n4610), .A3(n4611), .A4(n4612), .ZN(n4608) );
  NOR2_X1 U3239 ( .A1(n3934), .A2(n3875), .ZN(n4612) );
  NOR4_X1 U3240 ( .A1(n4613), .A2(KEYINPUT100), .A3(KEYINPUT58), .A4(KEYINPUT165), .ZN(n4606) );
  NAND3_X1 U3241 ( .A1(n4614), .A2(n4615), .A3(n4616), .ZN(n4613) );
  NAND2_X1 U3242 ( .A1(KEYINPUT84), .A2(n4617), .ZN(n4616) );
  NAND3_X1 U3243 ( .A1(n4618), .A2(n4619), .A3(n4620), .ZN(n4615) );
  OR2_X1 U3244 ( .A1(n3891), .A2(n3935), .ZN(n4620) );
  NAND3_X1 U3245 ( .A1(n4621), .A2(n4622), .A3(n4623), .ZN(n4619) );
  NAND2_X1 U3246 ( .A1(n3889), .A2(n3937), .ZN(n4623) );
  NAND3_X1 U3247 ( .A1(n4624), .A2(n4625), .A3(n4626), .ZN(n4622) );
  OR2_X1 U3248 ( .A1(n3882), .A2(n3924), .ZN(n4626) );
  NAND3_X1 U3249 ( .A1(n4627), .A2(n4628), .A3(n4629), .ZN(n4625) );
  NAND2_X1 U3250 ( .A1(n3880), .A2(n3931), .ZN(n4629) );
  NAND2_X1 U3251 ( .A1(n4630), .A2(n4617), .ZN(n4628) );
  OR2_X1 U3252 ( .A1(n3881), .A2(n3930), .ZN(n4630) );
  NAND2_X1 U3253 ( .A1(n3881), .A2(n3930), .ZN(n4627) );
  NAND2_X1 U3254 ( .A1(n4631), .A2(n4632), .ZN(n3930) );
  OR2_X1 U3255 ( .A1(n3844), .A2(G2211), .ZN(n4632) );
  NAND2_X1 U3256 ( .A1(G65), .A2(n3844), .ZN(n4631) );
  NAND2_X1 U3257 ( .A1(n4633), .A2(n4634), .ZN(n3881) );
  NAND2_X1 U3258 ( .A1(G147), .A2(n3844), .ZN(n4634) );
  NAND2_X1 U3259 ( .A1(G171), .A2(G18), .ZN(n4633) );
  OR2_X1 U3260 ( .A1(n3880), .A2(n3931), .ZN(n4624) );
  NAND2_X1 U3261 ( .A1(n4635), .A2(n4636), .ZN(n3931) );
  OR2_X1 U3262 ( .A1(n3844), .A2(G2218), .ZN(n4636) );
  NAND2_X1 U3263 ( .A1(G83), .A2(n3844), .ZN(n4635) );
  NAND2_X1 U3264 ( .A1(n4637), .A2(n4638), .ZN(n3880) );
  NAND2_X1 U3265 ( .A1(G180), .A2(G18), .ZN(n4637) );
  NAND2_X1 U3266 ( .A1(n3882), .A2(n3924), .ZN(n4621) );
  NAND2_X1 U3267 ( .A1(n4639), .A2(n4640), .ZN(n3924) );
  OR2_X1 U3268 ( .A1(n3844), .A2(G2224), .ZN(n4640) );
  NAND2_X1 U3269 ( .A1(G84), .A2(n3844), .ZN(n4639) );
  NAND2_X1 U3270 ( .A1(n4641), .A2(n4642), .ZN(n3882) );
  NAND2_X1 U3271 ( .A1(G179), .A2(G18), .ZN(n4641) );
  OR2_X1 U3272 ( .A1(n3889), .A2(n3937), .ZN(n4618) );
  NAND2_X1 U3273 ( .A1(n4643), .A2(n4644), .ZN(n3937) );
  NAND2_X1 U3274 ( .A1(G18), .A2(n4645), .ZN(n4644) );
  NAND2_X1 U3275 ( .A1(G85), .A2(n3844), .ZN(n4643) );
  NAND2_X1 U3276 ( .A1(n4646), .A2(n4647), .ZN(n3889) );
  NAND2_X1 U3277 ( .A1(G178), .A2(G18), .ZN(n4646) );
  NAND2_X1 U3278 ( .A1(n3935), .A2(n3891), .ZN(n4614) );
  NAND2_X1 U3279 ( .A1(n4648), .A2(n4649), .ZN(n3891) );
  NAND2_X1 U3280 ( .A1(G177), .A2(n3860), .ZN(n4649) );
  NAND2_X1 U3281 ( .A1(n4650), .A2(n4651), .ZN(n3935) );
  NAND2_X1 U3282 ( .A1(G18), .A2(n4652), .ZN(n4651) );
  NAND2_X1 U3283 ( .A1(G64), .A2(n3844), .ZN(n4650) );
  NAND2_X1 U3284 ( .A1(n3922), .A2(n3874), .ZN(n4603) );
  NAND2_X1 U3285 ( .A1(n4653), .A2(n4654), .ZN(n4602) );
  INV_X1 U3286 ( .A(n4610), .ZN(n4654) );
  NOR2_X1 U3287 ( .A1(n3874), .A2(n3922), .ZN(n4610) );
  NAND2_X1 U3288 ( .A1(n4655), .A2(n4656), .ZN(n3922) );
  NAND2_X1 U3289 ( .A1(G18), .A2(n4657), .ZN(n4656) );
  NAND2_X1 U3290 ( .A1(G110), .A2(n3844), .ZN(n4655) );
  NAND2_X1 U3291 ( .A1(n4648), .A2(n4658), .ZN(n3874) );
  NAND2_X1 U3292 ( .A1(G173), .A2(n3860), .ZN(n4658) );
  NAND2_X1 U3293 ( .A1(n4659), .A2(n4660), .ZN(n4653) );
  NAND2_X1 U3294 ( .A1(n4661), .A2(n4662), .ZN(n4660) );
  INV_X1 U3295 ( .A(n4609), .ZN(n4662) );
  NOR2_X1 U3296 ( .A1(n3890), .A2(n3936), .ZN(n4609) );
  NAND2_X1 U3297 ( .A1(n4663), .A2(n4664), .ZN(n4661) );
  NAND3_X1 U3298 ( .A1(n4665), .A2(n3875), .A3(n3934), .ZN(n4664) );
  NAND2_X1 U3299 ( .A1(n4666), .A2(n4667), .ZN(n3934) );
  OR2_X1 U3300 ( .A1(n3844), .A2(G2239), .ZN(n4667) );
  NAND2_X1 U3301 ( .A1(G63), .A2(n3844), .ZN(n4666) );
  NAND2_X1 U3302 ( .A1(n4648), .A2(n4668), .ZN(n3875) );
  NAND2_X1 U3303 ( .A1(G176), .A2(n3860), .ZN(n4668) );
  INV_X1 U3304 ( .A(n4611), .ZN(n4665) );
  NOR2_X1 U3305 ( .A1(n3888), .A2(n3921), .ZN(n4611) );
  NAND2_X1 U3306 ( .A1(n3921), .A2(n3888), .ZN(n4663) );
  NAND2_X1 U3307 ( .A1(n4648), .A2(n4669), .ZN(n3888) );
  NAND2_X1 U3308 ( .A1(G175), .A2(n3860), .ZN(n4669) );
  NAND2_X1 U3309 ( .A1(n4670), .A2(n4671), .ZN(n3921) );
  NAND2_X1 U3310 ( .A1(G18), .A2(n4672), .ZN(n4671) );
  NAND2_X1 U3311 ( .A1(G86), .A2(n3844), .ZN(n4670) );
  NAND2_X1 U3312 ( .A1(n3936), .A2(n3890), .ZN(n4659) );
  NAND2_X1 U3313 ( .A1(n4648), .A2(n4673), .ZN(n3890) );
  NAND2_X1 U3314 ( .A1(G174), .A2(n3860), .ZN(n4673) );
  NAND2_X1 U3315 ( .A1(n4674), .A2(n4675), .ZN(n3936) );
  NAND2_X1 U3316 ( .A1(G18), .A2(n4676), .ZN(n4675) );
  NAND2_X1 U3317 ( .A1(G109), .A2(n3844), .ZN(n4674) );
  NAND2_X1 U3318 ( .A1(KEYINPUT31), .A2(n4617), .ZN(n4601) );
  OR4_X1 U3319 ( .A1(n4677), .A2(n4678), .A3(KEYINPUT69), .A4(n4679), .ZN(n4617) );
  NOR2_X1 U3320 ( .A1(n4680), .A2(n4681), .ZN(n4679) );
  NOR2_X1 U3321 ( .A1(n4682), .A2(KEYINPUT30), .ZN(n4681) );
  NOR2_X1 U3322 ( .A1(n4585), .A2(n4584), .ZN(n4682) );
  NOR2_X1 U3323 ( .A1(KEYINPUT83), .A2(n4683), .ZN(n4584) );
  NOR3_X1 U3324 ( .A1(n4684), .A2(n4685), .A3(n4686), .ZN(n4683) );
  NOR2_X1 U3325 ( .A1(n3979), .A2(n3904), .ZN(n4685) );
  NOR4_X1 U3326 ( .A1(KEYINPUT68), .A2(n4687), .A3(n4688), .A4(n4689), .ZN(n4680) );
  INV_X1 U3327 ( .A(n4578), .ZN(n4689) );
  NOR4_X1 U3328 ( .A1(n4690), .A2(n4691), .A3(KEYINPUT98), .A4(KEYINPUT162),  .ZN(n4578) );
  NOR2_X1 U3329 ( .A1(n4692), .A2(n4693), .ZN(n4691) );
  NOR2_X1 U3330 ( .A1(n4694), .A2(n4695), .ZN(n4692) );
  NOR2_X1 U3331 ( .A1(n4696), .A2(n4697), .ZN(n4695) );
  NOR2_X1 U3332 ( .A1(n4698), .A2(n4699), .ZN(n4696) );
  AND3_X1 U3333 ( .A1(n3846), .A2(n4700), .A3(n3945), .ZN(n4699) );
  NAND2_X1 U3334 ( .A1(n3957), .A2(n3835), .ZN(n4700) );
  NOR2_X1 U3335 ( .A1(n3957), .A2(n3835), .ZN(n4698) );
  NOR2_X1 U3336 ( .A1(n4701), .A2(n3850), .ZN(n4694) );
  NOR2_X1 U3337 ( .A1(n3958), .A2(n4702), .ZN(n4690) );
  AND2_X1 U3338 ( .A1(KEYINPUT36), .A2(G89), .ZN(n4688) );
  NOR2_X1 U3339 ( .A1(n4583), .A2(n4582), .ZN(n4687) );
  AND4_X1 U3340 ( .A1(n4703), .A2(n4704), .A3(n4705), .A4(n4706), .ZN(n4582) );
  NOR3_X1 U3341 ( .A1(KEYINPUT163), .A2(KEYINPUT99), .A3(KEYINPUT48), .ZN(n4706) );
  NAND2_X1 U3342 ( .A1(n3832), .A2(n3942), .ZN(n4705) );
  NAND2_X1 U3343 ( .A1(G89), .A2(n4707), .ZN(n4704) );
  OR2_X1 U3344 ( .A1(KEYINPUT119), .A2(n4708), .ZN(n4707) );
  NOR4_X1 U3345 ( .A1(n4709), .A2(n4710), .A3(n4711), .A4(n4712), .ZN(n4708) );
  NOR2_X1 U3346 ( .A1(n3942), .A2(n3832), .ZN(n4711) );
  NOR3_X1 U3347 ( .A1(n3840), .A2(G70), .A3(G18), .ZN(n4710) );
  NAND2_X1 U3348 ( .A1(n4713), .A2(n4714), .ZN(n4703) );
  NAND2_X1 U3349 ( .A1(n4715), .A2(n4716), .ZN(n4714) );
  NAND2_X1 U3350 ( .A1(n4717), .A2(n4718), .ZN(n4716) );
  NAND3_X1 U3351 ( .A1(n4719), .A2(n4720), .A3(n4721), .ZN(n4718) );
  NAND2_X1 U3352 ( .A1(n3852), .A2(n3953), .ZN(n4721) );
  NAND4_X1 U3353 ( .A1(G70), .A2(n3840), .A3(n4722), .A4(n3844), .ZN(n4720) );
  INV_X1 U3354 ( .A(n4709), .ZN(n4722) );
  NOR2_X1 U3355 ( .A1(n3852), .A2(n3953), .ZN(n4709) );
  NAND2_X1 U3356 ( .A1(n4723), .A2(n4724), .ZN(n3953) );
  OR2_X1 U3357 ( .A1(n3844), .A2(G3705), .ZN(n4724) );
  NAND2_X1 U3358 ( .A1(G74), .A2(n3844), .ZN(n4723) );
  NAND2_X1 U3359 ( .A1(n4725), .A2(n4726), .ZN(n3852) );
  NAND2_X1 U3360 ( .A1(G207), .A2(G18), .ZN(n4725) );
  NAND2_X1 U3361 ( .A1(n4727), .A2(n4728), .ZN(n3840) );
  NAND2_X1 U3362 ( .A1(G41), .A2(n3844), .ZN(n4728) );
  NAND2_X1 U3363 ( .A1(G198), .A2(G18), .ZN(n4727) );
  NAND2_X1 U3364 ( .A1(n3851), .A2(n3948), .ZN(n4719) );
  INV_X1 U3365 ( .A(n4712), .ZN(n4717) );
  NAND2_X1 U3366 ( .A1(n4729), .A2(n4730), .ZN(n4712) );
  OR2_X1 U3367 ( .A1(n3851), .A2(n3948), .ZN(n4730) );
  NAND2_X1 U3368 ( .A1(n4731), .A2(n4732), .ZN(n3948) );
  OR2_X1 U3369 ( .A1(n3844), .A2(G3711), .ZN(n4732) );
  NAND2_X1 U3370 ( .A1(G76), .A2(n3844), .ZN(n4731) );
  NAND2_X1 U3371 ( .A1(n4733), .A2(n4734), .ZN(n3851) );
  NAND2_X1 U3372 ( .A1(G26), .A2(n3844), .ZN(n4734) );
  NAND2_X1 U3373 ( .A1(G206), .A2(G18), .ZN(n4733) );
  OR2_X1 U3374 ( .A1(n3845), .A2(n3943), .ZN(n4729) );
  NAND2_X1 U3375 ( .A1(n3845), .A2(n3943), .ZN(n4715) );
  NAND2_X1 U3376 ( .A1(n4735), .A2(n4736), .ZN(n3943) );
  NAND2_X1 U3377 ( .A1(G18), .A2(n4737), .ZN(n4736) );
  NAND2_X1 U3378 ( .A1(G75), .A2(n3844), .ZN(n4735) );
  NAND2_X1 U3379 ( .A1(n4738), .A2(n4739), .ZN(n3845) );
  NAND2_X1 U3380 ( .A1(G205), .A2(G18), .ZN(n4738) );
  OR2_X1 U3381 ( .A1(n3832), .A2(n3942), .ZN(n4713) );
  NAND2_X1 U3382 ( .A1(n4740), .A2(n4741), .ZN(n3942) );
  NAND2_X1 U3383 ( .A1(G18), .A2(n4742), .ZN(n4741) );
  NAND2_X1 U3384 ( .A1(G73), .A2(n3844), .ZN(n4740) );
  NAND2_X1 U3385 ( .A1(n4743), .A2(n4744), .ZN(n3832) );
  NAND2_X1 U3386 ( .A1(G204), .A2(G18), .ZN(n4743) );
  NOR2_X1 U3387 ( .A1(KEYINPUT145), .A2(n4745), .ZN(n4583) );
  NOR4_X1 U3388 ( .A1(n4746), .A2(n4747), .A3(n4697), .A4(n4693), .ZN(n4745) );
  NOR2_X1 U3389 ( .A1(n4748), .A2(n3849), .ZN(n4693) );
  INV_X1 U3390 ( .A(n4702), .ZN(n3849) );
  NAND2_X1 U3391 ( .A1(n4749), .A2(n4750), .ZN(n4702) );
  OR2_X1 U3392 ( .A1(G200), .A2(n3844), .ZN(n4750) );
  INV_X1 U3393 ( .A(n3958), .ZN(n4748) );
  NAND2_X1 U3394 ( .A1(n4751), .A2(n4752), .ZN(n3958) );
  NAND2_X1 U3395 ( .A1(G3749), .A2(G18), .ZN(n4752) );
  OR2_X1 U3396 ( .A1(G56), .A2(G18), .ZN(n4751) );
  NOR2_X1 U3397 ( .A1(n3944), .A2(n4753), .ZN(n4697) );
  INV_X1 U3398 ( .A(n3850), .ZN(n4753) );
  NAND2_X1 U3399 ( .A1(n4754), .A2(n4755), .ZN(n3850) );
  OR2_X1 U3400 ( .A1(G201), .A2(n3844), .ZN(n4755) );
  INV_X1 U3401 ( .A(n4701), .ZN(n3944) );
  NAND2_X1 U3402 ( .A1(n4756), .A2(n4757), .ZN(n4701) );
  NAND2_X1 U3403 ( .A1(G3743), .A2(G18), .ZN(n4757) );
  OR2_X1 U3404 ( .A1(G55), .A2(G18), .ZN(n4756) );
  AND2_X1 U3405 ( .A1(n3957), .A2(n3835), .ZN(n4747) );
  NAND2_X1 U3406 ( .A1(n4758), .A2(n4759), .ZN(n3835) );
  OR2_X1 U3407 ( .A1(G202), .A2(n3844), .ZN(n4759) );
  OR2_X1 U3408 ( .A1(G127), .A2(G18), .ZN(n4758) );
  NAND2_X1 U3409 ( .A1(n4760), .A2(n4761), .ZN(n3957) );
  NAND2_X1 U3410 ( .A1(G3737), .A2(G18), .ZN(n4761) );
  OR2_X1 U3411 ( .A1(G54), .A2(G18), .ZN(n4760) );
  NOR2_X1 U3412 ( .A1(n3945), .A2(n3846), .ZN(n4746) );
  NAND2_X1 U3413 ( .A1(n4762), .A2(n4763), .ZN(n3846) );
  NAND2_X1 U3414 ( .A1(G130), .A2(n3844), .ZN(n4763) );
  NAND2_X1 U3415 ( .A1(G203), .A2(G18), .ZN(n4762) );
  NAND2_X1 U3416 ( .A1(n4764), .A2(n4765), .ZN(n3945) );
  OR2_X1 U3417 ( .A1(n3844), .A2(G3729), .ZN(n4765) );
  NAND2_X1 U3418 ( .A1(G53), .A2(n3844), .ZN(n4764) );
  INV_X1 U3419 ( .A(n4570), .ZN(n4678) );
  NOR4_X1 U3420 ( .A1(n4766), .A2(n4767), .A3(KEYINPUT96), .A4(KEYINPUT160),  .ZN(n4570) );
  AND2_X1 U3421 ( .A1(n4768), .A2(n4769), .ZN(n4767) );
  NOR2_X1 U3422 ( .A1(n4770), .A2(n3969), .ZN(n4766) );
  NOR2_X1 U3423 ( .A1(n4769), .A2(n4768), .ZN(n4770) );
  NAND2_X1 U3424 ( .A1(n4771), .A2(n4772), .ZN(n4768) );
  NAND2_X1 U3425 ( .A1(n4773), .A2(n3965), .ZN(n4772) );
  NAND2_X1 U3426 ( .A1(n4774), .A2(n4775), .ZN(n4771) );
  NAND2_X1 U3427 ( .A1(n4776), .A2(n4777), .ZN(n4775) );
  NAND2_X1 U3428 ( .A1(n3908), .A2(n3970), .ZN(n4777) );
  NAND3_X1 U3429 ( .A1(n3966), .A2(n4778), .A3(n3900), .ZN(n4776) );
  NAND2_X1 U3430 ( .A1(n4779), .A2(n4780), .ZN(n4778) );
  NAND2_X1 U3431 ( .A1(n3910), .A2(n4781), .ZN(n4774) );
  INV_X1 U3432 ( .A(n3893), .ZN(n4769) );
  NOR2_X1 U3433 ( .A1(n4585), .A2(n4574), .ZN(n4677) );
  AND3_X1 U3434 ( .A1(n4782), .A2(n4783), .A3(n4784), .ZN(n4574) );
  NOR3_X1 U3435 ( .A1(KEYINPUT161), .A2(KEYINPUT97), .A3(KEYINPUT57), .ZN(n4784) );
  NAND2_X1 U3436 ( .A1(n4785), .A2(n4786), .ZN(n4783) );
  NAND3_X1 U3437 ( .A1(n4787), .A2(n4788), .A3(n4789), .ZN(n4786) );
  NAND2_X1 U3438 ( .A1(n3895), .A2(n3964), .ZN(n4789) );
  NAND2_X1 U3439 ( .A1(n4790), .A2(n4791), .ZN(n4788) );
  NAND2_X1 U3440 ( .A1(n4792), .A2(n4793), .ZN(n4791) );
  NAND2_X1 U3441 ( .A1(n3905), .A2(n3978), .ZN(n4793) );
  NAND2_X1 U3442 ( .A1(n3904), .A2(n3979), .ZN(n4792) );
  NAND2_X1 U3443 ( .A1(n4794), .A2(n4795), .ZN(n3979) );
  OR2_X1 U3444 ( .A1(n3844), .A2(G4394), .ZN(n4795) );
  NAND2_X1 U3445 ( .A1(G77), .A2(n3844), .ZN(n4794) );
  NAND2_X1 U3446 ( .A1(n4796), .A2(n4797), .ZN(n3904) );
  NAND2_X1 U3447 ( .A1(G118), .A2(n3844), .ZN(n4797) );
  NAND2_X1 U3448 ( .A1(G187), .A2(G18), .ZN(n4796) );
  INV_X1 U3449 ( .A(n4686), .ZN(n4790) );
  NAND2_X1 U3450 ( .A1(n4798), .A2(n4799), .ZN(n4686) );
  OR2_X1 U3451 ( .A1(n3905), .A2(n3978), .ZN(n4799) );
  NAND2_X1 U3452 ( .A1(n4800), .A2(n4801), .ZN(n3978) );
  NAND2_X1 U3453 ( .A1(G18), .A2(n4802), .ZN(n4801) );
  NAND2_X1 U3454 ( .A1(G78), .A2(n3844), .ZN(n4800) );
  NAND2_X1 U3455 ( .A1(n4803), .A2(n4804), .ZN(n3905) );
  NAND2_X1 U3456 ( .A1(G196), .A2(G18), .ZN(n4803) );
  OR2_X1 U3457 ( .A1(n3909), .A2(n3972), .ZN(n4798) );
  NAND2_X1 U3458 ( .A1(n3909), .A2(n3972), .ZN(n4787) );
  NAND2_X1 U3459 ( .A1(n4805), .A2(n4806), .ZN(n3972) );
  OR2_X1 U3460 ( .A1(n3844), .A2(G4405), .ZN(n4806) );
  NAND2_X1 U3461 ( .A1(G59), .A2(n3844), .ZN(n4805) );
  NAND2_X1 U3462 ( .A1(n4807), .A2(n4808), .ZN(n3909) );
  NAND2_X1 U3463 ( .A1(G94), .A2(n3844), .ZN(n4808) );
  NAND2_X1 U3464 ( .A1(G195), .A2(G18), .ZN(n4807) );
  INV_X1 U3465 ( .A(n4684), .ZN(n4785) );
  NAND2_X1 U3466 ( .A1(n4809), .A2(n4810), .ZN(n4684) );
  OR2_X1 U3467 ( .A1(n3895), .A2(n3964), .ZN(n4810) );
  NAND2_X1 U3468 ( .A1(n4811), .A2(n4812), .ZN(n3964) );
  OR2_X1 U3469 ( .A1(n3844), .A2(G4410), .ZN(n4812) );
  NAND2_X1 U3470 ( .A1(G81), .A2(n3844), .ZN(n4811) );
  NAND2_X1 U3471 ( .A1(n4813), .A2(n4814), .ZN(n3895) );
  NAND2_X1 U3472 ( .A1(G121), .A2(n3844), .ZN(n4814) );
  NAND2_X1 U3473 ( .A1(G194), .A2(G18), .ZN(n4813) );
  OR2_X1 U3474 ( .A1(n3911), .A2(n3963), .ZN(n4809) );
  NAND2_X1 U3475 ( .A1(n3911), .A2(n3963), .ZN(n4782) );
  NAND2_X1 U3476 ( .A1(n4815), .A2(n4816), .ZN(n3963) );
  NAND2_X1 U3477 ( .A1(G18), .A2(n4817), .ZN(n4816) );
  NAND2_X1 U3478 ( .A1(G80), .A2(n3844), .ZN(n4815) );
  NAND2_X1 U3479 ( .A1(n4818), .A2(n4819), .ZN(n3911) );
  NAND2_X1 U3480 ( .A1(G193), .A2(G18), .ZN(n4818) );
  NOR2_X1 U3481 ( .A1(KEYINPUT144), .A2(n4820), .ZN(n4585) );
  NOR4_X1 U3482 ( .A1(n4821), .A2(n4822), .A3(n4823), .A4(n4824), .ZN(n4820) );
  AND2_X1 U3483 ( .A1(n3969), .A2(n3893), .ZN(n4824) );
  NAND2_X1 U3484 ( .A1(n4825), .A2(n4826), .ZN(n3893) );
  OR2_X1 U3485 ( .A1(G189), .A2(n3844), .ZN(n4826) );
  OR2_X1 U3486 ( .A1(G18), .A2(G66), .ZN(n4825) );
  NAND2_X1 U3487 ( .A1(n4827), .A2(n4828), .ZN(n3969) );
  NAND2_X1 U3488 ( .A1(G4437), .A2(G18), .ZN(n4828) );
  OR2_X1 U3489 ( .A1(G62), .A2(G18), .ZN(n4827) );
  NOR2_X1 U3490 ( .A1(n3965), .A2(n4773), .ZN(n4823) );
  INV_X1 U3491 ( .A(n3910), .ZN(n4773) );
  NAND2_X1 U3492 ( .A1(n4829), .A2(n4830), .ZN(n3910) );
  OR2_X1 U3493 ( .A1(G190), .A2(n3844), .ZN(n4830) );
  OR2_X1 U3494 ( .A1(G18), .A2(G50), .ZN(n4829) );
  INV_X1 U3495 ( .A(n4781), .ZN(n3965) );
  NAND2_X1 U3496 ( .A1(n4831), .A2(n4832), .ZN(n4781) );
  NAND2_X1 U3497 ( .A1(G4432), .A2(G18), .ZN(n4832) );
  OR2_X1 U3498 ( .A1(G61), .A2(G18), .ZN(n4831) );
  NOR2_X1 U3499 ( .A1(n3970), .A2(n3908), .ZN(n4822) );
  INV_X1 U3500 ( .A(n4779), .ZN(n3908) );
  NAND2_X1 U3501 ( .A1(n4833), .A2(n4834), .ZN(n4779) );
  OR2_X1 U3502 ( .A1(G191), .A2(n3844), .ZN(n4834) );
  OR2_X1 U3503 ( .A1(G18), .A2(G32), .ZN(n4833) );
  INV_X1 U3504 ( .A(n4780), .ZN(n3970) );
  NAND2_X1 U3505 ( .A1(n4835), .A2(n4836), .ZN(n4780) );
  NAND2_X1 U3506 ( .A1(G4427), .A2(G18), .ZN(n4836) );
  OR2_X1 U3507 ( .A1(G60), .A2(G18), .ZN(n4835) );
  NOR2_X1 U3508 ( .A1(n3966), .A2(n3900), .ZN(n4821) );
  NAND2_X1 U3509 ( .A1(n4837), .A2(n4838), .ZN(n3900) );
  NAND2_X1 U3510 ( .A1(G35), .A2(n3844), .ZN(n4838) );
  NAND2_X1 U3511 ( .A1(G192), .A2(G18), .ZN(n4837) );
  NAND2_X1 U3512 ( .A1(n4839), .A2(n4840), .ZN(n3966) );
  OR2_X1 U3513 ( .A1(n3844), .A2(G4420), .ZN(n4840) );
  NAND2_X1 U3514 ( .A1(G79), .A2(n3844), .ZN(n4839) );
  NAND2_X1 U3515 ( .A1(n4841), .A2(n4842), .ZN(n4590) );
  INV_X1 U3516 ( .A(KEYINPUT86), .ZN(n4842) );
  NAND4_X1 U3517 ( .A1(n4843), .A2(n4844), .A3(n4845), .A4(n4846), .ZN(n4841) );
  NOR2_X1 U3518 ( .A1(n4847), .A2(n4848), .ZN(n4846) );
  NOR2_X1 U3519 ( .A1(n3865), .A2(n4000), .ZN(n4848) );
  NOR2_X1 U3520 ( .A1(n4849), .A2(n3999), .ZN(n4847) );
  INV_X1 U3521 ( .A(n3871), .ZN(n4849) );
  NAND2_X1 U3522 ( .A1(n3982), .A2(n3870), .ZN(n4845) );
  NAND2_X1 U3523 ( .A1(n3992), .A2(n3857), .ZN(n4843) );
  NOR2_X1 U3524 ( .A1(KEYINPUT74), .A2(KEYINPUT118), .ZN(n4599) );
  NAND2_X1 U3525 ( .A1(n4850), .A2(n4851), .ZN(n4598) );
  NAND2_X1 U3526 ( .A1(n3857), .A2(n4852), .ZN(n4851) );
  INV_X1 U3527 ( .A(n3992), .ZN(n4850) );
  NAND2_X1 U3528 ( .A1(n4853), .A2(n4854), .ZN(n3992) );
  NAND2_X1 U3529 ( .A1(G1486), .A2(G18), .ZN(n4854) );
  OR2_X1 U3530 ( .A1(G88), .A2(G18), .ZN(n4853) );
  OR2_X1 U3531 ( .A1(n4852), .A2(n3857), .ZN(n4597) );
  NAND2_X1 U3532 ( .A1(n4855), .A2(n3860), .ZN(n3857) );
  OR2_X1 U3533 ( .A1(n3866), .A2(G166), .ZN(n4855) );
  NAND2_X1 U3534 ( .A1(n4856), .A2(n4857), .ZN(n4852) );
  NAND2_X1 U3535 ( .A1(n3982), .A2(n4858), .ZN(n4857) );
  OR2_X1 U3536 ( .A1(n4859), .A2(n3870), .ZN(n4858) );
  NAND2_X1 U3537 ( .A1(n4860), .A2(n4861), .ZN(n3982) );
  NAND2_X1 U3538 ( .A1(G18), .A2(G1480), .ZN(n4861) );
  OR2_X1 U3539 ( .A1(G18), .A2(G112), .ZN(n4860) );
  NAND2_X1 U3540 ( .A1(n4859), .A2(n3870), .ZN(n4856) );
  NAND2_X1 U3541 ( .A1(n3860), .A2(n4862), .ZN(n3870) );
  OR2_X1 U3542 ( .A1(G167), .A2(n3866), .ZN(n4862) );
  NAND2_X1 U3543 ( .A1(n4863), .A2(n4864), .ZN(n4859) );
  NAND2_X1 U3544 ( .A1(n4865), .A2(n3871), .ZN(n4864) );
  NAND2_X1 U3545 ( .A1(n3860), .A2(n4866), .ZN(n3871) );
  OR2_X1 U3546 ( .A1(G168), .A2(n3866), .ZN(n4866) );
  NAND2_X1 U3547 ( .A1(n3999), .A2(n4867), .ZN(n4865) );
  OR2_X1 U3548 ( .A1(n4867), .A2(n3999), .ZN(n4863) );
  AND2_X1 U3549 ( .A1(n4868), .A2(n4869), .ZN(n3999) );
  NAND2_X1 U3550 ( .A1(G18), .A2(G106), .ZN(n4869) );
  OR2_X1 U3551 ( .A1(G87), .A2(G18), .ZN(n4868) );
  NAND2_X1 U3552 ( .A1(n4870), .A2(n4871), .ZN(n4867) );
  NAND3_X1 U3553 ( .A1(n4000), .A2(n4844), .A3(n3865), .ZN(n4871) );
  INV_X1 U3554 ( .A(n3869), .ZN(n3865) );
  NAND2_X1 U3555 ( .A1(KEYINPUT0), .A2(n3860), .ZN(n3869) );
  NAND2_X1 U3556 ( .A1(n3858), .A2(n3987), .ZN(n4844) );
  NAND2_X1 U3557 ( .A1(n4872), .A2(n4873), .ZN(n4000) );
  OR2_X1 U3558 ( .A1(n3844), .A2(G1462), .ZN(n4873) );
  NAND2_X1 U3559 ( .A1(G113), .A2(n3844), .ZN(n4872) );
  OR2_X1 U3560 ( .A1(n3987), .A2(n3858), .ZN(n4870) );
  AND2_X1 U3561 ( .A1(n4874), .A2(n4648), .ZN(n3858) );
  NAND2_X1 U3562 ( .A1(G169), .A2(n3860), .ZN(n4874) );
  NAND2_X1 U3563 ( .A1(n4875), .A2(n4876), .ZN(n3987) );
  NAND2_X1 U3564 ( .A1(G1469), .A2(G18), .ZN(n4876) );
  OR2_X1 U3565 ( .A1(G18), .A2(G111), .ZN(n4875) );
  NAND3_X1 U3566 ( .A1(n4877), .A2(n4359), .A3(G4528), .ZN(n4588) );
  NAND2_X1 U3567 ( .A1(G1455), .A2(G2204), .ZN(n4877) );
  NAND4_X1 U3568 ( .A1(n4878), .A2(n4510), .A3(n4879), .A4(n4880), .ZN(G246) );
  NOR4_X1 U3569 ( .A1(KEYINPUT41), .A2(KEYINPUT4), .A3(KEYINPUT22), .A4(KEYINPUT11), .ZN(n4880) );
  NAND2_X1 U3570 ( .A1(KEYINPUT46), .A2(n4523), .ZN(n4879) );
  NAND2_X1 U3571 ( .A1(G38), .A2(n4881), .ZN(n4510) );
  NAND2_X1 U3572 ( .A1(G1496), .A2(n4358), .ZN(n4881) );
  NAND2_X1 U3573 ( .A1(n4512), .A2(n4882), .ZN(n4878) );
  OR4_X1 U3574 ( .A1(n4524), .A2(n4883), .A3(KEYINPUT126), .A4(KEYINPUT64),  .ZN(n4882) );
  AND2_X1 U3575 ( .A1(n4522), .A2(n4523), .ZN(n4883) );
  NAND3_X1 U3576 ( .A1(n4530), .A2(n4884), .A3(n4885), .ZN(n4523) );
  NOR3_X1 U3577 ( .A1(n4886), .A2(KEYINPUT82), .A3(KEYINPUT129), .ZN(n4885) );
  NOR2_X1 U3578 ( .A1(n4887), .A2(n4888), .ZN(n4886) );
  NOR2_X1 U3579 ( .A1(n4889), .A2(KEYINPUT33), .ZN(n4888) );
  NOR2_X1 U3580 ( .A1(n4890), .A2(n4505), .ZN(n4889) );
  NOR2_X1 U3581 ( .A1(n4459), .A2(KEYINPUT89), .ZN(n4505) );
  NOR2_X1 U3582 ( .A1(n4416), .A2(n4489), .ZN(n4459) );
  INV_X1 U3583 ( .A(n4441), .ZN(n4489) );
  NAND2_X1 U3584 ( .A1(n4413), .A2(n4478), .ZN(n4416) );
  NOR2_X1 U3585 ( .A1(n4437), .A2(n4479), .ZN(n4478) );
  NAND2_X1 U3586 ( .A1(n4434), .A2(n4401), .ZN(n4479) );
  NAND2_X1 U3587 ( .A1(G2211), .A2(n4023), .ZN(n4401) );
  INV_X1 U3588 ( .A(n4432), .ZN(n4434) );
  INV_X1 U3589 ( .A(n4508), .ZN(n4887) );
  NAND4_X1 U3590 ( .A1(n4891), .A2(n4892), .A3(n4540), .A4(n4893), .ZN(n4508) );
  NOR3_X1 U3591 ( .A1(KEYINPUT108), .A2(KEYINPUT77), .A3(KEYINPUT183), .ZN(n4893) );
  AND2_X1 U3592 ( .A1(n4894), .A2(n4895), .ZN(n4540) );
  NAND2_X1 U3593 ( .A1(n4274), .A2(n4272), .ZN(n4895) );
  OR2_X1 U3594 ( .A1(n4243), .A2(n4896), .ZN(n4272) );
  NOR2_X1 U3595 ( .A1(n4075), .A2(G4432), .ZN(n4896) );
  INV_X1 U3596 ( .A(n4897), .ZN(n4075) );
  NOR2_X1 U3597 ( .A1(n4248), .A2(n4270), .ZN(n4243) );
  INV_X1 U3598 ( .A(n4245), .ZN(n4270) );
  NAND2_X1 U3599 ( .A1(n4898), .A2(n4899), .ZN(n4245) );
  NAND2_X1 U3600 ( .A1(n4264), .A2(n4277), .ZN(n4899) );
  OR2_X1 U3601 ( .A1(n4073), .A2(G4427), .ZN(n4898) );
  NAND2_X1 U3602 ( .A1(n4074), .A2(n4900), .ZN(n4894) );
  INV_X1 U3603 ( .A(G4437), .ZN(n4900) );
  NAND2_X1 U3604 ( .A1(n4901), .A2(n4902), .ZN(n4892) );
  OR3_X1 U3605 ( .A1(KEYINPUT109), .A2(KEYINPUT59), .A3(n4252), .ZN(n4902) );
  NAND2_X1 U3606 ( .A1(n4903), .A2(n4904), .ZN(n4252) );
  NAND2_X1 U3607 ( .A1(n4231), .A2(n4226), .ZN(n4904) );
  NAND2_X1 U3608 ( .A1(n4905), .A2(n4906), .ZN(n4226) );
  OR2_X1 U3609 ( .A1(n4213), .A2(n4214), .ZN(n4906) );
  AND2_X1 U3610 ( .A1(n4292), .A2(n4907), .ZN(n4214) );
  NAND2_X1 U3611 ( .A1(n4281), .A2(n4298), .ZN(n4907) );
  NAND2_X1 U3612 ( .A1(n4908), .A2(n4909), .ZN(n4298) );
  NAND2_X1 U3613 ( .A1(n4224), .A2(n4232), .ZN(n4909) );
  NAND2_X1 U3614 ( .A1(n4081), .A2(n4802), .ZN(n4908) );
  INV_X1 U3615 ( .A(G4400), .ZN(n4802) );
  INV_X1 U3616 ( .A(n4910), .ZN(n4231) );
  NAND2_X1 U3617 ( .A1(n4079), .A2(n4817), .ZN(n4903) );
  INV_X1 U3618 ( .A(G4415), .ZN(n4817) );
  OR2_X1 U3619 ( .A1(n4550), .A2(KEYINPUT152), .ZN(n4901) );
  NAND2_X1 U3620 ( .A1(n4911), .A2(n4912), .ZN(n4891) );
  OR2_X1 U3621 ( .A1(KEYINPUT34), .A2(n4913), .ZN(n4912) );
  NOR2_X1 U3622 ( .A1(n4914), .A2(n4915), .ZN(n4913) );
  NOR2_X1 U3623 ( .A1(KEYINPUT152), .A2(n4550), .ZN(n4915) );
  AND2_X1 U3624 ( .A1(n4244), .A2(n4274), .ZN(n4550) );
  XNOR2_X1 U3625 ( .A(G4437), .B(n4074), .ZN(n4274) );
  NAND2_X1 U3626 ( .A1(n4916), .A2(n4917), .ZN(n4074) );
  NAND2_X1 U3627 ( .A1(G66), .A2(n3844), .ZN(n4917) );
  NAND2_X1 U3628 ( .A1(G219), .A2(G18), .ZN(n4916) );
  NOR2_X1 U3629 ( .A1(n4275), .A2(n4248), .ZN(n4244) );
  XOR2_X1 U3630 ( .A(G4432), .B(n4897), .Z(n4248) );
  NAND2_X1 U3631 ( .A1(n4918), .A2(n4919), .ZN(n4897) );
  NAND2_X1 U3632 ( .A1(G50), .A2(n3844), .ZN(n4919) );
  NAND2_X1 U3633 ( .A1(G220), .A2(G18), .ZN(n4918) );
  NAND2_X1 U3634 ( .A1(n4278), .A2(n4277), .ZN(n4275) );
  XOR2_X1 U3635 ( .A(G4427), .B(n4073), .Z(n4277) );
  AND2_X1 U3636 ( .A1(n4920), .A2(n4921), .ZN(n4073) );
  NAND2_X1 U3637 ( .A1(G32), .A2(n3844), .ZN(n4921) );
  NAND2_X1 U3638 ( .A1(G221), .A2(G18), .ZN(n4920) );
  NOR2_X1 U3639 ( .A1(n4264), .A2(n4249), .ZN(n4278) );
  AND2_X1 U3640 ( .A1(G4420), .A2(n4065), .ZN(n4249) );
  NOR2_X1 U3641 ( .A1(n4065), .A2(G4420), .ZN(n4264) );
  NAND2_X1 U3642 ( .A1(n4922), .A2(n4923), .ZN(n4065) );
  OR2_X1 U3643 ( .A1(G222), .A2(n3844), .ZN(n4923) );
  OR2_X1 U3644 ( .A1(G18), .A2(G35), .ZN(n4922) );
  NOR2_X1 U3645 ( .A1(KEYINPUT91), .A2(n4262), .ZN(n4914) );
  NOR3_X1 U3646 ( .A1(n4910), .A2(n4213), .A3(n4215), .ZN(n4262) );
  NAND3_X1 U3647 ( .A1(n4232), .A2(n4281), .A3(n4279), .ZN(n4215) );
  AND2_X1 U3648 ( .A1(n4283), .A2(n4216), .ZN(n4279) );
  NAND2_X1 U3649 ( .A1(G4394), .A2(n4072), .ZN(n4216) );
  INV_X1 U3650 ( .A(n4224), .ZN(n4283) );
  NOR2_X1 U3651 ( .A1(n4072), .A2(G4394), .ZN(n4224) );
  NAND2_X1 U3652 ( .A1(n4924), .A2(n4925), .ZN(n4072) );
  OR2_X1 U3653 ( .A1(G217), .A2(n3844), .ZN(n4925) );
  OR2_X1 U3654 ( .A1(G118), .A2(G18), .ZN(n4924) );
  INV_X1 U3655 ( .A(n4294), .ZN(n4281) );
  NAND2_X1 U3656 ( .A1(n4292), .A2(n4926), .ZN(n4294) );
  NAND2_X1 U3657 ( .A1(G4405), .A2(n4080), .ZN(n4926) );
  OR2_X1 U3658 ( .A1(n4080), .A2(G4405), .ZN(n4292) );
  NAND2_X1 U3659 ( .A1(n4927), .A2(n4928), .ZN(n4080) );
  OR2_X1 U3660 ( .A1(G225), .A2(n3844), .ZN(n4928) );
  OR2_X1 U3661 ( .A1(G18), .A2(G94), .ZN(n4927) );
  XNOR2_X1 U3662 ( .A(G4400), .B(n4081), .ZN(n4232) );
  NAND2_X1 U3663 ( .A1(n4929), .A2(n4804), .ZN(n4081) );
  NAND2_X1 U3664 ( .A1(G97), .A2(n3844), .ZN(n4804) );
  NAND2_X1 U3665 ( .A1(G226), .A2(G18), .ZN(n4929) );
  NAND2_X1 U3666 ( .A1(n4905), .A2(n4930), .ZN(n4213) );
  NAND2_X1 U3667 ( .A1(G4410), .A2(n4078), .ZN(n4930) );
  INV_X1 U3668 ( .A(n4212), .ZN(n4905) );
  NOR2_X1 U3669 ( .A1(n4078), .A2(G4410), .ZN(n4212) );
  NAND2_X1 U3670 ( .A1(n4931), .A2(n4932), .ZN(n4078) );
  OR2_X1 U3671 ( .A1(G224), .A2(n3844), .ZN(n4932) );
  OR2_X1 U3672 ( .A1(G121), .A2(G18), .ZN(n4931) );
  XOR2_X1 U3673 ( .A(G4415), .B(n4079), .Z(n4910) );
  NAND2_X1 U3674 ( .A1(n4933), .A2(n4819), .ZN(n4079) );
  NAND2_X1 U3675 ( .A1(G47), .A2(n3844), .ZN(n4819) );
  NAND2_X1 U3676 ( .A1(G223), .A2(G18), .ZN(n4933) );
  NAND4_X1 U3677 ( .A1(n4934), .A2(n4935), .A3(n4553), .A4(n4936), .ZN(n4911) );
  NOR4_X1 U3678 ( .A1(KEYINPUT75), .A2(KEYINPUT167), .A3(KEYINPUT101), .A4(n4937), .ZN(n4936) );
  NOR2_X1 U3679 ( .A1(n4317), .A2(n4938), .ZN(n4937) );
  AND2_X1 U3680 ( .A1(n4314), .A2(n4259), .ZN(n4938) );
  NOR4_X1 U3681 ( .A1(KEYINPUT102), .A2(n4561), .A3(KEYINPUT50), .A4(KEYINPUT170), .ZN(n4317) );
  NAND2_X1 U3682 ( .A1(n4939), .A2(n4940), .ZN(n4561) );
  NAND2_X1 U3683 ( .A1(n4941), .A2(n4114), .ZN(n4940) );
  NAND2_X1 U3684 ( .A1(n4100), .A2(n4942), .ZN(n4114) );
  NAND2_X1 U3685 ( .A1(n4107), .A2(n4943), .ZN(n4942) );
  INV_X1 U3686 ( .A(n4098), .ZN(n4943) );
  NOR2_X1 U3687 ( .A1(n4097), .A2(n4944), .ZN(n4098) );
  NOR2_X1 U3688 ( .A1(n4180), .A2(n4179), .ZN(n4097) );
  AND2_X1 U3689 ( .A1(n4945), .A2(n4946), .ZN(n4100) );
  NAND2_X1 U3690 ( .A1(n4093), .A2(n4104), .ZN(n4946) );
  INV_X1 U3691 ( .A(n4173), .ZN(n4104) );
  NAND2_X1 U3692 ( .A1(n4060), .A2(n4737), .ZN(n4945) );
  INV_X1 U3693 ( .A(G3717), .ZN(n4737) );
  INV_X1 U3694 ( .A(n4123), .ZN(n4941) );
  NAND2_X1 U3695 ( .A1(n4058), .A2(n4742), .ZN(n4939) );
  INV_X1 U3696 ( .A(G3723), .ZN(n4742) );
  INV_X1 U3697 ( .A(n4255), .ZN(n4553) );
  NAND2_X1 U3698 ( .A1(n4947), .A2(n4948), .ZN(n4255) );
  NAND2_X1 U3699 ( .A1(n4165), .A2(n4143), .ZN(n4948) );
  NAND2_X1 U3700 ( .A1(n4134), .A2(n4949), .ZN(n4143) );
  NAND2_X1 U3701 ( .A1(n4053), .A2(n4950), .ZN(n4949) );
  OR2_X1 U3702 ( .A1(n4137), .A2(n4139), .ZN(n4134) );
  INV_X1 U3703 ( .A(n4162), .ZN(n4139) );
  NAND2_X1 U3704 ( .A1(n4951), .A2(n4952), .ZN(n4162) );
  OR2_X1 U3705 ( .A1(n4152), .A2(n4167), .ZN(n4952) );
  NAND2_X1 U3706 ( .A1(n4054), .A2(n4953), .ZN(n4951) );
  INV_X1 U3707 ( .A(G3737), .ZN(n4953) );
  OR2_X1 U3708 ( .A1(n4057), .A2(G3749), .ZN(n4947) );
  NAND2_X1 U3709 ( .A1(n4315), .A2(n4954), .ZN(n4935) );
  NAND2_X1 U3710 ( .A1(n4314), .A2(n4259), .ZN(n4954) );
  NAND2_X1 U3711 ( .A1(n4140), .A2(n4165), .ZN(n4259) );
  XOR2_X1 U3712 ( .A(n4057), .B(G3749), .Z(n4165) );
  NAND2_X1 U3713 ( .A1(n4749), .A2(n4955), .ZN(n4057) );
  OR2_X1 U3714 ( .A1(G231), .A2(n3844), .ZN(n4955) );
  NAND2_X1 U3715 ( .A1(n4956), .A2(n3844), .ZN(n4749) );
  INV_X1 U3716 ( .A(G100), .ZN(n4956) );
  NOR2_X1 U3717 ( .A1(n4138), .A2(n4137), .ZN(n4140) );
  XNOR2_X1 U3718 ( .A(n4053), .B(n4950), .ZN(n4137) );
  INV_X1 U3719 ( .A(G3743), .ZN(n4950) );
  AND2_X1 U3720 ( .A1(n4754), .A2(n4957), .ZN(n4053) );
  OR2_X1 U3721 ( .A1(G232), .A2(n3844), .ZN(n4957) );
  NAND2_X1 U3722 ( .A1(n4958), .A2(n3844), .ZN(n4754) );
  INV_X1 U3723 ( .A(G124), .ZN(n4958) );
  OR2_X1 U3724 ( .A1(n4168), .A2(n4167), .ZN(n4138) );
  XOR2_X1 U3725 ( .A(G3737), .B(n4054), .Z(n4167) );
  NAND2_X1 U3726 ( .A1(n4959), .A2(n4960), .ZN(n4054) );
  NAND2_X1 U3727 ( .A1(G127), .A2(n3844), .ZN(n4960) );
  NAND2_X1 U3728 ( .A1(G233), .A2(G18), .ZN(n4959) );
  NAND2_X1 U3729 ( .A1(n4152), .A2(n4141), .ZN(n4168) );
  NAND2_X1 U3730 ( .A1(G3729), .A2(n4046), .ZN(n4141) );
  INV_X1 U3731 ( .A(n4159), .ZN(n4152) );
  NOR2_X1 U3732 ( .A1(n4046), .A2(G3729), .ZN(n4159) );
  NAND2_X1 U3733 ( .A1(n4961), .A2(n4962), .ZN(n4046) );
  OR2_X1 U3734 ( .A1(G234), .A2(n3844), .ZN(n4962) );
  OR2_X1 U3735 ( .A1(G130), .A2(G18), .ZN(n4961) );
  INV_X1 U3736 ( .A(KEYINPUT149), .ZN(n4314) );
  AND2_X1 U3737 ( .A1(G4526), .A2(n4963), .ZN(n4315) );
  OR2_X1 U3738 ( .A1(KEYINPUT121), .A2(n4560), .ZN(n4963) );
  NOR2_X1 U3739 ( .A1(n4123), .A2(n4115), .ZN(n4560) );
  NAND3_X1 U3740 ( .A1(n4107), .A2(n4176), .A3(n4177), .ZN(n4115) );
  NOR2_X1 U3741 ( .A1(n4091), .A2(n4111), .ZN(n4177) );
  NOR3_X1 U3742 ( .A1(n4051), .A2(G18), .A3(n4964), .ZN(n4111) );
  INV_X1 U3743 ( .A(n4180), .ZN(n4091) );
  NAND3_X1 U3744 ( .A1(n3844), .A2(n4964), .A3(n4051), .ZN(n4180) );
  AND2_X1 U3745 ( .A1(n4965), .A2(n4966), .ZN(n4051) );
  OR2_X1 U3746 ( .A1(G229), .A2(n3844), .ZN(n4966) );
  OR2_X1 U3747 ( .A1(G18), .A2(G41), .ZN(n4965) );
  INV_X1 U3748 ( .A(G3701), .ZN(n4964) );
  INV_X1 U3749 ( .A(n4179), .ZN(n4176) );
  NAND2_X1 U3750 ( .A1(n4105), .A2(n4967), .ZN(n4179) );
  NAND2_X1 U3751 ( .A1(G3705), .A2(n4040), .ZN(n4967) );
  INV_X1 U3752 ( .A(n4944), .ZN(n4105) );
  NOR2_X1 U3753 ( .A1(n4040), .A2(G3705), .ZN(n4944) );
  AND2_X1 U3754 ( .A1(n4968), .A2(n4726), .ZN(n4040) );
  NAND2_X1 U3755 ( .A1(G29), .A2(n3844), .ZN(n4726) );
  NAND2_X1 U3756 ( .A1(G238), .A2(G18), .ZN(n4968) );
  NOR2_X1 U3757 ( .A1(n4106), .A2(n4173), .ZN(n4107) );
  XOR2_X1 U3758 ( .A(G3717), .B(n4060), .Z(n4173) );
  NAND2_X1 U3759 ( .A1(n4969), .A2(n4739), .ZN(n4060) );
  NAND2_X1 U3760 ( .A1(G23), .A2(n3844), .ZN(n4739) );
  NAND2_X1 U3761 ( .A1(G236), .A2(G18), .ZN(n4969) );
  INV_X1 U3762 ( .A(n4096), .ZN(n4106) );
  NOR2_X1 U3763 ( .A1(n4093), .A2(n4970), .ZN(n4096) );
  AND2_X1 U3764 ( .A1(G3711), .A2(n4059), .ZN(n4970) );
  NOR2_X1 U3765 ( .A1(n4059), .A2(G3711), .ZN(n4093) );
  NAND2_X1 U3766 ( .A1(n4971), .A2(n4972), .ZN(n4059) );
  OR2_X1 U3767 ( .A1(G237), .A2(n3844), .ZN(n4972) );
  OR2_X1 U3768 ( .A1(G18), .A2(G26), .ZN(n4971) );
  XOR2_X1 U3769 ( .A(G3723), .B(n4058), .Z(n4123) );
  NAND2_X1 U3770 ( .A1(n4973), .A2(n4744), .ZN(n4058) );
  NAND2_X1 U3771 ( .A1(G103), .A2(n3844), .ZN(n4744) );
  NAND2_X1 U3772 ( .A1(G235), .A2(G18), .ZN(n4973) );
  NAND2_X1 U3773 ( .A1(KEYINPUT37), .A2(G4526), .ZN(n4934) );
  NAND2_X1 U3774 ( .A1(n4504), .A2(n4974), .ZN(n4884) );
  INV_X1 U3775 ( .A(n4890), .ZN(n4974) );
  NOR2_X1 U3776 ( .A1(KEYINPUT159), .A2(n4539), .ZN(n4890) );
  NOR3_X1 U3777 ( .A1(n4475), .A2(n4465), .A3(n4470), .ZN(n4539) );
  NAND2_X1 U3778 ( .A1(n4472), .A2(n4473), .ZN(n4470) );
  XNOR2_X1 U3779 ( .A(G2239), .B(n4975), .ZN(n4472) );
  OR3_X1 U3780 ( .A1(KEYINPUT62), .A2(KEYINPUT116), .A3(n4456), .ZN(n4504) );
  NAND2_X1 U3781 ( .A1(n4976), .A2(n4977), .ZN(n4456) );
  NAND2_X1 U3782 ( .A1(n4441), .A2(n4418), .ZN(n4977) );
  NAND2_X1 U3783 ( .A1(n4427), .A2(n4978), .ZN(n4418) );
  NAND2_X1 U3784 ( .A1(n4413), .A2(n4493), .ZN(n4978) );
  NAND2_X1 U3785 ( .A1(n4438), .A2(n4979), .ZN(n4493) );
  NAND2_X1 U3786 ( .A1(n4432), .A2(n4431), .ZN(n4979) );
  INV_X1 U3787 ( .A(n4437), .ZN(n4431) );
  NAND2_X1 U3788 ( .A1(n4438), .A2(n4980), .ZN(n4437) );
  NAND2_X1 U3789 ( .A1(G2218), .A2(n4024), .ZN(n4980) );
  NOR2_X1 U3790 ( .A1(n4023), .A2(G2211), .ZN(n4432) );
  NAND2_X1 U3791 ( .A1(n4981), .A2(n4982), .ZN(n4023) );
  OR2_X1 U3792 ( .A1(G151), .A2(n3844), .ZN(n4982) );
  OR2_X1 U3793 ( .A1(G147), .A2(G18), .ZN(n4981) );
  OR2_X1 U3794 ( .A1(n4024), .A2(G2218), .ZN(n4438) );
  AND2_X1 U3795 ( .A1(n4983), .A2(n4638), .ZN(n4024) );
  NAND2_X1 U3796 ( .A1(G138), .A2(n3844), .ZN(n4638) );
  NAND2_X1 U3797 ( .A1(G160), .A2(G18), .ZN(n4983) );
  NOR2_X1 U3798 ( .A1(n4411), .A2(n4409), .ZN(n4413) );
  INV_X1 U3799 ( .A(n4400), .ZN(n4411) );
  NOR2_X1 U3800 ( .A1(n4397), .A2(n4984), .ZN(n4400) );
  AND2_X1 U3801 ( .A1(G2224), .A2(n4016), .ZN(n4984) );
  AND2_X1 U3802 ( .A1(n4985), .A2(n4986), .ZN(n4427) );
  NAND2_X1 U3803 ( .A1(n4397), .A2(n4410), .ZN(n4986) );
  INV_X1 U3804 ( .A(n4409), .ZN(n4410) );
  XOR2_X1 U3805 ( .A(G2230), .B(n4025), .Z(n4409) );
  NOR2_X1 U3806 ( .A1(n4016), .A2(G2224), .ZN(n4397) );
  AND2_X1 U3807 ( .A1(n4987), .A2(n4642), .ZN(n4016) );
  NAND2_X1 U3808 ( .A1(G144), .A2(n3844), .ZN(n4642) );
  NAND2_X1 U3809 ( .A1(G159), .A2(G18), .ZN(n4987) );
  NAND2_X1 U3810 ( .A1(n4025), .A2(n4645), .ZN(n4985) );
  INV_X1 U3811 ( .A(G2230), .ZN(n4645) );
  NAND2_X1 U3812 ( .A1(n4988), .A2(n4647), .ZN(n4025) );
  NAND2_X1 U3813 ( .A1(G135), .A2(n3844), .ZN(n4647) );
  NAND2_X1 U3814 ( .A1(G158), .A2(G18), .ZN(n4988) );
  XOR2_X1 U3815 ( .A(n4652), .B(n4026), .Z(n4441) );
  NAND2_X1 U3816 ( .A1(n4026), .A2(n4652), .ZN(n4976) );
  INV_X1 U3817 ( .A(G2236), .ZN(n4652) );
  NAND2_X1 U3818 ( .A1(n4648), .A2(n4989), .ZN(n4026) );
  NAND2_X1 U3819 ( .A1(G157), .A2(n3860), .ZN(n4989) );
  AND2_X1 U3820 ( .A1(n4990), .A2(n4991), .ZN(n4530) );
  NAND2_X1 U3821 ( .A1(n4468), .A2(n4507), .ZN(n4991) );
  NAND2_X1 U3822 ( .A1(n4992), .A2(n4993), .ZN(n4507) );
  NAND2_X1 U3823 ( .A1(n4498), .A2(n4454), .ZN(n4993) );
  NAND2_X1 U3824 ( .A1(n4994), .A2(n4995), .ZN(n4454) );
  NAND2_X1 U3825 ( .A1(n4497), .A2(n4473), .ZN(n4995) );
  XNOR2_X1 U3826 ( .A(G2247), .B(n4010), .ZN(n4473) );
  NOR2_X1 U3827 ( .A1(n4011), .A2(G2239), .ZN(n4497) );
  INV_X1 U3828 ( .A(n4975), .ZN(n4011) );
  NAND2_X1 U3829 ( .A1(n4648), .A2(n4996), .ZN(n4975) );
  NAND2_X1 U3830 ( .A1(G156), .A2(n3860), .ZN(n4996) );
  NAND2_X1 U3831 ( .A1(n4010), .A2(n4672), .ZN(n4994) );
  INV_X1 U3832 ( .A(G2247), .ZN(n4672) );
  NAND2_X1 U3833 ( .A1(n4648), .A2(n4997), .ZN(n4010) );
  NAND2_X1 U3834 ( .A1(G155), .A2(n3860), .ZN(n4997) );
  INV_X1 U3835 ( .A(n4465), .ZN(n4498) );
  XOR2_X1 U3836 ( .A(G2253), .B(n4013), .Z(n4465) );
  NAND2_X1 U3837 ( .A1(n4013), .A2(n4676), .ZN(n4992) );
  INV_X1 U3838 ( .A(G2253), .ZN(n4676) );
  NAND2_X1 U3839 ( .A1(n4648), .A2(n4998), .ZN(n4013) );
  NAND2_X1 U3840 ( .A1(G154), .A2(n3860), .ZN(n4998) );
  INV_X1 U3841 ( .A(n4475), .ZN(n4468) );
  XOR2_X1 U3842 ( .A(G2256), .B(n4012), .Z(n4475) );
  NAND2_X1 U3843 ( .A1(n4012), .A2(n4657), .ZN(n4990) );
  INV_X1 U3844 ( .A(G2256), .ZN(n4657) );
  NAND2_X1 U3845 ( .A1(n4648), .A2(n4999), .ZN(n4012) );
  NAND2_X1 U3846 ( .A1(G153), .A2(n3860), .ZN(n4999) );
  NAND2_X1 U3847 ( .A1(n5000), .A2(n4562), .ZN(n4522) );
  NAND3_X1 U3848 ( .A1(n4374), .A2(n4349), .A3(n4334), .ZN(n4562) );
  NOR3_X1 U3849 ( .A1(n4368), .A2(n4343), .A3(n4385), .ZN(n4334) );
  NAND2_X1 U3850 ( .A1(n4326), .A2(n4369), .ZN(n4385) );
  INV_X1 U3851 ( .A(n4365), .ZN(n4369) );
  NAND2_X1 U3852 ( .A1(G1462), .A2(n4038), .ZN(n4326) );
  INV_X1 U3853 ( .A(KEYINPUT95), .ZN(n5000) );
  NAND2_X1 U3854 ( .A1(n5001), .A2(n5002), .ZN(n4524) );
  NAND2_X1 U3855 ( .A1(n4349), .A2(n4340), .ZN(n5002) );
  NAND2_X1 U3856 ( .A1(n5003), .A2(n5004), .ZN(n4340) );
  NAND2_X1 U3857 ( .A1(n4374), .A2(n4333), .ZN(n5004) );
  NAND2_X1 U3858 ( .A1(n4379), .A2(n5005), .ZN(n4333) );
  NAND2_X1 U3859 ( .A1(n4372), .A2(n4366), .ZN(n5005) );
  NAND2_X1 U3860 ( .A1(n5006), .A2(n5007), .ZN(n4366) );
  NAND2_X1 U3861 ( .A1(n4365), .A2(n4347), .ZN(n5007) );
  INV_X1 U3862 ( .A(n4368), .ZN(n4347) );
  XNOR2_X1 U3863 ( .A(n4031), .B(G1469), .ZN(n4368) );
  NOR2_X1 U3864 ( .A1(n4038), .A2(G1462), .ZN(n4365) );
  NAND2_X1 U3865 ( .A1(n5008), .A2(n3860), .ZN(n4038) );
  OR2_X1 U3866 ( .A1(n3866), .A2(G209), .ZN(n5008) );
  OR2_X1 U3867 ( .A1(n4031), .A2(G1469), .ZN(n5006) );
  NAND2_X1 U3868 ( .A1(n3860), .A2(n5009), .ZN(n4031) );
  OR2_X1 U3869 ( .A1(G216), .A2(n3866), .ZN(n5009) );
  INV_X1 U3870 ( .A(n4343), .ZN(n4372) );
  NAND2_X1 U3871 ( .A1(n4379), .A2(n5010), .ZN(n4343) );
  NAND2_X1 U3872 ( .A1(G106), .A2(n4032), .ZN(n5010) );
  OR2_X1 U3873 ( .A1(n4032), .A2(G106), .ZN(n4379) );
  NAND2_X1 U3874 ( .A1(n3860), .A2(n5011), .ZN(n4032) );
  OR2_X1 U3875 ( .A1(G215), .A2(n3866), .ZN(n5011) );
  INV_X1 U3876 ( .A(n4648), .ZN(n3866) );
  INV_X1 U3877 ( .A(n4332), .ZN(n4374) );
  NAND2_X1 U3878 ( .A1(n5003), .A2(n5012), .ZN(n4332) );
  NAND2_X1 U3879 ( .A1(G1480), .A2(n4036), .ZN(n5012) );
  INV_X1 U3880 ( .A(n4331), .ZN(n5003) );
  NOR2_X1 U3881 ( .A1(n4036), .A2(G1480), .ZN(n4331) );
  AND2_X1 U3882 ( .A1(n4648), .A2(n5013), .ZN(n4036) );
  NAND2_X1 U3883 ( .A1(G214), .A2(n3860), .ZN(n5013) );
  XNOR2_X1 U3884 ( .A(G1486), .B(n4039), .ZN(n4349) );
  NAND2_X1 U3885 ( .A1(n4039), .A2(n5014), .ZN(n5001) );
  INV_X1 U3886 ( .A(G1486), .ZN(n5014) );
  NAND2_X1 U3887 ( .A1(n5015), .A2(n4648), .ZN(n4039) );
  NAND2_X1 U3888 ( .A1(n3844), .A2(n3860), .ZN(n4648) );
  NAND2_X1 U3889 ( .A1(G213), .A2(n3860), .ZN(n5015) );
  NAND2_X1 U3890 ( .A1(G9), .A2(G12), .ZN(n3860) );
  NOR2_X1 U3891 ( .A1(n3812), .A2(n3807), .ZN(n4512) );
  NAND2_X1 U3892 ( .A1(n3814), .A2(n5016), .ZN(n3807) );
  NAND2_X1 U3893 ( .A1(G38), .A2(n5017), .ZN(n5016) );
  NAND2_X1 U3894 ( .A1(n4358), .A2(n4359), .ZN(n3814) );
  INV_X1 U3895 ( .A(n5017), .ZN(n4358) );
  NAND2_X1 U3896 ( .A1(G4528), .A2(G1492), .ZN(n5017) );
  XOR2_X1 U3897 ( .A(n5018), .B(n4359), .Z(n3812) );
  INV_X1 U3898 ( .A(G38), .ZN(n4359) );
  NAND2_X1 U3899 ( .A1(G1496), .A2(G4528), .ZN(n5018) );
endmodule

