//Key = 0100010011001100010010010010110110010011100110010100100010101110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314;

XNOR2_X1 U726 ( .A(G107), .B(n1009), .ZN(G9) );
NAND4_X1 U727 ( .A1(n1010), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1009) );
NOR2_X1 U728 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
XOR2_X1 U729 ( .A(n1016), .B(KEYINPUT6), .Z(n1015) );
NOR2_X1 U730 ( .A1(n1017), .A2(n1018), .ZN(G75) );
NOR4_X1 U731 ( .A1(G953), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1018) );
NOR2_X1 U732 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U733 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U734 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR2_X1 U735 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NOR2_X1 U736 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR3_X1 U737 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1030) );
NOR2_X1 U738 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U739 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U740 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR3_X1 U741 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1033) );
NOR2_X1 U742 ( .A1(n1044), .A2(n1045), .ZN(n1032) );
XOR2_X1 U743 ( .A(KEYINPUT20), .B(n1046), .Z(n1045) );
NOR3_X1 U744 ( .A1(n1041), .A2(n1047), .A3(n1036), .ZN(n1028) );
NOR2_X1 U745 ( .A1(n1048), .A2(n1010), .ZN(n1047) );
NOR2_X1 U746 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR4_X1 U747 ( .A1(n1051), .A2(n1036), .A3(n1041), .A4(n1031), .ZN(n1024) );
NOR3_X1 U748 ( .A1(n1019), .A2(G953), .A3(G952), .ZN(n1017) );
AND4_X1 U749 ( .A1(n1052), .A2(n1042), .A3(n1053), .A4(n1054), .ZN(n1019) );
NOR4_X1 U750 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
XNOR2_X1 U751 ( .A(n1059), .B(n1060), .ZN(n1058) );
XNOR2_X1 U752 ( .A(n1061), .B(n1062), .ZN(n1057) );
XOR2_X1 U753 ( .A(n1063), .B(KEYINPUT55), .Z(n1062) );
AND2_X1 U754 ( .A1(n1031), .A2(KEYINPUT58), .ZN(n1056) );
INV_X1 U755 ( .A(n1064), .ZN(n1031) );
NOR2_X1 U756 ( .A1(KEYINPUT58), .A2(n1010), .ZN(n1055) );
NOR2_X1 U757 ( .A1(n1065), .A2(n1066), .ZN(n1053) );
XOR2_X1 U758 ( .A(n1067), .B(n1068), .Z(n1066) );
XNOR2_X1 U759 ( .A(KEYINPUT26), .B(KEYINPUT15), .ZN(n1067) );
INV_X1 U760 ( .A(n1040), .ZN(n1065) );
XNOR2_X1 U761 ( .A(n1069), .B(G478), .ZN(n1052) );
XOR2_X1 U762 ( .A(n1070), .B(n1071), .Z(G72) );
NOR2_X1 U763 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U764 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NAND2_X1 U765 ( .A1(n1076), .A2(n1077), .ZN(n1070) );
NAND2_X1 U766 ( .A1(n1078), .A2(n1073), .ZN(n1077) );
XOR2_X1 U767 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND2_X1 U768 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
XNOR2_X1 U769 ( .A(KEYINPUT61), .B(n1083), .ZN(n1082) );
NAND3_X1 U770 ( .A1(n1080), .A2(G900), .A3(G953), .ZN(n1076) );
AND3_X1 U771 ( .A1(n1084), .A2(n1085), .A3(KEYINPUT23), .ZN(n1080) );
NAND2_X1 U772 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U773 ( .A(KEYINPUT49), .B(n1088), .Z(n1084) );
NOR2_X1 U774 ( .A1(n1089), .A2(n1087), .ZN(n1088) );
XOR2_X1 U775 ( .A(n1090), .B(n1091), .Z(n1087) );
NAND3_X1 U776 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1090) );
NAND2_X1 U777 ( .A1(KEYINPUT46), .A2(n1095), .ZN(n1094) );
NAND3_X1 U778 ( .A1(n1096), .A2(n1097), .A3(G131), .ZN(n1093) );
INV_X1 U779 ( .A(KEYINPUT46), .ZN(n1097) );
OR2_X1 U780 ( .A1(n1096), .A2(G131), .ZN(n1092) );
NOR2_X1 U781 ( .A1(KEYINPUT41), .A2(n1095), .ZN(n1096) );
XOR2_X1 U782 ( .A(n1098), .B(n1099), .Z(n1095) );
NOR2_X1 U783 ( .A1(G134), .A2(KEYINPUT0), .ZN(n1099) );
XOR2_X1 U784 ( .A(n1086), .B(KEYINPUT53), .Z(n1089) );
XOR2_X1 U785 ( .A(n1100), .B(n1101), .Z(G69) );
NOR2_X1 U786 ( .A1(n1102), .A2(n1073), .ZN(n1101) );
AND2_X1 U787 ( .A1(G898), .A2(G224), .ZN(n1102) );
NOR3_X1 U788 ( .A1(KEYINPUT37), .A2(n1103), .A3(n1104), .ZN(n1100) );
NOR2_X1 U789 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NOR2_X1 U790 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
XOR2_X1 U791 ( .A(n1109), .B(KEYINPUT43), .Z(n1108) );
NOR2_X1 U792 ( .A1(G898), .A2(n1073), .ZN(n1107) );
AND2_X1 U793 ( .A1(n1109), .A2(n1106), .ZN(n1103) );
XOR2_X1 U794 ( .A(n1110), .B(n1111), .Z(n1106) );
XOR2_X1 U795 ( .A(n1112), .B(n1113), .Z(n1110) );
NAND2_X1 U796 ( .A1(n1073), .A2(n1114), .ZN(n1109) );
NOR2_X1 U797 ( .A1(n1115), .A2(n1116), .ZN(G66) );
XOR2_X1 U798 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NOR2_X1 U800 ( .A1(n1115), .A2(n1121), .ZN(G63) );
NOR3_X1 U801 ( .A1(n1069), .A2(n1122), .A3(n1123), .ZN(n1121) );
AND3_X1 U802 ( .A1(n1124), .A2(G478), .A3(n1125), .ZN(n1123) );
NOR2_X1 U803 ( .A1(n1126), .A2(n1124), .ZN(n1122) );
AND2_X1 U804 ( .A1(n1021), .A2(G478), .ZN(n1126) );
NOR2_X1 U805 ( .A1(n1115), .A2(n1127), .ZN(G60) );
XNOR2_X1 U806 ( .A(n1128), .B(n1129), .ZN(n1127) );
AND2_X1 U807 ( .A1(G475), .A2(n1125), .ZN(n1129) );
NAND3_X1 U808 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(G6) );
NAND2_X1 U809 ( .A1(KEYINPUT51), .A2(n1133), .ZN(n1132) );
OR3_X1 U810 ( .A1(n1133), .A2(KEYINPUT51), .A3(G104), .ZN(n1131) );
NAND2_X1 U811 ( .A1(G104), .A2(n1134), .ZN(n1130) );
NAND2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
INV_X1 U813 ( .A(KEYINPUT51), .ZN(n1136) );
XNOR2_X1 U814 ( .A(KEYINPUT10), .B(n1133), .ZN(n1135) );
NOR2_X1 U815 ( .A1(n1115), .A2(n1137), .ZN(G57) );
XOR2_X1 U816 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U817 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR3_X1 U818 ( .A1(n1120), .A2(KEYINPUT50), .A3(n1063), .ZN(n1141) );
INV_X1 U819 ( .A(G472), .ZN(n1063) );
XNOR2_X1 U820 ( .A(n1142), .B(n1143), .ZN(n1138) );
NOR2_X1 U821 ( .A1(n1115), .A2(n1144), .ZN(G54) );
XOR2_X1 U822 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U823 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U824 ( .A(n1149), .B(n1150), .ZN(n1145) );
AND2_X1 U825 ( .A1(G469), .A2(n1125), .ZN(n1150) );
INV_X1 U826 ( .A(n1120), .ZN(n1125) );
NOR2_X1 U827 ( .A1(n1115), .A2(n1151), .ZN(G51) );
XOR2_X1 U828 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U829 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U830 ( .A1(n1060), .A2(n1120), .ZN(n1155) );
NAND2_X1 U831 ( .A1(G902), .A2(n1021), .ZN(n1120) );
NAND3_X1 U832 ( .A1(n1156), .A2(n1083), .A3(n1081), .ZN(n1021) );
AND4_X1 U833 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1081) );
NOR4_X1 U834 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1160) );
INV_X1 U835 ( .A(n1165), .ZN(n1162) );
NAND3_X1 U836 ( .A1(n1011), .A2(n1038), .A3(n1166), .ZN(n1159) );
INV_X1 U837 ( .A(n1114), .ZN(n1156) );
NAND4_X1 U838 ( .A1(n1167), .A2(n1133), .A3(n1168), .A4(n1169), .ZN(n1114) );
NOR4_X1 U839 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1169) );
NAND2_X1 U840 ( .A1(n1174), .A2(n1175), .ZN(n1168) );
INV_X1 U841 ( .A(n1051), .ZN(n1175) );
NOR2_X1 U842 ( .A1(n1176), .A2(n1011), .ZN(n1051) );
NAND4_X1 U843 ( .A1(n1177), .A2(n1176), .A3(n1010), .A4(n1013), .ZN(n1133) );
NAND4_X1 U844 ( .A1(n1177), .A2(n1010), .A3(n1011), .A4(n1013), .ZN(n1167) );
INV_X1 U845 ( .A(n1036), .ZN(n1013) );
NAND2_X1 U846 ( .A1(n1178), .A2(KEYINPUT5), .ZN(n1154) );
XOR2_X1 U847 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U848 ( .A1(KEYINPUT27), .A2(n1181), .ZN(n1180) );
XNOR2_X1 U849 ( .A(G125), .B(n1182), .ZN(n1179) );
NOR2_X1 U850 ( .A1(n1073), .A2(G952), .ZN(n1115) );
XNOR2_X1 U851 ( .A(n1157), .B(n1183), .ZN(G48) );
XOR2_X1 U852 ( .A(KEYINPUT25), .B(G146), .Z(n1183) );
NAND3_X1 U853 ( .A1(n1176), .A2(n1038), .A3(n1166), .ZN(n1157) );
XNOR2_X1 U854 ( .A(n1158), .B(n1184), .ZN(G45) );
NOR2_X1 U855 ( .A1(KEYINPUT48), .A2(n1185), .ZN(n1184) );
NAND4_X1 U856 ( .A1(n1186), .A2(n1038), .A3(n1187), .A4(n1068), .ZN(n1158) );
XOR2_X1 U857 ( .A(G140), .B(n1164), .Z(G42) );
AND3_X1 U858 ( .A1(n1046), .A2(n1010), .A3(n1188), .ZN(n1164) );
XOR2_X1 U859 ( .A(n1189), .B(n1163), .Z(G39) );
AND3_X1 U860 ( .A1(n1166), .A2(n1046), .A3(n1190), .ZN(n1163) );
NAND2_X1 U861 ( .A1(KEYINPUT28), .A2(n1098), .ZN(n1189) );
XNOR2_X1 U862 ( .A(G134), .B(n1083), .ZN(G36) );
NAND3_X1 U863 ( .A1(n1186), .A2(n1011), .A3(n1046), .ZN(n1083) );
XOR2_X1 U864 ( .A(n1191), .B(n1165), .Z(G33) );
NAND3_X1 U865 ( .A1(n1046), .A2(n1186), .A3(n1176), .ZN(n1165) );
AND3_X1 U866 ( .A1(n1010), .A2(n1192), .A3(n1193), .ZN(n1186) );
INV_X1 U867 ( .A(n1041), .ZN(n1046) );
NAND2_X1 U868 ( .A1(n1194), .A2(n1040), .ZN(n1041) );
XOR2_X1 U869 ( .A(G128), .B(n1195), .Z(G30) );
NOR3_X1 U870 ( .A1(n1016), .A2(KEYINPUT18), .A3(n1196), .ZN(n1195) );
XOR2_X1 U871 ( .A(n1197), .B(KEYINPUT54), .Z(n1196) );
NAND2_X1 U872 ( .A1(n1166), .A2(n1011), .ZN(n1197) );
AND4_X1 U873 ( .A1(n1010), .A2(n1198), .A3(n1199), .A4(n1192), .ZN(n1166) );
XOR2_X1 U874 ( .A(G101), .B(n1172), .Z(G3) );
AND4_X1 U875 ( .A1(n1177), .A2(n1190), .A3(n1193), .A4(n1010), .ZN(n1172) );
XNOR2_X1 U876 ( .A(n1161), .B(n1200), .ZN(G27) );
NAND2_X1 U877 ( .A1(KEYINPUT44), .A2(G125), .ZN(n1200) );
AND3_X1 U878 ( .A1(n1188), .A2(n1038), .A3(n1064), .ZN(n1161) );
AND4_X1 U879 ( .A1(n1201), .A2(n1176), .A3(n1199), .A4(n1192), .ZN(n1188) );
NAND2_X1 U880 ( .A1(n1202), .A2(n1023), .ZN(n1192) );
NAND3_X1 U881 ( .A1(n1203), .A2(n1075), .A3(n1204), .ZN(n1202) );
XOR2_X1 U882 ( .A(n1073), .B(KEYINPUT52), .Z(n1204) );
INV_X1 U883 ( .A(G900), .ZN(n1075) );
XOR2_X1 U884 ( .A(G122), .B(n1173), .Z(G24) );
AND3_X1 U885 ( .A1(n1177), .A2(n1064), .A3(n1205), .ZN(n1173) );
NOR3_X1 U886 ( .A1(n1036), .A2(n1206), .A3(n1207), .ZN(n1205) );
NAND2_X1 U887 ( .A1(n1042), .A2(n1201), .ZN(n1036) );
XNOR2_X1 U888 ( .A(G119), .B(n1208), .ZN(G21) );
NAND2_X1 U889 ( .A1(KEYINPUT32), .A2(n1171), .ZN(n1208) );
AND3_X1 U890 ( .A1(n1064), .A2(n1198), .A3(n1209), .ZN(n1171) );
XNOR2_X1 U891 ( .A(n1210), .B(n1211), .ZN(G18) );
NAND2_X1 U892 ( .A1(KEYINPUT39), .A2(n1212), .ZN(n1210) );
NAND2_X1 U893 ( .A1(n1174), .A2(n1011), .ZN(n1212) );
NOR2_X1 U894 ( .A1(n1068), .A2(n1207), .ZN(n1011) );
INV_X1 U895 ( .A(n1206), .ZN(n1068) );
AND3_X1 U896 ( .A1(n1064), .A2(n1193), .A3(n1177), .ZN(n1174) );
XOR2_X1 U897 ( .A(n1213), .B(n1214), .Z(G15) );
NAND4_X1 U898 ( .A1(n1064), .A2(n1176), .A3(n1215), .A4(n1193), .ZN(n1214) );
INV_X1 U899 ( .A(n1044), .ZN(n1193) );
NAND2_X1 U900 ( .A1(n1042), .A2(n1198), .ZN(n1044) );
XOR2_X1 U901 ( .A(n1043), .B(KEYINPUT30), .Z(n1198) );
INV_X1 U902 ( .A(n1201), .ZN(n1043) );
NOR2_X1 U903 ( .A1(n1014), .A2(n1216), .ZN(n1215) );
XOR2_X1 U904 ( .A(n1016), .B(KEYINPUT59), .Z(n1216) );
NOR2_X1 U905 ( .A1(n1217), .A2(n1218), .ZN(n1014) );
INV_X1 U906 ( .A(n1023), .ZN(n1218) );
INV_X1 U907 ( .A(n1219), .ZN(n1217) );
NOR2_X1 U908 ( .A1(n1187), .A2(n1206), .ZN(n1176) );
NOR2_X1 U909 ( .A1(n1049), .A2(n1220), .ZN(n1064) );
INV_X1 U910 ( .A(n1050), .ZN(n1220) );
XOR2_X1 U911 ( .A(n1170), .B(n1221), .Z(G12) );
XOR2_X1 U912 ( .A(KEYINPUT22), .B(G110), .Z(n1221) );
AND3_X1 U913 ( .A1(n1201), .A2(n1010), .A3(n1209), .ZN(n1170) );
AND3_X1 U914 ( .A1(n1190), .A2(n1199), .A3(n1177), .ZN(n1209) );
AND2_X1 U915 ( .A1(n1038), .A2(n1222), .ZN(n1177) );
NAND2_X1 U916 ( .A1(n1219), .A2(n1023), .ZN(n1222) );
NAND3_X1 U917 ( .A1(n1223), .A2(n1073), .A3(G952), .ZN(n1023) );
NAND3_X1 U918 ( .A1(n1203), .A2(n1224), .A3(G953), .ZN(n1219) );
XOR2_X1 U919 ( .A(KEYINPUT1), .B(G898), .Z(n1224) );
AND2_X1 U920 ( .A1(n1225), .A2(n1223), .ZN(n1203) );
NAND2_X1 U921 ( .A1(G237), .A2(G234), .ZN(n1223) );
XOR2_X1 U922 ( .A(n1226), .B(KEYINPUT29), .Z(n1225) );
INV_X1 U923 ( .A(n1016), .ZN(n1038) );
NAND2_X1 U924 ( .A1(n1039), .A2(n1040), .ZN(n1016) );
NAND2_X1 U925 ( .A1(G214), .A2(n1227), .ZN(n1040) );
INV_X1 U926 ( .A(n1194), .ZN(n1039) );
XNOR2_X1 U927 ( .A(n1228), .B(n1060), .ZN(n1194) );
NAND2_X1 U928 ( .A1(G210), .A2(n1227), .ZN(n1060) );
NAND2_X1 U929 ( .A1(n1229), .A2(n1226), .ZN(n1227) );
INV_X1 U930 ( .A(G237), .ZN(n1229) );
NAND2_X1 U931 ( .A1(KEYINPUT40), .A2(n1059), .ZN(n1228) );
AND3_X1 U932 ( .A1(n1230), .A2(n1231), .A3(n1226), .ZN(n1059) );
OR2_X1 U933 ( .A1(n1152), .A2(n1232), .ZN(n1231) );
NAND2_X1 U934 ( .A1(n1232), .A2(n1233), .ZN(n1230) );
XOR2_X1 U935 ( .A(n1152), .B(KEYINPUT2), .Z(n1233) );
XOR2_X1 U936 ( .A(n1112), .B(n1234), .Z(n1152) );
XNOR2_X1 U937 ( .A(n1235), .B(KEYINPUT16), .ZN(n1234) );
NAND2_X1 U938 ( .A1(KEYINPUT35), .A2(n1236), .ZN(n1235) );
XNOR2_X1 U939 ( .A(n1237), .B(n1113), .ZN(n1236) );
XNOR2_X1 U940 ( .A(n1238), .B(n1239), .ZN(n1113) );
XNOR2_X1 U941 ( .A(G101), .B(G107), .ZN(n1238) );
NAND2_X1 U942 ( .A1(KEYINPUT38), .A2(n1111), .ZN(n1237) );
XOR2_X1 U943 ( .A(G113), .B(n1240), .Z(n1111) );
XOR2_X1 U944 ( .A(n1241), .B(G122), .Z(n1112) );
XNOR2_X1 U945 ( .A(n1242), .B(KEYINPUT9), .ZN(n1232) );
NAND2_X1 U946 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
NAND2_X1 U947 ( .A1(KEYINPUT63), .A2(n1245), .ZN(n1244) );
XOR2_X1 U948 ( .A(n1246), .B(n1182), .Z(n1243) );
AND2_X1 U949 ( .A1(G224), .A2(n1073), .ZN(n1182) );
OR2_X1 U950 ( .A1(n1245), .A2(KEYINPUT63), .ZN(n1246) );
XNOR2_X1 U951 ( .A(G125), .B(n1181), .ZN(n1245) );
INV_X1 U952 ( .A(n1042), .ZN(n1199) );
XNOR2_X1 U953 ( .A(n1247), .B(n1119), .ZN(n1042) );
NAND2_X1 U954 ( .A1(G217), .A2(n1248), .ZN(n1119) );
OR2_X1 U955 ( .A1(n1118), .A2(G902), .ZN(n1247) );
XNOR2_X1 U956 ( .A(n1249), .B(n1250), .ZN(n1118) );
XOR2_X1 U957 ( .A(n1251), .B(n1252), .Z(n1250) );
XOR2_X1 U958 ( .A(n1253), .B(KEYINPUT11), .Z(n1252) );
NAND2_X1 U959 ( .A1(n1254), .A2(G221), .ZN(n1253) );
NAND2_X1 U960 ( .A1(KEYINPUT12), .A2(n1098), .ZN(n1251) );
INV_X1 U961 ( .A(G137), .ZN(n1098) );
XOR2_X1 U962 ( .A(n1147), .B(n1255), .Z(n1249) );
XNOR2_X1 U963 ( .A(n1256), .B(n1257), .ZN(n1255) );
NOR2_X1 U964 ( .A1(G119), .A2(KEYINPUT24), .ZN(n1257) );
NAND2_X1 U965 ( .A1(KEYINPUT31), .A2(n1258), .ZN(n1256) );
XOR2_X1 U966 ( .A(G140), .B(n1259), .Z(n1258) );
NOR2_X1 U967 ( .A1(G125), .A2(KEYINPUT36), .ZN(n1259) );
XOR2_X1 U968 ( .A(n1241), .B(n1260), .Z(n1147) );
INV_X1 U969 ( .A(G110), .ZN(n1241) );
INV_X1 U970 ( .A(n1027), .ZN(n1190) );
NAND2_X1 U971 ( .A1(n1206), .A2(n1207), .ZN(n1027) );
INV_X1 U972 ( .A(n1187), .ZN(n1207) );
XNOR2_X1 U973 ( .A(n1069), .B(n1261), .ZN(n1187) );
NOR2_X1 U974 ( .A1(G478), .A2(KEYINPUT57), .ZN(n1261) );
NOR2_X1 U975 ( .A1(n1124), .A2(G902), .ZN(n1069) );
XNOR2_X1 U976 ( .A(n1262), .B(n1263), .ZN(n1124) );
XOR2_X1 U977 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U978 ( .A(G107), .B(n1266), .Z(n1265) );
NOR3_X1 U979 ( .A1(n1267), .A2(KEYINPUT45), .A3(n1268), .ZN(n1266) );
NOR2_X1 U980 ( .A1(G122), .A2(n1211), .ZN(n1268) );
XOR2_X1 U981 ( .A(KEYINPUT19), .B(n1269), .Z(n1267) );
NOR2_X1 U982 ( .A1(G116), .A2(n1270), .ZN(n1269) );
XOR2_X1 U983 ( .A(KEYINPUT47), .B(G122), .Z(n1270) );
AND2_X1 U984 ( .A1(n1254), .A2(G217), .ZN(n1264) );
AND2_X1 U985 ( .A1(G234), .A2(n1073), .ZN(n1254) );
INV_X1 U986 ( .A(G953), .ZN(n1073) );
XOR2_X1 U987 ( .A(n1271), .B(n1272), .Z(n1262) );
XOR2_X1 U988 ( .A(G143), .B(G134), .Z(n1272) );
INV_X1 U989 ( .A(G128), .ZN(n1271) );
XOR2_X1 U990 ( .A(n1273), .B(G475), .Z(n1206) );
NAND2_X1 U991 ( .A1(n1128), .A2(n1226), .ZN(n1273) );
XNOR2_X1 U992 ( .A(n1274), .B(n1275), .ZN(n1128) );
XOR2_X1 U993 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U994 ( .A(n1278), .B(n1279), .Z(n1277) );
NOR2_X1 U995 ( .A1(KEYINPUT33), .A2(n1239), .ZN(n1279) );
NOR2_X1 U996 ( .A1(n1280), .A2(n1281), .ZN(n1278) );
XOR2_X1 U997 ( .A(n1282), .B(KEYINPUT17), .Z(n1281) );
NAND2_X1 U998 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NOR2_X1 U999 ( .A1(n1283), .A2(n1284), .ZN(n1280) );
XOR2_X1 U1000 ( .A(KEYINPUT21), .B(G131), .Z(n1284) );
XOR2_X1 U1001 ( .A(n1285), .B(G143), .Z(n1283) );
NAND2_X1 U1002 ( .A1(G214), .A2(n1286), .ZN(n1285) );
NOR2_X1 U1003 ( .A1(KEYINPUT3), .A2(n1086), .ZN(n1276) );
XNOR2_X1 U1004 ( .A(G125), .B(G140), .ZN(n1086) );
XOR2_X1 U1005 ( .A(n1213), .B(n1287), .Z(n1274) );
XOR2_X1 U1006 ( .A(G146), .B(G122), .Z(n1287) );
AND2_X1 U1007 ( .A1(n1049), .A2(n1050), .ZN(n1010) );
NAND2_X1 U1008 ( .A1(G221), .A2(n1248), .ZN(n1050) );
NAND2_X1 U1009 ( .A1(G234), .A2(n1226), .ZN(n1248) );
XNOR2_X1 U1010 ( .A(n1288), .B(G469), .ZN(n1049) );
NAND2_X1 U1011 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XOR2_X1 U1012 ( .A(n1291), .B(n1292), .Z(n1290) );
XOR2_X1 U1013 ( .A(n1293), .B(n1148), .Z(n1292) );
XOR2_X1 U1014 ( .A(n1294), .B(n1295), .Z(n1148) );
XOR2_X1 U1015 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U1016 ( .A(G140), .B(G101), .Z(n1297) );
NOR2_X1 U1017 ( .A1(G953), .A2(n1074), .ZN(n1296) );
INV_X1 U1018 ( .A(G227), .ZN(n1074) );
XOR2_X1 U1019 ( .A(n1298), .B(n1299), .Z(n1294) );
XOR2_X1 U1020 ( .A(n1300), .B(n1239), .Z(n1298) );
XOR2_X1 U1021 ( .A(G104), .B(KEYINPUT42), .Z(n1239) );
NAND2_X1 U1022 ( .A1(KEYINPUT62), .A2(G107), .ZN(n1300) );
NAND2_X1 U1023 ( .A1(KEYINPUT56), .A2(n1091), .ZN(n1293) );
XOR2_X1 U1024 ( .A(n1149), .B(n1260), .Z(n1091) );
NAND2_X1 U1025 ( .A1(KEYINPUT8), .A2(n1185), .ZN(n1149) );
INV_X1 U1026 ( .A(G143), .ZN(n1185) );
XOR2_X1 U1027 ( .A(KEYINPUT4), .B(G110), .Z(n1291) );
XOR2_X1 U1028 ( .A(n1226), .B(KEYINPUT14), .Z(n1289) );
XOR2_X1 U1029 ( .A(n1301), .B(G472), .Z(n1201) );
NAND2_X1 U1030 ( .A1(KEYINPUT60), .A2(n1061), .ZN(n1301) );
AND2_X1 U1031 ( .A1(n1302), .A2(n1226), .ZN(n1061) );
INV_X1 U1032 ( .A(G902), .ZN(n1226) );
XOR2_X1 U1033 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U1034 ( .A(KEYINPUT34), .B(n1140), .Z(n1304) );
AND2_X1 U1035 ( .A1(n1305), .A2(n1306), .ZN(n1140) );
NAND2_X1 U1036 ( .A1(n1240), .A2(n1213), .ZN(n1306) );
XOR2_X1 U1037 ( .A(n1307), .B(KEYINPUT7), .Z(n1305) );
OR2_X1 U1038 ( .A1(n1213), .A2(n1240), .ZN(n1307) );
XOR2_X1 U1039 ( .A(G119), .B(n1211), .Z(n1240) );
INV_X1 U1040 ( .A(G116), .ZN(n1211) );
INV_X1 U1041 ( .A(G113), .ZN(n1213) );
XOR2_X1 U1042 ( .A(n1308), .B(n1143), .Z(n1303) );
XNOR2_X1 U1043 ( .A(n1309), .B(G101), .ZN(n1143) );
NAND2_X1 U1044 ( .A1(G210), .A2(n1286), .ZN(n1309) );
NOR2_X1 U1045 ( .A1(G953), .A2(G237), .ZN(n1286) );
NAND2_X1 U1046 ( .A1(n1310), .A2(n1311), .ZN(n1308) );
NAND3_X1 U1047 ( .A1(n1299), .A2(n1181), .A3(n1312), .ZN(n1311) );
INV_X1 U1048 ( .A(KEYINPUT13), .ZN(n1312) );
INV_X1 U1049 ( .A(n1313), .ZN(n1299) );
NAND2_X1 U1050 ( .A1(n1142), .A2(KEYINPUT13), .ZN(n1310) );
XNOR2_X1 U1051 ( .A(n1313), .B(n1181), .ZN(n1142) );
XOR2_X1 U1052 ( .A(G143), .B(n1260), .Z(n1181) );
XOR2_X1 U1053 ( .A(G128), .B(G146), .Z(n1260) );
XOR2_X1 U1054 ( .A(n1191), .B(n1314), .Z(n1313) );
XOR2_X1 U1055 ( .A(G137), .B(G134), .Z(n1314) );
INV_X1 U1056 ( .A(G131), .ZN(n1191) );
endmodule


