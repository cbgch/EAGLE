//Key = 0111101111010111011011110101011001101110100110010011010001110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372;

XNOR2_X1 U761 ( .A(G107), .B(n1051), .ZN(G9) );
NOR2_X1 U762 ( .A1(n1052), .A2(n1053), .ZN(G75) );
XOR2_X1 U763 ( .A(KEYINPUT41), .B(n1054), .Z(n1053) );
NOR3_X1 U764 ( .A1(n1055), .A2(G953), .A3(G952), .ZN(n1054) );
NOR4_X1 U765 ( .A1(n1056), .A2(n1057), .A3(G953), .A4(n1058), .ZN(n1052) );
NOR4_X1 U766 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1058) );
NOR2_X1 U767 ( .A1(n1063), .A2(n1064), .ZN(n1059) );
NOR2_X1 U768 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1063) );
XOR2_X1 U770 ( .A(n1066), .B(KEYINPUT48), .Z(n1067) );
NOR3_X1 U771 ( .A1(n1066), .A2(n1069), .A3(n1070), .ZN(n1057) );
NOR2_X1 U772 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR2_X1 U773 ( .A1(n1073), .A2(n1060), .ZN(n1072) );
NOR2_X1 U774 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U775 ( .A1(n1076), .A2(n1062), .ZN(n1075) );
NOR2_X1 U776 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XNOR2_X1 U777 ( .A(n1079), .B(KEYINPUT15), .ZN(n1078) );
NOR2_X1 U778 ( .A1(n1080), .A2(n1061), .ZN(n1074) );
NOR2_X1 U779 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U780 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NOR3_X1 U781 ( .A1(n1062), .A2(n1085), .A3(n1061), .ZN(n1071) );
NOR2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NAND2_X1 U784 ( .A1(KEYINPUT25), .A2(n1090), .ZN(n1066) );
NAND3_X1 U785 ( .A1(n1091), .A2(G952), .A3(n1092), .ZN(n1056) );
XNOR2_X1 U786 ( .A(n1055), .B(KEYINPUT63), .ZN(n1092) );
AND4_X1 U787 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1055) );
NOR4_X1 U788 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
XOR2_X1 U789 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U790 ( .A1(G478), .A2(KEYINPUT26), .ZN(n1102) );
INV_X1 U791 ( .A(n1103), .ZN(n1099) );
NOR3_X1 U792 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1095) );
NOR2_X1 U793 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U794 ( .A(G472), .B(KEYINPUT5), .ZN(n1108) );
NOR2_X1 U795 ( .A1(G472), .A2(n1109), .ZN(n1105) );
XOR2_X1 U796 ( .A(n1110), .B(n1111), .Z(n1104) );
NOR2_X1 U797 ( .A1(KEYINPUT39), .A2(n1112), .ZN(n1111) );
XNOR2_X1 U798 ( .A(n1113), .B(n1114), .ZN(n1093) );
NAND2_X1 U799 ( .A1(KEYINPUT3), .A2(n1115), .ZN(n1113) );
NAND3_X1 U800 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(G72) );
XOR2_X1 U801 ( .A(n1119), .B(KEYINPUT19), .Z(n1118) );
NAND2_X1 U802 ( .A1(G953), .A2(n1120), .ZN(n1119) );
NAND2_X1 U803 ( .A1(G900), .A2(n1121), .ZN(n1120) );
OR2_X1 U804 ( .A1(n1122), .A2(G227), .ZN(n1121) );
NAND2_X1 U805 ( .A1(n1123), .A2(n1124), .ZN(n1117) );
XNOR2_X1 U806 ( .A(n1125), .B(n1122), .ZN(n1123) );
NAND4_X1 U807 ( .A1(G227), .A2(n1122), .A3(G900), .A4(G953), .ZN(n1116) );
XNOR2_X1 U808 ( .A(n1126), .B(n1127), .ZN(n1122) );
XNOR2_X1 U809 ( .A(n1128), .B(KEYINPUT0), .ZN(n1126) );
NAND2_X1 U810 ( .A1(n1129), .A2(n1130), .ZN(G69) );
NAND2_X1 U811 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U812 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
NAND2_X1 U813 ( .A1(n1135), .A2(n1134), .ZN(n1129) );
NAND2_X1 U814 ( .A1(G953), .A2(n1136), .ZN(n1134) );
INV_X1 U815 ( .A(n1132), .ZN(n1135) );
NAND2_X1 U816 ( .A1(KEYINPUT37), .A2(n1137), .ZN(n1132) );
XOR2_X1 U817 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U818 ( .A1(n1140), .A2(n1133), .ZN(n1139) );
INV_X1 U819 ( .A(n1141), .ZN(n1133) );
XOR2_X1 U820 ( .A(n1142), .B(n1143), .Z(n1140) );
NOR3_X1 U821 ( .A1(n1144), .A2(KEYINPUT12), .A3(n1145), .ZN(n1142) );
NOR2_X1 U822 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U823 ( .A(n1148), .B(KEYINPUT59), .Z(n1144) );
NAND2_X1 U824 ( .A1(n1146), .A2(n1147), .ZN(n1148) );
INV_X1 U825 ( .A(n1149), .ZN(n1146) );
NAND2_X1 U826 ( .A1(n1150), .A2(n1124), .ZN(n1138) );
NAND2_X1 U827 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U828 ( .A(n1153), .B(KEYINPUT55), .Z(n1151) );
NOR2_X1 U829 ( .A1(n1154), .A2(n1155), .ZN(G66) );
XOR2_X1 U830 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U831 ( .A1(KEYINPUT33), .A2(n1158), .ZN(n1157) );
NAND2_X1 U832 ( .A1(n1159), .A2(n1160), .ZN(n1156) );
INV_X1 U833 ( .A(n1112), .ZN(n1160) );
NOR2_X1 U834 ( .A1(n1154), .A2(n1161), .ZN(G63) );
XOR2_X1 U835 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U836 ( .A1(n1159), .A2(G478), .ZN(n1162) );
NOR2_X1 U837 ( .A1(n1154), .A2(n1164), .ZN(G60) );
XNOR2_X1 U838 ( .A(n1165), .B(n1166), .ZN(n1164) );
NAND2_X1 U839 ( .A1(n1159), .A2(G475), .ZN(n1165) );
XOR2_X1 U840 ( .A(n1153), .B(n1167), .Z(G6) );
NAND2_X1 U841 ( .A1(KEYINPUT2), .A2(G104), .ZN(n1167) );
NOR2_X1 U842 ( .A1(n1154), .A2(n1168), .ZN(G57) );
XOR2_X1 U843 ( .A(n1169), .B(n1170), .Z(n1168) );
XNOR2_X1 U844 ( .A(n1171), .B(n1172), .ZN(n1170) );
XOR2_X1 U845 ( .A(n1173), .B(n1174), .Z(n1169) );
XNOR2_X1 U846 ( .A(n1175), .B(KEYINPUT18), .ZN(n1174) );
NAND2_X1 U847 ( .A1(KEYINPUT43), .A2(n1176), .ZN(n1175) );
NAND2_X1 U848 ( .A1(n1159), .A2(G472), .ZN(n1173) );
NOR2_X1 U849 ( .A1(n1154), .A2(n1177), .ZN(G54) );
XOR2_X1 U850 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U851 ( .A(n1180), .B(n1181), .Z(n1179) );
NAND2_X1 U852 ( .A1(n1159), .A2(G469), .ZN(n1181) );
NAND2_X1 U853 ( .A1(n1182), .A2(n1183), .ZN(n1180) );
NAND2_X1 U854 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NAND2_X1 U855 ( .A1(KEYINPUT27), .A2(n1186), .ZN(n1185) );
NAND2_X1 U856 ( .A1(KEYINPUT62), .A2(n1187), .ZN(n1186) );
INV_X1 U857 ( .A(n1188), .ZN(n1187) );
NAND2_X1 U858 ( .A1(n1188), .A2(n1189), .ZN(n1182) );
NAND2_X1 U859 ( .A1(KEYINPUT62), .A2(n1190), .ZN(n1189) );
NAND2_X1 U860 ( .A1(n1191), .A2(KEYINPUT27), .ZN(n1190) );
INV_X1 U861 ( .A(n1184), .ZN(n1191) );
XNOR2_X1 U862 ( .A(n1192), .B(n1193), .ZN(n1184) );
NAND2_X1 U863 ( .A1(KEYINPUT50), .A2(n1194), .ZN(n1178) );
NOR2_X1 U864 ( .A1(n1154), .A2(n1195), .ZN(G51) );
XOR2_X1 U865 ( .A(n1196), .B(n1197), .Z(n1195) );
XNOR2_X1 U866 ( .A(n1198), .B(n1199), .ZN(n1197) );
NOR4_X1 U867 ( .A1(n1200), .A2(n1201), .A3(KEYINPUT56), .A4(n1202), .ZN(n1199) );
NOR2_X1 U868 ( .A1(KEYINPUT34), .A2(n1203), .ZN(n1201) );
NOR2_X1 U869 ( .A1(G902), .A2(n1091), .ZN(n1203) );
NOR2_X1 U870 ( .A1(n1159), .A2(n1204), .ZN(n1200) );
INV_X1 U871 ( .A(KEYINPUT34), .ZN(n1204) );
NOR2_X1 U872 ( .A1(n1205), .A2(n1091), .ZN(n1159) );
AND3_X1 U873 ( .A1(n1152), .A2(n1153), .A3(n1125), .ZN(n1091) );
AND4_X1 U874 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1125) );
NOR4_X1 U875 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1209) );
NAND2_X1 U876 ( .A1(n1214), .A2(n1215), .ZN(n1208) );
NAND2_X1 U877 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND3_X1 U878 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1217) );
NAND2_X1 U879 ( .A1(KEYINPUT1), .A2(n1221), .ZN(n1219) );
NAND2_X1 U880 ( .A1(n1222), .A2(n1223), .ZN(n1218) );
INV_X1 U881 ( .A(KEYINPUT1), .ZN(n1223) );
NAND2_X1 U882 ( .A1(n1224), .A2(n1225), .ZN(n1222) );
XNOR2_X1 U883 ( .A(KEYINPUT22), .B(n1226), .ZN(n1216) );
NAND3_X1 U884 ( .A1(n1227), .A2(n1228), .A3(n1079), .ZN(n1153) );
AND4_X1 U885 ( .A1(n1051), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1152) );
NOR3_X1 U886 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1231) );
NOR3_X1 U887 ( .A1(n1235), .A2(n1236), .A3(n1065), .ZN(n1234) );
XNOR2_X1 U888 ( .A(KEYINPUT40), .B(n1061), .ZN(n1235) );
NOR2_X1 U889 ( .A1(n1237), .A2(n1238), .ZN(n1232) );
NOR2_X1 U890 ( .A1(n1239), .A2(n1220), .ZN(n1237) );
NAND3_X1 U891 ( .A1(n1077), .A2(n1228), .A3(n1227), .ZN(n1051) );
INV_X1 U892 ( .A(n1236), .ZN(n1227) );
INV_X1 U893 ( .A(n1070), .ZN(n1228) );
NAND2_X1 U894 ( .A1(n1240), .A2(KEYINPUT20), .ZN(n1198) );
XNOR2_X1 U895 ( .A(G125), .B(n1241), .ZN(n1240) );
NOR2_X1 U896 ( .A1(KEYINPUT35), .A2(n1176), .ZN(n1241) );
NOR2_X1 U897 ( .A1(n1242), .A2(G952), .ZN(n1154) );
XNOR2_X1 U898 ( .A(KEYINPUT49), .B(G953), .ZN(n1242) );
XNOR2_X1 U899 ( .A(G146), .B(n1206), .ZN(G48) );
NAND2_X1 U900 ( .A1(n1243), .A2(n1079), .ZN(n1206) );
NAND2_X1 U901 ( .A1(n1244), .A2(n1245), .ZN(G45) );
OR2_X1 U902 ( .A1(n1246), .A2(G143), .ZN(n1245) );
NAND2_X1 U903 ( .A1(G143), .A2(n1247), .ZN(n1244) );
NAND2_X1 U904 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
OR2_X1 U905 ( .A1(n1207), .A2(KEYINPUT51), .ZN(n1249) );
NAND2_X1 U906 ( .A1(KEYINPUT51), .A2(n1246), .ZN(n1248) );
NAND2_X1 U907 ( .A1(KEYINPUT21), .A2(n1250), .ZN(n1246) );
INV_X1 U908 ( .A(n1207), .ZN(n1250) );
NAND3_X1 U909 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1207) );
NOR3_X1 U910 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1253) );
XOR2_X1 U911 ( .A(G140), .B(n1213), .Z(G42) );
NOR4_X1 U912 ( .A1(n1062), .A2(n1221), .A3(n1065), .A4(n1257), .ZN(n1213) );
NAND2_X1 U913 ( .A1(n1258), .A2(n1259), .ZN(G39) );
NAND2_X1 U914 ( .A1(n1212), .A2(n1260), .ZN(n1259) );
XOR2_X1 U915 ( .A(KEYINPUT29), .B(n1261), .Z(n1258) );
NOR2_X1 U916 ( .A1(n1212), .A2(n1260), .ZN(n1261) );
AND3_X1 U917 ( .A1(n1239), .A2(n1252), .A3(n1214), .ZN(n1212) );
XNOR2_X1 U918 ( .A(G134), .B(n1262), .ZN(G36) );
NOR2_X1 U919 ( .A1(n1263), .A2(KEYINPUT60), .ZN(n1262) );
NOR3_X1 U920 ( .A1(n1264), .A2(n1221), .A3(n1062), .ZN(n1263) );
XOR2_X1 U921 ( .A(G131), .B(n1265), .Z(G33) );
NOR2_X1 U922 ( .A1(n1062), .A2(n1226), .ZN(n1265) );
NAND3_X1 U923 ( .A1(n1252), .A2(n1079), .A3(n1251), .ZN(n1226) );
INV_X1 U924 ( .A(n1221), .ZN(n1252) );
INV_X1 U925 ( .A(n1214), .ZN(n1062) );
NOR2_X1 U926 ( .A1(n1083), .A2(n1098), .ZN(n1214) );
INV_X1 U927 ( .A(n1084), .ZN(n1098) );
XOR2_X1 U928 ( .A(n1211), .B(n1266), .Z(G30) );
NOR2_X1 U929 ( .A1(KEYINPUT54), .A2(n1267), .ZN(n1266) );
AND2_X1 U930 ( .A1(n1243), .A2(n1077), .ZN(n1211) );
NOR4_X1 U931 ( .A1(n1221), .A2(n1254), .A3(n1268), .A4(n1269), .ZN(n1243) );
NAND2_X1 U932 ( .A1(n1087), .A2(n1224), .ZN(n1221) );
XNOR2_X1 U933 ( .A(n1270), .B(n1233), .ZN(G3) );
NOR3_X1 U934 ( .A1(n1061), .A2(n1236), .A3(n1068), .ZN(n1233) );
XOR2_X1 U935 ( .A(G125), .B(n1210), .Z(G27) );
AND4_X1 U936 ( .A1(n1082), .A2(n1224), .A3(n1079), .A4(n1271), .ZN(n1210) );
NOR2_X1 U937 ( .A1(n1060), .A2(n1065), .ZN(n1271) );
INV_X1 U938 ( .A(n1094), .ZN(n1060) );
INV_X1 U939 ( .A(n1257), .ZN(n1079) );
NAND2_X1 U940 ( .A1(n1272), .A2(n1273), .ZN(n1224) );
NAND4_X1 U941 ( .A1(G902), .A2(G953), .A3(n1090), .A4(n1274), .ZN(n1273) );
INV_X1 U942 ( .A(G900), .ZN(n1274) );
XNOR2_X1 U943 ( .A(G122), .B(n1230), .ZN(G24) );
OR4_X1 U944 ( .A1(n1238), .A2(n1070), .A3(n1256), .A4(n1255), .ZN(n1230) );
NAND2_X1 U945 ( .A1(n1269), .A2(n1268), .ZN(n1070) );
NAND3_X1 U946 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(G21) );
NAND2_X1 U947 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NAND2_X1 U948 ( .A1(n1280), .A2(n1281), .ZN(n1276) );
INV_X1 U949 ( .A(KEYINPUT38), .ZN(n1281) );
NAND2_X1 U950 ( .A1(n1282), .A2(G119), .ZN(n1280) );
XNOR2_X1 U951 ( .A(n1278), .B(KEYINPUT32), .ZN(n1282) );
NAND2_X1 U952 ( .A1(KEYINPUT38), .A2(n1283), .ZN(n1275) );
NAND2_X1 U953 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
OR3_X1 U954 ( .A1(n1279), .A2(n1278), .A3(KEYINPUT32), .ZN(n1285) );
NAND2_X1 U955 ( .A1(KEYINPUT32), .A2(n1278), .ZN(n1284) );
AND3_X1 U956 ( .A1(n1286), .A2(n1287), .A3(n1239), .ZN(n1278) );
NOR3_X1 U957 ( .A1(n1268), .A2(n1269), .A3(n1061), .ZN(n1239) );
INV_X1 U958 ( .A(n1288), .ZN(n1269) );
NAND2_X1 U959 ( .A1(KEYINPUT6), .A2(n1238), .ZN(n1287) );
NAND2_X1 U960 ( .A1(n1289), .A2(n1290), .ZN(n1286) );
INV_X1 U961 ( .A(KEYINPUT6), .ZN(n1290) );
NAND3_X1 U962 ( .A1(n1254), .A2(n1291), .A3(n1094), .ZN(n1289) );
XNOR2_X1 U963 ( .A(G116), .B(n1292), .ZN(G18) );
NAND4_X1 U964 ( .A1(n1220), .A2(n1094), .A3(n1082), .A4(n1293), .ZN(n1292) );
XNOR2_X1 U965 ( .A(KEYINPUT14), .B(n1291), .ZN(n1293) );
INV_X1 U966 ( .A(n1264), .ZN(n1220) );
NAND2_X1 U967 ( .A1(n1251), .A2(n1077), .ZN(n1264) );
NOR2_X1 U968 ( .A1(n1294), .A2(n1256), .ZN(n1077) );
INV_X1 U969 ( .A(n1068), .ZN(n1251) );
XNOR2_X1 U970 ( .A(G113), .B(n1229), .ZN(G15) );
OR3_X1 U971 ( .A1(n1068), .A2(n1257), .A3(n1238), .ZN(n1229) );
NAND3_X1 U972 ( .A1(n1082), .A2(n1291), .A3(n1094), .ZN(n1238) );
NOR2_X1 U973 ( .A1(n1088), .A2(n1295), .ZN(n1094) );
INV_X1 U974 ( .A(n1089), .ZN(n1295) );
NAND2_X1 U975 ( .A1(n1256), .A2(n1294), .ZN(n1257) );
NAND2_X1 U976 ( .A1(n1268), .A2(n1288), .ZN(n1068) );
XOR2_X1 U977 ( .A(G110), .B(n1296), .Z(G12) );
NOR3_X1 U978 ( .A1(n1297), .A2(n1236), .A3(n1061), .ZN(n1296) );
NAND2_X1 U979 ( .A1(n1256), .A2(n1255), .ZN(n1061) );
INV_X1 U980 ( .A(n1294), .ZN(n1255) );
NAND3_X1 U981 ( .A1(n1298), .A2(n1299), .A3(n1103), .ZN(n1294) );
NAND2_X1 U982 ( .A1(G475), .A2(n1300), .ZN(n1103) );
OR2_X1 U983 ( .A1(n1166), .A2(G902), .ZN(n1300) );
NAND2_X1 U984 ( .A1(n1097), .A2(n1301), .ZN(n1299) );
INV_X1 U985 ( .A(KEYINPUT42), .ZN(n1301) );
NOR3_X1 U986 ( .A1(G475), .A2(G902), .A3(n1166), .ZN(n1097) );
XOR2_X1 U987 ( .A(n1302), .B(n1303), .Z(n1166) );
XOR2_X1 U988 ( .A(G104), .B(n1304), .Z(n1303) );
XOR2_X1 U989 ( .A(G146), .B(G122), .Z(n1304) );
XOR2_X1 U990 ( .A(n1305), .B(n1128), .Z(n1302) );
XOR2_X1 U991 ( .A(G125), .B(n1306), .Z(n1128) );
XOR2_X1 U992 ( .A(n1307), .B(n1308), .Z(n1305) );
NOR2_X1 U993 ( .A1(KEYINPUT16), .A2(n1309), .ZN(n1308) );
INV_X1 U994 ( .A(G113), .ZN(n1309) );
NAND2_X1 U995 ( .A1(n1310), .A2(n1311), .ZN(n1307) );
NAND2_X1 U996 ( .A1(n1312), .A2(G131), .ZN(n1311) );
XOR2_X1 U997 ( .A(n1313), .B(KEYINPUT46), .Z(n1310) );
OR2_X1 U998 ( .A1(n1312), .A2(G131), .ZN(n1313) );
XOR2_X1 U999 ( .A(n1314), .B(G143), .Z(n1312) );
NAND2_X1 U1000 ( .A1(n1315), .A2(G214), .ZN(n1314) );
NAND2_X1 U1001 ( .A1(KEYINPUT42), .A2(G475), .ZN(n1298) );
XOR2_X1 U1002 ( .A(n1101), .B(G478), .Z(n1256) );
NAND2_X1 U1003 ( .A1(n1163), .A2(n1316), .ZN(n1101) );
XNOR2_X1 U1004 ( .A(KEYINPUT58), .B(n1205), .ZN(n1316) );
XOR2_X1 U1005 ( .A(n1317), .B(n1318), .Z(n1163) );
XNOR2_X1 U1006 ( .A(n1319), .B(n1320), .ZN(n1318) );
XOR2_X1 U1007 ( .A(n1321), .B(n1322), .Z(n1320) );
AND3_X1 U1008 ( .A1(n1323), .A2(G234), .A3(G217), .ZN(n1322) );
XNOR2_X1 U1009 ( .A(KEYINPUT31), .B(G953), .ZN(n1323) );
NAND2_X1 U1010 ( .A1(KEYINPUT11), .A2(n1324), .ZN(n1321) );
INV_X1 U1011 ( .A(G134), .ZN(n1324) );
XOR2_X1 U1012 ( .A(n1325), .B(n1326), .Z(n1317) );
XOR2_X1 U1013 ( .A(KEYINPUT61), .B(G122), .Z(n1326) );
XNOR2_X1 U1014 ( .A(G107), .B(G116), .ZN(n1325) );
NAND3_X1 U1015 ( .A1(n1082), .A2(n1291), .A3(n1087), .ZN(n1236) );
INV_X1 U1016 ( .A(n1225), .ZN(n1087) );
NAND2_X1 U1017 ( .A1(n1088), .A2(n1089), .ZN(n1225) );
NAND2_X1 U1018 ( .A1(G221), .A2(n1327), .ZN(n1089) );
XNOR2_X1 U1019 ( .A(n1328), .B(G469), .ZN(n1088) );
NAND2_X1 U1020 ( .A1(n1329), .A2(n1205), .ZN(n1328) );
XOR2_X1 U1021 ( .A(n1330), .B(n1331), .Z(n1329) );
XOR2_X1 U1022 ( .A(n1127), .B(n1194), .Z(n1331) );
XOR2_X1 U1023 ( .A(n1306), .B(n1332), .Z(n1194) );
XOR2_X1 U1024 ( .A(G110), .B(n1333), .Z(n1332) );
AND2_X1 U1025 ( .A1(n1124), .A2(G227), .ZN(n1333) );
XNOR2_X1 U1026 ( .A(n1334), .B(n1193), .ZN(n1127) );
XOR2_X1 U1027 ( .A(n1176), .B(KEYINPUT17), .Z(n1193) );
XNOR2_X1 U1028 ( .A(KEYINPUT23), .B(n1335), .ZN(n1330) );
NAND2_X1 U1029 ( .A1(KEYINPUT36), .A2(n1192), .ZN(n1335) );
XOR2_X1 U1030 ( .A(n1336), .B(n1337), .Z(n1192) );
NAND2_X1 U1031 ( .A1(KEYINPUT8), .A2(n1270), .ZN(n1336) );
INV_X1 U1032 ( .A(G101), .ZN(n1270) );
NAND2_X1 U1033 ( .A1(n1272), .A2(n1338), .ZN(n1291) );
NAND3_X1 U1034 ( .A1(n1141), .A2(n1090), .A3(n1339), .ZN(n1338) );
XNOR2_X1 U1035 ( .A(G902), .B(KEYINPUT53), .ZN(n1339) );
NOR2_X1 U1036 ( .A1(G898), .A2(n1124), .ZN(n1141) );
NAND3_X1 U1037 ( .A1(n1090), .A2(n1124), .A3(n1340), .ZN(n1272) );
XNOR2_X1 U1038 ( .A(G952), .B(KEYINPUT4), .ZN(n1340) );
NAND2_X1 U1039 ( .A1(G237), .A2(G234), .ZN(n1090) );
INV_X1 U1040 ( .A(n1254), .ZN(n1082) );
NAND2_X1 U1041 ( .A1(n1083), .A2(n1084), .ZN(n1254) );
NAND2_X1 U1042 ( .A1(G214), .A2(n1341), .ZN(n1084) );
XOR2_X1 U1043 ( .A(n1114), .B(n1342), .Z(n1083) );
NOR2_X1 U1044 ( .A1(n1115), .A2(KEYINPUT52), .ZN(n1342) );
INV_X1 U1045 ( .A(n1202), .ZN(n1115) );
NAND2_X1 U1046 ( .A1(G210), .A2(n1341), .ZN(n1202) );
NAND2_X1 U1047 ( .A1(n1343), .A2(n1205), .ZN(n1341) );
INV_X1 U1048 ( .A(G237), .ZN(n1343) );
NAND2_X1 U1049 ( .A1(n1344), .A2(n1205), .ZN(n1114) );
XOR2_X1 U1050 ( .A(n1345), .B(n1346), .Z(n1344) );
XOR2_X1 U1051 ( .A(n1176), .B(n1196), .Z(n1346) );
XNOR2_X1 U1052 ( .A(n1347), .B(n1348), .ZN(n1196) );
XOR2_X1 U1053 ( .A(n1349), .B(n1350), .Z(n1348) );
NOR2_X1 U1054 ( .A1(KEYINPUT24), .A2(n1149), .ZN(n1350) );
XOR2_X1 U1055 ( .A(G113), .B(n1351), .Z(n1149) );
NOR2_X1 U1056 ( .A1(G953), .A2(n1136), .ZN(n1349) );
INV_X1 U1057 ( .A(G224), .ZN(n1136) );
XNOR2_X1 U1058 ( .A(n1143), .B(n1147), .ZN(n1347) );
XNOR2_X1 U1059 ( .A(n1352), .B(n1337), .ZN(n1147) );
XOR2_X1 U1060 ( .A(G104), .B(G107), .Z(n1337) );
XNOR2_X1 U1061 ( .A(G101), .B(KEYINPUT13), .ZN(n1352) );
XOR2_X1 U1062 ( .A(G110), .B(n1353), .Z(n1143) );
NOR2_X1 U1063 ( .A1(G122), .A2(KEYINPUT45), .ZN(n1353) );
XNOR2_X1 U1064 ( .A(G125), .B(KEYINPUT10), .ZN(n1345) );
XNOR2_X1 U1065 ( .A(KEYINPUT44), .B(n1065), .ZN(n1297) );
OR2_X1 U1066 ( .A1(n1288), .A2(n1268), .ZN(n1065) );
XOR2_X1 U1067 ( .A(n1110), .B(n1112), .Z(n1268) );
NAND2_X1 U1068 ( .A1(G217), .A2(n1327), .ZN(n1112) );
NAND2_X1 U1069 ( .A1(G234), .A2(n1205), .ZN(n1327) );
NOR2_X1 U1070 ( .A1(n1158), .A2(G902), .ZN(n1110) );
XOR2_X1 U1071 ( .A(n1354), .B(n1355), .Z(n1158) );
XOR2_X1 U1072 ( .A(n1356), .B(n1357), .Z(n1355) );
XNOR2_X1 U1073 ( .A(n1267), .B(G125), .ZN(n1357) );
XNOR2_X1 U1074 ( .A(G146), .B(n1260), .ZN(n1356) );
XOR2_X1 U1075 ( .A(n1358), .B(n1359), .Z(n1354) );
XOR2_X1 U1076 ( .A(n1360), .B(n1361), .Z(n1359) );
AND3_X1 U1077 ( .A1(G221), .A2(n1124), .A3(G234), .ZN(n1361) );
INV_X1 U1078 ( .A(G953), .ZN(n1124) );
NOR2_X1 U1079 ( .A1(G110), .A2(KEYINPUT28), .ZN(n1360) );
XNOR2_X1 U1080 ( .A(n1362), .B(n1279), .ZN(n1358) );
INV_X1 U1081 ( .A(G119), .ZN(n1279) );
NAND2_X1 U1082 ( .A1(n1363), .A2(n1306), .ZN(n1362) );
XOR2_X1 U1083 ( .A(G140), .B(KEYINPUT57), .Z(n1306) );
XNOR2_X1 U1084 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n1363) );
XOR2_X1 U1085 ( .A(n1107), .B(G472), .Z(n1288) );
INV_X1 U1086 ( .A(n1109), .ZN(n1107) );
NAND2_X1 U1087 ( .A1(n1364), .A2(n1205), .ZN(n1109) );
INV_X1 U1088 ( .A(G902), .ZN(n1205) );
XNOR2_X1 U1089 ( .A(n1365), .B(n1366), .ZN(n1364) );
XOR2_X1 U1090 ( .A(n1172), .B(n1176), .Z(n1366) );
XOR2_X1 U1091 ( .A(G146), .B(n1319), .Z(n1176) );
XNOR2_X1 U1092 ( .A(n1267), .B(G143), .ZN(n1319) );
INV_X1 U1093 ( .A(G128), .ZN(n1267) );
XNOR2_X1 U1094 ( .A(n1367), .B(G101), .ZN(n1172) );
NAND2_X1 U1095 ( .A1(n1315), .A2(G210), .ZN(n1367) );
NOR2_X1 U1096 ( .A1(G953), .A2(G237), .ZN(n1315) );
INV_X1 U1097 ( .A(n1171), .ZN(n1365) );
XOR2_X1 U1098 ( .A(n1188), .B(n1368), .Z(n1171) );
XNOR2_X1 U1099 ( .A(G113), .B(n1369), .ZN(n1368) );
NAND2_X1 U1100 ( .A1(KEYINPUT47), .A2(n1351), .ZN(n1369) );
XNOR2_X1 U1101 ( .A(n1370), .B(G119), .ZN(n1351) );
INV_X1 U1102 ( .A(G116), .ZN(n1370) );
XNOR2_X1 U1103 ( .A(KEYINPUT23), .B(n1334), .ZN(n1188) );
XOR2_X1 U1104 ( .A(n1371), .B(n1372), .Z(n1334) );
XNOR2_X1 U1105 ( .A(KEYINPUT30), .B(n1260), .ZN(n1372) );
INV_X1 U1106 ( .A(G137), .ZN(n1260) );
XNOR2_X1 U1107 ( .A(G134), .B(G131), .ZN(n1371) );
endmodule


