//Key = 1000101111001001001111111101100101101001001110010010111101011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371;

XOR2_X1 U749 ( .A(n1036), .B(n1037), .Z(G9) );
NOR2_X1 U750 ( .A1(KEYINPUT29), .A2(n1038), .ZN(n1037) );
INV_X1 U751 ( .A(n1039), .ZN(n1038) );
XNOR2_X1 U752 ( .A(G107), .B(KEYINPUT26), .ZN(n1036) );
NAND4_X1 U753 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(G75) );
INV_X1 U754 ( .A(n1044), .ZN(n1043) );
NAND4_X1 U755 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1042) );
NOR4_X1 U756 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
XOR2_X1 U757 ( .A(n1053), .B(n1054), .Z(n1052) );
XNOR2_X1 U758 ( .A(KEYINPUT44), .B(n1055), .ZN(n1054) );
XNOR2_X1 U759 ( .A(n1056), .B(KEYINPUT32), .ZN(n1047) );
XOR2_X1 U760 ( .A(n1057), .B(n1058), .Z(n1045) );
NAND2_X1 U761 ( .A1(G952), .A2(n1059), .ZN(n1041) );
NAND3_X1 U762 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NAND2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NAND2_X1 U764 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND4_X1 U765 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
NAND2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NAND2_X1 U767 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U768 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U769 ( .A1(n1046), .A2(n1077), .ZN(n1071) );
NAND2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U771 ( .A1(n1049), .A2(n1080), .ZN(n1079) );
NAND3_X1 U772 ( .A1(n1046), .A2(n1081), .A3(n1073), .ZN(n1065) );
NAND2_X1 U773 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND3_X1 U774 ( .A1(n1084), .A2(n1085), .A3(n1067), .ZN(n1083) );
NAND2_X1 U775 ( .A1(n1050), .A2(n1086), .ZN(n1085) );
NAND2_X1 U776 ( .A1(n1068), .A2(n1087), .ZN(n1086) );
INV_X1 U777 ( .A(KEYINPUT10), .ZN(n1087) );
NAND4_X1 U778 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1070), .ZN(n1084) );
NAND2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U780 ( .A1(KEYINPUT10), .A2(n1068), .ZN(n1088) );
NAND2_X1 U781 ( .A1(n1068), .A2(n1093), .ZN(n1082) );
INV_X1 U782 ( .A(n1094), .ZN(n1063) );
OR2_X1 U783 ( .A1(G953), .A2(KEYINPUT4), .ZN(n1060) );
NAND2_X1 U784 ( .A1(KEYINPUT4), .A2(G953), .ZN(n1040) );
XOR2_X1 U785 ( .A(n1095), .B(n1096), .Z(G72) );
XOR2_X1 U786 ( .A(n1097), .B(n1098), .Z(n1096) );
NAND2_X1 U787 ( .A1(G953), .A2(n1099), .ZN(n1098) );
NAND2_X1 U788 ( .A1(G900), .A2(G227), .ZN(n1099) );
NAND2_X1 U789 ( .A1(n1100), .A2(n1101), .ZN(n1097) );
XOR2_X1 U790 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U791 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U792 ( .A(n1106), .B(KEYINPUT49), .Z(n1100) );
OR2_X1 U793 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U794 ( .A1(n1109), .A2(G953), .ZN(n1095) );
XOR2_X1 U795 ( .A(n1110), .B(n1111), .Z(G69) );
NOR2_X1 U796 ( .A1(n1112), .A2(G953), .ZN(n1111) );
NAND2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
NAND2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U799 ( .A1(G953), .A2(n1117), .ZN(n1116) );
INV_X1 U800 ( .A(n1118), .ZN(n1115) );
NAND3_X1 U801 ( .A1(G953), .A2(n1119), .A3(n1118), .ZN(n1113) );
NAND2_X1 U802 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
NAND2_X1 U803 ( .A1(G953), .A2(n1122), .ZN(n1121) );
XOR2_X1 U804 ( .A(n1123), .B(n1124), .Z(n1120) );
NOR2_X1 U805 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
XOR2_X1 U806 ( .A(n1127), .B(KEYINPUT36), .Z(n1126) );
NAND2_X1 U807 ( .A1(G898), .A2(G224), .ZN(n1119) );
NOR2_X1 U808 ( .A1(n1044), .A2(n1128), .ZN(G66) );
NOR3_X1 U809 ( .A1(n1057), .A2(n1129), .A3(n1130), .ZN(n1128) );
NOR3_X1 U810 ( .A1(n1131), .A2(n1058), .A3(n1132), .ZN(n1130) );
NOR2_X1 U811 ( .A1(n1133), .A2(n1134), .ZN(n1129) );
NOR2_X1 U812 ( .A1(n1062), .A2(n1058), .ZN(n1133) );
NOR2_X1 U813 ( .A1(n1044), .A2(n1135), .ZN(G63) );
XNOR2_X1 U814 ( .A(n1136), .B(n1137), .ZN(n1135) );
AND2_X1 U815 ( .A1(G478), .A2(n1138), .ZN(n1137) );
NOR2_X1 U816 ( .A1(n1044), .A2(n1139), .ZN(G60) );
NOR2_X1 U817 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U818 ( .A(n1142), .B(KEYINPUT61), .Z(n1141) );
NAND2_X1 U819 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NOR2_X1 U820 ( .A1(n1143), .A2(n1144), .ZN(n1140) );
AND2_X1 U821 ( .A1(n1138), .A2(G475), .ZN(n1144) );
INV_X1 U822 ( .A(n1145), .ZN(n1143) );
NAND2_X1 U823 ( .A1(n1146), .A2(n1147), .ZN(G6) );
OR2_X1 U824 ( .A1(n1148), .A2(G104), .ZN(n1147) );
NAND2_X1 U825 ( .A1(G104), .A2(n1149), .ZN(n1146) );
NAND2_X1 U826 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND2_X1 U827 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
INV_X1 U828 ( .A(KEYINPUT42), .ZN(n1153) );
NAND2_X1 U829 ( .A1(KEYINPUT42), .A2(n1148), .ZN(n1150) );
NAND2_X1 U830 ( .A1(KEYINPUT53), .A2(n1152), .ZN(n1148) );
NOR2_X1 U831 ( .A1(n1044), .A2(n1154), .ZN(G57) );
XOR2_X1 U832 ( .A(n1155), .B(n1156), .Z(n1154) );
XNOR2_X1 U833 ( .A(n1157), .B(n1158), .ZN(n1156) );
XOR2_X1 U834 ( .A(KEYINPUT45), .B(n1159), .Z(n1155) );
AND2_X1 U835 ( .A1(G472), .A2(n1138), .ZN(n1159) );
NOR3_X1 U836 ( .A1(n1160), .A2(n1044), .A3(n1161), .ZN(G54) );
NOR4_X1 U837 ( .A1(n1162), .A2(n1163), .A3(n1055), .A4(n1164), .ZN(n1161) );
XOR2_X1 U838 ( .A(n1165), .B(KEYINPUT63), .Z(n1163) );
NOR2_X1 U839 ( .A1(n1166), .A2(n1167), .ZN(n1160) );
XOR2_X1 U840 ( .A(n1165), .B(KEYINPUT59), .Z(n1167) );
XOR2_X1 U841 ( .A(n1168), .B(n1169), .Z(n1165) );
XOR2_X1 U842 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND3_X1 U843 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1171) );
NAND2_X1 U844 ( .A1(KEYINPUT58), .A2(G140), .ZN(n1174) );
NAND3_X1 U845 ( .A1(n1175), .A2(n1176), .A3(G110), .ZN(n1173) );
NAND2_X1 U846 ( .A1(n1177), .A2(n1178), .ZN(n1172) );
NAND2_X1 U847 ( .A1(n1179), .A2(n1176), .ZN(n1177) );
INV_X1 U848 ( .A(KEYINPUT58), .ZN(n1176) );
XNOR2_X1 U849 ( .A(KEYINPUT31), .B(n1175), .ZN(n1179) );
NAND2_X1 U850 ( .A1(KEYINPUT21), .A2(n1180), .ZN(n1168) );
XNOR2_X1 U851 ( .A(n1104), .B(n1181), .ZN(n1180) );
NOR3_X1 U852 ( .A1(n1164), .A2(n1162), .A3(n1055), .ZN(n1166) );
INV_X1 U853 ( .A(G469), .ZN(n1055) );
XNOR2_X1 U854 ( .A(n1062), .B(KEYINPUT25), .ZN(n1162) );
NOR2_X1 U855 ( .A1(n1044), .A2(n1182), .ZN(G51) );
XOR2_X1 U856 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U857 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U858 ( .A1(n1187), .A2(n1132), .ZN(n1186) );
INV_X1 U859 ( .A(n1138), .ZN(n1132) );
NOR2_X1 U860 ( .A1(n1164), .A2(n1062), .ZN(n1138) );
AND2_X1 U861 ( .A1(n1112), .A2(n1109), .ZN(n1062) );
AND4_X1 U862 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1109) );
NOR4_X1 U863 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
NOR2_X1 U864 ( .A1(n1196), .A2(n1197), .ZN(n1190) );
NOR2_X1 U865 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XNOR2_X1 U866 ( .A(n1200), .B(KEYINPUT37), .ZN(n1198) );
AND4_X1 U867 ( .A1(n1039), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1112) );
NOR4_X1 U868 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203) );
NOR3_X1 U869 ( .A1(n1089), .A2(n1076), .A3(n1208), .ZN(n1207) );
NOR4_X1 U870 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1089), .ZN(n1206) );
NOR2_X1 U871 ( .A1(KEYINPUT18), .A2(n1212), .ZN(n1210) );
NOR2_X1 U872 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NOR2_X1 U873 ( .A1(n1215), .A2(n1216), .ZN(n1209) );
INV_X1 U874 ( .A(KEYINPUT18), .ZN(n1216) );
NOR2_X1 U875 ( .A1(n1152), .A2(n1217), .ZN(n1202) );
AND3_X1 U876 ( .A1(n1215), .A2(n1068), .A3(n1200), .ZN(n1152) );
NAND3_X1 U877 ( .A1(n1218), .A2(n1068), .A3(n1215), .ZN(n1039) );
NAND2_X1 U878 ( .A1(KEYINPUT9), .A2(n1219), .ZN(n1185) );
NOR2_X1 U879 ( .A1(n1108), .A2(G952), .ZN(n1044) );
XNOR2_X1 U880 ( .A(G146), .B(n1220), .ZN(G48) );
OR2_X1 U881 ( .A1(n1199), .A2(n1075), .ZN(n1220) );
XOR2_X1 U882 ( .A(n1189), .B(n1221), .Z(G45) );
XNOR2_X1 U883 ( .A(KEYINPUT12), .B(n1222), .ZN(n1221) );
NAND4_X1 U884 ( .A1(n1213), .A2(n1093), .A3(n1223), .A4(n1224), .ZN(n1189) );
NOR3_X1 U885 ( .A1(n1225), .A2(n1226), .A3(n1227), .ZN(n1224) );
XNOR2_X1 U886 ( .A(G140), .B(n1228), .ZN(G42) );
NOR2_X1 U887 ( .A1(n1195), .A2(KEYINPUT46), .ZN(n1228) );
AND4_X1 U888 ( .A1(n1091), .A2(n1229), .A3(n1200), .A4(n1092), .ZN(n1195) );
XNOR2_X1 U889 ( .A(n1230), .B(n1196), .ZN(G39) );
AND2_X1 U890 ( .A1(n1229), .A2(n1231), .ZN(n1196) );
XOR2_X1 U891 ( .A(G134), .B(n1194), .Z(G36) );
AND3_X1 U892 ( .A1(n1223), .A2(n1218), .A3(n1229), .ZN(n1194) );
XNOR2_X1 U893 ( .A(G131), .B(n1232), .ZN(G33) );
NAND2_X1 U894 ( .A1(KEYINPUT33), .A2(n1193), .ZN(n1232) );
AND3_X1 U895 ( .A1(n1223), .A2(n1200), .A3(n1229), .ZN(n1193) );
NOR4_X1 U896 ( .A1(n1056), .A2(n1078), .A3(n1050), .A4(n1226), .ZN(n1229) );
XOR2_X1 U897 ( .A(G128), .B(n1192), .Z(G30) );
NOR2_X1 U898 ( .A1(n1199), .A2(n1076), .ZN(n1192) );
NAND3_X1 U899 ( .A1(n1051), .A2(n1213), .A3(n1233), .ZN(n1199) );
XOR2_X1 U900 ( .A(G101), .B(n1234), .Z(G3) );
NOR2_X1 U901 ( .A1(n1235), .A2(n1089), .ZN(n1234) );
XNOR2_X1 U902 ( .A(G125), .B(n1188), .ZN(G27) );
NAND4_X1 U903 ( .A1(n1233), .A2(n1200), .A3(n1073), .A4(n1092), .ZN(n1188) );
NOR3_X1 U904 ( .A1(n1236), .A2(n1226), .A3(n1237), .ZN(n1233) );
AND2_X1 U905 ( .A1(n1238), .A2(n1094), .ZN(n1226) );
XOR2_X1 U906 ( .A(KEYINPUT23), .B(n1239), .Z(n1238) );
NOR4_X1 U907 ( .A1(n1240), .A2(n1164), .A3(n1108), .A4(n1107), .ZN(n1239) );
XOR2_X1 U908 ( .A(G900), .B(KEYINPUT51), .Z(n1107) );
INV_X1 U909 ( .A(n1241), .ZN(n1240) );
XOR2_X1 U910 ( .A(n1242), .B(n1243), .Z(G24) );
XOR2_X1 U911 ( .A(KEYINPUT24), .B(G122), .Z(n1243) );
NAND2_X1 U912 ( .A1(KEYINPUT22), .A2(n1244), .ZN(n1242) );
INV_X1 U913 ( .A(n1201), .ZN(n1244) );
NAND4_X1 U914 ( .A1(n1245), .A2(n1068), .A3(n1246), .A4(n1247), .ZN(n1201) );
NOR2_X1 U915 ( .A1(n1051), .A2(n1091), .ZN(n1068) );
XNOR2_X1 U916 ( .A(n1248), .B(n1205), .ZN(G21) );
AND2_X1 U917 ( .A1(n1231), .A2(n1245), .ZN(n1205) );
INV_X1 U918 ( .A(n1208), .ZN(n1245) );
NOR3_X1 U919 ( .A1(n1237), .A2(n1211), .A3(n1092), .ZN(n1231) );
INV_X1 U920 ( .A(n1046), .ZN(n1211) );
XOR2_X1 U921 ( .A(n1249), .B(n1250), .Z(G18) );
XOR2_X1 U922 ( .A(KEYINPUT0), .B(G116), .Z(n1250) );
NAND4_X1 U923 ( .A1(n1223), .A2(n1073), .A3(n1251), .A4(n1252), .ZN(n1249) );
NOR3_X1 U924 ( .A1(n1076), .A2(KEYINPUT14), .A3(n1253), .ZN(n1252) );
INV_X1 U925 ( .A(n1218), .ZN(n1076) );
NOR2_X1 U926 ( .A1(n1247), .A2(n1225), .ZN(n1218) );
INV_X1 U927 ( .A(n1246), .ZN(n1225) );
XNOR2_X1 U928 ( .A(n1093), .B(KEYINPUT27), .ZN(n1251) );
XNOR2_X1 U929 ( .A(n1204), .B(n1254), .ZN(G15) );
XNOR2_X1 U930 ( .A(G113), .B(KEYINPUT5), .ZN(n1254) );
NOR3_X1 U931 ( .A1(n1075), .A2(n1208), .A3(n1089), .ZN(n1204) );
INV_X1 U932 ( .A(n1223), .ZN(n1089) );
NOR2_X1 U933 ( .A1(n1092), .A2(n1091), .ZN(n1223) );
INV_X1 U934 ( .A(n1237), .ZN(n1091) );
NAND2_X1 U935 ( .A1(n1073), .A2(n1255), .ZN(n1208) );
NOR2_X1 U936 ( .A1(n1256), .A2(n1049), .ZN(n1073) );
INV_X1 U937 ( .A(n1200), .ZN(n1075) );
NOR2_X1 U938 ( .A1(n1246), .A2(n1227), .ZN(n1200) );
INV_X1 U939 ( .A(n1247), .ZN(n1227) );
XNOR2_X1 U940 ( .A(n1178), .B(n1217), .ZN(G12) );
NOR3_X1 U941 ( .A1(n1237), .A2(n1051), .A3(n1235), .ZN(n1217) );
NAND2_X1 U942 ( .A1(n1046), .A2(n1215), .ZN(n1235) );
NOR2_X1 U943 ( .A1(n1078), .A2(n1214), .ZN(n1215) );
INV_X1 U944 ( .A(n1255), .ZN(n1214) );
NOR2_X1 U945 ( .A1(n1236), .A2(n1253), .ZN(n1255) );
AND2_X1 U946 ( .A1(n1094), .A2(n1257), .ZN(n1253) );
NAND4_X1 U947 ( .A1(G953), .A2(G902), .A3(n1241), .A4(n1122), .ZN(n1257) );
INV_X1 U948 ( .A(G898), .ZN(n1122) );
NAND3_X1 U949 ( .A1(n1241), .A2(n1108), .A3(G952), .ZN(n1094) );
NAND2_X1 U950 ( .A1(G237), .A2(G234), .ZN(n1241) );
INV_X1 U951 ( .A(n1093), .ZN(n1236) );
NOR2_X1 U952 ( .A1(n1067), .A2(n1050), .ZN(n1093) );
INV_X1 U953 ( .A(n1070), .ZN(n1050) );
NAND2_X1 U954 ( .A1(G214), .A2(n1258), .ZN(n1070) );
INV_X1 U955 ( .A(n1056), .ZN(n1067) );
XOR2_X1 U956 ( .A(n1259), .B(n1187), .Z(n1056) );
NAND2_X1 U957 ( .A1(G210), .A2(n1258), .ZN(n1187) );
NAND2_X1 U958 ( .A1(n1260), .A2(n1164), .ZN(n1258) );
INV_X1 U959 ( .A(G237), .ZN(n1260) );
NAND2_X1 U960 ( .A1(n1261), .A2(n1164), .ZN(n1259) );
XNOR2_X1 U961 ( .A(G125), .B(n1183), .ZN(n1261) );
XNOR2_X1 U962 ( .A(n1262), .B(n1263), .ZN(n1183) );
XOR2_X1 U963 ( .A(n1264), .B(n1265), .Z(n1262) );
NOR2_X1 U964 ( .A1(G953), .A2(n1117), .ZN(n1265) );
INV_X1 U965 ( .A(G224), .ZN(n1117) );
NAND2_X1 U966 ( .A1(n1266), .A2(n1267), .ZN(n1264) );
NAND3_X1 U967 ( .A1(n1124), .A2(n1127), .A3(n1268), .ZN(n1267) );
NAND2_X1 U968 ( .A1(n1269), .A2(n1270), .ZN(n1266) );
NAND2_X1 U969 ( .A1(n1268), .A2(n1127), .ZN(n1270) );
NAND2_X1 U970 ( .A1(n1271), .A2(n1272), .ZN(n1127) );
XNOR2_X1 U971 ( .A(KEYINPUT43), .B(n1273), .ZN(n1271) );
XNOR2_X1 U972 ( .A(n1125), .B(KEYINPUT2), .ZN(n1268) );
AND2_X1 U973 ( .A1(n1274), .A2(n1275), .ZN(n1125) );
XOR2_X1 U974 ( .A(KEYINPUT43), .B(n1273), .Z(n1275) );
XNOR2_X1 U975 ( .A(n1124), .B(KEYINPUT17), .ZN(n1269) );
XNOR2_X1 U976 ( .A(G110), .B(n1276), .ZN(n1124) );
INV_X1 U977 ( .A(n1213), .ZN(n1078) );
NOR2_X1 U978 ( .A1(n1080), .A2(n1049), .ZN(n1213) );
AND2_X1 U979 ( .A1(G221), .A2(n1277), .ZN(n1049) );
INV_X1 U980 ( .A(n1256), .ZN(n1080) );
XOR2_X1 U981 ( .A(n1278), .B(n1053), .Z(n1256) );
NAND2_X1 U982 ( .A1(n1279), .A2(n1164), .ZN(n1053) );
XOR2_X1 U983 ( .A(n1104), .B(n1280), .Z(n1279) );
XOR2_X1 U984 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR2_X1 U985 ( .A1(KEYINPUT35), .A2(n1181), .ZN(n1282) );
XNOR2_X1 U986 ( .A(n1102), .B(n1273), .ZN(n1181) );
XNOR2_X1 U987 ( .A(n1283), .B(n1284), .ZN(n1273) );
XOR2_X1 U988 ( .A(KEYINPUT13), .B(G107), .Z(n1284) );
XNOR2_X1 U989 ( .A(G101), .B(G104), .ZN(n1283) );
XNOR2_X1 U990 ( .A(n1285), .B(n1286), .ZN(n1102) );
XNOR2_X1 U991 ( .A(n1287), .B(n1288), .ZN(n1285) );
NAND2_X1 U992 ( .A1(KEYINPUT55), .A2(n1222), .ZN(n1287) );
NOR2_X1 U993 ( .A1(n1289), .A2(n1290), .ZN(n1281) );
NOR2_X1 U994 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XNOR2_X1 U995 ( .A(G110), .B(G140), .ZN(n1292) );
XOR2_X1 U996 ( .A(n1170), .B(KEYINPUT20), .Z(n1291) );
NOR2_X1 U997 ( .A1(n1293), .A2(n1294), .ZN(n1289) );
XNOR2_X1 U998 ( .A(n1175), .B(G110), .ZN(n1294) );
XOR2_X1 U999 ( .A(n1170), .B(KEYINPUT1), .Z(n1293) );
NAND2_X1 U1000 ( .A1(G227), .A2(n1108), .ZN(n1170) );
NAND2_X1 U1001 ( .A1(KEYINPUT19), .A2(G469), .ZN(n1278) );
NOR2_X1 U1002 ( .A1(n1246), .A2(n1247), .ZN(n1046) );
XNOR2_X1 U1003 ( .A(n1295), .B(G475), .ZN(n1247) );
NAND2_X1 U1004 ( .A1(n1164), .A2(n1145), .ZN(n1295) );
NAND3_X1 U1005 ( .A1(n1296), .A2(n1297), .A3(n1298), .ZN(n1145) );
OR2_X1 U1006 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
NAND2_X1 U1007 ( .A1(n1301), .A2(n1302), .ZN(n1297) );
INV_X1 U1008 ( .A(KEYINPUT6), .ZN(n1302) );
NAND2_X1 U1009 ( .A1(n1303), .A2(n1300), .ZN(n1301) );
XNOR2_X1 U1010 ( .A(KEYINPUT7), .B(n1299), .ZN(n1303) );
NAND2_X1 U1011 ( .A1(KEYINPUT6), .A2(n1304), .ZN(n1296) );
NAND2_X1 U1012 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
OR2_X1 U1013 ( .A1(n1299), .A2(KEYINPUT7), .ZN(n1306) );
NAND3_X1 U1014 ( .A1(n1300), .A2(n1299), .A3(KEYINPUT7), .ZN(n1305) );
XOR2_X1 U1015 ( .A(G104), .B(n1307), .Z(n1299) );
NOR2_X1 U1016 ( .A1(KEYINPUT3), .A2(n1308), .ZN(n1307) );
XNOR2_X1 U1017 ( .A(G113), .B(n1276), .ZN(n1308) );
XNOR2_X1 U1018 ( .A(n1309), .B(n1310), .ZN(n1300) );
XNOR2_X1 U1019 ( .A(n1219), .B(n1311), .ZN(n1310) );
XNOR2_X1 U1020 ( .A(n1288), .B(G131), .ZN(n1311) );
INV_X1 U1021 ( .A(G125), .ZN(n1219) );
XOR2_X1 U1022 ( .A(n1312), .B(n1313), .Z(n1309) );
XOR2_X1 U1023 ( .A(n1314), .B(n1315), .Z(n1313) );
NAND2_X1 U1024 ( .A1(n1316), .A2(G214), .ZN(n1315) );
NAND2_X1 U1025 ( .A1(KEYINPUT54), .A2(G140), .ZN(n1314) );
NAND2_X1 U1026 ( .A1(KEYINPUT15), .A2(n1222), .ZN(n1312) );
XNOR2_X1 U1027 ( .A(n1317), .B(G478), .ZN(n1246) );
NAND2_X1 U1028 ( .A1(n1164), .A2(n1136), .ZN(n1317) );
NAND2_X1 U1029 ( .A1(n1318), .A2(n1319), .ZN(n1136) );
NAND4_X1 U1030 ( .A1(G217), .A2(n1320), .A3(n1321), .A4(n1322), .ZN(n1319) );
NAND2_X1 U1031 ( .A1(n1323), .A2(n1324), .ZN(n1318) );
NAND2_X1 U1032 ( .A1(G217), .A2(n1320), .ZN(n1324) );
INV_X1 U1033 ( .A(n1325), .ZN(n1320) );
NAND2_X1 U1034 ( .A1(n1321), .A2(n1322), .ZN(n1323) );
NAND2_X1 U1035 ( .A1(n1326), .A2(n1327), .ZN(n1322) );
XOR2_X1 U1036 ( .A(n1328), .B(G107), .Z(n1327) );
XNOR2_X1 U1037 ( .A(n1329), .B(KEYINPUT41), .ZN(n1326) );
XOR2_X1 U1038 ( .A(n1330), .B(KEYINPUT11), .Z(n1321) );
NAND2_X1 U1039 ( .A1(n1331), .A2(n1329), .ZN(n1330) );
XNOR2_X1 U1040 ( .A(n1332), .B(n1333), .ZN(n1329) );
XNOR2_X1 U1041 ( .A(KEYINPUT57), .B(n1222), .ZN(n1333) );
INV_X1 U1042 ( .A(G143), .ZN(n1222) );
XNOR2_X1 U1043 ( .A(G134), .B(n1334), .ZN(n1332) );
XNOR2_X1 U1044 ( .A(G107), .B(n1328), .ZN(n1331) );
NAND3_X1 U1045 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1328) );
NAND2_X1 U1046 ( .A1(KEYINPUT56), .A2(n1276), .ZN(n1337) );
INV_X1 U1047 ( .A(n1338), .ZN(n1276) );
OR3_X1 U1048 ( .A1(n1339), .A2(KEYINPUT56), .A3(G116), .ZN(n1336) );
NAND2_X1 U1049 ( .A1(G116), .A2(n1339), .ZN(n1335) );
NAND2_X1 U1050 ( .A1(KEYINPUT52), .A2(n1338), .ZN(n1339) );
XOR2_X1 U1051 ( .A(G122), .B(KEYINPUT62), .Z(n1338) );
INV_X1 U1052 ( .A(n1092), .ZN(n1051) );
XNOR2_X1 U1053 ( .A(n1340), .B(n1341), .ZN(n1092) );
XOR2_X1 U1054 ( .A(KEYINPUT28), .B(G472), .Z(n1341) );
NAND2_X1 U1055 ( .A1(n1342), .A2(n1164), .ZN(n1340) );
XOR2_X1 U1056 ( .A(n1157), .B(n1343), .Z(n1342) );
XNOR2_X1 U1057 ( .A(KEYINPUT34), .B(n1344), .ZN(n1343) );
NOR2_X1 U1058 ( .A1(KEYINPUT40), .A2(n1263), .ZN(n1344) );
INV_X1 U1059 ( .A(n1158), .ZN(n1263) );
XOR2_X1 U1060 ( .A(n1345), .B(n1286), .Z(n1158) );
INV_X1 U1061 ( .A(n1334), .ZN(n1286) );
NAND2_X1 U1062 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
NAND2_X1 U1063 ( .A1(n1348), .A2(n1288), .ZN(n1347) );
XOR2_X1 U1064 ( .A(KEYINPUT50), .B(n1349), .Z(n1346) );
NOR2_X1 U1065 ( .A1(n1348), .A2(n1288), .ZN(n1349) );
XNOR2_X1 U1066 ( .A(KEYINPUT60), .B(G143), .ZN(n1348) );
XOR2_X1 U1067 ( .A(n1350), .B(n1351), .Z(n1157) );
XNOR2_X1 U1068 ( .A(G101), .B(n1352), .ZN(n1351) );
NAND2_X1 U1069 ( .A1(n1316), .A2(G210), .ZN(n1352) );
NOR2_X1 U1070 ( .A1(G953), .A2(G237), .ZN(n1316) );
XNOR2_X1 U1071 ( .A(n1104), .B(n1274), .ZN(n1350) );
INV_X1 U1072 ( .A(n1272), .ZN(n1274) );
XOR2_X1 U1073 ( .A(G113), .B(n1353), .Z(n1272) );
XNOR2_X1 U1074 ( .A(n1248), .B(G116), .ZN(n1353) );
INV_X1 U1075 ( .A(G119), .ZN(n1248) );
XNOR2_X1 U1076 ( .A(G131), .B(n1354), .ZN(n1104) );
XNOR2_X1 U1077 ( .A(n1230), .B(G134), .ZN(n1354) );
XNOR2_X1 U1078 ( .A(n1355), .B(n1057), .ZN(n1237) );
NOR2_X1 U1079 ( .A1(n1134), .A2(G902), .ZN(n1057) );
INV_X1 U1080 ( .A(n1131), .ZN(n1134) );
XNOR2_X1 U1081 ( .A(n1356), .B(n1357), .ZN(n1131) );
XNOR2_X1 U1082 ( .A(n1358), .B(n1334), .ZN(n1357) );
XOR2_X1 U1083 ( .A(G128), .B(KEYINPUT38), .Z(n1334) );
NAND3_X1 U1084 ( .A1(n1359), .A2(n1360), .A3(n1361), .ZN(n1358) );
OR2_X1 U1085 ( .A1(n1105), .A2(KEYINPUT47), .ZN(n1361) );
NAND3_X1 U1086 ( .A1(KEYINPUT47), .A2(n1362), .A3(n1288), .ZN(n1360) );
INV_X1 U1087 ( .A(G146), .ZN(n1288) );
INV_X1 U1088 ( .A(n1363), .ZN(n1362) );
NAND2_X1 U1089 ( .A1(G146), .A2(n1363), .ZN(n1359) );
NAND2_X1 U1090 ( .A1(KEYINPUT8), .A2(n1105), .ZN(n1363) );
XNOR2_X1 U1091 ( .A(G125), .B(n1175), .ZN(n1105) );
INV_X1 U1092 ( .A(G140), .ZN(n1175) );
XOR2_X1 U1093 ( .A(n1364), .B(n1365), .Z(n1356) );
NOR3_X1 U1094 ( .A1(n1366), .A2(KEYINPUT16), .A3(n1367), .ZN(n1365) );
NOR3_X1 U1095 ( .A1(n1368), .A2(n1369), .A3(n1325), .ZN(n1367) );
XNOR2_X1 U1096 ( .A(G137), .B(n1370), .ZN(n1368) );
XNOR2_X1 U1097 ( .A(KEYINPUT48), .B(KEYINPUT30), .ZN(n1370) );
NOR2_X1 U1098 ( .A1(n1371), .A2(n1230), .ZN(n1366) );
INV_X1 U1099 ( .A(G137), .ZN(n1230) );
NOR2_X1 U1100 ( .A1(n1369), .A2(n1325), .ZN(n1371) );
NAND2_X1 U1101 ( .A1(G234), .A2(n1108), .ZN(n1325) );
INV_X1 U1102 ( .A(G953), .ZN(n1108) );
INV_X1 U1103 ( .A(G221), .ZN(n1369) );
XNOR2_X1 U1104 ( .A(G119), .B(G110), .ZN(n1364) );
NAND2_X1 U1105 ( .A1(KEYINPUT39), .A2(n1058), .ZN(n1355) );
NAND2_X1 U1106 ( .A1(G217), .A2(n1277), .ZN(n1058) );
NAND2_X1 U1107 ( .A1(G234), .A2(n1164), .ZN(n1277) );
INV_X1 U1108 ( .A(G902), .ZN(n1164) );
INV_X1 U1109 ( .A(G110), .ZN(n1178) );
endmodule


