//Key = 0101110000101001110101001011111011111110110010000010010111110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407;

XNOR2_X1 U770 ( .A(n1071), .B(n1072), .ZN(G9) );
NOR2_X1 U771 ( .A1(n1073), .A2(n1074), .ZN(G75) );
NOR4_X1 U772 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
INV_X1 U773 ( .A(G952), .ZN(n1078) );
XOR2_X1 U774 ( .A(n1079), .B(KEYINPUT39), .Z(n1077) );
NAND2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND3_X1 U776 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NAND2_X1 U777 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NAND2_X1 U778 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND3_X1 U780 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
NAND3_X1 U781 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1089) );
NAND3_X1 U782 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1085) );
NAND2_X1 U783 ( .A1(n1100), .A2(n1101), .ZN(n1080) );
INV_X1 U784 ( .A(n1102), .ZN(n1076) );
NAND4_X1 U785 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1075) );
NAND3_X1 U786 ( .A1(n1082), .A2(n1107), .A3(n1084), .ZN(n1104) );
INV_X1 U787 ( .A(n1108), .ZN(n1084) );
NAND2_X1 U788 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
NAND2_X1 U789 ( .A1(n1087), .A2(n1111), .ZN(n1110) );
NAND2_X1 U790 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U791 ( .A1(n1091), .A2(n1114), .ZN(n1113) );
NAND2_X1 U792 ( .A1(n1115), .A2(n1096), .ZN(n1112) );
NAND2_X1 U793 ( .A1(n1098), .A2(n1116), .ZN(n1109) );
INV_X1 U794 ( .A(n1117), .ZN(n1098) );
NAND2_X1 U795 ( .A1(n1100), .A2(n1118), .ZN(n1103) );
NOR3_X1 U796 ( .A1(n1119), .A2(n1117), .A3(n1108), .ZN(n1100) );
NOR3_X1 U797 ( .A1(n1120), .A2(G953), .A3(n1121), .ZN(n1073) );
INV_X1 U798 ( .A(n1105), .ZN(n1121) );
NAND4_X1 U799 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1105) );
NOR4_X1 U800 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n1125) );
XNOR2_X1 U801 ( .A(G469), .B(n1130), .ZN(n1129) );
XNOR2_X1 U802 ( .A(n1131), .B(n1132), .ZN(n1128) );
NOR3_X1 U803 ( .A1(n1099), .A2(n1133), .A3(n1093), .ZN(n1124) );
NAND2_X1 U804 ( .A1(G475), .A2(n1134), .ZN(n1123) );
XNOR2_X1 U805 ( .A(n1135), .B(n1136), .ZN(n1122) );
NAND2_X1 U806 ( .A1(KEYINPUT10), .A2(n1137), .ZN(n1136) );
XNOR2_X1 U807 ( .A(G952), .B(KEYINPUT28), .ZN(n1120) );
NAND2_X1 U808 ( .A1(n1138), .A2(n1139), .ZN(G72) );
NAND2_X1 U809 ( .A1(n1140), .A2(n1106), .ZN(n1139) );
XOR2_X1 U810 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U811 ( .A1(KEYINPUT40), .A2(n1143), .ZN(n1142) );
NAND2_X1 U812 ( .A1(n1144), .A2(G953), .ZN(n1138) );
XOR2_X1 U813 ( .A(n1141), .B(n1145), .Z(n1144) );
AND2_X1 U814 ( .A1(G227), .A2(G900), .ZN(n1145) );
NAND2_X1 U815 ( .A1(n1146), .A2(n1147), .ZN(n1141) );
NAND2_X1 U816 ( .A1(G953), .A2(n1148), .ZN(n1147) );
XOR2_X1 U817 ( .A(n1149), .B(n1150), .Z(n1146) );
XOR2_X1 U818 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U819 ( .A1(KEYINPUT16), .A2(n1153), .ZN(n1152) );
NAND3_X1 U820 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1151) );
OR2_X1 U821 ( .A1(n1157), .A2(KEYINPUT37), .ZN(n1156) );
NAND3_X1 U822 ( .A1(KEYINPUT37), .A2(G125), .A3(G140), .ZN(n1155) );
NAND2_X1 U823 ( .A1(n1158), .A2(n1159), .ZN(n1154) );
XNOR2_X1 U824 ( .A(KEYINPUT15), .B(n1160), .ZN(n1158) );
XOR2_X1 U825 ( .A(n1161), .B(n1162), .Z(G69) );
XOR2_X1 U826 ( .A(n1163), .B(n1164), .Z(n1162) );
NAND2_X1 U827 ( .A1(KEYINPUT19), .A2(n1165), .ZN(n1164) );
NAND2_X1 U828 ( .A1(G953), .A2(n1166), .ZN(n1165) );
NAND2_X1 U829 ( .A1(n1167), .A2(G224), .ZN(n1166) );
XNOR2_X1 U830 ( .A(G898), .B(KEYINPUT4), .ZN(n1167) );
NAND2_X1 U831 ( .A1(n1168), .A2(n1169), .ZN(n1163) );
NAND2_X1 U832 ( .A1(G953), .A2(n1170), .ZN(n1169) );
XNOR2_X1 U833 ( .A(KEYINPUT41), .B(n1171), .ZN(n1170) );
XOR2_X1 U834 ( .A(n1172), .B(n1173), .Z(n1168) );
XNOR2_X1 U835 ( .A(KEYINPUT54), .B(n1174), .ZN(n1173) );
NOR2_X1 U836 ( .A1(KEYINPUT48), .A2(n1175), .ZN(n1174) );
XNOR2_X1 U837 ( .A(n1176), .B(n1177), .ZN(n1175) );
NAND2_X1 U838 ( .A1(n1106), .A2(n1178), .ZN(n1161) );
NOR2_X1 U839 ( .A1(n1179), .A2(n1180), .ZN(G66) );
XNOR2_X1 U840 ( .A(n1181), .B(n1182), .ZN(n1180) );
NOR2_X1 U841 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NOR2_X1 U842 ( .A1(n1179), .A2(n1185), .ZN(G63) );
NOR3_X1 U843 ( .A1(n1135), .A2(n1186), .A3(n1187), .ZN(n1185) );
AND3_X1 U844 ( .A1(n1188), .A2(G478), .A3(n1189), .ZN(n1187) );
NOR2_X1 U845 ( .A1(n1190), .A2(n1188), .ZN(n1186) );
NOR2_X1 U846 ( .A1(n1102), .A2(n1137), .ZN(n1190) );
NOR2_X1 U847 ( .A1(n1179), .A2(n1191), .ZN(G60) );
XNOR2_X1 U848 ( .A(n1192), .B(n1193), .ZN(n1191) );
NOR2_X1 U849 ( .A1(n1194), .A2(n1184), .ZN(n1193) );
XNOR2_X1 U850 ( .A(G104), .B(n1195), .ZN(G6) );
NOR2_X1 U851 ( .A1(n1196), .A2(n1197), .ZN(G57) );
XNOR2_X1 U852 ( .A(n1179), .B(KEYINPUT30), .ZN(n1197) );
XNOR2_X1 U853 ( .A(n1198), .B(n1199), .ZN(n1196) );
XOR2_X1 U854 ( .A(n1200), .B(n1201), .Z(n1199) );
AND2_X1 U855 ( .A1(G472), .A2(n1189), .ZN(n1201) );
NOR3_X1 U856 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1200) );
NOR2_X1 U857 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XOR2_X1 U858 ( .A(n1207), .B(KEYINPUT63), .Z(n1206) );
AND3_X1 U859 ( .A1(n1205), .A2(n1208), .A3(n1209), .ZN(n1203) );
INV_X1 U860 ( .A(KEYINPUT49), .ZN(n1205) );
NOR2_X1 U861 ( .A1(n1209), .A2(n1208), .ZN(n1202) );
XOR2_X1 U862 ( .A(G101), .B(KEYINPUT35), .Z(n1208) );
NOR2_X1 U863 ( .A1(KEYINPUT9), .A2(n1210), .ZN(n1209) );
XNOR2_X1 U864 ( .A(KEYINPUT63), .B(n1207), .ZN(n1210) );
NOR2_X1 U865 ( .A1(n1179), .A2(n1211), .ZN(G54) );
NOR2_X1 U866 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NOR2_X1 U867 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XNOR2_X1 U868 ( .A(n1216), .B(n1217), .ZN(n1215) );
NOR2_X1 U869 ( .A1(n1218), .A2(n1219), .ZN(n1214) );
NOR3_X1 U870 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1212) );
NOR2_X1 U871 ( .A1(n1222), .A2(n1216), .ZN(n1221) );
NOR2_X1 U872 ( .A1(n1217), .A2(n1218), .ZN(n1222) );
NOR2_X1 U873 ( .A1(n1223), .A2(n1224), .ZN(n1220) );
AND2_X1 U874 ( .A1(n1217), .A2(n1225), .ZN(n1224) );
INV_X1 U875 ( .A(n1216), .ZN(n1223) );
NAND2_X1 U876 ( .A1(n1189), .A2(G469), .ZN(n1216) );
INV_X1 U877 ( .A(KEYINPUT59), .ZN(n1219) );
NOR2_X1 U878 ( .A1(n1226), .A2(n1227), .ZN(G51) );
XOR2_X1 U879 ( .A(n1228), .B(n1229), .Z(n1227) );
XNOR2_X1 U880 ( .A(n1230), .B(n1231), .ZN(n1229) );
NOR2_X1 U881 ( .A1(n1131), .A2(n1184), .ZN(n1231) );
INV_X1 U882 ( .A(n1189), .ZN(n1184) );
NOR2_X1 U883 ( .A1(n1232), .A2(n1102), .ZN(n1189) );
NOR2_X1 U884 ( .A1(n1178), .A2(n1143), .ZN(n1102) );
NAND4_X1 U885 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1143) );
NOR4_X1 U886 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1236) );
NOR2_X1 U887 ( .A1(n1241), .A2(n1242), .ZN(n1235) );
INV_X1 U888 ( .A(n1243), .ZN(n1241) );
OR2_X1 U889 ( .A1(n1244), .A2(n1119), .ZN(n1233) );
NAND4_X1 U890 ( .A1(n1245), .A2(n1195), .A3(n1246), .A4(n1247), .ZN(n1178) );
NOR4_X1 U891 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1072), .ZN(n1247) );
AND3_X1 U892 ( .A1(n1101), .A2(n1091), .A3(n1251), .ZN(n1072) );
NOR3_X1 U893 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1246) );
NOR2_X1 U894 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
INV_X1 U895 ( .A(KEYINPUT12), .ZN(n1255) );
NOR4_X1 U896 ( .A1(KEYINPUT12), .A2(n1257), .A3(n1258), .A4(n1117), .ZN(n1253) );
NAND2_X1 U897 ( .A1(n1096), .A2(n1091), .ZN(n1117) );
NAND3_X1 U898 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1257) );
INV_X1 U899 ( .A(n1116), .ZN(n1260) );
NAND3_X1 U900 ( .A1(n1251), .A2(n1091), .A3(n1118), .ZN(n1195) );
XNOR2_X1 U901 ( .A(KEYINPUT23), .B(n1262), .ZN(n1228) );
NOR2_X1 U902 ( .A1(KEYINPUT62), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U903 ( .A(n1264), .B(n1160), .ZN(n1263) );
XNOR2_X1 U904 ( .A(n1179), .B(KEYINPUT34), .ZN(n1226) );
AND2_X1 U905 ( .A1(n1265), .A2(G953), .ZN(n1179) );
XNOR2_X1 U906 ( .A(G952), .B(KEYINPUT42), .ZN(n1265) );
XNOR2_X1 U907 ( .A(n1266), .B(n1240), .ZN(G48) );
AND3_X1 U908 ( .A1(n1118), .A2(n1116), .A3(n1267), .ZN(n1240) );
NAND2_X1 U909 ( .A1(n1268), .A2(n1269), .ZN(G45) );
OR2_X1 U910 ( .A1(n1234), .A2(G143), .ZN(n1269) );
XOR2_X1 U911 ( .A(n1270), .B(KEYINPUT0), .Z(n1268) );
NAND2_X1 U912 ( .A1(G143), .A2(n1234), .ZN(n1270) );
NAND4_X1 U913 ( .A1(n1271), .A2(n1116), .A3(n1272), .A4(n1261), .ZN(n1234) );
XNOR2_X1 U914 ( .A(n1159), .B(n1242), .ZN(G42) );
AND3_X1 U915 ( .A1(n1087), .A2(n1114), .A3(n1273), .ZN(n1242) );
XNOR2_X1 U916 ( .A(G137), .B(n1274), .ZN(G39) );
NAND2_X1 U917 ( .A1(KEYINPUT27), .A2(n1239), .ZN(n1274) );
AND3_X1 U918 ( .A1(n1267), .A2(n1082), .A3(n1087), .ZN(n1239) );
XOR2_X1 U919 ( .A(n1238), .B(n1275), .Z(G36) );
NOR2_X1 U920 ( .A1(KEYINPUT22), .A2(n1276), .ZN(n1275) );
AND3_X1 U921 ( .A1(n1271), .A2(n1101), .A3(n1087), .ZN(n1238) );
INV_X1 U922 ( .A(n1119), .ZN(n1087) );
XOR2_X1 U923 ( .A(G131), .B(n1277), .Z(G33) );
NOR2_X1 U924 ( .A1(n1278), .A2(n1119), .ZN(n1277) );
NAND2_X1 U925 ( .A1(n1097), .A2(n1279), .ZN(n1119) );
XOR2_X1 U926 ( .A(n1244), .B(KEYINPUT51), .Z(n1278) );
NAND2_X1 U927 ( .A1(n1271), .A2(n1118), .ZN(n1244) );
AND3_X1 U928 ( .A1(n1114), .A2(n1280), .A3(n1115), .ZN(n1271) );
XOR2_X1 U929 ( .A(n1237), .B(n1281), .Z(G30) );
NOR2_X1 U930 ( .A1(KEYINPUT7), .A2(n1282), .ZN(n1281) );
AND3_X1 U931 ( .A1(n1101), .A2(n1116), .A3(n1267), .ZN(n1237) );
AND4_X1 U932 ( .A1(n1283), .A2(n1094), .A3(n1114), .A4(n1280), .ZN(n1267) );
XNOR2_X1 U933 ( .A(n1284), .B(n1250), .ZN(G3) );
AND3_X1 U934 ( .A1(n1082), .A2(n1251), .A3(n1115), .ZN(n1250) );
XNOR2_X1 U935 ( .A(G125), .B(n1243), .ZN(G27) );
NAND3_X1 U936 ( .A1(n1096), .A2(n1116), .A3(n1273), .ZN(n1243) );
AND4_X1 U937 ( .A1(n1094), .A2(n1118), .A3(n1095), .A4(n1280), .ZN(n1273) );
NAND2_X1 U938 ( .A1(n1108), .A2(n1285), .ZN(n1280) );
NAND4_X1 U939 ( .A1(G953), .A2(G902), .A3(n1286), .A4(n1148), .ZN(n1285) );
INV_X1 U940 ( .A(G900), .ZN(n1148) );
XOR2_X1 U941 ( .A(n1256), .B(n1287), .Z(G24) );
XNOR2_X1 U942 ( .A(KEYINPUT58), .B(n1288), .ZN(n1287) );
NAND4_X1 U943 ( .A1(n1289), .A2(n1091), .A3(n1272), .A4(n1261), .ZN(n1256) );
NOR2_X1 U944 ( .A1(n1290), .A2(n1094), .ZN(n1091) );
INV_X1 U945 ( .A(n1095), .ZN(n1290) );
NAND3_X1 U946 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(G21) );
NAND2_X1 U947 ( .A1(n1252), .A2(n1294), .ZN(n1293) );
NAND2_X1 U948 ( .A1(n1295), .A2(n1296), .ZN(n1292) );
INV_X1 U949 ( .A(KEYINPUT36), .ZN(n1296) );
NAND2_X1 U950 ( .A1(n1297), .A2(n1298), .ZN(n1295) );
XNOR2_X1 U951 ( .A(KEYINPUT31), .B(n1294), .ZN(n1297) );
NAND2_X1 U952 ( .A1(KEYINPUT36), .A2(n1299), .ZN(n1291) );
NAND2_X1 U953 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
OR3_X1 U954 ( .A1(n1294), .A2(n1252), .A3(KEYINPUT31), .ZN(n1301) );
INV_X1 U955 ( .A(n1298), .ZN(n1252) );
NAND4_X1 U956 ( .A1(n1283), .A2(n1289), .A3(n1094), .A4(n1082), .ZN(n1298) );
INV_X1 U957 ( .A(n1302), .ZN(n1283) );
NAND2_X1 U958 ( .A1(KEYINPUT31), .A2(n1294), .ZN(n1300) );
XNOR2_X1 U959 ( .A(G116), .B(n1245), .ZN(G18) );
NAND3_X1 U960 ( .A1(n1115), .A2(n1101), .A3(n1289), .ZN(n1245) );
NOR2_X1 U961 ( .A1(n1261), .A2(n1258), .ZN(n1101) );
XNOR2_X1 U962 ( .A(n1303), .B(n1249), .ZN(G15) );
AND3_X1 U963 ( .A1(n1289), .A2(n1115), .A3(n1118), .ZN(n1249) );
AND2_X1 U964 ( .A1(n1304), .A2(n1261), .ZN(n1118) );
XNOR2_X1 U965 ( .A(n1272), .B(KEYINPUT60), .ZN(n1304) );
NOR2_X1 U966 ( .A1(n1302), .A2(n1094), .ZN(n1115) );
XOR2_X1 U967 ( .A(n1095), .B(KEYINPUT18), .Z(n1302) );
AND3_X1 U968 ( .A1(n1116), .A2(n1259), .A3(n1096), .ZN(n1289) );
AND2_X1 U969 ( .A1(n1092), .A2(n1305), .ZN(n1096) );
XNOR2_X1 U970 ( .A(n1306), .B(KEYINPUT17), .ZN(n1092) );
XNOR2_X1 U971 ( .A(n1248), .B(n1307), .ZN(G12) );
NAND2_X1 U972 ( .A1(KEYINPUT29), .A2(G110), .ZN(n1307) );
AND4_X1 U973 ( .A1(n1094), .A2(n1082), .A3(n1251), .A4(n1095), .ZN(n1248) );
XOR2_X1 U974 ( .A(n1127), .B(KEYINPUT56), .Z(n1095) );
XNOR2_X1 U975 ( .A(n1308), .B(G472), .ZN(n1127) );
NAND2_X1 U976 ( .A1(n1309), .A2(n1232), .ZN(n1308) );
XOR2_X1 U977 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U978 ( .A(G101), .B(n1207), .ZN(n1311) );
NAND2_X1 U979 ( .A1(n1312), .A2(G210), .ZN(n1207) );
NOR2_X1 U980 ( .A1(KEYINPUT20), .A2(n1198), .ZN(n1310) );
XNOR2_X1 U981 ( .A(n1313), .B(n1314), .ZN(n1198) );
XOR2_X1 U982 ( .A(n1153), .B(n1315), .Z(n1314) );
XOR2_X1 U983 ( .A(G137), .B(G131), .Z(n1315) );
XNOR2_X1 U984 ( .A(n1264), .B(n1316), .ZN(n1313) );
AND3_X1 U985 ( .A1(n1116), .A2(n1259), .A3(n1114), .ZN(n1251) );
NOR2_X1 U986 ( .A1(n1306), .A2(n1093), .ZN(n1114) );
INV_X1 U987 ( .A(n1305), .ZN(n1093) );
NAND2_X1 U988 ( .A1(G221), .A2(n1317), .ZN(n1305) );
NAND3_X1 U989 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1306) );
OR2_X1 U990 ( .A1(n1321), .A2(G469), .ZN(n1320) );
NAND3_X1 U991 ( .A1(G469), .A2(n1321), .A3(KEYINPUT3), .ZN(n1319) );
NOR2_X1 U992 ( .A1(KEYINPUT47), .A2(n1130), .ZN(n1321) );
NAND2_X1 U993 ( .A1(n1130), .A2(n1322), .ZN(n1318) );
INV_X1 U994 ( .A(KEYINPUT3), .ZN(n1322) );
NAND2_X1 U995 ( .A1(n1323), .A2(n1232), .ZN(n1130) );
XNOR2_X1 U996 ( .A(n1217), .B(n1324), .ZN(n1323) );
XNOR2_X1 U997 ( .A(KEYINPUT52), .B(n1325), .ZN(n1324) );
NOR2_X1 U998 ( .A1(KEYINPUT25), .A2(n1225), .ZN(n1325) );
INV_X1 U999 ( .A(n1218), .ZN(n1225) );
XNOR2_X1 U1000 ( .A(n1326), .B(n1327), .ZN(n1218) );
XNOR2_X1 U1001 ( .A(n1159), .B(G110), .ZN(n1327) );
NAND2_X1 U1002 ( .A1(G227), .A2(n1106), .ZN(n1326) );
XNOR2_X1 U1003 ( .A(n1328), .B(n1329), .ZN(n1217) );
XOR2_X1 U1004 ( .A(n1330), .B(n1331), .Z(n1329) );
XNOR2_X1 U1005 ( .A(G104), .B(G107), .ZN(n1331) );
NAND2_X1 U1006 ( .A1(KEYINPUT24), .A2(n1284), .ZN(n1330) );
INV_X1 U1007 ( .A(G101), .ZN(n1284) );
XNOR2_X1 U1008 ( .A(n1149), .B(n1153), .ZN(n1328) );
XNOR2_X1 U1009 ( .A(n1276), .B(KEYINPUT50), .ZN(n1153) );
XNOR2_X1 U1010 ( .A(n1332), .B(n1333), .ZN(n1149) );
XOR2_X1 U1011 ( .A(n1334), .B(n1335), .Z(n1333) );
NOR2_X1 U1012 ( .A1(KEYINPUT14), .A2(n1282), .ZN(n1334) );
INV_X1 U1013 ( .A(G128), .ZN(n1282) );
NAND2_X1 U1014 ( .A1(n1108), .A2(n1336), .ZN(n1259) );
NAND4_X1 U1015 ( .A1(G953), .A2(G902), .A3(n1286), .A4(n1171), .ZN(n1336) );
INV_X1 U1016 ( .A(G898), .ZN(n1171) );
NAND3_X1 U1017 ( .A1(n1286), .A2(n1106), .A3(G952), .ZN(n1108) );
NAND2_X1 U1018 ( .A1(G237), .A2(G234), .ZN(n1286) );
NOR2_X1 U1019 ( .A1(n1097), .A2(n1099), .ZN(n1116) );
INV_X1 U1020 ( .A(n1279), .ZN(n1099) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1337), .ZN(n1279) );
XNOR2_X1 U1022 ( .A(n1338), .B(n1131), .ZN(n1097) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1337), .ZN(n1131) );
NAND2_X1 U1024 ( .A1(n1339), .A2(n1232), .ZN(n1337) );
INV_X1 U1025 ( .A(G237), .ZN(n1339) );
NAND2_X1 U1026 ( .A1(KEYINPUT26), .A2(n1132), .ZN(n1338) );
AND2_X1 U1027 ( .A1(n1340), .A2(n1232), .ZN(n1132) );
XNOR2_X1 U1028 ( .A(n1341), .B(n1342), .ZN(n1340) );
INV_X1 U1029 ( .A(n1230), .ZN(n1342) );
XNOR2_X1 U1030 ( .A(n1343), .B(n1344), .ZN(n1230) );
XOR2_X1 U1031 ( .A(n1345), .B(n1346), .Z(n1344) );
NAND2_X1 U1032 ( .A1(KEYINPUT21), .A2(n1316), .ZN(n1346) );
INV_X1 U1033 ( .A(n1176), .ZN(n1316) );
XOR2_X1 U1034 ( .A(G113), .B(n1347), .Z(n1176) );
XNOR2_X1 U1035 ( .A(n1294), .B(G116), .ZN(n1347) );
INV_X1 U1036 ( .A(G119), .ZN(n1294) );
NAND2_X1 U1037 ( .A1(G224), .A2(n1106), .ZN(n1345) );
XNOR2_X1 U1038 ( .A(n1177), .B(n1172), .ZN(n1343) );
NAND2_X1 U1039 ( .A1(n1348), .A2(n1349), .ZN(n1172) );
NAND2_X1 U1040 ( .A1(n1350), .A2(G110), .ZN(n1349) );
XOR2_X1 U1041 ( .A(KEYINPUT61), .B(n1351), .Z(n1348) );
NOR2_X1 U1042 ( .A1(G110), .A2(n1350), .ZN(n1351) );
XNOR2_X1 U1043 ( .A(KEYINPUT11), .B(G122), .ZN(n1350) );
XOR2_X1 U1044 ( .A(n1352), .B(n1353), .Z(n1177) );
XNOR2_X1 U1045 ( .A(n1354), .B(G101), .ZN(n1353) );
INV_X1 U1046 ( .A(G104), .ZN(n1354) );
NAND2_X1 U1047 ( .A1(KEYINPUT32), .A2(n1071), .ZN(n1352) );
XNOR2_X1 U1048 ( .A(G125), .B(n1355), .ZN(n1341) );
NOR2_X1 U1049 ( .A1(KEYINPUT46), .A2(n1264), .ZN(n1355) );
XNOR2_X1 U1050 ( .A(G128), .B(n1356), .ZN(n1264) );
NOR2_X1 U1051 ( .A1(KEYINPUT2), .A2(n1357), .ZN(n1356) );
XOR2_X1 U1052 ( .A(G143), .B(n1358), .Z(n1357) );
NOR2_X1 U1053 ( .A1(G146), .A2(KEYINPUT13), .ZN(n1358) );
NOR2_X1 U1054 ( .A1(n1272), .A2(n1261), .ZN(n1082) );
NAND3_X1 U1055 ( .A1(n1359), .A2(n1360), .A3(n1361), .ZN(n1261) );
INV_X1 U1056 ( .A(n1133), .ZN(n1361) );
NOR2_X1 U1057 ( .A1(n1134), .A2(G475), .ZN(n1133) );
NAND3_X1 U1058 ( .A1(G475), .A2(n1134), .A3(n1362), .ZN(n1360) );
INV_X1 U1059 ( .A(KEYINPUT8), .ZN(n1362) );
NAND2_X1 U1060 ( .A1(n1192), .A2(n1232), .ZN(n1134) );
XNOR2_X1 U1061 ( .A(n1363), .B(n1364), .ZN(n1192) );
XOR2_X1 U1062 ( .A(n1365), .B(n1332), .Z(n1364) );
XNOR2_X1 U1063 ( .A(G131), .B(G143), .ZN(n1332) );
NAND2_X1 U1064 ( .A1(n1312), .A2(G214), .ZN(n1365) );
NOR2_X1 U1065 ( .A1(G953), .A2(G237), .ZN(n1312) );
XOR2_X1 U1066 ( .A(n1366), .B(n1367), .Z(n1363) );
XNOR2_X1 U1067 ( .A(G104), .B(n1368), .ZN(n1367) );
NAND3_X1 U1068 ( .A1(n1369), .A2(n1370), .A3(n1371), .ZN(n1368) );
NAND2_X1 U1069 ( .A1(G122), .A2(n1303), .ZN(n1371) );
INV_X1 U1070 ( .A(G113), .ZN(n1303) );
NAND2_X1 U1071 ( .A1(n1372), .A2(n1373), .ZN(n1370) );
INV_X1 U1072 ( .A(KEYINPUT33), .ZN(n1373) );
NAND2_X1 U1073 ( .A1(n1374), .A2(n1288), .ZN(n1372) );
XNOR2_X1 U1074 ( .A(KEYINPUT1), .B(G113), .ZN(n1374) );
NAND2_X1 U1075 ( .A1(KEYINPUT33), .A2(n1375), .ZN(n1369) );
NAND2_X1 U1076 ( .A1(n1376), .A2(n1377), .ZN(n1375) );
OR2_X1 U1077 ( .A1(G113), .A2(KEYINPUT1), .ZN(n1377) );
NAND3_X1 U1078 ( .A1(G113), .A2(n1288), .A3(KEYINPUT1), .ZN(n1376) );
INV_X1 U1079 ( .A(G122), .ZN(n1288) );
NAND3_X1 U1080 ( .A1(n1378), .A2(n1379), .A3(KEYINPUT57), .ZN(n1366) );
NAND2_X1 U1081 ( .A1(n1380), .A2(n1266), .ZN(n1379) );
NAND2_X1 U1082 ( .A1(n1157), .A2(n1381), .ZN(n1380) );
NAND2_X1 U1083 ( .A1(G125), .A2(n1159), .ZN(n1381) );
INV_X1 U1084 ( .A(n1382), .ZN(n1157) );
NAND2_X1 U1085 ( .A1(G146), .A2(n1383), .ZN(n1378) );
XNOR2_X1 U1086 ( .A(G125), .B(G140), .ZN(n1383) );
NAND2_X1 U1087 ( .A1(KEYINPUT8), .A2(n1194), .ZN(n1359) );
INV_X1 U1088 ( .A(G475), .ZN(n1194) );
INV_X1 U1089 ( .A(n1258), .ZN(n1272) );
XOR2_X1 U1090 ( .A(n1135), .B(n1137), .Z(n1258) );
INV_X1 U1091 ( .A(G478), .ZN(n1137) );
NOR2_X1 U1092 ( .A1(n1188), .A2(G902), .ZN(n1135) );
XNOR2_X1 U1093 ( .A(n1384), .B(n1385), .ZN(n1188) );
AND2_X1 U1094 ( .A1(n1386), .A2(G217), .ZN(n1385) );
NAND2_X1 U1095 ( .A1(n1387), .A2(n1388), .ZN(n1384) );
NAND2_X1 U1096 ( .A1(n1389), .A2(n1390), .ZN(n1388) );
XOR2_X1 U1097 ( .A(KEYINPUT53), .B(n1391), .Z(n1387) );
NOR2_X1 U1098 ( .A1(n1389), .A2(n1390), .ZN(n1391) );
XOR2_X1 U1099 ( .A(n1392), .B(n1393), .Z(n1390) );
XNOR2_X1 U1100 ( .A(n1071), .B(n1394), .ZN(n1393) );
NOR2_X1 U1101 ( .A1(G116), .A2(KEYINPUT43), .ZN(n1394) );
INV_X1 U1102 ( .A(G107), .ZN(n1071) );
XNOR2_X1 U1103 ( .A(G122), .B(KEYINPUT45), .ZN(n1392) );
XNOR2_X1 U1104 ( .A(G128), .B(n1395), .ZN(n1389) );
XNOR2_X1 U1105 ( .A(G143), .B(n1276), .ZN(n1395) );
INV_X1 U1106 ( .A(G134), .ZN(n1276) );
XNOR2_X1 U1107 ( .A(n1126), .B(KEYINPUT44), .ZN(n1094) );
XOR2_X1 U1108 ( .A(n1396), .B(n1183), .Z(n1126) );
NAND2_X1 U1109 ( .A1(G217), .A2(n1317), .ZN(n1183) );
NAND2_X1 U1110 ( .A1(n1397), .A2(n1232), .ZN(n1317) );
XNOR2_X1 U1111 ( .A(G234), .B(KEYINPUT5), .ZN(n1397) );
NAND2_X1 U1112 ( .A1(n1181), .A2(n1232), .ZN(n1396) );
INV_X1 U1113 ( .A(G902), .ZN(n1232) );
XNOR2_X1 U1114 ( .A(n1398), .B(n1399), .ZN(n1181) );
XOR2_X1 U1115 ( .A(n1400), .B(n1401), .Z(n1399) );
XNOR2_X1 U1116 ( .A(G110), .B(n1402), .ZN(n1401) );
NAND2_X1 U1117 ( .A1(n1403), .A2(KEYINPUT38), .ZN(n1402) );
XNOR2_X1 U1118 ( .A(G128), .B(G119), .ZN(n1403) );
NOR2_X1 U1119 ( .A1(n1382), .A2(n1404), .ZN(n1400) );
XOR2_X1 U1120 ( .A(KEYINPUT6), .B(n1405), .Z(n1404) );
NOR2_X1 U1121 ( .A1(G140), .A2(n1406), .ZN(n1405) );
XNOR2_X1 U1122 ( .A(KEYINPUT55), .B(n1160), .ZN(n1406) );
INV_X1 U1123 ( .A(G125), .ZN(n1160) );
NOR2_X1 U1124 ( .A1(n1159), .A2(G125), .ZN(n1382) );
INV_X1 U1125 ( .A(G140), .ZN(n1159) );
XOR2_X1 U1126 ( .A(n1407), .B(n1335), .Z(n1398) );
XNOR2_X1 U1127 ( .A(G137), .B(n1266), .ZN(n1335) );
INV_X1 U1128 ( .A(G146), .ZN(n1266) );
NAND2_X1 U1129 ( .A1(n1386), .A2(G221), .ZN(n1407) );
AND2_X1 U1130 ( .A1(G234), .A2(n1106), .ZN(n1386) );
INV_X1 U1131 ( .A(G953), .ZN(n1106) );
endmodule


