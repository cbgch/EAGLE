//Key = 1111011000000111000000110111010101011100001010100000111001000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263;

AND3_X1 U711 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n960) );
XNOR2_X1 U712 ( .A(G107), .B(n961), .ZN(G9) );
NAND4_X1 U713 ( .A1(KEYINPUT23), .A2(n962), .A3(n963), .A4(n964), .ZN(n961) );
XOR2_X1 U714 ( .A(KEYINPUT12), .B(n965), .Z(n964) );
NOR2_X1 U715 ( .A1(n966), .A2(n967), .ZN(G75) );
NOR4_X1 U716 ( .A1(n968), .A2(n969), .A3(n970), .A4(n971), .ZN(n967) );
XNOR2_X1 U717 ( .A(KEYINPUT27), .B(n972), .ZN(n969) );
NAND3_X1 U718 ( .A1(n973), .A2(n974), .A3(n975), .ZN(n968) );
NAND4_X1 U719 ( .A1(n976), .A2(n977), .A3(n978), .A4(n979), .ZN(n975) );
NOR2_X1 U720 ( .A1(n980), .A2(n981), .ZN(n979) );
NAND2_X1 U721 ( .A1(n982), .A2(n983), .ZN(n977) );
NAND2_X1 U722 ( .A1(n984), .A2(n962), .ZN(n983) );
NAND4_X1 U723 ( .A1(n985), .A2(n986), .A3(n987), .A4(n988), .ZN(n976) );
NAND2_X1 U724 ( .A1(n989), .A2(n990), .ZN(n987) );
XOR2_X1 U725 ( .A(n991), .B(KEYINPUT14), .Z(n989) );
NAND3_X1 U726 ( .A1(n984), .A2(n992), .A3(n960), .ZN(n986) );
NAND2_X1 U727 ( .A1(n962), .A2(n993), .ZN(n985) );
NAND2_X1 U728 ( .A1(n994), .A2(n995), .ZN(n993) );
NAND2_X1 U729 ( .A1(n996), .A2(n997), .ZN(n995) );
NAND4_X1 U730 ( .A1(n962), .A2(n998), .A3(n984), .A4(n999), .ZN(n973) );
NOR3_X1 U731 ( .A1(n982), .A2(n1000), .A3(n1001), .ZN(n999) );
NOR2_X1 U732 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NOR2_X1 U733 ( .A1(n1004), .A2(n981), .ZN(n1002) );
NOR2_X1 U734 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NOR2_X1 U735 ( .A1(n980), .A2(n1007), .ZN(n1000) );
AND2_X1 U736 ( .A1(n1008), .A2(n978), .ZN(n1007) );
INV_X1 U737 ( .A(n1005), .ZN(n978) );
NAND2_X1 U738 ( .A1(n1005), .A2(n1006), .ZN(n998) );
INV_X1 U739 ( .A(KEYINPUT17), .ZN(n1006) );
NOR3_X1 U740 ( .A1(n971), .A2(G952), .A3(n1009), .ZN(n966) );
INV_X1 U741 ( .A(n974), .ZN(n1009) );
NAND2_X1 U742 ( .A1(n1010), .A2(n1011), .ZN(n974) );
NOR4_X1 U743 ( .A1(n980), .A2(n1012), .A3(n1013), .A4(n1014), .ZN(n1011) );
XOR2_X1 U744 ( .A(n1015), .B(n1016), .Z(n1014) );
XNOR2_X1 U745 ( .A(n1017), .B(KEYINPUT62), .ZN(n1015) );
NOR2_X1 U746 ( .A1(n1018), .A2(n1019), .ZN(n1012) );
NOR4_X1 U747 ( .A1(n1020), .A2(n1021), .A3(n991), .A4(n1022), .ZN(n1010) );
XOR2_X1 U748 ( .A(G469), .B(n1023), .Z(n1022) );
NOR2_X1 U749 ( .A1(KEYINPUT10), .A2(n1024), .ZN(n1023) );
XOR2_X1 U750 ( .A(n1025), .B(KEYINPUT44), .Z(n1020) );
INV_X1 U751 ( .A(n1026), .ZN(n971) );
NAND3_X1 U752 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(G72) );
NAND2_X1 U753 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
INV_X1 U754 ( .A(KEYINPUT0), .ZN(n1031) );
OR2_X1 U755 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NAND3_X1 U756 ( .A1(KEYINPUT0), .A2(n1034), .A3(n1035), .ZN(n1028) );
NAND2_X1 U757 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NAND2_X1 U758 ( .A1(G953), .A2(n1038), .ZN(n1037) );
INV_X1 U759 ( .A(n1039), .ZN(n1036) );
NAND2_X1 U760 ( .A1(n1033), .A2(n1032), .ZN(n1027) );
NAND2_X1 U761 ( .A1(G953), .A2(n1040), .ZN(n1032) );
NAND2_X1 U762 ( .A1(G900), .A2(G227), .ZN(n1040) );
INV_X1 U763 ( .A(n1035), .ZN(n1033) );
XOR2_X1 U764 ( .A(n1041), .B(n1042), .Z(n1035) );
NOR3_X1 U765 ( .A1(n1043), .A2(n1039), .A3(n1044), .ZN(n1042) );
NOR2_X1 U766 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
XOR2_X1 U767 ( .A(n1047), .B(KEYINPUT2), .Z(n1043) );
NAND2_X1 U768 ( .A1(n1045), .A2(n1048), .ZN(n1047) );
XOR2_X1 U769 ( .A(KEYINPUT55), .B(n1046), .Z(n1048) );
XNOR2_X1 U770 ( .A(n1049), .B(n1050), .ZN(n1046) );
XOR2_X1 U771 ( .A(n1051), .B(G131), .Z(n1049) );
NAND2_X1 U772 ( .A1(KEYINPUT26), .A2(n1052), .ZN(n1051) );
NAND2_X1 U773 ( .A1(n1053), .A2(n970), .ZN(n1041) );
XOR2_X1 U774 ( .A(n1054), .B(n1055), .Z(G69) );
XOR2_X1 U775 ( .A(n1056), .B(n1057), .Z(n1055) );
NAND2_X1 U776 ( .A1(KEYINPUT25), .A2(n1058), .ZN(n1057) );
NAND2_X1 U777 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U778 ( .A1(G953), .A2(n1061), .ZN(n1060) );
XOR2_X1 U779 ( .A(n1062), .B(n1063), .Z(n1059) );
XNOR2_X1 U780 ( .A(n1064), .B(n1065), .ZN(n1062) );
NOR2_X1 U781 ( .A1(KEYINPUT34), .A2(n1066), .ZN(n1065) );
XOR2_X1 U782 ( .A(n1067), .B(G113), .Z(n1066) );
NAND2_X1 U783 ( .A1(n1053), .A2(n972), .ZN(n1056) );
NAND2_X1 U784 ( .A1(G953), .A2(n1068), .ZN(n1054) );
NAND2_X1 U785 ( .A1(G898), .A2(G224), .ZN(n1068) );
NOR2_X1 U786 ( .A1(n1069), .A2(n1070), .ZN(G66) );
NOR3_X1 U787 ( .A1(n1071), .A2(n1017), .A3(n1072), .ZN(n1070) );
NOR2_X1 U788 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U789 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NOR2_X1 U790 ( .A1(n972), .A2(n970), .ZN(n1075) );
XOR2_X1 U791 ( .A(n1077), .B(KEYINPUT46), .Z(n1071) );
NAND3_X1 U792 ( .A1(n1016), .A2(n1074), .A3(n1078), .ZN(n1077) );
NOR2_X1 U793 ( .A1(n1069), .A2(n1079), .ZN(G63) );
XOR2_X1 U794 ( .A(n1080), .B(n1081), .Z(n1079) );
AND2_X1 U795 ( .A1(G478), .A2(n1078), .ZN(n1080) );
NOR2_X1 U796 ( .A1(n1069), .A2(n1082), .ZN(G60) );
XNOR2_X1 U797 ( .A(n1083), .B(n1084), .ZN(n1082) );
AND2_X1 U798 ( .A1(G475), .A2(n1078), .ZN(n1084) );
XNOR2_X1 U799 ( .A(G104), .B(n1085), .ZN(G6) );
NAND3_X1 U800 ( .A1(n1086), .A2(n963), .A3(n1087), .ZN(n1085) );
XNOR2_X1 U801 ( .A(n962), .B(KEYINPUT6), .ZN(n1087) );
NOR2_X1 U802 ( .A1(n1069), .A2(n1088), .ZN(G57) );
XOR2_X1 U803 ( .A(n1089), .B(n1090), .Z(n1088) );
XNOR2_X1 U804 ( .A(n1091), .B(n1092), .ZN(n1090) );
NOR2_X1 U805 ( .A1(KEYINPUT4), .A2(n1093), .ZN(n1092) );
NOR3_X1 U806 ( .A1(n1094), .A2(KEYINPUT7), .A3(n1019), .ZN(n1091) );
NOR2_X1 U807 ( .A1(n1069), .A2(n1095), .ZN(G54) );
XOR2_X1 U808 ( .A(n1096), .B(n1097), .Z(n1095) );
XOR2_X1 U809 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND2_X1 U810 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NAND2_X1 U811 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U812 ( .A(KEYINPUT47), .B(n1104), .Z(n1102) );
NAND2_X1 U813 ( .A1(n1105), .A2(n1106), .ZN(n1100) );
INV_X1 U814 ( .A(n1103), .ZN(n1106) );
XNOR2_X1 U815 ( .A(G110), .B(G140), .ZN(n1103) );
XNOR2_X1 U816 ( .A(n1104), .B(n1107), .ZN(n1105) );
XNOR2_X1 U817 ( .A(KEYINPUT36), .B(KEYINPUT19), .ZN(n1107) );
XOR2_X1 U818 ( .A(n1108), .B(n1109), .Z(n1096) );
NOR2_X1 U819 ( .A1(n1110), .A2(KEYINPUT51), .ZN(n1109) );
AND2_X1 U820 ( .A1(G469), .A2(n1078), .ZN(n1110) );
INV_X1 U821 ( .A(n1094), .ZN(n1078) );
XOR2_X1 U822 ( .A(n1111), .B(KEYINPUT9), .Z(n1108) );
NAND2_X1 U823 ( .A1(n1112), .A2(KEYINPUT35), .ZN(n1111) );
XNOR2_X1 U824 ( .A(n1052), .B(n1113), .ZN(n1112) );
XNOR2_X1 U825 ( .A(n1114), .B(KEYINPUT40), .ZN(n1052) );
NOR2_X1 U826 ( .A1(n1115), .A2(n1116), .ZN(G51) );
XOR2_X1 U827 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U828 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U829 ( .A1(KEYINPUT33), .A2(n1121), .ZN(n1119) );
XNOR2_X1 U830 ( .A(n1122), .B(n1123), .ZN(n1117) );
NOR2_X1 U831 ( .A1(n1124), .A2(n1094), .ZN(n1123) );
NAND2_X1 U832 ( .A1(G902), .A2(n1125), .ZN(n1094) );
OR2_X1 U833 ( .A1(n970), .A2(n972), .ZN(n1125) );
NAND4_X1 U834 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n972) );
AND4_X1 U835 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1129) );
NAND3_X1 U836 ( .A1(n963), .A2(n1008), .A3(n962), .ZN(n1128) );
NAND2_X1 U837 ( .A1(n1134), .A2(n1135), .ZN(n1008) );
NAND4_X1 U838 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n970) );
NOR4_X1 U839 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1139) );
NOR2_X1 U840 ( .A1(n1144), .A2(n1145), .ZN(n1138) );
NOR2_X1 U841 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NOR2_X1 U842 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
NOR2_X1 U843 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XOR2_X1 U844 ( .A(n1134), .B(KEYINPUT49), .Z(n1150) );
NOR3_X1 U845 ( .A1(n1152), .A2(KEYINPUT54), .A3(n1153), .ZN(n1148) );
NAND2_X1 U846 ( .A1(KEYINPUT54), .A2(n1154), .ZN(n1137) );
OR2_X1 U847 ( .A1(n1155), .A2(n994), .ZN(n1136) );
XOR2_X1 U848 ( .A(n1156), .B(KEYINPUT50), .Z(n1115) );
NAND2_X1 U849 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND2_X1 U850 ( .A1(n1069), .A2(n1159), .ZN(n1158) );
INV_X1 U851 ( .A(KEYINPUT18), .ZN(n1159) );
NOR2_X1 U852 ( .A1(n1160), .A2(n1053), .ZN(n1069) );
NAND3_X1 U853 ( .A1(G953), .A2(n1160), .A3(KEYINPUT18), .ZN(n1157) );
XOR2_X1 U854 ( .A(G952), .B(KEYINPUT63), .Z(n1160) );
XNOR2_X1 U855 ( .A(G146), .B(n1161), .ZN(G48) );
NOR2_X1 U856 ( .A1(KEYINPUT32), .A2(n1162), .ZN(n1161) );
NOR4_X1 U857 ( .A1(n1163), .A2(n994), .A3(n980), .A4(n988), .ZN(n1162) );
INV_X1 U858 ( .A(n1003), .ZN(n980) );
NAND3_X1 U859 ( .A1(n1086), .A2(n1164), .A3(n1165), .ZN(n1163) );
XOR2_X1 U860 ( .A(n1166), .B(KEYINPUT16), .Z(n1165) );
XOR2_X1 U861 ( .A(G143), .B(n1144), .Z(G45) );
NOR4_X1 U862 ( .A1(n1167), .A2(n1151), .A3(n1168), .A4(n1169), .ZN(n1144) );
XOR2_X1 U863 ( .A(G140), .B(n1170), .Z(G42) );
NOR2_X1 U864 ( .A1(KEYINPUT11), .A2(n1171), .ZN(n1170) );
INV_X1 U865 ( .A(n1143), .ZN(n1171) );
NOR2_X1 U866 ( .A1(n1172), .A2(n1152), .ZN(n1143) );
XOR2_X1 U867 ( .A(n1173), .B(n1154), .Z(G39) );
NOR3_X1 U868 ( .A1(n1152), .A2(n1147), .A3(n981), .ZN(n1154) );
XNOR2_X1 U869 ( .A(G137), .B(KEYINPUT29), .ZN(n1173) );
XOR2_X1 U870 ( .A(G134), .B(n1142), .Z(G36) );
NOR3_X1 U871 ( .A1(n1152), .A2(n1135), .A3(n1167), .ZN(n1142) );
XOR2_X1 U872 ( .A(G131), .B(n1141), .Z(G33) );
NOR3_X1 U873 ( .A1(n1134), .A2(n1152), .A3(n1167), .ZN(n1141) );
INV_X1 U874 ( .A(n990), .ZN(n1167) );
NAND4_X1 U875 ( .A1(n984), .A2(n982), .A3(n1166), .A4(n1003), .ZN(n1152) );
INV_X1 U876 ( .A(n991), .ZN(n984) );
NAND2_X1 U877 ( .A1(n997), .A2(n1174), .ZN(n991) );
XOR2_X1 U878 ( .A(G128), .B(n1140), .Z(G30) );
NOR3_X1 U879 ( .A1(n1147), .A2(n1135), .A3(n1151), .ZN(n1140) );
NAND4_X1 U880 ( .A1(n1175), .A2(n982), .A3(n1166), .A4(n1003), .ZN(n1151) );
XNOR2_X1 U881 ( .A(G101), .B(n1126), .ZN(G3) );
NAND3_X1 U882 ( .A1(n990), .A2(n963), .A3(n1153), .ZN(n1126) );
XOR2_X1 U883 ( .A(G125), .B(n1176), .Z(G27) );
NOR2_X1 U884 ( .A1(n1177), .A2(n994), .ZN(n1176) );
INV_X1 U885 ( .A(n1175), .ZN(n994) );
XOR2_X1 U886 ( .A(n1155), .B(KEYINPUT48), .Z(n1177) );
NAND4_X1 U887 ( .A1(n988), .A2(n1178), .A3(n1166), .A4(n1003), .ZN(n1155) );
NAND2_X1 U888 ( .A1(n1005), .A2(n1179), .ZN(n1166) );
NAND3_X1 U889 ( .A1(G902), .A2(n1180), .A3(n1039), .ZN(n1179) );
NOR2_X1 U890 ( .A1(n1053), .A2(G900), .ZN(n1039) );
INV_X1 U891 ( .A(n1172), .ZN(n1178) );
NAND3_X1 U892 ( .A1(n960), .A2(n992), .A3(n1086), .ZN(n1172) );
XNOR2_X1 U893 ( .A(n1127), .B(n1181), .ZN(G24) );
NOR2_X1 U894 ( .A1(KEYINPUT59), .A2(n1182), .ZN(n1181) );
INV_X1 U895 ( .A(G122), .ZN(n1182) );
NAND4_X1 U896 ( .A1(n1183), .A2(n962), .A3(n1013), .A4(n1021), .ZN(n1127) );
NOR2_X1 U897 ( .A1(n1184), .A2(n960), .ZN(n962) );
XOR2_X1 U898 ( .A(n1185), .B(n1133), .Z(G21) );
NAND3_X1 U899 ( .A1(n1153), .A2(n1164), .A3(n1183), .ZN(n1133) );
INV_X1 U900 ( .A(n1147), .ZN(n1164) );
NAND2_X1 U901 ( .A1(n960), .A2(n1184), .ZN(n1147) );
XNOR2_X1 U902 ( .A(G116), .B(n1132), .ZN(G18) );
NAND3_X1 U903 ( .A1(n990), .A2(n965), .A3(n1183), .ZN(n1132) );
INV_X1 U904 ( .A(n1135), .ZN(n965) );
NAND2_X1 U905 ( .A1(n1169), .A2(n1013), .ZN(n1135) );
XNOR2_X1 U906 ( .A(G113), .B(n1131), .ZN(G15) );
NAND3_X1 U907 ( .A1(n990), .A2(n1086), .A3(n1183), .ZN(n1131) );
AND2_X1 U908 ( .A1(n988), .A2(n1186), .ZN(n1183) );
INV_X1 U909 ( .A(n1134), .ZN(n1086) );
NAND2_X1 U910 ( .A1(n1168), .A2(n1021), .ZN(n1134) );
INV_X1 U911 ( .A(n1169), .ZN(n1021) );
NOR2_X1 U912 ( .A1(n992), .A2(n960), .ZN(n990) );
XOR2_X1 U913 ( .A(n1130), .B(n1187), .Z(G12) );
XNOR2_X1 U914 ( .A(G110), .B(KEYINPUT28), .ZN(n1187) );
NAND4_X1 U915 ( .A1(n1153), .A2(n960), .A3(n963), .A4(n992), .ZN(n1130) );
INV_X1 U916 ( .A(n1184), .ZN(n992) );
NAND2_X1 U917 ( .A1(n1025), .A2(n1188), .ZN(n1184) );
NAND2_X1 U918 ( .A1(G472), .A2(n1189), .ZN(n1188) );
NAND2_X1 U919 ( .A1(n1018), .A2(n1019), .ZN(n1025) );
INV_X1 U920 ( .A(G472), .ZN(n1019) );
INV_X1 U921 ( .A(n1189), .ZN(n1018) );
NAND2_X1 U922 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
XOR2_X1 U923 ( .A(n1093), .B(n1192), .Z(n1190) );
INV_X1 U924 ( .A(n1089), .ZN(n1192) );
XOR2_X1 U925 ( .A(n1193), .B(n1194), .Z(n1089) );
XOR2_X1 U926 ( .A(n1195), .B(G101), .Z(n1193) );
NAND3_X1 U927 ( .A1(n1196), .A2(n1053), .A3(G210), .ZN(n1195) );
XOR2_X1 U928 ( .A(KEYINPUT57), .B(G237), .Z(n1196) );
XOR2_X1 U929 ( .A(n1197), .B(n1198), .Z(n1093) );
XOR2_X1 U930 ( .A(G113), .B(n1199), .Z(n1198) );
NOR2_X1 U931 ( .A1(G116), .A2(KEYINPUT56), .ZN(n1199) );
XOR2_X1 U932 ( .A(n1185), .B(KEYINPUT20), .Z(n1197) );
AND2_X1 U933 ( .A1(n1186), .A2(n982), .ZN(n963) );
INV_X1 U934 ( .A(n988), .ZN(n982) );
XOR2_X1 U935 ( .A(n1024), .B(G469), .Z(n988) );
NAND2_X1 U936 ( .A1(n1200), .A2(n1191), .ZN(n1024) );
XOR2_X1 U937 ( .A(n1201), .B(n1202), .Z(n1200) );
XOR2_X1 U938 ( .A(n1203), .B(n1204), .Z(n1202) );
XOR2_X1 U939 ( .A(KEYINPUT40), .B(G140), .Z(n1204) );
NOR2_X1 U940 ( .A1(G110), .A2(KEYINPUT38), .ZN(n1203) );
XOR2_X1 U941 ( .A(n1205), .B(n1194), .Z(n1201) );
XNOR2_X1 U942 ( .A(n1114), .B(n1099), .ZN(n1194) );
XOR2_X1 U943 ( .A(G131), .B(n1206), .Z(n1099) );
NOR2_X1 U944 ( .A1(KEYINPUT58), .A2(n1207), .ZN(n1206) );
XNOR2_X1 U945 ( .A(n1050), .B(KEYINPUT45), .ZN(n1207) );
XOR2_X1 U946 ( .A(G134), .B(G137), .Z(n1050) );
XNOR2_X1 U947 ( .A(n1113), .B(n1104), .ZN(n1205) );
NOR2_X1 U948 ( .A1(n1038), .A2(G953), .ZN(n1104) );
INV_X1 U949 ( .A(G227), .ZN(n1038) );
XOR2_X1 U950 ( .A(G104), .B(n1208), .Z(n1113) );
AND3_X1 U951 ( .A1(n1209), .A2(n1003), .A3(n1175), .ZN(n1186) );
NOR2_X1 U952 ( .A1(n997), .A2(n996), .ZN(n1175) );
INV_X1 U953 ( .A(n1174), .ZN(n996) );
NAND2_X1 U954 ( .A1(G214), .A2(n1210), .ZN(n1174) );
XNOR2_X1 U955 ( .A(n1211), .B(n1124), .ZN(n997) );
NAND2_X1 U956 ( .A1(G210), .A2(n1210), .ZN(n1124) );
NAND2_X1 U957 ( .A1(n1212), .A2(n1213), .ZN(n1210) );
NAND2_X1 U958 ( .A1(n1214), .A2(n1191), .ZN(n1211) );
XOR2_X1 U959 ( .A(n1215), .B(n1120), .Z(n1214) );
XOR2_X1 U960 ( .A(n1216), .B(n1217), .Z(n1120) );
XOR2_X1 U961 ( .A(n1063), .B(n1218), .Z(n1217) );
INV_X1 U962 ( .A(n1067), .ZN(n1218) );
XOR2_X1 U963 ( .A(n1219), .B(G116), .Z(n1067) );
NAND2_X1 U964 ( .A1(KEYINPUT13), .A2(n1185), .ZN(n1219) );
INV_X1 U965 ( .A(G119), .ZN(n1185) );
XNOR2_X1 U966 ( .A(n1220), .B(n1208), .ZN(n1063) );
XOR2_X1 U967 ( .A(G101), .B(G107), .Z(n1208) );
XNOR2_X1 U968 ( .A(G110), .B(KEYINPUT37), .ZN(n1220) );
XOR2_X1 U969 ( .A(n1221), .B(KEYINPUT52), .Z(n1216) );
NAND2_X1 U970 ( .A1(n1222), .A2(n1223), .ZN(n1215) );
NAND2_X1 U971 ( .A1(n1121), .A2(n1122), .ZN(n1223) );
XOR2_X1 U972 ( .A(n1224), .B(KEYINPUT41), .Z(n1222) );
OR2_X1 U973 ( .A1(n1122), .A2(n1121), .ZN(n1224) );
XOR2_X1 U974 ( .A(n1114), .B(n1225), .Z(n1121) );
XOR2_X1 U975 ( .A(KEYINPUT61), .B(G125), .Z(n1225) );
XOR2_X1 U976 ( .A(n1226), .B(n1227), .Z(n1114) );
NAND2_X1 U977 ( .A1(G224), .A2(n1053), .ZN(n1122) );
NAND2_X1 U978 ( .A1(G221), .A2(n1228), .ZN(n1003) );
NAND2_X1 U979 ( .A1(n1005), .A2(n1229), .ZN(n1209) );
NAND4_X1 U980 ( .A1(G953), .A2(G902), .A3(n1180), .A4(n1061), .ZN(n1229) );
INV_X1 U981 ( .A(G898), .ZN(n1061) );
NAND3_X1 U982 ( .A1(n1026), .A2(n1180), .A3(G952), .ZN(n1005) );
NAND2_X1 U983 ( .A1(G237), .A2(G234), .ZN(n1180) );
XOR2_X1 U984 ( .A(n1053), .B(KEYINPUT39), .Z(n1026) );
NAND2_X1 U985 ( .A1(n1017), .A2(n1233), .ZN(n1232) );
OR3_X1 U986 ( .A1(n1233), .A2(n1017), .A3(KEYINPUT60), .ZN(n1231) );
NOR2_X1 U987 ( .A1(n1074), .A2(G902), .ZN(n1017) );
XNOR2_X1 U988 ( .A(n1234), .B(n1235), .ZN(n1074) );
XNOR2_X1 U989 ( .A(n1236), .B(n1237), .ZN(n1235) );
XOR2_X1 U990 ( .A(n1238), .B(n1239), .Z(n1237) );
NOR2_X1 U991 ( .A1(KEYINPUT43), .A2(n1240), .ZN(n1239) );
XOR2_X1 U992 ( .A(n1241), .B(G110), .Z(n1240) );
NAND2_X1 U993 ( .A1(KEYINPUT22), .A2(n1242), .ZN(n1241) );
XOR2_X1 U994 ( .A(G128), .B(G119), .Z(n1242) );
NAND2_X1 U995 ( .A1(G221), .A2(n1243), .ZN(n1238) );
XNOR2_X1 U996 ( .A(G137), .B(n1244), .ZN(n1234) );
XOR2_X1 U997 ( .A(KEYINPUT24), .B(G146), .Z(n1244) );
NAND2_X1 U998 ( .A1(KEYINPUT15), .A2(n1076), .ZN(n1233) );
NAND2_X1 U999 ( .A1(KEYINPUT60), .A2(n1016), .ZN(n1230) );
INV_X1 U1000 ( .A(n1076), .ZN(n1016) );
NAND2_X1 U1001 ( .A1(G217), .A2(n1228), .ZN(n1076) );
NAND2_X1 U1002 ( .A1(G234), .A2(n1245), .ZN(n1228) );
XOR2_X1 U1003 ( .A(KEYINPUT21), .B(n1212), .Z(n1245) );
XOR2_X1 U1004 ( .A(G902), .B(KEYINPUT42), .Z(n1212) );
INV_X1 U1005 ( .A(n981), .ZN(n1153) );
NAND2_X1 U1006 ( .A1(n1246), .A2(n1168), .ZN(n981) );
INV_X1 U1007 ( .A(n1013), .ZN(n1168) );
XOR2_X1 U1008 ( .A(n1247), .B(n1248), .Z(n1013) );
XOR2_X1 U1009 ( .A(KEYINPUT53), .B(G478), .Z(n1248) );
OR2_X1 U1010 ( .A1(n1081), .A2(G902), .ZN(n1247) );
XNOR2_X1 U1011 ( .A(n1249), .B(n1250), .ZN(n1081) );
XOR2_X1 U1012 ( .A(n1251), .B(n1252), .Z(n1250) );
NAND2_X1 U1013 ( .A1(n1243), .A2(G217), .ZN(n1252) );
AND2_X1 U1014 ( .A1(G234), .A2(n1053), .ZN(n1243) );
NAND2_X1 U1015 ( .A1(n1253), .A2(KEYINPUT3), .ZN(n1251) );
XNOR2_X1 U1016 ( .A(G107), .B(n1254), .ZN(n1253) );
XOR2_X1 U1017 ( .A(G122), .B(G116), .Z(n1254) );
XOR2_X1 U1018 ( .A(n1226), .B(n1255), .Z(n1249) );
XOR2_X1 U1019 ( .A(G143), .B(G134), .Z(n1255) );
INV_X1 U1020 ( .A(G128), .ZN(n1226) );
XOR2_X1 U1021 ( .A(n1169), .B(KEYINPUT30), .Z(n1246) );
XOR2_X1 U1022 ( .A(n1256), .B(G475), .Z(n1169) );
NAND2_X1 U1023 ( .A1(n1257), .A2(n1083), .ZN(n1256) );
XNOR2_X1 U1024 ( .A(n1258), .B(n1259), .ZN(n1083) );
XOR2_X1 U1025 ( .A(n1221), .B(n1260), .Z(n1259) );
XNOR2_X1 U1026 ( .A(n1261), .B(n1262), .ZN(n1260) );
NAND2_X1 U1027 ( .A1(KEYINPUT1), .A2(n1263), .ZN(n1262) );
INV_X1 U1028 ( .A(G131), .ZN(n1263) );
NAND4_X1 U1029 ( .A1(KEYINPUT5), .A2(G214), .A3(n1213), .A4(n1053), .ZN(n1261) );
INV_X1 U1030 ( .A(G953), .ZN(n1053) );
INV_X1 U1031 ( .A(G237), .ZN(n1213) );
XNOR2_X1 U1032 ( .A(G113), .B(n1064), .ZN(n1221) );
XOR2_X1 U1033 ( .A(G104), .B(G122), .Z(n1064) );
XNOR2_X1 U1034 ( .A(n1227), .B(n1236), .ZN(n1258) );
XNOR2_X1 U1035 ( .A(n1045), .B(KEYINPUT31), .ZN(n1236) );
XNOR2_X1 U1036 ( .A(G125), .B(G140), .ZN(n1045) );
XOR2_X1 U1037 ( .A(G143), .B(G146), .Z(n1227) );
XOR2_X1 U1038 ( .A(n1191), .B(KEYINPUT8), .Z(n1257) );
INV_X1 U1039 ( .A(G902), .ZN(n1191) );
endmodule


