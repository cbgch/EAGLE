//Key = 0010010011010000001101011001000011010000100001101011011011011101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;

XOR2_X1 U727 ( .A(n998), .B(n999), .Z(G9) );
XNOR2_X1 U728 ( .A(KEYINPUT38), .B(n1000), .ZN(n999) );
NOR3_X1 U729 ( .A1(n1001), .A2(KEYINPUT41), .A3(n1002), .ZN(n998) );
NOR2_X1 U730 ( .A1(n1003), .A2(n1004), .ZN(G75) );
NOR4_X1 U731 ( .A1(G953), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n1004) );
INV_X1 U732 ( .A(n1008), .ZN(n1007) );
NOR2_X1 U733 ( .A1(n1009), .A2(n1010), .ZN(n1006) );
NOR2_X1 U734 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR2_X1 U735 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NOR2_X1 U736 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U737 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NOR2_X1 U738 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR2_X1 U739 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U740 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U741 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U742 ( .A1(n1027), .A2(n1028), .ZN(n1019) );
NOR2_X1 U743 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
AND3_X1 U744 ( .A1(n1031), .A2(n1032), .A3(G221), .ZN(n1029) );
INV_X1 U745 ( .A(n1033), .ZN(n1031) );
NOR3_X1 U746 ( .A1(n1022), .A2(n1034), .A3(n1028), .ZN(n1015) );
NOR2_X1 U747 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR4_X1 U748 ( .A1(n1037), .A2(n1028), .A3(n1022), .A4(n1018), .ZN(n1011) );
INV_X1 U749 ( .A(n1038), .ZN(n1018) );
INV_X1 U750 ( .A(n1039), .ZN(n1028) );
NOR2_X1 U751 ( .A1(n1040), .A2(n1041), .ZN(n1037) );
NOR2_X1 U752 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR3_X1 U753 ( .A1(n1005), .A2(G953), .A3(G952), .ZN(n1003) );
AND4_X1 U754 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1005) );
NOR4_X1 U755 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1022), .ZN(n1047) );
XNOR2_X1 U756 ( .A(n1051), .B(KEYINPUT5), .ZN(n1050) );
XOR2_X1 U757 ( .A(n1052), .B(n1053), .Z(n1049) );
NAND2_X1 U758 ( .A1(KEYINPUT51), .A2(n1054), .ZN(n1052) );
XNOR2_X1 U759 ( .A(n1042), .B(KEYINPUT17), .ZN(n1046) );
XNOR2_X1 U760 ( .A(n1026), .B(KEYINPUT14), .ZN(n1045) );
XNOR2_X1 U761 ( .A(n1055), .B(n1056), .ZN(n1044) );
XNOR2_X1 U762 ( .A(n1057), .B(KEYINPUT4), .ZN(n1055) );
XOR2_X1 U763 ( .A(n1058), .B(n1059), .Z(G72) );
NAND2_X1 U764 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U765 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
XOR2_X1 U766 ( .A(n1064), .B(n1065), .Z(n1062) );
NAND3_X1 U767 ( .A1(n1065), .A2(G900), .A3(G953), .ZN(n1060) );
NOR3_X1 U768 ( .A1(n1066), .A2(n1067), .A3(KEYINPUT29), .ZN(n1065) );
NOR2_X1 U769 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U770 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U771 ( .A1(G140), .A2(n1072), .ZN(n1071) );
NOR2_X1 U772 ( .A1(n1073), .A2(n1074), .ZN(n1070) );
NOR2_X1 U773 ( .A1(n1075), .A2(n1076), .ZN(n1066) );
NOR2_X1 U774 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR2_X1 U775 ( .A1(n1073), .A2(n1072), .ZN(n1078) );
XOR2_X1 U776 ( .A(n1074), .B(KEYINPUT19), .Z(n1072) );
NOR2_X1 U777 ( .A1(G140), .A2(n1074), .ZN(n1077) );
XNOR2_X1 U778 ( .A(n1079), .B(n1080), .ZN(n1074) );
NAND2_X1 U779 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NAND3_X1 U780 ( .A1(KEYINPUT59), .A2(n1083), .A3(n1084), .ZN(n1082) );
XOR2_X1 U781 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U782 ( .A1(KEYINPUT46), .A2(G137), .ZN(n1085) );
NAND2_X1 U783 ( .A1(n1087), .A2(n1088), .ZN(n1081) );
NAND2_X1 U784 ( .A1(KEYINPUT59), .A2(n1083), .ZN(n1088) );
XOR2_X1 U785 ( .A(n1089), .B(n1086), .Z(n1087) );
NAND2_X1 U786 ( .A1(KEYINPUT46), .A2(n1090), .ZN(n1089) );
INV_X1 U787 ( .A(G137), .ZN(n1090) );
INV_X1 U788 ( .A(n1069), .ZN(n1075) );
NAND2_X1 U789 ( .A1(KEYINPUT11), .A2(G125), .ZN(n1069) );
NAND2_X1 U790 ( .A1(KEYINPUT54), .A2(n1091), .ZN(n1058) );
NAND2_X1 U791 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U792 ( .A1(G900), .A2(G227), .ZN(n1093) );
XOR2_X1 U793 ( .A(n1094), .B(n1095), .Z(G69) );
XOR2_X1 U794 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U795 ( .A1(n1092), .A2(n1098), .ZN(n1097) );
NAND2_X1 U796 ( .A1(G898), .A2(G224), .ZN(n1098) );
XNOR2_X1 U797 ( .A(KEYINPUT45), .B(G953), .ZN(n1092) );
NAND4_X1 U798 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1096) );
NAND3_X1 U799 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
NAND2_X1 U800 ( .A1(n1106), .A2(n1107), .ZN(n1101) );
NAND2_X1 U801 ( .A1(n1108), .A2(n1104), .ZN(n1107) );
XNOR2_X1 U802 ( .A(KEYINPUT18), .B(n1103), .ZN(n1108) );
NAND2_X1 U803 ( .A1(G953), .A2(n1109), .ZN(n1100) );
OR2_X1 U804 ( .A1(n1104), .A2(n1103), .ZN(n1099) );
XOR2_X1 U805 ( .A(n1110), .B(n1111), .Z(n1103) );
XOR2_X1 U806 ( .A(KEYINPUT62), .B(KEYINPUT33), .Z(n1111) );
INV_X1 U807 ( .A(KEYINPUT3), .ZN(n1104) );
AND2_X1 U808 ( .A1(n1112), .A2(n1063), .ZN(n1094) );
NOR2_X1 U809 ( .A1(n1113), .A2(n1114), .ZN(G66) );
NOR3_X1 U810 ( .A1(n1057), .A2(n1115), .A3(n1116), .ZN(n1114) );
NOR3_X1 U811 ( .A1(n1117), .A2(n1056), .A3(n1118), .ZN(n1116) );
INV_X1 U812 ( .A(n1119), .ZN(n1118) );
NOR2_X1 U813 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
NOR2_X1 U814 ( .A1(n1008), .A2(n1056), .ZN(n1120) );
NOR2_X1 U815 ( .A1(n1113), .A2(n1122), .ZN(G63) );
NOR3_X1 U816 ( .A1(n1053), .A2(n1123), .A3(n1124), .ZN(n1122) );
AND3_X1 U817 ( .A1(n1125), .A2(n1119), .A3(G478), .ZN(n1124) );
NOR2_X1 U818 ( .A1(n1126), .A2(n1125), .ZN(n1123) );
NOR2_X1 U819 ( .A1(n1008), .A2(n1054), .ZN(n1126) );
INV_X1 U820 ( .A(G478), .ZN(n1054) );
NOR2_X1 U821 ( .A1(n1113), .A2(n1127), .ZN(G60) );
XOR2_X1 U822 ( .A(n1128), .B(n1129), .Z(n1127) );
AND2_X1 U823 ( .A1(G475), .A2(n1119), .ZN(n1128) );
XOR2_X1 U824 ( .A(G104), .B(n1130), .Z(G6) );
NOR2_X1 U825 ( .A1(n1113), .A2(n1131), .ZN(G57) );
XOR2_X1 U826 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U827 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U828 ( .A1(KEYINPUT34), .A2(n1136), .ZN(n1135) );
AND2_X1 U829 ( .A1(G472), .A2(n1119), .ZN(n1134) );
NOR2_X1 U830 ( .A1(n1113), .A2(n1137), .ZN(G54) );
XOR2_X1 U831 ( .A(n1138), .B(n1139), .Z(n1137) );
AND2_X1 U832 ( .A1(G469), .A2(n1119), .ZN(n1139) );
NOR2_X1 U833 ( .A1(KEYINPUT16), .A2(n1140), .ZN(n1138) );
XOR2_X1 U834 ( .A(n1141), .B(n1142), .Z(n1140) );
XNOR2_X1 U835 ( .A(G140), .B(n1143), .ZN(n1142) );
NAND2_X1 U836 ( .A1(KEYINPUT60), .A2(G110), .ZN(n1143) );
XOR2_X1 U837 ( .A(n1144), .B(n1145), .Z(n1141) );
NOR2_X1 U838 ( .A1(KEYINPUT55), .A2(n1146), .ZN(n1145) );
NOR2_X1 U839 ( .A1(n1113), .A2(n1147), .ZN(G51) );
XOR2_X1 U840 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U841 ( .A(n1150), .B(n1151), .ZN(n1149) );
NAND3_X1 U842 ( .A1(n1119), .A2(n1152), .A3(KEYINPUT24), .ZN(n1151) );
NOR2_X1 U843 ( .A1(n1153), .A2(n1008), .ZN(n1119) );
NOR2_X1 U844 ( .A1(n1064), .A2(n1112), .ZN(n1008) );
NAND2_X1 U845 ( .A1(n1154), .A2(n1155), .ZN(n1112) );
NOR4_X1 U846 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1130), .ZN(n1155) );
NOR2_X1 U847 ( .A1(n1159), .A2(n1002), .ZN(n1130) );
NOR4_X1 U848 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1154) );
NOR2_X1 U849 ( .A1(n1002), .A2(n1001), .ZN(n1163) );
NAND3_X1 U850 ( .A1(n1164), .A2(n1165), .A3(n1039), .ZN(n1002) );
NOR2_X1 U851 ( .A1(n1166), .A2(n1167), .ZN(n1162) );
XOR2_X1 U852 ( .A(n1168), .B(KEYINPUT43), .Z(n1166) );
NAND4_X1 U853 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1064) );
AND3_X1 U854 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1172) );
NAND2_X1 U855 ( .A1(n1176), .A2(n1177), .ZN(n1171) );
NAND2_X1 U856 ( .A1(n1178), .A2(n1001), .ZN(n1177) );
XNOR2_X1 U857 ( .A(n1036), .B(KEYINPUT58), .ZN(n1178) );
INV_X1 U858 ( .A(n1179), .ZN(n1176) );
NAND2_X1 U859 ( .A1(n1024), .A2(n1180), .ZN(n1169) );
NAND2_X1 U860 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND4_X1 U861 ( .A1(n1183), .A2(n1164), .A3(n1051), .A4(n1184), .ZN(n1182) );
NAND3_X1 U862 ( .A1(n1185), .A2(n1186), .A3(n1035), .ZN(n1181) );
OR2_X1 U863 ( .A1(n1187), .A2(KEYINPUT36), .ZN(n1186) );
NAND2_X1 U864 ( .A1(KEYINPUT36), .A2(n1188), .ZN(n1185) );
NAND3_X1 U865 ( .A1(n1014), .A2(n1184), .A3(n1030), .ZN(n1188) );
INV_X1 U866 ( .A(n1189), .ZN(n1014) );
NAND2_X1 U867 ( .A1(n1190), .A2(KEYINPUT48), .ZN(n1150) );
XOR2_X1 U868 ( .A(n1191), .B(n1192), .Z(n1190) );
NOR2_X1 U869 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XOR2_X1 U870 ( .A(n1195), .B(KEYINPUT2), .Z(n1194) );
NAND2_X1 U871 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NOR2_X1 U872 ( .A1(n1198), .A2(n1196), .ZN(n1193) );
XOR2_X1 U873 ( .A(G125), .B(KEYINPUT30), .Z(n1196) );
XOR2_X1 U874 ( .A(n1197), .B(KEYINPUT25), .Z(n1198) );
NOR2_X1 U875 ( .A1(n1063), .A2(G952), .ZN(n1113) );
XNOR2_X1 U876 ( .A(n1199), .B(n1200), .ZN(G48) );
NOR3_X1 U877 ( .A1(n1179), .A2(KEYINPUT10), .A3(n1159), .ZN(n1200) );
XNOR2_X1 U878 ( .A(G143), .B(n1201), .ZN(G45) );
NAND4_X1 U879 ( .A1(n1202), .A2(n1024), .A3(n1203), .A4(n1164), .ZN(n1201) );
NOR2_X1 U880 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
XOR2_X1 U881 ( .A(n1184), .B(KEYINPUT1), .Z(n1202) );
XNOR2_X1 U882 ( .A(n1170), .B(n1206), .ZN(G42) );
XNOR2_X1 U883 ( .A(KEYINPUT44), .B(n1073), .ZN(n1206) );
NAND2_X1 U884 ( .A1(n1187), .A2(n1207), .ZN(n1170) );
XNOR2_X1 U885 ( .A(G137), .B(n1173), .ZN(G39) );
NAND4_X1 U886 ( .A1(n1038), .A2(n1187), .A3(n1026), .A4(n1208), .ZN(n1173) );
XNOR2_X1 U887 ( .A(G134), .B(n1209), .ZN(G36) );
NAND2_X1 U888 ( .A1(n1210), .A2(n1035), .ZN(n1209) );
XOR2_X1 U889 ( .A(n1175), .B(n1211), .Z(G33) );
XNOR2_X1 U890 ( .A(G131), .B(KEYINPUT49), .ZN(n1211) );
NAND2_X1 U891 ( .A1(n1210), .A2(n1036), .ZN(n1175) );
AND2_X1 U892 ( .A1(n1024), .A2(n1187), .ZN(n1210) );
AND3_X1 U893 ( .A1(n1030), .A2(n1184), .A3(n1189), .ZN(n1187) );
NOR2_X1 U894 ( .A1(n1042), .A2(n1048), .ZN(n1189) );
XOR2_X1 U895 ( .A(G128), .B(n1212), .Z(G30) );
NOR2_X1 U896 ( .A1(n1001), .A2(n1179), .ZN(n1212) );
NAND4_X1 U897 ( .A1(n1164), .A2(n1026), .A3(n1208), .A4(n1184), .ZN(n1179) );
INV_X1 U898 ( .A(n1035), .ZN(n1001) );
XOR2_X1 U899 ( .A(G101), .B(n1161), .Z(G3) );
AND4_X1 U900 ( .A1(n1038), .A2(n1024), .A3(n1164), .A4(n1165), .ZN(n1161) );
AND2_X1 U901 ( .A1(n1041), .A2(n1030), .ZN(n1164) );
XNOR2_X1 U902 ( .A(G125), .B(n1174), .ZN(G27) );
NAND4_X1 U903 ( .A1(n1207), .A2(n1213), .A3(n1041), .A4(n1184), .ZN(n1174) );
NAND2_X1 U904 ( .A1(n1214), .A2(n1215), .ZN(n1184) );
NAND4_X1 U905 ( .A1(G902), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1215) );
INV_X1 U906 ( .A(G900), .ZN(n1218) );
XNOR2_X1 U907 ( .A(KEYINPUT28), .B(n1063), .ZN(n1216) );
NOR3_X1 U908 ( .A1(n1026), .A2(n1025), .A3(n1159), .ZN(n1207) );
INV_X1 U909 ( .A(n1036), .ZN(n1159) );
XOR2_X1 U910 ( .A(G122), .B(n1160), .Z(G24) );
AND4_X1 U911 ( .A1(n1219), .A2(n1039), .A3(n1183), .A4(n1051), .ZN(n1160) );
NOR2_X1 U912 ( .A1(n1208), .A2(n1026), .ZN(n1039) );
XOR2_X1 U913 ( .A(G119), .B(n1158), .Z(G21) );
AND4_X1 U914 ( .A1(n1219), .A2(n1038), .A3(n1026), .A4(n1208), .ZN(n1158) );
XNOR2_X1 U915 ( .A(n1220), .B(n1157), .ZN(G18) );
AND3_X1 U916 ( .A1(n1024), .A2(n1035), .A3(n1219), .ZN(n1157) );
NOR2_X1 U917 ( .A1(n1051), .A2(n1205), .ZN(n1035) );
XOR2_X1 U918 ( .A(G113), .B(n1156), .Z(G15) );
AND3_X1 U919 ( .A1(n1024), .A2(n1036), .A3(n1219), .ZN(n1156) );
NOR3_X1 U920 ( .A1(n1167), .A2(n1221), .A3(n1022), .ZN(n1219) );
INV_X1 U921 ( .A(n1213), .ZN(n1022) );
NOR2_X1 U922 ( .A1(n1033), .A2(n1222), .ZN(n1213) );
AND2_X1 U923 ( .A1(G221), .A2(n1032), .ZN(n1222) );
NOR2_X1 U924 ( .A1(n1183), .A2(n1204), .ZN(n1036) );
INV_X1 U925 ( .A(n1051), .ZN(n1204) );
AND2_X1 U926 ( .A1(n1223), .A2(n1026), .ZN(n1024) );
XNOR2_X1 U927 ( .A(KEYINPUT22), .B(n1208), .ZN(n1223) );
XNOR2_X1 U928 ( .A(n1224), .B(n1225), .ZN(G12) );
NOR2_X1 U929 ( .A1(n1167), .A2(n1168), .ZN(n1225) );
NAND4_X1 U930 ( .A1(n1038), .A2(n1030), .A3(n1226), .A4(n1227), .ZN(n1168) );
INV_X1 U931 ( .A(n1026), .ZN(n1227) );
XNOR2_X1 U932 ( .A(n1228), .B(G472), .ZN(n1026) );
NAND2_X1 U933 ( .A1(n1229), .A2(n1153), .ZN(n1228) );
XNOR2_X1 U934 ( .A(n1230), .B(n1136), .ZN(n1229) );
XOR2_X1 U935 ( .A(n1231), .B(n1232), .Z(n1136) );
XNOR2_X1 U936 ( .A(G116), .B(G119), .ZN(n1231) );
XNOR2_X1 U937 ( .A(n1132), .B(KEYINPUT0), .ZN(n1230) );
XNOR2_X1 U938 ( .A(n1233), .B(n1234), .ZN(n1132) );
XNOR2_X1 U939 ( .A(G101), .B(n1197), .ZN(n1234) );
XOR2_X1 U940 ( .A(n1235), .B(n1236), .Z(n1233) );
AND2_X1 U941 ( .A1(n1237), .A2(G210), .ZN(n1236) );
NOR2_X1 U942 ( .A1(n1025), .A2(n1221), .ZN(n1226) );
INV_X1 U943 ( .A(n1165), .ZN(n1221) );
NAND2_X1 U944 ( .A1(n1238), .A2(n1214), .ZN(n1165) );
NAND2_X1 U945 ( .A1(n1239), .A2(n1063), .ZN(n1214) );
INV_X1 U946 ( .A(n1010), .ZN(n1239) );
NAND2_X1 U947 ( .A1(G952), .A2(n1217), .ZN(n1010) );
NAND4_X1 U948 ( .A1(n1217), .A2(n1109), .A3(G902), .A4(G953), .ZN(n1238) );
INV_X1 U949 ( .A(G898), .ZN(n1109) );
NAND2_X1 U950 ( .A1(G237), .A2(n1240), .ZN(n1217) );
INV_X1 U951 ( .A(n1208), .ZN(n1025) );
NAND2_X1 U952 ( .A1(n1241), .A2(n1242), .ZN(n1208) );
NAND2_X1 U953 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
INV_X1 U954 ( .A(n1057), .ZN(n1244) );
XNOR2_X1 U955 ( .A(KEYINPUT37), .B(n1056), .ZN(n1243) );
NAND2_X1 U956 ( .A1(n1245), .A2(n1057), .ZN(n1241) );
NOR2_X1 U957 ( .A1(n1121), .A2(G902), .ZN(n1057) );
INV_X1 U958 ( .A(n1117), .ZN(n1121) );
XNOR2_X1 U959 ( .A(n1246), .B(n1247), .ZN(n1117) );
XNOR2_X1 U960 ( .A(n1248), .B(n1249), .ZN(n1247) );
XOR2_X1 U961 ( .A(n1250), .B(n1251), .Z(n1249) );
NOR2_X1 U962 ( .A1(KEYINPUT7), .A2(n1252), .ZN(n1251) );
XNOR2_X1 U963 ( .A(n1073), .B(G125), .ZN(n1252) );
NAND2_X1 U964 ( .A1(G221), .A2(n1253), .ZN(n1250) );
XOR2_X1 U965 ( .A(n1254), .B(n1255), .Z(n1246) );
XNOR2_X1 U966 ( .A(n1199), .B(G137), .ZN(n1255) );
XNOR2_X1 U967 ( .A(G119), .B(G110), .ZN(n1254) );
XNOR2_X1 U968 ( .A(KEYINPUT9), .B(n1056), .ZN(n1245) );
NAND2_X1 U969 ( .A1(G217), .A2(n1032), .ZN(n1056) );
AND2_X1 U970 ( .A1(n1033), .A2(n1256), .ZN(n1030) );
NAND2_X1 U971 ( .A1(G221), .A2(n1032), .ZN(n1256) );
NAND2_X1 U972 ( .A1(n1240), .A2(n1153), .ZN(n1032) );
XOR2_X1 U973 ( .A(G234), .B(KEYINPUT13), .Z(n1240) );
XNOR2_X1 U974 ( .A(n1257), .B(G469), .ZN(n1033) );
NAND2_X1 U975 ( .A1(n1258), .A2(n1153), .ZN(n1257) );
XOR2_X1 U976 ( .A(n1259), .B(n1260), .Z(n1258) );
XNOR2_X1 U977 ( .A(n1144), .B(n1146), .ZN(n1260) );
XOR2_X1 U978 ( .A(n1235), .B(n1261), .Z(n1144) );
XNOR2_X1 U979 ( .A(n1262), .B(n1080), .ZN(n1261) );
XOR2_X1 U980 ( .A(n1248), .B(n1263), .Z(n1080) );
NOR2_X1 U981 ( .A1(KEYINPUT20), .A2(n1264), .ZN(n1263) );
XNOR2_X1 U982 ( .A(G143), .B(G146), .ZN(n1264) );
NAND2_X1 U983 ( .A1(G227), .A2(n1063), .ZN(n1262) );
XOR2_X1 U984 ( .A(n1265), .B(n1266), .Z(n1235) );
NOR2_X1 U985 ( .A1(KEYINPUT31), .A2(n1086), .ZN(n1266) );
XNOR2_X1 U986 ( .A(n1267), .B(KEYINPUT52), .ZN(n1086) );
INV_X1 U987 ( .A(G131), .ZN(n1267) );
XNOR2_X1 U988 ( .A(G134), .B(G137), .ZN(n1265) );
XNOR2_X1 U989 ( .A(n1268), .B(KEYINPUT26), .ZN(n1259) );
NAND3_X1 U990 ( .A1(n1269), .A2(n1270), .A3(KEYINPUT63), .ZN(n1268) );
NAND2_X1 U991 ( .A1(KEYINPUT23), .A2(n1271), .ZN(n1270) );
XNOR2_X1 U992 ( .A(G110), .B(G140), .ZN(n1271) );
OR3_X1 U993 ( .A1(n1224), .A2(G140), .A3(KEYINPUT23), .ZN(n1269) );
NOR2_X1 U994 ( .A1(n1051), .A2(n1183), .ZN(n1038) );
INV_X1 U995 ( .A(n1205), .ZN(n1183) );
XOR2_X1 U996 ( .A(n1053), .B(n1272), .Z(n1205) );
NOR2_X1 U997 ( .A1(G478), .A2(KEYINPUT42), .ZN(n1272) );
NOR2_X1 U998 ( .A1(n1125), .A2(G902), .ZN(n1053) );
XOR2_X1 U999 ( .A(n1273), .B(n1274), .Z(n1125) );
AND2_X1 U1000 ( .A1(n1253), .A2(G217), .ZN(n1274) );
AND2_X1 U1001 ( .A1(G234), .A2(n1063), .ZN(n1253) );
NAND2_X1 U1002 ( .A1(KEYINPUT21), .A2(n1275), .ZN(n1273) );
XOR2_X1 U1003 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U1004 ( .A(n1278), .B(n1279), .ZN(n1277) );
NAND2_X1 U1005 ( .A1(KEYINPUT56), .A2(n1280), .ZN(n1278) );
XNOR2_X1 U1006 ( .A(n1281), .B(n1282), .ZN(n1280) );
XNOR2_X1 U1007 ( .A(G143), .B(n1083), .ZN(n1282) );
INV_X1 U1008 ( .A(G134), .ZN(n1083) );
XNOR2_X1 U1009 ( .A(n1220), .B(n1283), .ZN(n1276) );
NOR2_X1 U1010 ( .A1(KEYINPUT6), .A2(n1000), .ZN(n1283) );
XNOR2_X1 U1011 ( .A(n1284), .B(G475), .ZN(n1051) );
OR2_X1 U1012 ( .A1(n1129), .A2(G902), .ZN(n1284) );
XNOR2_X1 U1013 ( .A(n1285), .B(n1286), .ZN(n1129) );
XOR2_X1 U1014 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U1015 ( .A(G113), .B(G104), .Z(n1288) );
XNOR2_X1 U1016 ( .A(n1199), .B(G125), .ZN(n1287) );
XNOR2_X1 U1017 ( .A(n1279), .B(n1289), .ZN(n1285) );
XNOR2_X1 U1018 ( .A(n1290), .B(n1291), .ZN(n1289) );
NOR2_X1 U1019 ( .A1(KEYINPUT47), .A2(n1073), .ZN(n1291) );
INV_X1 U1020 ( .A(G140), .ZN(n1073) );
NAND2_X1 U1021 ( .A1(KEYINPUT27), .A2(n1292), .ZN(n1290) );
XOR2_X1 U1022 ( .A(n1293), .B(n1294), .Z(n1292) );
XNOR2_X1 U1023 ( .A(G131), .B(G143), .ZN(n1294) );
NAND2_X1 U1024 ( .A1(G214), .A2(n1237), .ZN(n1293) );
NOR2_X1 U1025 ( .A1(G953), .A2(G237), .ZN(n1237) );
INV_X1 U1026 ( .A(n1041), .ZN(n1167) );
NOR2_X1 U1027 ( .A1(n1295), .A2(n1048), .ZN(n1041) );
INV_X1 U1028 ( .A(n1043), .ZN(n1048) );
NAND2_X1 U1029 ( .A1(G214), .A2(n1296), .ZN(n1043) );
INV_X1 U1030 ( .A(n1042), .ZN(n1295) );
XNOR2_X1 U1031 ( .A(n1297), .B(n1152), .ZN(n1042) );
AND2_X1 U1032 ( .A1(G210), .A2(n1296), .ZN(n1152) );
NAND2_X1 U1033 ( .A1(n1298), .A2(n1299), .ZN(n1296) );
INV_X1 U1034 ( .A(G237), .ZN(n1299) );
XNOR2_X1 U1035 ( .A(KEYINPUT40), .B(n1153), .ZN(n1298) );
NAND2_X1 U1036 ( .A1(n1300), .A2(n1301), .ZN(n1297) );
XOR2_X1 U1037 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U1038 ( .A(n1304), .B(n1191), .ZN(n1303) );
NAND2_X1 U1039 ( .A1(G224), .A2(n1063), .ZN(n1191) );
INV_X1 U1040 ( .A(G953), .ZN(n1063) );
NAND2_X1 U1041 ( .A1(KEYINPUT57), .A2(n1148), .ZN(n1304) );
XOR2_X1 U1042 ( .A(n1110), .B(n1305), .Z(n1148) );
XNOR2_X1 U1043 ( .A(KEYINPUT35), .B(n1105), .ZN(n1305) );
INV_X1 U1044 ( .A(n1106), .ZN(n1105) );
XOR2_X1 U1045 ( .A(G110), .B(n1279), .Z(n1106) );
XOR2_X1 U1046 ( .A(G122), .B(KEYINPUT32), .Z(n1279) );
XOR2_X1 U1047 ( .A(n1306), .B(n1232), .Z(n1110) );
XOR2_X1 U1048 ( .A(G113), .B(KEYINPUT12), .Z(n1232) );
XNOR2_X1 U1049 ( .A(n1307), .B(n1308), .ZN(n1306) );
INV_X1 U1050 ( .A(n1146), .ZN(n1308) );
XOR2_X1 U1051 ( .A(G101), .B(n1309), .Z(n1146) );
XNOR2_X1 U1052 ( .A(n1000), .B(G104), .ZN(n1309) );
INV_X1 U1053 ( .A(G107), .ZN(n1000) );
NAND2_X1 U1054 ( .A1(KEYINPUT8), .A2(n1310), .ZN(n1307) );
XNOR2_X1 U1055 ( .A(G119), .B(n1311), .ZN(n1310) );
NAND2_X1 U1056 ( .A1(KEYINPUT61), .A2(n1220), .ZN(n1311) );
INV_X1 U1057 ( .A(G116), .ZN(n1220) );
XOR2_X1 U1058 ( .A(n1197), .B(G125), .Z(n1302) );
NAND2_X1 U1059 ( .A1(n1312), .A2(n1313), .ZN(n1197) );
OR2_X1 U1060 ( .A1(n1314), .A2(n1281), .ZN(n1313) );
XOR2_X1 U1061 ( .A(n1315), .B(KEYINPUT15), .Z(n1312) );
NAND2_X1 U1062 ( .A1(n1281), .A2(n1314), .ZN(n1315) );
XOR2_X1 U1063 ( .A(G143), .B(n1316), .Z(n1314) );
NOR2_X1 U1064 ( .A1(KEYINPUT39), .A2(n1199), .ZN(n1316) );
INV_X1 U1065 ( .A(G146), .ZN(n1199) );
INV_X1 U1066 ( .A(n1248), .ZN(n1281) );
XOR2_X1 U1067 ( .A(G128), .B(KEYINPUT50), .Z(n1248) );
XNOR2_X1 U1068 ( .A(KEYINPUT53), .B(n1153), .ZN(n1300) );
INV_X1 U1069 ( .A(G902), .ZN(n1153) );
INV_X1 U1070 ( .A(G110), .ZN(n1224) );
endmodule


