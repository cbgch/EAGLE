//Key = 0101111010110000101001001001010110100000000010111110011100001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369;

XNOR2_X1 U759 ( .A(G107), .B(n1053), .ZN(G9) );
NAND3_X1 U760 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NOR2_X1 U761 ( .A1(n1057), .A2(n1058), .ZN(G75) );
XOR2_X1 U762 ( .A(KEYINPUT56), .B(n1059), .Z(n1058) );
AND3_X1 U763 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NOR4_X1 U764 ( .A1(n1063), .A2(n1064), .A3(n1062), .A4(n1065), .ZN(n1057) );
NAND4_X1 U765 ( .A1(n1066), .A2(n1067), .A3(n1060), .A4(n1061), .ZN(n1063) );
NAND4_X1 U766 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1060) );
NOR2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XNOR2_X1 U768 ( .A(KEYINPUT47), .B(n1074), .ZN(n1070) );
XOR2_X1 U769 ( .A(KEYINPUT35), .B(n1075), .Z(n1069) );
NOR4_X1 U770 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1075) );
XOR2_X1 U771 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U772 ( .A1(G469), .A2(KEYINPUT61), .ZN(n1081) );
NOR2_X1 U773 ( .A1(KEYINPUT28), .A2(n1082), .ZN(n1077) );
AND2_X1 U774 ( .A1(n1083), .A2(KEYINPUT28), .ZN(n1076) );
XOR2_X1 U775 ( .A(KEYINPUT42), .B(n1084), .Z(n1068) );
NOR3_X1 U776 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
NOR3_X1 U777 ( .A1(n1088), .A2(KEYINPUT9), .A3(n1089), .ZN(n1087) );
AND2_X1 U778 ( .A1(n1088), .A2(KEYINPUT9), .ZN(n1086) );
INV_X1 U779 ( .A(n1090), .ZN(n1085) );
NAND4_X1 U780 ( .A1(n1091), .A2(n1092), .A3(n1082), .A4(n1055), .ZN(n1067) );
XOR2_X1 U781 ( .A(n1093), .B(KEYINPUT31), .Z(n1091) );
NAND2_X1 U782 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND4_X1 U783 ( .A1(n1096), .A2(n1097), .A3(n1095), .A4(n1094), .ZN(n1066) );
INV_X1 U784 ( .A(KEYINPUT52), .ZN(n1094) );
NAND2_X1 U785 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND4_X1 U786 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1099) );
NAND2_X1 U787 ( .A1(n1078), .A2(n1104), .ZN(n1103) );
NAND2_X1 U788 ( .A1(n1092), .A2(n1082), .ZN(n1104) );
NAND4_X1 U789 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1102) );
NAND2_X1 U790 ( .A1(n1092), .A2(n1109), .ZN(n1107) );
NAND3_X1 U791 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1106) );
XNOR2_X1 U792 ( .A(n1092), .B(KEYINPUT16), .ZN(n1112) );
NAND2_X1 U793 ( .A1(n1082), .A2(n1113), .ZN(n1105) );
OR2_X1 U794 ( .A1(n1114), .A2(n1056), .ZN(n1113) );
NAND3_X1 U795 ( .A1(n1115), .A2(n1108), .A3(n1092), .ZN(n1098) );
NAND2_X1 U796 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U797 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XOR2_X1 U798 ( .A(KEYINPUT15), .B(n1082), .Z(n1119) );
NAND2_X1 U799 ( .A1(n1120), .A2(n1082), .ZN(n1116) );
XOR2_X1 U800 ( .A(n1121), .B(n1122), .Z(G72) );
XOR2_X1 U801 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U802 ( .A1(G953), .A2(n1125), .ZN(n1124) );
NAND2_X1 U803 ( .A1(G900), .A2(G227), .ZN(n1125) );
NAND3_X1 U804 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1123) );
XOR2_X1 U805 ( .A(n1129), .B(KEYINPUT20), .Z(n1128) );
NAND2_X1 U806 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XNOR2_X1 U807 ( .A(n1132), .B(n1133), .ZN(n1131) );
XNOR2_X1 U808 ( .A(n1134), .B(n1135), .ZN(n1130) );
NAND2_X1 U809 ( .A1(n1136), .A2(n1137), .ZN(n1127) );
XNOR2_X1 U810 ( .A(G125), .B(n1132), .ZN(n1137) );
NAND2_X1 U811 ( .A1(KEYINPUT46), .A2(n1138), .ZN(n1132) );
XNOR2_X1 U812 ( .A(n1135), .B(n1139), .ZN(n1136) );
INV_X1 U813 ( .A(n1134), .ZN(n1139) );
NAND2_X1 U814 ( .A1(G953), .A2(n1140), .ZN(n1126) );
AND2_X1 U815 ( .A1(n1064), .A2(n1061), .ZN(n1121) );
XOR2_X1 U816 ( .A(n1141), .B(n1142), .Z(G69) );
NAND2_X1 U817 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U818 ( .A1(G898), .A2(G224), .ZN(n1144) );
XNOR2_X1 U819 ( .A(KEYINPUT57), .B(n1061), .ZN(n1143) );
NAND3_X1 U820 ( .A1(n1145), .A2(n1146), .A3(KEYINPUT5), .ZN(n1141) );
NAND2_X1 U821 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
INV_X1 U822 ( .A(KEYINPUT37), .ZN(n1148) );
XNOR2_X1 U823 ( .A(n1149), .B(n1150), .ZN(n1147) );
NAND2_X1 U824 ( .A1(n1061), .A2(n1065), .ZN(n1149) );
NAND4_X1 U825 ( .A1(n1065), .A2(n1061), .A3(n1150), .A4(KEYINPUT37), .ZN(n1145) );
NAND3_X1 U826 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
XOR2_X1 U827 ( .A(KEYINPUT4), .B(n1154), .Z(n1153) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND2_X1 U829 ( .A1(n1155), .A2(n1156), .ZN(n1152) );
XOR2_X1 U830 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U831 ( .A1(KEYINPUT45), .A2(n1159), .ZN(n1157) );
NAND2_X1 U832 ( .A1(G953), .A2(n1160), .ZN(n1151) );
NOR2_X1 U833 ( .A1(n1161), .A2(n1162), .ZN(G66) );
XOR2_X1 U834 ( .A(n1163), .B(n1164), .Z(n1162) );
OR2_X1 U835 ( .A1(n1165), .A2(n1088), .ZN(n1163) );
NOR2_X1 U836 ( .A1(n1161), .A2(n1166), .ZN(G63) );
XOR2_X1 U837 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U838 ( .A1(n1169), .A2(KEYINPUT41), .ZN(n1167) );
AND2_X1 U839 ( .A1(G478), .A2(n1170), .ZN(n1169) );
NOR2_X1 U840 ( .A1(n1161), .A2(n1171), .ZN(G60) );
NOR2_X1 U841 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XOR2_X1 U842 ( .A(n1174), .B(KEYINPUT34), .Z(n1173) );
NAND2_X1 U843 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NOR2_X1 U844 ( .A1(n1175), .A2(n1176), .ZN(n1172) );
AND2_X1 U845 ( .A1(n1170), .A2(G475), .ZN(n1175) );
XNOR2_X1 U846 ( .A(n1177), .B(n1178), .ZN(G6) );
NOR2_X1 U847 ( .A1(G104), .A2(KEYINPUT12), .ZN(n1178) );
NOR2_X1 U848 ( .A1(n1179), .A2(n1180), .ZN(G57) );
XOR2_X1 U849 ( .A(n1181), .B(n1182), .Z(n1180) );
XNOR2_X1 U850 ( .A(n1183), .B(n1184), .ZN(n1182) );
NAND2_X1 U851 ( .A1(n1170), .A2(G472), .ZN(n1183) );
XNOR2_X1 U852 ( .A(G101), .B(n1185), .ZN(n1181) );
NOR2_X1 U853 ( .A1(KEYINPUT36), .A2(n1186), .ZN(n1185) );
XNOR2_X1 U854 ( .A(n1187), .B(n1188), .ZN(n1186) );
XNOR2_X1 U855 ( .A(n1189), .B(n1190), .ZN(n1187) );
NOR2_X1 U856 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U857 ( .A(KEYINPUT7), .B(KEYINPUT17), .Z(n1192) );
XNOR2_X1 U858 ( .A(n1161), .B(KEYINPUT54), .ZN(n1179) );
NOR2_X1 U859 ( .A1(n1161), .A2(n1193), .ZN(G54) );
XOR2_X1 U860 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U861 ( .A(n1196), .B(n1197), .Z(n1195) );
NAND2_X1 U862 ( .A1(n1170), .A2(G469), .ZN(n1197) );
NAND2_X1 U863 ( .A1(KEYINPUT50), .A2(n1198), .ZN(n1196) );
XNOR2_X1 U864 ( .A(n1199), .B(n1200), .ZN(n1198) );
NOR2_X1 U865 ( .A1(KEYINPUT13), .A2(n1201), .ZN(n1199) );
XOR2_X1 U866 ( .A(n1202), .B(n1203), .Z(n1194) );
NAND2_X1 U867 ( .A1(KEYINPUT10), .A2(n1204), .ZN(n1203) );
NOR2_X1 U868 ( .A1(n1161), .A2(n1205), .ZN(G51) );
XNOR2_X1 U869 ( .A(n1206), .B(n1207), .ZN(n1205) );
XOR2_X1 U870 ( .A(n1208), .B(n1209), .Z(n1206) );
NAND2_X1 U871 ( .A1(n1170), .A2(G210), .ZN(n1208) );
INV_X1 U872 ( .A(n1165), .ZN(n1170) );
NAND2_X1 U873 ( .A1(G902), .A2(n1210), .ZN(n1165) );
NAND2_X1 U874 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
INV_X1 U875 ( .A(n1065), .ZN(n1212) );
NAND4_X1 U876 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1065) );
NOR4_X1 U877 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1177), .ZN(n1216) );
AND3_X1 U878 ( .A1(n1054), .A2(n1055), .A3(n1114), .ZN(n1177) );
NOR2_X1 U879 ( .A1(n1220), .A2(n1221), .ZN(n1215) );
INV_X1 U880 ( .A(n1222), .ZN(n1220) );
NAND4_X1 U881 ( .A1(n1056), .A2(n1055), .A3(n1223), .A4(n1224), .ZN(n1213) );
OR2_X1 U882 ( .A1(n1054), .A2(KEYINPUT2), .ZN(n1224) );
NAND2_X1 U883 ( .A1(KEYINPUT2), .A2(n1225), .ZN(n1223) );
NAND3_X1 U884 ( .A1(n1095), .A2(n1083), .A3(n1226), .ZN(n1225) );
INV_X1 U885 ( .A(n1109), .ZN(n1083) );
NOR4_X1 U886 ( .A1(n1072), .A2(n1227), .A3(n1096), .A4(n1078), .ZN(n1055) );
XOR2_X1 U887 ( .A(n1064), .B(KEYINPUT27), .Z(n1211) );
NAND4_X1 U888 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1064) );
NOR4_X1 U889 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1231) );
NAND2_X1 U890 ( .A1(n1114), .A2(n1236), .ZN(n1230) );
NAND2_X1 U891 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NAND3_X1 U892 ( .A1(n1118), .A2(n1239), .A3(n1096), .ZN(n1238) );
AND2_X1 U893 ( .A1(n1240), .A2(n1062), .ZN(n1161) );
INV_X1 U894 ( .A(G952), .ZN(n1062) );
XNOR2_X1 U895 ( .A(G953), .B(KEYINPUT48), .ZN(n1240) );
XNOR2_X1 U896 ( .A(G146), .B(n1229), .ZN(G48) );
NAND3_X1 U897 ( .A1(n1241), .A2(n1242), .A3(n1114), .ZN(n1229) );
XNOR2_X1 U898 ( .A(G143), .B(n1228), .ZN(G45) );
NAND3_X1 U899 ( .A1(n1120), .A2(n1241), .A3(n1243), .ZN(n1228) );
XNOR2_X1 U900 ( .A(n1138), .B(n1235), .ZN(G42) );
AND3_X1 U901 ( .A1(n1118), .A2(n1244), .A3(n1114), .ZN(n1235) );
XNOR2_X1 U902 ( .A(n1245), .B(n1234), .ZN(G39) );
AND3_X1 U903 ( .A1(n1244), .A2(n1242), .A3(n1092), .ZN(n1234) );
XOR2_X1 U904 ( .A(G134), .B(n1233), .Z(G36) );
AND2_X1 U905 ( .A1(n1246), .A2(n1056), .ZN(n1233) );
XNOR2_X1 U906 ( .A(G131), .B(n1247), .ZN(G33) );
NAND2_X1 U907 ( .A1(n1248), .A2(n1246), .ZN(n1247) );
INV_X1 U908 ( .A(n1237), .ZN(n1246) );
NAND2_X1 U909 ( .A1(n1120), .A2(n1244), .ZN(n1237) );
AND4_X1 U910 ( .A1(n1082), .A2(n1249), .A3(n1250), .A4(n1108), .ZN(n1244) );
NOR2_X1 U911 ( .A1(n1251), .A2(n1110), .ZN(n1082) );
XNOR2_X1 U912 ( .A(n1114), .B(KEYINPUT44), .ZN(n1248) );
NAND2_X1 U913 ( .A1(n1252), .A2(n1253), .ZN(G30) );
NAND2_X1 U914 ( .A1(n1232), .A2(n1254), .ZN(n1253) );
XOR2_X1 U915 ( .A(KEYINPUT8), .B(n1255), .Z(n1252) );
NOR2_X1 U916 ( .A1(n1232), .A2(n1254), .ZN(n1255) );
AND3_X1 U917 ( .A1(n1242), .A2(n1056), .A3(n1241), .ZN(n1232) );
AND2_X1 U918 ( .A1(n1239), .A2(n1250), .ZN(n1241) );
XNOR2_X1 U919 ( .A(n1256), .B(n1219), .ZN(G3) );
AND2_X1 U920 ( .A1(n1257), .A2(n1120), .ZN(n1219) );
XNOR2_X1 U921 ( .A(G125), .B(n1258), .ZN(G27) );
NAND4_X1 U922 ( .A1(n1259), .A2(n1096), .A3(n1114), .A4(n1239), .ZN(n1258) );
AND3_X1 U923 ( .A1(n1109), .A2(n1108), .A3(n1249), .ZN(n1239) );
AND2_X1 U924 ( .A1(n1260), .A2(n1095), .ZN(n1249) );
NAND2_X1 U925 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
NAND3_X1 U926 ( .A1(G902), .A2(n1140), .A3(n1263), .ZN(n1262) );
XNOR2_X1 U927 ( .A(G953), .B(KEYINPUT49), .ZN(n1263) );
INV_X1 U928 ( .A(G900), .ZN(n1140) );
INV_X1 U929 ( .A(n1250), .ZN(n1096) );
XNOR2_X1 U930 ( .A(n1118), .B(KEYINPUT21), .ZN(n1259) );
XNOR2_X1 U931 ( .A(G122), .B(n1214), .ZN(G24) );
NAND4_X1 U932 ( .A1(n1264), .A2(n1243), .A3(n1100), .A4(n1101), .ZN(n1214) );
AND2_X1 U933 ( .A1(n1265), .A2(n1073), .ZN(n1243) );
XNOR2_X1 U934 ( .A(n1266), .B(KEYINPUT11), .ZN(n1265) );
XNOR2_X1 U935 ( .A(n1267), .B(n1221), .ZN(G21) );
AND3_X1 U936 ( .A1(n1092), .A2(n1242), .A3(n1264), .ZN(n1221) );
NOR2_X1 U937 ( .A1(n1100), .A2(n1101), .ZN(n1242) );
NAND2_X1 U938 ( .A1(n1268), .A2(n1269), .ZN(G18) );
NAND2_X1 U939 ( .A1(G116), .A2(n1222), .ZN(n1269) );
XOR2_X1 U940 ( .A(KEYINPUT1), .B(n1270), .Z(n1268) );
NOR2_X1 U941 ( .A1(G116), .A2(n1222), .ZN(n1270) );
NAND3_X1 U942 ( .A1(n1120), .A2(n1056), .A3(n1264), .ZN(n1222) );
NOR2_X1 U943 ( .A1(n1073), .A2(n1074), .ZN(n1056) );
XNOR2_X1 U944 ( .A(n1271), .B(n1218), .ZN(G15) );
AND3_X1 U945 ( .A1(n1114), .A2(n1120), .A3(n1264), .ZN(n1218) );
NOR3_X1 U946 ( .A1(n1272), .A2(n1078), .A3(n1250), .ZN(n1264) );
INV_X1 U947 ( .A(n1108), .ZN(n1078) );
NOR2_X1 U948 ( .A1(n1227), .A2(n1100), .ZN(n1120) );
INV_X1 U949 ( .A(n1072), .ZN(n1100) );
AND2_X1 U950 ( .A1(n1074), .A2(n1073), .ZN(n1114) );
INV_X1 U951 ( .A(n1266), .ZN(n1074) );
XNOR2_X1 U952 ( .A(n1273), .B(n1217), .ZN(G12) );
AND2_X1 U953 ( .A1(n1257), .A2(n1118), .ZN(n1217) );
NOR2_X1 U954 ( .A1(n1072), .A2(n1101), .ZN(n1118) );
INV_X1 U955 ( .A(n1227), .ZN(n1101) );
NAND3_X1 U956 ( .A1(n1274), .A2(n1275), .A3(n1090), .ZN(n1227) );
NAND2_X1 U957 ( .A1(n1089), .A2(n1088), .ZN(n1090) );
NAND2_X1 U958 ( .A1(KEYINPUT39), .A2(n1088), .ZN(n1275) );
OR3_X1 U959 ( .A1(n1089), .A2(KEYINPUT39), .A3(n1088), .ZN(n1274) );
NAND2_X1 U960 ( .A1(G217), .A2(n1276), .ZN(n1088) );
AND2_X1 U961 ( .A1(n1164), .A2(n1277), .ZN(n1089) );
XOR2_X1 U962 ( .A(n1278), .B(n1279), .Z(n1164) );
XNOR2_X1 U963 ( .A(n1273), .B(n1280), .ZN(n1279) );
XNOR2_X1 U964 ( .A(KEYINPUT38), .B(n1267), .ZN(n1280) );
XOR2_X1 U965 ( .A(n1281), .B(n1282), .Z(n1278) );
XOR2_X1 U966 ( .A(n1283), .B(n1284), .Z(n1281) );
NOR3_X1 U967 ( .A1(n1285), .A2(KEYINPUT63), .A3(n1286), .ZN(n1284) );
NOR4_X1 U968 ( .A1(G953), .A2(n1287), .A3(n1288), .A4(n1289), .ZN(n1286) );
XNOR2_X1 U969 ( .A(G137), .B(KEYINPUT59), .ZN(n1287) );
NOR2_X1 U970 ( .A1(n1290), .A2(G137), .ZN(n1285) );
NOR3_X1 U971 ( .A1(n1289), .A2(G953), .A3(n1288), .ZN(n1290) );
INV_X1 U972 ( .A(G234), .ZN(n1288) );
XOR2_X1 U973 ( .A(G221), .B(KEYINPUT18), .Z(n1289) );
NAND2_X1 U974 ( .A1(n1291), .A2(n1292), .ZN(n1283) );
NAND2_X1 U975 ( .A1(G140), .A2(n1133), .ZN(n1292) );
INV_X1 U976 ( .A(G125), .ZN(n1133) );
XOR2_X1 U977 ( .A(n1293), .B(KEYINPUT33), .Z(n1291) );
NAND2_X1 U978 ( .A1(G125), .A2(n1138), .ZN(n1293) );
XNOR2_X1 U979 ( .A(n1294), .B(G472), .ZN(n1072) );
NAND2_X1 U980 ( .A1(n1295), .A2(n1277), .ZN(n1294) );
XOR2_X1 U981 ( .A(n1296), .B(n1297), .Z(n1295) );
XNOR2_X1 U982 ( .A(n1200), .B(n1191), .ZN(n1297) );
XNOR2_X1 U983 ( .A(n1298), .B(n1299), .ZN(n1191) );
NOR2_X1 U984 ( .A1(KEYINPUT30), .A2(n1300), .ZN(n1299) );
XNOR2_X1 U985 ( .A(G113), .B(G119), .ZN(n1298) );
XOR2_X1 U986 ( .A(n1301), .B(n1302), .Z(n1296) );
XOR2_X1 U987 ( .A(n1184), .B(n1303), .Z(n1302) );
NOR2_X1 U988 ( .A1(KEYINPUT23), .A2(n1188), .ZN(n1303) );
NAND3_X1 U989 ( .A1(n1304), .A2(n1061), .A3(G210), .ZN(n1184) );
NAND2_X1 U990 ( .A1(KEYINPUT3), .A2(G101), .ZN(n1301) );
AND4_X1 U991 ( .A1(n1092), .A2(n1054), .A3(n1250), .A4(n1108), .ZN(n1257) );
NAND2_X1 U992 ( .A1(G221), .A2(n1276), .ZN(n1108) );
NAND2_X1 U993 ( .A1(G234), .A2(n1277), .ZN(n1276) );
XNOR2_X1 U994 ( .A(n1080), .B(G469), .ZN(n1250) );
NAND2_X1 U995 ( .A1(n1305), .A2(n1277), .ZN(n1080) );
XOR2_X1 U996 ( .A(n1306), .B(n1307), .Z(n1305) );
XNOR2_X1 U997 ( .A(n1202), .B(n1308), .ZN(n1307) );
NOR2_X1 U998 ( .A1(KEYINPUT22), .A2(n1309), .ZN(n1308) );
XNOR2_X1 U999 ( .A(n1204), .B(KEYINPUT26), .ZN(n1309) );
XNOR2_X1 U1000 ( .A(G110), .B(n1138), .ZN(n1204) );
INV_X1 U1001 ( .A(G140), .ZN(n1138) );
NAND2_X1 U1002 ( .A1(G227), .A2(n1061), .ZN(n1202) );
XNOR2_X1 U1003 ( .A(n1201), .B(n1200), .ZN(n1306) );
INV_X1 U1004 ( .A(n1189), .ZN(n1200) );
XOR2_X1 U1005 ( .A(n1135), .B(KEYINPUT25), .Z(n1189) );
XOR2_X1 U1006 ( .A(G131), .B(n1310), .Z(n1135) );
XNOR2_X1 U1007 ( .A(n1245), .B(G134), .ZN(n1310) );
INV_X1 U1008 ( .A(G137), .ZN(n1245) );
XOR2_X1 U1009 ( .A(n1311), .B(n1312), .Z(n1201) );
XOR2_X1 U1010 ( .A(KEYINPUT62), .B(n1313), .Z(n1312) );
NOR2_X1 U1011 ( .A1(G107), .A2(KEYINPUT40), .ZN(n1313) );
XNOR2_X1 U1012 ( .A(n1134), .B(n1314), .ZN(n1311) );
XOR2_X1 U1013 ( .A(G143), .B(n1282), .Z(n1134) );
XNOR2_X1 U1014 ( .A(n1254), .B(G146), .ZN(n1282) );
INV_X1 U1015 ( .A(n1272), .ZN(n1054) );
NAND3_X1 U1016 ( .A1(n1226), .A2(n1095), .A3(n1109), .ZN(n1272) );
NOR2_X1 U1017 ( .A1(n1111), .A2(n1110), .ZN(n1109) );
AND2_X1 U1018 ( .A1(G214), .A2(n1315), .ZN(n1110) );
NAND2_X1 U1019 ( .A1(n1277), .A2(n1304), .ZN(n1315) );
INV_X1 U1020 ( .A(n1251), .ZN(n1111) );
NAND3_X1 U1021 ( .A1(n1316), .A2(n1317), .A3(n1318), .ZN(n1251) );
NAND2_X1 U1022 ( .A1(G902), .A2(G210), .ZN(n1318) );
NAND3_X1 U1023 ( .A1(n1319), .A2(n1277), .A3(n1320), .ZN(n1317) );
OR2_X1 U1024 ( .A1(n1320), .A2(n1319), .ZN(n1316) );
AND2_X1 U1025 ( .A1(n1321), .A2(n1322), .ZN(n1319) );
NAND2_X1 U1026 ( .A1(n1323), .A2(n1209), .ZN(n1322) );
XOR2_X1 U1027 ( .A(KEYINPUT6), .B(n1324), .Z(n1321) );
NOR2_X1 U1028 ( .A1(n1209), .A2(n1323), .ZN(n1324) );
XNOR2_X1 U1029 ( .A(KEYINPUT51), .B(n1207), .ZN(n1323) );
XNOR2_X1 U1030 ( .A(n1325), .B(n1188), .ZN(n1207) );
XOR2_X1 U1031 ( .A(n1326), .B(n1327), .Z(n1188) );
XNOR2_X1 U1032 ( .A(n1328), .B(n1329), .ZN(n1327) );
NOR2_X1 U1033 ( .A1(G128), .A2(KEYINPUT14), .ZN(n1329) );
NAND2_X1 U1034 ( .A1(KEYINPUT32), .A2(G146), .ZN(n1326) );
XNOR2_X1 U1035 ( .A(G125), .B(n1330), .ZN(n1325) );
AND2_X1 U1036 ( .A1(n1061), .A2(G224), .ZN(n1330) );
XNOR2_X1 U1037 ( .A(n1331), .B(n1158), .ZN(n1209) );
XOR2_X1 U1038 ( .A(n1332), .B(n1300), .Z(n1158) );
XNOR2_X1 U1039 ( .A(G116), .B(KEYINPUT60), .ZN(n1300) );
XNOR2_X1 U1040 ( .A(n1333), .B(n1271), .ZN(n1332) );
INV_X1 U1041 ( .A(G113), .ZN(n1271) );
NAND2_X1 U1042 ( .A1(KEYINPUT29), .A2(n1267), .ZN(n1333) );
INV_X1 U1043 ( .A(G119), .ZN(n1267) );
XOR2_X1 U1044 ( .A(n1155), .B(n1159), .Z(n1331) );
XNOR2_X1 U1045 ( .A(G107), .B(n1314), .ZN(n1159) );
XNOR2_X1 U1046 ( .A(n1256), .B(G104), .ZN(n1314) );
INV_X1 U1047 ( .A(G101), .ZN(n1256) );
AND2_X1 U1048 ( .A1(n1334), .A2(n1335), .ZN(n1155) );
NAND2_X1 U1049 ( .A1(G110), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1050 ( .A(n1337), .B(KEYINPUT43), .Z(n1334) );
NAND2_X1 U1051 ( .A1(G122), .A2(n1273), .ZN(n1337) );
NAND2_X1 U1052 ( .A1(G237), .A2(G210), .ZN(n1320) );
NAND2_X1 U1053 ( .A1(n1338), .A2(G237), .ZN(n1095) );
XNOR2_X1 U1054 ( .A(G234), .B(KEYINPUT55), .ZN(n1338) );
NAND2_X1 U1055 ( .A1(n1339), .A2(n1261), .ZN(n1226) );
NAND2_X1 U1056 ( .A1(G952), .A2(n1061), .ZN(n1261) );
NAND3_X1 U1057 ( .A1(G902), .A2(n1160), .A3(G953), .ZN(n1339) );
INV_X1 U1058 ( .A(G898), .ZN(n1160) );
NOR2_X1 U1059 ( .A1(n1266), .A2(n1073), .ZN(n1092) );
XNOR2_X1 U1060 ( .A(n1340), .B(G475), .ZN(n1073) );
OR2_X1 U1061 ( .A1(n1176), .A2(G902), .ZN(n1340) );
XNOR2_X1 U1062 ( .A(n1341), .B(n1342), .ZN(n1176) );
XOR2_X1 U1063 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1064 ( .A(G125), .B(n1345), .ZN(n1344) );
AND3_X1 U1065 ( .A1(G214), .A2(n1061), .A3(n1304), .ZN(n1345) );
INV_X1 U1066 ( .A(G237), .ZN(n1304) );
NAND3_X1 U1067 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1343) );
NAND2_X1 U1068 ( .A1(KEYINPUT0), .A2(G104), .ZN(n1348) );
NAND3_X1 U1069 ( .A1(n1349), .A2(n1350), .A3(n1351), .ZN(n1347) );
INV_X1 U1070 ( .A(KEYINPUT0), .ZN(n1350) );
OR2_X1 U1071 ( .A1(n1351), .A2(n1349), .ZN(n1346) );
NOR2_X1 U1072 ( .A1(n1352), .A2(G104), .ZN(n1349) );
INV_X1 U1073 ( .A(KEYINPUT24), .ZN(n1352) );
XNOR2_X1 U1074 ( .A(G113), .B(n1336), .ZN(n1351) );
XOR2_X1 U1075 ( .A(n1353), .B(n1354), .Z(n1341) );
XNOR2_X1 U1076 ( .A(G146), .B(n1328), .ZN(n1354) );
XNOR2_X1 U1077 ( .A(G131), .B(G140), .ZN(n1353) );
XNOR2_X1 U1078 ( .A(n1355), .B(G478), .ZN(n1266) );
NAND2_X1 U1079 ( .A1(n1168), .A2(n1277), .ZN(n1355) );
INV_X1 U1080 ( .A(G902), .ZN(n1277) );
XNOR2_X1 U1081 ( .A(n1356), .B(n1357), .ZN(n1168) );
NOR2_X1 U1082 ( .A1(KEYINPUT58), .A2(n1358), .ZN(n1357) );
XOR2_X1 U1083 ( .A(n1359), .B(n1360), .Z(n1358) );
XNOR2_X1 U1084 ( .A(n1254), .B(n1361), .ZN(n1360) );
XNOR2_X1 U1085 ( .A(n1328), .B(G134), .ZN(n1361) );
INV_X1 U1086 ( .A(G143), .ZN(n1328) );
INV_X1 U1087 ( .A(G128), .ZN(n1254) );
XNOR2_X1 U1088 ( .A(n1362), .B(n1363), .ZN(n1359) );
INV_X1 U1089 ( .A(G107), .ZN(n1363) );
NAND3_X1 U1090 ( .A1(n1364), .A2(n1365), .A3(n1366), .ZN(n1362) );
NAND2_X1 U1091 ( .A1(KEYINPUT19), .A2(G116), .ZN(n1366) );
NAND3_X1 U1092 ( .A1(n1367), .A2(n1368), .A3(n1336), .ZN(n1365) );
INV_X1 U1093 ( .A(KEYINPUT19), .ZN(n1368) );
OR2_X1 U1094 ( .A1(n1336), .A2(n1367), .ZN(n1364) );
NOR2_X1 U1095 ( .A1(n1369), .A2(G116), .ZN(n1367) );
INV_X1 U1096 ( .A(KEYINPUT53), .ZN(n1369) );
INV_X1 U1097 ( .A(G122), .ZN(n1336) );
NAND3_X1 U1098 ( .A1(G217), .A2(n1061), .A3(G234), .ZN(n1356) );
INV_X1 U1099 ( .A(G953), .ZN(n1061) );
INV_X1 U1100 ( .A(G110), .ZN(n1273) );
endmodule


