//Key = 1001111100110111000111111100110111011010011010110010001001110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;

XOR2_X1 U723 ( .A(n998), .B(n999), .Z(G9) );
NAND4_X1 U724 ( .A1(KEYINPUT15), .A2(n1000), .A3(n1001), .A4(n1002), .ZN(n999) );
NAND4_X1 U725 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(G75) );
NAND3_X1 U726 ( .A1(n1007), .A2(n1008), .A3(G952), .ZN(n1006) );
NAND2_X1 U727 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NAND3_X1 U728 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1010) );
NAND2_X1 U729 ( .A1(n1014), .A2(n1015), .ZN(n1009) );
NAND2_X1 U730 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND3_X1 U731 ( .A1(n1001), .A2(n1018), .A3(n1011), .ZN(n1017) );
NAND2_X1 U732 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND2_X1 U733 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U734 ( .A1(n1012), .A2(n1023), .ZN(n1016) );
NAND2_X1 U735 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND2_X1 U736 ( .A1(n1011), .A2(n1026), .ZN(n1025) );
NAND2_X1 U737 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U738 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND2_X1 U739 ( .A1(n1001), .A2(n1031), .ZN(n1024) );
NAND3_X1 U740 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NAND3_X1 U741 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1033) );
INV_X1 U742 ( .A(KEYINPUT27), .ZN(n1037) );
NAND2_X1 U743 ( .A1(KEYINPUT27), .A2(n1011), .ZN(n1032) );
NOR2_X1 U744 ( .A1(G953), .A2(n1038), .ZN(n1005) );
NOR4_X1 U745 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1038) );
XNOR2_X1 U746 ( .A(n1043), .B(n1044), .ZN(n1042) );
XNOR2_X1 U747 ( .A(KEYINPUT60), .B(n1045), .ZN(n1043) );
NOR2_X1 U748 ( .A1(KEYINPUT1), .A2(n1046), .ZN(n1045) );
AND2_X1 U749 ( .A1(n1047), .A2(n1048), .ZN(n1041) );
NAND3_X1 U750 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1040) );
NAND4_X1 U751 ( .A1(n1052), .A2(n1053), .A3(n1029), .A4(n1054), .ZN(n1039) );
NOR3_X1 U752 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NOR2_X1 U753 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
INV_X1 U754 ( .A(KEYINPUT57), .ZN(n1058) );
NOR2_X1 U755 ( .A1(KEYINPUT57), .A2(G469), .ZN(n1056) );
XOR2_X1 U756 ( .A(KEYINPUT17), .B(n1060), .Z(n1055) );
NOR2_X1 U757 ( .A1(n1048), .A2(n1047), .ZN(n1060) );
XNOR2_X1 U758 ( .A(n1061), .B(KEYINPUT41), .ZN(n1047) );
XOR2_X1 U759 ( .A(n1062), .B(n1063), .Z(n1053) );
NAND2_X1 U760 ( .A1(KEYINPUT44), .A2(n1064), .ZN(n1063) );
XOR2_X1 U761 ( .A(n1065), .B(n1066), .Z(G72) );
NOR2_X1 U762 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U763 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NAND2_X1 U764 ( .A1(n1071), .A2(n1072), .ZN(n1065) );
NAND3_X1 U765 ( .A1(n1073), .A2(n1068), .A3(n1074), .ZN(n1072) );
NAND3_X1 U766 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1071) );
INV_X1 U767 ( .A(n1074), .ZN(n1077) );
NAND2_X1 U768 ( .A1(n1078), .A2(n1079), .ZN(n1074) );
NAND2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U770 ( .A(KEYINPUT42), .B(n1082), .Z(n1078) );
NOR2_X1 U771 ( .A1(n1080), .A2(n1081), .ZN(n1082) );
XOR2_X1 U772 ( .A(n1083), .B(G125), .Z(n1081) );
AND2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1080) );
NAND2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U775 ( .A(KEYINPUT38), .B(n1088), .Z(n1087) );
XOR2_X1 U776 ( .A(n1089), .B(KEYINPUT53), .Z(n1084) );
NAND2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XNOR2_X1 U778 ( .A(n1088), .B(KEYINPUT38), .ZN(n1090) );
NAND2_X1 U779 ( .A1(G953), .A2(n1070), .ZN(n1076) );
XOR2_X1 U780 ( .A(KEYINPUT34), .B(n1003), .Z(n1075) );
XOR2_X1 U781 ( .A(n1092), .B(n1093), .Z(G69) );
NOR2_X1 U782 ( .A1(n1094), .A2(n1068), .ZN(n1093) );
AND2_X1 U783 ( .A1(G224), .A2(G898), .ZN(n1094) );
NAND2_X1 U784 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
NAND3_X1 U785 ( .A1(n1097), .A2(n1068), .A3(n1098), .ZN(n1096) );
XOR2_X1 U786 ( .A(n1099), .B(KEYINPUT26), .Z(n1095) );
OR3_X1 U787 ( .A1(n1098), .A2(n1100), .A3(n1097), .ZN(n1099) );
NOR2_X1 U788 ( .A1(n1101), .A2(n1102), .ZN(G66) );
XOR2_X1 U789 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR2_X1 U790 ( .A1(n1064), .A2(n1105), .ZN(n1103) );
NOR2_X1 U791 ( .A1(n1101), .A2(n1106), .ZN(G63) );
NOR3_X1 U792 ( .A1(n1048), .A2(n1107), .A3(n1108), .ZN(n1106) );
AND3_X1 U793 ( .A1(n1109), .A2(G478), .A3(n1110), .ZN(n1108) );
NOR2_X1 U794 ( .A1(n1111), .A2(n1109), .ZN(n1107) );
NOR2_X1 U795 ( .A1(n1112), .A2(n1061), .ZN(n1111) );
INV_X1 U796 ( .A(G478), .ZN(n1061) );
NOR2_X1 U797 ( .A1(n1097), .A2(n1073), .ZN(n1112) );
NOR2_X1 U798 ( .A1(n1101), .A2(n1113), .ZN(G60) );
XNOR2_X1 U799 ( .A(n1114), .B(n1115), .ZN(n1113) );
NOR2_X1 U800 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NOR2_X1 U801 ( .A1(KEYINPUT37), .A2(n1118), .ZN(n1117) );
INV_X1 U802 ( .A(n1119), .ZN(n1118) );
NOR2_X1 U803 ( .A1(KEYINPUT19), .A2(n1119), .ZN(n1116) );
NAND2_X1 U804 ( .A1(n1110), .A2(G475), .ZN(n1119) );
XOR2_X1 U805 ( .A(n1120), .B(G104), .Z(G6) );
NAND2_X1 U806 ( .A1(KEYINPUT31), .A2(n1121), .ZN(n1120) );
NAND3_X1 U807 ( .A1(n1001), .A2(n1002), .A3(n1122), .ZN(n1121) );
NOR2_X1 U808 ( .A1(n1101), .A2(n1123), .ZN(G57) );
XOR2_X1 U809 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U810 ( .A(G101), .B(n1126), .Z(n1125) );
AND2_X1 U811 ( .A1(G472), .A2(n1110), .ZN(n1126) );
INV_X1 U812 ( .A(n1105), .ZN(n1110) );
NOR2_X1 U813 ( .A1(n1101), .A2(n1127), .ZN(G54) );
XOR2_X1 U814 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U815 ( .A1(n1130), .A2(n1105), .ZN(n1129) );
NAND2_X1 U816 ( .A1(n1131), .A2(n1132), .ZN(n1128) );
NAND4_X1 U817 ( .A1(n1133), .A2(KEYINPUT54), .A3(n1134), .A4(n1135), .ZN(n1132) );
NAND2_X1 U818 ( .A1(n1136), .A2(n1137), .ZN(n1131) );
NAND2_X1 U819 ( .A1(n1134), .A2(n1138), .ZN(n1137) );
OR2_X1 U820 ( .A1(n1133), .A2(KEYINPUT54), .ZN(n1138) );
XOR2_X1 U821 ( .A(n1139), .B(n1140), .Z(n1134) );
NAND2_X1 U822 ( .A1(KEYINPUT47), .A2(n1141), .ZN(n1139) );
NAND2_X1 U823 ( .A1(n1133), .A2(n1135), .ZN(n1136) );
INV_X1 U824 ( .A(KEYINPUT9), .ZN(n1135) );
XOR2_X1 U825 ( .A(n1142), .B(n1143), .Z(n1133) );
NOR2_X1 U826 ( .A1(n1101), .A2(n1144), .ZN(G51) );
XOR2_X1 U827 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U828 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U829 ( .A(G125), .B(n1149), .Z(n1148) );
NOR2_X1 U830 ( .A1(KEYINPUT39), .A2(n1150), .ZN(n1147) );
XOR2_X1 U831 ( .A(n1086), .B(n1151), .Z(n1145) );
NOR2_X1 U832 ( .A1(n1044), .A2(n1105), .ZN(n1151) );
NAND2_X1 U833 ( .A1(G902), .A2(n1152), .ZN(n1105) );
NAND2_X1 U834 ( .A1(n1003), .A2(n1004), .ZN(n1152) );
INV_X1 U835 ( .A(n1097), .ZN(n1004) );
NAND4_X1 U836 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1097) );
NOR3_X1 U837 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1156) );
NOR2_X1 U838 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U839 ( .A(KEYINPUT11), .B(n1162), .Z(n1161) );
INV_X1 U840 ( .A(n1163), .ZN(n1158) );
NOR2_X1 U841 ( .A1(n1164), .A2(n1165), .ZN(n1157) );
NOR2_X1 U842 ( .A1(n1166), .A2(n1013), .ZN(n1164) );
AND2_X1 U843 ( .A1(n1001), .A2(n1167), .ZN(n1013) );
NAND2_X1 U844 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U845 ( .A1(n1170), .A2(n1027), .ZN(n1166) );
XOR2_X1 U846 ( .A(n1171), .B(KEYINPUT52), .Z(n1170) );
INV_X1 U847 ( .A(n1073), .ZN(n1003) );
NAND4_X1 U848 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1073) );
NOR4_X1 U849 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1175) );
INV_X1 U850 ( .A(n1180), .ZN(n1178) );
NOR3_X1 U851 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1174) );
NOR2_X1 U852 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
AND4_X1 U853 ( .A1(n1184), .A2(n1186), .A3(n1019), .A4(n1187), .ZN(n1182) );
INV_X1 U854 ( .A(n1188), .ZN(n1019) );
INV_X1 U855 ( .A(KEYINPUT29), .ZN(n1184) );
NOR3_X1 U856 ( .A1(n1189), .A2(n1190), .A3(n1171), .ZN(n1181) );
XOR2_X1 U857 ( .A(KEYINPUT59), .B(n1011), .Z(n1189) );
NOR2_X1 U858 ( .A1(n1068), .A2(G952), .ZN(n1101) );
XNOR2_X1 U859 ( .A(n1177), .B(n1191), .ZN(G48) );
NAND2_X1 U860 ( .A1(KEYINPUT7), .A2(G146), .ZN(n1191) );
NOR3_X1 U861 ( .A1(n1190), .A2(n1034), .A3(n1168), .ZN(n1177) );
XNOR2_X1 U862 ( .A(G143), .B(n1185), .ZN(G45) );
NAND3_X1 U863 ( .A1(n1188), .A2(n1187), .A3(n1186), .ZN(n1185) );
NOR4_X1 U864 ( .A1(n1027), .A2(n1034), .A3(n1192), .A4(n1052), .ZN(n1186) );
XOR2_X1 U865 ( .A(n1172), .B(n1193), .Z(G42) );
XOR2_X1 U866 ( .A(n1083), .B(KEYINPUT43), .Z(n1193) );
NAND2_X1 U867 ( .A1(n1194), .A2(n1195), .ZN(n1172) );
XOR2_X1 U868 ( .A(G137), .B(n1196), .Z(G39) );
NOR3_X1 U869 ( .A1(n1171), .A2(n1190), .A3(n1197), .ZN(n1196) );
XOR2_X1 U870 ( .A(n1198), .B(n1173), .Z(G36) );
NAND3_X1 U871 ( .A1(n1194), .A2(n1000), .A3(n1199), .ZN(n1173) );
XOR2_X1 U872 ( .A(G131), .B(n1179), .Z(G33) );
AND3_X1 U873 ( .A1(n1194), .A2(n1122), .A3(n1199), .ZN(n1179) );
AND3_X1 U874 ( .A1(n1188), .A2(n1187), .A3(n1011), .ZN(n1194) );
INV_X1 U875 ( .A(n1197), .ZN(n1011) );
NAND2_X1 U876 ( .A1(n1036), .A2(n1051), .ZN(n1197) );
XOR2_X1 U877 ( .A(G128), .B(n1176), .Z(G30) );
NOR3_X1 U878 ( .A1(n1169), .A2(n1034), .A3(n1190), .ZN(n1176) );
NAND4_X1 U879 ( .A1(n1188), .A2(n1030), .A3(n1200), .A4(n1187), .ZN(n1190) );
INV_X1 U880 ( .A(n1000), .ZN(n1169) );
XOR2_X1 U881 ( .A(n1201), .B(n1202), .Z(G3) );
NOR3_X1 U882 ( .A1(n1171), .A2(n1165), .A3(n1027), .ZN(n1202) );
NOR2_X1 U883 ( .A1(KEYINPUT12), .A2(n1203), .ZN(n1201) );
INV_X1 U884 ( .A(G101), .ZN(n1203) );
XOR2_X1 U885 ( .A(n1204), .B(n1180), .Z(G27) );
NAND4_X1 U886 ( .A1(n1012), .A2(n1195), .A3(n1162), .A4(n1187), .ZN(n1180) );
NAND2_X1 U887 ( .A1(n1205), .A2(n1206), .ZN(n1187) );
NAND4_X1 U888 ( .A1(G902), .A2(G953), .A3(n1008), .A4(n1070), .ZN(n1206) );
INV_X1 U889 ( .A(G900), .ZN(n1070) );
NOR3_X1 U890 ( .A1(n1200), .A2(n1207), .A3(n1168), .ZN(n1195) );
XOR2_X1 U891 ( .A(n1208), .B(n1163), .Z(G24) );
NAND3_X1 U892 ( .A1(n1209), .A2(n1001), .A3(n1210), .ZN(n1163) );
NOR3_X1 U893 ( .A1(n1034), .A2(n1052), .A3(n1192), .ZN(n1210) );
NOR2_X1 U894 ( .A1(n1200), .A2(n1030), .ZN(n1001) );
XOR2_X1 U895 ( .A(n1211), .B(n1212), .Z(G21) );
NAND2_X1 U896 ( .A1(KEYINPUT10), .A2(n1213), .ZN(n1212) );
INV_X1 U897 ( .A(n1155), .ZN(n1213) );
NAND3_X1 U898 ( .A1(n1209), .A2(n1014), .A3(n1214), .ZN(n1155) );
NOR3_X1 U899 ( .A1(n1034), .A2(n1029), .A3(n1207), .ZN(n1214) );
INV_X1 U900 ( .A(n1162), .ZN(n1034) );
XOR2_X1 U901 ( .A(n1153), .B(n1215), .Z(G18) );
NAND2_X1 U902 ( .A1(KEYINPUT24), .A2(G116), .ZN(n1215) );
NAND4_X1 U903 ( .A1(n1209), .A2(n1199), .A3(n1000), .A4(n1162), .ZN(n1153) );
NOR2_X1 U904 ( .A1(n1216), .A2(n1192), .ZN(n1000) );
XNOR2_X1 U905 ( .A(G113), .B(n1217), .ZN(G15) );
NAND2_X1 U906 ( .A1(n1218), .A2(n1162), .ZN(n1217) );
XOR2_X1 U907 ( .A(n1160), .B(KEYINPUT23), .Z(n1218) );
NAND3_X1 U908 ( .A1(n1199), .A2(n1122), .A3(n1209), .ZN(n1160) );
AND2_X1 U909 ( .A1(n1012), .A2(n1219), .ZN(n1209) );
AND2_X1 U910 ( .A1(n1021), .A2(n1220), .ZN(n1012) );
XOR2_X1 U911 ( .A(KEYINPUT14), .B(n1022), .Z(n1220) );
INV_X1 U912 ( .A(n1168), .ZN(n1122) );
NAND2_X1 U913 ( .A1(n1192), .A2(n1221), .ZN(n1168) );
XOR2_X1 U914 ( .A(KEYINPUT49), .B(n1216), .Z(n1221) );
INV_X1 U915 ( .A(n1027), .ZN(n1199) );
NAND2_X1 U916 ( .A1(n1207), .A2(n1200), .ZN(n1027) );
INV_X1 U917 ( .A(n1029), .ZN(n1200) );
XNOR2_X1 U918 ( .A(G110), .B(n1154), .ZN(G12) );
NAND4_X1 U919 ( .A1(n1014), .A2(n1002), .A3(n1029), .A4(n1030), .ZN(n1154) );
INV_X1 U920 ( .A(n1207), .ZN(n1030) );
XNOR2_X1 U921 ( .A(n1062), .B(n1064), .ZN(n1207) );
NAND2_X1 U922 ( .A1(G217), .A2(n1222), .ZN(n1064) );
NAND2_X1 U923 ( .A1(n1223), .A2(n1224), .ZN(n1062) );
XOR2_X1 U924 ( .A(KEYINPUT5), .B(n1104), .Z(n1223) );
XNOR2_X1 U925 ( .A(n1225), .B(n1226), .ZN(n1104) );
XOR2_X1 U926 ( .A(n1227), .B(n1228), .Z(n1226) );
XNOR2_X1 U927 ( .A(G146), .B(KEYINPUT3), .ZN(n1228) );
NAND2_X1 U928 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
NAND2_X1 U929 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND3_X1 U930 ( .A1(G234), .A2(n1068), .A3(G221), .ZN(n1232) );
XOR2_X1 U931 ( .A(n1233), .B(KEYINPUT63), .Z(n1229) );
NAND4_X1 U932 ( .A1(n1234), .A2(G221), .A3(G234), .A4(n1068), .ZN(n1233) );
XOR2_X1 U933 ( .A(n1231), .B(KEYINPUT32), .Z(n1234) );
INV_X1 U934 ( .A(G137), .ZN(n1231) );
XNOR2_X1 U935 ( .A(n1140), .B(n1235), .ZN(n1225) );
XNOR2_X1 U936 ( .A(n1236), .B(n1237), .ZN(n1235) );
NOR2_X1 U937 ( .A1(KEYINPUT48), .A2(n1238), .ZN(n1237) );
XOR2_X1 U938 ( .A(n1211), .B(n1239), .Z(n1238) );
NAND2_X1 U939 ( .A1(KEYINPUT33), .A2(n1240), .ZN(n1239) );
INV_X1 U940 ( .A(G128), .ZN(n1240) );
NAND2_X1 U941 ( .A1(KEYINPUT13), .A2(G125), .ZN(n1236) );
XOR2_X1 U942 ( .A(n1241), .B(G472), .Z(n1029) );
NAND2_X1 U943 ( .A1(n1242), .A2(n1224), .ZN(n1241) );
XOR2_X1 U944 ( .A(n1124), .B(n1243), .Z(n1242) );
XOR2_X1 U945 ( .A(KEYINPUT55), .B(n1244), .Z(n1243) );
NOR2_X1 U946 ( .A1(G101), .A2(KEYINPUT40), .ZN(n1244) );
XOR2_X1 U947 ( .A(n1245), .B(n1246), .Z(n1124) );
XOR2_X1 U948 ( .A(n1247), .B(n1248), .Z(n1246) );
NAND2_X1 U949 ( .A1(G210), .A2(n1249), .ZN(n1247) );
XOR2_X1 U950 ( .A(n1142), .B(n1250), .Z(n1245) );
NOR2_X1 U951 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NOR2_X1 U952 ( .A1(n1211), .A2(n1253), .ZN(n1252) );
XNOR2_X1 U953 ( .A(G116), .B(KEYINPUT50), .ZN(n1253) );
INV_X1 U954 ( .A(G119), .ZN(n1211) );
NOR2_X1 U955 ( .A1(G119), .A2(n1254), .ZN(n1251) );
XNOR2_X1 U956 ( .A(G116), .B(KEYINPUT30), .ZN(n1254) );
XOR2_X1 U957 ( .A(n1255), .B(n1091), .Z(n1142) );
INV_X1 U958 ( .A(n1165), .ZN(n1002) );
NAND3_X1 U959 ( .A1(n1162), .A2(n1219), .A3(n1188), .ZN(n1165) );
NOR2_X1 U960 ( .A1(n1022), .A2(n1021), .ZN(n1188) );
AND2_X1 U961 ( .A1(n1256), .A2(n1049), .ZN(n1021) );
NAND3_X1 U962 ( .A1(n1130), .A2(n1224), .A3(n1257), .ZN(n1049) );
INV_X1 U963 ( .A(G469), .ZN(n1130) );
XNOR2_X1 U964 ( .A(KEYINPUT21), .B(n1059), .ZN(n1256) );
NAND2_X1 U965 ( .A1(G469), .A2(n1258), .ZN(n1059) );
NAND2_X1 U966 ( .A1(n1257), .A2(n1224), .ZN(n1258) );
XNOR2_X1 U967 ( .A(n1259), .B(n1260), .ZN(n1257) );
XNOR2_X1 U968 ( .A(n1255), .B(n1140), .ZN(n1260) );
XOR2_X1 U969 ( .A(G110), .B(G140), .Z(n1140) );
XNOR2_X1 U970 ( .A(n1088), .B(KEYINPUT2), .ZN(n1255) );
XOR2_X1 U971 ( .A(G131), .B(n1261), .Z(n1088) );
XOR2_X1 U972 ( .A(G137), .B(G134), .Z(n1261) );
XOR2_X1 U973 ( .A(n1262), .B(n1141), .Z(n1259) );
NOR2_X1 U974 ( .A1(n1069), .A2(G953), .ZN(n1141) );
INV_X1 U975 ( .A(G227), .ZN(n1069) );
NAND2_X1 U976 ( .A1(KEYINPUT61), .A2(n1263), .ZN(n1262) );
XOR2_X1 U977 ( .A(n1091), .B(n1143), .Z(n1263) );
INV_X1 U978 ( .A(n1050), .ZN(n1022) );
NAND2_X1 U979 ( .A1(G221), .A2(n1222), .ZN(n1050) );
NAND2_X1 U980 ( .A1(G234), .A2(n1224), .ZN(n1222) );
NAND2_X1 U981 ( .A1(n1205), .A2(n1264), .ZN(n1219) );
NAND3_X1 U982 ( .A1(n1100), .A2(n1008), .A3(G902), .ZN(n1264) );
NOR2_X1 U983 ( .A1(n1068), .A2(G898), .ZN(n1100) );
NAND3_X1 U984 ( .A1(n1008), .A2(n1068), .A3(G952), .ZN(n1205) );
NAND2_X1 U985 ( .A1(n1265), .A2(G237), .ZN(n1008) );
XNOR2_X1 U986 ( .A(G234), .B(KEYINPUT28), .ZN(n1265) );
NOR2_X1 U987 ( .A1(n1036), .A2(n1035), .ZN(n1162) );
INV_X1 U988 ( .A(n1051), .ZN(n1035) );
NAND2_X1 U989 ( .A1(G214), .A2(n1266), .ZN(n1051) );
XOR2_X1 U990 ( .A(n1267), .B(n1044), .Z(n1036) );
NAND2_X1 U991 ( .A1(G210), .A2(n1266), .ZN(n1044) );
NAND2_X1 U992 ( .A1(n1268), .A2(n1224), .ZN(n1266) );
INV_X1 U993 ( .A(G237), .ZN(n1268) );
XNOR2_X1 U994 ( .A(n1046), .B(KEYINPUT58), .ZN(n1267) );
AND2_X1 U995 ( .A1(n1269), .A2(n1224), .ZN(n1046) );
XOR2_X1 U996 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U997 ( .A(n1272), .B(n1149), .Z(n1271) );
AND2_X1 U998 ( .A1(G224), .A2(n1068), .ZN(n1149) );
NAND2_X1 U999 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
OR2_X1 U1000 ( .A1(n1275), .A2(n1091), .ZN(n1274) );
XOR2_X1 U1001 ( .A(n1276), .B(KEYINPUT16), .Z(n1273) );
NAND2_X1 U1002 ( .A1(n1275), .A2(n1091), .ZN(n1276) );
INV_X1 U1003 ( .A(n1086), .ZN(n1091) );
XNOR2_X1 U1004 ( .A(G146), .B(n1277), .ZN(n1086) );
XNOR2_X1 U1005 ( .A(n1204), .B(KEYINPUT36), .ZN(n1275) );
NAND2_X1 U1006 ( .A1(KEYINPUT46), .A2(n1150), .ZN(n1270) );
INV_X1 U1007 ( .A(n1098), .ZN(n1150) );
XOR2_X1 U1008 ( .A(n1278), .B(n1279), .Z(n1098) );
XOR2_X1 U1009 ( .A(n1143), .B(n1280), .Z(n1279) );
XNOR2_X1 U1010 ( .A(n1281), .B(n1282), .ZN(n1280) );
NOR2_X1 U1011 ( .A1(KEYINPUT56), .A2(n1283), .ZN(n1282) );
INV_X1 U1012 ( .A(n1248), .ZN(n1283) );
NAND2_X1 U1013 ( .A1(KEYINPUT25), .A2(n1208), .ZN(n1281) );
XOR2_X1 U1014 ( .A(G101), .B(n1284), .Z(n1143) );
XOR2_X1 U1015 ( .A(G107), .B(G104), .Z(n1284) );
XNOR2_X1 U1016 ( .A(G110), .B(n1285), .ZN(n1278) );
XOR2_X1 U1017 ( .A(G119), .B(G116), .Z(n1285) );
INV_X1 U1018 ( .A(n1171), .ZN(n1014) );
NAND2_X1 U1019 ( .A1(n1192), .A2(n1052), .ZN(n1171) );
INV_X1 U1020 ( .A(n1216), .ZN(n1052) );
XNOR2_X1 U1021 ( .A(n1286), .B(G475), .ZN(n1216) );
NAND2_X1 U1022 ( .A1(n1224), .A2(n1114), .ZN(n1286) );
NAND2_X1 U1023 ( .A1(n1287), .A2(n1288), .ZN(n1114) );
NAND2_X1 U1024 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XOR2_X1 U1025 ( .A(KEYINPUT6), .B(n1291), .Z(n1287) );
NOR2_X1 U1026 ( .A1(n1289), .A2(n1290), .ZN(n1291) );
XNOR2_X1 U1027 ( .A(n1292), .B(n1293), .ZN(n1290) );
NOR2_X1 U1028 ( .A1(KEYINPUT18), .A2(n1248), .ZN(n1293) );
XNOR2_X1 U1029 ( .A(G113), .B(KEYINPUT22), .ZN(n1248) );
XOR2_X1 U1030 ( .A(G104), .B(n1208), .Z(n1292) );
INV_X1 U1031 ( .A(G122), .ZN(n1208) );
XOR2_X1 U1032 ( .A(n1294), .B(n1295), .Z(n1289) );
XOR2_X1 U1033 ( .A(n1296), .B(n1297), .Z(n1295) );
XNOR2_X1 U1034 ( .A(G131), .B(G146), .ZN(n1297) );
NAND3_X1 U1035 ( .A1(n1298), .A2(n1299), .A3(KEYINPUT4), .ZN(n1296) );
NAND2_X1 U1036 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
INV_X1 U1037 ( .A(KEYINPUT51), .ZN(n1301) );
XOR2_X1 U1038 ( .A(G140), .B(n1302), .Z(n1300) );
AND2_X1 U1039 ( .A1(n1204), .A2(KEYINPUT0), .ZN(n1302) );
NAND3_X1 U1040 ( .A1(n1303), .A2(n1204), .A3(KEYINPUT51), .ZN(n1298) );
INV_X1 U1041 ( .A(G125), .ZN(n1204) );
XOR2_X1 U1042 ( .A(KEYINPUT0), .B(n1083), .Z(n1303) );
INV_X1 U1043 ( .A(G140), .ZN(n1083) );
XOR2_X1 U1044 ( .A(n1304), .B(n1305), .Z(n1294) );
NOR2_X1 U1045 ( .A1(G143), .A2(KEYINPUT62), .ZN(n1305) );
NAND2_X1 U1046 ( .A1(G214), .A2(n1249), .ZN(n1304) );
NOR2_X1 U1047 ( .A1(G953), .A2(G237), .ZN(n1249) );
INV_X1 U1048 ( .A(G902), .ZN(n1224) );
XNOR2_X1 U1049 ( .A(n1048), .B(G478), .ZN(n1192) );
NOR2_X1 U1050 ( .A1(n1109), .A2(G902), .ZN(n1048) );
XOR2_X1 U1051 ( .A(n1306), .B(n1307), .Z(n1109) );
NOR4_X1 U1052 ( .A1(n1308), .A2(n1309), .A3(KEYINPUT8), .A4(n1310), .ZN(n1307) );
NOR2_X1 U1053 ( .A1(KEYINPUT35), .A2(n1311), .ZN(n1310) );
NOR2_X1 U1054 ( .A1(n1312), .A2(n1313), .ZN(n1309) );
AND2_X1 U1055 ( .A1(n1314), .A2(n1311), .ZN(n1312) );
AND4_X1 U1056 ( .A1(n1313), .A2(KEYINPUT35), .A3(n1314), .A4(n1311), .ZN(n1308) );
XNOR2_X1 U1057 ( .A(n1315), .B(n1277), .ZN(n1311) );
XOR2_X1 U1058 ( .A(G128), .B(G143), .Z(n1277) );
NAND2_X1 U1059 ( .A1(KEYINPUT20), .A2(n1198), .ZN(n1315) );
INV_X1 U1060 ( .A(G134), .ZN(n1198) );
INV_X1 U1061 ( .A(KEYINPUT45), .ZN(n1314) );
XOR2_X1 U1062 ( .A(n998), .B(n1316), .Z(n1313) );
XOR2_X1 U1063 ( .A(G122), .B(G116), .Z(n1316) );
INV_X1 U1064 ( .A(G107), .ZN(n998) );
NAND3_X1 U1065 ( .A1(G217), .A2(n1068), .A3(G234), .ZN(n1306) );
INV_X1 U1066 ( .A(G953), .ZN(n1068) );
endmodule


