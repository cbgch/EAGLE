//Key = 1001110001101000101101010010110110010100100010001100001001100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424;

XNOR2_X1 U773 ( .A(n1075), .B(n1076), .ZN(G9) );
NOR2_X1 U774 ( .A1(n1077), .A2(n1078), .ZN(G75) );
NOR4_X1 U775 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1082), .ZN(n1078) );
NAND2_X1 U776 ( .A1(n1083), .A2(n1084), .ZN(n1080) );
NOR3_X1 U777 ( .A1(n1085), .A2(KEYINPUT1), .A3(n1086), .ZN(n1079) );
NOR2_X1 U778 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR3_X1 U779 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
NOR3_X1 U780 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1090) );
NOR2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR3_X1 U782 ( .A1(n1097), .A2(n1098), .A3(n1095), .ZN(n1087) );
NOR3_X1 U783 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
NOR3_X1 U784 ( .A1(n1102), .A2(n1103), .A3(n1089), .ZN(n1101) );
NOR2_X1 U785 ( .A1(n1104), .A2(n1091), .ZN(n1099) );
NOR2_X1 U786 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
AND2_X1 U787 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
NOR3_X1 U788 ( .A1(n1109), .A2(G953), .A3(G952), .ZN(n1077) );
INV_X1 U789 ( .A(n1083), .ZN(n1109) );
NAND4_X1 U790 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1083) );
NOR4_X1 U791 ( .A1(n1091), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1113) );
XNOR2_X1 U792 ( .A(G475), .B(n1117), .ZN(n1116) );
XOR2_X1 U793 ( .A(KEYINPUT22), .B(n1118), .Z(n1115) );
NOR3_X1 U794 ( .A1(n1119), .A2(n1120), .A3(n1108), .ZN(n1112) );
NOR2_X1 U795 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
XOR2_X1 U796 ( .A(KEYINPUT48), .B(G472), .Z(n1122) );
INV_X1 U797 ( .A(n1123), .ZN(n1121) );
NAND2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1111) );
XNOR2_X1 U799 ( .A(KEYINPUT38), .B(n1126), .ZN(n1110) );
XOR2_X1 U800 ( .A(n1127), .B(n1128), .Z(G72) );
XOR2_X1 U801 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U802 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U803 ( .A1(G900), .A2(G227), .ZN(n1132) );
NAND2_X1 U804 ( .A1(n1133), .A2(n1134), .ZN(n1129) );
NAND2_X1 U805 ( .A1(G953), .A2(n1135), .ZN(n1134) );
XOR2_X1 U806 ( .A(n1136), .B(n1137), .Z(n1133) );
XNOR2_X1 U807 ( .A(n1138), .B(G140), .ZN(n1137) );
XOR2_X1 U808 ( .A(n1139), .B(n1140), .Z(n1136) );
NAND2_X1 U809 ( .A1(KEYINPUT32), .A2(n1141), .ZN(n1139) );
NAND2_X1 U810 ( .A1(KEYINPUT16), .A2(n1142), .ZN(n1127) );
NAND2_X1 U811 ( .A1(n1082), .A2(n1084), .ZN(n1142) );
XOR2_X1 U812 ( .A(n1143), .B(n1144), .Z(G69) );
NOR2_X1 U813 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
INV_X1 U814 ( .A(n1131), .ZN(n1146) );
XOR2_X1 U815 ( .A(G953), .B(KEYINPUT55), .Z(n1131) );
AND2_X1 U816 ( .A1(G224), .A2(G898), .ZN(n1145) );
NAND2_X1 U817 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
NAND2_X1 U818 ( .A1(n1149), .A2(n1084), .ZN(n1148) );
XOR2_X1 U819 ( .A(n1081), .B(n1150), .Z(n1149) );
NAND3_X1 U820 ( .A1(n1151), .A2(n1150), .A3(G953), .ZN(n1147) );
XNOR2_X1 U821 ( .A(n1152), .B(n1153), .ZN(n1150) );
XOR2_X1 U822 ( .A(KEYINPUT35), .B(n1154), .Z(n1153) );
XNOR2_X1 U823 ( .A(KEYINPUT34), .B(n1155), .ZN(n1151) );
NOR2_X1 U824 ( .A1(n1156), .A2(n1157), .ZN(G66) );
XOR2_X1 U825 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U826 ( .A(n1160), .B(KEYINPUT4), .Z(n1158) );
NAND2_X1 U827 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U828 ( .A1(n1156), .A2(n1163), .ZN(G63) );
XOR2_X1 U829 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U830 ( .A1(n1161), .A2(G478), .ZN(n1164) );
NOR2_X1 U831 ( .A1(n1156), .A2(n1166), .ZN(G60) );
XOR2_X1 U832 ( .A(n1167), .B(n1168), .Z(n1166) );
NAND2_X1 U833 ( .A1(n1161), .A2(G475), .ZN(n1167) );
XNOR2_X1 U834 ( .A(G104), .B(n1169), .ZN(G6) );
NAND3_X1 U835 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1169) );
XNOR2_X1 U836 ( .A(n1173), .B(KEYINPUT61), .ZN(n1172) );
NOR2_X1 U837 ( .A1(n1156), .A2(n1174), .ZN(G57) );
XOR2_X1 U838 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U839 ( .A(n1177), .B(n1178), .Z(n1176) );
XNOR2_X1 U840 ( .A(G101), .B(KEYINPUT30), .ZN(n1178) );
XOR2_X1 U841 ( .A(n1179), .B(n1180), .Z(n1175) );
XOR2_X1 U842 ( .A(n1181), .B(n1182), .Z(n1179) );
NAND2_X1 U843 ( .A1(n1161), .A2(G472), .ZN(n1181) );
NOR2_X1 U844 ( .A1(n1156), .A2(n1183), .ZN(G54) );
XOR2_X1 U845 ( .A(n1184), .B(n1185), .Z(n1183) );
XOR2_X1 U846 ( .A(n1186), .B(n1187), .Z(n1184) );
NOR2_X1 U847 ( .A1(KEYINPUT24), .A2(n1188), .ZN(n1187) );
NAND3_X1 U848 ( .A1(G469), .A2(n1189), .A3(n1190), .ZN(n1186) );
XNOR2_X1 U849 ( .A(KEYINPUT3), .B(G902), .ZN(n1190) );
XOR2_X1 U850 ( .A(KEYINPUT9), .B(n1191), .Z(n1189) );
NOR2_X1 U851 ( .A1(n1156), .A2(n1192), .ZN(G51) );
XOR2_X1 U852 ( .A(n1193), .B(n1194), .Z(n1192) );
XNOR2_X1 U853 ( .A(n1195), .B(n1196), .ZN(n1194) );
NAND2_X1 U854 ( .A1(n1197), .A2(n1198), .ZN(n1195) );
INV_X1 U855 ( .A(n1199), .ZN(n1197) );
XOR2_X1 U856 ( .A(n1200), .B(KEYINPUT41), .Z(n1193) );
NAND3_X1 U857 ( .A1(G210), .A2(n1201), .A3(n1161), .ZN(n1200) );
NOR2_X1 U858 ( .A1(n1202), .A2(n1191), .ZN(n1161) );
NOR2_X1 U859 ( .A1(n1082), .A2(n1203), .ZN(n1191) );
XOR2_X1 U860 ( .A(KEYINPUT43), .B(n1081), .Z(n1203) );
NAND4_X1 U861 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1081) );
NOR3_X1 U862 ( .A1(n1208), .A2(n1209), .A3(n1076), .ZN(n1207) );
NOR3_X1 U863 ( .A1(n1096), .A2(n1095), .A3(n1210), .ZN(n1076) );
INV_X1 U864 ( .A(n1211), .ZN(n1208) );
NAND2_X1 U865 ( .A1(n1170), .A2(n1212), .ZN(n1206) );
NAND3_X1 U866 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1212) );
INV_X1 U867 ( .A(n1092), .ZN(n1215) );
NAND2_X1 U868 ( .A1(n1216), .A2(n1217), .ZN(n1092) );
NAND2_X1 U869 ( .A1(n1173), .A2(n1171), .ZN(n1217) );
NAND2_X1 U870 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
NAND3_X1 U871 ( .A1(n1220), .A2(n1097), .A3(n1221), .ZN(n1214) );
INV_X1 U872 ( .A(KEYINPUT44), .ZN(n1221) );
NAND2_X1 U873 ( .A1(KEYINPUT44), .A2(n1093), .ZN(n1213) );
NAND3_X1 U874 ( .A1(n1222), .A2(n1223), .A3(KEYINPUT33), .ZN(n1205) );
NAND3_X1 U875 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1223) );
INV_X1 U876 ( .A(n1089), .ZN(n1224) );
NAND2_X1 U877 ( .A1(n1227), .A2(n1228), .ZN(n1204) );
NAND2_X1 U878 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NAND2_X1 U879 ( .A1(n1226), .A2(n1231), .ZN(n1230) );
INV_X1 U880 ( .A(KEYINPUT33), .ZN(n1231) );
NAND4_X1 U881 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1082) );
NOR4_X1 U882 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235) );
NOR3_X1 U883 ( .A1(n1240), .A2(n1241), .A3(n1096), .ZN(n1239) );
NOR3_X1 U884 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1234) );
NOR2_X1 U885 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND4_X1 U886 ( .A1(n1100), .A2(n1173), .A3(n1247), .A4(n1248), .ZN(n1246) );
INV_X1 U887 ( .A(KEYINPUT36), .ZN(n1245) );
NOR2_X1 U888 ( .A1(KEYINPUT36), .A2(n1249), .ZN(n1243) );
NOR2_X1 U889 ( .A1(KEYINPUT50), .A2(n1250), .ZN(n1242) );
NAND2_X1 U890 ( .A1(n1251), .A2(n1252), .ZN(n1233) );
XOR2_X1 U891 ( .A(KEYINPUT59), .B(n1106), .Z(n1252) );
INV_X1 U892 ( .A(n1253), .ZN(n1251) );
NAND2_X1 U893 ( .A1(n1254), .A2(n1255), .ZN(n1232) );
NAND2_X1 U894 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND4_X1 U895 ( .A1(KEYINPUT50), .A2(n1258), .A3(n1259), .A4(n1106), .ZN(n1257) );
XOR2_X1 U896 ( .A(n1260), .B(KEYINPUT11), .Z(n1256) );
XNOR2_X1 U897 ( .A(KEYINPUT3), .B(n1261), .ZN(n1202) );
NOR2_X1 U898 ( .A1(n1084), .A2(G952), .ZN(n1156) );
XOR2_X1 U899 ( .A(G146), .B(n1262), .Z(G48) );
NOR2_X1 U900 ( .A1(KEYINPUT46), .A2(n1263), .ZN(n1262) );
INV_X1 U901 ( .A(n1238), .ZN(n1263) );
NOR3_X1 U902 ( .A1(n1240), .A2(n1241), .A3(n1264), .ZN(n1238) );
XNOR2_X1 U903 ( .A(n1265), .B(n1266), .ZN(G45) );
NOR2_X1 U904 ( .A1(n1267), .A2(n1253), .ZN(n1266) );
NAND3_X1 U905 ( .A1(n1126), .A2(n1220), .A3(n1268), .ZN(n1253) );
NOR3_X1 U906 ( .A1(n1269), .A2(n1259), .A3(n1241), .ZN(n1268) );
XNOR2_X1 U907 ( .A(n1106), .B(KEYINPUT13), .ZN(n1267) );
XOR2_X1 U908 ( .A(n1237), .B(n1270), .Z(G42) );
XNOR2_X1 U909 ( .A(KEYINPUT7), .B(n1271), .ZN(n1270) );
AND3_X1 U910 ( .A1(n1254), .A2(n1106), .A3(n1272), .ZN(n1237) );
XOR2_X1 U911 ( .A(G137), .B(n1236), .Z(G39) );
NOR3_X1 U912 ( .A1(n1097), .A2(n1091), .A3(n1240), .ZN(n1236) );
INV_X1 U913 ( .A(n1219), .ZN(n1097) );
XOR2_X1 U914 ( .A(n1273), .B(n1274), .Z(G36) );
NOR2_X1 U915 ( .A1(KEYINPUT2), .A2(n1275), .ZN(n1274) );
NOR2_X1 U916 ( .A1(n1091), .A2(n1260), .ZN(n1273) );
NAND2_X1 U917 ( .A1(n1276), .A2(n1277), .ZN(n1260) );
INV_X1 U918 ( .A(n1254), .ZN(n1091) );
XNOR2_X1 U919 ( .A(G131), .B(n1250), .ZN(G33) );
NAND3_X1 U920 ( .A1(n1173), .A2(n1254), .A3(n1276), .ZN(n1250) );
AND3_X1 U921 ( .A1(n1106), .A2(n1247), .A3(n1220), .ZN(n1276) );
NOR2_X1 U922 ( .A1(n1103), .A2(n1278), .ZN(n1254) );
INV_X1 U923 ( .A(n1102), .ZN(n1278) );
XNOR2_X1 U924 ( .A(G128), .B(n1279), .ZN(G30) );
NAND2_X1 U925 ( .A1(n1222), .A2(n1280), .ZN(n1279) );
XOR2_X1 U926 ( .A(KEYINPUT17), .B(n1281), .Z(n1280) );
NOR2_X1 U927 ( .A1(n1096), .A2(n1240), .ZN(n1281) );
NAND4_X1 U928 ( .A1(n1106), .A2(n1114), .A3(n1247), .A4(n1282), .ZN(n1240) );
NAND2_X1 U929 ( .A1(n1283), .A2(n1284), .ZN(G3) );
NAND3_X1 U930 ( .A1(n1285), .A2(n1286), .A3(KEYINPUT40), .ZN(n1284) );
NAND2_X1 U931 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
NAND2_X1 U932 ( .A1(KEYINPUT0), .A2(n1289), .ZN(n1285) );
NAND3_X1 U933 ( .A1(n1170), .A2(n1287), .A3(n1093), .ZN(n1289) );
NAND2_X1 U934 ( .A1(n1290), .A2(n1291), .ZN(n1283) );
NAND2_X1 U935 ( .A1(n1292), .A2(n1287), .ZN(n1291) );
OR2_X1 U936 ( .A1(n1288), .A2(KEYINPUT40), .ZN(n1292) );
INV_X1 U937 ( .A(KEYINPUT0), .ZN(n1288) );
NAND2_X1 U938 ( .A1(n1093), .A2(n1170), .ZN(n1290) );
AND2_X1 U939 ( .A1(n1220), .A2(n1219), .ZN(n1093) );
NAND2_X1 U940 ( .A1(n1293), .A2(n1294), .ZN(G27) );
NAND2_X1 U941 ( .A1(n1295), .A2(n1141), .ZN(n1294) );
XOR2_X1 U942 ( .A(KEYINPUT28), .B(n1296), .Z(n1293) );
NOR2_X1 U943 ( .A1(n1295), .A2(n1141), .ZN(n1296) );
INV_X1 U944 ( .A(n1249), .ZN(n1295) );
NAND2_X1 U945 ( .A1(n1100), .A2(n1272), .ZN(n1249) );
NOR3_X1 U946 ( .A1(n1248), .A2(n1259), .A3(n1264), .ZN(n1272) );
INV_X1 U947 ( .A(n1173), .ZN(n1264) );
INV_X1 U948 ( .A(n1247), .ZN(n1259) );
NAND2_X1 U949 ( .A1(n1297), .A2(n1298), .ZN(n1247) );
NAND2_X1 U950 ( .A1(n1299), .A2(n1135), .ZN(n1297) );
INV_X1 U951 ( .A(G900), .ZN(n1135) );
XOR2_X1 U952 ( .A(G122), .B(n1209), .Z(G24) );
AND4_X1 U953 ( .A1(n1227), .A2(n1171), .A3(n1126), .A4(n1300), .ZN(n1209) );
INV_X1 U954 ( .A(n1095), .ZN(n1171) );
NAND2_X1 U955 ( .A1(n1301), .A2(n1302), .ZN(n1095) );
XOR2_X1 U956 ( .A(KEYINPUT37), .B(n1303), .Z(n1302) );
XNOR2_X1 U957 ( .A(n1304), .B(n1305), .ZN(G21) );
NAND2_X1 U958 ( .A1(KEYINPUT21), .A2(n1306), .ZN(n1304) );
NAND2_X1 U959 ( .A1(n1226), .A2(n1227), .ZN(n1306) );
AND3_X1 U960 ( .A1(n1114), .A2(n1282), .A3(n1219), .ZN(n1226) );
INV_X1 U961 ( .A(n1301), .ZN(n1282) );
NAND2_X1 U962 ( .A1(n1307), .A2(n1308), .ZN(G18) );
NAND2_X1 U963 ( .A1(G116), .A2(n1211), .ZN(n1308) );
XOR2_X1 U964 ( .A(n1309), .B(KEYINPUT47), .Z(n1307) );
OR2_X1 U965 ( .A1(n1211), .A2(G116), .ZN(n1309) );
NAND3_X1 U966 ( .A1(n1220), .A2(n1277), .A3(n1227), .ZN(n1211) );
AND2_X1 U967 ( .A1(n1100), .A2(n1225), .ZN(n1227) );
INV_X1 U968 ( .A(n1096), .ZN(n1277) );
NAND2_X1 U969 ( .A1(n1310), .A2(n1126), .ZN(n1096) );
XNOR2_X1 U970 ( .A(n1269), .B(KEYINPUT26), .ZN(n1310) );
XNOR2_X1 U971 ( .A(G113), .B(n1311), .ZN(G15) );
NAND3_X1 U972 ( .A1(n1258), .A2(n1312), .A3(n1100), .ZN(n1311) );
NOR2_X1 U973 ( .A1(n1089), .A2(n1241), .ZN(n1100) );
NAND2_X1 U974 ( .A1(n1107), .A2(n1313), .ZN(n1089) );
XNOR2_X1 U975 ( .A(KEYINPUT5), .B(n1225), .ZN(n1312) );
INV_X1 U976 ( .A(n1229), .ZN(n1258) );
NAND2_X1 U977 ( .A1(n1220), .A2(n1173), .ZN(n1229) );
NOR2_X1 U978 ( .A1(n1269), .A2(n1126), .ZN(n1173) );
NOR2_X1 U979 ( .A1(n1303), .A2(n1301), .ZN(n1220) );
XOR2_X1 U980 ( .A(n1114), .B(KEYINPUT39), .Z(n1303) );
NAND3_X1 U981 ( .A1(n1314), .A2(n1315), .A3(n1316), .ZN(G12) );
NAND2_X1 U982 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND3_X1 U983 ( .A1(n1170), .A2(n1319), .A3(n1218), .ZN(n1318) );
NAND2_X1 U984 ( .A1(KEYINPUT29), .A2(n1320), .ZN(n1317) );
XNOR2_X1 U985 ( .A(KEYINPUT58), .B(n1321), .ZN(n1320) );
NAND4_X1 U986 ( .A1(KEYINPUT29), .A2(n1218), .A3(n1322), .A4(n1321), .ZN(n1315) );
AND2_X1 U987 ( .A1(n1319), .A2(n1170), .ZN(n1322) );
INV_X1 U988 ( .A(n1210), .ZN(n1170) );
NAND3_X1 U989 ( .A1(n1222), .A2(n1225), .A3(n1106), .ZN(n1210) );
NOR2_X1 U990 ( .A1(n1108), .A2(n1107), .ZN(n1106) );
NOR2_X1 U991 ( .A1(n1323), .A2(n1120), .ZN(n1107) );
NOR2_X1 U992 ( .A1(n1125), .A2(n1124), .ZN(n1120) );
AND2_X1 U993 ( .A1(n1324), .A2(n1125), .ZN(n1323) );
NAND2_X1 U994 ( .A1(n1325), .A2(n1261), .ZN(n1125) );
XNOR2_X1 U995 ( .A(n1188), .B(n1185), .ZN(n1325) );
XNOR2_X1 U996 ( .A(n1326), .B(n1327), .ZN(n1185) );
XNOR2_X1 U997 ( .A(n1271), .B(G110), .ZN(n1327) );
NAND2_X1 U998 ( .A1(G227), .A2(n1084), .ZN(n1326) );
XOR2_X1 U999 ( .A(n1328), .B(n1329), .Z(n1188) );
NOR2_X1 U1000 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
NOR2_X1 U1001 ( .A1(n1332), .A2(n1138), .ZN(n1331) );
INV_X1 U1002 ( .A(KEYINPUT23), .ZN(n1138) );
XNOR2_X1 U1003 ( .A(n1075), .B(G104), .ZN(n1332) );
NOR2_X1 U1004 ( .A1(KEYINPUT23), .A2(n1333), .ZN(n1330) );
NOR2_X1 U1005 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
XNOR2_X1 U1006 ( .A(n1180), .B(G101), .ZN(n1328) );
XOR2_X1 U1007 ( .A(KEYINPUT56), .B(n1124), .Z(n1324) );
XOR2_X1 U1008 ( .A(G469), .B(KEYINPUT45), .Z(n1124) );
INV_X1 U1009 ( .A(n1313), .ZN(n1108) );
NAND2_X1 U1010 ( .A1(G221), .A2(n1336), .ZN(n1313) );
NAND2_X1 U1011 ( .A1(n1337), .A2(n1298), .ZN(n1225) );
NAND3_X1 U1012 ( .A1(n1338), .A2(n1084), .A3(G952), .ZN(n1298) );
NAND2_X1 U1013 ( .A1(n1299), .A2(n1155), .ZN(n1337) );
XNOR2_X1 U1014 ( .A(G898), .B(KEYINPUT52), .ZN(n1155) );
NOR3_X1 U1015 ( .A1(n1261), .A2(n1086), .A3(n1084), .ZN(n1299) );
INV_X1 U1016 ( .A(n1338), .ZN(n1086) );
NAND2_X1 U1017 ( .A1(G237), .A2(G234), .ZN(n1338) );
INV_X1 U1018 ( .A(n1241), .ZN(n1222) );
NAND2_X1 U1019 ( .A1(n1103), .A2(n1102), .ZN(n1241) );
NAND2_X1 U1020 ( .A1(G214), .A2(n1201), .ZN(n1102) );
NAND2_X1 U1021 ( .A1(n1339), .A2(n1261), .ZN(n1201) );
NAND2_X1 U1022 ( .A1(n1340), .A2(n1341), .ZN(n1103) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1342), .ZN(n1341) );
NAND2_X1 U1024 ( .A1(n1261), .A2(n1343), .ZN(n1342) );
OR2_X1 U1025 ( .A1(n1339), .A2(n1344), .ZN(n1343) );
INV_X1 U1026 ( .A(G237), .ZN(n1339) );
NAND3_X1 U1027 ( .A1(n1345), .A2(n1261), .A3(n1344), .ZN(n1340) );
XOR2_X1 U1028 ( .A(n1346), .B(n1347), .Z(n1344) );
INV_X1 U1029 ( .A(n1196), .ZN(n1347) );
XOR2_X1 U1030 ( .A(n1348), .B(n1152), .Z(n1196) );
XNOR2_X1 U1031 ( .A(G122), .B(G110), .ZN(n1152) );
NAND2_X1 U1032 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1033 ( .A1(n1154), .A2(n1351), .ZN(n1350) );
INV_X1 U1034 ( .A(KEYINPUT27), .ZN(n1351) );
XOR2_X1 U1035 ( .A(n1182), .B(n1352), .Z(n1154) );
NAND3_X1 U1036 ( .A1(n1352), .A2(n1182), .A3(KEYINPUT27), .ZN(n1349) );
AND2_X1 U1037 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
NAND2_X1 U1038 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
XOR2_X1 U1039 ( .A(KEYINPUT19), .B(n1357), .Z(n1353) );
NOR2_X1 U1040 ( .A1(n1355), .A2(n1356), .ZN(n1357) );
XNOR2_X1 U1041 ( .A(n1287), .B(KEYINPUT31), .ZN(n1356) );
INV_X1 U1042 ( .A(G101), .ZN(n1287) );
NOR2_X1 U1043 ( .A1(n1358), .A2(n1335), .ZN(n1355) );
NOR2_X1 U1044 ( .A1(n1359), .A2(G107), .ZN(n1335) );
INV_X1 U1045 ( .A(G104), .ZN(n1359) );
XNOR2_X1 U1046 ( .A(KEYINPUT63), .B(n1334), .ZN(n1358) );
NOR2_X1 U1047 ( .A1(n1075), .A2(G104), .ZN(n1334) );
NAND3_X1 U1048 ( .A1(n1360), .A2(n1361), .A3(n1198), .ZN(n1346) );
NAND2_X1 U1049 ( .A1(n1362), .A2(n1363), .ZN(n1198) );
NAND2_X1 U1050 ( .A1(n1364), .A2(n1365), .ZN(n1361) );
INV_X1 U1051 ( .A(KEYINPUT54), .ZN(n1365) );
NAND3_X1 U1052 ( .A1(n1366), .A2(n1367), .A3(n1368), .ZN(n1364) );
INV_X1 U1053 ( .A(n1362), .ZN(n1368) );
NOR2_X1 U1054 ( .A1(n1141), .A2(n1369), .ZN(n1362) );
NAND2_X1 U1055 ( .A1(n1363), .A2(n1370), .ZN(n1367) );
INV_X1 U1056 ( .A(n1371), .ZN(n1363) );
NAND3_X1 U1057 ( .A1(n1371), .A2(n1141), .A3(n1369), .ZN(n1366) );
NAND2_X1 U1058 ( .A1(KEYINPUT54), .A2(n1199), .ZN(n1360) );
NAND2_X1 U1059 ( .A1(n1372), .A2(n1373), .ZN(n1199) );
NAND2_X1 U1060 ( .A1(n1374), .A2(n1141), .ZN(n1373) );
XNOR2_X1 U1061 ( .A(n1370), .B(n1371), .ZN(n1374) );
NAND3_X1 U1062 ( .A1(n1369), .A2(n1371), .A3(G125), .ZN(n1372) );
XOR2_X1 U1063 ( .A(G143), .B(n1375), .Z(n1371) );
INV_X1 U1064 ( .A(n1370), .ZN(n1369) );
NAND2_X1 U1065 ( .A1(G224), .A2(n1084), .ZN(n1370) );
NAND2_X1 U1066 ( .A1(G210), .A2(G237), .ZN(n1345) );
XOR2_X1 U1067 ( .A(n1219), .B(KEYINPUT51), .Z(n1319) );
NOR2_X1 U1068 ( .A1(n1300), .A2(n1126), .ZN(n1219) );
XOR2_X1 U1069 ( .A(n1376), .B(n1377), .Z(n1126) );
XOR2_X1 U1070 ( .A(KEYINPUT10), .B(G478), .Z(n1377) );
NAND2_X1 U1071 ( .A1(n1165), .A2(n1261), .ZN(n1376) );
XNOR2_X1 U1072 ( .A(n1378), .B(n1379), .ZN(n1165) );
XOR2_X1 U1073 ( .A(n1380), .B(n1381), .Z(n1379) );
XNOR2_X1 U1074 ( .A(G116), .B(n1075), .ZN(n1381) );
INV_X1 U1075 ( .A(G107), .ZN(n1075) );
XNOR2_X1 U1076 ( .A(n1275), .B(G128), .ZN(n1380) );
INV_X1 U1077 ( .A(G134), .ZN(n1275) );
XOR2_X1 U1078 ( .A(n1382), .B(n1383), .Z(n1378) );
XNOR2_X1 U1079 ( .A(n1384), .B(n1385), .ZN(n1383) );
NOR2_X1 U1080 ( .A1(G122), .A2(KEYINPUT15), .ZN(n1385) );
NAND2_X1 U1081 ( .A1(KEYINPUT12), .A2(n1265), .ZN(n1384) );
NAND2_X1 U1082 ( .A1(G217), .A2(n1386), .ZN(n1382) );
INV_X1 U1083 ( .A(n1269), .ZN(n1300) );
XNOR2_X1 U1084 ( .A(n1117), .B(n1387), .ZN(n1269) );
NOR2_X1 U1085 ( .A1(G475), .A2(KEYINPUT53), .ZN(n1387) );
NAND2_X1 U1086 ( .A1(n1168), .A2(n1261), .ZN(n1117) );
XNOR2_X1 U1087 ( .A(n1388), .B(n1389), .ZN(n1168) );
XNOR2_X1 U1088 ( .A(n1390), .B(n1391), .ZN(n1389) );
NAND2_X1 U1089 ( .A1(n1392), .A2(G214), .ZN(n1390) );
XNOR2_X1 U1090 ( .A(n1393), .B(n1394), .ZN(n1388) );
NAND2_X1 U1091 ( .A1(n1395), .A2(KEYINPUT57), .ZN(n1394) );
XNOR2_X1 U1092 ( .A(G104), .B(n1396), .ZN(n1395) );
XOR2_X1 U1093 ( .A(G122), .B(G113), .Z(n1396) );
NAND2_X1 U1094 ( .A1(KEYINPUT62), .A2(n1397), .ZN(n1393) );
XOR2_X1 U1095 ( .A(n1398), .B(n1399), .Z(n1397) );
XNOR2_X1 U1096 ( .A(G146), .B(G125), .ZN(n1399) );
NAND2_X1 U1097 ( .A1(KEYINPUT18), .A2(n1271), .ZN(n1398) );
INV_X1 U1098 ( .A(n1248), .ZN(n1218) );
NAND2_X1 U1099 ( .A1(n1301), .A2(n1114), .ZN(n1248) );
XNOR2_X1 U1100 ( .A(n1400), .B(n1162), .ZN(n1114) );
AND2_X1 U1101 ( .A1(G217), .A2(n1336), .ZN(n1162) );
NAND2_X1 U1102 ( .A1(G234), .A2(n1261), .ZN(n1336) );
OR2_X1 U1103 ( .A1(n1159), .A2(G902), .ZN(n1400) );
XNOR2_X1 U1104 ( .A(n1401), .B(n1402), .ZN(n1159) );
XOR2_X1 U1105 ( .A(G137), .B(n1403), .Z(n1402) );
NOR2_X1 U1106 ( .A1(KEYINPUT20), .A2(n1404), .ZN(n1403) );
XOR2_X1 U1107 ( .A(n1405), .B(n1406), .Z(n1404) );
XNOR2_X1 U1108 ( .A(n1141), .B(n1407), .ZN(n1406) );
XNOR2_X1 U1109 ( .A(KEYINPUT49), .B(n1271), .ZN(n1407) );
INV_X1 U1110 ( .A(G140), .ZN(n1271) );
INV_X1 U1111 ( .A(G125), .ZN(n1141) );
XOR2_X1 U1112 ( .A(n1408), .B(n1375), .Z(n1405) );
XNOR2_X1 U1113 ( .A(G119), .B(G110), .ZN(n1408) );
NAND2_X1 U1114 ( .A1(n1386), .A2(G221), .ZN(n1401) );
AND2_X1 U1115 ( .A1(G234), .A2(n1084), .ZN(n1386) );
INV_X1 U1116 ( .A(G953), .ZN(n1084) );
NOR2_X1 U1117 ( .A1(n1409), .A2(n1118), .ZN(n1301) );
NOR2_X1 U1118 ( .A1(n1123), .A2(G472), .ZN(n1118) );
AND2_X1 U1119 ( .A1(G472), .A2(n1123), .ZN(n1409) );
NAND2_X1 U1120 ( .A1(n1410), .A2(n1261), .ZN(n1123) );
INV_X1 U1121 ( .A(G902), .ZN(n1261) );
NAND2_X1 U1122 ( .A1(n1411), .A2(n1412), .ZN(n1410) );
OR2_X1 U1123 ( .A1(n1413), .A2(n1414), .ZN(n1412) );
XOR2_X1 U1124 ( .A(n1415), .B(KEYINPUT8), .Z(n1411) );
NAND2_X1 U1125 ( .A1(n1414), .A2(n1413), .ZN(n1415) );
NAND2_X1 U1126 ( .A1(n1416), .A2(n1417), .ZN(n1413) );
OR2_X1 U1127 ( .A1(n1418), .A2(n1182), .ZN(n1417) );
XOR2_X1 U1128 ( .A(n1419), .B(KEYINPUT6), .Z(n1416) );
NAND2_X1 U1129 ( .A1(n1418), .A2(n1182), .ZN(n1419) );
XOR2_X1 U1130 ( .A(G113), .B(n1420), .Z(n1182) );
XNOR2_X1 U1131 ( .A(n1305), .B(G116), .ZN(n1420) );
INV_X1 U1132 ( .A(G119), .ZN(n1305) );
XOR2_X1 U1133 ( .A(n1180), .B(KEYINPUT42), .Z(n1418) );
XOR2_X1 U1134 ( .A(n1140), .B(KEYINPUT60), .Z(n1180) );
XNOR2_X1 U1135 ( .A(n1421), .B(n1422), .ZN(n1140) );
XOR2_X1 U1136 ( .A(n1375), .B(n1391), .Z(n1422) );
XNOR2_X1 U1137 ( .A(G131), .B(n1265), .ZN(n1391) );
INV_X1 U1138 ( .A(G143), .ZN(n1265) );
XOR2_X1 U1139 ( .A(G128), .B(G146), .Z(n1375) );
XNOR2_X1 U1140 ( .A(G134), .B(G137), .ZN(n1421) );
XNOR2_X1 U1141 ( .A(n1423), .B(n1424), .ZN(n1414) );
NOR2_X1 U1142 ( .A1(KEYINPUT25), .A2(n1177), .ZN(n1424) );
NAND2_X1 U1143 ( .A1(n1392), .A2(G210), .ZN(n1177) );
NOR2_X1 U1144 ( .A1(G953), .A2(G237), .ZN(n1392) );
XNOR2_X1 U1145 ( .A(G101), .B(KEYINPUT14), .ZN(n1423) );
OR2_X1 U1146 ( .A1(n1321), .A2(KEYINPUT29), .ZN(n1314) );
INV_X1 U1147 ( .A(G110), .ZN(n1321) );
endmodule


