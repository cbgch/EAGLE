//Key = 0010011001011111100000011100101010101100100001111011010001111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346;

XOR2_X1 U738 ( .A(G107), .B(n1024), .Z(G9) );
NOR2_X1 U739 ( .A1(n1025), .A2(n1026), .ZN(G75) );
NOR4_X1 U740 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
NOR2_X1 U741 ( .A1(n1031), .A2(n1032), .ZN(n1028) );
NOR2_X1 U742 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U743 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
INV_X1 U744 ( .A(n1037), .ZN(n1036) );
NOR2_X1 U745 ( .A1(n1038), .A2(n1039), .ZN(n1035) );
NOR2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR3_X1 U747 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1040) );
AND3_X1 U748 ( .A1(n1045), .A2(n1046), .A3(KEYINPUT44), .ZN(n1044) );
NOR2_X1 U749 ( .A1(n1047), .A2(n1045), .ZN(n1043) );
NOR3_X1 U750 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
NOR3_X1 U751 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1050) );
INV_X1 U752 ( .A(KEYINPUT9), .ZN(n1051) );
NOR2_X1 U753 ( .A1(KEYINPUT9), .A2(n1054), .ZN(n1049) );
NOR2_X1 U754 ( .A1(KEYINPUT44), .A2(n1055), .ZN(n1048) );
NOR3_X1 U755 ( .A1(n1054), .A2(n1056), .A3(n1057), .ZN(n1042) );
NOR2_X1 U756 ( .A1(n1058), .A2(n1054), .ZN(n1038) );
NOR2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR2_X1 U758 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
XOR2_X1 U759 ( .A(KEYINPUT37), .B(n1063), .Z(n1062) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1045), .ZN(n1059) );
NOR2_X1 U761 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR4_X1 U762 ( .A1(n1067), .A2(n1041), .A3(n1054), .A4(n1045), .ZN(n1033) );
INV_X1 U763 ( .A(n1063), .ZN(n1041) );
NOR2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR3_X1 U765 ( .A1(n1029), .A2(G952), .A3(n1027), .ZN(n1025) );
AND3_X1 U766 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1027) );
AND3_X1 U767 ( .A1(n1073), .A2(n1056), .A3(n1053), .ZN(n1072) );
XOR2_X1 U768 ( .A(n1074), .B(KEYINPUT51), .Z(n1071) );
NAND4_X1 U769 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
NOR2_X1 U770 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
XOR2_X1 U771 ( .A(n1081), .B(n1082), .Z(n1080) );
NOR2_X1 U772 ( .A1(n1083), .A2(KEYINPUT55), .ZN(n1082) );
NOR2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1079) );
XOR2_X1 U774 ( .A(n1086), .B(KEYINPUT63), .Z(n1076) );
NAND2_X1 U775 ( .A1(n1085), .A2(n1084), .ZN(n1086) );
INV_X1 U776 ( .A(G472), .ZN(n1084) );
XNOR2_X1 U777 ( .A(n1087), .B(KEYINPUT1), .ZN(n1085) );
XNOR2_X1 U778 ( .A(n1088), .B(G475), .ZN(n1075) );
XNOR2_X1 U779 ( .A(n1089), .B(G469), .ZN(n1070) );
XOR2_X1 U780 ( .A(n1090), .B(n1091), .Z(G72) );
XOR2_X1 U781 ( .A(n1092), .B(n1093), .Z(n1091) );
NOR2_X1 U782 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NOR2_X1 U783 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NAND2_X1 U784 ( .A1(n1098), .A2(n1099), .ZN(n1092) );
NAND2_X1 U785 ( .A1(G953), .A2(n1097), .ZN(n1099) );
XOR2_X1 U786 ( .A(n1100), .B(n1101), .Z(n1098) );
XOR2_X1 U787 ( .A(G125), .B(n1102), .Z(n1101) );
XOR2_X1 U788 ( .A(KEYINPUT62), .B(G140), .Z(n1102) );
XOR2_X1 U789 ( .A(n1103), .B(n1104), .Z(n1100) );
NAND2_X1 U790 ( .A1(n1095), .A2(n1105), .ZN(n1090) );
NAND2_X1 U791 ( .A1(n1106), .A2(n1107), .ZN(G69) );
NAND2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U793 ( .A1(G953), .A2(n1110), .ZN(n1109) );
NAND3_X1 U794 ( .A1(G953), .A2(n1111), .A3(n1112), .ZN(n1106) );
XNOR2_X1 U795 ( .A(n1108), .B(KEYINPUT8), .ZN(n1112) );
XNOR2_X1 U796 ( .A(n1113), .B(n1114), .ZN(n1108) );
AND2_X1 U797 ( .A1(n1095), .A2(n1115), .ZN(n1114) );
NAND2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1113) );
NAND2_X1 U799 ( .A1(G953), .A2(n1118), .ZN(n1117) );
XOR2_X1 U800 ( .A(n1119), .B(n1120), .Z(n1116) );
XNOR2_X1 U801 ( .A(n1121), .B(n1122), .ZN(n1120) );
NOR2_X1 U802 ( .A1(KEYINPUT52), .A2(n1123), .ZN(n1119) );
NAND2_X1 U803 ( .A1(G898), .A2(G224), .ZN(n1111) );
NOR2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XOR2_X1 U805 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U806 ( .A(n1128), .B(KEYINPUT4), .Z(n1126) );
NAND2_X1 U807 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XOR2_X1 U808 ( .A(KEYINPUT54), .B(n1083), .Z(n1130) );
NOR2_X1 U809 ( .A1(G952), .A2(n1131), .ZN(n1124) );
XOR2_X1 U810 ( .A(KEYINPUT47), .B(G953), .Z(n1131) );
NOR2_X1 U811 ( .A1(n1132), .A2(n1133), .ZN(G63) );
XOR2_X1 U812 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U813 ( .A(n1136), .B(KEYINPUT45), .Z(n1134) );
NAND2_X1 U814 ( .A1(n1129), .A2(G478), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1132), .A2(n1137), .ZN(G60) );
NOR3_X1 U816 ( .A1(n1088), .A2(n1138), .A3(n1139), .ZN(n1137) );
AND3_X1 U817 ( .A1(n1140), .A2(G475), .A3(n1129), .ZN(n1139) );
NOR2_X1 U818 ( .A1(n1141), .A2(n1140), .ZN(n1138) );
AND2_X1 U819 ( .A1(n1030), .A2(G475), .ZN(n1141) );
XOR2_X1 U820 ( .A(G104), .B(n1142), .Z(G6) );
NOR2_X1 U821 ( .A1(n1132), .A2(n1143), .ZN(G57) );
NOR2_X1 U822 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U823 ( .A(KEYINPUT56), .B(n1146), .Z(n1145) );
NOR2_X1 U824 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XNOR2_X1 U825 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR2_X1 U826 ( .A1(n1151), .A2(n1152), .ZN(n1144) );
INV_X1 U827 ( .A(n1147), .ZN(n1152) );
XOR2_X1 U828 ( .A(n1153), .B(G101), .Z(n1147) );
XOR2_X1 U829 ( .A(n1149), .B(n1150), .Z(n1151) );
NOR2_X1 U830 ( .A1(KEYINPUT27), .A2(n1154), .ZN(n1150) );
XOR2_X1 U831 ( .A(KEYINPUT40), .B(n1155), .Z(n1154) );
NAND2_X1 U832 ( .A1(n1129), .A2(G472), .ZN(n1149) );
NOR2_X1 U833 ( .A1(n1132), .A2(n1156), .ZN(G54) );
XOR2_X1 U834 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U835 ( .A1(KEYINPUT61), .A2(n1159), .ZN(n1158) );
NOR2_X1 U836 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U837 ( .A(n1162), .B(KEYINPUT59), .Z(n1161) );
NAND2_X1 U838 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U839 ( .A1(n1163), .A2(n1164), .ZN(n1160) );
XNOR2_X1 U840 ( .A(n1165), .B(n1166), .ZN(n1164) );
NAND2_X1 U841 ( .A1(KEYINPUT11), .A2(n1167), .ZN(n1165) );
XNOR2_X1 U842 ( .A(n1168), .B(n1169), .ZN(n1167) );
XOR2_X1 U843 ( .A(n1103), .B(KEYINPUT19), .Z(n1169) );
NAND2_X1 U844 ( .A1(n1129), .A2(G469), .ZN(n1157) );
INV_X1 U845 ( .A(n1170), .ZN(n1129) );
NOR2_X1 U846 ( .A1(n1132), .A2(n1171), .ZN(G51) );
XOR2_X1 U847 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U848 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U849 ( .A(KEYINPUT57), .B(n1176), .Z(n1175) );
NOR2_X1 U850 ( .A1(n1170), .A2(n1177), .ZN(n1176) );
XOR2_X1 U851 ( .A(KEYINPUT28), .B(G210), .Z(n1177) );
NAND2_X1 U852 ( .A1(G902), .A2(n1030), .ZN(n1170) );
OR2_X1 U853 ( .A1(n1105), .A2(n1115), .ZN(n1030) );
NAND4_X1 U854 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1115) );
NOR4_X1 U855 ( .A1(n1142), .A2(n1024), .A3(n1182), .A4(n1183), .ZN(n1181) );
INV_X1 U856 ( .A(n1184), .ZN(n1182) );
AND2_X1 U857 ( .A1(n1068), .A2(n1185), .ZN(n1024) );
AND2_X1 U858 ( .A1(n1069), .A2(n1185), .ZN(n1142) );
AND3_X1 U859 ( .A1(n1063), .A2(n1186), .A3(n1187), .ZN(n1185) );
NOR2_X1 U860 ( .A1(n1188), .A2(n1189), .ZN(n1180) );
NOR2_X1 U861 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U862 ( .A1(n1061), .A2(n1192), .ZN(n1188) );
NAND3_X1 U863 ( .A1(n1193), .A2(n1186), .A3(n1066), .ZN(n1178) );
NAND2_X1 U864 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NAND4_X1 U865 ( .A1(n1069), .A2(n1196), .A3(n1061), .A4(n1191), .ZN(n1195) );
INV_X1 U866 ( .A(KEYINPUT60), .ZN(n1191) );
NAND2_X1 U867 ( .A1(n1037), .A2(n1187), .ZN(n1194) );
NAND2_X1 U868 ( .A1(n1197), .A2(n1198), .ZN(n1105) );
AND4_X1 U869 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1198) );
NOR4_X1 U870 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1197) );
NOR2_X1 U871 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
AND2_X1 U872 ( .A1(n1209), .A2(n1210), .ZN(n1205) );
XNOR2_X1 U873 ( .A(n1211), .B(n1212), .ZN(n1172) );
NOR2_X1 U874 ( .A1(n1095), .A2(G952), .ZN(n1132) );
XOR2_X1 U875 ( .A(G146), .B(n1204), .Z(G48) );
AND2_X1 U876 ( .A1(n1213), .A2(n1069), .ZN(n1204) );
XOR2_X1 U877 ( .A(G143), .B(n1214), .Z(G45) );
NOR2_X1 U878 ( .A1(n1208), .A2(n1215), .ZN(n1214) );
XOR2_X1 U879 ( .A(KEYINPUT24), .B(n1066), .Z(n1215) );
NAND4_X1 U880 ( .A1(n1216), .A2(n1187), .A3(n1217), .A4(n1218), .ZN(n1208) );
XOR2_X1 U881 ( .A(G140), .B(n1203), .Z(G42) );
AND3_X1 U882 ( .A1(n1069), .A2(n1065), .A3(n1209), .ZN(n1203) );
XOR2_X1 U883 ( .A(n1219), .B(n1220), .Z(G39) );
XNOR2_X1 U884 ( .A(G137), .B(KEYINPUT26), .ZN(n1220) );
NAND4_X1 U885 ( .A1(n1210), .A2(n1221), .A3(n1222), .A4(n1218), .ZN(n1219) );
XOR2_X1 U886 ( .A(KEYINPUT3), .B(n1046), .Z(n1222) );
INV_X1 U887 ( .A(n1045), .ZN(n1221) );
XNOR2_X1 U888 ( .A(G134), .B(n1202), .ZN(G36) );
NAND3_X1 U889 ( .A1(n1209), .A2(n1068), .A3(n1066), .ZN(n1202) );
XOR2_X1 U890 ( .A(n1223), .B(n1201), .Z(G33) );
NAND3_X1 U891 ( .A1(n1209), .A2(n1069), .A3(n1066), .ZN(n1201) );
NOR3_X1 U892 ( .A1(n1055), .A2(n1224), .A3(n1045), .ZN(n1209) );
NAND2_X1 U893 ( .A1(n1073), .A2(n1225), .ZN(n1045) );
INV_X1 U894 ( .A(n1057), .ZN(n1073) );
XOR2_X1 U895 ( .A(n1226), .B(n1200), .Z(G30) );
NAND2_X1 U896 ( .A1(n1213), .A2(n1068), .ZN(n1200) );
AND4_X1 U897 ( .A1(n1187), .A2(n1227), .A3(n1228), .A4(n1218), .ZN(n1213) );
XOR2_X1 U898 ( .A(n1229), .B(n1230), .Z(G3) );
NAND4_X1 U899 ( .A1(n1037), .A2(n1066), .A3(n1231), .A4(n1046), .ZN(n1230) );
INV_X1 U900 ( .A(n1055), .ZN(n1046) );
NOR2_X1 U901 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
XOR2_X1 U902 ( .A(n1061), .B(KEYINPUT38), .Z(n1233) );
XNOR2_X1 U903 ( .A(G125), .B(n1199), .ZN(G27) );
NAND4_X1 U904 ( .A1(n1069), .A2(n1196), .A3(n1234), .A4(n1065), .ZN(n1199) );
NOR2_X1 U905 ( .A1(n1224), .A2(n1061), .ZN(n1234) );
INV_X1 U906 ( .A(n1218), .ZN(n1224) );
NAND2_X1 U907 ( .A1(n1032), .A2(n1235), .ZN(n1218) );
NAND4_X1 U908 ( .A1(G953), .A2(G902), .A3(n1236), .A4(n1097), .ZN(n1235) );
INV_X1 U909 ( .A(G900), .ZN(n1097) );
XOR2_X1 U910 ( .A(n1237), .B(n1179), .Z(G24) );
NAND4_X1 U911 ( .A1(n1216), .A2(n1238), .A3(n1063), .A4(n1217), .ZN(n1179) );
NOR2_X1 U912 ( .A1(n1228), .A2(n1227), .ZN(n1063) );
XOR2_X1 U913 ( .A(G119), .B(n1183), .Z(G21) );
AND2_X1 U914 ( .A1(n1238), .A2(n1210), .ZN(n1183) );
AND3_X1 U915 ( .A1(n1227), .A2(n1228), .A3(n1037), .ZN(n1210) );
INV_X1 U916 ( .A(n1239), .ZN(n1227) );
XNOR2_X1 U917 ( .A(G116), .B(n1240), .ZN(G18) );
NOR2_X1 U918 ( .A1(KEYINPUT10), .A2(n1241), .ZN(n1240) );
NOR2_X1 U919 ( .A1(n1242), .A2(n1061), .ZN(n1241) );
XOR2_X1 U920 ( .A(n1192), .B(KEYINPUT33), .Z(n1242) );
NAND4_X1 U921 ( .A1(n1066), .A2(n1196), .A3(n1068), .A4(n1186), .ZN(n1192) );
NOR2_X1 U922 ( .A1(n1078), .A2(n1216), .ZN(n1068) );
XNOR2_X1 U923 ( .A(G113), .B(n1190), .ZN(G15) );
NAND3_X1 U924 ( .A1(n1066), .A2(n1069), .A3(n1238), .ZN(n1190) );
NOR3_X1 U925 ( .A1(n1061), .A2(n1232), .A3(n1054), .ZN(n1238) );
INV_X1 U926 ( .A(n1196), .ZN(n1054) );
NOR2_X1 U927 ( .A1(n1052), .A2(n1243), .ZN(n1196) );
INV_X1 U928 ( .A(n1053), .ZN(n1243) );
INV_X1 U929 ( .A(n1186), .ZN(n1232) );
AND2_X1 U930 ( .A1(n1216), .A2(n1078), .ZN(n1069) );
INV_X1 U931 ( .A(n1207), .ZN(n1066) );
NAND2_X1 U932 ( .A1(n1239), .A2(n1228), .ZN(n1207) );
XOR2_X1 U933 ( .A(n1244), .B(n1184), .Z(G12) );
NAND4_X1 U934 ( .A1(n1037), .A2(n1065), .A3(n1187), .A4(n1186), .ZN(n1184) );
NAND2_X1 U935 ( .A1(n1032), .A2(n1245), .ZN(n1186) );
NAND4_X1 U936 ( .A1(G953), .A2(G902), .A3(n1236), .A4(n1118), .ZN(n1245) );
INV_X1 U937 ( .A(G898), .ZN(n1118) );
NAND3_X1 U938 ( .A1(n1246), .A2(n1236), .A3(G952), .ZN(n1032) );
NAND2_X1 U939 ( .A1(G237), .A2(G234), .ZN(n1236) );
INV_X1 U940 ( .A(n1029), .ZN(n1246) );
XOR2_X1 U941 ( .A(n1095), .B(KEYINPUT25), .Z(n1029) );
NOR2_X1 U942 ( .A1(n1055), .A2(n1061), .ZN(n1187) );
NAND2_X1 U943 ( .A1(n1225), .A2(n1057), .ZN(n1061) );
NAND3_X1 U944 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(n1057) );
OR2_X1 U945 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NAND3_X1 U946 ( .A1(n1251), .A2(n1250), .A3(n1252), .ZN(n1248) );
NAND2_X1 U947 ( .A1(G237), .A2(G210), .ZN(n1250) );
XNOR2_X1 U948 ( .A(n1211), .B(n1253), .ZN(n1251) );
XNOR2_X1 U949 ( .A(n1254), .B(KEYINPUT39), .ZN(n1253) );
NAND4_X1 U950 ( .A1(KEYINPUT46), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1254) );
NAND2_X1 U951 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
INV_X1 U952 ( .A(KEYINPUT34), .ZN(n1259) );
NAND2_X1 U953 ( .A1(n1174), .A2(n1260), .ZN(n1258) );
XNOR2_X1 U954 ( .A(KEYINPUT15), .B(n1212), .ZN(n1260) );
NAND2_X1 U955 ( .A1(KEYINPUT34), .A2(n1261), .ZN(n1256) );
NAND2_X1 U956 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NAND3_X1 U957 ( .A1(KEYINPUT15), .A2(n1174), .A3(n1212), .ZN(n1263) );
OR2_X1 U958 ( .A1(n1212), .A2(KEYINPUT15), .ZN(n1262) );
OR2_X1 U959 ( .A1(n1212), .A2(n1174), .ZN(n1255) );
NOR2_X1 U960 ( .A1(n1110), .A2(G953), .ZN(n1174) );
INV_X1 U961 ( .A(G224), .ZN(n1110) );
XNOR2_X1 U962 ( .A(n1264), .B(n1265), .ZN(n1212) );
XOR2_X1 U963 ( .A(n1266), .B(n1267), .Z(n1211) );
XNOR2_X1 U964 ( .A(n1268), .B(n1123), .ZN(n1267) );
XNOR2_X1 U965 ( .A(n1229), .B(n1269), .ZN(n1123) );
NOR2_X1 U966 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NOR2_X1 U967 ( .A1(KEYINPUT48), .A2(n1272), .ZN(n1271) );
INV_X1 U968 ( .A(n1273), .ZN(n1272) );
NOR2_X1 U969 ( .A1(KEYINPUT17), .A2(n1273), .ZN(n1270) );
NAND2_X1 U970 ( .A1(KEYINPUT12), .A2(n1121), .ZN(n1268) );
AND2_X1 U971 ( .A1(n1274), .A2(n1275), .ZN(n1121) );
NAND2_X1 U972 ( .A1(G110), .A2(n1237), .ZN(n1275) );
XOR2_X1 U973 ( .A(n1276), .B(KEYINPUT0), .Z(n1274) );
NAND2_X1 U974 ( .A1(G122), .A2(n1244), .ZN(n1276) );
XOR2_X1 U975 ( .A(n1122), .B(KEYINPUT13), .Z(n1266) );
NAND2_X1 U976 ( .A1(n1277), .A2(n1278), .ZN(n1122) );
NAND2_X1 U977 ( .A1(G113), .A2(n1279), .ZN(n1278) );
XOR2_X1 U978 ( .A(KEYINPUT30), .B(n1280), .Z(n1277) );
NOR2_X1 U979 ( .A1(G113), .A2(n1279), .ZN(n1280) );
NAND2_X1 U980 ( .A1(G902), .A2(G210), .ZN(n1247) );
XNOR2_X1 U981 ( .A(n1056), .B(KEYINPUT14), .ZN(n1225) );
NAND2_X1 U982 ( .A1(G214), .A2(n1281), .ZN(n1056) );
NAND2_X1 U983 ( .A1(n1252), .A2(n1282), .ZN(n1281) );
NAND2_X1 U984 ( .A1(n1052), .A2(n1053), .ZN(n1055) );
NAND2_X1 U985 ( .A1(G221), .A2(n1283), .ZN(n1053) );
XNOR2_X1 U986 ( .A(n1284), .B(G469), .ZN(n1052) );
NAND2_X1 U987 ( .A1(KEYINPUT58), .A2(n1089), .ZN(n1284) );
AND2_X1 U988 ( .A1(n1285), .A2(n1252), .ZN(n1089) );
XOR2_X1 U989 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U990 ( .A(n1288), .B(n1289), .ZN(n1287) );
NOR2_X1 U991 ( .A1(KEYINPUT7), .A2(n1163), .ZN(n1289) );
AND2_X1 U992 ( .A1(n1290), .A2(n1291), .ZN(n1163) );
NAND2_X1 U993 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND2_X1 U994 ( .A1(G227), .A2(n1095), .ZN(n1293) );
OR3_X1 U995 ( .A1(n1096), .A2(G953), .A3(n1292), .ZN(n1290) );
INV_X1 U996 ( .A(G227), .ZN(n1096) );
NAND2_X1 U997 ( .A1(KEYINPUT6), .A2(n1103), .ZN(n1288) );
XOR2_X1 U998 ( .A(n1294), .B(n1295), .Z(n1103) );
XOR2_X1 U999 ( .A(KEYINPUT5), .B(G128), .Z(n1295) );
NAND3_X1 U1000 ( .A1(n1296), .A2(n1297), .A3(n1298), .ZN(n1294) );
OR2_X1 U1001 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
NAND3_X1 U1002 ( .A1(n1300), .A2(n1299), .A3(KEYINPUT32), .ZN(n1297) );
NOR2_X1 U1003 ( .A1(KEYINPUT43), .A2(n1301), .ZN(n1300) );
NAND2_X1 U1004 ( .A1(n1301), .A2(n1302), .ZN(n1296) );
INV_X1 U1005 ( .A(KEYINPUT32), .ZN(n1302) );
XOR2_X1 U1006 ( .A(n1303), .B(KEYINPUT2), .Z(n1301) );
INV_X1 U1007 ( .A(G143), .ZN(n1303) );
XNOR2_X1 U1008 ( .A(n1166), .B(n1168), .ZN(n1286) );
XOR2_X1 U1009 ( .A(n1229), .B(n1273), .Z(n1168) );
XNOR2_X1 U1010 ( .A(G104), .B(G107), .ZN(n1273) );
NOR2_X1 U1011 ( .A1(n1228), .A2(n1239), .ZN(n1065) );
XOR2_X1 U1012 ( .A(n1304), .B(n1083), .Z(n1239) );
AND2_X1 U1013 ( .A1(G217), .A2(n1283), .ZN(n1083) );
NAND2_X1 U1014 ( .A1(G234), .A2(n1252), .ZN(n1283) );
XOR2_X1 U1015 ( .A(n1081), .B(KEYINPUT42), .Z(n1304) );
NAND2_X1 U1016 ( .A1(n1127), .A2(n1252), .ZN(n1081) );
XNOR2_X1 U1017 ( .A(n1305), .B(n1306), .ZN(n1127) );
XOR2_X1 U1018 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U1019 ( .A(G119), .B(G137), .ZN(n1308) );
NAND2_X1 U1020 ( .A1(G221), .A2(n1309), .ZN(n1307) );
XNOR2_X1 U1021 ( .A(n1292), .B(n1310), .ZN(n1305) );
XOR2_X1 U1022 ( .A(n1311), .B(n1265), .Z(n1310) );
XOR2_X1 U1023 ( .A(G125), .B(G146), .Z(n1265) );
NOR2_X1 U1024 ( .A1(KEYINPUT29), .A2(n1226), .ZN(n1311) );
XNOR2_X1 U1025 ( .A(n1244), .B(G140), .ZN(n1292) );
XNOR2_X1 U1026 ( .A(n1087), .B(G472), .ZN(n1228) );
NAND2_X1 U1027 ( .A1(n1312), .A2(n1252), .ZN(n1087) );
INV_X1 U1028 ( .A(G902), .ZN(n1252) );
XOR2_X1 U1029 ( .A(n1313), .B(n1314), .Z(n1312) );
XNOR2_X1 U1030 ( .A(n1315), .B(KEYINPUT22), .ZN(n1314) );
NAND2_X1 U1031 ( .A1(KEYINPUT50), .A2(n1229), .ZN(n1315) );
INV_X1 U1032 ( .A(G101), .ZN(n1229) );
XOR2_X1 U1033 ( .A(n1155), .B(n1153), .Z(n1313) );
NAND3_X1 U1034 ( .A1(G210), .A2(n1095), .A3(n1316), .ZN(n1153) );
XOR2_X1 U1035 ( .A(n1282), .B(KEYINPUT20), .Z(n1316) );
XNOR2_X1 U1036 ( .A(n1317), .B(n1318), .ZN(n1155) );
XOR2_X1 U1037 ( .A(n1319), .B(n1320), .Z(n1318) );
XOR2_X1 U1038 ( .A(G113), .B(n1299), .Z(n1320) );
INV_X1 U1039 ( .A(G146), .ZN(n1299) );
NAND2_X1 U1040 ( .A1(KEYINPUT23), .A2(n1321), .ZN(n1319) );
INV_X1 U1041 ( .A(n1279), .ZN(n1321) );
XOR2_X1 U1042 ( .A(G119), .B(G116), .Z(n1279) );
XNOR2_X1 U1043 ( .A(n1166), .B(n1264), .ZN(n1317) );
XOR2_X1 U1044 ( .A(n1104), .B(KEYINPUT53), .Z(n1166) );
XNOR2_X1 U1045 ( .A(n1223), .B(n1322), .ZN(n1104) );
XOR2_X1 U1046 ( .A(G137), .B(G134), .Z(n1322) );
NOR2_X1 U1047 ( .A1(n1217), .A2(n1216), .ZN(n1037) );
XNOR2_X1 U1048 ( .A(n1088), .B(n1323), .ZN(n1216) );
NOR2_X1 U1049 ( .A1(G475), .A2(KEYINPUT21), .ZN(n1323) );
NOR2_X1 U1050 ( .A1(n1140), .A2(G902), .ZN(n1088) );
XOR2_X1 U1051 ( .A(n1324), .B(G125), .Z(n1140) );
XOR2_X1 U1052 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1053 ( .A(n1327), .B(n1328), .Z(n1326) );
XOR2_X1 U1054 ( .A(G143), .B(G104), .Z(n1328) );
XOR2_X1 U1055 ( .A(KEYINPUT18), .B(G146), .Z(n1327) );
XOR2_X1 U1056 ( .A(n1329), .B(n1330), .Z(n1325) );
XNOR2_X1 U1057 ( .A(n1331), .B(n1332), .ZN(n1330) );
NOR2_X1 U1058 ( .A1(G140), .A2(KEYINPUT35), .ZN(n1332) );
NAND2_X1 U1059 ( .A1(KEYINPUT16), .A2(n1223), .ZN(n1331) );
INV_X1 U1060 ( .A(G131), .ZN(n1223) );
XOR2_X1 U1061 ( .A(n1333), .B(n1334), .Z(n1329) );
NOR2_X1 U1062 ( .A1(KEYINPUT41), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1063 ( .A(G113), .B(n1237), .Z(n1335) );
NAND3_X1 U1064 ( .A1(n1282), .A2(n1095), .A3(G214), .ZN(n1333) );
INV_X1 U1065 ( .A(G237), .ZN(n1282) );
INV_X1 U1066 ( .A(n1078), .ZN(n1217) );
XOR2_X1 U1067 ( .A(n1336), .B(G478), .Z(n1078) );
OR2_X1 U1068 ( .A1(n1135), .A2(G902), .ZN(n1336) );
XNOR2_X1 U1069 ( .A(n1337), .B(n1338), .ZN(n1135) );
XOR2_X1 U1070 ( .A(G134), .B(n1339), .Z(n1338) );
NOR2_X1 U1071 ( .A1(KEYINPUT49), .A2(n1340), .ZN(n1339) );
XOR2_X1 U1072 ( .A(G107), .B(n1341), .Z(n1340) );
NOR3_X1 U1073 ( .A1(KEYINPUT31), .A2(n1342), .A3(n1343), .ZN(n1341) );
NOR3_X1 U1074 ( .A1(KEYINPUT36), .A2(G116), .A3(n1237), .ZN(n1343) );
INV_X1 U1075 ( .A(G122), .ZN(n1237) );
NOR2_X1 U1076 ( .A1(n1344), .A2(n1345), .ZN(n1342) );
INV_X1 U1077 ( .A(KEYINPUT36), .ZN(n1345) );
XOR2_X1 U1078 ( .A(G122), .B(G116), .Z(n1344) );
XOR2_X1 U1079 ( .A(n1346), .B(n1264), .Z(n1337) );
XNOR2_X1 U1080 ( .A(n1226), .B(G143), .ZN(n1264) );
INV_X1 U1081 ( .A(G128), .ZN(n1226) );
NAND2_X1 U1082 ( .A1(G217), .A2(n1309), .ZN(n1346) );
AND2_X1 U1083 ( .A1(G234), .A2(n1095), .ZN(n1309) );
INV_X1 U1084 ( .A(G953), .ZN(n1095) );
INV_X1 U1085 ( .A(G110), .ZN(n1244) );
endmodule


