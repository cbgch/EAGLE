//Key = 1110000000001100111111001111011111001110111001111100001000000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307;

XOR2_X1 U720 ( .A(G107), .B(n997), .Z(G9) );
NOR2_X1 U721 ( .A1(n998), .A2(n999), .ZN(G75) );
NOR4_X1 U722 ( .A1(n1000), .A2(n1001), .A3(G953), .A4(n1002), .ZN(n999) );
AND3_X1 U723 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1001) );
NAND3_X1 U724 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n1000) );
XOR2_X1 U725 ( .A(n1009), .B(KEYINPUT46), .Z(n1008) );
NAND2_X1 U726 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND3_X1 U727 ( .A1(n1012), .A2(n1013), .A3(n1003), .ZN(n1011) );
NAND2_X1 U728 ( .A1(n1005), .A2(n1014), .ZN(n1010) );
NAND2_X1 U729 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U730 ( .A1(n1003), .A2(n1017), .ZN(n1016) );
AND3_X1 U731 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1003) );
NAND3_X1 U732 ( .A1(n1013), .A2(n1021), .A3(n1020), .ZN(n1015) );
NAND2_X1 U733 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND3_X1 U734 ( .A1(n1024), .A2(n1018), .A3(n1025), .ZN(n1023) );
NAND2_X1 U735 ( .A1(n1026), .A2(n1019), .ZN(n1022) );
XOR2_X1 U736 ( .A(n1027), .B(KEYINPUT13), .Z(n1026) );
NAND2_X1 U737 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND3_X1 U738 ( .A1(n1013), .A2(n1030), .A3(n1020), .ZN(n1007) );
INV_X1 U739 ( .A(n1031), .ZN(n1020) );
NAND2_X1 U740 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NAND3_X1 U741 ( .A1(n1034), .A2(n1019), .A3(n1035), .ZN(n1033) );
XNOR2_X1 U742 ( .A(n1018), .B(KEYINPUT24), .ZN(n1035) );
NAND2_X1 U743 ( .A1(n1005), .A2(n1036), .ZN(n1032) );
NAND2_X1 U744 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U745 ( .A1(n1018), .A2(n1039), .ZN(n1038) );
XNOR2_X1 U746 ( .A(KEYINPUT7), .B(n1040), .ZN(n1039) );
NAND2_X1 U747 ( .A1(n1019), .A2(n1041), .ZN(n1037) );
NOR3_X1 U748 ( .A1(n1002), .A2(G953), .A3(G952), .ZN(n998) );
AND4_X1 U749 ( .A1(n1042), .A2(n1019), .A3(n1018), .A4(n1043), .ZN(n1002) );
NOR4_X1 U750 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
XOR2_X1 U751 ( .A(n1048), .B(KEYINPUT40), .Z(n1046) );
XOR2_X1 U752 ( .A(n1049), .B(n1050), .Z(G72) );
XOR2_X1 U753 ( .A(n1051), .B(n1052), .Z(n1050) );
NAND2_X1 U754 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U755 ( .A1(G953), .A2(n1055), .ZN(n1054) );
XOR2_X1 U756 ( .A(n1056), .B(n1057), .Z(n1053) );
XOR2_X1 U757 ( .A(n1058), .B(n1059), .Z(n1057) );
NOR2_X1 U758 ( .A1(G140), .A2(KEYINPUT22), .ZN(n1058) );
XNOR2_X1 U759 ( .A(n1060), .B(n1061), .ZN(n1056) );
NOR2_X1 U760 ( .A1(KEYINPUT44), .A2(n1062), .ZN(n1061) );
XNOR2_X1 U761 ( .A(n1063), .B(G131), .ZN(n1062) );
NAND2_X1 U762 ( .A1(n1064), .A2(G953), .ZN(n1051) );
XOR2_X1 U763 ( .A(n1065), .B(KEYINPUT28), .Z(n1064) );
NAND2_X1 U764 ( .A1(G900), .A2(G227), .ZN(n1065) );
NOR2_X1 U765 ( .A1(n1066), .A2(G953), .ZN(n1049) );
XOR2_X1 U766 ( .A(n1067), .B(n1068), .Z(G69) );
XOR2_X1 U767 ( .A(n1069), .B(n1070), .Z(n1068) );
NOR2_X1 U768 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
AND2_X1 U769 ( .A1(G224), .A2(G898), .ZN(n1071) );
NAND2_X1 U770 ( .A1(n1073), .A2(n1074), .ZN(n1069) );
NAND2_X1 U771 ( .A1(G953), .A2(n1075), .ZN(n1074) );
XOR2_X1 U772 ( .A(n1076), .B(n1077), .Z(n1073) );
XNOR2_X1 U773 ( .A(n1078), .B(n1079), .ZN(n1077) );
NOR2_X1 U774 ( .A1(KEYINPUT59), .A2(n1080), .ZN(n1079) );
XNOR2_X1 U775 ( .A(KEYINPUT5), .B(KEYINPUT49), .ZN(n1076) );
NAND2_X1 U776 ( .A1(n1072), .A2(n1081), .ZN(n1067) );
NAND2_X1 U777 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U778 ( .A1(n1084), .A2(n1085), .ZN(G66) );
XOR2_X1 U779 ( .A(n1086), .B(n1087), .Z(n1085) );
XOR2_X1 U780 ( .A(KEYINPUT38), .B(n1088), .Z(n1087) );
NOR2_X1 U781 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR2_X1 U782 ( .A1(n1084), .A2(n1091), .ZN(G63) );
XOR2_X1 U783 ( .A(n1092), .B(n1093), .Z(n1091) );
AND2_X1 U784 ( .A1(G478), .A2(n1094), .ZN(n1092) );
NOR2_X1 U785 ( .A1(n1084), .A2(n1095), .ZN(G60) );
XOR2_X1 U786 ( .A(n1096), .B(n1097), .Z(n1095) );
XOR2_X1 U787 ( .A(KEYINPUT63), .B(n1098), .Z(n1097) );
AND2_X1 U788 ( .A1(G475), .A2(n1094), .ZN(n1098) );
XOR2_X1 U789 ( .A(G104), .B(n1099), .Z(G6) );
NOR3_X1 U790 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
XNOR2_X1 U791 ( .A(n1013), .B(KEYINPUT55), .ZN(n1101) );
NOR2_X1 U792 ( .A1(n1084), .A2(n1103), .ZN(G57) );
XOR2_X1 U793 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U794 ( .A(n1106), .B(n1107), .Z(n1104) );
AND2_X1 U795 ( .A1(G472), .A2(n1094), .ZN(n1107) );
NAND3_X1 U796 ( .A1(n1108), .A2(n1109), .A3(KEYINPUT31), .ZN(n1106) );
NAND2_X1 U797 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U798 ( .A(KEYINPUT16), .B(n1112), .Z(n1108) );
NOR2_X1 U799 ( .A1(n1110), .A2(n1111), .ZN(n1112) );
XNOR2_X1 U800 ( .A(n1113), .B(KEYINPUT17), .ZN(n1111) );
XNOR2_X1 U801 ( .A(KEYINPUT3), .B(n1114), .ZN(n1110) );
NOR2_X1 U802 ( .A1(n1084), .A2(n1115), .ZN(G54) );
XOR2_X1 U803 ( .A(n1116), .B(n1117), .Z(n1115) );
XNOR2_X1 U804 ( .A(n1118), .B(n1119), .ZN(n1116) );
NAND2_X1 U805 ( .A1(KEYINPUT21), .A2(n1120), .ZN(n1119) );
NAND2_X1 U806 ( .A1(KEYINPUT48), .A2(n1121), .ZN(n1118) );
NAND2_X1 U807 ( .A1(n1094), .A2(G469), .ZN(n1121) );
NOR2_X1 U808 ( .A1(n1084), .A2(n1122), .ZN(G51) );
XNOR2_X1 U809 ( .A(n1123), .B(n1124), .ZN(n1122) );
XOR2_X1 U810 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U811 ( .A1(n1127), .A2(n1090), .ZN(n1126) );
INV_X1 U812 ( .A(n1094), .ZN(n1090) );
NOR2_X1 U813 ( .A1(n1128), .A2(n1006), .ZN(n1094) );
AND3_X1 U814 ( .A1(n1082), .A2(n1129), .A3(n1066), .ZN(n1006) );
AND2_X1 U815 ( .A1(n1130), .A2(n1131), .ZN(n1066) );
NOR4_X1 U816 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1131) );
NOR2_X1 U817 ( .A1(n1100), .A2(n1136), .ZN(n1135) );
INV_X1 U818 ( .A(n1034), .ZN(n1100) );
AND4_X1 U819 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1130) );
NAND2_X1 U820 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XNOR2_X1 U821 ( .A(KEYINPUT26), .B(n1083), .ZN(n1129) );
AND4_X1 U822 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1082) );
NOR4_X1 U823 ( .A1(n1147), .A2(n1148), .A3(n997), .A4(n1149), .ZN(n1146) );
AND3_X1 U824 ( .A1(n1012), .A2(n1013), .A3(n1150), .ZN(n997) );
NAND3_X1 U825 ( .A1(n1150), .A2(n1013), .A3(n1034), .ZN(n1145) );
NAND2_X1 U826 ( .A1(n1151), .A2(n1152), .ZN(n1144) );
XNOR2_X1 U827 ( .A(n1004), .B(KEYINPUT20), .ZN(n1151) );
NAND2_X1 U828 ( .A1(n1153), .A2(n1154), .ZN(n1143) );
NOR2_X1 U829 ( .A1(KEYINPUT14), .A2(n1155), .ZN(n1125) );
NOR2_X1 U830 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U831 ( .A(KEYINPUT58), .B(n1158), .Z(n1157) );
NOR2_X1 U832 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U833 ( .A(n1060), .B(n1114), .ZN(n1160) );
NOR2_X1 U834 ( .A1(n1161), .A2(n1162), .ZN(n1156) );
XNOR2_X1 U835 ( .A(G125), .B(n1114), .ZN(n1162) );
INV_X1 U836 ( .A(n1159), .ZN(n1161) );
NOR2_X1 U837 ( .A1(n1072), .A2(G952), .ZN(n1084) );
XNOR2_X1 U838 ( .A(G146), .B(n1163), .ZN(G48) );
NAND4_X1 U839 ( .A1(KEYINPUT27), .A2(n1142), .A3(n1041), .A4(n1164), .ZN(n1163) );
XNOR2_X1 U840 ( .A(KEYINPUT36), .B(n1165), .ZN(n1164) );
AND3_X1 U841 ( .A1(n1166), .A2(n1167), .A3(n1034), .ZN(n1142) );
XNOR2_X1 U842 ( .A(G143), .B(n1139), .ZN(G45) );
NAND3_X1 U843 ( .A1(n1141), .A2(n1004), .A3(n1168), .ZN(n1139) );
NOR3_X1 U844 ( .A1(n1040), .A2(n1169), .A3(n1170), .ZN(n1168) );
XNOR2_X1 U845 ( .A(G140), .B(n1138), .ZN(G42) );
NAND4_X1 U846 ( .A1(n1141), .A2(n1034), .A3(n1017), .A4(n1019), .ZN(n1138) );
XNOR2_X1 U847 ( .A(G137), .B(n1137), .ZN(G39) );
NAND3_X1 U848 ( .A1(n1141), .A2(n1019), .A3(n1154), .ZN(n1137) );
XNOR2_X1 U849 ( .A(n1134), .B(n1171), .ZN(G36) );
NOR2_X1 U850 ( .A1(G134), .A2(KEYINPUT60), .ZN(n1171) );
NOR2_X1 U851 ( .A1(n1136), .A2(n1172), .ZN(n1134) );
INV_X1 U852 ( .A(n1012), .ZN(n1172) );
NAND3_X1 U853 ( .A1(n1004), .A2(n1019), .A3(n1141), .ZN(n1136) );
XNOR2_X1 U854 ( .A(G131), .B(n1173), .ZN(G33) );
NAND4_X1 U855 ( .A1(n1141), .A2(n1004), .A3(n1034), .A4(n1174), .ZN(n1173) );
XOR2_X1 U856 ( .A(KEYINPUT4), .B(n1019), .Z(n1174) );
NOR2_X1 U857 ( .A1(n1175), .A2(n1025), .ZN(n1019) );
XOR2_X1 U858 ( .A(G128), .B(n1133), .Z(G30) );
AND4_X1 U859 ( .A1(n1141), .A2(n1012), .A3(n1166), .A4(n1167), .ZN(n1133) );
AND2_X1 U860 ( .A1(n1041), .A2(n1165), .ZN(n1141) );
XNOR2_X1 U861 ( .A(G101), .B(n1176), .ZN(G3) );
NAND2_X1 U862 ( .A1(n1152), .A2(n1004), .ZN(n1176) );
XNOR2_X1 U863 ( .A(n1177), .B(n1060), .ZN(G27) );
NAND2_X1 U864 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND3_X1 U865 ( .A1(n1180), .A2(n1040), .A3(n1181), .ZN(n1179) );
INV_X1 U866 ( .A(KEYINPUT12), .ZN(n1181) );
INV_X1 U867 ( .A(n1166), .ZN(n1040) );
NAND2_X1 U868 ( .A1(n1132), .A2(KEYINPUT12), .ZN(n1178) );
AND2_X1 U869 ( .A1(n1180), .A2(n1166), .ZN(n1132) );
AND4_X1 U870 ( .A1(n1034), .A2(n1017), .A3(n1018), .A4(n1165), .ZN(n1180) );
NAND2_X1 U871 ( .A1(n1182), .A2(n1031), .ZN(n1165) );
NAND4_X1 U872 ( .A1(G953), .A2(G902), .A3(n1183), .A4(n1055), .ZN(n1182) );
INV_X1 U873 ( .A(G900), .ZN(n1055) );
XOR2_X1 U874 ( .A(G122), .B(n1148), .Z(G24) );
AND4_X1 U875 ( .A1(n1153), .A2(n1013), .A3(n1184), .A4(n1047), .ZN(n1148) );
NOR2_X1 U876 ( .A1(n1185), .A2(n1186), .ZN(n1013) );
XNOR2_X1 U877 ( .A(G119), .B(n1187), .ZN(G21) );
NAND4_X1 U878 ( .A1(n1188), .A2(n1154), .A3(n1166), .A4(n1189), .ZN(n1187) );
AND2_X1 U879 ( .A1(n1005), .A2(n1167), .ZN(n1154) );
NAND2_X1 U880 ( .A1(n1190), .A2(n1191), .ZN(n1167) );
NAND3_X1 U881 ( .A1(n1186), .A2(n1185), .A3(n1192), .ZN(n1191) );
INV_X1 U882 ( .A(KEYINPUT10), .ZN(n1192) );
NAND2_X1 U883 ( .A1(KEYINPUT10), .A2(n1004), .ZN(n1190) );
XNOR2_X1 U884 ( .A(n1018), .B(KEYINPUT42), .ZN(n1188) );
XNOR2_X1 U885 ( .A(G116), .B(n1193), .ZN(G18) );
NAND2_X1 U886 ( .A1(KEYINPUT45), .A2(n1147), .ZN(n1193) );
AND3_X1 U887 ( .A1(n1004), .A2(n1012), .A3(n1153), .ZN(n1147) );
NOR2_X1 U888 ( .A1(n1047), .A2(n1170), .ZN(n1012) );
INV_X1 U889 ( .A(n1184), .ZN(n1170) );
NAND2_X1 U890 ( .A1(n1194), .A2(n1195), .ZN(G15) );
NAND2_X1 U891 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND2_X1 U892 ( .A1(n1198), .A2(G113), .ZN(n1194) );
NAND2_X1 U893 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND2_X1 U894 ( .A1(KEYINPUT34), .A2(n1201), .ZN(n1200) );
INV_X1 U895 ( .A(n1083), .ZN(n1201) );
OR2_X1 U896 ( .A1(n1196), .A2(KEYINPUT34), .ZN(n1199) );
NOR2_X1 U897 ( .A1(KEYINPUT35), .A2(n1083), .ZN(n1196) );
NAND3_X1 U898 ( .A1(n1004), .A2(n1034), .A3(n1153), .ZN(n1083) );
AND3_X1 U899 ( .A1(n1166), .A2(n1189), .A3(n1018), .ZN(n1153) );
NOR2_X1 U900 ( .A1(n1202), .A2(n1028), .ZN(n1018) );
NOR2_X1 U901 ( .A1(n1184), .A2(n1169), .ZN(n1034) );
INV_X1 U902 ( .A(n1047), .ZN(n1169) );
NOR2_X1 U903 ( .A1(n1185), .A2(n1042), .ZN(n1004) );
NAND3_X1 U904 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(G12) );
NAND2_X1 U905 ( .A1(G110), .A2(n1206), .ZN(n1205) );
NAND2_X1 U906 ( .A1(n1207), .A2(n1208), .ZN(n1204) );
INV_X1 U907 ( .A(KEYINPUT1), .ZN(n1208) );
NAND2_X1 U908 ( .A1(n1209), .A2(n1149), .ZN(n1207) );
INV_X1 U909 ( .A(n1206), .ZN(n1149) );
XNOR2_X1 U910 ( .A(KEYINPUT53), .B(G110), .ZN(n1209) );
NAND2_X1 U911 ( .A1(KEYINPUT1), .A2(n1210), .ZN(n1203) );
NAND2_X1 U912 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
OR3_X1 U913 ( .A1(n1206), .A2(G110), .A3(KEYINPUT53), .ZN(n1212) );
NAND2_X1 U914 ( .A1(n1152), .A2(n1017), .ZN(n1206) );
AND2_X1 U915 ( .A1(n1042), .A2(n1185), .ZN(n1017) );
NAND3_X1 U916 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1185) );
XOR2_X1 U917 ( .A(KEYINPUT29), .B(n1044), .Z(n1215) );
AND2_X1 U918 ( .A1(n1216), .A2(n1089), .ZN(n1044) );
NAND2_X1 U919 ( .A1(n1045), .A2(n1217), .ZN(n1214) );
INV_X1 U920 ( .A(KEYINPUT9), .ZN(n1217) );
NOR2_X1 U921 ( .A1(n1089), .A2(n1216), .ZN(n1045) );
INV_X1 U922 ( .A(n1218), .ZN(n1216) );
NAND3_X1 U923 ( .A1(n1218), .A2(n1089), .A3(KEYINPUT9), .ZN(n1213) );
NAND2_X1 U924 ( .A1(G217), .A2(n1219), .ZN(n1089) );
NAND2_X1 U925 ( .A1(n1086), .A2(n1128), .ZN(n1218) );
XNOR2_X1 U926 ( .A(n1220), .B(n1221), .ZN(n1086) );
XOR2_X1 U927 ( .A(n1222), .B(n1223), .Z(n1221) );
NAND2_X1 U928 ( .A1(n1224), .A2(G221), .ZN(n1223) );
NAND2_X1 U929 ( .A1(KEYINPUT30), .A2(n1225), .ZN(n1222) );
XOR2_X1 U930 ( .A(n1226), .B(n1227), .Z(n1225) );
XOR2_X1 U931 ( .A(n1228), .B(n1229), .Z(n1227) );
XOR2_X1 U932 ( .A(G119), .B(G110), .Z(n1226) );
INV_X1 U933 ( .A(n1186), .ZN(n1042) );
XNOR2_X1 U934 ( .A(n1230), .B(G472), .ZN(n1186) );
NAND2_X1 U935 ( .A1(n1231), .A2(n1128), .ZN(n1230) );
XNOR2_X1 U936 ( .A(n1105), .B(n1232), .ZN(n1231) );
NOR2_X1 U937 ( .A1(KEYINPUT8), .A2(n1233), .ZN(n1232) );
XNOR2_X1 U938 ( .A(n1113), .B(n1114), .ZN(n1233) );
INV_X1 U939 ( .A(n1234), .ZN(n1113) );
XNOR2_X1 U940 ( .A(n1235), .B(n1236), .ZN(n1105) );
XNOR2_X1 U941 ( .A(n1237), .B(n1238), .ZN(n1236) );
NAND2_X1 U942 ( .A1(KEYINPUT54), .A2(G116), .ZN(n1237) );
XNOR2_X1 U943 ( .A(n1239), .B(n1197), .ZN(n1235) );
NAND3_X1 U944 ( .A1(n1240), .A2(n1072), .A3(n1241), .ZN(n1239) );
XOR2_X1 U945 ( .A(KEYINPUT23), .B(G210), .Z(n1241) );
AND2_X1 U946 ( .A1(n1005), .A2(n1150), .ZN(n1152) );
INV_X1 U947 ( .A(n1102), .ZN(n1150) );
NAND3_X1 U948 ( .A1(n1041), .A2(n1189), .A3(n1166), .ZN(n1102) );
NOR2_X1 U949 ( .A1(n1024), .A2(n1025), .ZN(n1166) );
AND2_X1 U950 ( .A1(G214), .A2(n1242), .ZN(n1025) );
INV_X1 U951 ( .A(n1175), .ZN(n1024) );
XOR2_X1 U952 ( .A(n1243), .B(n1127), .Z(n1175) );
NAND2_X1 U953 ( .A1(G210), .A2(n1242), .ZN(n1127) );
NAND2_X1 U954 ( .A1(n1128), .A2(n1240), .ZN(n1242) );
NAND2_X1 U955 ( .A1(n1244), .A2(n1128), .ZN(n1243) );
XOR2_X1 U956 ( .A(n1245), .B(n1246), .Z(n1244) );
NOR2_X1 U957 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NOR2_X1 U958 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
XNOR2_X1 U959 ( .A(KEYINPUT32), .B(n1159), .ZN(n1249) );
AND2_X1 U960 ( .A1(n1159), .A2(n1250), .ZN(n1247) );
NAND3_X1 U961 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1250) );
OR2_X1 U962 ( .A1(n1060), .A2(KEYINPUT18), .ZN(n1253) );
NAND3_X1 U963 ( .A1(KEYINPUT18), .A2(n1060), .A3(n1114), .ZN(n1252) );
NAND2_X1 U964 ( .A1(n1254), .A2(n1255), .ZN(n1251) );
NAND2_X1 U965 ( .A1(n1256), .A2(KEYINPUT18), .ZN(n1255) );
XNOR2_X1 U966 ( .A(n1257), .B(n1060), .ZN(n1256) );
INV_X1 U967 ( .A(G125), .ZN(n1060) );
XNOR2_X1 U968 ( .A(KEYINPUT6), .B(KEYINPUT11), .ZN(n1257) );
INV_X1 U969 ( .A(n1114), .ZN(n1254) );
XOR2_X1 U970 ( .A(G143), .B(n1228), .Z(n1114) );
XOR2_X1 U971 ( .A(G128), .B(G146), .Z(n1228) );
NAND2_X1 U972 ( .A1(G224), .A2(n1072), .ZN(n1159) );
NOR2_X1 U973 ( .A1(KEYINPUT57), .A2(n1123), .ZN(n1245) );
XOR2_X1 U974 ( .A(n1258), .B(n1259), .Z(n1123) );
INV_X1 U975 ( .A(n1078), .ZN(n1259) );
XOR2_X1 U976 ( .A(G110), .B(n1260), .Z(n1078) );
XOR2_X1 U977 ( .A(KEYINPUT37), .B(G122), .Z(n1260) );
NAND2_X1 U978 ( .A1(KEYINPUT47), .A2(n1261), .ZN(n1258) );
INV_X1 U979 ( .A(n1080), .ZN(n1261) );
XNOR2_X1 U980 ( .A(n1262), .B(n1263), .ZN(n1080) );
XOR2_X1 U981 ( .A(n1238), .B(n1264), .Z(n1263) );
XNOR2_X1 U982 ( .A(n1265), .B(G119), .ZN(n1238) );
XNOR2_X1 U983 ( .A(G116), .B(n1266), .ZN(n1262) );
NOR2_X1 U984 ( .A1(KEYINPUT15), .A2(n1197), .ZN(n1266) );
INV_X1 U985 ( .A(G113), .ZN(n1197) );
NAND2_X1 U986 ( .A1(n1031), .A2(n1267), .ZN(n1189) );
NAND4_X1 U987 ( .A1(G953), .A2(G902), .A3(n1183), .A4(n1075), .ZN(n1267) );
INV_X1 U988 ( .A(G898), .ZN(n1075) );
NAND3_X1 U989 ( .A1(n1183), .A2(n1072), .A3(n1268), .ZN(n1031) );
XOR2_X1 U990 ( .A(KEYINPUT52), .B(G952), .Z(n1268) );
NAND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1183) );
NOR2_X1 U992 ( .A1(n1029), .A2(n1028), .ZN(n1041) );
AND2_X1 U993 ( .A1(G221), .A2(n1219), .ZN(n1028) );
NAND2_X1 U994 ( .A1(G234), .A2(n1128), .ZN(n1219) );
INV_X1 U995 ( .A(n1202), .ZN(n1029) );
XNOR2_X1 U996 ( .A(n1269), .B(G469), .ZN(n1202) );
NAND2_X1 U997 ( .A1(n1270), .A2(n1128), .ZN(n1269) );
XNOR2_X1 U998 ( .A(n1117), .B(n1271), .ZN(n1270) );
XOR2_X1 U999 ( .A(n1272), .B(KEYINPUT62), .Z(n1271) );
NAND2_X1 U1000 ( .A1(KEYINPUT33), .A2(n1120), .ZN(n1272) );
XNOR2_X1 U1001 ( .A(n1273), .B(n1274), .ZN(n1117) );
XOR2_X1 U1002 ( .A(n1275), .B(n1276), .Z(n1274) );
XNOR2_X1 U1003 ( .A(G110), .B(n1277), .ZN(n1276) );
AND2_X1 U1004 ( .A1(n1072), .A2(G227), .ZN(n1277) );
NAND2_X1 U1005 ( .A1(KEYINPUT25), .A2(n1265), .ZN(n1275) );
INV_X1 U1006 ( .A(G101), .ZN(n1265) );
XOR2_X1 U1007 ( .A(n1278), .B(n1264), .Z(n1273) );
XOR2_X1 U1008 ( .A(G104), .B(G107), .Z(n1264) );
XNOR2_X1 U1009 ( .A(n1234), .B(n1059), .ZN(n1278) );
XNOR2_X1 U1010 ( .A(n1279), .B(n1280), .ZN(n1059) );
NOR2_X1 U1011 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XOR2_X1 U1012 ( .A(n1283), .B(KEYINPUT19), .Z(n1282) );
NAND2_X1 U1013 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NOR2_X1 U1014 ( .A1(n1286), .A2(n1285), .ZN(n1281) );
XOR2_X1 U1015 ( .A(n1284), .B(KEYINPUT43), .Z(n1286) );
XNOR2_X1 U1016 ( .A(G146), .B(KEYINPUT2), .ZN(n1284) );
NAND2_X1 U1017 ( .A1(KEYINPUT41), .A2(G128), .ZN(n1279) );
XOR2_X1 U1018 ( .A(n1287), .B(n1288), .Z(n1234) );
INV_X1 U1019 ( .A(n1063), .ZN(n1288) );
XOR2_X1 U1020 ( .A(G134), .B(n1220), .Z(n1063) );
XOR2_X1 U1021 ( .A(G137), .B(KEYINPUT61), .Z(n1220) );
NAND2_X1 U1022 ( .A1(KEYINPUT0), .A2(n1289), .ZN(n1287) );
INV_X1 U1023 ( .A(G131), .ZN(n1289) );
NOR2_X1 U1024 ( .A1(n1184), .A2(n1047), .ZN(n1005) );
XNOR2_X1 U1025 ( .A(n1290), .B(G475), .ZN(n1047) );
NAND2_X1 U1026 ( .A1(n1096), .A2(n1128), .ZN(n1290) );
INV_X1 U1027 ( .A(G902), .ZN(n1128) );
XOR2_X1 U1028 ( .A(n1291), .B(n1292), .Z(n1096) );
XOR2_X1 U1029 ( .A(n1229), .B(n1293), .Z(n1292) );
XOR2_X1 U1030 ( .A(G104), .B(n1294), .Z(n1293) );
NOR2_X1 U1031 ( .A1(KEYINPUT50), .A2(n1295), .ZN(n1294) );
XOR2_X1 U1032 ( .A(n1296), .B(n1297), .Z(n1295) );
XNOR2_X1 U1033 ( .A(G131), .B(G143), .ZN(n1297) );
NAND3_X1 U1034 ( .A1(n1240), .A2(n1072), .A3(n1298), .ZN(n1296) );
XOR2_X1 U1035 ( .A(KEYINPUT39), .B(G214), .Z(n1298) );
INV_X1 U1036 ( .A(G237), .ZN(n1240) );
XNOR2_X1 U1037 ( .A(n1120), .B(G125), .ZN(n1229) );
INV_X1 U1038 ( .A(G140), .ZN(n1120) );
XNOR2_X1 U1039 ( .A(G113), .B(n1299), .ZN(n1291) );
XOR2_X1 U1040 ( .A(G146), .B(G122), .Z(n1299) );
XNOR2_X1 U1041 ( .A(n1048), .B(KEYINPUT56), .ZN(n1184) );
XOR2_X1 U1042 ( .A(n1300), .B(G478), .Z(n1048) );
OR2_X1 U1043 ( .A1(n1093), .A2(G902), .ZN(n1300) );
XNOR2_X1 U1044 ( .A(n1301), .B(n1302), .ZN(n1093) );
XOR2_X1 U1045 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U1046 ( .A(G122), .B(G116), .Z(n1304) );
XNOR2_X1 U1047 ( .A(n1285), .B(G134), .ZN(n1303) );
INV_X1 U1048 ( .A(G143), .ZN(n1285) );
XOR2_X1 U1049 ( .A(n1305), .B(n1306), .Z(n1301) );
NOR2_X1 U1050 ( .A1(G128), .A2(KEYINPUT51), .ZN(n1306) );
XOR2_X1 U1051 ( .A(n1307), .B(G107), .Z(n1305) );
NAND2_X1 U1052 ( .A1(G217), .A2(n1224), .ZN(n1307) );
AND2_X1 U1053 ( .A1(G234), .A2(n1072), .ZN(n1224) );
INV_X1 U1054 ( .A(G953), .ZN(n1072) );
NAND2_X1 U1055 ( .A1(KEYINPUT53), .A2(G110), .ZN(n1211) );
endmodule


