//Key = 0001110100000110010010000101111000001111100111010101011011001010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282;

XNOR2_X1 U716 ( .A(G107), .B(n975), .ZN(G9) );
NOR2_X1 U717 ( .A1(n976), .A2(n977), .ZN(G75) );
NOR4_X1 U718 ( .A1(n978), .A2(n979), .A3(n980), .A4(n981), .ZN(n977) );
XOR2_X1 U719 ( .A(n982), .B(KEYINPUT56), .Z(n980) );
NAND3_X1 U720 ( .A1(n983), .A2(n984), .A3(KEYINPUT25), .ZN(n982) );
NAND2_X1 U721 ( .A1(n985), .A2(n986), .ZN(n983) );
NAND3_X1 U722 ( .A1(n987), .A2(n988), .A3(n989), .ZN(n986) );
NAND2_X1 U723 ( .A1(n990), .A2(n991), .ZN(n985) );
NAND2_X1 U724 ( .A1(n992), .A2(n993), .ZN(n991) );
NAND2_X1 U725 ( .A1(n988), .A2(n994), .ZN(n993) );
NAND2_X1 U726 ( .A1(n995), .A2(n996), .ZN(n994) );
NAND2_X1 U727 ( .A1(n997), .A2(n998), .ZN(n996) );
XNOR2_X1 U728 ( .A(n999), .B(KEYINPUT7), .ZN(n997) );
NAND2_X1 U729 ( .A1(n1000), .A2(n1001), .ZN(n995) );
NAND2_X1 U730 ( .A1(n989), .A2(n1002), .ZN(n992) );
NAND4_X1 U731 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n978) );
NAND4_X1 U732 ( .A1(n1007), .A2(n1008), .A3(KEYINPUT25), .A4(n1009), .ZN(n1004) );
NOR2_X1 U733 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND2_X1 U734 ( .A1(n1012), .A2(n1013), .ZN(n1008) );
NAND2_X1 U735 ( .A1(n989), .A2(n988), .ZN(n1013) );
NAND3_X1 U736 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1007) );
NAND3_X1 U737 ( .A1(n1017), .A2(n1018), .A3(n989), .ZN(n1015) );
AND2_X1 U738 ( .A1(n1000), .A2(n999), .ZN(n989) );
NAND2_X1 U739 ( .A1(n988), .A2(n1019), .ZN(n1014) );
NAND2_X1 U740 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND3_X1 U741 ( .A1(n1000), .A2(n1022), .A3(n1023), .ZN(n1021) );
NAND2_X1 U742 ( .A1(n1024), .A2(n1025), .ZN(n1020) );
XNOR2_X1 U743 ( .A(n999), .B(KEYINPUT40), .ZN(n1024) );
XNOR2_X1 U744 ( .A(KEYINPUT19), .B(n1026), .ZN(n1003) );
NOR3_X1 U745 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n976) );
XOR2_X1 U746 ( .A(n981), .B(KEYINPUT54), .Z(n1029) );
INV_X1 U747 ( .A(G952), .ZN(n981) );
INV_X1 U748 ( .A(n1005), .ZN(n1028) );
NAND4_X1 U749 ( .A1(n999), .A2(n988), .A3(n1030), .A4(n1031), .ZN(n1005) );
NOR3_X1 U750 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
XNOR2_X1 U751 ( .A(n1035), .B(n1036), .ZN(n1034) );
NAND2_X1 U752 ( .A1(n1037), .A2(KEYINPUT57), .ZN(n1035) );
XOR2_X1 U753 ( .A(n1038), .B(KEYINPUT48), .Z(n1037) );
XNOR2_X1 U754 ( .A(n1039), .B(n1040), .ZN(n1033) );
XNOR2_X1 U755 ( .A(KEYINPUT41), .B(n1041), .ZN(n1039) );
NOR2_X1 U756 ( .A1(KEYINPUT55), .A2(n1042), .ZN(n1041) );
XNOR2_X1 U757 ( .A(n1043), .B(G475), .ZN(n1030) );
XOR2_X1 U758 ( .A(KEYINPUT42), .B(G953), .Z(n1027) );
XOR2_X1 U759 ( .A(n1044), .B(n1045), .Z(G72) );
NOR2_X1 U760 ( .A1(KEYINPUT59), .A2(n1046), .ZN(n1045) );
XOR2_X1 U761 ( .A(n1047), .B(n1048), .Z(n1046) );
AND2_X1 U762 ( .A1(n1026), .A2(n1006), .ZN(n1048) );
NAND2_X1 U763 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
XOR2_X1 U764 ( .A(n1051), .B(n1052), .Z(n1049) );
XOR2_X1 U765 ( .A(n1053), .B(KEYINPUT46), .Z(n1052) );
NAND2_X1 U766 ( .A1(KEYINPUT30), .A2(n1054), .ZN(n1053) );
NOR2_X1 U767 ( .A1(n1006), .A2(n1055), .ZN(n1044) );
XOR2_X1 U768 ( .A(KEYINPUT0), .B(n1056), .Z(n1055) );
NOR2_X1 U769 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
XOR2_X1 U770 ( .A(n1059), .B(n1060), .Z(G69) );
XOR2_X1 U771 ( .A(n1061), .B(n1062), .Z(n1060) );
NOR2_X1 U772 ( .A1(G953), .A2(n1063), .ZN(n1062) );
XNOR2_X1 U773 ( .A(KEYINPUT52), .B(n979), .ZN(n1063) );
NAND3_X1 U774 ( .A1(KEYINPUT4), .A2(n1064), .A3(n1065), .ZN(n1061) );
XOR2_X1 U775 ( .A(n1066), .B(n1067), .Z(n1065) );
XOR2_X1 U776 ( .A(n1068), .B(n1069), .Z(n1067) );
XOR2_X1 U777 ( .A(n1070), .B(n1071), .Z(n1066) );
NAND2_X1 U778 ( .A1(n1072), .A2(n1073), .ZN(n1064) );
XNOR2_X1 U779 ( .A(KEYINPUT49), .B(n1074), .ZN(n1072) );
NAND2_X1 U780 ( .A1(G953), .A2(n1075), .ZN(n1059) );
NAND2_X1 U781 ( .A1(G224), .A2(G898), .ZN(n1075) );
NOR2_X1 U782 ( .A1(n1076), .A2(n1077), .ZN(G66) );
NOR3_X1 U783 ( .A1(n1042), .A2(n1078), .A3(n1079), .ZN(n1077) );
NOR4_X1 U784 ( .A1(n1080), .A2(n1081), .A3(KEYINPUT15), .A4(n1040), .ZN(n1079) );
INV_X1 U785 ( .A(n1082), .ZN(n1080) );
NOR2_X1 U786 ( .A1(n1083), .A2(n1082), .ZN(n1078) );
NOR3_X1 U787 ( .A1(n1040), .A2(KEYINPUT15), .A3(n1084), .ZN(n1083) );
NOR2_X1 U788 ( .A1(n1076), .A2(n1085), .ZN(G63) );
XNOR2_X1 U789 ( .A(n1086), .B(n1087), .ZN(n1085) );
NAND3_X1 U790 ( .A1(n1088), .A2(n1089), .A3(G478), .ZN(n1086) );
XOR2_X1 U791 ( .A(KEYINPUT12), .B(G902), .Z(n1088) );
NOR2_X1 U792 ( .A1(n1076), .A2(n1090), .ZN(G60) );
NOR3_X1 U793 ( .A1(n1043), .A2(n1091), .A3(n1092), .ZN(n1090) );
AND3_X1 U794 ( .A1(n1093), .A2(G475), .A3(n1094), .ZN(n1092) );
NOR2_X1 U795 ( .A1(n1095), .A2(n1093), .ZN(n1091) );
AND2_X1 U796 ( .A1(n1089), .A2(G475), .ZN(n1095) );
NAND2_X1 U797 ( .A1(n1096), .A2(n1097), .ZN(G6) );
NAND2_X1 U798 ( .A1(G104), .A2(n1098), .ZN(n1097) );
XOR2_X1 U799 ( .A(n1099), .B(KEYINPUT31), .Z(n1096) );
OR2_X1 U800 ( .A1(n1098), .A2(G104), .ZN(n1099) );
NOR2_X1 U801 ( .A1(n1076), .A2(n1100), .ZN(G57) );
XOR2_X1 U802 ( .A(n1101), .B(n1102), .Z(n1100) );
XOR2_X1 U803 ( .A(n1103), .B(n1104), .Z(n1102) );
INV_X1 U804 ( .A(n1105), .ZN(n1103) );
XOR2_X1 U805 ( .A(n1106), .B(n1107), .Z(n1101) );
XOR2_X1 U806 ( .A(KEYINPUT60), .B(n1108), .Z(n1107) );
NOR2_X1 U807 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U808 ( .A(KEYINPUT44), .B(KEYINPUT37), .Z(n1110) );
NOR2_X1 U809 ( .A1(n1038), .A2(n1081), .ZN(n1106) );
INV_X1 U810 ( .A(G472), .ZN(n1038) );
NOR2_X1 U811 ( .A1(n1076), .A2(n1111), .ZN(G54) );
XOR2_X1 U812 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U813 ( .A(n1105), .B(n1114), .Z(n1113) );
NAND2_X1 U814 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U815 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U816 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NAND2_X1 U817 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U818 ( .A1(n1123), .A2(n1124), .ZN(n1119) );
NAND2_X1 U819 ( .A1(G110), .A2(n1125), .ZN(n1115) );
NAND2_X1 U820 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U821 ( .A1(n1121), .A2(n1124), .ZN(n1127) );
INV_X1 U822 ( .A(n1122), .ZN(n1124) );
NAND2_X1 U823 ( .A1(n1122), .A2(n1123), .ZN(n1126) );
XOR2_X1 U824 ( .A(n1128), .B(n1121), .Z(n1123) );
XNOR2_X1 U825 ( .A(KEYINPUT29), .B(KEYINPUT14), .ZN(n1128) );
NOR2_X1 U826 ( .A1(G140), .A2(KEYINPUT21), .ZN(n1122) );
XOR2_X1 U827 ( .A(n1129), .B(n1130), .Z(n1112) );
AND2_X1 U828 ( .A1(G469), .A2(n1094), .ZN(n1130) );
NAND3_X1 U829 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1129) );
NAND2_X1 U830 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
OR3_X1 U831 ( .A1(n1135), .A2(n1134), .A3(KEYINPUT9), .ZN(n1132) );
NAND2_X1 U832 ( .A1(KEYINPUT51), .A2(n1136), .ZN(n1135) );
NAND2_X1 U833 ( .A1(KEYINPUT9), .A2(n1137), .ZN(n1131) );
INV_X1 U834 ( .A(n1136), .ZN(n1137) );
XOR2_X1 U835 ( .A(KEYINPUT32), .B(n1109), .Z(n1136) );
NOR2_X1 U836 ( .A1(n1076), .A2(n1138), .ZN(G51) );
XOR2_X1 U837 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U838 ( .A1(KEYINPUT63), .A2(n1141), .ZN(n1140) );
XNOR2_X1 U839 ( .A(n1142), .B(KEYINPUT61), .ZN(n1141) );
NAND2_X1 U840 ( .A1(n1094), .A2(G210), .ZN(n1139) );
INV_X1 U841 ( .A(n1081), .ZN(n1094) );
NAND2_X1 U842 ( .A1(G902), .A2(n1089), .ZN(n1081) );
INV_X1 U843 ( .A(n1084), .ZN(n1089) );
NOR2_X1 U844 ( .A1(n979), .A2(n1026), .ZN(n1084) );
NAND4_X1 U845 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1026) );
NOR4_X1 U846 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1146) );
INV_X1 U847 ( .A(n1151), .ZN(n1149) );
NOR2_X1 U848 ( .A1(n1152), .A2(n1153), .ZN(n1145) );
NAND2_X1 U849 ( .A1(n1154), .A2(n999), .ZN(n1143) );
XOR2_X1 U850 ( .A(KEYINPUT47), .B(n1155), .Z(n1154) );
NOR2_X1 U851 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NOR2_X1 U852 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
AND4_X1 U853 ( .A1(n1158), .A2(n1160), .A3(n1161), .A4(n1000), .ZN(n1156) );
INV_X1 U854 ( .A(KEYINPUT38), .ZN(n1158) );
NAND2_X1 U855 ( .A1(n1162), .A2(n1163), .ZN(n979) );
AND4_X1 U856 ( .A1(n1164), .A2(n975), .A3(n1165), .A4(n1166), .ZN(n1163) );
NAND3_X1 U857 ( .A1(n990), .A2(n1167), .A3(n1025), .ZN(n975) );
AND4_X1 U858 ( .A1(n1168), .A2(n1169), .A3(n1098), .A4(n1170), .ZN(n1162) );
NAND3_X1 U859 ( .A1(n987), .A2(n1167), .A3(n1000), .ZN(n1170) );
NAND3_X1 U860 ( .A1(n990), .A2(n1167), .A3(n998), .ZN(n1098) );
NOR2_X1 U861 ( .A1(n1006), .A2(G952), .ZN(n1076) );
XOR2_X1 U862 ( .A(n1171), .B(n1144), .Z(G48) );
NAND4_X1 U863 ( .A1(n1160), .A2(n998), .A3(n1001), .A4(n1002), .ZN(n1144) );
XOR2_X1 U864 ( .A(G143), .B(n1153), .Z(G45) );
AND4_X1 U865 ( .A1(n1001), .A2(n1172), .A3(n987), .A4(n1173), .ZN(n1153) );
NOR3_X1 U866 ( .A1(n1161), .A2(n1174), .A3(n1175), .ZN(n1173) );
XOR2_X1 U867 ( .A(G140), .B(n1152), .Z(G42) );
AND3_X1 U868 ( .A1(n999), .A2(n1002), .A3(n1176), .ZN(n1152) );
XNOR2_X1 U869 ( .A(G137), .B(n1177), .ZN(G39) );
NAND2_X1 U870 ( .A1(n1178), .A2(n999), .ZN(n1177) );
XOR2_X1 U871 ( .A(n1159), .B(KEYINPUT53), .Z(n1178) );
NAND3_X1 U872 ( .A1(n1000), .A2(n1002), .A3(n1160), .ZN(n1159) );
XOR2_X1 U873 ( .A(G134), .B(n1148), .Z(G36) );
AND2_X1 U874 ( .A1(n1179), .A2(n1025), .ZN(n1148) );
XOR2_X1 U875 ( .A(G131), .B(n1147), .Z(G33) );
AND2_X1 U876 ( .A1(n1179), .A2(n998), .ZN(n1147) );
AND4_X1 U877 ( .A1(n987), .A2(n999), .A3(n1002), .A4(n1180), .ZN(n1179) );
NOR2_X1 U878 ( .A1(n1181), .A2(n1023), .ZN(n999) );
XOR2_X1 U879 ( .A(n1150), .B(n1182), .Z(G30) );
NOR2_X1 U880 ( .A1(KEYINPUT6), .A2(n1183), .ZN(n1182) );
INV_X1 U881 ( .A(G128), .ZN(n1183) );
AND4_X1 U882 ( .A1(n1001), .A2(n1160), .A3(n1184), .A4(n1025), .ZN(n1150) );
NOR3_X1 U883 ( .A1(n1185), .A2(n1174), .A3(n1016), .ZN(n1160) );
INV_X1 U884 ( .A(n1180), .ZN(n1174) );
XNOR2_X1 U885 ( .A(G101), .B(n1186), .ZN(G3) );
NAND3_X1 U886 ( .A1(n1167), .A2(n1187), .A3(n1000), .ZN(n1186) );
XOR2_X1 U887 ( .A(KEYINPUT1), .B(n987), .Z(n1187) );
XOR2_X1 U888 ( .A(n1188), .B(n1151), .Z(G27) );
NAND3_X1 U889 ( .A1(n1001), .A2(n988), .A3(n1176), .ZN(n1151) );
AND4_X1 U890 ( .A1(n1185), .A2(n998), .A3(n1012), .A4(n1180), .ZN(n1176) );
NAND2_X1 U891 ( .A1(n1189), .A2(n1190), .ZN(n1180) );
OR3_X1 U892 ( .A1(n1191), .A2(n1010), .A3(n1050), .ZN(n1190) );
NAND2_X1 U893 ( .A1(n1073), .A2(n1058), .ZN(n1050) );
INV_X1 U894 ( .A(G900), .ZN(n1058) );
INV_X1 U895 ( .A(n984), .ZN(n1010) );
XNOR2_X1 U896 ( .A(G122), .B(n1164), .ZN(G24) );
NAND4_X1 U897 ( .A1(n1001), .A2(n988), .A3(n1172), .A4(n1192), .ZN(n1164) );
AND3_X1 U898 ( .A1(n990), .A2(n1193), .A3(n1032), .ZN(n1192) );
NOR2_X1 U899 ( .A1(n1011), .A2(n1012), .ZN(n990) );
XNOR2_X1 U900 ( .A(G119), .B(n1169), .ZN(G21) );
NAND4_X1 U901 ( .A1(n1001), .A2(n988), .A3(n1000), .A4(n1194), .ZN(n1169) );
AND3_X1 U902 ( .A1(n1012), .A2(n1193), .A3(n1011), .ZN(n1194) );
INV_X1 U903 ( .A(n1185), .ZN(n1011) );
XOR2_X1 U904 ( .A(n1195), .B(n1168), .Z(G18) );
NAND3_X1 U905 ( .A1(n1001), .A2(n1025), .A3(n1196), .ZN(n1168) );
NOR2_X1 U906 ( .A1(n1172), .A2(n1175), .ZN(n1025) );
XNOR2_X1 U907 ( .A(n1197), .B(KEYINPUT39), .ZN(n1001) );
XOR2_X1 U908 ( .A(G113), .B(n1198), .Z(G15) );
NOR2_X1 U909 ( .A1(KEYINPUT10), .A2(n1166), .ZN(n1198) );
NAND3_X1 U910 ( .A1(n1196), .A2(n1197), .A3(n998), .ZN(n1166) );
AND2_X1 U911 ( .A1(n1172), .A2(n1175), .ZN(n998) );
AND3_X1 U912 ( .A1(n988), .A2(n1193), .A3(n987), .ZN(n1196) );
NOR2_X1 U913 ( .A1(n1012), .A2(n1185), .ZN(n987) );
NOR2_X1 U914 ( .A1(n1199), .A2(n1018), .ZN(n988) );
INV_X1 U915 ( .A(n1017), .ZN(n1199) );
XOR2_X1 U916 ( .A(n1118), .B(n1165), .Z(G12) );
NAND4_X1 U917 ( .A1(n1000), .A2(n1167), .A3(n1185), .A4(n1012), .ZN(n1165) );
INV_X1 U918 ( .A(n1016), .ZN(n1012) );
XOR2_X1 U919 ( .A(n1042), .B(n1040), .Z(n1016) );
NAND2_X1 U920 ( .A1(G217), .A2(n1200), .ZN(n1040) );
NOR2_X1 U921 ( .A1(n1082), .A2(G902), .ZN(n1042) );
XOR2_X1 U922 ( .A(n1201), .B(n1202), .Z(n1082) );
XOR2_X1 U923 ( .A(n1203), .B(n1204), .Z(n1202) );
XOR2_X1 U924 ( .A(G110), .B(n1205), .Z(n1204) );
NOR2_X1 U925 ( .A1(KEYINPUT22), .A2(n1206), .ZN(n1205) );
XOR2_X1 U926 ( .A(G146), .B(n1054), .Z(n1206) );
XOR2_X1 U927 ( .A(n1188), .B(G140), .Z(n1054) );
INV_X1 U928 ( .A(G125), .ZN(n1188) );
AND3_X1 U929 ( .A1(G221), .A2(n1006), .A3(G234), .ZN(n1203) );
XNOR2_X1 U930 ( .A(G119), .B(n1207), .ZN(n1201) );
XOR2_X1 U931 ( .A(G137), .B(G128), .Z(n1207) );
XOR2_X1 U932 ( .A(n1036), .B(G472), .Z(n1185) );
NAND2_X1 U933 ( .A1(n1208), .A2(n1191), .ZN(n1036) );
XOR2_X1 U934 ( .A(n1209), .B(n1104), .Z(n1208) );
XNOR2_X1 U935 ( .A(n1070), .B(n1210), .ZN(n1104) );
XOR2_X1 U936 ( .A(n1211), .B(n1212), .Z(n1210) );
NAND2_X1 U937 ( .A1(KEYINPUT5), .A2(n1195), .ZN(n1212) );
INV_X1 U938 ( .A(G116), .ZN(n1195) );
NAND2_X1 U939 ( .A1(G210), .A2(n1213), .ZN(n1211) );
XNOR2_X1 U940 ( .A(G101), .B(n1214), .ZN(n1070) );
XNOR2_X1 U941 ( .A(n1109), .B(n1215), .ZN(n1209) );
NOR2_X1 U942 ( .A1(KEYINPUT35), .A2(n1105), .ZN(n1215) );
AND3_X1 U943 ( .A1(n1184), .A2(n1193), .A3(n1197), .ZN(n1167) );
NOR2_X1 U944 ( .A1(n1022), .A2(n1023), .ZN(n1197) );
AND2_X1 U945 ( .A1(G214), .A2(n1216), .ZN(n1023) );
OR2_X1 U946 ( .A1(G902), .A2(G237), .ZN(n1216) );
INV_X1 U947 ( .A(n1181), .ZN(n1022) );
NAND3_X1 U948 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1181) );
OR2_X1 U949 ( .A1(n1220), .A2(n1142), .ZN(n1219) );
NAND3_X1 U950 ( .A1(n1142), .A2(n1220), .A3(n1191), .ZN(n1218) );
NAND2_X1 U951 ( .A1(G237), .A2(G210), .ZN(n1220) );
XNOR2_X1 U952 ( .A(n1221), .B(n1222), .ZN(n1142) );
XOR2_X1 U953 ( .A(n1223), .B(n1109), .Z(n1222) );
AND2_X1 U954 ( .A1(n1006), .A2(G224), .ZN(n1223) );
XOR2_X1 U955 ( .A(n1224), .B(n1225), .Z(n1221) );
XOR2_X1 U956 ( .A(G125), .B(n1069), .Z(n1225) );
AND2_X1 U957 ( .A1(n1226), .A2(n1227), .ZN(n1069) );
NAND2_X1 U958 ( .A1(G122), .A2(n1228), .ZN(n1227) );
XOR2_X1 U959 ( .A(KEYINPUT13), .B(n1229), .Z(n1228) );
XOR2_X1 U960 ( .A(KEYINPUT43), .B(n1230), .Z(n1226) );
NOR2_X1 U961 ( .A1(G122), .A2(n1231), .ZN(n1230) );
XNOR2_X1 U962 ( .A(n1229), .B(KEYINPUT50), .ZN(n1231) );
XNOR2_X1 U963 ( .A(n1118), .B(KEYINPUT23), .ZN(n1229) );
NAND2_X1 U964 ( .A1(n1232), .A2(KEYINPUT45), .ZN(n1224) );
XOR2_X1 U965 ( .A(n1233), .B(n1234), .Z(n1232) );
XOR2_X1 U966 ( .A(n1071), .B(n1214), .Z(n1234) );
XOR2_X1 U967 ( .A(G113), .B(G119), .Z(n1214) );
XNOR2_X1 U968 ( .A(n1235), .B(G116), .ZN(n1071) );
XNOR2_X1 U969 ( .A(KEYINPUT20), .B(KEYINPUT18), .ZN(n1235) );
XNOR2_X1 U970 ( .A(KEYINPUT28), .B(n1236), .ZN(n1233) );
NOR2_X1 U971 ( .A1(KEYINPUT26), .A2(n1237), .ZN(n1236) );
XNOR2_X1 U972 ( .A(G101), .B(n1068), .ZN(n1237) );
NOR2_X1 U973 ( .A1(KEYINPUT16), .A2(n1238), .ZN(n1068) );
NAND2_X1 U974 ( .A1(G902), .A2(G210), .ZN(n1217) );
NAND2_X1 U975 ( .A1(n1189), .A2(n1239), .ZN(n1193) );
NAND4_X1 U976 ( .A1(n1074), .A2(n1240), .A3(n1073), .A4(n984), .ZN(n1239) );
XOR2_X1 U977 ( .A(G953), .B(KEYINPUT8), .Z(n1073) );
XOR2_X1 U978 ( .A(KEYINPUT2), .B(G902), .Z(n1240) );
XNOR2_X1 U979 ( .A(G898), .B(KEYINPUT34), .ZN(n1074) );
NAND3_X1 U980 ( .A1(n984), .A2(n1006), .A3(G952), .ZN(n1189) );
NAND2_X1 U981 ( .A1(G237), .A2(G234), .ZN(n984) );
XOR2_X1 U982 ( .A(n1161), .B(KEYINPUT62), .Z(n1184) );
INV_X1 U983 ( .A(n1002), .ZN(n1161) );
NOR2_X1 U984 ( .A1(n1017), .A2(n1018), .ZN(n1002) );
AND2_X1 U985 ( .A1(G221), .A2(n1200), .ZN(n1018) );
NAND2_X1 U986 ( .A1(G234), .A2(n1191), .ZN(n1200) );
XOR2_X1 U987 ( .A(n1241), .B(G469), .Z(n1017) );
NAND2_X1 U988 ( .A1(n1242), .A2(n1191), .ZN(n1241) );
INV_X1 U989 ( .A(G902), .ZN(n1191) );
XOR2_X1 U990 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U991 ( .A(n1051), .B(n1245), .Z(n1244) );
XNOR2_X1 U992 ( .A(n1134), .B(n1121), .ZN(n1245) );
NOR2_X1 U993 ( .A1(n1057), .A2(G953), .ZN(n1121) );
INV_X1 U994 ( .A(G227), .ZN(n1057) );
XNOR2_X1 U995 ( .A(G101), .B(n1238), .ZN(n1134) );
XOR2_X1 U996 ( .A(G107), .B(n1246), .Z(n1238) );
XOR2_X1 U997 ( .A(n1105), .B(n1109), .Z(n1051) );
XNOR2_X1 U998 ( .A(n1171), .B(n1247), .ZN(n1109) );
INV_X1 U999 ( .A(G146), .ZN(n1171) );
XOR2_X1 U1000 ( .A(n1248), .B(n1249), .Z(n1105) );
XOR2_X1 U1001 ( .A(G137), .B(G134), .Z(n1249) );
XOR2_X1 U1002 ( .A(G110), .B(n1250), .Z(n1243) );
XOR2_X1 U1003 ( .A(KEYINPUT32), .B(G140), .Z(n1250) );
NOR2_X1 U1004 ( .A1(n1032), .A2(n1172), .ZN(n1000) );
XNOR2_X1 U1005 ( .A(n1043), .B(n1251), .ZN(n1172) );
NOR2_X1 U1006 ( .A1(G475), .A2(KEYINPUT58), .ZN(n1251) );
NOR2_X1 U1007 ( .A1(n1093), .A2(G902), .ZN(n1043) );
XOR2_X1 U1008 ( .A(n1252), .B(n1253), .Z(n1093) );
XOR2_X1 U1009 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U1010 ( .A(G125), .B(G122), .Z(n1255) );
XOR2_X1 U1011 ( .A(KEYINPUT36), .B(G146), .Z(n1254) );
XOR2_X1 U1012 ( .A(n1256), .B(n1257), .Z(n1252) );
XNOR2_X1 U1013 ( .A(n1258), .B(n1259), .ZN(n1257) );
NOR2_X1 U1014 ( .A1(G140), .A2(KEYINPUT24), .ZN(n1259) );
NAND2_X1 U1015 ( .A1(KEYINPUT3), .A2(n1246), .ZN(n1258) );
INV_X1 U1016 ( .A(G104), .ZN(n1246) );
XOR2_X1 U1017 ( .A(n1260), .B(G113), .Z(n1256) );
NAND3_X1 U1018 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1260) );
OR2_X1 U1019 ( .A1(n1248), .A2(n1264), .ZN(n1263) );
NAND2_X1 U1020 ( .A1(KEYINPUT33), .A2(n1265), .ZN(n1262) );
NAND2_X1 U1021 ( .A1(n1266), .A2(n1264), .ZN(n1265) );
XOR2_X1 U1022 ( .A(KEYINPUT27), .B(G131), .Z(n1266) );
NAND2_X1 U1023 ( .A1(n1267), .A2(n1268), .ZN(n1261) );
INV_X1 U1024 ( .A(KEYINPUT33), .ZN(n1268) );
NAND2_X1 U1025 ( .A1(n1269), .A2(n1270), .ZN(n1267) );
NAND3_X1 U1026 ( .A1(KEYINPUT27), .A2(n1264), .A3(n1248), .ZN(n1270) );
XNOR2_X1 U1027 ( .A(n1271), .B(G143), .ZN(n1264) );
NAND2_X1 U1028 ( .A1(G214), .A2(n1213), .ZN(n1271) );
NOR2_X1 U1029 ( .A1(G953), .A2(G237), .ZN(n1213) );
OR2_X1 U1030 ( .A1(n1248), .A2(KEYINPUT27), .ZN(n1269) );
INV_X1 U1031 ( .A(G131), .ZN(n1248) );
INV_X1 U1032 ( .A(n1175), .ZN(n1032) );
XNOR2_X1 U1033 ( .A(G478), .B(n1272), .ZN(n1175) );
NOR2_X1 U1034 ( .A1(G902), .A2(n1087), .ZN(n1272) );
NAND3_X1 U1035 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1087) );
NAND2_X1 U1036 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
OR3_X1 U1037 ( .A1(n1277), .A2(n1276), .A3(KEYINPUT11), .ZN(n1274) );
XOR2_X1 U1038 ( .A(n1278), .B(n1279), .Z(n1276) );
XOR2_X1 U1039 ( .A(G116), .B(n1280), .Z(n1279) );
XOR2_X1 U1040 ( .A(G134), .B(G122), .Z(n1280) );
XNOR2_X1 U1041 ( .A(G107), .B(n1247), .ZN(n1278) );
XOR2_X1 U1042 ( .A(G128), .B(G143), .Z(n1247) );
NAND2_X1 U1043 ( .A1(KEYINPUT17), .A2(n1281), .ZN(n1277) );
INV_X1 U1044 ( .A(n1282), .ZN(n1281) );
NAND2_X1 U1045 ( .A1(KEYINPUT11), .A2(n1282), .ZN(n1273) );
NAND3_X1 U1046 ( .A1(G217), .A2(n1006), .A3(G234), .ZN(n1282) );
INV_X1 U1047 ( .A(G953), .ZN(n1006) );
INV_X1 U1048 ( .A(G110), .ZN(n1118) );
endmodule


