//Key = 1000100100001011111110010011011111101011001010101010011101111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357;

XNOR2_X1 U748 ( .A(n1032), .B(n1033), .ZN(G9) );
NOR2_X1 U749 ( .A1(n1034), .A2(n1035), .ZN(G75) );
NOR3_X1 U750 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NAND3_X1 U751 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1036) );
NAND2_X1 U752 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND4_X1 U754 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1045) );
NAND3_X1 U755 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1048) );
NAND2_X1 U756 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U758 ( .A1(n1057), .A2(n1058), .ZN(n1051) );
NAND2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U760 ( .A1(KEYINPUT54), .A2(n1061), .ZN(n1060) );
NAND2_X1 U761 ( .A1(KEYINPUT26), .A2(n1062), .ZN(n1059) );
NAND2_X1 U762 ( .A1(n1063), .A2(n1064), .ZN(n1050) );
NAND2_X1 U763 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
OR2_X1 U764 ( .A1(n1067), .A2(KEYINPUT54), .ZN(n1066) );
NAND2_X1 U765 ( .A1(n1062), .A2(n1068), .ZN(n1065) );
INV_X1 U766 ( .A(KEYINPUT26), .ZN(n1068) );
NAND3_X1 U767 ( .A1(n1053), .A2(n1069), .A3(n1057), .ZN(n1044) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND3_X1 U769 ( .A1(n1072), .A2(n1073), .A3(n1046), .ZN(n1071) );
NAND2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND3_X1 U771 ( .A1(n1076), .A2(n1077), .A3(n1049), .ZN(n1072) );
NAND2_X1 U772 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NAND2_X1 U773 ( .A1(n1047), .A2(n1080), .ZN(n1070) );
INV_X1 U774 ( .A(n1081), .ZN(n1042) );
NOR3_X1 U775 ( .A1(n1082), .A2(G953), .A3(n1083), .ZN(n1034) );
INV_X1 U776 ( .A(n1039), .ZN(n1083) );
NAND4_X1 U777 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1039) );
NOR4_X1 U778 ( .A1(n1088), .A2(n1074), .A3(n1089), .A4(n1090), .ZN(n1087) );
XNOR2_X1 U779 ( .A(n1091), .B(n1092), .ZN(n1090) );
NAND2_X1 U780 ( .A1(KEYINPUT29), .A2(n1093), .ZN(n1091) );
NOR2_X1 U781 ( .A1(n1094), .A2(n1095), .ZN(n1089) );
INV_X1 U782 ( .A(n1096), .ZN(n1088) );
NOR2_X1 U783 ( .A1(n1075), .A2(n1097), .ZN(n1086) );
XOR2_X1 U784 ( .A(n1098), .B(n1099), .Z(n1097) );
XNOR2_X1 U785 ( .A(KEYINPUT57), .B(KEYINPUT48), .ZN(n1099) );
XNOR2_X1 U786 ( .A(n1100), .B(n1101), .ZN(n1085) );
XOR2_X1 U787 ( .A(KEYINPUT30), .B(n1102), .Z(n1101) );
XNOR2_X1 U788 ( .A(KEYINPUT41), .B(n1037), .ZN(n1082) );
XOR2_X1 U789 ( .A(n1103), .B(n1104), .Z(G72) );
XOR2_X1 U790 ( .A(n1105), .B(n1106), .Z(n1104) );
NAND2_X1 U791 ( .A1(n1040), .A2(n1107), .ZN(n1106) );
NAND4_X1 U792 ( .A1(KEYINPUT7), .A2(n1108), .A3(n1109), .A4(n1110), .ZN(n1105) );
NAND2_X1 U793 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U794 ( .A1(G953), .A2(n1113), .ZN(n1109) );
XOR2_X1 U795 ( .A(KEYINPUT17), .B(n1114), .Z(n1108) );
NOR2_X1 U796 ( .A1(n1111), .A2(n1112), .ZN(n1114) );
XNOR2_X1 U797 ( .A(n1115), .B(n1116), .ZN(n1111) );
XNOR2_X1 U798 ( .A(n1117), .B(n1118), .ZN(n1116) );
NAND2_X1 U799 ( .A1(KEYINPUT20), .A2(n1119), .ZN(n1117) );
NOR2_X1 U800 ( .A1(n1120), .A2(n1121), .ZN(n1103) );
AND2_X1 U801 ( .A1(G227), .A2(G900), .ZN(n1120) );
XOR2_X1 U802 ( .A(n1122), .B(n1123), .Z(G69) );
XOR2_X1 U803 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND2_X1 U804 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U805 ( .A1(G953), .A2(n1128), .ZN(n1127) );
XNOR2_X1 U806 ( .A(KEYINPUT19), .B(n1129), .ZN(n1126) );
NAND2_X1 U807 ( .A1(n1130), .A2(n1040), .ZN(n1124) );
NAND2_X1 U808 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U809 ( .A(n1133), .B(KEYINPUT3), .Z(n1131) );
NOR2_X1 U810 ( .A1(n1134), .A2(n1121), .ZN(n1122) );
XNOR2_X1 U811 ( .A(n1040), .B(KEYINPUT33), .ZN(n1121) );
AND2_X1 U812 ( .A1(G224), .A2(G898), .ZN(n1134) );
NOR2_X1 U813 ( .A1(n1135), .A2(n1136), .ZN(G66) );
XOR2_X1 U814 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
XOR2_X1 U816 ( .A(n1141), .B(KEYINPUT62), .Z(n1135) );
NAND2_X1 U817 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U818 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
INV_X1 U819 ( .A(KEYINPUT2), .ZN(n1145) );
NAND3_X1 U820 ( .A1(G952), .A2(G953), .A3(KEYINPUT2), .ZN(n1142) );
NOR2_X1 U821 ( .A1(n1144), .A2(n1146), .ZN(G63) );
XNOR2_X1 U822 ( .A(n1147), .B(n1148), .ZN(n1146) );
NOR2_X1 U823 ( .A1(n1149), .A2(n1140), .ZN(n1148) );
NOR2_X1 U824 ( .A1(n1150), .A2(n1151), .ZN(G60) );
XOR2_X1 U825 ( .A(KEYINPUT56), .B(n1144), .Z(n1151) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1150) );
NOR2_X1 U827 ( .A1(n1095), .A2(n1140), .ZN(n1153) );
XOR2_X1 U828 ( .A(G104), .B(n1154), .Z(G6) );
NOR2_X1 U829 ( .A1(n1155), .A2(n1055), .ZN(n1154) );
NOR2_X1 U830 ( .A1(n1144), .A2(n1156), .ZN(G57) );
XOR2_X1 U831 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U832 ( .A(n1159), .B(n1160), .ZN(n1158) );
NOR2_X1 U833 ( .A1(n1161), .A2(n1140), .ZN(n1160) );
XNOR2_X1 U834 ( .A(G101), .B(n1162), .ZN(n1157) );
NAND2_X1 U835 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NAND2_X1 U836 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
INV_X1 U837 ( .A(n1167), .ZN(n1166) );
NAND2_X1 U838 ( .A1(KEYINPUT42), .A2(n1168), .ZN(n1165) );
OR2_X1 U839 ( .A1(n1169), .A2(KEYINPUT8), .ZN(n1168) );
NAND2_X1 U840 ( .A1(n1169), .A2(n1170), .ZN(n1163) );
NAND2_X1 U841 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
INV_X1 U842 ( .A(KEYINPUT8), .ZN(n1172) );
NAND2_X1 U843 ( .A1(n1167), .A2(KEYINPUT42), .ZN(n1171) );
NOR2_X1 U844 ( .A1(n1173), .A2(n1174), .ZN(n1167) );
AND2_X1 U845 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NOR2_X1 U846 ( .A1(n1144), .A2(n1177), .ZN(G54) );
XOR2_X1 U847 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U848 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U849 ( .A(n1182), .B(n1183), .Z(n1178) );
XNOR2_X1 U850 ( .A(n1184), .B(n1185), .ZN(n1183) );
NOR2_X1 U851 ( .A1(n1186), .A2(n1140), .ZN(n1185) );
NOR3_X1 U852 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(G51) );
AND2_X1 U853 ( .A1(n1144), .A2(KEYINPUT23), .ZN(n1189) );
NOR2_X1 U854 ( .A1(n1040), .A2(G952), .ZN(n1144) );
NOR3_X1 U855 ( .A1(KEYINPUT23), .A2(n1040), .A3(n1037), .ZN(n1188) );
INV_X1 U856 ( .A(G952), .ZN(n1037) );
NOR2_X1 U857 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
XOR2_X1 U858 ( .A(n1192), .B(n1193), .Z(n1191) );
NOR2_X1 U859 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NOR2_X1 U860 ( .A1(n1093), .A2(n1140), .ZN(n1192) );
NAND2_X1 U861 ( .A1(G902), .A2(n1038), .ZN(n1140) );
NAND3_X1 U862 ( .A1(n1132), .A2(n1133), .A3(n1196), .ZN(n1038) );
INV_X1 U863 ( .A(n1107), .ZN(n1196) );
NAND4_X1 U864 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1107) );
AND4_X1 U865 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
OR3_X1 U866 ( .A1(n1205), .A2(n1056), .A3(n1206), .ZN(n1204) );
XNOR2_X1 U867 ( .A(KEYINPUT0), .B(n1067), .ZN(n1205) );
NOR2_X1 U868 ( .A1(n1207), .A2(n1208), .ZN(n1199) );
AND4_X1 U869 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1132) );
AND4_X1 U870 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1212) );
INV_X1 U871 ( .A(n1033), .ZN(n1213) );
NOR2_X1 U872 ( .A1(n1056), .A2(n1155), .ZN(n1033) );
NAND2_X1 U873 ( .A1(n1053), .A2(n1217), .ZN(n1155) );
NAND4_X1 U874 ( .A1(n1061), .A2(n1057), .A3(n1218), .A4(n1219), .ZN(n1211) );
NAND2_X1 U875 ( .A1(KEYINPUT58), .A2(n1220), .ZN(n1219) );
NAND2_X1 U876 ( .A1(n1221), .A2(n1222), .ZN(n1218) );
INV_X1 U877 ( .A(KEYINPUT58), .ZN(n1222) );
NAND3_X1 U878 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1221) );
NAND3_X1 U879 ( .A1(n1217), .A2(n1226), .A3(n1227), .ZN(n1209) );
XOR2_X1 U880 ( .A(KEYINPUT1), .B(n1053), .Z(n1226) );
AND2_X1 U881 ( .A1(n1195), .A2(n1194), .ZN(n1190) );
XOR2_X1 U882 ( .A(n1228), .B(n1129), .Z(n1194) );
XOR2_X1 U883 ( .A(n1229), .B(n1230), .Z(n1228) );
NOR2_X1 U884 ( .A1(KEYINPUT13), .A2(n1231), .ZN(n1230) );
XNOR2_X1 U885 ( .A(G125), .B(n1176), .ZN(n1231) );
INV_X1 U886 ( .A(KEYINPUT16), .ZN(n1195) );
XNOR2_X1 U887 ( .A(G146), .B(n1197), .ZN(G48) );
OR3_X1 U888 ( .A1(n1232), .A2(n1233), .A3(n1055), .ZN(n1197) );
XNOR2_X1 U889 ( .A(n1234), .B(n1235), .ZN(G45) );
NOR2_X1 U890 ( .A1(KEYINPUT45), .A2(n1203), .ZN(n1235) );
NAND4_X1 U891 ( .A1(n1236), .A2(n1223), .A3(n1061), .A4(n1237), .ZN(n1203) );
NOR3_X1 U892 ( .A1(n1238), .A2(n1239), .A3(n1233), .ZN(n1237) );
XNOR2_X1 U893 ( .A(n1184), .B(n1240), .ZN(G42) );
NOR2_X1 U894 ( .A1(KEYINPUT9), .A2(n1202), .ZN(n1240) );
NAND3_X1 U895 ( .A1(n1241), .A2(n1062), .A3(n1227), .ZN(n1202) );
XNOR2_X1 U896 ( .A(G137), .B(n1198), .ZN(G39) );
NAND4_X1 U897 ( .A1(n1242), .A2(n1241), .A3(n1057), .A4(n1243), .ZN(n1198) );
XOR2_X1 U898 ( .A(n1244), .B(n1245), .Z(G36) );
NOR2_X1 U899 ( .A1(KEYINPUT43), .A2(n1246), .ZN(n1245) );
AND2_X1 U900 ( .A1(n1241), .A2(n1247), .ZN(n1246) );
INV_X1 U901 ( .A(n1206), .ZN(n1241) );
XNOR2_X1 U902 ( .A(G134), .B(KEYINPUT21), .ZN(n1244) );
XNOR2_X1 U903 ( .A(n1119), .B(n1208), .ZN(G33) );
NOR3_X1 U904 ( .A1(n1055), .A2(n1206), .A3(n1067), .ZN(n1208) );
NAND4_X1 U905 ( .A1(n1046), .A2(n1223), .A3(n1248), .A4(n1049), .ZN(n1206) );
INV_X1 U906 ( .A(n1227), .ZN(n1055) );
XOR2_X1 U907 ( .A(G128), .B(n1207), .Z(G30) );
NOR3_X1 U908 ( .A1(n1056), .A2(n1233), .A3(n1232), .ZN(n1207) );
NAND4_X1 U909 ( .A1(n1242), .A2(n1223), .A3(n1080), .A4(n1243), .ZN(n1232) );
XOR2_X1 U910 ( .A(n1249), .B(n1250), .Z(G3) );
NOR3_X1 U911 ( .A1(n1067), .A2(n1220), .A3(n1064), .ZN(n1250) );
INV_X1 U912 ( .A(n1057), .ZN(n1064) );
INV_X1 U913 ( .A(n1217), .ZN(n1220) );
NOR2_X1 U914 ( .A1(KEYINPUT28), .A2(n1251), .ZN(n1249) );
NAND2_X1 U915 ( .A1(n1252), .A2(n1253), .ZN(G27) );
NAND2_X1 U916 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U917 ( .A1(G125), .A2(n1256), .ZN(n1252) );
NAND2_X1 U918 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND2_X1 U919 ( .A1(KEYINPUT35), .A2(n1259), .ZN(n1258) );
INV_X1 U920 ( .A(n1201), .ZN(n1259) );
OR2_X1 U921 ( .A1(n1254), .A2(KEYINPUT35), .ZN(n1257) );
NOR2_X1 U922 ( .A1(KEYINPUT47), .A2(n1201), .ZN(n1254) );
NAND4_X1 U923 ( .A1(n1227), .A2(n1062), .A3(n1260), .A4(n1047), .ZN(n1201) );
NOR2_X1 U924 ( .A1(n1233), .A2(n1238), .ZN(n1260) );
INV_X1 U925 ( .A(n1248), .ZN(n1233) );
NAND2_X1 U926 ( .A1(n1081), .A2(n1261), .ZN(n1248) );
NAND4_X1 U927 ( .A1(G902), .A2(G953), .A3(n1262), .A4(n1113), .ZN(n1261) );
INV_X1 U928 ( .A(G900), .ZN(n1113) );
XNOR2_X1 U929 ( .A(G122), .B(n1210), .ZN(G24) );
NAND4_X1 U930 ( .A1(n1263), .A2(n1053), .A3(n1236), .A4(n1264), .ZN(n1210) );
NOR2_X1 U931 ( .A1(n1243), .A2(n1242), .ZN(n1053) );
XOR2_X1 U932 ( .A(G119), .B(n1265), .Z(G21) );
NOR2_X1 U933 ( .A1(KEYINPUT37), .A2(n1216), .ZN(n1265) );
NAND4_X1 U934 ( .A1(n1242), .A2(n1263), .A3(n1057), .A4(n1243), .ZN(n1216) );
NAND3_X1 U935 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(G18) );
NAND2_X1 U936 ( .A1(KEYINPUT40), .A2(n1269), .ZN(n1268) );
NAND3_X1 U937 ( .A1(G116), .A2(n1270), .A3(n1215), .ZN(n1267) );
NAND2_X1 U938 ( .A1(n1271), .A2(n1272), .ZN(n1266) );
NAND2_X1 U939 ( .A1(n1273), .A2(n1270), .ZN(n1272) );
INV_X1 U940 ( .A(KEYINPUT40), .ZN(n1270) );
XNOR2_X1 U941 ( .A(KEYINPUT6), .B(n1269), .ZN(n1273) );
INV_X1 U942 ( .A(n1215), .ZN(n1271) );
NAND2_X1 U943 ( .A1(n1263), .A2(n1247), .ZN(n1215) );
NOR2_X1 U944 ( .A1(n1067), .A2(n1056), .ZN(n1247) );
NAND2_X1 U945 ( .A1(n1239), .A2(n1236), .ZN(n1056) );
NOR3_X1 U946 ( .A1(n1238), .A2(n1225), .A3(n1075), .ZN(n1263) );
INV_X1 U947 ( .A(n1080), .ZN(n1238) );
XOR2_X1 U948 ( .A(n1224), .B(KEYINPUT5), .Z(n1080) );
XNOR2_X1 U949 ( .A(G113), .B(n1214), .ZN(G15) );
NAND4_X1 U950 ( .A1(n1061), .A2(n1227), .A3(n1274), .A4(n1047), .ZN(n1214) );
INV_X1 U951 ( .A(n1075), .ZN(n1047) );
NAND2_X1 U952 ( .A1(n1079), .A2(n1275), .ZN(n1075) );
NOR2_X1 U953 ( .A1(n1225), .A2(n1276), .ZN(n1274) );
NOR2_X1 U954 ( .A1(n1236), .A2(n1239), .ZN(n1227) );
INV_X1 U955 ( .A(n1264), .ZN(n1239) );
INV_X1 U956 ( .A(n1067), .ZN(n1061) );
NAND2_X1 U957 ( .A1(n1242), .A2(n1084), .ZN(n1067) );
XNOR2_X1 U958 ( .A(G110), .B(n1133), .ZN(G12) );
NAND3_X1 U959 ( .A1(n1062), .A2(n1217), .A3(n1057), .ZN(n1133) );
NOR2_X1 U960 ( .A1(n1264), .A2(n1236), .ZN(n1057) );
XOR2_X1 U961 ( .A(n1098), .B(KEYINPUT39), .Z(n1236) );
XNOR2_X1 U962 ( .A(n1277), .B(n1149), .ZN(n1098) );
INV_X1 U963 ( .A(G478), .ZN(n1149) );
NAND2_X1 U964 ( .A1(n1147), .A2(n1278), .ZN(n1277) );
XNOR2_X1 U965 ( .A(n1279), .B(n1280), .ZN(n1147) );
AND3_X1 U966 ( .A1(G234), .A2(n1040), .A3(G217), .ZN(n1280) );
NAND2_X1 U967 ( .A1(KEYINPUT55), .A2(n1281), .ZN(n1279) );
XOR2_X1 U968 ( .A(n1282), .B(n1283), .Z(n1281) );
XNOR2_X1 U969 ( .A(n1032), .B(n1284), .ZN(n1283) );
XNOR2_X1 U970 ( .A(n1269), .B(n1285), .ZN(n1282) );
XOR2_X1 U971 ( .A(G134), .B(G122), .Z(n1285) );
INV_X1 U972 ( .A(G116), .ZN(n1269) );
NAND2_X1 U973 ( .A1(n1286), .A2(n1096), .ZN(n1264) );
NAND2_X1 U974 ( .A1(n1094), .A2(n1095), .ZN(n1096) );
INV_X1 U975 ( .A(G475), .ZN(n1095) );
NAND2_X1 U976 ( .A1(G475), .A2(n1287), .ZN(n1286) );
XOR2_X1 U977 ( .A(KEYINPUT18), .B(n1094), .Z(n1287) );
NOR2_X1 U978 ( .A1(n1152), .A2(G902), .ZN(n1094) );
XOR2_X1 U979 ( .A(n1288), .B(n1289), .Z(n1152) );
XNOR2_X1 U980 ( .A(n1112), .B(n1290), .ZN(n1289) );
XOR2_X1 U981 ( .A(n1291), .B(n1292), .Z(n1290) );
NAND2_X1 U982 ( .A1(KEYINPUT44), .A2(n1234), .ZN(n1291) );
XNOR2_X1 U983 ( .A(G125), .B(n1184), .ZN(n1112) );
XOR2_X1 U984 ( .A(n1293), .B(n1294), .Z(n1288) );
XNOR2_X1 U985 ( .A(n1119), .B(G104), .ZN(n1294) );
XOR2_X1 U986 ( .A(n1295), .B(n1296), .Z(n1293) );
AND3_X1 U987 ( .A1(G214), .A2(n1040), .A3(n1297), .ZN(n1296) );
NAND2_X1 U988 ( .A1(KEYINPUT60), .A2(n1298), .ZN(n1295) );
NOR3_X1 U989 ( .A1(n1276), .A2(n1225), .A3(n1077), .ZN(n1217) );
INV_X1 U990 ( .A(n1223), .ZN(n1077) );
NOR2_X1 U991 ( .A1(n1079), .A2(n1078), .ZN(n1223) );
INV_X1 U992 ( .A(n1275), .ZN(n1078) );
NAND2_X1 U993 ( .A1(G221), .A2(n1299), .ZN(n1275) );
XNOR2_X1 U994 ( .A(n1300), .B(n1186), .ZN(n1079) );
INV_X1 U995 ( .A(G469), .ZN(n1186) );
NAND2_X1 U996 ( .A1(n1301), .A2(n1278), .ZN(n1300) );
XOR2_X1 U997 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U998 ( .A(n1304), .B(n1181), .ZN(n1303) );
XOR2_X1 U999 ( .A(n1305), .B(n1175), .Z(n1181) );
NAND2_X1 U1000 ( .A1(G227), .A2(n1040), .ZN(n1305) );
NAND2_X1 U1001 ( .A1(KEYINPUT36), .A2(n1184), .ZN(n1304) );
XNOR2_X1 U1002 ( .A(G110), .B(n1306), .ZN(n1302) );
NAND2_X1 U1003 ( .A1(KEYINPUT31), .A2(n1307), .ZN(n1306) );
XNOR2_X1 U1004 ( .A(n1251), .B(n1180), .ZN(n1307) );
XNOR2_X1 U1005 ( .A(n1308), .B(n1118), .ZN(n1180) );
XNOR2_X1 U1006 ( .A(n1309), .B(KEYINPUT61), .ZN(n1118) );
NAND2_X1 U1007 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NAND2_X1 U1008 ( .A1(n1312), .A2(n1298), .ZN(n1311) );
XNOR2_X1 U1009 ( .A(n1284), .B(KEYINPUT49), .ZN(n1312) );
XNOR2_X1 U1010 ( .A(G104), .B(G107), .ZN(n1308) );
AND2_X1 U1011 ( .A1(n1081), .A2(n1313), .ZN(n1225) );
NAND4_X1 U1012 ( .A1(G902), .A2(G953), .A3(n1262), .A4(n1128), .ZN(n1313) );
INV_X1 U1013 ( .A(G898), .ZN(n1128) );
NAND3_X1 U1014 ( .A1(n1262), .A2(n1040), .A3(G952), .ZN(n1081) );
NAND2_X1 U1015 ( .A1(G237), .A2(G234), .ZN(n1262) );
INV_X1 U1016 ( .A(n1224), .ZN(n1276) );
NOR2_X1 U1017 ( .A1(n1046), .A2(n1074), .ZN(n1224) );
INV_X1 U1018 ( .A(n1049), .ZN(n1074) );
NAND2_X1 U1019 ( .A1(n1314), .A2(n1315), .ZN(n1049) );
XNOR2_X1 U1020 ( .A(G214), .B(KEYINPUT50), .ZN(n1314) );
XNOR2_X1 U1021 ( .A(n1092), .B(n1093), .ZN(n1046) );
NAND2_X1 U1022 ( .A1(G210), .A2(n1315), .ZN(n1093) );
NAND2_X1 U1023 ( .A1(n1316), .A2(n1278), .ZN(n1315) );
XNOR2_X1 U1024 ( .A(G237), .B(KEYINPUT22), .ZN(n1316) );
NAND2_X1 U1025 ( .A1(n1317), .A2(n1278), .ZN(n1092) );
XOR2_X1 U1026 ( .A(n1318), .B(n1319), .Z(n1317) );
XNOR2_X1 U1027 ( .A(n1176), .B(n1320), .ZN(n1319) );
NOR2_X1 U1028 ( .A1(KEYINPUT24), .A2(n1129), .ZN(n1320) );
XOR2_X1 U1029 ( .A(n1321), .B(n1322), .Z(n1129) );
XOR2_X1 U1030 ( .A(n1182), .B(n1292), .Z(n1322) );
XOR2_X1 U1031 ( .A(G113), .B(G122), .Z(n1292) );
XNOR2_X1 U1032 ( .A(n1251), .B(G110), .ZN(n1182) );
XOR2_X1 U1033 ( .A(n1323), .B(n1324), .Z(n1321) );
XNOR2_X1 U1034 ( .A(G104), .B(n1325), .ZN(n1324) );
NAND2_X1 U1035 ( .A1(KEYINPUT53), .A2(n1032), .ZN(n1325) );
INV_X1 U1036 ( .A(G107), .ZN(n1032) );
NAND2_X1 U1037 ( .A1(KEYINPUT63), .A2(n1326), .ZN(n1323) );
XNOR2_X1 U1038 ( .A(n1327), .B(n1328), .ZN(n1318) );
NOR2_X1 U1039 ( .A1(KEYINPUT52), .A2(n1229), .ZN(n1328) );
NAND2_X1 U1040 ( .A1(G224), .A2(n1329), .ZN(n1229) );
XNOR2_X1 U1041 ( .A(KEYINPUT46), .B(n1040), .ZN(n1329) );
NOR2_X1 U1042 ( .A1(G125), .A2(KEYINPUT51), .ZN(n1327) );
NOR2_X1 U1043 ( .A1(n1242), .A2(n1084), .ZN(n1062) );
INV_X1 U1044 ( .A(n1243), .ZN(n1084) );
XOR2_X1 U1045 ( .A(n1330), .B(n1139), .Z(n1243) );
NAND2_X1 U1046 ( .A1(G217), .A2(n1299), .ZN(n1139) );
NAND2_X1 U1047 ( .A1(G234), .A2(n1278), .ZN(n1299) );
OR2_X1 U1048 ( .A1(n1138), .A2(G902), .ZN(n1330) );
XNOR2_X1 U1049 ( .A(n1331), .B(n1332), .ZN(n1138) );
XOR2_X1 U1050 ( .A(n1333), .B(n1334), .Z(n1332) );
XOR2_X1 U1051 ( .A(n1335), .B(n1336), .Z(n1334) );
AND3_X1 U1052 ( .A1(G221), .A2(n1040), .A3(G234), .ZN(n1336) );
NAND2_X1 U1053 ( .A1(KEYINPUT27), .A2(G110), .ZN(n1335) );
NAND2_X1 U1054 ( .A1(n1337), .A2(n1338), .ZN(n1333) );
NAND2_X1 U1055 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
XNOR2_X1 U1056 ( .A(G140), .B(n1341), .ZN(n1340) );
XNOR2_X1 U1057 ( .A(KEYINPUT34), .B(n1342), .ZN(n1339) );
NAND2_X1 U1058 ( .A1(n1343), .A2(n1344), .ZN(n1337) );
XNOR2_X1 U1059 ( .A(n1345), .B(n1342), .ZN(n1344) );
XNOR2_X1 U1060 ( .A(KEYINPUT38), .B(KEYINPUT10), .ZN(n1345) );
XNOR2_X1 U1061 ( .A(n1341), .B(n1184), .ZN(n1343) );
INV_X1 U1062 ( .A(G140), .ZN(n1184) );
NAND2_X1 U1063 ( .A1(KEYINPUT4), .A2(n1255), .ZN(n1341) );
INV_X1 U1064 ( .A(G125), .ZN(n1255) );
XOR2_X1 U1065 ( .A(n1346), .B(n1347), .Z(n1331) );
XOR2_X1 U1066 ( .A(KEYINPUT25), .B(G137), .Z(n1347) );
XNOR2_X1 U1067 ( .A(G119), .B(G128), .ZN(n1346) );
XOR2_X1 U1068 ( .A(n1348), .B(n1102), .Z(n1242) );
AND2_X1 U1069 ( .A1(n1349), .A2(n1278), .ZN(n1102) );
INV_X1 U1070 ( .A(G902), .ZN(n1278) );
XOR2_X1 U1071 ( .A(n1350), .B(n1351), .Z(n1349) );
XOR2_X1 U1072 ( .A(n1352), .B(n1159), .Z(n1351) );
NAND3_X1 U1073 ( .A1(n1297), .A2(n1040), .A3(G210), .ZN(n1159) );
INV_X1 U1074 ( .A(G953), .ZN(n1040) );
INV_X1 U1075 ( .A(G237), .ZN(n1297) );
NAND2_X1 U1076 ( .A1(KEYINPUT12), .A2(n1251), .ZN(n1352) );
INV_X1 U1077 ( .A(G101), .ZN(n1251) );
XOR2_X1 U1078 ( .A(n1169), .B(n1353), .Z(n1350) );
NOR2_X1 U1079 ( .A1(n1173), .A2(n1354), .ZN(n1353) );
XOR2_X1 U1080 ( .A(n1355), .B(KEYINPUT14), .Z(n1354) );
NAND2_X1 U1081 ( .A1(n1175), .A2(n1176), .ZN(n1355) );
NOR2_X1 U1082 ( .A1(n1176), .A2(n1175), .ZN(n1173) );
XOR2_X1 U1083 ( .A(n1119), .B(n1115), .Z(n1175) );
XOR2_X1 U1084 ( .A(G134), .B(G137), .Z(n1115) );
INV_X1 U1085 ( .A(G131), .ZN(n1119) );
NAND2_X1 U1086 ( .A1(n1310), .A2(n1356), .ZN(n1176) );
NAND2_X1 U1087 ( .A1(n1357), .A2(n1298), .ZN(n1356) );
XOR2_X1 U1088 ( .A(KEYINPUT15), .B(n1284), .Z(n1357) );
NAND2_X1 U1089 ( .A1(n1342), .A2(n1284), .ZN(n1310) );
XNOR2_X1 U1090 ( .A(G128), .B(n1234), .ZN(n1284) );
INV_X1 U1091 ( .A(G143), .ZN(n1234) );
INV_X1 U1092 ( .A(n1298), .ZN(n1342) );
XOR2_X1 U1093 ( .A(G146), .B(KEYINPUT32), .Z(n1298) );
XOR2_X1 U1094 ( .A(G113), .B(n1326), .Z(n1169) );
XNOR2_X1 U1095 ( .A(G119), .B(G116), .ZN(n1326) );
NAND2_X1 U1096 ( .A1(KEYINPUT59), .A2(n1100), .ZN(n1348) );
XOR2_X1 U1097 ( .A(n1161), .B(KEYINPUT11), .Z(n1100) );
INV_X1 U1098 ( .A(G472), .ZN(n1161) );
endmodule


