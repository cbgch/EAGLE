//Key = 1101100101101100100100011010001110101000110111010010000010110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345;

XNOR2_X1 U731 ( .A(G107), .B(n1020), .ZN(G9) );
NAND4_X1 U732 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1020) );
XNOR2_X1 U733 ( .A(n1025), .B(KEYINPUT56), .ZN(n1021) );
NOR2_X1 U734 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR3_X1 U735 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
NAND3_X1 U736 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1028) );
NAND2_X1 U737 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U738 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND4_X1 U739 ( .A1(n1024), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1037) );
NAND2_X1 U740 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NAND2_X1 U741 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U742 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U743 ( .A1(n1047), .A2(n1048), .ZN(n1041) );
NAND2_X1 U744 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U745 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XNOR2_X1 U746 ( .A(KEYINPUT27), .B(n1053), .ZN(n1052) );
NAND4_X1 U747 ( .A1(n1054), .A2(n1055), .A3(n1043), .A4(n1056), .ZN(n1036) );
NOR2_X1 U748 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
INV_X1 U749 ( .A(n1047), .ZN(n1058) );
NOR2_X1 U750 ( .A1(n1059), .A2(n1038), .ZN(n1057) );
NOR2_X1 U751 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U752 ( .A1(n1062), .A2(n1061), .ZN(n1055) );
INV_X1 U753 ( .A(n1024), .ZN(n1061) );
NAND4_X1 U754 ( .A1(n1060), .A2(n1063), .A3(n1064), .A4(n1040), .ZN(n1054) );
INV_X1 U755 ( .A(n1065), .ZN(n1034) );
NOR3_X1 U756 ( .A1(n1066), .A2(G953), .A3(G952), .ZN(n1026) );
INV_X1 U757 ( .A(n1031), .ZN(n1066) );
NAND4_X1 U758 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1031) );
NOR4_X1 U759 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1070) );
NOR3_X1 U760 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1074) );
INV_X1 U761 ( .A(KEYINPUT40), .ZN(n1075) );
NOR2_X1 U762 ( .A1(KEYINPUT40), .A2(G478), .ZN(n1073) );
XNOR2_X1 U763 ( .A(G469), .B(n1078), .ZN(n1072) );
NAND3_X1 U764 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1071) );
XOR2_X1 U765 ( .A(n1082), .B(n1083), .Z(n1080) );
XOR2_X1 U766 ( .A(n1084), .B(KEYINPUT23), .Z(n1083) );
XOR2_X1 U767 ( .A(n1085), .B(n1086), .Z(n1079) );
NAND2_X1 U768 ( .A1(KEYINPUT59), .A2(n1087), .ZN(n1086) );
NOR3_X1 U769 ( .A1(n1062), .A2(n1088), .A3(n1089), .ZN(n1069) );
INV_X1 U770 ( .A(n1090), .ZN(n1088) );
XOR2_X1 U771 ( .A(n1091), .B(n1092), .Z(G72) );
NOR2_X1 U772 ( .A1(KEYINPUT63), .A2(n1093), .ZN(n1092) );
XOR2_X1 U773 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U774 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U775 ( .A1(G953), .A2(n1098), .ZN(n1097) );
XOR2_X1 U776 ( .A(n1099), .B(n1100), .Z(n1096) );
XNOR2_X1 U777 ( .A(n1101), .B(n1102), .ZN(n1100) );
XOR2_X1 U778 ( .A(n1103), .B(n1104), .Z(n1099) );
NOR2_X1 U779 ( .A1(KEYINPUT51), .A2(n1105), .ZN(n1104) );
XOR2_X1 U780 ( .A(G128), .B(n1106), .Z(n1105) );
XNOR2_X1 U781 ( .A(KEYINPUT24), .B(KEYINPUT19), .ZN(n1103) );
NAND2_X1 U782 ( .A1(n1029), .A2(n1032), .ZN(n1094) );
NAND2_X1 U783 ( .A1(G953), .A2(n1107), .ZN(n1091) );
NAND2_X1 U784 ( .A1(G900), .A2(G227), .ZN(n1107) );
XOR2_X1 U785 ( .A(n1108), .B(n1109), .Z(G69) );
NOR2_X1 U786 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR3_X1 U787 ( .A1(n1032), .A2(n1112), .A3(n1113), .ZN(n1111) );
NOR2_X1 U788 ( .A1(G953), .A2(n1114), .ZN(n1110) );
NOR2_X1 U789 ( .A1(n1115), .A2(KEYINPUT17), .ZN(n1114) );
INV_X1 U790 ( .A(n1030), .ZN(n1115) );
NOR2_X1 U791 ( .A1(n1116), .A2(n1117), .ZN(n1108) );
XOR2_X1 U792 ( .A(n1118), .B(n1119), .Z(n1117) );
XNOR2_X1 U793 ( .A(n1120), .B(KEYINPUT43), .ZN(n1118) );
NOR2_X1 U794 ( .A1(G898), .A2(n1032), .ZN(n1116) );
NOR2_X1 U795 ( .A1(n1121), .A2(n1122), .ZN(G66) );
XNOR2_X1 U796 ( .A(n1123), .B(n1124), .ZN(n1122) );
NOR2_X1 U797 ( .A1(n1082), .A2(n1125), .ZN(n1124) );
NOR2_X1 U798 ( .A1(n1121), .A2(n1126), .ZN(G63) );
XOR2_X1 U799 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U800 ( .A1(n1077), .A2(n1125), .ZN(n1127) );
NOR2_X1 U801 ( .A1(n1121), .A2(n1129), .ZN(G60) );
XNOR2_X1 U802 ( .A(n1130), .B(n1131), .ZN(n1129) );
XOR2_X1 U803 ( .A(KEYINPUT62), .B(n1132), .Z(n1131) );
AND2_X1 U804 ( .A1(G475), .A2(n1133), .ZN(n1132) );
XOR2_X1 U805 ( .A(n1134), .B(n1135), .Z(G6) );
NOR2_X1 U806 ( .A1(KEYINPUT53), .A2(n1136), .ZN(n1135) );
NOR3_X1 U807 ( .A1(n1121), .A2(n1137), .A3(n1138), .ZN(G57) );
NOR2_X1 U808 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U809 ( .A(n1141), .B(n1142), .Z(n1140) );
OR2_X1 U810 ( .A1(n1143), .A2(KEYINPUT21), .ZN(n1141) );
INV_X1 U811 ( .A(n1144), .ZN(n1139) );
NOR2_X1 U812 ( .A1(n1144), .A2(n1145), .ZN(n1137) );
XOR2_X1 U813 ( .A(n1146), .B(n1142), .Z(n1145) );
XNOR2_X1 U814 ( .A(n1147), .B(n1148), .ZN(n1142) );
XOR2_X1 U815 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U816 ( .A1(n1087), .A2(n1125), .ZN(n1150) );
INV_X1 U817 ( .A(G472), .ZN(n1087) );
NAND2_X1 U818 ( .A1(n1143), .A2(n1151), .ZN(n1146) );
INV_X1 U819 ( .A(KEYINPUT21), .ZN(n1151) );
NOR2_X1 U820 ( .A1(n1121), .A2(n1152), .ZN(G54) );
XOR2_X1 U821 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR3_X1 U822 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1154) );
NOR2_X1 U823 ( .A1(KEYINPUT29), .A2(n1158), .ZN(n1157) );
NOR2_X1 U824 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
AND2_X1 U825 ( .A1(n1161), .A2(KEYINPUT11), .ZN(n1160) );
NOR3_X1 U826 ( .A1(KEYINPUT11), .A2(n1162), .A3(n1161), .ZN(n1159) );
NOR2_X1 U827 ( .A1(n1163), .A2(n1164), .ZN(n1156) );
INV_X1 U828 ( .A(KEYINPUT29), .ZN(n1164) );
NOR2_X1 U829 ( .A1(n1162), .A2(n1165), .ZN(n1163) );
XNOR2_X1 U830 ( .A(KEYINPUT11), .B(n1166), .ZN(n1165) );
NOR2_X1 U831 ( .A1(n1167), .A2(n1166), .ZN(n1155) );
XOR2_X1 U832 ( .A(n1168), .B(n1169), .Z(n1153) );
NOR2_X1 U833 ( .A1(n1170), .A2(n1125), .ZN(n1169) );
NAND2_X1 U834 ( .A1(n1171), .A2(KEYINPUT58), .ZN(n1168) );
XNOR2_X1 U835 ( .A(n1172), .B(n1173), .ZN(n1171) );
NOR2_X1 U836 ( .A1(n1121), .A2(n1174), .ZN(G51) );
XOR2_X1 U837 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U838 ( .A1(KEYINPUT10), .A2(n1177), .ZN(n1176) );
XOR2_X1 U839 ( .A(n1178), .B(n1179), .Z(n1177) );
XNOR2_X1 U840 ( .A(n1180), .B(n1181), .ZN(n1179) );
NOR2_X1 U841 ( .A1(n1182), .A2(KEYINPUT55), .ZN(n1180) );
NAND2_X1 U842 ( .A1(n1133), .A2(n1183), .ZN(n1175) );
XOR2_X1 U843 ( .A(KEYINPUT42), .B(G210), .Z(n1183) );
INV_X1 U844 ( .A(n1125), .ZN(n1133) );
NAND2_X1 U845 ( .A1(G902), .A2(n1184), .ZN(n1125) );
OR2_X1 U846 ( .A1(n1030), .A2(n1029), .ZN(n1184) );
NAND4_X1 U847 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1029) );
NOR4_X1 U848 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1188) );
NOR2_X1 U849 ( .A1(n1193), .A2(n1194), .ZN(n1187) );
NOR3_X1 U850 ( .A1(n1195), .A2(n1045), .A3(n1063), .ZN(n1194) );
INV_X1 U851 ( .A(n1196), .ZN(n1193) );
NAND4_X1 U852 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1030) );
NOR4_X1 U853 ( .A1(n1201), .A2(n1134), .A3(n1202), .A4(n1203), .ZN(n1200) );
INV_X1 U854 ( .A(n1204), .ZN(n1203) );
INV_X1 U855 ( .A(n1205), .ZN(n1202) );
AND4_X1 U856 ( .A1(n1206), .A2(n1022), .A3(n1024), .A4(n1025), .ZN(n1134) );
NOR2_X1 U857 ( .A1(n1207), .A2(n1208), .ZN(n1199) );
NOR2_X1 U858 ( .A1(n1209), .A2(n1060), .ZN(n1208) );
XOR2_X1 U859 ( .A(n1210), .B(KEYINPUT18), .Z(n1209) );
NOR3_X1 U860 ( .A1(n1045), .A2(n1211), .A3(n1064), .ZN(n1207) );
NAND4_X1 U861 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1197) );
NOR2_X1 U862 ( .A1(n1032), .A2(G952), .ZN(n1121) );
XNOR2_X1 U863 ( .A(G146), .B(n1196), .ZN(G48) );
NAND3_X1 U864 ( .A1(n1212), .A2(n1206), .A3(n1213), .ZN(n1196) );
XNOR2_X1 U865 ( .A(G143), .B(n1185), .ZN(G45) );
NAND4_X1 U866 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1185) );
XNOR2_X1 U867 ( .A(n1217), .B(n1218), .ZN(G42) );
NOR3_X1 U868 ( .A1(n1219), .A2(n1045), .A3(n1195), .ZN(n1218) );
XNOR2_X1 U869 ( .A(KEYINPUT1), .B(n1063), .ZN(n1219) );
XNOR2_X1 U870 ( .A(G137), .B(n1186), .ZN(G39) );
NAND3_X1 U871 ( .A1(n1212), .A2(n1047), .A3(n1220), .ZN(n1186) );
INV_X1 U872 ( .A(n1195), .ZN(n1220) );
XOR2_X1 U873 ( .A(G134), .B(n1192), .Z(G36) );
NOR3_X1 U874 ( .A1(n1064), .A2(n1046), .A3(n1195), .ZN(n1192) );
XOR2_X1 U875 ( .A(G131), .B(n1191), .Z(G33) );
NOR3_X1 U876 ( .A1(n1045), .A2(n1064), .A3(n1195), .ZN(n1191) );
NAND4_X1 U877 ( .A1(n1025), .A2(n1038), .A3(n1221), .A4(n1040), .ZN(n1195) );
XOR2_X1 U878 ( .A(G128), .B(n1190), .Z(G30) );
AND3_X1 U879 ( .A1(n1212), .A2(n1023), .A3(n1213), .ZN(n1190) );
AND3_X1 U880 ( .A1(n1222), .A2(n1221), .A3(n1025), .ZN(n1213) );
INV_X1 U881 ( .A(n1046), .ZN(n1023) );
XOR2_X1 U882 ( .A(G101), .B(n1223), .Z(G3) );
NOR2_X1 U883 ( .A1(n1060), .A2(n1210), .ZN(n1223) );
NAND4_X1 U884 ( .A1(n1214), .A2(n1025), .A3(n1047), .A4(n1224), .ZN(n1210) );
INV_X1 U885 ( .A(n1064), .ZN(n1214) );
INV_X1 U886 ( .A(n1222), .ZN(n1060) );
XOR2_X1 U887 ( .A(G125), .B(n1189), .Z(G27) );
AND4_X1 U888 ( .A1(n1222), .A2(n1221), .A3(n1043), .A4(n1225), .ZN(n1189) );
NOR2_X1 U889 ( .A1(n1045), .A2(n1063), .ZN(n1225) );
INV_X1 U890 ( .A(n1226), .ZN(n1063) );
NAND2_X1 U891 ( .A1(n1065), .A2(n1227), .ZN(n1221) );
NAND4_X1 U892 ( .A1(G902), .A2(n1228), .A3(n1229), .A4(n1098), .ZN(n1227) );
INV_X1 U893 ( .A(G900), .ZN(n1098) );
XNOR2_X1 U894 ( .A(KEYINPUT61), .B(n1032), .ZN(n1228) );
XNOR2_X1 U895 ( .A(G122), .B(n1198), .ZN(G24) );
NAND4_X1 U896 ( .A1(n1230), .A2(n1024), .A3(n1215), .A4(n1216), .ZN(n1198) );
NOR2_X1 U897 ( .A1(n1231), .A2(n1232), .ZN(n1024) );
NAND2_X1 U898 ( .A1(n1233), .A2(n1234), .ZN(G21) );
NAND2_X1 U899 ( .A1(G119), .A2(n1204), .ZN(n1234) );
XOR2_X1 U900 ( .A(n1235), .B(KEYINPUT20), .Z(n1233) );
OR2_X1 U901 ( .A1(n1204), .A2(G119), .ZN(n1235) );
NAND3_X1 U902 ( .A1(n1230), .A2(n1047), .A3(n1212), .ZN(n1204) );
AND2_X1 U903 ( .A1(n1232), .A2(n1231), .ZN(n1212) );
INV_X1 U904 ( .A(n1236), .ZN(n1232) );
INV_X1 U905 ( .A(n1211), .ZN(n1230) );
XOR2_X1 U906 ( .A(G116), .B(n1201), .Z(G18) );
NOR3_X1 U907 ( .A1(n1211), .A2(n1046), .A3(n1064), .ZN(n1201) );
NAND2_X1 U908 ( .A1(n1237), .A2(n1216), .ZN(n1046) );
XOR2_X1 U909 ( .A(KEYINPUT14), .B(n1238), .Z(n1237) );
XOR2_X1 U910 ( .A(G113), .B(n1239), .Z(G15) );
NOR3_X1 U911 ( .A1(n1240), .A2(n1211), .A3(n1045), .ZN(n1239) );
INV_X1 U912 ( .A(n1206), .ZN(n1045) );
NAND2_X1 U913 ( .A1(n1043), .A2(n1022), .ZN(n1211) );
NOR2_X1 U914 ( .A1(n1053), .A2(n1051), .ZN(n1043) );
INV_X1 U915 ( .A(n1068), .ZN(n1051) );
XNOR2_X1 U916 ( .A(KEYINPUT32), .B(n1064), .ZN(n1240) );
NAND2_X1 U917 ( .A1(n1231), .A2(n1236), .ZN(n1064) );
XNOR2_X1 U918 ( .A(G110), .B(n1205), .ZN(G12) );
NAND4_X1 U919 ( .A1(n1226), .A2(n1022), .A3(n1025), .A4(n1047), .ZN(n1205) );
NAND2_X1 U920 ( .A1(n1241), .A2(n1242), .ZN(n1047) );
OR3_X1 U921 ( .A1(n1216), .A2(n1215), .A3(KEYINPUT14), .ZN(n1242) );
NAND2_X1 U922 ( .A1(KEYINPUT14), .A2(n1206), .ZN(n1241) );
NOR2_X1 U923 ( .A1(n1216), .A2(n1238), .ZN(n1206) );
INV_X1 U924 ( .A(n1215), .ZN(n1238) );
NAND2_X1 U925 ( .A1(n1243), .A2(n1067), .ZN(n1215) );
NAND2_X1 U926 ( .A1(G475), .A2(n1244), .ZN(n1067) );
XNOR2_X1 U927 ( .A(n1089), .B(KEYINPUT22), .ZN(n1243) );
NOR2_X1 U928 ( .A1(n1244), .A2(G475), .ZN(n1089) );
NAND2_X1 U929 ( .A1(n1130), .A2(n1245), .ZN(n1244) );
XNOR2_X1 U930 ( .A(n1246), .B(n1247), .ZN(n1130) );
XOR2_X1 U931 ( .A(n1248), .B(n1249), .Z(n1247) );
XNOR2_X1 U932 ( .A(n1250), .B(n1251), .ZN(n1249) );
NAND3_X1 U933 ( .A1(n1252), .A2(n1032), .A3(n1253), .ZN(n1250) );
XOR2_X1 U934 ( .A(KEYINPUT48), .B(G214), .Z(n1253) );
NAND2_X1 U935 ( .A1(KEYINPUT0), .A2(n1254), .ZN(n1248) );
XNOR2_X1 U936 ( .A(n1255), .B(n1256), .ZN(n1246) );
INV_X1 U937 ( .A(n1101), .ZN(n1256) );
XNOR2_X1 U938 ( .A(n1257), .B(n1258), .ZN(n1101) );
NAND2_X1 U939 ( .A1(KEYINPUT4), .A2(n1259), .ZN(n1255) );
XNOR2_X1 U940 ( .A(n1136), .B(n1260), .ZN(n1259) );
XOR2_X1 U941 ( .A(G122), .B(G113), .Z(n1260) );
NAND2_X1 U942 ( .A1(n1261), .A2(n1090), .ZN(n1216) );
NAND2_X1 U943 ( .A1(n1076), .A2(n1077), .ZN(n1090) );
INV_X1 U944 ( .A(G478), .ZN(n1077) );
XOR2_X1 U945 ( .A(KEYINPUT7), .B(n1262), .Z(n1261) );
NOR2_X1 U946 ( .A1(n1076), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U947 ( .A(G478), .B(KEYINPUT28), .ZN(n1263) );
NOR2_X1 U948 ( .A1(n1128), .A2(n1264), .ZN(n1076) );
XNOR2_X1 U949 ( .A(n1265), .B(n1266), .ZN(n1128) );
XOR2_X1 U950 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U951 ( .A(G116), .B(n1269), .Z(n1268) );
AND3_X1 U952 ( .A1(G217), .A2(n1032), .A3(G234), .ZN(n1269) );
XOR2_X1 U953 ( .A(n1270), .B(n1271), .Z(n1265) );
XNOR2_X1 U954 ( .A(KEYINPUT9), .B(n1254), .ZN(n1271) );
XNOR2_X1 U955 ( .A(G134), .B(G122), .ZN(n1270) );
INV_X1 U956 ( .A(n1049), .ZN(n1025) );
NAND2_X1 U957 ( .A1(n1053), .A2(n1068), .ZN(n1049) );
NAND2_X1 U958 ( .A1(G221), .A2(n1272), .ZN(n1068) );
NAND3_X1 U959 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1053) );
NAND2_X1 U960 ( .A1(G469), .A2(n1078), .ZN(n1275) );
NAND2_X1 U961 ( .A1(KEYINPUT39), .A2(n1276), .ZN(n1274) );
NAND2_X1 U962 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
XNOR2_X1 U963 ( .A(KEYINPUT13), .B(n1170), .ZN(n1278) );
NAND2_X1 U964 ( .A1(n1279), .A2(n1280), .ZN(n1273) );
INV_X1 U965 ( .A(KEYINPUT39), .ZN(n1280) );
NAND2_X1 U966 ( .A1(n1281), .A2(n1282), .ZN(n1279) );
NAND3_X1 U967 ( .A1(KEYINPUT13), .A2(n1277), .A3(n1170), .ZN(n1282) );
INV_X1 U968 ( .A(n1078), .ZN(n1277) );
NAND2_X1 U969 ( .A1(n1283), .A2(n1245), .ZN(n1078) );
XOR2_X1 U970 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U971 ( .A(n1172), .B(n1161), .ZN(n1285) );
INV_X1 U972 ( .A(n1166), .ZN(n1161) );
XNOR2_X1 U973 ( .A(G110), .B(n1217), .ZN(n1166) );
XOR2_X1 U974 ( .A(n1286), .B(n1287), .Z(n1284) );
XNOR2_X1 U975 ( .A(n1162), .B(KEYINPUT60), .ZN(n1287) );
INV_X1 U976 ( .A(n1167), .ZN(n1162) );
NAND2_X1 U977 ( .A1(n1288), .A2(G227), .ZN(n1167) );
XNOR2_X1 U978 ( .A(G953), .B(KEYINPUT15), .ZN(n1288) );
NAND2_X1 U979 ( .A1(KEYINPUT47), .A2(n1173), .ZN(n1286) );
XNOR2_X1 U980 ( .A(n1289), .B(n1290), .ZN(n1173) );
XOR2_X1 U981 ( .A(n1267), .B(n1106), .Z(n1290) );
XNOR2_X1 U982 ( .A(n1251), .B(n1291), .ZN(n1106) );
NOR2_X1 U983 ( .A1(KEYINPUT37), .A2(n1292), .ZN(n1291) );
INV_X1 U984 ( .A(G146), .ZN(n1251) );
XOR2_X1 U985 ( .A(G107), .B(G128), .Z(n1267) );
XNOR2_X1 U986 ( .A(n1293), .B(n1294), .ZN(n1289) );
NAND2_X1 U987 ( .A1(KEYINPUT41), .A2(n1136), .ZN(n1293) );
INV_X1 U988 ( .A(G104), .ZN(n1136) );
OR2_X1 U989 ( .A1(n1170), .A2(KEYINPUT13), .ZN(n1281) );
INV_X1 U990 ( .A(G469), .ZN(n1170) );
AND2_X1 U991 ( .A1(n1222), .A2(n1224), .ZN(n1022) );
NAND2_X1 U992 ( .A1(n1065), .A2(n1295), .ZN(n1224) );
NAND4_X1 U993 ( .A1(G953), .A2(G902), .A3(n1229), .A4(n1113), .ZN(n1295) );
INV_X1 U994 ( .A(G898), .ZN(n1113) );
NAND3_X1 U995 ( .A1(n1229), .A2(n1032), .A3(G952), .ZN(n1065) );
NAND2_X1 U996 ( .A1(G237), .A2(G234), .ZN(n1229) );
NOR2_X1 U997 ( .A1(n1038), .A2(n1062), .ZN(n1222) );
INV_X1 U998 ( .A(n1040), .ZN(n1062) );
NAND2_X1 U999 ( .A1(G214), .A2(n1296), .ZN(n1040) );
XNOR2_X1 U1000 ( .A(n1081), .B(KEYINPUT36), .ZN(n1038) );
XOR2_X1 U1001 ( .A(n1297), .B(n1298), .Z(n1081) );
AND2_X1 U1002 ( .A1(n1296), .A2(G210), .ZN(n1298) );
NAND2_X1 U1003 ( .A1(n1299), .A2(n1252), .ZN(n1296) );
NAND2_X1 U1004 ( .A1(n1300), .A2(n1245), .ZN(n1297) );
XOR2_X1 U1005 ( .A(n1178), .B(n1301), .Z(n1300) );
XNOR2_X1 U1006 ( .A(n1182), .B(n1181), .ZN(n1301) );
XOR2_X1 U1007 ( .A(n1302), .B(n1303), .Z(n1178) );
NOR2_X1 U1008 ( .A1(G953), .A2(n1112), .ZN(n1303) );
INV_X1 U1009 ( .A(G224), .ZN(n1112) );
NAND2_X1 U1010 ( .A1(n1304), .A2(n1305), .ZN(n1302) );
NAND2_X1 U1011 ( .A1(n1119), .A2(n1306), .ZN(n1305) );
INV_X1 U1012 ( .A(n1120), .ZN(n1306) );
NAND2_X1 U1013 ( .A1(n1120), .A2(n1307), .ZN(n1304) );
XNOR2_X1 U1014 ( .A(n1119), .B(KEYINPUT38), .ZN(n1307) );
XNOR2_X1 U1015 ( .A(n1308), .B(n1309), .ZN(n1119) );
XOR2_X1 U1016 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U1017 ( .A(G104), .B(n1312), .ZN(n1311) );
NOR2_X1 U1018 ( .A1(KEYINPUT46), .A2(n1313), .ZN(n1312) );
XNOR2_X1 U1019 ( .A(KEYINPUT12), .B(n1294), .ZN(n1313) );
NAND2_X1 U1020 ( .A1(KEYINPUT44), .A2(n1314), .ZN(n1310) );
XNOR2_X1 U1021 ( .A(G107), .B(n1315), .ZN(n1308) );
XOR2_X1 U1022 ( .A(KEYINPUT33), .B(G122), .Z(n1315) );
NOR2_X1 U1023 ( .A1(n1236), .A2(n1231), .ZN(n1226) );
XOR2_X1 U1024 ( .A(n1316), .B(n1085), .Z(n1231) );
NAND2_X1 U1025 ( .A1(n1317), .A2(n1245), .ZN(n1085) );
XOR2_X1 U1026 ( .A(n1318), .B(n1319), .Z(n1317) );
XNOR2_X1 U1027 ( .A(n1143), .B(n1320), .ZN(n1319) );
NOR2_X1 U1028 ( .A1(KEYINPUT54), .A2(n1294), .ZN(n1320) );
INV_X1 U1029 ( .A(n1147), .ZN(n1294) );
XOR2_X1 U1030 ( .A(G101), .B(KEYINPUT31), .Z(n1147) );
XNOR2_X1 U1031 ( .A(n1182), .B(n1321), .ZN(n1143) );
INV_X1 U1032 ( .A(n1172), .ZN(n1321) );
XOR2_X1 U1033 ( .A(n1102), .B(n1322), .Z(n1172) );
NOR2_X1 U1034 ( .A1(KEYINPUT52), .A2(n1323), .ZN(n1322) );
XOR2_X1 U1035 ( .A(KEYINPUT24), .B(n1257), .Z(n1323) );
XOR2_X1 U1036 ( .A(G131), .B(KEYINPUT50), .Z(n1257) );
XOR2_X1 U1037 ( .A(G134), .B(G137), .Z(n1102) );
AND2_X1 U1038 ( .A1(n1324), .A2(n1325), .ZN(n1182) );
NAND2_X1 U1039 ( .A1(G128), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1040 ( .A(n1327), .B(KEYINPUT8), .Z(n1324) );
OR2_X1 U1041 ( .A1(n1326), .A2(G128), .ZN(n1327) );
XOR2_X1 U1042 ( .A(G146), .B(n1292), .Z(n1326) );
XNOR2_X1 U1043 ( .A(n1254), .B(KEYINPUT57), .ZN(n1292) );
INV_X1 U1044 ( .A(G143), .ZN(n1254) );
XOR2_X1 U1045 ( .A(n1328), .B(n1149), .Z(n1318) );
AND3_X1 U1046 ( .A1(n1252), .A2(n1032), .A3(G210), .ZN(n1149) );
INV_X1 U1047 ( .A(G237), .ZN(n1252) );
NAND2_X1 U1048 ( .A1(KEYINPUT30), .A2(n1144), .ZN(n1328) );
XOR2_X1 U1049 ( .A(n1120), .B(KEYINPUT25), .Z(n1144) );
XOR2_X1 U1050 ( .A(G113), .B(n1329), .Z(n1120) );
XOR2_X1 U1051 ( .A(G119), .B(G116), .Z(n1329) );
NAND2_X1 U1052 ( .A1(KEYINPUT45), .A2(G472), .ZN(n1316) );
XNOR2_X1 U1053 ( .A(n1084), .B(n1330), .ZN(n1236) );
XOR2_X1 U1054 ( .A(KEYINPUT2), .B(n1331), .Z(n1330) );
NOR2_X1 U1055 ( .A1(KEYINPUT6), .A2(n1332), .ZN(n1331) );
XNOR2_X1 U1056 ( .A(KEYINPUT5), .B(n1082), .ZN(n1332) );
NAND2_X1 U1057 ( .A1(G217), .A2(n1272), .ZN(n1082) );
NAND2_X1 U1058 ( .A1(G234), .A2(n1299), .ZN(n1272) );
NAND2_X1 U1059 ( .A1(n1123), .A2(n1245), .ZN(n1084) );
INV_X1 U1060 ( .A(n1264), .ZN(n1245) );
XOR2_X1 U1061 ( .A(n1299), .B(KEYINPUT34), .Z(n1264) );
INV_X1 U1062 ( .A(G902), .ZN(n1299) );
XNOR2_X1 U1063 ( .A(n1333), .B(n1334), .ZN(n1123) );
XOR2_X1 U1064 ( .A(n1335), .B(n1336), .Z(n1334) );
XOR2_X1 U1065 ( .A(n1337), .B(n1338), .Z(n1336) );
AND3_X1 U1066 ( .A1(G221), .A2(n1032), .A3(G234), .ZN(n1338) );
INV_X1 U1067 ( .A(G953), .ZN(n1032) );
NAND2_X1 U1068 ( .A1(KEYINPUT16), .A2(G146), .ZN(n1337) );
NAND2_X1 U1069 ( .A1(n1339), .A2(n1340), .ZN(n1335) );
NAND2_X1 U1070 ( .A1(KEYINPUT3), .A2(n1258), .ZN(n1340) );
XNOR2_X1 U1071 ( .A(n1217), .B(n1181), .ZN(n1258) );
INV_X1 U1072 ( .A(n1341), .ZN(n1181) );
OR3_X1 U1073 ( .A1(n1217), .A2(n1341), .A3(KEYINPUT3), .ZN(n1339) );
XOR2_X1 U1074 ( .A(G125), .B(KEYINPUT49), .Z(n1341) );
INV_X1 U1075 ( .A(G140), .ZN(n1217) );
XOR2_X1 U1076 ( .A(n1342), .B(n1343), .Z(n1333) );
XNOR2_X1 U1077 ( .A(G137), .B(n1314), .ZN(n1343) );
INV_X1 U1078 ( .A(G110), .ZN(n1314) );
NAND2_X1 U1079 ( .A1(n1344), .A2(n1345), .ZN(n1342) );
XOR2_X1 U1080 ( .A(G128), .B(G119), .Z(n1345) );
XOR2_X1 U1081 ( .A(KEYINPUT35), .B(KEYINPUT26), .Z(n1344) );
endmodule


