//Key = 0001010100000100011001000000111100000110011010110111010100000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281;

XNOR2_X1 U699 ( .A(G107), .B(n966), .ZN(G9) );
NAND4_X1 U700 ( .A1(n967), .A2(n968), .A3(n969), .A4(n970), .ZN(n966) );
NOR2_X1 U701 ( .A1(n971), .A2(n972), .ZN(n969) );
XNOR2_X1 U702 ( .A(n973), .B(KEYINPUT3), .ZN(n972) );
INV_X1 U703 ( .A(n974), .ZN(n971) );
NOR2_X1 U704 ( .A1(n975), .A2(n976), .ZN(G75) );
NOR4_X1 U705 ( .A1(n977), .A2(n978), .A3(G953), .A4(n979), .ZN(n976) );
NOR4_X1 U706 ( .A1(n980), .A2(n981), .A3(n982), .A4(n983), .ZN(n978) );
NOR2_X1 U707 ( .A1(n984), .A2(n985), .ZN(n980) );
NOR2_X1 U708 ( .A1(n986), .A2(n987), .ZN(n985) );
NOR2_X1 U709 ( .A1(n988), .A2(n967), .ZN(n986) );
NOR2_X1 U710 ( .A1(n989), .A2(n990), .ZN(n988) );
NOR3_X1 U711 ( .A1(n991), .A2(n992), .A3(n993), .ZN(n984) );
NAND2_X1 U712 ( .A1(n994), .A2(n995), .ZN(n977) );
NAND2_X1 U713 ( .A1(n996), .A2(n997), .ZN(n995) );
NAND2_X1 U714 ( .A1(n998), .A2(n999), .ZN(n997) );
NAND2_X1 U715 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NAND2_X1 U716 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NAND3_X1 U717 ( .A1(n970), .A2(n1004), .A3(n1005), .ZN(n1003) );
NAND2_X1 U718 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
OR2_X1 U719 ( .A1(n1008), .A2(KEYINPUT23), .ZN(n1007) );
NAND2_X1 U720 ( .A1(n1009), .A2(n1010), .ZN(n1002) );
NAND2_X1 U721 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND2_X1 U722 ( .A1(n1005), .A2(n1013), .ZN(n1012) );
NAND2_X1 U723 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND2_X1 U724 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U725 ( .A1(n970), .A2(n1018), .ZN(n1011) );
NAND2_X1 U726 ( .A1(KEYINPUT23), .A2(n1019), .ZN(n998) );
NAND4_X1 U727 ( .A1(n1000), .A2(n1020), .A3(n1005), .A4(n970), .ZN(n1019) );
INV_X1 U728 ( .A(n983), .ZN(n1000) );
NOR3_X1 U729 ( .A1(n979), .A2(G953), .A3(G952), .ZN(n975) );
AND4_X1 U730 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n979) );
NOR4_X1 U731 ( .A1(n987), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1024) );
XNOR2_X1 U732 ( .A(n1028), .B(n1029), .ZN(n1027) );
XOR2_X1 U733 ( .A(KEYINPUT43), .B(n1030), .Z(n1026) );
NOR2_X1 U734 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
XOR2_X1 U735 ( .A(KEYINPUT54), .B(G472), .Z(n1032) );
XNOR2_X1 U736 ( .A(n1033), .B(KEYINPUT26), .ZN(n1031) );
NOR3_X1 U737 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1023) );
AND2_X1 U738 ( .A1(n1037), .A2(G472), .ZN(n1036) );
NOR2_X1 U739 ( .A1(n1038), .A2(n1039), .ZN(n1034) );
XOR2_X1 U740 ( .A(KEYINPUT50), .B(n1040), .Z(n1022) );
AND2_X1 U741 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
XOR2_X1 U742 ( .A(n1041), .B(n1042), .Z(G72) );
XOR2_X1 U743 ( .A(n1043), .B(n1044), .Z(n1042) );
NOR3_X1 U744 ( .A1(n1045), .A2(KEYINPUT20), .A3(G953), .ZN(n1044) );
INV_X1 U745 ( .A(n1046), .ZN(n1045) );
NOR3_X1 U746 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1043) );
NOR2_X1 U747 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
XNOR2_X1 U748 ( .A(n1052), .B(n1053), .ZN(n1051) );
XOR2_X1 U749 ( .A(KEYINPUT63), .B(n1054), .Z(n1047) );
NOR2_X1 U750 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XOR2_X1 U751 ( .A(KEYINPUT18), .B(n1050), .Z(n1056) );
XNOR2_X1 U752 ( .A(n1052), .B(n1057), .ZN(n1055) );
INV_X1 U753 ( .A(n1053), .ZN(n1057) );
NAND2_X1 U754 ( .A1(n1058), .A2(KEYINPUT46), .ZN(n1052) );
XNOR2_X1 U755 ( .A(n1059), .B(KEYINPUT16), .ZN(n1058) );
NOR2_X1 U756 ( .A1(n1060), .A2(n1061), .ZN(n1041) );
AND2_X1 U757 ( .A1(G227), .A2(G900), .ZN(n1060) );
XOR2_X1 U758 ( .A(n1062), .B(n1063), .Z(G69) );
NOR2_X1 U759 ( .A1(n1064), .A2(n1061), .ZN(n1063) );
NOR2_X1 U760 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND3_X1 U761 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1062) );
NAND3_X1 U762 ( .A1(n1070), .A2(n1061), .A3(n1071), .ZN(n1069) );
NAND2_X1 U763 ( .A1(KEYINPUT51), .A2(n1072), .ZN(n1071) );
NAND2_X1 U764 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
OR2_X1 U765 ( .A1(n1075), .A2(KEYINPUT51), .ZN(n1068) );
NAND3_X1 U766 ( .A1(n1075), .A2(n1076), .A3(KEYINPUT51), .ZN(n1067) );
NAND3_X1 U767 ( .A1(n1070), .A2(n1061), .A3(n1073), .ZN(n1076) );
XOR2_X1 U768 ( .A(KEYINPUT53), .B(KEYINPUT39), .Z(n1073) );
INV_X1 U769 ( .A(n1074), .ZN(n1075) );
NAND2_X1 U770 ( .A1(n1077), .A2(n1078), .ZN(n1074) );
NAND2_X1 U771 ( .A1(G953), .A2(n1066), .ZN(n1078) );
XOR2_X1 U772 ( .A(n1079), .B(n1080), .Z(n1077) );
XOR2_X1 U773 ( .A(n1081), .B(KEYINPUT34), .Z(n1079) );
NOR2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(G66) );
XOR2_X1 U775 ( .A(n1084), .B(n1085), .Z(n1083) );
NAND2_X1 U776 ( .A1(n1086), .A2(n1038), .ZN(n1084) );
INV_X1 U777 ( .A(n1087), .ZN(n1038) );
NOR2_X1 U778 ( .A1(n1082), .A2(n1088), .ZN(G63) );
XOR2_X1 U779 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U780 ( .A1(KEYINPUT33), .A2(n1091), .ZN(n1090) );
XOR2_X1 U781 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND2_X1 U782 ( .A1(n1086), .A2(G478), .ZN(n1089) );
NOR2_X1 U783 ( .A1(n1082), .A2(n1094), .ZN(G60) );
XOR2_X1 U784 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND2_X1 U785 ( .A1(n1086), .A2(G475), .ZN(n1095) );
XNOR2_X1 U786 ( .A(n1097), .B(n1098), .ZN(G6) );
NOR2_X1 U787 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NOR2_X1 U788 ( .A1(n1082), .A2(n1101), .ZN(G57) );
XOR2_X1 U789 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U790 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U791 ( .A1(n1086), .A2(G472), .ZN(n1105) );
NAND2_X1 U792 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NAND2_X1 U793 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
XNOR2_X1 U794 ( .A(G101), .B(KEYINPUT24), .ZN(n1108) );
XOR2_X1 U795 ( .A(n1110), .B(n1111), .Z(n1102) );
NOR2_X1 U796 ( .A1(n1082), .A2(n1112), .ZN(G54) );
XOR2_X1 U797 ( .A(n1113), .B(n1114), .Z(n1112) );
AND2_X1 U798 ( .A1(G469), .A2(n1086), .ZN(n1114) );
NAND2_X1 U799 ( .A1(n1115), .A2(KEYINPUT55), .ZN(n1113) );
XOR2_X1 U800 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U801 ( .A1(G110), .A2(KEYINPUT58), .ZN(n1117) );
NOR2_X1 U802 ( .A1(n1061), .A2(G952), .ZN(n1082) );
NOR2_X1 U803 ( .A1(n1118), .A2(n1119), .ZN(G51) );
XOR2_X1 U804 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U805 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR3_X1 U806 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
INV_X1 U807 ( .A(KEYINPUT35), .ZN(n1124) );
NOR2_X1 U808 ( .A1(KEYINPUT35), .A2(n1127), .ZN(n1122) );
NAND2_X1 U809 ( .A1(n1086), .A2(n1029), .ZN(n1120) );
NOR2_X1 U810 ( .A1(n1128), .A2(n994), .ZN(n1086) );
NOR2_X1 U811 ( .A1(n1046), .A2(n1070), .ZN(n994) );
NAND4_X1 U812 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1070) );
AND3_X1 U813 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
NAND2_X1 U814 ( .A1(n967), .A2(n1136), .ZN(n1131) );
NAND3_X1 U815 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
XNOR2_X1 U816 ( .A(KEYINPUT7), .B(n1100), .ZN(n1139) );
NAND4_X1 U817 ( .A1(n1020), .A2(n970), .A3(n974), .A4(n1140), .ZN(n1100) );
NAND4_X1 U818 ( .A1(n968), .A2(n970), .A3(n974), .A4(n1140), .ZN(n1138) );
XOR2_X1 U819 ( .A(KEYINPUT38), .B(n1141), .Z(n1137) );
NAND2_X1 U820 ( .A1(n1142), .A2(n1143), .ZN(n1046) );
NOR4_X1 U821 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1143) );
NOR4_X1 U822 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1142) );
NOR3_X1 U823 ( .A1(n992), .A2(n1008), .A3(n1152), .ZN(n1151) );
INV_X1 U824 ( .A(n1153), .ZN(n1148) );
NOR2_X1 U825 ( .A1(G952), .A2(n1154), .ZN(n1118) );
XNOR2_X1 U826 ( .A(KEYINPUT29), .B(n1061), .ZN(n1154) );
XOR2_X1 U827 ( .A(n1147), .B(n1155), .Z(G48) );
NOR2_X1 U828 ( .A1(KEYINPUT19), .A2(n1156), .ZN(n1155) );
INV_X1 U829 ( .A(G146), .ZN(n1156) );
AND4_X1 U830 ( .A1(n1157), .A2(n1158), .A3(n1020), .A4(n1018), .ZN(n1147) );
XNOR2_X1 U831 ( .A(n1159), .B(n1150), .ZN(G45) );
NOR2_X1 U832 ( .A1(n1160), .A2(n1152), .ZN(n1150) );
XOR2_X1 U833 ( .A(G140), .B(n1149), .Z(G42) );
AND3_X1 U834 ( .A1(n1020), .A2(n1017), .A3(n1161), .ZN(n1149) );
XOR2_X1 U835 ( .A(G137), .B(n1146), .Z(G39) );
AND3_X1 U836 ( .A1(n1157), .A2(n1161), .A3(n1009), .ZN(n1146) );
AND4_X1 U837 ( .A1(n1016), .A2(n996), .A3(n1018), .A4(n1162), .ZN(n1161) );
XOR2_X1 U838 ( .A(G134), .B(n1145), .Z(G36) );
NOR3_X1 U839 ( .A1(n1152), .A2(n1006), .A3(n992), .ZN(n1145) );
INV_X1 U840 ( .A(n996), .ZN(n992) );
XNOR2_X1 U841 ( .A(n1163), .B(n1164), .ZN(G33) );
NOR3_X1 U842 ( .A1(n1152), .A2(n1165), .A3(n1008), .ZN(n1164) );
INV_X1 U843 ( .A(n1020), .ZN(n1008) );
XNOR2_X1 U844 ( .A(n996), .B(KEYINPUT12), .ZN(n1165) );
NOR2_X1 U845 ( .A1(n989), .A2(n1035), .ZN(n996) );
INV_X1 U846 ( .A(n1166), .ZN(n989) );
NAND3_X1 U847 ( .A1(n1018), .A2(n1162), .A3(n1167), .ZN(n1152) );
XOR2_X1 U848 ( .A(n1168), .B(G128), .Z(G30) );
NAND2_X1 U849 ( .A1(KEYINPUT47), .A2(n1153), .ZN(n1168) );
NAND4_X1 U850 ( .A1(n1157), .A2(n1158), .A3(n968), .A4(n974), .ZN(n1153) );
XNOR2_X1 U851 ( .A(G101), .B(n1129), .ZN(G3) );
NAND3_X1 U852 ( .A1(n1167), .A2(n974), .A3(n1169), .ZN(n1129) );
XNOR2_X1 U853 ( .A(n1144), .B(n1170), .ZN(G27) );
NAND2_X1 U854 ( .A1(KEYINPUT28), .A2(G125), .ZN(n1170) );
AND4_X1 U855 ( .A1(n1158), .A2(n1020), .A3(n1005), .A4(n1017), .ZN(n1144) );
AND3_X1 U856 ( .A1(n967), .A2(n1162), .A3(n1016), .ZN(n1158) );
NAND2_X1 U857 ( .A1(n1171), .A2(n983), .ZN(n1162) );
XOR2_X1 U858 ( .A(n1172), .B(KEYINPUT4), .Z(n1171) );
NAND3_X1 U859 ( .A1(G902), .A2(n1173), .A3(n1048), .ZN(n1172) );
AND2_X1 U860 ( .A1(G953), .A2(n1174), .ZN(n1048) );
XOR2_X1 U861 ( .A(KEYINPUT31), .B(G900), .Z(n1174) );
XNOR2_X1 U862 ( .A(n1130), .B(n1175), .ZN(G24) );
NOR2_X1 U863 ( .A1(KEYINPUT48), .A2(n1176), .ZN(n1175) );
OR4_X1 U864 ( .A1(n1160), .A2(n987), .A3(n981), .A4(n973), .ZN(n1130) );
INV_X1 U865 ( .A(n970), .ZN(n981) );
NOR2_X1 U866 ( .A1(n1157), .A2(n1016), .ZN(n970) );
NAND3_X1 U867 ( .A1(n1025), .A2(n1177), .A3(n967), .ZN(n1160) );
XNOR2_X1 U868 ( .A(n1178), .B(n1179), .ZN(G21) );
NOR2_X1 U869 ( .A1(KEYINPUT45), .A2(n1133), .ZN(n1179) );
NAND4_X1 U870 ( .A1(n1157), .A2(n1169), .A3(n1016), .A4(n1005), .ZN(n1133) );
INV_X1 U871 ( .A(n1017), .ZN(n1157) );
XOR2_X1 U872 ( .A(n1180), .B(G116), .Z(G18) );
NAND2_X1 U873 ( .A1(KEYINPUT21), .A2(n1181), .ZN(n1180) );
NAND2_X1 U874 ( .A1(n1141), .A2(n967), .ZN(n1181) );
NOR4_X1 U875 ( .A1(n1014), .A2(n987), .A3(n1006), .A4(n973), .ZN(n1141) );
INV_X1 U876 ( .A(n968), .ZN(n1006) );
NOR2_X1 U877 ( .A1(n1177), .A2(n1182), .ZN(n968) );
INV_X1 U878 ( .A(n1025), .ZN(n1182) );
INV_X1 U879 ( .A(n1167), .ZN(n1014) );
XOR2_X1 U880 ( .A(n1135), .B(n1183), .Z(G15) );
XNOR2_X1 U881 ( .A(G113), .B(KEYINPUT10), .ZN(n1183) );
NAND4_X1 U882 ( .A1(n1167), .A2(n1020), .A3(n1184), .A4(n1005), .ZN(n1135) );
INV_X1 U883 ( .A(n987), .ZN(n1005) );
NAND2_X1 U884 ( .A1(n1185), .A2(n991), .ZN(n987) );
INV_X1 U885 ( .A(n993), .ZN(n1185) );
NOR2_X1 U886 ( .A1(n973), .A2(n1099), .ZN(n1184) );
NOR2_X1 U887 ( .A1(n1025), .A2(n1186), .ZN(n1020) );
INV_X1 U888 ( .A(n1177), .ZN(n1186) );
NOR2_X1 U889 ( .A1(n1017), .A2(n1016), .ZN(n1167) );
XNOR2_X1 U890 ( .A(G110), .B(n1134), .ZN(G12) );
NAND4_X1 U891 ( .A1(n1016), .A2(n1169), .A3(n974), .A4(n1017), .ZN(n1134) );
XNOR2_X1 U892 ( .A(n1187), .B(n1188), .ZN(n1017) );
NOR2_X1 U893 ( .A1(KEYINPUT11), .A2(n1033), .ZN(n1188) );
INV_X1 U894 ( .A(n1037), .ZN(n1033) );
NAND2_X1 U895 ( .A1(n1189), .A2(n1190), .ZN(n1037) );
XOR2_X1 U896 ( .A(n1191), .B(n1192), .Z(n1189) );
XNOR2_X1 U897 ( .A(n1053), .B(n1111), .ZN(n1192) );
XNOR2_X1 U898 ( .A(n1193), .B(n1194), .ZN(n1111) );
XNOR2_X1 U899 ( .A(n1178), .B(G116), .ZN(n1194) );
XOR2_X1 U900 ( .A(n1195), .B(n1196), .Z(n1191) );
NOR2_X1 U901 ( .A1(KEYINPUT36), .A2(n1059), .ZN(n1196) );
XOR2_X1 U902 ( .A(n1197), .B(KEYINPUT5), .Z(n1195) );
NAND2_X1 U903 ( .A1(n1107), .A2(n1198), .ZN(n1197) );
NAND2_X1 U904 ( .A1(n1109), .A2(n1199), .ZN(n1198) );
NAND2_X1 U905 ( .A1(n1200), .A2(G210), .ZN(n1109) );
NAND3_X1 U906 ( .A1(G210), .A2(G101), .A3(n1200), .ZN(n1107) );
XNOR2_X1 U907 ( .A(G472), .B(KEYINPUT56), .ZN(n1187) );
XOR2_X1 U908 ( .A(n1018), .B(KEYINPUT6), .Z(n974) );
AND2_X1 U909 ( .A1(n993), .A2(n991), .ZN(n1018) );
NAND2_X1 U910 ( .A1(G221), .A2(n1201), .ZN(n991) );
XNOR2_X1 U911 ( .A(n1202), .B(G469), .ZN(n993) );
NAND2_X1 U912 ( .A1(n1203), .A2(n1190), .ZN(n1202) );
XOR2_X1 U913 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U914 ( .A(KEYINPUT42), .B(KEYINPUT40), .Z(n1205) );
XOR2_X1 U915 ( .A(n1116), .B(G110), .Z(n1204) );
XOR2_X1 U916 ( .A(n1206), .B(n1207), .Z(n1116) );
XOR2_X1 U917 ( .A(n1110), .B(n1208), .Z(n1207) );
XNOR2_X1 U918 ( .A(n1209), .B(n1210), .ZN(n1208) );
NAND2_X1 U919 ( .A1(G227), .A2(n1061), .ZN(n1209) );
XNOR2_X1 U920 ( .A(n1053), .B(n1059), .ZN(n1110) );
XNOR2_X1 U921 ( .A(n1211), .B(n1212), .ZN(n1053) );
XOR2_X1 U922 ( .A(KEYINPUT62), .B(G137), .Z(n1212) );
XNOR2_X1 U923 ( .A(G131), .B(n1213), .ZN(n1211) );
XNOR2_X1 U924 ( .A(G101), .B(n1214), .ZN(n1206) );
XOR2_X1 U925 ( .A(KEYINPUT16), .B(G140), .Z(n1214) );
NOR3_X1 U926 ( .A1(n1099), .A2(n973), .A3(n982), .ZN(n1169) );
INV_X1 U927 ( .A(n1009), .ZN(n982) );
NOR2_X1 U928 ( .A1(n1025), .A2(n1177), .ZN(n1009) );
XNOR2_X1 U929 ( .A(n1021), .B(KEYINPUT52), .ZN(n1177) );
XOR2_X1 U930 ( .A(n1215), .B(G475), .Z(n1021) );
NAND2_X1 U931 ( .A1(n1096), .A2(n1190), .ZN(n1215) );
XNOR2_X1 U932 ( .A(n1216), .B(n1217), .ZN(n1096) );
XOR2_X1 U933 ( .A(n1218), .B(n1050), .Z(n1217) );
XOR2_X1 U934 ( .A(n1219), .B(n1220), .Z(n1216) );
AND2_X1 U935 ( .A1(G214), .A2(n1200), .ZN(n1220) );
NOR2_X1 U936 ( .A1(G953), .A2(G237), .ZN(n1200) );
XNOR2_X1 U937 ( .A(n1221), .B(n1163), .ZN(n1219) );
INV_X1 U938 ( .A(G131), .ZN(n1163) );
NAND3_X1 U939 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1221) );
NAND2_X1 U940 ( .A1(n1225), .A2(n1097), .ZN(n1224) );
NAND2_X1 U941 ( .A1(KEYINPUT57), .A2(n1226), .ZN(n1223) );
NAND2_X1 U942 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
XNOR2_X1 U943 ( .A(KEYINPUT9), .B(n1097), .ZN(n1227) );
NAND2_X1 U944 ( .A1(n1229), .A2(n1230), .ZN(n1222) );
INV_X1 U945 ( .A(KEYINPUT57), .ZN(n1230) );
NAND2_X1 U946 ( .A1(n1231), .A2(n1232), .ZN(n1229) );
NAND2_X1 U947 ( .A1(KEYINPUT9), .A2(n1097), .ZN(n1232) );
OR3_X1 U948 ( .A1(n1225), .A2(KEYINPUT9), .A3(n1097), .ZN(n1231) );
INV_X1 U949 ( .A(n1228), .ZN(n1225) );
XNOR2_X1 U950 ( .A(G113), .B(n1176), .ZN(n1228) );
XNOR2_X1 U951 ( .A(n1233), .B(G478), .ZN(n1025) );
NAND2_X1 U952 ( .A1(n1234), .A2(n1190), .ZN(n1233) );
XNOR2_X1 U953 ( .A(n1092), .B(n1093), .ZN(n1234) );
XNOR2_X1 U954 ( .A(n1235), .B(n1236), .ZN(n1093) );
XNOR2_X1 U955 ( .A(G128), .B(n1176), .ZN(n1236) );
XNOR2_X1 U956 ( .A(G143), .B(KEYINPUT2), .ZN(n1235) );
XOR2_X1 U957 ( .A(n1237), .B(n1238), .Z(n1092) );
XOR2_X1 U958 ( .A(G116), .B(G107), .Z(n1238) );
XOR2_X1 U959 ( .A(n1239), .B(n1213), .Z(n1237) );
XOR2_X1 U960 ( .A(G134), .B(KEYINPUT27), .Z(n1213) );
NAND2_X1 U961 ( .A1(G217), .A2(n1240), .ZN(n1239) );
INV_X1 U962 ( .A(n1140), .ZN(n973) );
NAND2_X1 U963 ( .A1(n983), .A2(n1241), .ZN(n1140) );
NAND4_X1 U964 ( .A1(G953), .A2(G902), .A3(n1173), .A4(n1066), .ZN(n1241) );
INV_X1 U965 ( .A(G898), .ZN(n1066) );
NAND3_X1 U966 ( .A1(n1173), .A2(n1061), .A3(G952), .ZN(n983) );
NAND2_X1 U967 ( .A1(G237), .A2(n1242), .ZN(n1173) );
XOR2_X1 U968 ( .A(KEYINPUT25), .B(G234), .Z(n1242) );
INV_X1 U969 ( .A(n967), .ZN(n1099) );
NOR2_X1 U970 ( .A1(n1166), .A2(n1035), .ZN(n967) );
INV_X1 U971 ( .A(n990), .ZN(n1035) );
NAND2_X1 U972 ( .A1(G214), .A2(n1243), .ZN(n990) );
NAND3_X1 U973 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1166) );
OR2_X1 U974 ( .A1(n1247), .A2(KEYINPUT37), .ZN(n1246) );
NAND3_X1 U975 ( .A1(KEYINPUT37), .A2(n1248), .A3(n1028), .ZN(n1245) );
OR2_X1 U976 ( .A1(n1028), .A2(n1248), .ZN(n1244) );
NOR2_X1 U977 ( .A1(n1029), .A2(KEYINPUT22), .ZN(n1248) );
INV_X1 U978 ( .A(n1247), .ZN(n1029) );
NAND2_X1 U979 ( .A1(G210), .A2(n1243), .ZN(n1247) );
NAND2_X1 U980 ( .A1(n1249), .A2(n1128), .ZN(n1243) );
INV_X1 U981 ( .A(G237), .ZN(n1249) );
NAND2_X1 U982 ( .A1(n1127), .A2(n1190), .ZN(n1028) );
XNOR2_X1 U983 ( .A(n1125), .B(n1126), .ZN(n1127) );
XOR2_X1 U984 ( .A(n1081), .B(n1250), .Z(n1126) );
NOR2_X1 U985 ( .A1(KEYINPUT15), .A2(n1251), .ZN(n1250) );
XOR2_X1 U986 ( .A(KEYINPUT1), .B(n1080), .Z(n1251) );
XNOR2_X1 U987 ( .A(n1193), .B(n1252), .ZN(n1080) );
NOR2_X1 U988 ( .A1(KEYINPUT32), .A2(n1253), .ZN(n1252) );
XNOR2_X1 U989 ( .A(n1178), .B(n1254), .ZN(n1253) );
NOR2_X1 U990 ( .A1(G116), .A2(KEYINPUT60), .ZN(n1254) );
INV_X1 U991 ( .A(G119), .ZN(n1178) );
INV_X1 U992 ( .A(G113), .ZN(n1193) );
XOR2_X1 U993 ( .A(n1255), .B(n1256), .Z(n1081) );
XNOR2_X1 U994 ( .A(KEYINPUT13), .B(n1176), .ZN(n1256) );
INV_X1 U995 ( .A(G122), .ZN(n1176) );
XOR2_X1 U996 ( .A(n1257), .B(G110), .Z(n1255) );
NAND3_X1 U997 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1257) );
NAND2_X1 U998 ( .A1(KEYINPUT14), .A2(n1261), .ZN(n1260) );
NAND3_X1 U999 ( .A1(n1262), .A2(n1263), .A3(n1199), .ZN(n1259) );
INV_X1 U1000 ( .A(KEYINPUT14), .ZN(n1263) );
OR2_X1 U1001 ( .A1(n1199), .A2(n1262), .ZN(n1258) );
NOR2_X1 U1002 ( .A1(n1264), .A2(n1261), .ZN(n1262) );
NAND2_X1 U1003 ( .A1(n1265), .A2(n1266), .ZN(n1261) );
NAND2_X1 U1004 ( .A1(KEYINPUT44), .A2(n1210), .ZN(n1266) );
XNOR2_X1 U1005 ( .A(G107), .B(G104), .ZN(n1210) );
OR3_X1 U1006 ( .A1(n1097), .A2(G107), .A3(KEYINPUT44), .ZN(n1265) );
INV_X1 U1007 ( .A(G104), .ZN(n1097) );
INV_X1 U1008 ( .A(KEYINPUT49), .ZN(n1264) );
INV_X1 U1009 ( .A(G101), .ZN(n1199) );
XNOR2_X1 U1010 ( .A(n1267), .B(n1268), .ZN(n1125) );
INV_X1 U1011 ( .A(n1059), .ZN(n1268) );
XOR2_X1 U1012 ( .A(G128), .B(n1218), .Z(n1059) );
XNOR2_X1 U1013 ( .A(n1159), .B(G146), .ZN(n1218) );
INV_X1 U1014 ( .A(G143), .ZN(n1159) );
XNOR2_X1 U1015 ( .A(G125), .B(n1269), .ZN(n1267) );
NOR2_X1 U1016 ( .A1(G953), .A2(n1065), .ZN(n1269) );
INV_X1 U1017 ( .A(G224), .ZN(n1065) );
XNOR2_X1 U1018 ( .A(n1270), .B(n1039), .ZN(n1016) );
NAND2_X1 U1019 ( .A1(n1271), .A2(n1190), .ZN(n1039) );
XNOR2_X1 U1020 ( .A(n1128), .B(KEYINPUT30), .ZN(n1190) );
XOR2_X1 U1021 ( .A(n1085), .B(KEYINPUT0), .Z(n1271) );
XOR2_X1 U1022 ( .A(n1272), .B(n1273), .Z(n1085) );
AND2_X1 U1023 ( .A1(n1240), .A2(G221), .ZN(n1273) );
AND2_X1 U1024 ( .A1(G234), .A2(n1061), .ZN(n1240) );
INV_X1 U1025 ( .A(G953), .ZN(n1061) );
XOR2_X1 U1026 ( .A(n1274), .B(G137), .Z(n1272) );
NAND2_X1 U1027 ( .A1(n1275), .A2(KEYINPUT17), .ZN(n1274) );
XOR2_X1 U1028 ( .A(n1276), .B(n1277), .Z(n1275) );
NOR2_X1 U1029 ( .A1(KEYINPUT59), .A2(n1278), .ZN(n1277) );
XNOR2_X1 U1030 ( .A(G146), .B(n1050), .ZN(n1278) );
XOR2_X1 U1031 ( .A(G125), .B(G140), .Z(n1050) );
XNOR2_X1 U1032 ( .A(G110), .B(n1279), .ZN(n1276) );
NOR2_X1 U1033 ( .A1(KEYINPUT61), .A2(n1280), .ZN(n1279) );
XNOR2_X1 U1034 ( .A(G119), .B(n1281), .ZN(n1280) );
XOR2_X1 U1035 ( .A(KEYINPUT8), .B(G128), .Z(n1281) );
NAND2_X1 U1036 ( .A1(KEYINPUT41), .A2(n1087), .ZN(n1270) );
NAND2_X1 U1037 ( .A1(G217), .A2(n1201), .ZN(n1087) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1128), .ZN(n1201) );
INV_X1 U1039 ( .A(G902), .ZN(n1128) );
endmodule


