//Key = 1110100011000010011101000110001011101001010011111110010101100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396;

XOR2_X1 U759 ( .A(n1057), .B(n1058), .Z(G9) );
NAND2_X1 U760 ( .A1(KEYINPUT17), .A2(G107), .ZN(n1058) );
NAND3_X1 U761 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1057) );
XNOR2_X1 U762 ( .A(KEYINPUT3), .B(n1062), .ZN(n1060) );
NOR2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(G75) );
NOR4_X1 U764 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1064) );
NOR2_X1 U765 ( .A1(KEYINPUT1), .A2(n1069), .ZN(n1067) );
NOR4_X1 U766 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1062), .ZN(n1069) );
NAND2_X1 U767 ( .A1(n1073), .A2(n1074), .ZN(n1070) );
XNOR2_X1 U768 ( .A(KEYINPUT47), .B(n1075), .ZN(n1066) );
NAND4_X1 U769 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1065) );
NAND4_X1 U770 ( .A1(n1073), .A2(n1074), .A3(n1080), .A4(n1081), .ZN(n1077) );
NAND3_X1 U771 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NAND2_X1 U772 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U773 ( .A1(n1087), .A2(n1088), .ZN(n1083) );
NAND2_X1 U774 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U775 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XNOR2_X1 U776 ( .A(n1093), .B(KEYINPUT6), .ZN(n1091) );
NAND2_X1 U777 ( .A1(KEYINPUT1), .A2(n1094), .ZN(n1089) );
NAND2_X1 U778 ( .A1(n1095), .A2(n1096), .ZN(n1082) );
XOR2_X1 U779 ( .A(KEYINPUT28), .B(n1085), .Z(n1096) );
NAND2_X1 U780 ( .A1(n1085), .A2(n1097), .ZN(n1076) );
NAND2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND3_X1 U782 ( .A1(n1087), .A2(n1100), .A3(n1073), .ZN(n1099) );
INV_X1 U783 ( .A(n1101), .ZN(n1073) );
NAND2_X1 U784 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NAND3_X1 U785 ( .A1(n1104), .A2(n1105), .A3(n1074), .ZN(n1103) );
NAND2_X1 U786 ( .A1(n1080), .A2(n1106), .ZN(n1102) );
OR2_X1 U787 ( .A1(n1107), .A2(n1059), .ZN(n1106) );
XOR2_X1 U788 ( .A(n1108), .B(KEYINPUT43), .Z(n1098) );
NAND4_X1 U789 ( .A1(n1109), .A2(n1087), .A3(n1074), .A4(n1110), .ZN(n1108) );
NOR2_X1 U790 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XNOR2_X1 U791 ( .A(KEYINPUT32), .B(n1105), .ZN(n1112) );
XNOR2_X1 U792 ( .A(KEYINPUT48), .B(n1101), .ZN(n1111) );
NOR3_X1 U793 ( .A1(n1113), .A2(G953), .A3(G952), .ZN(n1063) );
INV_X1 U794 ( .A(n1078), .ZN(n1113) );
NAND4_X1 U795 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1078) );
NOR4_X1 U796 ( .A1(n1118), .A2(n1092), .A3(n1119), .A4(n1120), .ZN(n1117) );
NOR2_X1 U797 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
NOR2_X1 U798 ( .A1(n1123), .A2(G902), .ZN(n1121) );
NOR2_X1 U799 ( .A1(n1071), .A2(n1124), .ZN(n1116) );
XOR2_X1 U800 ( .A(n1125), .B(n1126), .Z(n1124) );
XNOR2_X1 U801 ( .A(KEYINPUT58), .B(n1127), .ZN(n1126) );
NOR2_X1 U802 ( .A1(KEYINPUT52), .A2(n1128), .ZN(n1127) );
INV_X1 U803 ( .A(n1129), .ZN(n1128) );
XNOR2_X1 U804 ( .A(n1130), .B(KEYINPUT42), .ZN(n1115) );
XOR2_X1 U805 ( .A(n1131), .B(n1132), .Z(n1114) );
XOR2_X1 U806 ( .A(n1133), .B(n1134), .Z(G72) );
XOR2_X1 U807 ( .A(n1135), .B(n1136), .Z(n1134) );
NAND2_X1 U808 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U809 ( .A1(G953), .A2(n1139), .ZN(n1138) );
XOR2_X1 U810 ( .A(n1140), .B(n1141), .Z(n1137) );
XNOR2_X1 U811 ( .A(G140), .B(n1142), .ZN(n1141) );
XNOR2_X1 U812 ( .A(KEYINPUT63), .B(KEYINPUT27), .ZN(n1142) );
XOR2_X1 U813 ( .A(n1143), .B(n1144), .Z(n1140) );
XNOR2_X1 U814 ( .A(G125), .B(n1145), .ZN(n1143) );
NAND2_X1 U815 ( .A1(n1146), .A2(n1147), .ZN(n1135) );
NAND2_X1 U816 ( .A1(G900), .A2(G227), .ZN(n1147) );
XNOR2_X1 U817 ( .A(KEYINPUT23), .B(n1079), .ZN(n1146) );
NOR2_X1 U818 ( .A1(n1148), .A2(G953), .ZN(n1133) );
NAND3_X1 U819 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(G69) );
NAND3_X1 U820 ( .A1(n1152), .A2(n1153), .A3(G953), .ZN(n1151) );
NAND3_X1 U821 ( .A1(G898), .A2(G224), .A3(KEYINPUT2), .ZN(n1152) );
NAND2_X1 U822 ( .A1(n1154), .A2(n1155), .ZN(n1150) );
INV_X1 U823 ( .A(KEYINPUT2), .ZN(n1155) );
NAND2_X1 U824 ( .A1(n1156), .A2(n1157), .ZN(n1154) );
NAND2_X1 U825 ( .A1(n1158), .A2(n1153), .ZN(n1157) );
NAND3_X1 U826 ( .A1(n1075), .A2(n1079), .A3(n1159), .ZN(n1156) );
NAND2_X1 U827 ( .A1(n1160), .A2(KEYINPUT2), .ZN(n1149) );
NAND2_X1 U828 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U829 ( .A1(n1163), .A2(n1079), .ZN(n1162) );
XNOR2_X1 U830 ( .A(n1158), .B(n1159), .ZN(n1163) );
NAND3_X1 U831 ( .A1(n1159), .A2(G224), .A3(G953), .ZN(n1161) );
INV_X1 U832 ( .A(n1153), .ZN(n1159) );
NAND3_X1 U833 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1153) );
XOR2_X1 U834 ( .A(n1167), .B(KEYINPUT10), .Z(n1166) );
NAND2_X1 U835 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
OR2_X1 U836 ( .A1(n1168), .A2(n1169), .ZN(n1165) );
XOR2_X1 U837 ( .A(n1170), .B(n1171), .Z(n1168) );
OR2_X1 U838 ( .A1(n1079), .A2(G898), .ZN(n1164) );
NOR2_X1 U839 ( .A1(n1172), .A2(n1173), .ZN(G66) );
NOR3_X1 U840 ( .A1(n1174), .A2(n1131), .A3(n1175), .ZN(n1173) );
NOR2_X1 U841 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NOR2_X1 U842 ( .A1(n1178), .A2(n1132), .ZN(n1176) );
NOR2_X1 U843 ( .A1(n1075), .A2(n1068), .ZN(n1178) );
XOR2_X1 U844 ( .A(KEYINPUT40), .B(n1179), .Z(n1174) );
NOR3_X1 U845 ( .A1(n1180), .A2(n1181), .A3(n1132), .ZN(n1179) );
NOR2_X1 U846 ( .A1(n1172), .A2(n1182), .ZN(G63) );
XNOR2_X1 U847 ( .A(n1183), .B(n1184), .ZN(n1182) );
NOR2_X1 U848 ( .A1(n1185), .A2(n1180), .ZN(n1184) );
NOR2_X1 U849 ( .A1(n1172), .A2(n1186), .ZN(G60) );
NOR2_X1 U850 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U851 ( .A(KEYINPUT29), .B(n1189), .Z(n1188) );
AND2_X1 U852 ( .A1(n1190), .A2(n1123), .ZN(n1189) );
NOR2_X1 U853 ( .A1(n1123), .A2(n1190), .ZN(n1187) );
NOR2_X1 U854 ( .A1(n1180), .A2(n1122), .ZN(n1190) );
INV_X1 U855 ( .A(G475), .ZN(n1122) );
XNOR2_X1 U856 ( .A(n1191), .B(n1192), .ZN(G6) );
NOR2_X1 U857 ( .A1(n1172), .A2(n1193), .ZN(G57) );
XOR2_X1 U858 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U859 ( .A(n1196), .B(n1197), .Z(n1195) );
XOR2_X1 U860 ( .A(n1198), .B(n1199), .Z(n1194) );
XOR2_X1 U861 ( .A(KEYINPUT15), .B(n1200), .Z(n1199) );
NOR2_X1 U862 ( .A1(n1201), .A2(n1180), .ZN(n1198) );
NOR2_X1 U863 ( .A1(n1172), .A2(n1202), .ZN(G54) );
XOR2_X1 U864 ( .A(n1203), .B(n1204), .Z(n1202) );
XOR2_X1 U865 ( .A(n1205), .B(n1144), .Z(n1204) );
XOR2_X1 U866 ( .A(n1206), .B(n1207), .Z(n1203) );
NOR2_X1 U867 ( .A1(n1208), .A2(n1180), .ZN(n1206) );
NOR2_X1 U868 ( .A1(n1172), .A2(n1209), .ZN(G51) );
XOR2_X1 U869 ( .A(n1210), .B(n1211), .Z(n1209) );
NOR2_X1 U870 ( .A1(n1129), .A2(n1180), .ZN(n1211) );
NAND2_X1 U871 ( .A1(G902), .A2(n1212), .ZN(n1180) );
NAND2_X1 U872 ( .A1(n1148), .A2(n1158), .ZN(n1212) );
INV_X1 U873 ( .A(n1075), .ZN(n1158) );
NAND4_X1 U874 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1075) );
NOR4_X1 U875 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1216) );
NOR2_X1 U876 ( .A1(n1192), .A2(n1221), .ZN(n1215) );
AND4_X1 U877 ( .A1(n1222), .A2(n1080), .A3(n1223), .A4(n1074), .ZN(n1221) );
AND3_X1 U878 ( .A1(n1061), .A2(n1087), .A3(n1107), .ZN(n1192) );
NAND3_X1 U879 ( .A1(n1059), .A2(n1087), .A3(n1061), .ZN(n1214) );
NAND2_X1 U880 ( .A1(n1224), .A2(n1094), .ZN(n1213) );
INV_X1 U881 ( .A(n1068), .ZN(n1148) );
NAND4_X1 U882 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1068) );
NOR4_X1 U883 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1228) );
INV_X1 U884 ( .A(n1233), .ZN(n1231) );
INV_X1 U885 ( .A(n1234), .ZN(n1230) );
NOR3_X1 U886 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1227) );
NOR2_X1 U887 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
INV_X1 U888 ( .A(KEYINPUT36), .ZN(n1238) );
NOR4_X1 U889 ( .A1(KEYINPUT36), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1236) );
NAND3_X1 U890 ( .A1(n1243), .A2(n1072), .A3(n1244), .ZN(n1240) );
INV_X1 U891 ( .A(n1245), .ZN(n1235) );
NAND2_X1 U892 ( .A1(KEYINPUT44), .A2(n1246), .ZN(n1210) );
XOR2_X1 U893 ( .A(n1247), .B(n1248), .Z(n1246) );
XNOR2_X1 U894 ( .A(n1249), .B(n1250), .ZN(n1248) );
XOR2_X1 U895 ( .A(n1251), .B(KEYINPUT50), .Z(n1247) );
NOR2_X1 U896 ( .A1(n1079), .A2(G952), .ZN(n1172) );
XNOR2_X1 U897 ( .A(G146), .B(n1239), .ZN(G48) );
NAND3_X1 U898 ( .A1(n1107), .A2(n1252), .A3(n1223), .ZN(n1239) );
XNOR2_X1 U899 ( .A(G143), .B(n1245), .ZN(G45) );
NAND4_X1 U900 ( .A1(n1253), .A2(n1094), .A3(n1130), .A4(n1254), .ZN(n1245) );
XOR2_X1 U901 ( .A(G140), .B(n1229), .Z(G42) );
AND4_X1 U902 ( .A1(n1085), .A2(n1086), .A3(n1107), .A4(n1252), .ZN(n1229) );
XOR2_X1 U903 ( .A(n1225), .B(n1255), .Z(G39) );
XNOR2_X1 U904 ( .A(G137), .B(KEYINPUT60), .ZN(n1255) );
NAND3_X1 U905 ( .A1(n1074), .A2(n1085), .A3(n1256), .ZN(n1225) );
NOR3_X1 U906 ( .A1(n1241), .A2(n1257), .A3(n1258), .ZN(n1256) );
INV_X1 U907 ( .A(n1252), .ZN(n1241) );
XNOR2_X1 U908 ( .A(G134), .B(n1226), .ZN(G36) );
NAND3_X1 U909 ( .A1(n1085), .A2(n1059), .A3(n1253), .ZN(n1226) );
XNOR2_X1 U910 ( .A(G131), .B(n1259), .ZN(G33) );
NOR2_X1 U911 ( .A1(n1232), .A2(KEYINPUT22), .ZN(n1259) );
AND3_X1 U912 ( .A1(n1085), .A2(n1107), .A3(n1253), .ZN(n1232) );
AND2_X1 U913 ( .A1(n1095), .A2(n1252), .ZN(n1253) );
NOR2_X1 U914 ( .A1(n1093), .A2(n1092), .ZN(n1085) );
XOR2_X1 U915 ( .A(n1260), .B(n1261), .Z(G30) );
XNOR2_X1 U916 ( .A(G128), .B(KEYINPUT49), .ZN(n1261) );
NAND2_X1 U917 ( .A1(KEYINPUT19), .A2(n1234), .ZN(n1260) );
NAND3_X1 U918 ( .A1(n1252), .A2(n1059), .A3(n1223), .ZN(n1234) );
NOR3_X1 U919 ( .A1(n1262), .A2(n1263), .A3(n1109), .ZN(n1252) );
INV_X1 U920 ( .A(n1104), .ZN(n1109) );
XOR2_X1 U921 ( .A(G101), .B(n1220), .Z(G3) );
AND3_X1 U922 ( .A1(n1095), .A2(n1061), .A3(n1074), .ZN(n1220) );
XNOR2_X1 U923 ( .A(G125), .B(n1233), .ZN(G27) );
NAND3_X1 U924 ( .A1(n1086), .A2(n1107), .A3(n1264), .ZN(n1233) );
NOR3_X1 U925 ( .A1(n1071), .A2(n1262), .A3(n1072), .ZN(n1264) );
AND2_X1 U926 ( .A1(n1101), .A2(n1265), .ZN(n1262) );
NAND4_X1 U927 ( .A1(G953), .A2(G902), .A3(n1266), .A4(n1139), .ZN(n1265) );
INV_X1 U928 ( .A(G900), .ZN(n1139) );
XNOR2_X1 U929 ( .A(G122), .B(n1267), .ZN(G24) );
NAND2_X1 U930 ( .A1(n1094), .A2(n1268), .ZN(n1267) );
XOR2_X1 U931 ( .A(KEYINPUT7), .B(n1224), .Z(n1268) );
AND4_X1 U932 ( .A1(n1222), .A2(n1254), .A3(n1130), .A4(n1269), .ZN(n1224) );
NOR2_X1 U933 ( .A1(n1062), .A2(n1071), .ZN(n1269) );
INV_X1 U934 ( .A(n1080), .ZN(n1071) );
INV_X1 U935 ( .A(n1087), .ZN(n1062) );
NOR2_X1 U936 ( .A1(n1244), .A2(n1243), .ZN(n1087) );
NAND2_X1 U937 ( .A1(n1270), .A2(n1271), .ZN(G21) );
OR2_X1 U938 ( .A1(n1272), .A2(KEYINPUT39), .ZN(n1271) );
XOR2_X1 U939 ( .A(n1273), .B(n1274), .Z(n1270) );
NAND4_X1 U940 ( .A1(n1275), .A2(n1074), .A3(n1223), .A4(n1222), .ZN(n1274) );
NOR3_X1 U941 ( .A1(n1072), .A2(n1257), .A3(n1258), .ZN(n1223) );
INV_X1 U942 ( .A(n1094), .ZN(n1072) );
XNOR2_X1 U943 ( .A(n1080), .B(KEYINPUT45), .ZN(n1275) );
NAND2_X1 U944 ( .A1(KEYINPUT39), .A2(n1272), .ZN(n1273) );
XNOR2_X1 U945 ( .A(n1276), .B(n1219), .ZN(G18) );
AND2_X1 U946 ( .A1(n1277), .A2(n1059), .ZN(n1219) );
NOR2_X1 U947 ( .A1(n1254), .A2(n1278), .ZN(n1059) );
XNOR2_X1 U948 ( .A(n1279), .B(n1218), .ZN(G15) );
AND2_X1 U949 ( .A1(n1277), .A2(n1107), .ZN(n1218) );
INV_X1 U950 ( .A(n1242), .ZN(n1107) );
NAND2_X1 U951 ( .A1(n1278), .A2(n1254), .ZN(n1242) );
INV_X1 U952 ( .A(n1130), .ZN(n1278) );
AND4_X1 U953 ( .A1(n1095), .A2(n1080), .A3(n1094), .A4(n1222), .ZN(n1277) );
NOR2_X1 U954 ( .A1(n1104), .A2(n1263), .ZN(n1080) );
INV_X1 U955 ( .A(n1105), .ZN(n1263) );
NOR2_X1 U956 ( .A1(n1243), .A2(n1257), .ZN(n1095) );
INV_X1 U957 ( .A(n1244), .ZN(n1257) );
INV_X1 U958 ( .A(n1258), .ZN(n1243) );
NAND2_X1 U959 ( .A1(n1280), .A2(n1281), .ZN(G12) );
NAND2_X1 U960 ( .A1(n1217), .A2(n1282), .ZN(n1281) );
XOR2_X1 U961 ( .A(KEYINPUT30), .B(n1283), .Z(n1280) );
NOR2_X1 U962 ( .A1(n1217), .A2(n1282), .ZN(n1283) );
AND3_X1 U963 ( .A1(n1086), .A2(n1061), .A3(n1074), .ZN(n1217) );
NOR2_X1 U964 ( .A1(n1130), .A2(n1254), .ZN(n1074) );
OR2_X1 U965 ( .A1(n1284), .A2(n1118), .ZN(n1254) );
NOR3_X1 U966 ( .A1(G475), .A2(G902), .A3(n1123), .ZN(n1118) );
INV_X1 U967 ( .A(n1285), .ZN(n1123) );
AND2_X1 U968 ( .A1(n1286), .A2(n1287), .ZN(n1284) );
NAND2_X1 U969 ( .A1(n1285), .A2(n1288), .ZN(n1287) );
NAND2_X1 U970 ( .A1(n1289), .A2(n1290), .ZN(n1285) );
NAND2_X1 U971 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XOR2_X1 U972 ( .A(KEYINPUT57), .B(n1293), .Z(n1289) );
NOR2_X1 U973 ( .A1(n1292), .A2(n1291), .ZN(n1293) );
XOR2_X1 U974 ( .A(n1294), .B(n1295), .Z(n1291) );
XNOR2_X1 U975 ( .A(n1296), .B(n1297), .ZN(n1295) );
NOR3_X1 U976 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1297) );
NOR2_X1 U977 ( .A1(KEYINPUT35), .A2(n1301), .ZN(n1300) );
NOR2_X1 U978 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NOR3_X1 U979 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n1303) );
NOR2_X1 U980 ( .A1(KEYINPUT46), .A2(G131), .ZN(n1302) );
NOR2_X1 U981 ( .A1(n1307), .A2(n1308), .ZN(n1299) );
INV_X1 U982 ( .A(KEYINPUT35), .ZN(n1308) );
NOR2_X1 U983 ( .A1(n1305), .A2(n1309), .ZN(n1307) );
XNOR2_X1 U984 ( .A(n1304), .B(G131), .ZN(n1309) );
INV_X1 U985 ( .A(KEYINPUT46), .ZN(n1304) );
AND2_X1 U986 ( .A1(n1306), .A2(n1305), .ZN(n1298) );
XOR2_X1 U987 ( .A(G143), .B(n1310), .Z(n1305) );
AND3_X1 U988 ( .A1(G214), .A2(n1079), .A3(n1311), .ZN(n1310) );
INV_X1 U989 ( .A(G131), .ZN(n1306) );
NAND2_X1 U990 ( .A1(KEYINPUT18), .A2(n1312), .ZN(n1296) );
INV_X1 U991 ( .A(G125), .ZN(n1312) );
XNOR2_X1 U992 ( .A(G140), .B(n1313), .ZN(n1294) );
XOR2_X1 U993 ( .A(KEYINPUT25), .B(G146), .Z(n1313) );
XNOR2_X1 U994 ( .A(G104), .B(n1314), .ZN(n1292) );
XNOR2_X1 U995 ( .A(G122), .B(n1279), .ZN(n1314) );
XNOR2_X1 U996 ( .A(G475), .B(KEYINPUT26), .ZN(n1286) );
XOR2_X1 U997 ( .A(n1315), .B(n1185), .Z(n1130) );
INV_X1 U998 ( .A(G478), .ZN(n1185) );
NAND2_X1 U999 ( .A1(n1183), .A2(n1288), .ZN(n1315) );
XNOR2_X1 U1000 ( .A(n1316), .B(n1317), .ZN(n1183) );
XOR2_X1 U1001 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1002 ( .A(G128), .B(G122), .Z(n1319) );
XNOR2_X1 U1003 ( .A(n1320), .B(G134), .ZN(n1318) );
XOR2_X1 U1004 ( .A(n1321), .B(n1322), .Z(n1316) );
XNOR2_X1 U1005 ( .A(n1276), .B(G107), .ZN(n1322) );
NAND2_X1 U1006 ( .A1(G217), .A2(n1323), .ZN(n1321) );
AND4_X1 U1007 ( .A1(n1094), .A2(n1104), .A3(n1222), .A4(n1105), .ZN(n1061) );
NAND2_X1 U1008 ( .A1(G221), .A2(n1324), .ZN(n1105) );
NAND2_X1 U1009 ( .A1(n1101), .A2(n1325), .ZN(n1222) );
NAND4_X1 U1010 ( .A1(G953), .A2(G902), .A3(n1326), .A4(n1266), .ZN(n1325) );
XOR2_X1 U1011 ( .A(KEYINPUT53), .B(G898), .Z(n1326) );
NAND3_X1 U1012 ( .A1(n1266), .A2(n1079), .A3(G952), .ZN(n1101) );
NAND2_X1 U1013 ( .A1(G237), .A2(G234), .ZN(n1266) );
XNOR2_X1 U1014 ( .A(n1327), .B(n1328), .ZN(n1104) );
XNOR2_X1 U1015 ( .A(KEYINPUT59), .B(n1208), .ZN(n1328) );
INV_X1 U1016 ( .A(G469), .ZN(n1208) );
NAND3_X1 U1017 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1327) );
XNOR2_X1 U1018 ( .A(G902), .B(KEYINPUT13), .ZN(n1331) );
NAND2_X1 U1019 ( .A1(KEYINPUT62), .A2(n1332), .ZN(n1330) );
XNOR2_X1 U1020 ( .A(n1333), .B(n1334), .ZN(n1332) );
NAND2_X1 U1021 ( .A1(KEYINPUT33), .A2(n1335), .ZN(n1333) );
OR3_X1 U1022 ( .A1(n1334), .A2(n1335), .A3(KEYINPUT62), .ZN(n1329) );
XNOR2_X1 U1023 ( .A(n1207), .B(KEYINPUT41), .ZN(n1335) );
XNOR2_X1 U1024 ( .A(n1336), .B(n1337), .ZN(n1207) );
NAND2_X1 U1025 ( .A1(G227), .A2(n1079), .ZN(n1336) );
XNOR2_X1 U1026 ( .A(n1205), .B(n1338), .ZN(n1334) );
NOR2_X1 U1027 ( .A1(KEYINPUT20), .A2(n1144), .ZN(n1338) );
XNOR2_X1 U1028 ( .A(n1339), .B(n1340), .ZN(n1144) );
NOR2_X1 U1029 ( .A1(KEYINPUT12), .A2(n1341), .ZN(n1340) );
XNOR2_X1 U1030 ( .A(KEYINPUT5), .B(n1320), .ZN(n1341) );
INV_X1 U1031 ( .A(G143), .ZN(n1320) );
XNOR2_X1 U1032 ( .A(n1342), .B(n1197), .ZN(n1205) );
XOR2_X1 U1033 ( .A(G101), .B(n1343), .Z(n1197) );
NAND2_X1 U1034 ( .A1(n1344), .A2(n1345), .ZN(n1342) );
NAND2_X1 U1035 ( .A1(G107), .A2(n1191), .ZN(n1345) );
XOR2_X1 U1036 ( .A(KEYINPUT14), .B(n1346), .Z(n1344) );
NOR2_X1 U1037 ( .A1(G107), .A2(n1191), .ZN(n1346) );
NOR2_X1 U1038 ( .A1(n1347), .A2(n1092), .ZN(n1094) );
AND2_X1 U1039 ( .A1(G214), .A2(n1348), .ZN(n1092) );
INV_X1 U1040 ( .A(n1093), .ZN(n1347) );
XOR2_X1 U1041 ( .A(n1125), .B(n1129), .Z(n1093) );
NAND2_X1 U1042 ( .A1(G210), .A2(n1348), .ZN(n1129) );
NAND2_X1 U1043 ( .A1(n1288), .A2(n1311), .ZN(n1348) );
NAND2_X1 U1044 ( .A1(n1349), .A2(n1288), .ZN(n1125) );
XOR2_X1 U1045 ( .A(n1350), .B(n1351), .Z(n1349) );
XNOR2_X1 U1046 ( .A(n1251), .B(n1250), .ZN(n1351) );
XOR2_X1 U1047 ( .A(G125), .B(n1352), .Z(n1250) );
AND2_X1 U1048 ( .A1(n1079), .A2(G224), .ZN(n1352) );
NAND2_X1 U1049 ( .A1(n1353), .A2(n1354), .ZN(n1251) );
NAND4_X1 U1050 ( .A1(n1170), .A2(KEYINPUT4), .A3(n1355), .A4(n1356), .ZN(n1354) );
NAND2_X1 U1051 ( .A1(n1357), .A2(n1171), .ZN(n1356) );
NAND2_X1 U1052 ( .A1(n1358), .A2(n1359), .ZN(n1355) );
NAND3_X1 U1053 ( .A1(n1360), .A2(n1361), .A3(n1362), .ZN(n1353) );
NAND2_X1 U1054 ( .A1(KEYINPUT4), .A2(n1170), .ZN(n1362) );
XOR2_X1 U1055 ( .A(n1363), .B(n1364), .Z(n1170) );
NOR2_X1 U1056 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
XOR2_X1 U1057 ( .A(n1367), .B(KEYINPUT21), .Z(n1366) );
NAND2_X1 U1058 ( .A1(n1368), .A2(n1272), .ZN(n1367) );
XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(n1276), .ZN(n1368) );
NAND2_X1 U1060 ( .A1(KEYINPUT34), .A2(n1279), .ZN(n1363) );
INV_X1 U1061 ( .A(G113), .ZN(n1279) );
NAND2_X1 U1062 ( .A1(n1359), .A2(n1171), .ZN(n1361) );
INV_X1 U1063 ( .A(n1358), .ZN(n1171) );
XNOR2_X1 U1064 ( .A(KEYINPUT11), .B(n1169), .ZN(n1359) );
NAND2_X1 U1065 ( .A1(n1357), .A2(n1358), .ZN(n1360) );
XNOR2_X1 U1066 ( .A(n1369), .B(n1370), .ZN(n1358) );
XOR2_X1 U1067 ( .A(G107), .B(G101), .Z(n1370) );
NAND2_X1 U1068 ( .A1(KEYINPUT9), .A2(n1191), .ZN(n1369) );
INV_X1 U1069 ( .A(G104), .ZN(n1191) );
XNOR2_X1 U1070 ( .A(KEYINPUT38), .B(n1371), .ZN(n1357) );
INV_X1 U1071 ( .A(n1169), .ZN(n1371) );
XOR2_X1 U1072 ( .A(G110), .B(G122), .Z(n1169) );
XOR2_X1 U1073 ( .A(KEYINPUT31), .B(n1372), .Z(n1350) );
NOR2_X1 U1074 ( .A1(KEYINPUT37), .A2(n1249), .ZN(n1372) );
NOR2_X1 U1075 ( .A1(n1258), .A2(n1244), .ZN(n1086) );
XOR2_X1 U1076 ( .A(n1120), .B(KEYINPUT51), .Z(n1244) );
XOR2_X1 U1077 ( .A(n1373), .B(n1201), .Z(n1120) );
INV_X1 U1078 ( .A(G472), .ZN(n1201) );
NAND2_X1 U1079 ( .A1(n1374), .A2(n1288), .ZN(n1373) );
XNOR2_X1 U1080 ( .A(n1343), .B(n1375), .ZN(n1374) );
XNOR2_X1 U1081 ( .A(n1376), .B(n1196), .ZN(n1375) );
XOR2_X1 U1082 ( .A(n1249), .B(n1377), .Z(n1196) );
NOR2_X1 U1083 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
XOR2_X1 U1084 ( .A(n1380), .B(KEYINPUT8), .Z(n1379) );
NAND2_X1 U1085 ( .A1(G113), .A2(n1381), .ZN(n1380) );
XNOR2_X1 U1086 ( .A(n1272), .B(G116), .ZN(n1381) );
NOR3_X1 U1087 ( .A1(n1382), .A2(G113), .A3(n1365), .ZN(n1378) );
NOR2_X1 U1088 ( .A1(n1272), .A2(G116), .ZN(n1365) );
NOR2_X1 U1089 ( .A1(G119), .A2(n1276), .ZN(n1382) );
INV_X1 U1090 ( .A(G116), .ZN(n1276) );
XNOR2_X1 U1091 ( .A(G143), .B(n1339), .ZN(n1249) );
NAND2_X1 U1092 ( .A1(n1383), .A2(n1384), .ZN(n1376) );
NAND2_X1 U1093 ( .A1(n1200), .A2(G101), .ZN(n1384) );
XOR2_X1 U1094 ( .A(KEYINPUT61), .B(n1385), .Z(n1383) );
NOR2_X1 U1095 ( .A1(n1200), .A2(G101), .ZN(n1385) );
AND3_X1 U1096 ( .A1(n1311), .A2(n1079), .A3(G210), .ZN(n1200) );
INV_X1 U1097 ( .A(G237), .ZN(n1311) );
XNOR2_X1 U1098 ( .A(n1386), .B(n1145), .ZN(n1343) );
XNOR2_X1 U1099 ( .A(n1387), .B(n1388), .ZN(n1145) );
XNOR2_X1 U1100 ( .A(G134), .B(G131), .ZN(n1387) );
XNOR2_X1 U1101 ( .A(KEYINPUT56), .B(KEYINPUT55), .ZN(n1386) );
XNOR2_X1 U1102 ( .A(n1389), .B(n1131), .ZN(n1258) );
NOR2_X1 U1103 ( .A1(n1177), .A2(G902), .ZN(n1131) );
INV_X1 U1104 ( .A(n1181), .ZN(n1177) );
XOR2_X1 U1105 ( .A(n1390), .B(n1391), .Z(n1181) );
XOR2_X1 U1106 ( .A(n1392), .B(n1393), .Z(n1391) );
XNOR2_X1 U1107 ( .A(n1394), .B(n1272), .ZN(n1393) );
INV_X1 U1108 ( .A(G119), .ZN(n1272) );
NAND2_X1 U1109 ( .A1(n1323), .A2(G221), .ZN(n1394) );
AND2_X1 U1110 ( .A1(G234), .A2(n1079), .ZN(n1323) );
INV_X1 U1111 ( .A(G953), .ZN(n1079) );
XNOR2_X1 U1112 ( .A(KEYINPUT25), .B(G125), .ZN(n1392) );
XNOR2_X1 U1113 ( .A(n1388), .B(n1395), .ZN(n1390) );
XNOR2_X1 U1114 ( .A(n1337), .B(n1339), .ZN(n1395) );
XNOR2_X1 U1115 ( .A(G128), .B(G146), .ZN(n1339) );
XNOR2_X1 U1116 ( .A(n1282), .B(G140), .ZN(n1337) );
INV_X1 U1117 ( .A(G110), .ZN(n1282) );
XOR2_X1 U1118 ( .A(G137), .B(KEYINPUT16), .Z(n1388) );
NAND2_X1 U1119 ( .A1(n1396), .A2(KEYINPUT0), .ZN(n1389) );
XOR2_X1 U1120 ( .A(n1132), .B(KEYINPUT24), .Z(n1396) );
NAND2_X1 U1121 ( .A1(G217), .A2(n1324), .ZN(n1132) );
NAND2_X1 U1122 ( .A1(G234), .A2(n1288), .ZN(n1324) );
INV_X1 U1123 ( .A(G902), .ZN(n1288) );
endmodule


