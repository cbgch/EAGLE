//Key = 1100001110000000111000110011101010010100101100000111011000111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332;

XNOR2_X1 U740 ( .A(G107), .B(n1016), .ZN(G9) );
NOR2_X1 U741 ( .A1(n1017), .A2(n1018), .ZN(G75) );
NOR4_X1 U742 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
XOR2_X1 U743 ( .A(n1023), .B(KEYINPUT11), .Z(n1022) );
NAND2_X1 U744 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
OR2_X1 U745 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND3_X1 U746 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1024) );
NAND3_X1 U747 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1029) );
NAND2_X1 U748 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND3_X1 U749 ( .A1(n1036), .A2(n1037), .A3(n1034), .ZN(n1032) );
NAND2_X1 U750 ( .A1(n1038), .A2(n1039), .ZN(n1031) );
NOR2_X1 U751 ( .A1(n1040), .A2(n1026), .ZN(n1021) );
NAND3_X1 U752 ( .A1(n1038), .A2(n1034), .A3(n1030), .ZN(n1026) );
INV_X1 U753 ( .A(n1041), .ZN(n1040) );
NAND3_X1 U754 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1019) );
NAND3_X1 U755 ( .A1(n1028), .A2(n1045), .A3(n1030), .ZN(n1044) );
INV_X1 U756 ( .A(n1046), .ZN(n1030) );
NAND3_X1 U757 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1045) );
NAND2_X1 U758 ( .A1(n1050), .A2(n1037), .ZN(n1049) );
NAND4_X1 U759 ( .A1(n1051), .A2(n1034), .A3(n1052), .A4(n1053), .ZN(n1048) );
NAND3_X1 U760 ( .A1(n1054), .A2(n1055), .A3(n1038), .ZN(n1047) );
NOR2_X1 U761 ( .A1(n1056), .A2(n1057), .ZN(n1038) );
INV_X1 U762 ( .A(n1058), .ZN(n1054) );
NOR3_X1 U763 ( .A1(n1059), .A2(G953), .A3(G952), .ZN(n1017) );
INV_X1 U764 ( .A(n1042), .ZN(n1059) );
NAND4_X1 U765 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1042) );
NOR4_X1 U766 ( .A1(n1064), .A2(n1065), .A3(n1056), .A4(n1066), .ZN(n1063) );
XNOR2_X1 U767 ( .A(n1067), .B(KEYINPUT17), .ZN(n1064) );
NOR2_X1 U768 ( .A1(n1068), .A2(n1055), .ZN(n1062) );
NAND2_X1 U769 ( .A1(G478), .A2(n1069), .ZN(n1061) );
XOR2_X1 U770 ( .A(n1070), .B(n1071), .Z(n1060) );
XNOR2_X1 U771 ( .A(KEYINPUT56), .B(n1072), .ZN(n1071) );
NOR2_X1 U772 ( .A1(n1073), .A2(KEYINPUT15), .ZN(n1070) );
XOR2_X1 U773 ( .A(n1074), .B(n1075), .Z(G72) );
XOR2_X1 U774 ( .A(n1076), .B(n1077), .Z(n1075) );
NOR2_X1 U775 ( .A1(n1078), .A2(G953), .ZN(n1077) );
AND2_X1 U776 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U777 ( .A1(n1081), .A2(n1082), .ZN(n1076) );
NAND2_X1 U778 ( .A1(G953), .A2(n1083), .ZN(n1082) );
XNOR2_X1 U779 ( .A(n1084), .B(n1085), .ZN(n1081) );
XOR2_X1 U780 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U781 ( .A1(KEYINPUT47), .A2(n1088), .ZN(n1087) );
NAND2_X1 U782 ( .A1(G953), .A2(n1089), .ZN(n1074) );
NAND2_X1 U783 ( .A1(G900), .A2(G227), .ZN(n1089) );
XOR2_X1 U784 ( .A(n1090), .B(n1091), .Z(G69) );
XOR2_X1 U785 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND2_X1 U786 ( .A1(G953), .A2(n1094), .ZN(n1093) );
NAND2_X1 U787 ( .A1(G898), .A2(G224), .ZN(n1094) );
NAND2_X1 U788 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
NAND2_X1 U789 ( .A1(G953), .A2(n1097), .ZN(n1096) );
XNOR2_X1 U790 ( .A(n1098), .B(n1099), .ZN(n1095) );
NOR2_X1 U791 ( .A1(n1100), .A2(G953), .ZN(n1090) );
NOR2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(G66) );
NOR2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XOR2_X1 U794 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U795 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U796 ( .A1(n1109), .A2(n1110), .ZN(n1105) );
NOR2_X1 U797 ( .A1(n1109), .A2(n1110), .ZN(n1103) );
INV_X1 U798 ( .A(KEYINPUT5), .ZN(n1110) );
NOR2_X1 U799 ( .A1(n1101), .A2(n1111), .ZN(G63) );
XNOR2_X1 U800 ( .A(n1112), .B(n1113), .ZN(n1111) );
XOR2_X1 U801 ( .A(KEYINPUT24), .B(n1114), .Z(n1113) );
NOR2_X1 U802 ( .A1(n1115), .A2(n1108), .ZN(n1114) );
NOR2_X1 U803 ( .A1(n1101), .A2(n1116), .ZN(G60) );
XNOR2_X1 U804 ( .A(n1117), .B(n1118), .ZN(n1116) );
AND2_X1 U805 ( .A1(G475), .A2(n1119), .ZN(n1118) );
XOR2_X1 U806 ( .A(G104), .B(n1120), .Z(G6) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NOR3_X1 U808 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(G57) );
AND2_X1 U809 ( .A1(KEYINPUT54), .A2(n1101), .ZN(n1125) );
NOR3_X1 U810 ( .A1(KEYINPUT54), .A2(n1126), .A3(n1043), .ZN(n1124) );
NOR2_X1 U811 ( .A1(n1127), .A2(n1128), .ZN(n1123) );
XOR2_X1 U812 ( .A(KEYINPUT12), .B(n1129), .Z(n1128) );
NOR2_X1 U813 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U814 ( .A(n1132), .B(KEYINPUT43), .Z(n1130) );
NOR2_X1 U815 ( .A1(n1133), .A2(n1132), .ZN(n1127) );
XNOR2_X1 U816 ( .A(n1134), .B(n1135), .ZN(n1132) );
XOR2_X1 U817 ( .A(n1136), .B(n1137), .Z(n1135) );
NOR2_X1 U818 ( .A1(KEYINPUT36), .A2(n1138), .ZN(n1137) );
AND2_X1 U819 ( .A1(G472), .A2(n1119), .ZN(n1136) );
NOR2_X1 U820 ( .A1(n1101), .A2(n1139), .ZN(G54) );
XOR2_X1 U821 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U822 ( .A1(KEYINPUT63), .A2(n1142), .ZN(n1141) );
XOR2_X1 U823 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U824 ( .A(n1145), .B(n1146), .Z(n1144) );
XNOR2_X1 U825 ( .A(G140), .B(n1147), .ZN(n1146) );
XOR2_X1 U826 ( .A(KEYINPUT38), .B(KEYINPUT32), .Z(n1145) );
XOR2_X1 U827 ( .A(n1148), .B(n1149), .Z(n1143) );
XNOR2_X1 U828 ( .A(n1150), .B(n1151), .ZN(n1148) );
NAND2_X1 U829 ( .A1(KEYINPUT6), .A2(n1152), .ZN(n1151) );
NAND2_X1 U830 ( .A1(KEYINPUT1), .A2(n1153), .ZN(n1150) );
NAND2_X1 U831 ( .A1(n1119), .A2(G469), .ZN(n1140) );
INV_X1 U832 ( .A(n1108), .ZN(n1119) );
NOR2_X1 U833 ( .A1(n1101), .A2(n1154), .ZN(G51) );
XOR2_X1 U834 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U835 ( .A1(n1072), .A2(n1108), .ZN(n1156) );
NAND2_X1 U836 ( .A1(G902), .A2(n1020), .ZN(n1108) );
NAND3_X1 U837 ( .A1(n1080), .A2(n1157), .A3(n1100), .ZN(n1020) );
AND4_X1 U838 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1100) );
AND4_X1 U839 ( .A1(n1016), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1161) );
NAND3_X1 U840 ( .A1(n1035), .A2(n1041), .A3(n1165), .ZN(n1016) );
INV_X1 U841 ( .A(n1121), .ZN(n1035) );
NAND2_X1 U842 ( .A1(n1166), .A2(n1053), .ZN(n1121) );
NOR2_X1 U843 ( .A1(n1167), .A2(n1168), .ZN(n1160) );
NOR3_X1 U844 ( .A1(n1169), .A2(n1057), .A3(n1122), .ZN(n1168) );
INV_X1 U845 ( .A(n1053), .ZN(n1057) );
XOR2_X1 U846 ( .A(KEYINPUT8), .B(n1166), .Z(n1169) );
XNOR2_X1 U847 ( .A(KEYINPUT37), .B(n1079), .ZN(n1157) );
AND3_X1 U848 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1080) );
AND3_X1 U849 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1172) );
NAND2_X1 U850 ( .A1(n1176), .A2(n1177), .ZN(n1170) );
NAND3_X1 U851 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1177) );
NAND2_X1 U852 ( .A1(n1181), .A2(n1039), .ZN(n1180) );
NAND3_X1 U853 ( .A1(n1166), .A2(n1182), .A3(n1050), .ZN(n1179) );
NAND2_X1 U854 ( .A1(n1034), .A2(n1183), .ZN(n1178) );
NOR2_X1 U855 ( .A1(n1184), .A2(n1185), .ZN(n1155) );
XOR2_X1 U856 ( .A(n1186), .B(KEYINPUT59), .Z(n1185) );
NAND2_X1 U857 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NOR2_X1 U858 ( .A1(n1188), .A2(n1187), .ZN(n1184) );
XOR2_X1 U859 ( .A(KEYINPUT48), .B(n1189), .Z(n1187) );
XOR2_X1 U860 ( .A(n1190), .B(n1191), .Z(n1188) );
XOR2_X1 U861 ( .A(KEYINPUT9), .B(n1192), .Z(n1191) );
NOR2_X1 U862 ( .A1(KEYINPUT34), .A2(n1193), .ZN(n1192) );
AND2_X1 U863 ( .A1(G953), .A2(n1126), .ZN(n1101) );
XOR2_X1 U864 ( .A(G952), .B(KEYINPUT50), .Z(n1126) );
XOR2_X1 U865 ( .A(n1194), .B(n1195), .Z(G48) );
NOR2_X1 U866 ( .A1(KEYINPUT31), .A2(n1196), .ZN(n1195) );
INV_X1 U867 ( .A(G146), .ZN(n1196) );
NOR4_X1 U868 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1027), .ZN(n1194) );
NOR2_X1 U869 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
INV_X1 U870 ( .A(KEYINPUT25), .ZN(n1201) );
NOR2_X1 U871 ( .A1(n1202), .A2(n1182), .ZN(n1200) );
NOR2_X1 U872 ( .A1(KEYINPUT25), .A2(n1181), .ZN(n1197) );
XOR2_X1 U873 ( .A(n1171), .B(n1203), .Z(G45) );
NAND2_X1 U874 ( .A1(KEYINPUT16), .A2(G143), .ZN(n1203) );
NAND4_X1 U875 ( .A1(n1183), .A2(n1039), .A3(n1066), .A4(n1204), .ZN(n1171) );
XOR2_X1 U876 ( .A(n1205), .B(G140), .Z(G42) );
NAND2_X1 U877 ( .A1(KEYINPUT60), .A2(n1206), .ZN(n1205) );
NAND4_X1 U878 ( .A1(n1050), .A2(n1176), .A3(n1166), .A4(n1207), .ZN(n1206) );
XNOR2_X1 U879 ( .A(KEYINPUT58), .B(n1182), .ZN(n1207) );
NOR3_X1 U880 ( .A1(n1065), .A2(n1208), .A3(n1209), .ZN(n1050) );
INV_X1 U881 ( .A(n1034), .ZN(n1209) );
XNOR2_X1 U882 ( .A(G137), .B(n1173), .ZN(G39) );
NAND3_X1 U883 ( .A1(n1034), .A2(n1028), .A3(n1181), .ZN(n1173) );
XNOR2_X1 U884 ( .A(G134), .B(n1175), .ZN(G36) );
NAND3_X1 U885 ( .A1(n1183), .A2(n1041), .A3(n1034), .ZN(n1175) );
INV_X1 U886 ( .A(n1210), .ZN(n1183) );
XNOR2_X1 U887 ( .A(n1211), .B(n1212), .ZN(G33) );
NOR3_X1 U888 ( .A1(n1210), .A2(n1213), .A3(n1027), .ZN(n1212) );
XNOR2_X1 U889 ( .A(n1034), .B(KEYINPUT52), .ZN(n1213) );
NOR2_X1 U890 ( .A1(n1058), .A2(n1055), .ZN(n1034) );
INV_X1 U891 ( .A(n1214), .ZN(n1055) );
NAND3_X1 U892 ( .A1(n1166), .A2(n1182), .A3(n1036), .ZN(n1210) );
XNOR2_X1 U893 ( .A(G128), .B(n1079), .ZN(G30) );
NAND3_X1 U894 ( .A1(n1039), .A2(n1041), .A3(n1181), .ZN(n1079) );
NOR2_X1 U895 ( .A1(n1202), .A2(n1215), .ZN(n1181) );
NAND3_X1 U896 ( .A1(n1067), .A2(n1065), .A3(n1166), .ZN(n1202) );
XNOR2_X1 U897 ( .A(n1216), .B(n1167), .ZN(G3) );
AND2_X1 U898 ( .A1(n1036), .A2(n1217), .ZN(n1167) );
XOR2_X1 U899 ( .A(n1174), .B(n1218), .Z(G27) );
NAND2_X1 U900 ( .A1(KEYINPUT35), .A2(G125), .ZN(n1218) );
NAND4_X1 U901 ( .A1(n1219), .A2(n1037), .A3(n1176), .A4(n1220), .ZN(n1174) );
NOR3_X1 U902 ( .A1(n1199), .A2(n1215), .A3(n1208), .ZN(n1220) );
INV_X1 U903 ( .A(n1067), .ZN(n1208) );
INV_X1 U904 ( .A(n1182), .ZN(n1215) );
NAND2_X1 U905 ( .A1(n1046), .A2(n1221), .ZN(n1182) );
NAND4_X1 U906 ( .A1(G953), .A2(G902), .A3(n1222), .A4(n1083), .ZN(n1221) );
INV_X1 U907 ( .A(G900), .ZN(n1083) );
XNOR2_X1 U908 ( .A(G122), .B(n1158), .ZN(G24) );
NAND4_X1 U909 ( .A1(n1223), .A2(n1053), .A3(n1066), .A4(n1204), .ZN(n1158) );
NOR2_X1 U910 ( .A1(n1065), .A2(n1067), .ZN(n1053) );
NAND2_X1 U911 ( .A1(n1224), .A2(n1225), .ZN(G21) );
NAND2_X1 U912 ( .A1(G119), .A2(n1159), .ZN(n1225) );
XOR2_X1 U913 ( .A(KEYINPUT26), .B(n1226), .Z(n1224) );
NOR2_X1 U914 ( .A1(G119), .A2(n1159), .ZN(n1226) );
NAND4_X1 U915 ( .A1(n1223), .A2(n1028), .A3(n1067), .A4(n1065), .ZN(n1159) );
XOR2_X1 U916 ( .A(n1164), .B(n1227), .Z(G18) );
NAND2_X1 U917 ( .A1(n1228), .A2(KEYINPUT62), .ZN(n1227) );
XNOR2_X1 U918 ( .A(G116), .B(KEYINPUT0), .ZN(n1228) );
NAND3_X1 U919 ( .A1(n1036), .A2(n1041), .A3(n1223), .ZN(n1164) );
AND2_X1 U920 ( .A1(n1037), .A2(n1165), .ZN(n1223) );
NAND2_X1 U921 ( .A1(n1229), .A2(n1230), .ZN(n1041) );
OR3_X1 U922 ( .A1(n1066), .A2(n1231), .A3(KEYINPUT20), .ZN(n1230) );
NAND2_X1 U923 ( .A1(KEYINPUT20), .A2(n1028), .ZN(n1229) );
XNOR2_X1 U924 ( .A(G113), .B(n1163), .ZN(G15) );
NAND3_X1 U925 ( .A1(n1232), .A2(n1037), .A3(n1036), .ZN(n1163) );
NOR2_X1 U926 ( .A1(n1067), .A2(n1219), .ZN(n1036) );
INV_X1 U927 ( .A(n1056), .ZN(n1037) );
NAND2_X1 U928 ( .A1(n1052), .A2(n1233), .ZN(n1056) );
INV_X1 U929 ( .A(n1122), .ZN(n1232) );
NAND2_X1 U930 ( .A1(n1176), .A2(n1165), .ZN(n1122) );
INV_X1 U931 ( .A(n1027), .ZN(n1176) );
NAND2_X1 U932 ( .A1(n1231), .A2(n1066), .ZN(n1027) );
XNOR2_X1 U933 ( .A(G110), .B(n1162), .ZN(G12) );
NAND3_X1 U934 ( .A1(n1219), .A2(n1067), .A3(n1217), .ZN(n1162) );
AND3_X1 U935 ( .A1(n1028), .A2(n1166), .A3(n1165), .ZN(n1217) );
AND2_X1 U936 ( .A1(n1039), .A2(n1234), .ZN(n1165) );
NAND2_X1 U937 ( .A1(n1235), .A2(n1046), .ZN(n1234) );
NAND3_X1 U938 ( .A1(n1222), .A2(n1043), .A3(G952), .ZN(n1046) );
NAND4_X1 U939 ( .A1(G953), .A2(G902), .A3(n1222), .A4(n1097), .ZN(n1235) );
INV_X1 U940 ( .A(G898), .ZN(n1097) );
NAND2_X1 U941 ( .A1(G237), .A2(G234), .ZN(n1222) );
INV_X1 U942 ( .A(n1199), .ZN(n1039) );
NAND2_X1 U943 ( .A1(n1236), .A2(n1058), .ZN(n1199) );
XNOR2_X1 U944 ( .A(n1073), .B(n1072), .ZN(n1058) );
NAND2_X1 U945 ( .A1(G210), .A2(n1237), .ZN(n1072) );
AND2_X1 U946 ( .A1(n1238), .A2(n1239), .ZN(n1073) );
XNOR2_X1 U947 ( .A(n1189), .B(n1240), .ZN(n1238) );
XNOR2_X1 U948 ( .A(n1193), .B(n1190), .ZN(n1240) );
XOR2_X1 U949 ( .A(G125), .B(n1241), .Z(n1190) );
NAND2_X1 U950 ( .A1(G224), .A2(n1043), .ZN(n1193) );
XNOR2_X1 U951 ( .A(n1242), .B(n1098), .ZN(n1189) );
XOR2_X1 U952 ( .A(G110), .B(G122), .Z(n1098) );
NAND2_X1 U953 ( .A1(KEYINPUT49), .A2(n1099), .ZN(n1242) );
XOR2_X1 U954 ( .A(n1243), .B(n1244), .Z(n1099) );
XNOR2_X1 U955 ( .A(G101), .B(n1245), .ZN(n1244) );
NAND2_X1 U956 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
OR2_X1 U957 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
XOR2_X1 U958 ( .A(n1250), .B(KEYINPUT29), .Z(n1246) );
NAND2_X1 U959 ( .A1(n1249), .A2(n1248), .ZN(n1250) );
INV_X1 U960 ( .A(G113), .ZN(n1248) );
XOR2_X1 U961 ( .A(G116), .B(n1251), .Z(n1249) );
NOR2_X1 U962 ( .A1(G119), .A2(KEYINPUT33), .ZN(n1251) );
XNOR2_X1 U963 ( .A(KEYINPUT7), .B(n1214), .ZN(n1236) );
NAND2_X1 U964 ( .A1(G214), .A2(n1237), .ZN(n1214) );
NAND2_X1 U965 ( .A1(n1252), .A2(n1239), .ZN(n1237) );
INV_X1 U966 ( .A(G237), .ZN(n1252) );
NOR2_X1 U967 ( .A1(n1052), .A2(n1051), .ZN(n1166) );
INV_X1 U968 ( .A(n1233), .ZN(n1051) );
NAND2_X1 U969 ( .A1(n1253), .A2(G221), .ZN(n1233) );
XOR2_X1 U970 ( .A(n1254), .B(KEYINPUT39), .Z(n1253) );
XOR2_X1 U971 ( .A(n1255), .B(G469), .Z(n1052) );
NAND3_X1 U972 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1255) );
XNOR2_X1 U973 ( .A(KEYINPUT27), .B(n1239), .ZN(n1258) );
NAND2_X1 U974 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
NAND2_X1 U975 ( .A1(n1149), .A2(n1261), .ZN(n1260) );
XNOR2_X1 U976 ( .A(n1262), .B(n1263), .ZN(n1259) );
NAND2_X1 U977 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
NAND2_X1 U978 ( .A1(KEYINPUT45), .A2(n1152), .ZN(n1265) );
OR2_X1 U979 ( .A1(n1152), .A2(KEYINPUT2), .ZN(n1264) );
NAND3_X1 U980 ( .A1(n1149), .A2(n1261), .A3(n1266), .ZN(n1256) );
XNOR2_X1 U981 ( .A(n1267), .B(n1268), .ZN(n1266) );
INV_X1 U982 ( .A(n1263), .ZN(n1268) );
XOR2_X1 U983 ( .A(n1153), .B(n1269), .Z(n1263) );
XOR2_X1 U984 ( .A(G140), .B(n1270), .Z(n1269) );
NOR2_X1 U985 ( .A1(KEYINPUT55), .A2(n1147), .ZN(n1270) );
AND2_X1 U986 ( .A1(G227), .A2(n1043), .ZN(n1153) );
NAND2_X1 U987 ( .A1(n1271), .A2(n1272), .ZN(n1267) );
NAND2_X1 U988 ( .A1(KEYINPUT2), .A2(n1152), .ZN(n1272) );
OR2_X1 U989 ( .A1(n1152), .A2(KEYINPUT45), .ZN(n1271) );
XNOR2_X1 U990 ( .A(n1273), .B(n1274), .ZN(n1152) );
XNOR2_X1 U991 ( .A(KEYINPUT53), .B(n1216), .ZN(n1274) );
XNOR2_X1 U992 ( .A(n1275), .B(n1276), .ZN(n1273) );
INV_X1 U993 ( .A(n1084), .ZN(n1276) );
XOR2_X1 U994 ( .A(n1277), .B(n1278), .Z(n1084) );
NAND2_X1 U995 ( .A1(KEYINPUT22), .A2(n1243), .ZN(n1275) );
XOR2_X1 U996 ( .A(G104), .B(G107), .Z(n1243) );
INV_X1 U997 ( .A(KEYINPUT13), .ZN(n1261) );
NOR2_X1 U998 ( .A1(n1204), .A2(n1066), .ZN(n1028) );
XNOR2_X1 U999 ( .A(n1279), .B(G475), .ZN(n1066) );
NAND2_X1 U1000 ( .A1(n1117), .A2(n1239), .ZN(n1279) );
XNOR2_X1 U1001 ( .A(n1280), .B(n1281), .ZN(n1117) );
XNOR2_X1 U1002 ( .A(n1282), .B(n1283), .ZN(n1280) );
NOR2_X1 U1003 ( .A1(KEYINPUT41), .A2(n1284), .ZN(n1283) );
XNOR2_X1 U1004 ( .A(G104), .B(n1285), .ZN(n1284) );
XNOR2_X1 U1005 ( .A(n1286), .B(G113), .ZN(n1285) );
INV_X1 U1006 ( .A(G122), .ZN(n1286) );
NOR2_X1 U1007 ( .A1(KEYINPUT10), .A2(n1287), .ZN(n1282) );
XOR2_X1 U1008 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U1009 ( .A(n1290), .B(G143), .Z(n1289) );
NAND2_X1 U1010 ( .A1(n1291), .A2(G214), .ZN(n1290) );
NAND2_X1 U1011 ( .A1(KEYINPUT42), .A2(n1211), .ZN(n1288) );
INV_X1 U1012 ( .A(G131), .ZN(n1211) );
INV_X1 U1013 ( .A(n1231), .ZN(n1204) );
NOR2_X1 U1014 ( .A1(n1292), .A2(n1068), .ZN(n1231) );
AND3_X1 U1015 ( .A1(n1115), .A2(n1239), .A3(n1112), .ZN(n1068) );
AND2_X1 U1016 ( .A1(n1293), .A2(n1069), .ZN(n1292) );
NAND2_X1 U1017 ( .A1(n1112), .A2(n1239), .ZN(n1069) );
XOR2_X1 U1018 ( .A(n1294), .B(n1295), .Z(n1112) );
NOR2_X1 U1019 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
XOR2_X1 U1020 ( .A(KEYINPUT46), .B(n1298), .Z(n1297) );
NOR2_X1 U1021 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
AND2_X1 U1022 ( .A1(n1300), .A2(n1299), .ZN(n1296) );
XNOR2_X1 U1023 ( .A(n1301), .B(n1278), .ZN(n1299) );
XOR2_X1 U1024 ( .A(G128), .B(G143), .Z(n1278) );
XNOR2_X1 U1025 ( .A(G134), .B(KEYINPUT19), .ZN(n1301) );
NAND2_X1 U1026 ( .A1(n1302), .A2(n1303), .ZN(n1300) );
NAND2_X1 U1027 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
XOR2_X1 U1028 ( .A(KEYINPUT61), .B(n1306), .Z(n1302) );
NOR2_X1 U1029 ( .A1(n1304), .A2(n1305), .ZN(n1306) );
XOR2_X1 U1030 ( .A(G107), .B(KEYINPUT51), .Z(n1305) );
XNOR2_X1 U1031 ( .A(G116), .B(G122), .ZN(n1304) );
NAND3_X1 U1032 ( .A1(G234), .A2(n1043), .A3(G217), .ZN(n1294) );
XNOR2_X1 U1033 ( .A(KEYINPUT4), .B(n1115), .ZN(n1293) );
INV_X1 U1034 ( .A(G478), .ZN(n1115) );
XOR2_X1 U1035 ( .A(n1307), .B(n1107), .Z(n1067) );
NAND2_X1 U1036 ( .A1(G217), .A2(n1254), .ZN(n1107) );
NAND2_X1 U1037 ( .A1(G234), .A2(n1239), .ZN(n1254) );
OR2_X1 U1038 ( .A1(n1109), .A2(G902), .ZN(n1307) );
XOR2_X1 U1039 ( .A(n1308), .B(n1309), .Z(n1109) );
NOR2_X1 U1040 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
XOR2_X1 U1041 ( .A(n1312), .B(KEYINPUT40), .Z(n1311) );
NAND2_X1 U1042 ( .A1(n1313), .A2(G137), .ZN(n1312) );
NOR2_X1 U1043 ( .A1(G137), .A2(n1313), .ZN(n1310) );
AND3_X1 U1044 ( .A1(G221), .A2(n1043), .A3(n1314), .ZN(n1313) );
XNOR2_X1 U1045 ( .A(G234), .B(KEYINPUT23), .ZN(n1314) );
INV_X1 U1046 ( .A(G953), .ZN(n1043) );
NAND2_X1 U1047 ( .A1(n1315), .A2(n1316), .ZN(n1308) );
NAND2_X1 U1048 ( .A1(KEYINPUT30), .A2(n1317), .ZN(n1316) );
INV_X1 U1049 ( .A(n1318), .ZN(n1317) );
NAND2_X1 U1050 ( .A1(KEYINPUT14), .A2(n1318), .ZN(n1315) );
XOR2_X1 U1051 ( .A(n1281), .B(n1319), .Z(n1318) );
XNOR2_X1 U1052 ( .A(n1147), .B(n1320), .ZN(n1319) );
NOR2_X1 U1053 ( .A1(KEYINPUT21), .A2(n1321), .ZN(n1320) );
XNOR2_X1 U1054 ( .A(G119), .B(G128), .ZN(n1321) );
INV_X1 U1055 ( .A(G110), .ZN(n1147) );
XOR2_X1 U1056 ( .A(n1088), .B(n1277), .Z(n1281) );
XOR2_X1 U1057 ( .A(G125), .B(G140), .Z(n1088) );
INV_X1 U1058 ( .A(n1065), .ZN(n1219) );
XNOR2_X1 U1059 ( .A(n1322), .B(G472), .ZN(n1065) );
NAND2_X1 U1060 ( .A1(n1323), .A2(n1239), .ZN(n1322) );
INV_X1 U1061 ( .A(G902), .ZN(n1239) );
XOR2_X1 U1062 ( .A(n1138), .B(n1324), .Z(n1323) );
XNOR2_X1 U1063 ( .A(n1133), .B(n1134), .ZN(n1324) );
XOR2_X1 U1064 ( .A(n1149), .B(n1241), .Z(n1134) );
XOR2_X1 U1065 ( .A(G128), .B(n1325), .Z(n1241) );
NOR3_X1 U1066 ( .A1(n1326), .A2(KEYINPUT57), .A3(n1327), .ZN(n1325) );
NOR2_X1 U1067 ( .A1(G143), .A2(n1328), .ZN(n1327) );
XOR2_X1 U1068 ( .A(n1329), .B(KEYINPUT18), .Z(n1326) );
NAND2_X1 U1069 ( .A1(G143), .A2(n1328), .ZN(n1329) );
XOR2_X1 U1070 ( .A(n1277), .B(KEYINPUT28), .Z(n1328) );
XOR2_X1 U1071 ( .A(G146), .B(KEYINPUT3), .Z(n1277) );
XNOR2_X1 U1072 ( .A(n1086), .B(KEYINPUT44), .ZN(n1149) );
XNOR2_X1 U1073 ( .A(G131), .B(n1330), .ZN(n1086) );
XOR2_X1 U1074 ( .A(G137), .B(G134), .Z(n1330) );
INV_X1 U1075 ( .A(n1131), .ZN(n1133) );
XOR2_X1 U1076 ( .A(n1331), .B(n1216), .Z(n1131) );
INV_X1 U1077 ( .A(G101), .ZN(n1216) );
NAND2_X1 U1078 ( .A1(n1291), .A2(G210), .ZN(n1331) );
NOR2_X1 U1079 ( .A1(G953), .A2(G237), .ZN(n1291) );
XNOR2_X1 U1080 ( .A(G113), .B(n1332), .ZN(n1138) );
XOR2_X1 U1081 ( .A(G119), .B(G116), .Z(n1332) );
endmodule


