//Key = 1100010110110100100000111000101011100000110110101101100010101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
n1425, n1426, n1427, n1428, n1429, n1430;

XOR2_X1 U785 ( .A(n1085), .B(n1086), .Z(G9) );
NOR2_X1 U786 ( .A1(KEYINPUT25), .A2(n1087), .ZN(n1086) );
NOR2_X1 U787 ( .A1(n1088), .A2(n1089), .ZN(G75) );
NOR3_X1 U788 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
NOR2_X1 U789 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NAND3_X1 U790 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1090) );
NAND3_X1 U791 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1097) );
NAND2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NAND3_X1 U793 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1101) );
NAND2_X1 U794 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND3_X1 U795 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1107) );
XNOR2_X1 U796 ( .A(n1111), .B(n1112), .ZN(n1110) );
NAND2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1106) );
NAND2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U799 ( .A1(n1109), .A2(n1117), .ZN(n1116) );
OR2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U801 ( .A1(n1108), .A2(n1120), .ZN(n1115) );
NAND2_X1 U802 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
INV_X1 U803 ( .A(KEYINPUT17), .ZN(n1104) );
NAND2_X1 U804 ( .A1(n1123), .A2(n1124), .ZN(n1098) );
XOR2_X1 U805 ( .A(n1094), .B(KEYINPUT57), .Z(n1124) );
NAND4_X1 U806 ( .A1(n1108), .A2(n1113), .A3(n1125), .A4(n1109), .ZN(n1094) );
NOR2_X1 U807 ( .A1(KEYINPUT17), .A2(n1126), .ZN(n1125) );
NOR3_X1 U808 ( .A1(n1127), .A2(G953), .A3(G952), .ZN(n1088) );
INV_X1 U809 ( .A(n1095), .ZN(n1127) );
NAND4_X1 U810 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1095) );
NOR3_X1 U811 ( .A1(n1132), .A2(n1123), .A3(n1133), .ZN(n1131) );
XOR2_X1 U812 ( .A(n1134), .B(KEYINPUT24), .Z(n1130) );
NAND4_X1 U813 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1134) );
NOR2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U815 ( .A(n1141), .B(n1142), .Z(n1139) );
XNOR2_X1 U816 ( .A(KEYINPUT7), .B(n1143), .ZN(n1142) );
NAND2_X1 U817 ( .A1(n1144), .A2(n1145), .ZN(n1136) );
NAND2_X1 U818 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
NAND2_X1 U819 ( .A1(KEYINPUT42), .A2(n1148), .ZN(n1147) );
NAND2_X1 U820 ( .A1(n1149), .A2(n1150), .ZN(n1146) );
INV_X1 U821 ( .A(KEYINPUT42), .ZN(n1150) );
OR2_X1 U822 ( .A1(n1149), .A2(n1145), .ZN(n1135) );
NAND2_X1 U823 ( .A1(KEYINPUT5), .A2(n1148), .ZN(n1149) );
NAND2_X1 U824 ( .A1(G469), .A2(n1151), .ZN(n1129) );
XNOR2_X1 U825 ( .A(n1152), .B(n1153), .ZN(n1128) );
NAND2_X1 U826 ( .A1(KEYINPUT13), .A2(n1154), .ZN(n1153) );
XOR2_X1 U827 ( .A(n1155), .B(n1156), .Z(G72) );
NOR2_X1 U828 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NOR2_X1 U829 ( .A1(KEYINPUT35), .A2(n1159), .ZN(n1158) );
INV_X1 U830 ( .A(n1160), .ZN(n1159) );
NOR2_X1 U831 ( .A1(KEYINPUT40), .A2(n1160), .ZN(n1157) );
NAND2_X1 U832 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U833 ( .A1(G953), .A2(n1163), .ZN(n1162) );
XOR2_X1 U834 ( .A(n1164), .B(n1165), .Z(n1161) );
NAND2_X1 U835 ( .A1(n1166), .A2(n1167), .ZN(n1164) );
NAND3_X1 U836 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1167) );
XOR2_X1 U837 ( .A(n1171), .B(KEYINPUT54), .Z(n1166) );
NAND2_X1 U838 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NAND2_X1 U839 ( .A1(n1168), .A2(n1169), .ZN(n1173) );
INV_X1 U840 ( .A(n1174), .ZN(n1169) );
INV_X1 U841 ( .A(n1170), .ZN(n1172) );
NAND2_X1 U842 ( .A1(n1175), .A2(n1176), .ZN(n1155) );
NAND2_X1 U843 ( .A1(n1177), .A2(n1096), .ZN(n1176) );
NAND2_X1 U844 ( .A1(G953), .A2(n1178), .ZN(n1175) );
NAND2_X1 U845 ( .A1(G900), .A2(G227), .ZN(n1178) );
XOR2_X1 U846 ( .A(n1179), .B(n1180), .Z(G69) );
XOR2_X1 U847 ( .A(n1181), .B(n1182), .Z(n1180) );
NAND2_X1 U848 ( .A1(n1096), .A2(n1183), .ZN(n1182) );
NAND3_X1 U849 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1183) );
XNOR2_X1 U850 ( .A(n1187), .B(KEYINPUT39), .ZN(n1186) );
XOR2_X1 U851 ( .A(KEYINPUT41), .B(n1085), .Z(n1185) );
INV_X1 U852 ( .A(n1188), .ZN(n1184) );
NAND2_X1 U853 ( .A1(n1189), .A2(n1190), .ZN(n1181) );
NAND2_X1 U854 ( .A1(G953), .A2(n1191), .ZN(n1190) );
XOR2_X1 U855 ( .A(n1192), .B(n1193), .Z(n1189) );
NOR3_X1 U856 ( .A1(n1096), .A2(KEYINPUT26), .A3(n1194), .ZN(n1179) );
NOR2_X1 U857 ( .A1(n1195), .A2(n1191), .ZN(n1194) );
NOR2_X1 U858 ( .A1(n1196), .A2(n1197), .ZN(G66) );
XNOR2_X1 U859 ( .A(n1198), .B(n1199), .ZN(n1197) );
NAND4_X1 U860 ( .A1(n1200), .A2(n1092), .A3(n1201), .A4(n1202), .ZN(n1198) );
NAND2_X1 U861 ( .A1(KEYINPUT21), .A2(G902), .ZN(n1202) );
NAND2_X1 U862 ( .A1(n1203), .A2(n1204), .ZN(n1201) );
NAND2_X1 U863 ( .A1(KEYINPUT21), .A2(n1205), .ZN(n1203) );
XNOR2_X1 U864 ( .A(G217), .B(KEYINPUT11), .ZN(n1200) );
NOR2_X1 U865 ( .A1(n1196), .A2(n1206), .ZN(G63) );
NOR2_X1 U866 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U867 ( .A(KEYINPUT37), .B(n1209), .Z(n1208) );
NOR2_X1 U868 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U869 ( .A(KEYINPUT51), .B(n1212), .Z(n1211) );
NOR2_X1 U870 ( .A1(n1212), .A2(n1213), .ZN(n1207) );
INV_X1 U871 ( .A(n1210), .ZN(n1213) );
AND2_X1 U872 ( .A1(n1214), .A2(G478), .ZN(n1212) );
NOR2_X1 U873 ( .A1(n1196), .A2(n1215), .ZN(G60) );
NOR3_X1 U874 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
AND3_X1 U875 ( .A1(n1219), .A2(G475), .A3(n1214), .ZN(n1218) );
NOR2_X1 U876 ( .A1(n1220), .A2(n1219), .ZN(n1217) );
NOR2_X1 U877 ( .A1(n1221), .A2(n1145), .ZN(n1220) );
XNOR2_X1 U878 ( .A(G104), .B(n1222), .ZN(G6) );
NOR2_X1 U879 ( .A1(n1196), .A2(n1223), .ZN(G57) );
XNOR2_X1 U880 ( .A(n1224), .B(n1225), .ZN(n1223) );
XOR2_X1 U881 ( .A(n1226), .B(n1227), .Z(n1225) );
AND2_X1 U882 ( .A1(G472), .A2(n1214), .ZN(n1227) );
NOR2_X1 U883 ( .A1(KEYINPUT61), .A2(n1228), .ZN(n1226) );
XOR2_X1 U884 ( .A(n1229), .B(n1230), .Z(n1228) );
NAND2_X1 U885 ( .A1(n1231), .A2(n1232), .ZN(n1229) );
NAND2_X1 U886 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
XOR2_X1 U887 ( .A(n1235), .B(KEYINPUT6), .Z(n1231) );
OR2_X1 U888 ( .A1(n1234), .A2(n1233), .ZN(n1235) );
NOR2_X1 U889 ( .A1(n1196), .A2(n1236), .ZN(G54) );
XOR2_X1 U890 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U891 ( .A(n1239), .B(n1240), .Z(n1238) );
AND2_X1 U892 ( .A1(G469), .A2(n1214), .ZN(n1240) );
NOR2_X1 U893 ( .A1(n1204), .A2(n1221), .ZN(n1214) );
NAND2_X1 U894 ( .A1(KEYINPUT60), .A2(n1241), .ZN(n1239) );
XOR2_X1 U895 ( .A(n1242), .B(n1243), .Z(n1237) );
NOR2_X1 U896 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XOR2_X1 U897 ( .A(n1246), .B(KEYINPUT10), .Z(n1245) );
NAND2_X1 U898 ( .A1(n1247), .A2(n1234), .ZN(n1246) );
NOR2_X1 U899 ( .A1(n1247), .A2(n1234), .ZN(n1244) );
XOR2_X1 U900 ( .A(n1248), .B(KEYINPUT18), .Z(n1247) );
XNOR2_X1 U901 ( .A(G140), .B(n1249), .ZN(n1242) );
NOR2_X1 U902 ( .A1(G110), .A2(KEYINPUT12), .ZN(n1249) );
NOR2_X1 U903 ( .A1(n1196), .A2(n1250), .ZN(G51) );
XOR2_X1 U904 ( .A(n1251), .B(n1252), .Z(n1250) );
XOR2_X1 U905 ( .A(n1253), .B(n1254), .Z(n1252) );
NAND3_X1 U906 ( .A1(n1255), .A2(n1092), .A3(n1152), .ZN(n1254) );
INV_X1 U907 ( .A(n1256), .ZN(n1152) );
INV_X1 U908 ( .A(n1221), .ZN(n1092) );
NOR4_X1 U909 ( .A1(n1177), .A2(n1188), .A3(n1187), .A4(n1085), .ZN(n1221) );
AND3_X1 U910 ( .A1(n1119), .A2(n1109), .A3(n1257), .ZN(n1085) );
NAND3_X1 U911 ( .A1(n1258), .A2(n1222), .A3(n1259), .ZN(n1188) );
NOR3_X1 U912 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1259) );
INV_X1 U913 ( .A(n1263), .ZN(n1260) );
NAND3_X1 U914 ( .A1(n1109), .A2(n1118), .A3(n1257), .ZN(n1222) );
NAND2_X1 U915 ( .A1(n1264), .A2(n1265), .ZN(n1258) );
NAND2_X1 U916 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XOR2_X1 U917 ( .A(KEYINPUT44), .B(n1268), .Z(n1266) );
NAND4_X1 U918 ( .A1(n1269), .A2(n1270), .A3(n1271), .A4(n1272), .ZN(n1177) );
NOR4_X1 U919 ( .A1(n1273), .A2(n1274), .A3(n1275), .A4(n1276), .ZN(n1272) );
AND3_X1 U920 ( .A1(n1277), .A2(n1108), .A3(n1278), .ZN(n1276) );
NOR4_X1 U921 ( .A1(n1279), .A2(n1280), .A3(n1121), .A4(n1281), .ZN(n1275) );
XNOR2_X1 U922 ( .A(n1264), .B(KEYINPUT9), .ZN(n1280) );
INV_X1 U923 ( .A(n1282), .ZN(n1279) );
NOR2_X1 U924 ( .A1(n1283), .A2(n1284), .ZN(n1271) );
XNOR2_X1 U925 ( .A(KEYINPUT15), .B(n1204), .ZN(n1255) );
NAND2_X1 U926 ( .A1(n1285), .A2(n1286), .ZN(n1253) );
NAND4_X1 U927 ( .A1(KEYINPUT23), .A2(n1287), .A3(n1288), .A4(n1289), .ZN(n1286) );
NAND2_X1 U928 ( .A1(n1290), .A2(n1291), .ZN(n1285) );
NAND2_X1 U929 ( .A1(n1288), .A2(n1292), .ZN(n1291) );
OR2_X1 U930 ( .A1(n1289), .A2(n1287), .ZN(n1292) );
INV_X1 U931 ( .A(KEYINPUT20), .ZN(n1289) );
NAND2_X1 U932 ( .A1(KEYINPUT23), .A2(n1287), .ZN(n1290) );
NOR2_X1 U933 ( .A1(n1096), .A2(G952), .ZN(n1196) );
XOR2_X1 U934 ( .A(G146), .B(n1274), .Z(G48) );
AND3_X1 U935 ( .A1(n1293), .A2(n1118), .A3(n1278), .ZN(n1274) );
XNOR2_X1 U936 ( .A(G143), .B(n1294), .ZN(G45) );
NAND3_X1 U937 ( .A1(n1295), .A2(n1282), .A3(n1293), .ZN(n1294) );
NAND3_X1 U938 ( .A1(n1296), .A2(n1297), .A3(n1298), .ZN(G42) );
NAND2_X1 U939 ( .A1(G140), .A2(n1299), .ZN(n1298) );
NAND2_X1 U940 ( .A1(n1300), .A2(KEYINPUT48), .ZN(n1299) );
XNOR2_X1 U941 ( .A(n1273), .B(KEYINPUT58), .ZN(n1300) );
NAND3_X1 U942 ( .A1(KEYINPUT48), .A2(n1301), .A3(n1273), .ZN(n1297) );
OR2_X1 U943 ( .A1(n1273), .A2(KEYINPUT48), .ZN(n1296) );
NOR3_X1 U944 ( .A1(n1122), .A2(n1302), .A3(n1303), .ZN(n1273) );
XOR2_X1 U945 ( .A(n1304), .B(n1305), .Z(G39) );
NOR2_X1 U946 ( .A1(KEYINPUT31), .A2(n1306), .ZN(n1305) );
XNOR2_X1 U947 ( .A(KEYINPUT36), .B(n1307), .ZN(n1306) );
NAND3_X1 U948 ( .A1(n1277), .A2(n1278), .A3(n1308), .ZN(n1304) );
XNOR2_X1 U949 ( .A(n1108), .B(KEYINPUT32), .ZN(n1308) );
XOR2_X1 U950 ( .A(G134), .B(n1284), .Z(G36) );
AND3_X1 U951 ( .A1(n1295), .A2(n1119), .A3(n1277), .ZN(n1284) );
XOR2_X1 U952 ( .A(G131), .B(n1283), .Z(G33) );
NOR3_X1 U953 ( .A1(n1121), .A2(n1302), .A3(n1303), .ZN(n1283) );
INV_X1 U954 ( .A(n1277), .ZN(n1303) );
NOR3_X1 U955 ( .A1(n1309), .A2(n1123), .A3(n1281), .ZN(n1277) );
INV_X1 U956 ( .A(n1102), .ZN(n1123) );
XNOR2_X1 U957 ( .A(G128), .B(n1269), .ZN(G30) );
NAND3_X1 U958 ( .A1(n1293), .A2(n1119), .A3(n1278), .ZN(n1269) );
NOR2_X1 U959 ( .A1(n1281), .A2(n1093), .ZN(n1293) );
NAND3_X1 U960 ( .A1(n1111), .A2(n1112), .A3(n1310), .ZN(n1281) );
XNOR2_X1 U961 ( .A(n1311), .B(n1261), .ZN(G3) );
AND3_X1 U962 ( .A1(n1108), .A2(n1257), .A3(n1295), .ZN(n1261) );
XNOR2_X1 U963 ( .A(G125), .B(n1270), .ZN(G27) );
NAND4_X1 U964 ( .A1(n1312), .A2(n1313), .A3(n1118), .A4(n1310), .ZN(n1270) );
NAND2_X1 U965 ( .A1(n1314), .A2(n1315), .ZN(n1310) );
NAND2_X1 U966 ( .A1(n1316), .A2(n1163), .ZN(n1315) );
INV_X1 U967 ( .A(G900), .ZN(n1163) );
XOR2_X1 U968 ( .A(G122), .B(n1317), .Z(G24) );
NOR3_X1 U969 ( .A1(n1318), .A2(KEYINPUT45), .A3(n1267), .ZN(n1317) );
NAND4_X1 U970 ( .A1(n1113), .A2(n1109), .A3(n1282), .A4(n1319), .ZN(n1267) );
NAND2_X1 U971 ( .A1(n1320), .A2(n1321), .ZN(n1282) );
NAND2_X1 U972 ( .A1(n1119), .A2(n1322), .ZN(n1321) );
NAND3_X1 U973 ( .A1(n1323), .A2(n1324), .A3(KEYINPUT52), .ZN(n1320) );
NOR2_X1 U974 ( .A1(n1325), .A2(n1140), .ZN(n1109) );
XNOR2_X1 U975 ( .A(KEYINPUT34), .B(n1093), .ZN(n1318) );
XNOR2_X1 U976 ( .A(G119), .B(n1263), .ZN(G21) );
NAND4_X1 U977 ( .A1(n1278), .A2(n1313), .A3(n1108), .A4(n1319), .ZN(n1263) );
AND2_X1 U978 ( .A1(n1325), .A2(n1140), .ZN(n1278) );
NAND2_X1 U979 ( .A1(n1326), .A2(n1327), .ZN(G18) );
NAND2_X1 U980 ( .A1(G116), .A2(n1328), .ZN(n1327) );
XOR2_X1 U981 ( .A(n1329), .B(KEYINPUT38), .Z(n1326) );
OR2_X1 U982 ( .A1(n1328), .A2(G116), .ZN(n1329) );
NAND2_X1 U983 ( .A1(n1268), .A2(n1264), .ZN(n1328) );
AND4_X1 U984 ( .A1(n1295), .A2(n1113), .A3(n1119), .A4(n1319), .ZN(n1268) );
NOR2_X1 U985 ( .A1(n1137), .A2(n1324), .ZN(n1119) );
XNOR2_X1 U986 ( .A(n1330), .B(n1331), .ZN(G15) );
NOR3_X1 U987 ( .A1(KEYINPUT14), .A2(n1332), .A3(n1333), .ZN(n1331) );
NOR2_X1 U988 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
INV_X1 U989 ( .A(KEYINPUT27), .ZN(n1335) );
NOR4_X1 U990 ( .A1(n1302), .A2(n1336), .A3(n1121), .A4(n1319), .ZN(n1334) );
INV_X1 U991 ( .A(n1295), .ZN(n1121) );
INV_X1 U992 ( .A(n1118), .ZN(n1302) );
NOR2_X1 U993 ( .A1(KEYINPUT27), .A2(n1187), .ZN(n1332) );
AND4_X1 U994 ( .A1(n1295), .A2(n1313), .A3(n1118), .A4(n1319), .ZN(n1187) );
NAND2_X1 U995 ( .A1(n1337), .A2(n1338), .ZN(n1118) );
NAND2_X1 U996 ( .A1(n1108), .A2(n1322), .ZN(n1338) );
INV_X1 U997 ( .A(KEYINPUT52), .ZN(n1322) );
NAND3_X1 U998 ( .A1(n1137), .A2(n1324), .A3(KEYINPUT52), .ZN(n1337) );
INV_X1 U999 ( .A(n1323), .ZN(n1137) );
INV_X1 U1000 ( .A(n1336), .ZN(n1313) );
NAND2_X1 U1001 ( .A1(n1113), .A2(n1264), .ZN(n1336) );
NOR2_X1 U1002 ( .A1(n1111), .A2(n1133), .ZN(n1113) );
INV_X1 U1003 ( .A(n1112), .ZN(n1133) );
NOR2_X1 U1004 ( .A1(n1140), .A2(n1339), .ZN(n1295) );
XNOR2_X1 U1005 ( .A(n1340), .B(n1262), .ZN(G12) );
AND3_X1 U1006 ( .A1(n1108), .A2(n1257), .A3(n1312), .ZN(n1262) );
INV_X1 U1007 ( .A(n1122), .ZN(n1312) );
NAND2_X1 U1008 ( .A1(n1339), .A2(n1140), .ZN(n1122) );
NAND3_X1 U1009 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1140) );
NAND2_X1 U1010 ( .A1(n1344), .A2(n1199), .ZN(n1343) );
OR3_X1 U1011 ( .A1(n1199), .A2(n1344), .A3(G902), .ZN(n1342) );
NOR2_X1 U1012 ( .A1(n1345), .A2(G234), .ZN(n1344) );
XNOR2_X1 U1013 ( .A(n1346), .B(n1347), .ZN(n1199) );
XNOR2_X1 U1014 ( .A(n1340), .B(n1348), .ZN(n1347) );
XNOR2_X1 U1015 ( .A(n1307), .B(G119), .ZN(n1348) );
XOR2_X1 U1016 ( .A(n1349), .B(n1350), .Z(n1346) );
XOR2_X1 U1017 ( .A(n1351), .B(n1352), .Z(n1349) );
AND3_X1 U1018 ( .A1(G221), .A2(n1096), .A3(G234), .ZN(n1352) );
NAND2_X1 U1019 ( .A1(KEYINPUT30), .A2(n1353), .ZN(n1351) );
XOR2_X1 U1020 ( .A(KEYINPUT33), .B(G128), .Z(n1353) );
NAND2_X1 U1021 ( .A1(G217), .A2(G902), .ZN(n1341) );
INV_X1 U1022 ( .A(n1325), .ZN(n1339) );
NAND2_X1 U1023 ( .A1(n1354), .A2(n1355), .ZN(n1325) );
OR2_X1 U1024 ( .A1(n1143), .A2(n1356), .ZN(n1355) );
XOR2_X1 U1025 ( .A(n1357), .B(KEYINPUT50), .Z(n1354) );
NAND2_X1 U1026 ( .A1(n1356), .A2(n1143), .ZN(n1357) );
INV_X1 U1027 ( .A(G472), .ZN(n1143) );
XNOR2_X1 U1028 ( .A(n1141), .B(KEYINPUT29), .ZN(n1356) );
NAND2_X1 U1029 ( .A1(n1358), .A2(n1204), .ZN(n1141) );
XNOR2_X1 U1030 ( .A(n1359), .B(n1360), .ZN(n1358) );
INV_X1 U1031 ( .A(n1224), .ZN(n1360) );
XOR2_X1 U1032 ( .A(n1361), .B(n1311), .Z(n1224) );
INV_X1 U1033 ( .A(G101), .ZN(n1311) );
NAND2_X1 U1034 ( .A1(n1362), .A2(G210), .ZN(n1361) );
XOR2_X1 U1035 ( .A(n1363), .B(n1230), .Z(n1359) );
AND3_X1 U1036 ( .A1(n1364), .A2(n1365), .A3(n1366), .ZN(n1230) );
NAND2_X1 U1037 ( .A1(n1367), .A2(n1330), .ZN(n1365) );
XNOR2_X1 U1038 ( .A(n1368), .B(n1369), .ZN(n1367) );
AND2_X1 U1039 ( .A1(n1370), .A2(KEYINPUT62), .ZN(n1369) );
NAND3_X1 U1040 ( .A1(n1371), .A2(n1370), .A3(G113), .ZN(n1364) );
XNOR2_X1 U1041 ( .A(KEYINPUT62), .B(G116), .ZN(n1371) );
NAND2_X1 U1042 ( .A1(KEYINPUT8), .A2(n1372), .ZN(n1363) );
XNOR2_X1 U1043 ( .A(n1234), .B(n1233), .ZN(n1372) );
AND4_X1 U1044 ( .A1(n1264), .A2(n1111), .A3(n1112), .A4(n1319), .ZN(n1257) );
NAND2_X1 U1045 ( .A1(n1373), .A2(n1374), .ZN(n1319) );
NAND2_X1 U1046 ( .A1(n1316), .A2(n1191), .ZN(n1374) );
INV_X1 U1047 ( .A(G898), .ZN(n1191) );
NOR3_X1 U1048 ( .A1(n1204), .A2(n1126), .A3(n1096), .ZN(n1316) );
XOR2_X1 U1049 ( .A(n1314), .B(KEYINPUT59), .Z(n1373) );
NAND3_X1 U1050 ( .A1(G952), .A2(n1103), .A3(n1375), .ZN(n1314) );
XNOR2_X1 U1051 ( .A(G953), .B(KEYINPUT3), .ZN(n1375) );
INV_X1 U1052 ( .A(n1126), .ZN(n1103) );
NOR2_X1 U1053 ( .A1(n1376), .A2(n1205), .ZN(n1126) );
NAND2_X1 U1054 ( .A1(G221), .A2(n1377), .ZN(n1112) );
NAND2_X1 U1055 ( .A1(G234), .A2(n1204), .ZN(n1377) );
OR2_X1 U1056 ( .A1(n1132), .A2(n1378), .ZN(n1111) );
AND2_X1 U1057 ( .A1(n1379), .A2(n1151), .ZN(n1378) );
XOR2_X1 U1058 ( .A(KEYINPUT55), .B(G469), .Z(n1379) );
NOR2_X1 U1059 ( .A1(n1151), .A2(G469), .ZN(n1132) );
NAND2_X1 U1060 ( .A1(n1380), .A2(n1204), .ZN(n1151) );
XOR2_X1 U1061 ( .A(n1381), .B(n1382), .Z(n1380) );
XOR2_X1 U1062 ( .A(n1234), .B(n1383), .Z(n1382) );
XNOR2_X1 U1063 ( .A(G110), .B(G140), .ZN(n1383) );
NAND3_X1 U1064 ( .A1(n1384), .A2(n1385), .A3(n1168), .ZN(n1234) );
NAND2_X1 U1065 ( .A1(n1386), .A2(n1307), .ZN(n1168) );
NAND2_X1 U1066 ( .A1(n1386), .A2(n1387), .ZN(n1385) );
INV_X1 U1067 ( .A(KEYINPUT63), .ZN(n1387) );
NAND2_X1 U1068 ( .A1(n1174), .A2(KEYINPUT63), .ZN(n1384) );
NOR2_X1 U1069 ( .A1(n1307), .A2(n1386), .ZN(n1174) );
XOR2_X1 U1070 ( .A(G131), .B(G134), .Z(n1386) );
INV_X1 U1071 ( .A(G137), .ZN(n1307) );
XOR2_X1 U1072 ( .A(n1388), .B(n1241), .Z(n1381) );
AND2_X1 U1073 ( .A1(G227), .A2(n1096), .ZN(n1241) );
INV_X1 U1074 ( .A(G953), .ZN(n1096) );
NAND2_X1 U1075 ( .A1(KEYINPUT1), .A2(n1248), .ZN(n1388) );
XOR2_X1 U1076 ( .A(n1389), .B(n1390), .Z(n1248) );
XNOR2_X1 U1077 ( .A(n1170), .B(G101), .ZN(n1389) );
XNOR2_X1 U1078 ( .A(n1391), .B(KEYINPUT49), .ZN(n1170) );
INV_X1 U1079 ( .A(n1093), .ZN(n1264) );
NAND2_X1 U1080 ( .A1(n1392), .A2(n1102), .ZN(n1093) );
NAND2_X1 U1081 ( .A1(G214), .A2(n1393), .ZN(n1102) );
XOR2_X1 U1082 ( .A(KEYINPUT46), .B(n1100), .Z(n1392) );
INV_X1 U1083 ( .A(n1309), .ZN(n1100) );
NAND2_X1 U1084 ( .A1(n1394), .A2(n1395), .ZN(n1309) );
NAND2_X1 U1085 ( .A1(n1396), .A2(n1256), .ZN(n1395) );
XOR2_X1 U1086 ( .A(KEYINPUT0), .B(n1397), .Z(n1394) );
NOR2_X1 U1087 ( .A1(n1396), .A2(n1256), .ZN(n1397) );
NAND2_X1 U1088 ( .A1(G210), .A2(n1393), .ZN(n1256) );
NAND2_X1 U1089 ( .A1(n1376), .A2(n1204), .ZN(n1393) );
INV_X1 U1090 ( .A(G237), .ZN(n1376) );
XOR2_X1 U1091 ( .A(n1154), .B(KEYINPUT43), .Z(n1396) );
NAND2_X1 U1092 ( .A1(n1398), .A2(n1204), .ZN(n1154) );
XOR2_X1 U1093 ( .A(n1399), .B(n1400), .Z(n1398) );
XOR2_X1 U1094 ( .A(n1251), .B(n1288), .Z(n1400) );
XOR2_X1 U1095 ( .A(G125), .B(n1233), .Z(n1288) );
XNOR2_X1 U1096 ( .A(n1391), .B(KEYINPUT47), .ZN(n1233) );
XNOR2_X1 U1097 ( .A(G146), .B(n1401), .ZN(n1391) );
XNOR2_X1 U1098 ( .A(n1402), .B(n1192), .ZN(n1251) );
XNOR2_X1 U1099 ( .A(n1403), .B(n1404), .ZN(n1192) );
XNOR2_X1 U1100 ( .A(G122), .B(n1340), .ZN(n1404) );
XNOR2_X1 U1101 ( .A(G101), .B(n1405), .ZN(n1403) );
NOR2_X1 U1102 ( .A1(n1406), .A2(n1407), .ZN(n1405) );
AND3_X1 U1103 ( .A1(n1408), .A2(n1087), .A3(G104), .ZN(n1407) );
NOR2_X1 U1104 ( .A1(n1390), .A2(n1408), .ZN(n1406) );
INV_X1 U1105 ( .A(KEYINPUT22), .ZN(n1408) );
XNOR2_X1 U1106 ( .A(G104), .B(n1087), .ZN(n1390) );
INV_X1 U1107 ( .A(G107), .ZN(n1087) );
NAND2_X1 U1108 ( .A1(KEYINPUT56), .A2(n1193), .ZN(n1402) );
NAND3_X1 U1109 ( .A1(n1409), .A2(n1410), .A3(n1366), .ZN(n1193) );
NAND3_X1 U1110 ( .A1(G113), .A2(n1368), .A3(G119), .ZN(n1366) );
NAND2_X1 U1111 ( .A1(n1411), .A2(n1370), .ZN(n1410) );
INV_X1 U1112 ( .A(G119), .ZN(n1370) );
XNOR2_X1 U1113 ( .A(G113), .B(G116), .ZN(n1411) );
NAND3_X1 U1114 ( .A1(G116), .A2(n1330), .A3(G119), .ZN(n1409) );
XNOR2_X1 U1115 ( .A(n1287), .B(KEYINPUT4), .ZN(n1399) );
NOR2_X1 U1116 ( .A1(n1195), .A2(G953), .ZN(n1287) );
INV_X1 U1117 ( .A(G224), .ZN(n1195) );
NOR2_X1 U1118 ( .A1(n1323), .A2(n1324), .ZN(n1108) );
XOR2_X1 U1119 ( .A(n1148), .B(n1412), .Z(n1324) );
XNOR2_X1 U1120 ( .A(KEYINPUT16), .B(n1145), .ZN(n1412) );
INV_X1 U1121 ( .A(G475), .ZN(n1145) );
INV_X1 U1122 ( .A(n1216), .ZN(n1148) );
NOR2_X1 U1123 ( .A1(n1219), .A2(G902), .ZN(n1216) );
XNOR2_X1 U1124 ( .A(n1413), .B(n1414), .ZN(n1219) );
XNOR2_X1 U1125 ( .A(n1330), .B(n1415), .ZN(n1414) );
XOR2_X1 U1126 ( .A(KEYINPUT19), .B(G122), .Z(n1415) );
INV_X1 U1127 ( .A(G113), .ZN(n1330) );
XOR2_X1 U1128 ( .A(n1416), .B(G104), .Z(n1413) );
NAND2_X1 U1129 ( .A1(KEYINPUT28), .A2(n1417), .ZN(n1416) );
XOR2_X1 U1130 ( .A(n1418), .B(n1419), .Z(n1417) );
XOR2_X1 U1131 ( .A(n1420), .B(n1421), .Z(n1419) );
NOR2_X1 U1132 ( .A1(KEYINPUT53), .A2(n1350), .ZN(n1421) );
XOR2_X1 U1133 ( .A(G146), .B(n1165), .Z(n1350) );
XNOR2_X1 U1134 ( .A(G125), .B(n1301), .ZN(n1165) );
INV_X1 U1135 ( .A(G140), .ZN(n1301) );
NAND2_X1 U1136 ( .A1(n1362), .A2(G214), .ZN(n1420) );
NOR2_X1 U1137 ( .A1(G953), .A2(G237), .ZN(n1362) );
XNOR2_X1 U1138 ( .A(G131), .B(G143), .ZN(n1418) );
XNOR2_X1 U1139 ( .A(n1422), .B(G478), .ZN(n1323) );
NAND2_X1 U1140 ( .A1(n1204), .A2(n1210), .ZN(n1422) );
NAND2_X1 U1141 ( .A1(n1423), .A2(n1424), .ZN(n1210) );
NAND2_X1 U1142 ( .A1(n1425), .A2(n1426), .ZN(n1424) );
XOR2_X1 U1143 ( .A(n1427), .B(KEYINPUT2), .Z(n1423) );
OR2_X1 U1144 ( .A1(n1426), .A2(n1425), .ZN(n1427) );
NOR3_X1 U1145 ( .A1(n1205), .A2(G953), .A3(n1345), .ZN(n1425) );
INV_X1 U1146 ( .A(G217), .ZN(n1345) );
INV_X1 U1147 ( .A(G234), .ZN(n1205) );
XOR2_X1 U1148 ( .A(n1428), .B(n1429), .Z(n1426) );
XNOR2_X1 U1149 ( .A(n1368), .B(n1430), .ZN(n1429) );
XOR2_X1 U1150 ( .A(G134), .B(G122), .Z(n1430) );
INV_X1 U1151 ( .A(G116), .ZN(n1368) );
XNOR2_X1 U1152 ( .A(G107), .B(n1401), .ZN(n1428) );
XOR2_X1 U1153 ( .A(G128), .B(G143), .Z(n1401) );
INV_X1 U1154 ( .A(G902), .ZN(n1204) );
INV_X1 U1155 ( .A(G110), .ZN(n1340) );
endmodule


