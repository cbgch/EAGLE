//Key = 1111101000100001000011000100110011000010011110100000000101111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302;

XNOR2_X1 U717 ( .A(n988), .B(n989), .ZN(G9) );
NAND2_X1 U718 ( .A1(n990), .A2(n991), .ZN(n988) );
OR2_X1 U719 ( .A1(n992), .A2(KEYINPUT5), .ZN(n991) );
NAND3_X1 U720 ( .A1(n993), .A2(n994), .A3(KEYINPUT5), .ZN(n990) );
NOR2_X1 U721 ( .A1(n995), .A2(n996), .ZN(G75) );
NOR3_X1 U722 ( .A1(n997), .A2(G953), .A3(G952), .ZN(n996) );
NOR4_X1 U723 ( .A1(n998), .A2(n999), .A3(n1000), .A4(n997), .ZN(n995) );
AND4_X1 U724 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n997) );
NOR4_X1 U725 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1004) );
XOR2_X1 U726 ( .A(n1009), .B(n1010), .Z(n1007) );
NOR2_X1 U727 ( .A1(G475), .A2(KEYINPUT56), .ZN(n1010) );
XOR2_X1 U728 ( .A(n1011), .B(KEYINPUT47), .Z(n1006) );
NAND2_X1 U729 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND2_X1 U730 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
INV_X1 U731 ( .A(n1016), .ZN(n1001) );
NAND3_X1 U732 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n998) );
NAND4_X1 U733 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1019) );
INV_X1 U734 ( .A(KEYINPUT54), .ZN(n1023) );
NAND2_X1 U735 ( .A1(n1024), .A2(n1025), .ZN(n1021) );
NAND3_X1 U736 ( .A1(n1003), .A2(n1026), .A3(n1027), .ZN(n1025) );
OR2_X1 U737 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NAND2_X1 U738 ( .A1(n1030), .A2(n1031), .ZN(n1024) );
NAND2_X1 U739 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U740 ( .A1(n1027), .A2(n1034), .ZN(n1033) );
NAND2_X1 U741 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U742 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U743 ( .A1(n1003), .A2(n1039), .ZN(n1032) );
NAND3_X1 U744 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
OR3_X1 U745 ( .A1(n1043), .A2(n1044), .A3(KEYINPUT35), .ZN(n1041) );
NAND2_X1 U746 ( .A1(KEYINPUT35), .A2(n1027), .ZN(n1040) );
NAND4_X1 U747 ( .A1(n1003), .A2(n1030), .A3(n1027), .A4(n1045), .ZN(n1017) );
NOR3_X1 U748 ( .A1(n1046), .A2(KEYINPUT54), .A3(n1047), .ZN(n1045) );
INV_X1 U749 ( .A(n1022), .ZN(n1047) );
XOR2_X1 U750 ( .A(n1048), .B(n1049), .Z(G72) );
NOR2_X1 U751 ( .A1(n1050), .A2(n1018), .ZN(n1049) );
NOR2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(n1048) );
NAND2_X1 U754 ( .A1(n1055), .A2(n1018), .ZN(n1054) );
XNOR2_X1 U755 ( .A(n1056), .B(n1057), .ZN(n1055) );
NOR3_X1 U756 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
XNOR2_X1 U757 ( .A(n1061), .B(KEYINPUT52), .ZN(n1060) );
INV_X1 U758 ( .A(n1062), .ZN(n1059) );
NAND3_X1 U759 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1058) );
NAND3_X1 U760 ( .A1(G900), .A2(n1056), .A3(G953), .ZN(n1053) );
XNOR2_X1 U761 ( .A(n1066), .B(n1067), .ZN(n1056) );
NAND2_X1 U762 ( .A1(KEYINPUT15), .A2(n1068), .ZN(n1066) );
XOR2_X1 U763 ( .A(KEYINPUT28), .B(n1069), .Z(n1068) );
XOR2_X1 U764 ( .A(n1070), .B(n1071), .Z(G69) );
NOR2_X1 U765 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U766 ( .A1(G224), .A2(n1018), .ZN(n1072) );
NAND2_X1 U767 ( .A1(KEYINPUT32), .A2(n1074), .ZN(n1070) );
XOR2_X1 U768 ( .A(n1075), .B(n1076), .Z(n1074) );
NOR2_X1 U769 ( .A1(n1077), .A2(G953), .ZN(n1076) );
NOR2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1075) );
XOR2_X1 U771 ( .A(KEYINPUT19), .B(n1073), .Z(n1079) );
XOR2_X1 U772 ( .A(n1080), .B(n1081), .Z(n1078) );
XOR2_X1 U773 ( .A(KEYINPUT53), .B(n1082), .Z(n1081) );
NOR2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(G66) );
XOR2_X1 U775 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND3_X1 U776 ( .A1(n1087), .A2(n1088), .A3(KEYINPUT59), .ZN(n1085) );
NOR2_X1 U777 ( .A1(n1083), .A2(n1089), .ZN(G63) );
XOR2_X1 U778 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND2_X1 U779 ( .A1(n1087), .A2(G478), .ZN(n1090) );
NOR2_X1 U780 ( .A1(n1092), .A2(n1093), .ZN(G60) );
XOR2_X1 U781 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U782 ( .A1(n1096), .A2(KEYINPUT61), .ZN(n1095) );
NOR2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1094) );
NOR2_X1 U784 ( .A1(n1099), .A2(n1100), .ZN(n1092) );
XOR2_X1 U785 ( .A(KEYINPUT9), .B(G952), .Z(n1100) );
XNOR2_X1 U786 ( .A(KEYINPUT63), .B(G953), .ZN(n1099) );
XNOR2_X1 U787 ( .A(G104), .B(n1101), .ZN(G6) );
NOR2_X1 U788 ( .A1(n1083), .A2(n1102), .ZN(G57) );
XOR2_X1 U789 ( .A(n1103), .B(n1104), .Z(n1102) );
XOR2_X1 U790 ( .A(n1105), .B(n1106), .Z(n1104) );
XNOR2_X1 U791 ( .A(n1107), .B(n1108), .ZN(n1106) );
XOR2_X1 U792 ( .A(n1109), .B(n1110), .Z(n1103) );
XNOR2_X1 U793 ( .A(n1111), .B(G101), .ZN(n1110) );
NAND2_X1 U794 ( .A1(n1087), .A2(G472), .ZN(n1109) );
NOR2_X1 U795 ( .A1(n1083), .A2(n1112), .ZN(G54) );
XOR2_X1 U796 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U797 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U798 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
AND3_X1 U799 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1118) );
NOR2_X1 U800 ( .A1(n1122), .A2(n1119), .ZN(n1117) );
INV_X1 U801 ( .A(KEYINPUT43), .ZN(n1119) );
NAND2_X1 U802 ( .A1(KEYINPUT44), .A2(n1123), .ZN(n1115) );
XOR2_X1 U803 ( .A(n1124), .B(n1125), .Z(n1113) );
NAND2_X1 U804 ( .A1(n1087), .A2(G469), .ZN(n1124) );
NOR2_X1 U805 ( .A1(n1083), .A2(n1126), .ZN(G51) );
XOR2_X1 U806 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND2_X1 U807 ( .A1(n1087), .A2(n1014), .ZN(n1127) );
INV_X1 U808 ( .A(n1129), .ZN(n1014) );
INV_X1 U809 ( .A(n1097), .ZN(n1087) );
NAND2_X1 U810 ( .A1(G902), .A2(n1130), .ZN(n1097) );
OR2_X1 U811 ( .A1(n999), .A2(n1000), .ZN(n1130) );
NAND3_X1 U812 ( .A1(n1061), .A2(n1077), .A3(n1131), .ZN(n999) );
AND3_X1 U813 ( .A1(n1062), .A2(n1063), .A3(n1065), .ZN(n1131) );
AND4_X1 U814 ( .A1(n1101), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1077) );
AND4_X1 U815 ( .A1(n992), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1134) );
OR2_X1 U816 ( .A1(n994), .A2(n1042), .ZN(n992) );
NAND4_X1 U817 ( .A1(n1138), .A2(n1029), .A3(n1020), .A4(n1139), .ZN(n994) );
NAND3_X1 U818 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1133) );
NAND2_X1 U819 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
INV_X1 U820 ( .A(KEYINPUT55), .ZN(n1144) );
NAND2_X1 U821 ( .A1(n1046), .A2(KEYINPUT55), .ZN(n1140) );
NOR2_X1 U822 ( .A1(n1143), .A2(n1145), .ZN(n1046) );
NAND3_X1 U823 ( .A1(n1028), .A2(n1020), .A3(n1146), .ZN(n1101) );
AND3_X1 U824 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1061) );
NAND2_X1 U825 ( .A1(n1027), .A2(n1150), .ZN(n1149) );
NAND2_X1 U826 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XNOR2_X1 U827 ( .A(KEYINPUT4), .B(n1153), .ZN(n1152) );
XNOR2_X1 U828 ( .A(n1154), .B(KEYINPUT27), .ZN(n1151) );
NOR2_X1 U829 ( .A1(n1155), .A2(G952), .ZN(n1083) );
XOR2_X1 U830 ( .A(KEYINPUT63), .B(n1018), .Z(n1155) );
XNOR2_X1 U831 ( .A(G146), .B(n1147), .ZN(G48) );
NAND3_X1 U832 ( .A1(n1028), .A2(n993), .A3(n1156), .ZN(n1147) );
XNOR2_X1 U833 ( .A(G143), .B(n1148), .ZN(G45) );
NAND4_X1 U834 ( .A1(n1157), .A2(n993), .A3(n1158), .A4(n1016), .ZN(n1148) );
XNOR2_X1 U835 ( .A(G140), .B(n1159), .ZN(G42) );
NOR2_X1 U836 ( .A1(n1160), .A2(KEYINPUT30), .ZN(n1159) );
NOR2_X1 U837 ( .A1(n1161), .A2(n1153), .ZN(n1160) );
NAND2_X1 U838 ( .A1(n1162), .A2(n1138), .ZN(n1153) );
INV_X1 U839 ( .A(n1027), .ZN(n1161) );
XNOR2_X1 U840 ( .A(G137), .B(n1163), .ZN(G39) );
NAND2_X1 U841 ( .A1(n1154), .A2(n1027), .ZN(n1163) );
AND2_X1 U842 ( .A1(n1156), .A2(n1030), .ZN(n1154) );
XNOR2_X1 U843 ( .A(G134), .B(n1062), .ZN(G36) );
NAND3_X1 U844 ( .A1(n1027), .A2(n1029), .A3(n1157), .ZN(n1062) );
XNOR2_X1 U845 ( .A(G131), .B(n1065), .ZN(G33) );
NAND3_X1 U846 ( .A1(n1027), .A2(n1028), .A3(n1157), .ZN(n1065) );
NOR3_X1 U847 ( .A1(n1035), .A2(n1164), .A3(n1165), .ZN(n1157) );
INV_X1 U848 ( .A(n1138), .ZN(n1035) );
NOR2_X1 U849 ( .A1(n1044), .A2(n1005), .ZN(n1027) );
INV_X1 U850 ( .A(n1043), .ZN(n1005) );
XNOR2_X1 U851 ( .A(G128), .B(n1063), .ZN(G30) );
NAND3_X1 U852 ( .A1(n993), .A2(n1029), .A3(n1156), .ZN(n1063) );
AND4_X1 U853 ( .A1(n1166), .A2(n1138), .A3(n1167), .A4(n1168), .ZN(n1156) );
XOR2_X1 U854 ( .A(G101), .B(n1169), .Z(G3) );
NOR2_X1 U855 ( .A1(n1165), .A2(n1170), .ZN(n1169) );
XNOR2_X1 U856 ( .A(n1171), .B(n1172), .ZN(G27) );
NAND2_X1 U857 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
NAND4_X1 U858 ( .A1(n1003), .A2(n1028), .A3(n1175), .A4(n1176), .ZN(n1174) );
INV_X1 U859 ( .A(KEYINPUT20), .ZN(n1176) );
NOR3_X1 U860 ( .A1(n1042), .A2(n1143), .A3(n1164), .ZN(n1175) );
INV_X1 U861 ( .A(n1168), .ZN(n1164) );
NAND2_X1 U862 ( .A1(n1000), .A2(KEYINPUT20), .ZN(n1173) );
INV_X1 U863 ( .A(n1064), .ZN(n1000) );
NAND3_X1 U864 ( .A1(n1003), .A2(n993), .A3(n1162), .ZN(n1064) );
AND3_X1 U865 ( .A1(n1028), .A2(n1168), .A3(n1143), .ZN(n1162) );
NAND2_X1 U866 ( .A1(n1177), .A2(n1178), .ZN(n1168) );
NAND4_X1 U867 ( .A1(G953), .A2(G902), .A3(n1022), .A4(n1052), .ZN(n1178) );
INV_X1 U868 ( .A(G900), .ZN(n1052) );
XOR2_X1 U869 ( .A(n1132), .B(n1179), .Z(G24) );
XOR2_X1 U870 ( .A(KEYINPUT33), .B(G122), .Z(n1179) );
NAND4_X1 U871 ( .A1(n1180), .A2(n1020), .A3(n1158), .A4(n1016), .ZN(n1132) );
NOR2_X1 U872 ( .A1(n1167), .A2(n1166), .ZN(n1020) );
XOR2_X1 U873 ( .A(n1137), .B(n1181), .Z(G21) );
XNOR2_X1 U874 ( .A(KEYINPUT6), .B(n1182), .ZN(n1181) );
NAND4_X1 U875 ( .A1(n1166), .A2(n1180), .A3(n1030), .A4(n1167), .ZN(n1137) );
XNOR2_X1 U876 ( .A(G116), .B(n1136), .ZN(G18) );
NAND3_X1 U877 ( .A1(n1145), .A2(n1029), .A3(n1180), .ZN(n1136) );
AND2_X1 U878 ( .A1(n1183), .A2(n1016), .ZN(n1029) );
XNOR2_X1 U879 ( .A(KEYINPUT14), .B(n1158), .ZN(n1183) );
XNOR2_X1 U880 ( .A(G113), .B(n1135), .ZN(G15) );
NAND3_X1 U881 ( .A1(n1145), .A2(n1028), .A3(n1180), .ZN(n1135) );
AND3_X1 U882 ( .A1(n993), .A2(n1139), .A3(n1003), .ZN(n1180) );
NOR2_X1 U883 ( .A1(n1184), .A2(n1037), .ZN(n1003) );
INV_X1 U884 ( .A(n1165), .ZN(n1145) );
NAND2_X1 U885 ( .A1(n1166), .A2(n1002), .ZN(n1165) );
XOR2_X1 U886 ( .A(n1185), .B(n1186), .Z(G12) );
NAND2_X1 U887 ( .A1(KEYINPUT29), .A2(G110), .ZN(n1186) );
NAND2_X1 U888 ( .A1(n1142), .A2(n1143), .ZN(n1185) );
NOR2_X1 U889 ( .A1(n1002), .A2(n1166), .ZN(n1143) );
XNOR2_X1 U890 ( .A(n1008), .B(KEYINPUT3), .ZN(n1166) );
XNOR2_X1 U891 ( .A(n1187), .B(n1188), .ZN(n1008) );
XOR2_X1 U892 ( .A(KEYINPUT8), .B(G472), .Z(n1188) );
NAND3_X1 U893 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1187) );
NAND2_X1 U894 ( .A1(KEYINPUT57), .A2(n1192), .ZN(n1190) );
XOR2_X1 U895 ( .A(n1193), .B(n1194), .Z(n1192) );
NAND3_X1 U896 ( .A1(n1194), .A2(n1193), .A3(n1195), .ZN(n1189) );
INV_X1 U897 ( .A(KEYINPUT57), .ZN(n1195) );
XOR2_X1 U898 ( .A(G101), .B(n1196), .Z(n1193) );
NOR2_X1 U899 ( .A1(n1111), .A2(KEYINPUT51), .ZN(n1196) );
AND3_X1 U900 ( .A1(n1197), .A2(n1018), .A3(G210), .ZN(n1111) );
XNOR2_X1 U901 ( .A(n1198), .B(n1199), .ZN(n1194) );
XNOR2_X1 U902 ( .A(n1200), .B(KEYINPUT31), .ZN(n1199) );
NAND2_X1 U903 ( .A1(KEYINPUT41), .A2(n1108), .ZN(n1200) );
XOR2_X1 U904 ( .A(n1105), .B(n1201), .Z(n1198) );
NOR2_X1 U905 ( .A1(KEYINPUT49), .A2(n1107), .ZN(n1201) );
XNOR2_X1 U906 ( .A(n1202), .B(n1203), .ZN(n1107) );
XNOR2_X1 U907 ( .A(KEYINPUT36), .B(n1182), .ZN(n1203) );
XNOR2_X1 U908 ( .A(G116), .B(n1204), .ZN(n1202) );
INV_X1 U909 ( .A(n1167), .ZN(n1002) );
XNOR2_X1 U910 ( .A(n1205), .B(n1088), .ZN(n1167) );
AND2_X1 U911 ( .A1(G217), .A2(n1206), .ZN(n1088) );
NAND2_X1 U912 ( .A1(n1191), .A2(n1086), .ZN(n1205) );
XNOR2_X1 U913 ( .A(n1207), .B(n1208), .ZN(n1086) );
XOR2_X1 U914 ( .A(n1209), .B(n1210), .Z(n1208) );
XNOR2_X1 U915 ( .A(n1211), .B(n1212), .ZN(n1210) );
NAND2_X1 U916 ( .A1(KEYINPUT46), .A2(n1213), .ZN(n1212) );
NAND2_X1 U917 ( .A1(KEYINPUT25), .A2(n1214), .ZN(n1211) );
NAND2_X1 U918 ( .A1(n1215), .A2(G221), .ZN(n1209) );
XOR2_X1 U919 ( .A(n1216), .B(n1217), .Z(n1207) );
XNOR2_X1 U920 ( .A(G146), .B(n1182), .ZN(n1217) );
XNOR2_X1 U921 ( .A(G110), .B(n1218), .ZN(n1216) );
NOR2_X1 U922 ( .A1(KEYINPUT24), .A2(n1219), .ZN(n1218) );
INV_X1 U923 ( .A(n1170), .ZN(n1142) );
NAND2_X1 U924 ( .A1(n1146), .A2(n1030), .ZN(n1170) );
NAND2_X1 U925 ( .A1(n1220), .A2(n1221), .ZN(n1030) );
OR3_X1 U926 ( .A1(n1158), .A2(n1016), .A3(KEYINPUT14), .ZN(n1221) );
INV_X1 U927 ( .A(n1222), .ZN(n1158) );
NAND2_X1 U928 ( .A1(KEYINPUT14), .A2(n1028), .ZN(n1220) );
NOR2_X1 U929 ( .A1(n1016), .A2(n1222), .ZN(n1028) );
XOR2_X1 U930 ( .A(n1223), .B(n1009), .Z(n1222) );
NAND2_X1 U931 ( .A1(n1096), .A2(n1191), .ZN(n1009) );
AND3_X1 U932 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1096) );
NAND2_X1 U933 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
OR2_X1 U934 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
OR4_X1 U935 ( .A1(n1227), .A2(n1230), .A3(n1229), .A4(KEYINPUT62), .ZN(n1225) );
INV_X1 U936 ( .A(KEYINPUT21), .ZN(n1229) );
XOR2_X1 U937 ( .A(G104), .B(n1231), .Z(n1227) );
XNOR2_X1 U938 ( .A(G122), .B(n1232), .ZN(n1231) );
INV_X1 U939 ( .A(G113), .ZN(n1232) );
NAND2_X1 U940 ( .A1(n1230), .A2(KEYINPUT62), .ZN(n1224) );
XNOR2_X1 U941 ( .A(n1233), .B(n1234), .ZN(n1230) );
XOR2_X1 U942 ( .A(G143), .B(n1235), .Z(n1234) );
XOR2_X1 U943 ( .A(KEYINPUT38), .B(G146), .Z(n1235) );
XNOR2_X1 U944 ( .A(n1236), .B(n1219), .ZN(n1233) );
XNOR2_X1 U945 ( .A(n1067), .B(KEYINPUT17), .ZN(n1219) );
XNOR2_X1 U946 ( .A(G125), .B(n1237), .ZN(n1067) );
INV_X1 U947 ( .A(G140), .ZN(n1237) );
XOR2_X1 U948 ( .A(n1238), .B(n1239), .Z(n1236) );
NOR2_X1 U949 ( .A1(G131), .A2(KEYINPUT40), .ZN(n1239) );
NAND3_X1 U950 ( .A1(n1197), .A2(n1018), .A3(G214), .ZN(n1238) );
NAND2_X1 U951 ( .A1(KEYINPUT10), .A2(n1098), .ZN(n1223) );
INV_X1 U952 ( .A(G475), .ZN(n1098) );
XNOR2_X1 U953 ( .A(n1240), .B(G478), .ZN(n1016) );
NAND2_X1 U954 ( .A1(n1241), .A2(n1191), .ZN(n1240) );
XOR2_X1 U955 ( .A(n1091), .B(KEYINPUT18), .Z(n1241) );
XOR2_X1 U956 ( .A(n1242), .B(n1243), .Z(n1091) );
XOR2_X1 U957 ( .A(n1244), .B(n1245), .Z(n1243) );
NAND3_X1 U958 ( .A1(n1215), .A2(n1246), .A3(KEYINPUT42), .ZN(n1245) );
XOR2_X1 U959 ( .A(KEYINPUT7), .B(G217), .Z(n1246) );
AND2_X1 U960 ( .A1(G234), .A2(n1018), .ZN(n1215) );
NAND3_X1 U961 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(n1244) );
NAND2_X1 U962 ( .A1(G128), .A2(n1250), .ZN(n1249) );
NAND2_X1 U963 ( .A1(KEYINPUT37), .A2(n1251), .ZN(n1248) );
NAND2_X1 U964 ( .A1(n1252), .A2(n1214), .ZN(n1251) );
XNOR2_X1 U965 ( .A(KEYINPUT50), .B(n1250), .ZN(n1252) );
NAND2_X1 U966 ( .A1(n1253), .A2(n1254), .ZN(n1247) );
INV_X1 U967 ( .A(KEYINPUT37), .ZN(n1254) );
NAND2_X1 U968 ( .A1(n1255), .A2(n1256), .ZN(n1253) );
OR3_X1 U969 ( .A1(n1250), .A2(G128), .A3(KEYINPUT50), .ZN(n1256) );
NAND2_X1 U970 ( .A1(KEYINPUT50), .A2(n1250), .ZN(n1255) );
XOR2_X1 U971 ( .A(G143), .B(KEYINPUT1), .Z(n1250) );
XOR2_X1 U972 ( .A(n1257), .B(G134), .Z(n1242) );
NAND2_X1 U973 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NAND2_X1 U974 ( .A1(G107), .A2(n1260), .ZN(n1259) );
XOR2_X1 U975 ( .A(n1261), .B(KEYINPUT16), .Z(n1258) );
OR2_X1 U976 ( .A1(n1260), .A2(G107), .ZN(n1261) );
XOR2_X1 U977 ( .A(G116), .B(n1262), .Z(n1260) );
XOR2_X1 U978 ( .A(KEYINPUT39), .B(G122), .Z(n1262) );
AND3_X1 U979 ( .A1(n1138), .A2(n1139), .A3(n993), .ZN(n1146) );
INV_X1 U980 ( .A(n1042), .ZN(n993) );
NAND2_X1 U981 ( .A1(n1044), .A2(n1043), .ZN(n1042) );
NAND2_X1 U982 ( .A1(G214), .A2(n1263), .ZN(n1043) );
NAND3_X1 U983 ( .A1(n1264), .A2(n1265), .A3(n1012), .ZN(n1044) );
NAND2_X1 U984 ( .A1(n1266), .A2(n1129), .ZN(n1012) );
NAND2_X1 U985 ( .A1(KEYINPUT26), .A2(n1129), .ZN(n1265) );
OR3_X1 U986 ( .A1(n1266), .A2(KEYINPUT26), .A3(n1129), .ZN(n1264) );
NAND2_X1 U987 ( .A1(G210), .A2(n1263), .ZN(n1129) );
NAND2_X1 U988 ( .A1(n1197), .A2(n1267), .ZN(n1263) );
INV_X1 U989 ( .A(G237), .ZN(n1197) );
INV_X1 U990 ( .A(n1015), .ZN(n1266) );
NAND2_X1 U991 ( .A1(n1128), .A2(n1191), .ZN(n1015) );
XNOR2_X1 U992 ( .A(n1268), .B(n1269), .ZN(n1128) );
XOR2_X1 U993 ( .A(n1080), .B(n1105), .Z(n1269) );
NAND2_X1 U994 ( .A1(n1270), .A2(n1271), .ZN(n1105) );
OR2_X1 U995 ( .A1(n1272), .A2(KEYINPUT12), .ZN(n1271) );
NAND3_X1 U996 ( .A1(G128), .A2(n1273), .A3(KEYINPUT12), .ZN(n1270) );
XNOR2_X1 U997 ( .A(G110), .B(G122), .ZN(n1080) );
XOR2_X1 U998 ( .A(n1274), .B(n1275), .Z(n1268) );
AND2_X1 U999 ( .A1(n1018), .A2(G224), .ZN(n1275) );
XNOR2_X1 U1000 ( .A(n1276), .B(n1172), .ZN(n1274) );
INV_X1 U1001 ( .A(G125), .ZN(n1172) );
NAND2_X1 U1002 ( .A1(KEYINPUT58), .A2(n1082), .ZN(n1276) );
XNOR2_X1 U1003 ( .A(n1277), .B(n1278), .ZN(n1082) );
XOR2_X1 U1004 ( .A(n1279), .B(n1280), .Z(n1278) );
NOR2_X1 U1005 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XOR2_X1 U1006 ( .A(KEYINPUT22), .B(n1283), .Z(n1282) );
NOR2_X1 U1007 ( .A1(n1204), .A2(n1284), .ZN(n1283) );
AND2_X1 U1008 ( .A1(n1284), .A2(n1204), .ZN(n1281) );
XOR2_X1 U1009 ( .A(G113), .B(KEYINPUT13), .Z(n1204) );
NAND3_X1 U1010 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(n1284) );
NAND2_X1 U1011 ( .A1(KEYINPUT45), .A2(G119), .ZN(n1287) );
NAND3_X1 U1012 ( .A1(n1182), .A2(n1288), .A3(G116), .ZN(n1286) );
NAND2_X1 U1013 ( .A1(n1289), .A2(n1290), .ZN(n1285) );
INV_X1 U1014 ( .A(G116), .ZN(n1290) );
NAND2_X1 U1015 ( .A1(n1291), .A2(n1288), .ZN(n1289) );
INV_X1 U1016 ( .A(KEYINPUT45), .ZN(n1288) );
XNOR2_X1 U1017 ( .A(KEYINPUT2), .B(n1182), .ZN(n1291) );
INV_X1 U1018 ( .A(G119), .ZN(n1182) );
NOR2_X1 U1019 ( .A1(KEYINPUT11), .A2(G101), .ZN(n1279) );
XNOR2_X1 U1020 ( .A(G104), .B(G107), .ZN(n1277) );
NAND2_X1 U1021 ( .A1(n1177), .A2(n1292), .ZN(n1139) );
NAND3_X1 U1022 ( .A1(G902), .A2(n1022), .A3(n1073), .ZN(n1292) );
NOR2_X1 U1023 ( .A1(G898), .A2(n1018), .ZN(n1073) );
NAND3_X1 U1024 ( .A1(n1022), .A2(n1018), .A3(G952), .ZN(n1177) );
INV_X1 U1025 ( .A(G953), .ZN(n1018) );
NAND2_X1 U1026 ( .A1(G237), .A2(G234), .ZN(n1022) );
NOR2_X1 U1027 ( .A1(n1038), .A2(n1037), .ZN(n1138) );
AND2_X1 U1028 ( .A1(G221), .A2(n1206), .ZN(n1037) );
NAND2_X1 U1029 ( .A1(G234), .A2(n1267), .ZN(n1206) );
INV_X1 U1030 ( .A(G902), .ZN(n1267) );
INV_X1 U1031 ( .A(n1184), .ZN(n1038) );
XNOR2_X1 U1032 ( .A(n1293), .B(G469), .ZN(n1184) );
NAND2_X1 U1033 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
XOR2_X1 U1034 ( .A(n1191), .B(KEYINPUT23), .Z(n1295) );
XNOR2_X1 U1035 ( .A(G902), .B(KEYINPUT34), .ZN(n1191) );
XOR2_X1 U1036 ( .A(n1296), .B(n1122), .Z(n1294) );
XNOR2_X1 U1037 ( .A(n1120), .B(n1121), .ZN(n1122) );
XOR2_X1 U1038 ( .A(G140), .B(KEYINPUT48), .Z(n1121) );
INV_X1 U1039 ( .A(G110), .ZN(n1120) );
XOR2_X1 U1040 ( .A(n1297), .B(n1123), .Z(n1296) );
XNOR2_X1 U1041 ( .A(n1298), .B(n1299), .ZN(n1123) );
XNOR2_X1 U1042 ( .A(n1300), .B(G101), .ZN(n1299) );
INV_X1 U1043 ( .A(G104), .ZN(n1300) );
XOR2_X1 U1044 ( .A(n1301), .B(n1069), .Z(n1298) );
XNOR2_X1 U1045 ( .A(n1272), .B(n1108), .ZN(n1069) );
XOR2_X1 U1046 ( .A(G131), .B(n1302), .Z(n1108) );
XNOR2_X1 U1047 ( .A(n1213), .B(G134), .ZN(n1302) );
INV_X1 U1048 ( .A(G137), .ZN(n1213) );
XOR2_X1 U1049 ( .A(n1214), .B(n1273), .Z(n1272) );
XOR2_X1 U1050 ( .A(G143), .B(G146), .Z(n1273) );
INV_X1 U1051 ( .A(G128), .ZN(n1214) );
NAND2_X1 U1052 ( .A1(KEYINPUT60), .A2(n989), .ZN(n1301) );
INV_X1 U1053 ( .A(G107), .ZN(n989) );
NAND2_X1 U1054 ( .A1(KEYINPUT0), .A2(n1125), .ZN(n1297) );
NOR2_X1 U1055 ( .A1(n1051), .A2(G953), .ZN(n1125) );
INV_X1 U1056 ( .A(G227), .ZN(n1051) );
endmodule


