//Key = 0010101000101101011010110100101010110111010000000101001110001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;

XNOR2_X1 U787 ( .A(G107), .B(n1090), .ZN(G9) );
NAND3_X1 U788 ( .A1(n1091), .A2(n1092), .A3(KEYINPUT2), .ZN(n1090) );
NOR2_X1 U789 ( .A1(n1093), .A2(n1094), .ZN(G75) );
NOR4_X1 U790 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1094) );
NOR2_X1 U791 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NOR2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
XOR2_X1 U793 ( .A(n1103), .B(KEYINPUT56), .Z(n1102) );
NAND3_X1 U794 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1103) );
NOR3_X1 U795 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1106) );
NOR4_X1 U796 ( .A1(n1110), .A2(n1107), .A3(n1111), .A4(n1112), .ZN(n1101) );
INV_X1 U797 ( .A(n1104), .ZN(n1112) );
NOR2_X1 U798 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
NAND3_X1 U799 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1095) );
NAND3_X1 U800 ( .A1(n1118), .A2(n1119), .A3(n1105), .ZN(n1117) );
NAND2_X1 U801 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND4_X1 U802 ( .A1(n1108), .A2(n1104), .A3(n1109), .A4(n1122), .ZN(n1121) );
INV_X1 U803 ( .A(n1123), .ZN(n1109) );
NAND2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1120) );
NAND3_X1 U805 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1125) );
NAND2_X1 U806 ( .A1(n1122), .A2(n1091), .ZN(n1128) );
NAND2_X1 U807 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
XNOR2_X1 U808 ( .A(KEYINPUT31), .B(n1100), .ZN(n1130) );
NAND2_X1 U809 ( .A1(n1104), .A2(n1131), .ZN(n1126) );
NAND2_X1 U810 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NAND2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
INV_X1 U812 ( .A(n1107), .ZN(n1118) );
AND3_X1 U813 ( .A1(n1115), .A2(n1116), .A3(n1136), .ZN(n1093) );
NAND4_X1 U814 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1115) );
NOR4_X1 U815 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1140) );
NOR2_X1 U816 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NOR2_X1 U817 ( .A1(G902), .A2(n1147), .ZN(n1145) );
NOR2_X1 U818 ( .A1(n1100), .A2(n1111), .ZN(n1139) );
XOR2_X1 U819 ( .A(n1148), .B(n1149), .Z(n1138) );
NAND2_X1 U820 ( .A1(KEYINPUT32), .A2(n1150), .ZN(n1149) );
INV_X1 U821 ( .A(n1151), .ZN(n1137) );
XOR2_X1 U822 ( .A(n1152), .B(n1153), .Z(G72) );
XOR2_X1 U823 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U824 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U825 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U826 ( .A(n1160), .B(KEYINPUT63), .Z(n1158) );
NAND2_X1 U827 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U828 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U829 ( .A(KEYINPUT25), .B(n1165), .Z(n1161) );
NOR2_X1 U830 ( .A1(n1164), .A2(n1163), .ZN(n1165) );
XNOR2_X1 U831 ( .A(n1166), .B(G131), .ZN(n1163) );
NAND2_X1 U832 ( .A1(KEYINPUT12), .A2(n1167), .ZN(n1166) );
NAND2_X1 U833 ( .A1(n1168), .A2(n1116), .ZN(n1154) );
XOR2_X1 U834 ( .A(n1096), .B(KEYINPUT44), .Z(n1168) );
NAND2_X1 U835 ( .A1(G953), .A2(n1169), .ZN(n1152) );
NAND2_X1 U836 ( .A1(G900), .A2(G227), .ZN(n1169) );
XOR2_X1 U837 ( .A(n1170), .B(n1171), .Z(G69) );
NOR2_X1 U838 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NAND3_X1 U839 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1170) );
INV_X1 U840 ( .A(n1172), .ZN(n1176) );
NAND2_X1 U841 ( .A1(G953), .A2(n1177), .ZN(n1175) );
NAND2_X1 U842 ( .A1(n1098), .A2(n1116), .ZN(n1174) );
NOR2_X1 U843 ( .A1(n1178), .A2(n1179), .ZN(G66) );
XNOR2_X1 U844 ( .A(n1180), .B(n1181), .ZN(n1179) );
NOR2_X1 U845 ( .A1(n1148), .A2(n1182), .ZN(n1180) );
NOR2_X1 U846 ( .A1(n1178), .A2(n1183), .ZN(G63) );
NOR2_X1 U847 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
XOR2_X1 U848 ( .A(KEYINPUT59), .B(n1186), .Z(n1185) );
NOR3_X1 U849 ( .A1(n1182), .A2(n1187), .A3(n1188), .ZN(n1186) );
XNOR2_X1 U850 ( .A(n1189), .B(KEYINPUT5), .ZN(n1187) );
NOR2_X1 U851 ( .A1(n1189), .A2(n1190), .ZN(n1184) );
NOR2_X1 U852 ( .A1(n1188), .A2(n1182), .ZN(n1190) );
INV_X1 U853 ( .A(G478), .ZN(n1188) );
NOR2_X1 U854 ( .A1(n1191), .A2(n1192), .ZN(G60) );
XOR2_X1 U855 ( .A(n1147), .B(n1193), .Z(n1192) );
XOR2_X1 U856 ( .A(KEYINPUT52), .B(n1194), .Z(n1193) );
NOR2_X1 U857 ( .A1(n1146), .A2(n1182), .ZN(n1194) );
INV_X1 U858 ( .A(G475), .ZN(n1146) );
NOR2_X1 U859 ( .A1(n1195), .A2(n1196), .ZN(n1191) );
XNOR2_X1 U860 ( .A(KEYINPUT45), .B(n1136), .ZN(n1196) );
XNOR2_X1 U861 ( .A(KEYINPUT24), .B(G953), .ZN(n1195) );
XNOR2_X1 U862 ( .A(G104), .B(n1197), .ZN(G6) );
NAND2_X1 U863 ( .A1(n1092), .A2(n1198), .ZN(n1197) );
XNOR2_X1 U864 ( .A(KEYINPUT53), .B(n1199), .ZN(n1198) );
NOR3_X1 U865 ( .A1(n1178), .A2(n1200), .A3(n1201), .ZN(G57) );
NOR2_X1 U866 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
INV_X1 U867 ( .A(n1204), .ZN(n1203) );
XNOR2_X1 U868 ( .A(n1205), .B(KEYINPUT42), .ZN(n1202) );
NOR2_X1 U869 ( .A1(n1204), .A2(n1206), .ZN(n1200) );
XNOR2_X1 U870 ( .A(KEYINPUT47), .B(n1207), .ZN(n1206) );
INV_X1 U871 ( .A(n1205), .ZN(n1207) );
XNOR2_X1 U872 ( .A(n1208), .B(n1209), .ZN(n1205) );
XOR2_X1 U873 ( .A(n1210), .B(n1211), .Z(n1209) );
NOR2_X1 U874 ( .A1(KEYINPUT14), .A2(n1212), .ZN(n1211) );
NOR2_X1 U875 ( .A1(n1213), .A2(n1182), .ZN(n1210) );
NOR2_X1 U876 ( .A1(n1178), .A2(n1214), .ZN(G54) );
XOR2_X1 U877 ( .A(n1215), .B(n1216), .Z(n1214) );
XNOR2_X1 U878 ( .A(n1164), .B(n1217), .ZN(n1216) );
XOR2_X1 U879 ( .A(n1218), .B(n1219), .Z(n1215) );
NOR2_X1 U880 ( .A1(n1220), .A2(n1182), .ZN(n1218) );
NOR2_X1 U881 ( .A1(n1178), .A2(n1221), .ZN(G51) );
XOR2_X1 U882 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR2_X1 U883 ( .A1(n1182), .A2(n1224), .ZN(n1223) );
XOR2_X1 U884 ( .A(KEYINPUT55), .B(n1225), .Z(n1224) );
NAND2_X1 U885 ( .A1(G902), .A2(n1226), .ZN(n1182) );
OR2_X1 U886 ( .A1(n1096), .A2(n1098), .ZN(n1226) );
NAND4_X1 U887 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1098) );
NOR4_X1 U888 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1230) );
NAND2_X1 U889 ( .A1(n1092), .A2(n1235), .ZN(n1229) );
NAND2_X1 U890 ( .A1(n1199), .A2(n1236), .ZN(n1235) );
AND2_X1 U891 ( .A1(n1237), .A2(n1105), .ZN(n1092) );
NAND4_X1 U892 ( .A1(n1238), .A2(n1239), .A3(n1105), .A4(n1240), .ZN(n1228) );
NOR2_X1 U893 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
OR2_X1 U894 ( .A1(n1243), .A2(KEYINPUT0), .ZN(n1239) );
NAND2_X1 U895 ( .A1(KEYINPUT0), .A2(n1244), .ZN(n1238) );
NAND2_X1 U896 ( .A1(n1245), .A2(n1111), .ZN(n1244) );
INV_X1 U897 ( .A(n1124), .ZN(n1111) );
NAND3_X1 U898 ( .A1(n1243), .A2(n1104), .A3(n1246), .ZN(n1227) );
XNOR2_X1 U899 ( .A(KEYINPUT34), .B(n1247), .ZN(n1246) );
NAND4_X1 U900 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1096) );
NOR4_X1 U901 ( .A1(n1252), .A2(n1253), .A3(n1254), .A4(n1255), .ZN(n1251) );
NOR3_X1 U902 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1250) );
NOR3_X1 U903 ( .A1(n1259), .A2(n1260), .A3(n1100), .ZN(n1258) );
INV_X1 U904 ( .A(KEYINPUT29), .ZN(n1259) );
NOR2_X1 U905 ( .A1(KEYINPUT29), .A2(n1261), .ZN(n1257) );
NOR3_X1 U906 ( .A1(n1262), .A2(n1132), .A3(n1263), .ZN(n1256) );
XNOR2_X1 U907 ( .A(n1264), .B(KEYINPUT38), .ZN(n1262) );
NAND2_X1 U908 ( .A1(n1265), .A2(KEYINPUT17), .ZN(n1222) );
XOR2_X1 U909 ( .A(n1266), .B(n1173), .Z(n1265) );
NAND3_X1 U910 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(n1266) );
INV_X1 U911 ( .A(n1270), .ZN(n1269) );
NAND2_X1 U912 ( .A1(n1271), .A2(n1272), .ZN(n1268) );
INV_X1 U913 ( .A(KEYINPUT60), .ZN(n1272) );
XNOR2_X1 U914 ( .A(n1273), .B(n1274), .ZN(n1271) );
NOR2_X1 U915 ( .A1(G125), .A2(n1275), .ZN(n1274) );
NAND2_X1 U916 ( .A1(KEYINPUT60), .A2(n1276), .ZN(n1267) );
AND2_X1 U917 ( .A1(n1277), .A2(n1136), .ZN(n1178) );
INV_X1 U918 ( .A(G952), .ZN(n1136) );
XNOR2_X1 U919 ( .A(KEYINPUT24), .B(n1116), .ZN(n1277) );
XNOR2_X1 U920 ( .A(n1278), .B(n1279), .ZN(G48) );
NOR3_X1 U921 ( .A1(n1132), .A2(KEYINPUT33), .A3(n1280), .ZN(n1279) );
XOR2_X1 U922 ( .A(n1281), .B(KEYINPUT48), .Z(n1280) );
NAND2_X1 U923 ( .A1(n1129), .A2(n1282), .ZN(n1281) );
XNOR2_X1 U924 ( .A(G143), .B(n1249), .ZN(G45) );
NAND4_X1 U925 ( .A1(n1283), .A2(n1284), .A3(n1114), .A4(n1285), .ZN(n1249) );
NOR2_X1 U926 ( .A1(n1132), .A2(n1286), .ZN(n1285) );
INV_X1 U927 ( .A(n1287), .ZN(n1132) );
XNOR2_X1 U928 ( .A(n1288), .B(n1255), .ZN(G42) );
AND3_X1 U929 ( .A1(n1113), .A2(n1122), .A3(n1289), .ZN(n1255) );
XNOR2_X1 U930 ( .A(G137), .B(n1290), .ZN(G39) );
NOR2_X1 U931 ( .A1(n1291), .A2(KEYINPUT3), .ZN(n1290) );
INV_X1 U932 ( .A(n1261), .ZN(n1291) );
NAND2_X1 U933 ( .A1(n1260), .A2(n1122), .ZN(n1261) );
INV_X1 U934 ( .A(n1100), .ZN(n1122) );
AND2_X1 U935 ( .A1(n1104), .A2(n1282), .ZN(n1260) );
XOR2_X1 U936 ( .A(n1254), .B(n1292), .Z(G36) );
NOR2_X1 U937 ( .A1(KEYINPUT58), .A2(n1293), .ZN(n1292) );
NOR4_X1 U938 ( .A1(n1286), .A2(n1100), .A3(n1236), .A4(n1294), .ZN(n1254) );
XOR2_X1 U939 ( .A(G131), .B(n1253), .Z(G33) );
NOR3_X1 U940 ( .A1(n1100), .A2(n1294), .A3(n1263), .ZN(n1253) );
INV_X1 U941 ( .A(n1289), .ZN(n1263) );
NOR2_X1 U942 ( .A1(n1199), .A2(n1286), .ZN(n1289) );
NAND2_X1 U943 ( .A1(n1135), .A2(n1295), .ZN(n1100) );
XNOR2_X1 U944 ( .A(G128), .B(n1296), .ZN(G30) );
NOR2_X1 U945 ( .A1(n1252), .A2(KEYINPUT11), .ZN(n1296) );
AND3_X1 U946 ( .A1(n1091), .A2(n1287), .A3(n1282), .ZN(n1252) );
NOR2_X1 U947 ( .A1(n1286), .A2(n1264), .ZN(n1282) );
INV_X1 U948 ( .A(n1247), .ZN(n1264) );
NAND3_X1 U949 ( .A1(n1297), .A2(n1298), .A3(n1123), .ZN(n1286) );
XNOR2_X1 U950 ( .A(G101), .B(n1299), .ZN(G3) );
NAND2_X1 U951 ( .A1(KEYINPUT6), .A2(n1234), .ZN(n1299) );
AND3_X1 U952 ( .A1(n1237), .A2(n1114), .A3(n1104), .ZN(n1234) );
XNOR2_X1 U953 ( .A(G125), .B(n1248), .ZN(G27) );
NAND4_X1 U954 ( .A1(n1129), .A2(n1113), .A3(n1300), .A4(n1124), .ZN(n1248) );
AND2_X1 U955 ( .A1(n1297), .A2(n1287), .ZN(n1300) );
NAND2_X1 U956 ( .A1(n1107), .A2(n1301), .ZN(n1297) );
NAND3_X1 U957 ( .A1(G902), .A2(n1302), .A3(n1156), .ZN(n1301) );
NOR2_X1 U958 ( .A1(n1116), .A2(G900), .ZN(n1156) );
XNOR2_X1 U959 ( .A(G122), .B(n1303), .ZN(G24) );
NAND4_X1 U960 ( .A1(n1243), .A2(n1105), .A3(n1283), .A4(n1284), .ZN(n1303) );
NAND3_X1 U961 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(G21) );
NAND2_X1 U962 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
INV_X1 U963 ( .A(KEYINPUT4), .ZN(n1308) );
NAND2_X1 U964 ( .A1(G119), .A2(n1309), .ZN(n1307) );
NAND3_X1 U965 ( .A1(KEYINPUT4), .A2(n1310), .A3(G119), .ZN(n1305) );
OR2_X1 U966 ( .A1(n1309), .A2(KEYINPUT40), .ZN(n1310) );
OR3_X1 U967 ( .A1(n1309), .A2(KEYINPUT40), .A3(G119), .ZN(n1304) );
NAND3_X1 U968 ( .A1(n1243), .A2(n1247), .A3(n1311), .ZN(n1309) );
XNOR2_X1 U969 ( .A(n1104), .B(KEYINPUT15), .ZN(n1311) );
NAND2_X1 U970 ( .A1(n1312), .A2(n1313), .ZN(n1247) );
NAND3_X1 U971 ( .A1(n1151), .A2(n1314), .A3(n1315), .ZN(n1313) );
NAND2_X1 U972 ( .A1(KEYINPUT26), .A2(n1113), .ZN(n1312) );
INV_X1 U973 ( .A(n1316), .ZN(n1243) );
XNOR2_X1 U974 ( .A(n1317), .B(n1233), .ZN(G18) );
NOR3_X1 U975 ( .A1(n1236), .A2(n1294), .A3(n1316), .ZN(n1233) );
INV_X1 U976 ( .A(n1091), .ZN(n1236) );
NOR2_X1 U977 ( .A1(n1283), .A2(n1241), .ZN(n1091) );
XOR2_X1 U978 ( .A(n1232), .B(n1318), .Z(G15) );
NOR2_X1 U979 ( .A1(KEYINPUT61), .A2(n1319), .ZN(n1318) );
XNOR2_X1 U980 ( .A(KEYINPUT10), .B(n1320), .ZN(n1319) );
NOR3_X1 U981 ( .A1(n1199), .A2(n1294), .A3(n1316), .ZN(n1232) );
NAND2_X1 U982 ( .A1(n1124), .A2(n1245), .ZN(n1316) );
NOR2_X1 U983 ( .A1(n1123), .A2(n1108), .ZN(n1124) );
INV_X1 U984 ( .A(n1298), .ZN(n1108) );
INV_X1 U985 ( .A(n1114), .ZN(n1294) );
NAND2_X1 U986 ( .A1(n1321), .A2(n1322), .ZN(n1114) );
NAND3_X1 U987 ( .A1(n1151), .A2(n1323), .A3(n1315), .ZN(n1322) );
INV_X1 U988 ( .A(KEYINPUT26), .ZN(n1315) );
NAND2_X1 U989 ( .A1(KEYINPUT26), .A2(n1105), .ZN(n1321) );
NOR2_X1 U990 ( .A1(n1314), .A2(n1151), .ZN(n1105) );
INV_X1 U991 ( .A(n1129), .ZN(n1199) );
NOR2_X1 U992 ( .A1(n1284), .A2(n1242), .ZN(n1129) );
XNOR2_X1 U993 ( .A(n1231), .B(n1324), .ZN(G12) );
NOR2_X1 U994 ( .A1(G110), .A2(KEYINPUT9), .ZN(n1324) );
AND3_X1 U995 ( .A1(n1113), .A2(n1237), .A3(n1104), .ZN(n1231) );
NOR2_X1 U996 ( .A1(n1284), .A2(n1283), .ZN(n1104) );
INV_X1 U997 ( .A(n1242), .ZN(n1283) );
NOR2_X1 U998 ( .A1(n1325), .A2(n1143), .ZN(n1242) );
NOR3_X1 U999 ( .A1(G475), .A2(G902), .A3(n1147), .ZN(n1143) );
XNOR2_X1 U1000 ( .A(n1326), .B(KEYINPUT57), .ZN(n1325) );
NAND2_X1 U1001 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
OR2_X1 U1002 ( .A1(n1147), .A2(G902), .ZN(n1328) );
XNOR2_X1 U1003 ( .A(n1329), .B(n1330), .ZN(n1147) );
XOR2_X1 U1004 ( .A(n1331), .B(n1332), .Z(n1330) );
XNOR2_X1 U1005 ( .A(n1333), .B(n1334), .ZN(n1332) );
NOR2_X1 U1006 ( .A1(KEYINPUT27), .A2(n1320), .ZN(n1334) );
INV_X1 U1007 ( .A(G113), .ZN(n1320) );
NOR2_X1 U1008 ( .A1(KEYINPUT1), .A2(n1335), .ZN(n1333) );
XNOR2_X1 U1009 ( .A(G131), .B(KEYINPUT51), .ZN(n1335) );
XNOR2_X1 U1010 ( .A(G104), .B(G122), .ZN(n1331) );
XOR2_X1 U1011 ( .A(n1336), .B(n1337), .Z(n1329) );
XOR2_X1 U1012 ( .A(n1338), .B(n1339), .Z(n1336) );
AND2_X1 U1013 ( .A1(n1340), .A2(G214), .ZN(n1339) );
NAND3_X1 U1014 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1338) );
NAND2_X1 U1015 ( .A1(G125), .A2(n1288), .ZN(n1343) );
NAND2_X1 U1016 ( .A1(n1344), .A2(n1345), .ZN(n1342) );
INV_X1 U1017 ( .A(KEYINPUT37), .ZN(n1345) );
NAND2_X1 U1018 ( .A1(n1346), .A2(G140), .ZN(n1344) );
XNOR2_X1 U1019 ( .A(KEYINPUT8), .B(G125), .ZN(n1346) );
NAND2_X1 U1020 ( .A1(KEYINPUT37), .A2(n1347), .ZN(n1341) );
NAND2_X1 U1021 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
OR3_X1 U1022 ( .A1(n1288), .A2(G125), .A3(KEYINPUT8), .ZN(n1349) );
NAND2_X1 U1023 ( .A1(KEYINPUT8), .A2(G125), .ZN(n1348) );
XNOR2_X1 U1024 ( .A(G475), .B(KEYINPUT41), .ZN(n1327) );
INV_X1 U1025 ( .A(n1241), .ZN(n1284) );
NOR2_X1 U1026 ( .A1(n1350), .A2(n1142), .ZN(n1241) );
NOR3_X1 U1027 ( .A1(G478), .A2(G902), .A3(n1189), .ZN(n1142) );
INV_X1 U1028 ( .A(n1351), .ZN(n1189) );
XOR2_X1 U1029 ( .A(n1141), .B(KEYINPUT21), .Z(n1350) );
AND2_X1 U1030 ( .A1(G478), .A2(n1352), .ZN(n1141) );
NAND2_X1 U1031 ( .A1(n1353), .A2(n1351), .ZN(n1352) );
NAND2_X1 U1032 ( .A1(n1354), .A2(n1355), .ZN(n1351) );
NAND4_X1 U1033 ( .A1(G234), .A2(G217), .A3(n1356), .A4(n1116), .ZN(n1355) );
INV_X1 U1034 ( .A(n1357), .ZN(n1356) );
XOR2_X1 U1035 ( .A(n1358), .B(KEYINPUT36), .Z(n1354) );
NAND2_X1 U1036 ( .A1(n1357), .A2(n1359), .ZN(n1358) );
NAND3_X1 U1037 ( .A1(G217), .A2(n1116), .A3(G234), .ZN(n1359) );
XNOR2_X1 U1038 ( .A(n1360), .B(n1361), .ZN(n1357) );
NOR2_X1 U1039 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
AND2_X1 U1040 ( .A1(n1364), .A2(G107), .ZN(n1363) );
NOR2_X1 U1041 ( .A1(n1364), .A2(n1365), .ZN(n1362) );
XNOR2_X1 U1042 ( .A(G107), .B(KEYINPUT22), .ZN(n1365) );
XNOR2_X1 U1043 ( .A(n1366), .B(G122), .ZN(n1364) );
NAND2_X1 U1044 ( .A1(KEYINPUT35), .A2(n1317), .ZN(n1366) );
NAND3_X1 U1045 ( .A1(n1367), .A2(n1368), .A3(n1369), .ZN(n1360) );
OR2_X1 U1046 ( .A1(n1370), .A2(KEYINPUT54), .ZN(n1369) );
NAND3_X1 U1047 ( .A1(KEYINPUT54), .A2(n1371), .A3(n1293), .ZN(n1368) );
OR2_X1 U1048 ( .A1(n1293), .A2(n1371), .ZN(n1367) );
NOR2_X1 U1049 ( .A1(KEYINPUT62), .A2(n1372), .ZN(n1371) );
AND3_X1 U1050 ( .A1(n1123), .A2(n1298), .A3(n1245), .ZN(n1237) );
AND2_X1 U1051 ( .A1(n1287), .A2(n1373), .ZN(n1245) );
NAND2_X1 U1052 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
NAND3_X1 U1053 ( .A1(n1172), .A2(n1302), .A3(G902), .ZN(n1375) );
NOR2_X1 U1054 ( .A1(G898), .A2(n1116), .ZN(n1172) );
XNOR2_X1 U1055 ( .A(KEYINPUT20), .B(n1107), .ZN(n1374) );
NAND3_X1 U1056 ( .A1(n1302), .A2(n1116), .A3(G952), .ZN(n1107) );
NAND2_X1 U1057 ( .A1(G237), .A2(G234), .ZN(n1302) );
NOR2_X1 U1058 ( .A1(n1135), .A2(n1134), .ZN(n1287) );
INV_X1 U1059 ( .A(n1295), .ZN(n1134) );
NAND2_X1 U1060 ( .A1(G214), .A2(n1376), .ZN(n1295) );
XOR2_X1 U1061 ( .A(n1377), .B(n1225), .Z(n1135) );
AND2_X1 U1062 ( .A1(G210), .A2(n1376), .ZN(n1225) );
NAND2_X1 U1063 ( .A1(n1378), .A2(n1353), .ZN(n1376) );
INV_X1 U1064 ( .A(G237), .ZN(n1378) );
NAND2_X1 U1065 ( .A1(n1379), .A2(n1353), .ZN(n1377) );
XOR2_X1 U1066 ( .A(n1173), .B(n1380), .Z(n1379) );
XOR2_X1 U1067 ( .A(KEYINPUT49), .B(n1381), .Z(n1380) );
NOR2_X1 U1068 ( .A1(n1270), .A2(n1276), .ZN(n1381) );
NAND2_X1 U1069 ( .A1(n1382), .A2(n1383), .ZN(n1276) );
NAND2_X1 U1070 ( .A1(n1384), .A2(n1385), .ZN(n1383) );
XNOR2_X1 U1071 ( .A(n1273), .B(n1275), .ZN(n1384) );
NAND3_X1 U1072 ( .A1(n1273), .A2(n1386), .A3(G125), .ZN(n1382) );
NOR3_X1 U1073 ( .A1(n1386), .A2(n1273), .A3(n1385), .ZN(n1270) );
NOR2_X1 U1074 ( .A1(n1177), .A2(G953), .ZN(n1273) );
INV_X1 U1075 ( .A(G224), .ZN(n1177) );
INV_X1 U1076 ( .A(n1275), .ZN(n1386) );
XOR2_X1 U1077 ( .A(n1387), .B(n1388), .Z(n1173) );
XOR2_X1 U1078 ( .A(G122), .B(G110), .Z(n1388) );
XOR2_X1 U1079 ( .A(n1389), .B(n1390), .Z(n1387) );
NAND2_X1 U1080 ( .A1(n1391), .A2(n1392), .ZN(n1389) );
NAND2_X1 U1081 ( .A1(n1393), .A2(n1394), .ZN(n1392) );
XOR2_X1 U1082 ( .A(n1395), .B(KEYINPUT30), .Z(n1393) );
NAND2_X1 U1083 ( .A1(G101), .A2(n1396), .ZN(n1391) );
XOR2_X1 U1084 ( .A(n1395), .B(KEYINPUT16), .Z(n1396) );
XNOR2_X1 U1085 ( .A(n1397), .B(n1398), .ZN(n1395) );
INV_X1 U1086 ( .A(G104), .ZN(n1398) );
NAND2_X1 U1087 ( .A1(KEYINPUT28), .A2(n1399), .ZN(n1397) );
NAND2_X1 U1088 ( .A1(G221), .A2(n1400), .ZN(n1298) );
XOR2_X1 U1089 ( .A(n1401), .B(n1220), .Z(n1123) );
INV_X1 U1090 ( .A(G469), .ZN(n1220) );
NAND2_X1 U1091 ( .A1(n1402), .A2(n1353), .ZN(n1401) );
XOR2_X1 U1092 ( .A(n1164), .B(n1403), .Z(n1402) );
XNOR2_X1 U1093 ( .A(n1404), .B(n1219), .ZN(n1403) );
XNOR2_X1 U1094 ( .A(n1405), .B(n1406), .ZN(n1219) );
XNOR2_X1 U1095 ( .A(n1288), .B(G110), .ZN(n1406) );
INV_X1 U1096 ( .A(G140), .ZN(n1288) );
XNOR2_X1 U1097 ( .A(n1407), .B(n1408), .ZN(n1405) );
AND2_X1 U1098 ( .A1(n1116), .A2(G227), .ZN(n1408) );
NAND2_X1 U1099 ( .A1(KEYINPUT13), .A2(n1217), .ZN(n1404) );
XOR2_X1 U1100 ( .A(n1394), .B(n1409), .Z(n1217) );
XNOR2_X1 U1101 ( .A(n1399), .B(G104), .ZN(n1409) );
INV_X1 U1102 ( .A(G107), .ZN(n1399) );
XNOR2_X1 U1103 ( .A(n1410), .B(n1337), .ZN(n1164) );
XNOR2_X1 U1104 ( .A(n1278), .B(n1411), .ZN(n1337) );
NOR2_X1 U1105 ( .A1(n1151), .A2(n1323), .ZN(n1113) );
INV_X1 U1106 ( .A(n1314), .ZN(n1323) );
XOR2_X1 U1107 ( .A(n1150), .B(n1148), .Z(n1314) );
NAND2_X1 U1108 ( .A1(G217), .A2(n1400), .ZN(n1148) );
NAND2_X1 U1109 ( .A1(G234), .A2(n1353), .ZN(n1400) );
NAND2_X1 U1110 ( .A1(n1412), .A2(n1181), .ZN(n1150) );
XOR2_X1 U1111 ( .A(n1413), .B(n1414), .Z(n1181) );
XNOR2_X1 U1112 ( .A(n1415), .B(n1159), .ZN(n1414) );
XNOR2_X1 U1113 ( .A(G140), .B(n1385), .ZN(n1159) );
INV_X1 U1114 ( .A(G125), .ZN(n1385) );
NAND3_X1 U1115 ( .A1(n1416), .A2(n1417), .A3(n1418), .ZN(n1415) );
NAND2_X1 U1116 ( .A1(KEYINPUT46), .A2(n1419), .ZN(n1418) );
NAND3_X1 U1117 ( .A1(n1420), .A2(n1421), .A3(n1422), .ZN(n1417) );
INV_X1 U1118 ( .A(KEYINPUT46), .ZN(n1421) );
OR2_X1 U1119 ( .A1(n1422), .A2(n1420), .ZN(n1416) );
NOR2_X1 U1120 ( .A1(KEYINPUT50), .A2(n1419), .ZN(n1420) );
NAND3_X1 U1121 ( .A1(G234), .A2(n1116), .A3(G221), .ZN(n1422) );
INV_X1 U1122 ( .A(G953), .ZN(n1116) );
XNOR2_X1 U1123 ( .A(n1423), .B(n1278), .ZN(n1413) );
NAND2_X1 U1124 ( .A1(n1424), .A2(n1425), .ZN(n1423) );
OR2_X1 U1125 ( .A1(n1426), .A2(G110), .ZN(n1425) );
XOR2_X1 U1126 ( .A(n1427), .B(KEYINPUT19), .Z(n1424) );
NAND2_X1 U1127 ( .A1(G110), .A2(n1426), .ZN(n1427) );
XNOR2_X1 U1128 ( .A(G119), .B(n1410), .ZN(n1426) );
INV_X1 U1129 ( .A(G128), .ZN(n1410) );
XNOR2_X1 U1130 ( .A(G902), .B(KEYINPUT7), .ZN(n1412) );
XOR2_X1 U1131 ( .A(n1428), .B(n1213), .Z(n1151) );
INV_X1 U1132 ( .A(G472), .ZN(n1213) );
NAND2_X1 U1133 ( .A1(n1429), .A2(n1353), .ZN(n1428) );
INV_X1 U1134 ( .A(G902), .ZN(n1353) );
XNOR2_X1 U1135 ( .A(n1430), .B(n1208), .ZN(n1429) );
NAND2_X1 U1136 ( .A1(n1431), .A2(n1432), .ZN(n1208) );
OR2_X1 U1137 ( .A1(n1390), .A2(KEYINPUT43), .ZN(n1432) );
XNOR2_X1 U1138 ( .A(n1433), .B(n1434), .ZN(n1390) );
NAND3_X1 U1139 ( .A1(n1434), .A2(n1433), .A3(KEYINPUT43), .ZN(n1431) );
XNOR2_X1 U1140 ( .A(G113), .B(KEYINPUT39), .ZN(n1433) );
XNOR2_X1 U1141 ( .A(n1317), .B(G119), .ZN(n1434) );
INV_X1 U1142 ( .A(G116), .ZN(n1317) );
XNOR2_X1 U1143 ( .A(n1204), .B(n1212), .ZN(n1430) );
XNOR2_X1 U1144 ( .A(n1275), .B(n1407), .ZN(n1212) );
XNOR2_X1 U1145 ( .A(G131), .B(n1167), .ZN(n1407) );
XNOR2_X1 U1146 ( .A(n1293), .B(n1419), .ZN(n1167) );
INV_X1 U1147 ( .A(G137), .ZN(n1419) );
INV_X1 U1148 ( .A(G134), .ZN(n1293) );
NAND2_X1 U1149 ( .A1(n1435), .A2(n1436), .ZN(n1275) );
NAND2_X1 U1150 ( .A1(G146), .A2(n1370), .ZN(n1436) );
INV_X1 U1151 ( .A(n1372), .ZN(n1370) );
NAND2_X1 U1152 ( .A1(n1437), .A2(n1278), .ZN(n1435) );
INV_X1 U1153 ( .A(G146), .ZN(n1278) );
XNOR2_X1 U1154 ( .A(n1372), .B(KEYINPUT23), .ZN(n1437) );
XOR2_X1 U1155 ( .A(G128), .B(n1411), .Z(n1372) );
XOR2_X1 U1156 ( .A(G143), .B(KEYINPUT18), .Z(n1411) );
XOR2_X1 U1157 ( .A(n1438), .B(n1394), .Z(n1204) );
INV_X1 U1158 ( .A(G101), .ZN(n1394) );
NAND2_X1 U1159 ( .A1(G210), .A2(n1340), .ZN(n1438) );
NOR2_X1 U1160 ( .A1(G953), .A2(G237), .ZN(n1340) );
endmodule


