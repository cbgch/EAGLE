//Key = 1111101000100001111011000101101010011000000100101010111110110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409;

XNOR2_X1 U764 ( .A(G107), .B(n1054), .ZN(G9) );
NAND4_X1 U765 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NOR2_X1 U766 ( .A1(n1059), .A2(n1060), .ZN(G75) );
NOR3_X1 U767 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NAND3_X1 U768 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1061) );
NAND2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U770 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND3_X1 U771 ( .A1(n1056), .A2(n1071), .A3(n1072), .ZN(n1070) );
NAND3_X1 U772 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1071) );
NAND2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
OR2_X1 U775 ( .A1(n1080), .A2(KEYINPUT37), .ZN(n1079) );
NAND2_X1 U776 ( .A1(n1081), .A2(n1082), .ZN(n1078) );
NAND2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(n1074) );
NAND2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U779 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
INV_X1 U780 ( .A(KEYINPUT45), .ZN(n1088) );
NAND3_X1 U781 ( .A1(KEYINPUT45), .A2(n1087), .A3(n1089), .ZN(n1073) );
INV_X1 U782 ( .A(n1083), .ZN(n1089) );
NAND2_X1 U783 ( .A1(n1076), .A2(n1090), .ZN(n1069) );
NAND2_X1 U784 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND3_X1 U785 ( .A1(n1056), .A2(n1093), .A3(n1083), .ZN(n1092) );
NAND2_X1 U786 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U787 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U788 ( .A1(n1072), .A2(n1098), .ZN(n1091) );
NAND2_X1 U789 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND3_X1 U790 ( .A1(n1101), .A2(n1102), .A3(KEYINPUT37), .ZN(n1100) );
NAND2_X1 U791 ( .A1(n1083), .A2(n1103), .ZN(n1099) );
OR2_X1 U792 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
INV_X1 U793 ( .A(n1106), .ZN(n1067) );
NOR3_X1 U794 ( .A1(n1107), .A2(G953), .A3(G952), .ZN(n1059) );
INV_X1 U795 ( .A(n1064), .ZN(n1107) );
NAND4_X1 U796 ( .A1(n1108), .A2(n1109), .A3(n1110), .A4(n1111), .ZN(n1064) );
NOR4_X1 U797 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1111) );
XOR2_X1 U798 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U799 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XNOR2_X1 U800 ( .A(n1120), .B(n1121), .ZN(n1113) );
NAND2_X1 U801 ( .A1(KEYINPUT1), .A2(n1122), .ZN(n1121) );
NAND3_X1 U802 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1112) );
XOR2_X1 U803 ( .A(n1126), .B(n1127), .Z(n1125) );
OR3_X1 U804 ( .A1(n1128), .A2(n1129), .A3(KEYINPUT31), .ZN(n1124) );
NAND2_X1 U805 ( .A1(KEYINPUT31), .A2(n1128), .ZN(n1123) );
NOR3_X1 U806 ( .A1(n1096), .A2(n1130), .A3(n1081), .ZN(n1110) );
OR2_X1 U807 ( .A1(n1119), .A2(n1118), .ZN(n1109) );
XOR2_X1 U808 ( .A(G475), .B(KEYINPUT41), .Z(n1118) );
INV_X1 U809 ( .A(KEYINPUT38), .ZN(n1119) );
XOR2_X1 U810 ( .A(KEYINPUT36), .B(n1131), .Z(n1108) );
XOR2_X1 U811 ( .A(n1132), .B(n1133), .Z(G72) );
NOR2_X1 U812 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U813 ( .A(n1065), .B(KEYINPUT11), .Z(n1135) );
AND2_X1 U814 ( .A1(G227), .A2(G900), .ZN(n1134) );
NAND2_X1 U815 ( .A1(n1136), .A2(n1137), .ZN(n1132) );
NAND2_X1 U816 ( .A1(n1138), .A2(n1065), .ZN(n1137) );
XOR2_X1 U817 ( .A(n1062), .B(n1139), .Z(n1138) );
NAND3_X1 U818 ( .A1(n1139), .A2(G900), .A3(G953), .ZN(n1136) );
AND2_X1 U819 ( .A1(n1140), .A2(KEYINPUT17), .ZN(n1139) );
XOR2_X1 U820 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U821 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U822 ( .A1(KEYINPUT24), .A2(n1145), .ZN(n1143) );
XOR2_X1 U823 ( .A(n1146), .B(n1147), .Z(n1141) );
NOR2_X1 U824 ( .A1(KEYINPUT33), .A2(n1148), .ZN(n1147) );
NOR2_X1 U825 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
XOR2_X1 U826 ( .A(n1151), .B(KEYINPUT25), .Z(n1150) );
NAND2_X1 U827 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NOR2_X1 U828 ( .A1(n1153), .A2(n1152), .ZN(n1149) );
XNOR2_X1 U829 ( .A(n1154), .B(G137), .ZN(n1152) );
NAND2_X1 U830 ( .A1(KEYINPUT6), .A2(n1155), .ZN(n1154) );
XOR2_X1 U831 ( .A(n1156), .B(n1157), .Z(G69) );
XOR2_X1 U832 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND2_X1 U833 ( .A1(G953), .A2(n1160), .ZN(n1159) );
NAND2_X1 U834 ( .A1(G898), .A2(G224), .ZN(n1160) );
NAND3_X1 U835 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1158) );
XOR2_X1 U836 ( .A(n1164), .B(KEYINPUT47), .Z(n1163) );
NAND2_X1 U837 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
OR2_X1 U838 ( .A1(n1166), .A2(n1165), .ZN(n1162) );
NAND2_X1 U839 ( .A1(G953), .A2(n1167), .ZN(n1161) );
AND2_X1 U840 ( .A1(n1063), .A2(n1065), .ZN(n1156) );
NOR2_X1 U841 ( .A1(n1168), .A2(n1169), .ZN(G66) );
XNOR2_X1 U842 ( .A(n1170), .B(n1171), .ZN(n1169) );
NOR2_X1 U843 ( .A1(n1128), .A2(n1172), .ZN(n1171) );
NOR2_X1 U844 ( .A1(n1168), .A2(n1173), .ZN(G63) );
NOR3_X1 U845 ( .A1(n1127), .A2(n1174), .A3(n1175), .ZN(n1173) );
AND3_X1 U846 ( .A1(n1176), .A2(G478), .A3(n1177), .ZN(n1175) );
NOR2_X1 U847 ( .A1(n1178), .A2(n1176), .ZN(n1174) );
NOR2_X1 U848 ( .A1(n1179), .A2(n1126), .ZN(n1178) );
NOR2_X1 U849 ( .A1(n1062), .A2(n1063), .ZN(n1179) );
NOR3_X1 U850 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(G60) );
AND2_X1 U851 ( .A1(KEYINPUT30), .A2(n1168), .ZN(n1182) );
NOR3_X1 U852 ( .A1(KEYINPUT30), .A2(G953), .A3(G952), .ZN(n1181) );
XOR2_X1 U853 ( .A(n1183), .B(n1184), .Z(n1180) );
NAND2_X1 U854 ( .A1(KEYINPUT50), .A2(n1185), .ZN(n1183) );
NAND2_X1 U855 ( .A1(n1177), .A2(G475), .ZN(n1185) );
NAND3_X1 U856 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(G6) );
NAND2_X1 U857 ( .A1(G104), .A2(n1189), .ZN(n1188) );
NAND2_X1 U858 ( .A1(KEYINPUT12), .A2(n1190), .ZN(n1187) );
NAND2_X1 U859 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
INV_X1 U860 ( .A(n1189), .ZN(n1192) );
XNOR2_X1 U861 ( .A(KEYINPUT34), .B(G104), .ZN(n1191) );
NAND2_X1 U862 ( .A1(n1193), .A2(n1194), .ZN(n1186) );
INV_X1 U863 ( .A(KEYINPUT12), .ZN(n1194) );
NAND2_X1 U864 ( .A1(n1195), .A2(n1196), .ZN(n1193) );
OR3_X1 U865 ( .A1(n1189), .A2(G104), .A3(KEYINPUT34), .ZN(n1196) );
NAND2_X1 U866 ( .A1(KEYINPUT34), .A2(G104), .ZN(n1195) );
NOR3_X1 U867 ( .A1(n1168), .A2(n1197), .A3(n1198), .ZN(G57) );
NOR2_X1 U868 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U869 ( .A(n1201), .B(KEYINPUT58), .Z(n1200) );
NOR2_X1 U870 ( .A1(n1202), .A2(n1203), .ZN(n1197) );
XOR2_X1 U871 ( .A(n1201), .B(KEYINPUT23), .Z(n1203) );
XOR2_X1 U872 ( .A(n1204), .B(n1205), .Z(n1201) );
AND2_X1 U873 ( .A1(G472), .A2(n1177), .ZN(n1205) );
XOR2_X1 U874 ( .A(n1206), .B(G101), .Z(n1204) );
NOR2_X1 U875 ( .A1(n1168), .A2(n1207), .ZN(G54) );
XOR2_X1 U876 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U877 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U878 ( .A(n1212), .B(n1213), .Z(n1211) );
XOR2_X1 U879 ( .A(n1214), .B(n1215), .Z(n1208) );
XNOR2_X1 U880 ( .A(KEYINPUT55), .B(n1216), .ZN(n1215) );
NOR2_X1 U881 ( .A1(n1217), .A2(KEYINPUT57), .ZN(n1216) );
AND2_X1 U882 ( .A1(G469), .A2(n1177), .ZN(n1217) );
INV_X1 U883 ( .A(n1172), .ZN(n1177) );
NOR2_X1 U884 ( .A1(n1168), .A2(n1218), .ZN(G51) );
XOR2_X1 U885 ( .A(n1219), .B(n1220), .Z(n1218) );
XOR2_X1 U886 ( .A(n1221), .B(n1222), .Z(n1220) );
NOR2_X1 U887 ( .A1(n1223), .A2(n1172), .ZN(n1222) );
NAND2_X1 U888 ( .A1(G902), .A2(n1224), .ZN(n1172) );
OR2_X1 U889 ( .A1(n1063), .A2(n1062), .ZN(n1224) );
NAND4_X1 U890 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1062) );
AND4_X1 U891 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1228) );
NAND2_X1 U892 ( .A1(n1233), .A2(n1234), .ZN(n1227) );
NAND2_X1 U893 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NAND3_X1 U894 ( .A1(n1237), .A2(n1238), .A3(n1105), .ZN(n1236) );
NAND2_X1 U895 ( .A1(n1055), .A2(n1239), .ZN(n1235) );
XOR2_X1 U896 ( .A(n1240), .B(KEYINPUT22), .Z(n1239) );
NAND4_X1 U897 ( .A1(n1241), .A2(n1189), .A3(n1242), .A4(n1243), .ZN(n1063) );
NOR4_X1 U898 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1247), .ZN(n1243) );
NOR3_X1 U899 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1247) );
XOR2_X1 U900 ( .A(n1058), .B(KEYINPUT59), .Z(n1249) );
NOR4_X1 U901 ( .A1(n1251), .A2(n1085), .A3(n1252), .A4(n1253), .ZN(n1246) );
NOR2_X1 U902 ( .A1(KEYINPUT48), .A2(n1254), .ZN(n1253) );
NOR2_X1 U903 ( .A1(n1255), .A2(n1080), .ZN(n1254) );
AND2_X1 U904 ( .A1(n1250), .A2(KEYINPUT48), .ZN(n1252) );
NAND2_X1 U905 ( .A1(n1056), .A2(n1058), .ZN(n1251) );
INV_X1 U906 ( .A(n1256), .ZN(n1245) );
NOR2_X1 U907 ( .A1(n1257), .A2(n1258), .ZN(n1242) );
INV_X1 U908 ( .A(n1259), .ZN(n1258) );
NAND4_X1 U909 ( .A1(n1087), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1189) );
NOR2_X1 U910 ( .A1(n1260), .A2(n1261), .ZN(n1221) );
XOR2_X1 U911 ( .A(n1262), .B(KEYINPUT28), .Z(n1261) );
NAND3_X1 U912 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1262) );
NOR2_X1 U913 ( .A1(n1266), .A2(n1264), .ZN(n1260) );
AND2_X1 U914 ( .A1(n1263), .A2(n1265), .ZN(n1266) );
NAND2_X1 U915 ( .A1(n1267), .A2(n1268), .ZN(n1265) );
INV_X1 U916 ( .A(KEYINPUT13), .ZN(n1268) );
NAND3_X1 U917 ( .A1(n1269), .A2(G125), .A3(KEYINPUT13), .ZN(n1263) );
NOR2_X1 U918 ( .A1(n1065), .A2(G952), .ZN(n1168) );
XOR2_X1 U919 ( .A(n1270), .B(n1225), .Z(G48) );
NAND3_X1 U920 ( .A1(n1087), .A2(n1240), .A3(n1233), .ZN(n1225) );
XOR2_X1 U921 ( .A(n1271), .B(n1272), .Z(G45) );
NAND4_X1 U922 ( .A1(n1237), .A2(n1233), .A3(n1273), .A4(n1238), .ZN(n1272) );
XOR2_X1 U923 ( .A(KEYINPUT39), .B(n1105), .Z(n1273) );
XOR2_X1 U924 ( .A(n1146), .B(n1226), .Z(G42) );
NAND3_X1 U925 ( .A1(n1104), .A2(n1087), .A3(n1274), .ZN(n1226) );
XNOR2_X1 U926 ( .A(G137), .B(n1232), .ZN(G39) );
NAND3_X1 U927 ( .A1(n1076), .A2(n1240), .A3(n1274), .ZN(n1232) );
XOR2_X1 U928 ( .A(n1231), .B(n1275), .Z(G36) );
NOR2_X1 U929 ( .A1(G134), .A2(KEYINPUT8), .ZN(n1275) );
NAND3_X1 U930 ( .A1(n1105), .A2(n1055), .A3(n1274), .ZN(n1231) );
XNOR2_X1 U931 ( .A(G131), .B(n1230), .ZN(G33) );
NAND3_X1 U932 ( .A1(n1105), .A2(n1087), .A3(n1274), .ZN(n1230) );
AND3_X1 U933 ( .A1(n1101), .A2(n1276), .A3(n1072), .ZN(n1274) );
NOR2_X1 U934 ( .A1(n1277), .A2(n1096), .ZN(n1072) );
INV_X1 U935 ( .A(n1097), .ZN(n1277) );
XOR2_X1 U936 ( .A(G128), .B(n1278), .Z(G30) );
NOR2_X1 U937 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NOR2_X1 U938 ( .A1(KEYINPUT19), .A2(n1281), .ZN(n1280) );
INV_X1 U939 ( .A(n1282), .ZN(n1281) );
NOR2_X1 U940 ( .A1(KEYINPUT52), .A2(n1282), .ZN(n1279) );
NAND3_X1 U941 ( .A1(n1055), .A2(n1240), .A3(n1233), .ZN(n1282) );
NOR2_X1 U942 ( .A1(n1250), .A2(n1283), .ZN(n1233) );
XOR2_X1 U943 ( .A(n1284), .B(n1256), .Z(G3) );
NAND4_X1 U944 ( .A1(n1076), .A2(n1105), .A3(n1057), .A4(n1058), .ZN(n1256) );
XOR2_X1 U945 ( .A(n1145), .B(n1229), .Z(G27) );
NAND4_X1 U946 ( .A1(n1104), .A2(n1083), .A3(n1285), .A4(n1087), .ZN(n1229) );
NOR2_X1 U947 ( .A1(n1283), .A2(n1094), .ZN(n1285) );
INV_X1 U948 ( .A(n1255), .ZN(n1094) );
INV_X1 U949 ( .A(n1276), .ZN(n1283) );
NAND2_X1 U950 ( .A1(n1106), .A2(n1286), .ZN(n1276) );
NAND4_X1 U951 ( .A1(G953), .A2(G902), .A3(n1287), .A4(n1288), .ZN(n1286) );
INV_X1 U952 ( .A(G900), .ZN(n1288) );
XOR2_X1 U953 ( .A(G122), .B(n1244), .Z(G24) );
AND4_X1 U954 ( .A1(n1237), .A2(n1289), .A3(n1056), .A4(n1238), .ZN(n1244) );
INV_X1 U955 ( .A(n1102), .ZN(n1056) );
NAND2_X1 U956 ( .A1(n1290), .A2(n1291), .ZN(n1102) );
XNOR2_X1 U957 ( .A(n1292), .B(KEYINPUT5), .ZN(n1290) );
NAND2_X1 U958 ( .A1(n1293), .A2(n1294), .ZN(G21) );
OR2_X1 U959 ( .A1(n1259), .A2(G119), .ZN(n1294) );
XOR2_X1 U960 ( .A(n1295), .B(KEYINPUT14), .Z(n1293) );
NAND2_X1 U961 ( .A1(G119), .A2(n1259), .ZN(n1295) );
NAND3_X1 U962 ( .A1(n1289), .A2(n1240), .A3(n1076), .ZN(n1259) );
NAND2_X1 U963 ( .A1(n1296), .A2(n1297), .ZN(n1240) );
OR3_X1 U964 ( .A1(n1298), .A2(n1291), .A3(KEYINPUT29), .ZN(n1297) );
INV_X1 U965 ( .A(n1292), .ZN(n1298) );
NAND2_X1 U966 ( .A1(KEYINPUT29), .A2(n1104), .ZN(n1296) );
XOR2_X1 U967 ( .A(G116), .B(n1257), .Z(G18) );
AND3_X1 U968 ( .A1(n1105), .A2(n1055), .A3(n1289), .ZN(n1257) );
INV_X1 U969 ( .A(n1085), .ZN(n1055) );
NAND2_X1 U970 ( .A1(n1299), .A2(n1238), .ZN(n1085) );
XNOR2_X1 U971 ( .A(G113), .B(n1241), .ZN(G15) );
NAND3_X1 U972 ( .A1(n1105), .A2(n1087), .A3(n1289), .ZN(n1241) );
AND3_X1 U973 ( .A1(n1255), .A2(n1058), .A3(n1083), .ZN(n1289) );
NOR2_X1 U974 ( .A1(n1131), .A2(n1081), .ZN(n1083) );
INV_X1 U975 ( .A(n1082), .ZN(n1131) );
NOR2_X1 U976 ( .A1(n1238), .A2(n1299), .ZN(n1087) );
INV_X1 U977 ( .A(n1237), .ZN(n1299) );
AND2_X1 U978 ( .A1(n1291), .A2(n1300), .ZN(n1105) );
XOR2_X1 U979 ( .A(KEYINPUT29), .B(n1292), .Z(n1300) );
NAND2_X1 U980 ( .A1(n1301), .A2(n1302), .ZN(G12) );
NAND4_X1 U981 ( .A1(n1303), .A2(n1304), .A3(n1058), .A4(n1305), .ZN(n1302) );
INV_X1 U982 ( .A(G110), .ZN(n1305) );
XOR2_X1 U983 ( .A(n1306), .B(KEYINPUT60), .Z(n1301) );
NAND2_X1 U984 ( .A1(G110), .A2(n1307), .ZN(n1306) );
NAND3_X1 U985 ( .A1(n1304), .A2(n1058), .A3(n1303), .ZN(n1307) );
INV_X1 U986 ( .A(n1248), .ZN(n1303) );
NAND2_X1 U987 ( .A1(n1076), .A2(n1104), .ZN(n1248) );
NOR2_X1 U988 ( .A1(n1292), .A2(n1291), .ZN(n1104) );
NOR2_X1 U989 ( .A1(n1130), .A2(n1308), .ZN(n1291) );
NOR2_X1 U990 ( .A1(n1128), .A2(n1129), .ZN(n1308) );
AND2_X1 U991 ( .A1(n1129), .A2(n1128), .ZN(n1130) );
NAND2_X1 U992 ( .A1(G217), .A2(n1309), .ZN(n1128) );
AND2_X1 U993 ( .A1(n1310), .A2(n1170), .ZN(n1129) );
NAND2_X1 U994 ( .A1(n1311), .A2(n1312), .ZN(n1170) );
NAND2_X1 U995 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U996 ( .A(n1315), .B(KEYINPUT9), .Z(n1311) );
OR2_X1 U997 ( .A1(n1314), .A2(n1313), .ZN(n1315) );
XOR2_X1 U998 ( .A(n1316), .B(n1317), .Z(n1313) );
XOR2_X1 U999 ( .A(G119), .B(G110), .Z(n1317) );
XOR2_X1 U1000 ( .A(n1318), .B(n1319), .Z(n1316) );
NAND2_X1 U1001 ( .A1(KEYINPUT3), .A2(n1320), .ZN(n1318) );
XOR2_X1 U1002 ( .A(n1270), .B(n1321), .Z(n1320) );
NAND2_X1 U1003 ( .A1(KEYINPUT46), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1004 ( .A(G140), .B(G125), .Z(n1322) );
XNOR2_X1 U1005 ( .A(n1323), .B(n1324), .ZN(n1314) );
XOR2_X1 U1006 ( .A(KEYINPUT2), .B(G137), .Z(n1324) );
NAND2_X1 U1007 ( .A1(G221), .A2(n1325), .ZN(n1323) );
XOR2_X1 U1008 ( .A(n1114), .B(KEYINPUT42), .Z(n1292) );
XNOR2_X1 U1009 ( .A(n1326), .B(G472), .ZN(n1114) );
NAND2_X1 U1010 ( .A1(n1327), .A2(n1310), .ZN(n1326) );
XOR2_X1 U1011 ( .A(n1328), .B(n1329), .Z(n1327) );
XOR2_X1 U1012 ( .A(n1206), .B(n1330), .Z(n1329) );
NOR2_X1 U1013 ( .A1(G101), .A2(KEYINPUT40), .ZN(n1330) );
NAND3_X1 U1014 ( .A1(n1331), .A2(n1065), .A3(G210), .ZN(n1206) );
NAND2_X1 U1015 ( .A1(KEYINPUT16), .A2(n1202), .ZN(n1328) );
INV_X1 U1016 ( .A(n1199), .ZN(n1202) );
XOR2_X1 U1017 ( .A(n1210), .B(n1332), .Z(n1199) );
XOR2_X1 U1018 ( .A(n1333), .B(n1334), .Z(n1332) );
NOR2_X1 U1019 ( .A1(n1238), .A2(n1237), .ZN(n1076) );
XOR2_X1 U1020 ( .A(n1116), .B(n1335), .Z(n1237) );
XOR2_X1 U1021 ( .A(KEYINPUT15), .B(G475), .Z(n1335) );
OR2_X1 U1022 ( .A1(n1184), .A2(G902), .ZN(n1116) );
XNOR2_X1 U1023 ( .A(n1336), .B(n1337), .ZN(n1184) );
XOR2_X1 U1024 ( .A(G113), .B(n1338), .Z(n1337) );
XOR2_X1 U1025 ( .A(KEYINPUT27), .B(G122), .Z(n1338) );
XOR2_X1 U1026 ( .A(n1339), .B(G104), .Z(n1336) );
NAND2_X1 U1027 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
NAND2_X1 U1028 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
XOR2_X1 U1029 ( .A(n1344), .B(KEYINPUT62), .Z(n1340) );
OR2_X1 U1030 ( .A1(n1343), .A2(n1342), .ZN(n1344) );
XNOR2_X1 U1031 ( .A(n1345), .B(n1270), .ZN(n1342) );
NAND2_X1 U1032 ( .A1(n1346), .A2(KEYINPUT53), .ZN(n1345) );
XOR2_X1 U1033 ( .A(n1146), .B(G125), .Z(n1346) );
INV_X1 U1034 ( .A(G140), .ZN(n1146) );
XNOR2_X1 U1035 ( .A(n1347), .B(n1348), .ZN(n1343) );
XOR2_X1 U1036 ( .A(G143), .B(G131), .Z(n1348) );
NAND3_X1 U1037 ( .A1(n1331), .A2(n1065), .A3(G214), .ZN(n1347) );
NAND3_X1 U1038 ( .A1(n1349), .A2(n1350), .A3(n1351), .ZN(n1238) );
NAND2_X1 U1039 ( .A1(n1352), .A2(n1126), .ZN(n1351) );
INV_X1 U1040 ( .A(G478), .ZN(n1126) );
NAND2_X1 U1041 ( .A1(n1353), .A2(n1354), .ZN(n1350) );
INV_X1 U1042 ( .A(KEYINPUT35), .ZN(n1354) );
NAND2_X1 U1043 ( .A1(G478), .A2(n1355), .ZN(n1353) );
XOR2_X1 U1044 ( .A(KEYINPUT43), .B(n1352), .Z(n1355) );
INV_X1 U1045 ( .A(n1356), .ZN(n1352) );
NAND2_X1 U1046 ( .A1(KEYINPUT35), .A2(n1357), .ZN(n1349) );
NAND2_X1 U1047 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
NAND3_X1 U1048 ( .A1(KEYINPUT43), .A2(G478), .A3(n1356), .ZN(n1359) );
OR2_X1 U1049 ( .A1(n1356), .A2(KEYINPUT43), .ZN(n1358) );
XNOR2_X1 U1050 ( .A(n1127), .B(KEYINPUT44), .ZN(n1356) );
NOR2_X1 U1051 ( .A1(n1176), .A2(G902), .ZN(n1127) );
XNOR2_X1 U1052 ( .A(n1360), .B(n1361), .ZN(n1176) );
AND2_X1 U1053 ( .A1(n1325), .A2(G217), .ZN(n1361) );
AND2_X1 U1054 ( .A1(G234), .A2(n1065), .ZN(n1325) );
NAND3_X1 U1055 ( .A1(n1362), .A2(n1363), .A3(n1364), .ZN(n1360) );
OR2_X1 U1056 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
NAND2_X1 U1057 ( .A1(n1367), .A2(n1368), .ZN(n1363) );
INV_X1 U1058 ( .A(KEYINPUT21), .ZN(n1368) );
NAND2_X1 U1059 ( .A1(n1369), .A2(n1365), .ZN(n1367) );
XNOR2_X1 U1060 ( .A(KEYINPUT18), .B(n1366), .ZN(n1369) );
NAND2_X1 U1061 ( .A1(KEYINPUT21), .A2(n1370), .ZN(n1362) );
NAND2_X1 U1062 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
NAND3_X1 U1063 ( .A1(KEYINPUT18), .A2(n1365), .A3(n1366), .ZN(n1372) );
XNOR2_X1 U1064 ( .A(n1155), .B(n1373), .ZN(n1365) );
NOR2_X1 U1065 ( .A1(KEYINPUT26), .A2(n1374), .ZN(n1373) );
OR2_X1 U1066 ( .A1(n1366), .A2(KEYINPUT18), .ZN(n1371) );
XNOR2_X1 U1067 ( .A(G107), .B(n1375), .ZN(n1366) );
XOR2_X1 U1068 ( .A(G122), .B(G116), .Z(n1375) );
NAND2_X1 U1069 ( .A1(n1106), .A2(n1376), .ZN(n1058) );
NAND4_X1 U1070 ( .A1(G953), .A2(G902), .A3(n1287), .A4(n1167), .ZN(n1376) );
INV_X1 U1071 ( .A(G898), .ZN(n1167) );
NAND3_X1 U1072 ( .A1(n1287), .A2(n1065), .A3(G952), .ZN(n1106) );
NAND2_X1 U1073 ( .A1(G237), .A2(G234), .ZN(n1287) );
NAND2_X1 U1074 ( .A1(n1377), .A2(n1378), .ZN(n1304) );
OR3_X1 U1075 ( .A1(n1080), .A2(n1255), .A3(KEYINPUT61), .ZN(n1378) );
INV_X1 U1076 ( .A(n1101), .ZN(n1080) );
NAND2_X1 U1077 ( .A1(KEYINPUT61), .A2(n1057), .ZN(n1377) );
INV_X1 U1078 ( .A(n1250), .ZN(n1057) );
NAND2_X1 U1079 ( .A1(n1101), .A2(n1255), .ZN(n1250) );
NOR2_X1 U1080 ( .A1(n1097), .A2(n1096), .ZN(n1255) );
AND2_X1 U1081 ( .A1(G214), .A2(n1379), .ZN(n1096) );
XOR2_X1 U1082 ( .A(n1380), .B(n1122), .Z(n1097) );
INV_X1 U1083 ( .A(n1223), .ZN(n1122) );
NAND2_X1 U1084 ( .A1(G210), .A2(n1379), .ZN(n1223) );
NAND2_X1 U1085 ( .A1(n1331), .A2(n1310), .ZN(n1379) );
INV_X1 U1086 ( .A(G237), .ZN(n1331) );
NAND2_X1 U1087 ( .A1(KEYINPUT10), .A2(n1120), .ZN(n1380) );
AND2_X1 U1088 ( .A1(n1381), .A2(n1310), .ZN(n1120) );
XOR2_X1 U1089 ( .A(n1267), .B(n1382), .Z(n1381) );
XOR2_X1 U1090 ( .A(n1219), .B(n1264), .Z(n1382) );
NAND2_X1 U1091 ( .A1(G224), .A2(n1065), .ZN(n1264) );
XNOR2_X1 U1092 ( .A(n1166), .B(n1165), .ZN(n1219) );
XNOR2_X1 U1093 ( .A(G110), .B(G122), .ZN(n1165) );
XNOR2_X1 U1094 ( .A(n1214), .B(n1333), .ZN(n1166) );
XOR2_X1 U1095 ( .A(G113), .B(n1383), .Z(n1333) );
XOR2_X1 U1096 ( .A(G119), .B(G116), .Z(n1383) );
XOR2_X1 U1097 ( .A(n1145), .B(n1334), .Z(n1267) );
INV_X1 U1098 ( .A(n1269), .ZN(n1334) );
XOR2_X1 U1099 ( .A(n1384), .B(n1319), .Z(n1269) );
NAND2_X1 U1100 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
NAND2_X1 U1101 ( .A1(n1387), .A2(n1271), .ZN(n1386) );
NAND2_X1 U1102 ( .A1(n1270), .A2(n1388), .ZN(n1387) );
NAND2_X1 U1103 ( .A1(KEYINPUT51), .A2(KEYINPUT4), .ZN(n1388) );
NAND3_X1 U1104 ( .A1(n1389), .A2(n1390), .A3(n1391), .ZN(n1385) );
INV_X1 U1105 ( .A(KEYINPUT51), .ZN(n1391) );
OR2_X1 U1106 ( .A1(G146), .A2(KEYINPUT4), .ZN(n1390) );
NAND2_X1 U1107 ( .A1(KEYINPUT4), .A2(n1392), .ZN(n1389) );
NAND2_X1 U1108 ( .A1(G143), .A2(n1270), .ZN(n1392) );
INV_X1 U1109 ( .A(G146), .ZN(n1270) );
INV_X1 U1110 ( .A(G125), .ZN(n1145) );
NOR2_X1 U1111 ( .A1(n1082), .A2(n1081), .ZN(n1101) );
AND2_X1 U1112 ( .A1(G221), .A2(n1309), .ZN(n1081) );
NAND2_X1 U1113 ( .A1(G234), .A2(n1310), .ZN(n1309) );
XOR2_X1 U1114 ( .A(n1393), .B(G469), .Z(n1082) );
NAND3_X1 U1115 ( .A1(n1394), .A2(n1310), .A3(n1395), .ZN(n1393) );
NAND2_X1 U1116 ( .A1(n1396), .A2(n1397), .ZN(n1395) );
XOR2_X1 U1117 ( .A(n1398), .B(n1399), .Z(n1397) );
INV_X1 U1118 ( .A(n1214), .ZN(n1398) );
XOR2_X1 U1119 ( .A(n1400), .B(n1401), .Z(n1396) );
XOR2_X1 U1120 ( .A(KEYINPUT63), .B(KEYINPUT49), .Z(n1401) );
INV_X1 U1121 ( .A(G902), .ZN(n1310) );
NAND2_X1 U1122 ( .A1(n1402), .A2(n1403), .ZN(n1394) );
XOR2_X1 U1123 ( .A(KEYINPUT0), .B(n1213), .Z(n1403) );
INV_X1 U1124 ( .A(n1400), .ZN(n1213) );
XOR2_X1 U1125 ( .A(n1404), .B(n1405), .Z(n1400) );
XOR2_X1 U1126 ( .A(G140), .B(G110), .Z(n1405) );
NAND2_X1 U1127 ( .A1(G227), .A2(n1065), .ZN(n1404) );
INV_X1 U1128 ( .A(G953), .ZN(n1065) );
XOR2_X1 U1129 ( .A(n1214), .B(n1399), .Z(n1402) );
XNOR2_X1 U1130 ( .A(n1406), .B(n1407), .ZN(n1399) );
NOR2_X1 U1131 ( .A1(KEYINPUT7), .A2(n1212), .ZN(n1407) );
XNOR2_X1 U1132 ( .A(n1144), .B(KEYINPUT54), .ZN(n1212) );
XOR2_X1 U1133 ( .A(n1374), .B(G146), .Z(n1144) );
XNOR2_X1 U1134 ( .A(n1271), .B(n1319), .ZN(n1374) );
XOR2_X1 U1135 ( .A(G128), .B(KEYINPUT32), .Z(n1319) );
INV_X1 U1136 ( .A(G143), .ZN(n1271) );
NAND2_X1 U1137 ( .A1(KEYINPUT56), .A2(n1210), .ZN(n1406) );
XOR2_X1 U1138 ( .A(n1408), .B(n1153), .Z(n1210) );
XOR2_X1 U1139 ( .A(G131), .B(KEYINPUT20), .Z(n1153) );
XOR2_X1 U1140 ( .A(n1155), .B(G137), .Z(n1408) );
INV_X1 U1141 ( .A(G134), .ZN(n1155) );
XOR2_X1 U1142 ( .A(n1284), .B(n1409), .Z(n1214) );
XOR2_X1 U1143 ( .A(G107), .B(G104), .Z(n1409) );
INV_X1 U1144 ( .A(G101), .ZN(n1284) );
endmodule


