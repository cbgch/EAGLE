//Key = 1001111101110011000000000101101001000101000010010001101101010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404;

XNOR2_X1 U763 ( .A(G107), .B(n1064), .ZN(G9) );
NOR2_X1 U764 ( .A1(n1065), .A2(n1066), .ZN(G75) );
NOR4_X1 U765 ( .A1(G953), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1066) );
NOR2_X1 U766 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR2_X1 U768 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U769 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U771 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR2_X1 U772 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NOR2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR2_X1 U775 ( .A1(n1088), .A2(n1089), .ZN(n1080) );
NOR2_X1 U776 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR3_X1 U777 ( .A1(n1089), .A2(n1092), .A3(n1083), .ZN(n1076) );
NOR2_X1 U778 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U779 ( .A(n1095), .B(KEYINPUT24), .Z(n1094) );
NOR2_X1 U780 ( .A1(n1096), .A2(n1097), .ZN(n1093) );
NOR4_X1 U781 ( .A1(n1098), .A2(n1083), .A3(n1089), .A4(n1079), .ZN(n1072) );
NOR2_X1 U782 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NOR3_X1 U783 ( .A1(n1067), .A2(G953), .A3(G952), .ZN(n1065) );
AND4_X1 U784 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1067) );
NOR4_X1 U785 ( .A1(n1105), .A2(n1106), .A3(n1089), .A4(n1107), .ZN(n1104) );
INV_X1 U786 ( .A(n1108), .ZN(n1089) );
XOR2_X1 U787 ( .A(n1109), .B(n1110), .Z(n1106) );
NOR2_X1 U788 ( .A1(G469), .A2(KEYINPUT20), .ZN(n1110) );
XOR2_X1 U789 ( .A(n1111), .B(n1112), .Z(n1105) );
NOR3_X1 U790 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1103) );
NOR2_X1 U791 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U792 ( .A(n1118), .B(KEYINPUT32), .Z(n1117) );
XOR2_X1 U793 ( .A(n1119), .B(n1120), .Z(G72) );
NOR2_X1 U794 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
AND2_X1 U795 ( .A1(G227), .A2(G900), .ZN(n1121) );
NAND3_X1 U796 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1119) );
NAND2_X1 U797 ( .A1(KEYINPUT46), .A2(n1126), .ZN(n1125) );
NAND2_X1 U798 ( .A1(n1127), .A2(n1128), .ZN(n1124) );
NAND2_X1 U799 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U800 ( .A1(G900), .A2(G953), .ZN(n1130) );
NAND2_X1 U801 ( .A1(n1131), .A2(n1122), .ZN(n1129) );
OR3_X1 U802 ( .A1(n1126), .A2(KEYINPUT46), .A3(n1127), .ZN(n1123) );
XOR2_X1 U803 ( .A(n1132), .B(n1133), .Z(n1127) );
XNOR2_X1 U804 ( .A(n1134), .B(n1135), .ZN(n1133) );
XOR2_X1 U805 ( .A(n1136), .B(n1137), .Z(n1132) );
NAND2_X1 U806 ( .A1(KEYINPUT54), .A2(n1138), .ZN(n1136) );
OR2_X1 U807 ( .A1(G953), .A2(n1131), .ZN(n1126) );
XOR2_X1 U808 ( .A(n1139), .B(n1140), .Z(G69) );
NOR2_X1 U809 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
AND3_X1 U810 ( .A1(G953), .A2(G224), .A3(G898), .ZN(n1142) );
NOR2_X1 U811 ( .A1(G953), .A2(n1143), .ZN(n1141) );
NOR2_X1 U812 ( .A1(n1144), .A2(KEYINPUT53), .ZN(n1143) );
NOR2_X1 U813 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NOR2_X1 U814 ( .A1(n1147), .A2(n1148), .ZN(n1139) );
NOR2_X1 U815 ( .A1(G898), .A2(n1122), .ZN(n1147) );
NOR2_X1 U816 ( .A1(n1149), .A2(n1150), .ZN(G66) );
XOR2_X1 U817 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U818 ( .A1(n1118), .A2(n1153), .ZN(n1152) );
NAND2_X1 U819 ( .A1(n1154), .A2(KEYINPUT59), .ZN(n1151) );
NOR2_X1 U820 ( .A1(n1149), .A2(n1155), .ZN(G63) );
XOR2_X1 U821 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U822 ( .A1(n1158), .A2(G478), .ZN(n1156) );
NOR2_X1 U823 ( .A1(n1149), .A2(n1159), .ZN(G60) );
XOR2_X1 U824 ( .A(n1160), .B(n1161), .Z(n1159) );
XNOR2_X1 U825 ( .A(KEYINPUT6), .B(n1162), .ZN(n1161) );
NOR2_X1 U826 ( .A1(n1163), .A2(KEYINPUT41), .ZN(n1162) );
NOR2_X1 U827 ( .A1(n1164), .A2(n1153), .ZN(n1163) );
XOR2_X1 U828 ( .A(G104), .B(n1165), .Z(G6) );
NOR4_X1 U829 ( .A1(KEYINPUT58), .A2(n1083), .A3(n1166), .A4(n1167), .ZN(n1165) );
NOR3_X1 U830 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(G57) );
AND2_X1 U831 ( .A1(KEYINPUT25), .A2(n1149), .ZN(n1170) );
NOR3_X1 U832 ( .A1(KEYINPUT25), .A2(G953), .A3(G952), .ZN(n1169) );
XOR2_X1 U833 ( .A(n1171), .B(n1172), .Z(n1168) );
XOR2_X1 U834 ( .A(n1173), .B(n1174), .Z(n1172) );
NAND2_X1 U835 ( .A1(KEYINPUT39), .A2(n1175), .ZN(n1174) );
NAND2_X1 U836 ( .A1(n1158), .A2(G472), .ZN(n1173) );
NOR2_X1 U837 ( .A1(n1149), .A2(n1176), .ZN(G54) );
NOR3_X1 U838 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1176) );
AND2_X1 U839 ( .A1(n1180), .A2(KEYINPUT48), .ZN(n1179) );
NOR3_X1 U840 ( .A1(KEYINPUT48), .A2(n1181), .A3(n1180), .ZN(n1178) );
INV_X1 U841 ( .A(n1182), .ZN(n1180) );
NOR3_X1 U842 ( .A1(n1153), .A2(KEYINPUT56), .A3(n1183), .ZN(n1181) );
NOR3_X1 U843 ( .A1(n1153), .A2(n1184), .A3(n1183), .ZN(n1177) );
INV_X1 U844 ( .A(G469), .ZN(n1183) );
NOR2_X1 U845 ( .A1(n1185), .A2(KEYINPUT48), .ZN(n1184) );
NOR2_X1 U846 ( .A1(KEYINPUT56), .A2(n1182), .ZN(n1185) );
XNOR2_X1 U847 ( .A(n1186), .B(n1187), .ZN(n1182) );
XNOR2_X1 U848 ( .A(n1188), .B(n1189), .ZN(n1187) );
NOR2_X1 U849 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U850 ( .A1(n1149), .A2(n1192), .ZN(G51) );
XOR2_X1 U851 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U852 ( .A(n1195), .B(n1148), .Z(n1194) );
XOR2_X1 U853 ( .A(n1196), .B(n1197), .Z(n1193) );
XOR2_X1 U854 ( .A(n1198), .B(n1199), .Z(n1197) );
NOR2_X1 U855 ( .A1(KEYINPUT13), .A2(n1200), .ZN(n1199) );
NAND2_X1 U856 ( .A1(n1158), .A2(n1201), .ZN(n1196) );
INV_X1 U857 ( .A(n1153), .ZN(n1158) );
NAND2_X1 U858 ( .A1(G902), .A2(n1069), .ZN(n1153) );
NAND3_X1 U859 ( .A1(n1202), .A2(n1203), .A3(n1131), .ZN(n1069) );
AND4_X1 U860 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1131) );
AND3_X1 U861 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1207) );
NAND2_X1 U862 ( .A1(n1108), .A2(n1211), .ZN(n1206) );
NAND2_X1 U863 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XNOR2_X1 U864 ( .A(n1214), .B(KEYINPUT2), .ZN(n1212) );
NAND2_X1 U865 ( .A1(n1095), .A2(n1215), .ZN(n1204) );
NAND2_X1 U866 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND4_X1 U867 ( .A1(n1218), .A2(n1090), .A3(n1219), .A4(n1220), .ZN(n1217) );
XOR2_X1 U868 ( .A(KEYINPUT44), .B(n1221), .Z(n1220) );
NOR2_X1 U869 ( .A1(n1222), .A2(n1223), .ZN(n1219) );
NAND3_X1 U870 ( .A1(n1224), .A2(n1100), .A3(n1225), .ZN(n1216) );
XOR2_X1 U871 ( .A(n1226), .B(KEYINPUT63), .Z(n1225) );
XNOR2_X1 U872 ( .A(KEYINPUT43), .B(n1145), .ZN(n1203) );
NAND4_X1 U873 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1145) );
NAND4_X1 U874 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1227) );
OR2_X1 U875 ( .A1(n1224), .A2(KEYINPUT19), .ZN(n1234) );
NAND2_X1 U876 ( .A1(KEYINPUT19), .A2(n1235), .ZN(n1233) );
NAND3_X1 U877 ( .A1(n1221), .A2(n1236), .A3(n1237), .ZN(n1235) );
INV_X1 U878 ( .A(n1085), .ZN(n1221) );
INV_X1 U879 ( .A(n1146), .ZN(n1202) );
NAND3_X1 U880 ( .A1(n1238), .A2(n1064), .A3(n1239), .ZN(n1146) );
NAND2_X1 U881 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NAND2_X1 U882 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND2_X1 U883 ( .A1(n1100), .A2(n1244), .ZN(n1243) );
NAND2_X1 U884 ( .A1(n1232), .A2(n1091), .ZN(n1242) );
NAND3_X1 U885 ( .A1(n1240), .A2(n1244), .A3(n1099), .ZN(n1064) );
NOR2_X1 U886 ( .A1(n1122), .A2(G952), .ZN(n1149) );
XOR2_X1 U887 ( .A(G146), .B(n1245), .Z(G48) );
NOR2_X1 U888 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XOR2_X1 U889 ( .A(n1248), .B(n1249), .Z(G45) );
NAND4_X1 U890 ( .A1(n1250), .A2(n1090), .A3(n1095), .A4(n1251), .ZN(n1249) );
XOR2_X1 U891 ( .A(KEYINPUT10), .B(n1222), .Z(n1251) );
NAND2_X1 U892 ( .A1(n1252), .A2(n1253), .ZN(G42) );
NAND2_X1 U893 ( .A1(G140), .A2(n1205), .ZN(n1253) );
XOR2_X1 U894 ( .A(KEYINPUT51), .B(n1254), .Z(n1252) );
NOR2_X1 U895 ( .A1(G140), .A2(n1205), .ZN(n1254) );
NAND3_X1 U896 ( .A1(n1091), .A2(n1108), .A3(n1255), .ZN(n1205) );
XOR2_X1 U897 ( .A(n1256), .B(n1257), .Z(G39) );
NOR2_X1 U898 ( .A1(G137), .A2(KEYINPUT31), .ZN(n1257) );
NAND2_X1 U899 ( .A1(n1214), .A2(n1108), .ZN(n1256) );
AND3_X1 U900 ( .A1(n1095), .A2(n1232), .A3(n1258), .ZN(n1214) );
NOR3_X1 U901 ( .A1(n1259), .A2(n1260), .A3(n1222), .ZN(n1258) );
INV_X1 U902 ( .A(n1226), .ZN(n1222) );
XNOR2_X1 U903 ( .A(G134), .B(n1208), .ZN(G36) );
NAND4_X1 U904 ( .A1(n1095), .A2(n1090), .A3(n1261), .A4(n1108), .ZN(n1208) );
AND2_X1 U905 ( .A1(n1226), .A2(n1099), .ZN(n1261) );
XOR2_X1 U906 ( .A(n1138), .B(n1262), .Z(G33) );
NAND2_X1 U907 ( .A1(n1108), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U908 ( .A(KEYINPUT23), .B(n1213), .ZN(n1263) );
NAND2_X1 U909 ( .A1(n1255), .A2(n1090), .ZN(n1213) );
INV_X1 U910 ( .A(n1247), .ZN(n1255) );
NAND3_X1 U911 ( .A1(n1100), .A2(n1226), .A3(n1095), .ZN(n1247) );
XNOR2_X1 U912 ( .A(n1264), .B(KEYINPUT5), .ZN(n1095) );
NOR2_X1 U913 ( .A1(n1086), .A2(n1265), .ZN(n1108) );
INV_X1 U914 ( .A(n1087), .ZN(n1265) );
NAND2_X1 U915 ( .A1(n1266), .A2(n1267), .ZN(G30) );
NAND2_X1 U916 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND2_X1 U917 ( .A1(G128), .A2(n1270), .ZN(n1266) );
NAND2_X1 U918 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND2_X1 U919 ( .A1(KEYINPUT8), .A2(n1273), .ZN(n1272) );
INV_X1 U920 ( .A(n1210), .ZN(n1273) );
OR2_X1 U921 ( .A1(n1268), .A2(KEYINPUT8), .ZN(n1271) );
NOR2_X1 U922 ( .A1(KEYINPUT35), .A2(n1210), .ZN(n1268) );
NAND4_X1 U923 ( .A1(n1224), .A2(n1099), .A3(n1264), .A4(n1226), .ZN(n1210) );
INV_X1 U924 ( .A(n1246), .ZN(n1224) );
XOR2_X1 U925 ( .A(n1274), .B(n1238), .Z(G3) );
NAND3_X1 U926 ( .A1(n1090), .A2(n1240), .A3(n1232), .ZN(n1238) );
INV_X1 U927 ( .A(n1166), .ZN(n1240) );
NAND3_X1 U928 ( .A1(n1264), .A2(n1275), .A3(n1276), .ZN(n1166) );
XOR2_X1 U929 ( .A(n1200), .B(n1209), .Z(G27) );
NAND4_X1 U930 ( .A1(n1085), .A2(n1226), .A3(n1091), .A4(n1277), .ZN(n1209) );
NOR2_X1 U931 ( .A1(n1079), .A2(n1167), .ZN(n1277) );
INV_X1 U932 ( .A(n1278), .ZN(n1079) );
NAND2_X1 U933 ( .A1(n1071), .A2(n1279), .ZN(n1226) );
NAND4_X1 U934 ( .A1(G902), .A2(G953), .A3(n1280), .A4(n1281), .ZN(n1279) );
INV_X1 U935 ( .A(G900), .ZN(n1281) );
XNOR2_X1 U936 ( .A(G122), .B(n1228), .ZN(G24) );
NAND3_X1 U937 ( .A1(n1231), .A2(n1244), .A3(n1250), .ZN(n1228) );
AND3_X1 U938 ( .A1(n1085), .A2(n1107), .A3(n1218), .ZN(n1250) );
XOR2_X1 U939 ( .A(n1282), .B(KEYINPUT18), .Z(n1218) );
INV_X1 U940 ( .A(n1223), .ZN(n1107) );
INV_X1 U941 ( .A(n1083), .ZN(n1244) );
NAND2_X1 U942 ( .A1(n1260), .A2(n1259), .ZN(n1083) );
XOR2_X1 U943 ( .A(G119), .B(n1283), .Z(G21) );
NOR3_X1 U944 ( .A1(n1284), .A2(n1246), .A3(n1075), .ZN(n1283) );
NAND3_X1 U945 ( .A1(n1085), .A2(n1236), .A3(n1237), .ZN(n1246) );
XNOR2_X1 U946 ( .A(G116), .B(n1229), .ZN(G18) );
NAND4_X1 U947 ( .A1(n1231), .A2(n1090), .A3(n1085), .A4(n1099), .ZN(n1229) );
NOR2_X1 U948 ( .A1(n1282), .A2(n1223), .ZN(n1099) );
XOR2_X1 U949 ( .A(n1285), .B(KEYINPUT0), .Z(n1085) );
XOR2_X1 U950 ( .A(n1286), .B(n1230), .Z(G15) );
NAND4_X1 U951 ( .A1(n1231), .A2(n1090), .A3(n1100), .A4(n1276), .ZN(n1230) );
INV_X1 U952 ( .A(n1167), .ZN(n1100) );
NAND2_X1 U953 ( .A1(n1223), .A2(n1282), .ZN(n1167) );
NOR2_X1 U954 ( .A1(n1259), .A2(n1236), .ZN(n1090) );
INV_X1 U955 ( .A(n1237), .ZN(n1259) );
INV_X1 U956 ( .A(n1284), .ZN(n1231) );
NAND2_X1 U957 ( .A1(n1278), .A2(n1275), .ZN(n1284) );
NOR2_X1 U958 ( .A1(n1096), .A2(n1114), .ZN(n1278) );
INV_X1 U959 ( .A(n1097), .ZN(n1114) );
XNOR2_X1 U960 ( .A(G110), .B(n1287), .ZN(G12) );
NAND4_X1 U961 ( .A1(n1288), .A2(n1275), .A3(n1264), .A4(n1289), .ZN(n1287) );
AND2_X1 U962 ( .A1(n1091), .A2(n1232), .ZN(n1289) );
INV_X1 U963 ( .A(n1075), .ZN(n1232) );
NAND2_X1 U964 ( .A1(n1223), .A2(n1290), .ZN(n1075) );
INV_X1 U965 ( .A(n1282), .ZN(n1290) );
NAND3_X1 U966 ( .A1(n1291), .A2(n1292), .A3(n1102), .ZN(n1282) );
NAND3_X1 U967 ( .A1(n1164), .A2(n1293), .A3(n1160), .ZN(n1102) );
NAND2_X1 U968 ( .A1(KEYINPUT26), .A2(n1164), .ZN(n1292) );
INV_X1 U969 ( .A(G475), .ZN(n1164) );
NAND2_X1 U970 ( .A1(n1113), .A2(n1294), .ZN(n1291) );
INV_X1 U971 ( .A(KEYINPUT26), .ZN(n1294) );
AND2_X1 U972 ( .A1(G475), .A2(n1295), .ZN(n1113) );
NAND2_X1 U973 ( .A1(n1160), .A2(n1293), .ZN(n1295) );
XOR2_X1 U974 ( .A(n1296), .B(n1297), .Z(n1160) );
XOR2_X1 U975 ( .A(G122), .B(G113), .Z(n1297) );
XNOR2_X1 U976 ( .A(n1298), .B(n1299), .ZN(n1296) );
NOR2_X1 U977 ( .A1(G104), .A2(KEYINPUT1), .ZN(n1299) );
NOR2_X1 U978 ( .A1(KEYINPUT49), .A2(n1300), .ZN(n1298) );
XOR2_X1 U979 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U980 ( .A(n1303), .B(n1304), .Z(n1302) );
NOR2_X1 U981 ( .A1(KEYINPUT45), .A2(n1305), .ZN(n1304) );
AND2_X1 U982 ( .A1(n1306), .A2(G214), .ZN(n1303) );
XOR2_X1 U983 ( .A(n1307), .B(G143), .Z(n1301) );
NAND2_X1 U984 ( .A1(n1308), .A2(n1138), .ZN(n1307) );
XNOR2_X1 U985 ( .A(KEYINPUT52), .B(KEYINPUT28), .ZN(n1308) );
XOR2_X1 U986 ( .A(n1309), .B(n1310), .Z(n1223) );
XOR2_X1 U987 ( .A(KEYINPUT36), .B(G478), .Z(n1310) );
NAND2_X1 U988 ( .A1(n1157), .A2(n1293), .ZN(n1309) );
XNOR2_X1 U989 ( .A(n1311), .B(n1312), .ZN(n1157) );
XNOR2_X1 U990 ( .A(n1313), .B(n1314), .ZN(n1312) );
NAND2_X1 U991 ( .A1(KEYINPUT37), .A2(n1315), .ZN(n1313) );
XOR2_X1 U992 ( .A(G128), .B(n1316), .Z(n1315) );
XOR2_X1 U993 ( .A(G143), .B(G134), .Z(n1316) );
XOR2_X1 U994 ( .A(n1317), .B(G122), .Z(n1311) );
NAND2_X1 U995 ( .A1(G217), .A2(n1318), .ZN(n1317) );
NOR2_X1 U996 ( .A1(n1237), .A2(n1260), .ZN(n1091) );
INV_X1 U997 ( .A(n1236), .ZN(n1260) );
NAND2_X1 U998 ( .A1(n1319), .A2(n1320), .ZN(n1236) );
NAND2_X1 U999 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NAND2_X1 U1000 ( .A1(n1116), .A2(n1323), .ZN(n1322) );
INV_X1 U1001 ( .A(KEYINPUT61), .ZN(n1323) );
INV_X1 U1002 ( .A(n1118), .ZN(n1321) );
OR2_X1 U1003 ( .A1(n1101), .A2(KEYINPUT61), .ZN(n1319) );
NAND2_X1 U1004 ( .A1(n1116), .A2(n1118), .ZN(n1101) );
NAND2_X1 U1005 ( .A1(G217), .A2(n1324), .ZN(n1118) );
AND2_X1 U1006 ( .A1(n1154), .A2(n1293), .ZN(n1116) );
XOR2_X1 U1007 ( .A(n1325), .B(n1326), .Z(n1154) );
XOR2_X1 U1008 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1009 ( .A(n1329), .B(n1305), .ZN(n1328) );
XNOR2_X1 U1010 ( .A(n1330), .B(n1134), .ZN(n1305) );
XOR2_X1 U1011 ( .A(G125), .B(G140), .Z(n1134) );
XNOR2_X1 U1012 ( .A(G146), .B(KEYINPUT29), .ZN(n1330) );
NAND2_X1 U1013 ( .A1(KEYINPUT33), .A2(n1331), .ZN(n1329) );
XNOR2_X1 U1014 ( .A(G137), .B(n1332), .ZN(n1331) );
NAND2_X1 U1015 ( .A1(G221), .A2(n1318), .ZN(n1332) );
AND2_X1 U1016 ( .A1(G234), .A2(n1122), .ZN(n1318) );
XOR2_X1 U1017 ( .A(n1333), .B(n1334), .Z(n1325) );
XOR2_X1 U1018 ( .A(KEYINPUT22), .B(G128), .Z(n1334) );
INV_X1 U1019 ( .A(G119), .ZN(n1333) );
XNOR2_X1 U1020 ( .A(n1335), .B(n1111), .ZN(n1237) );
NAND2_X1 U1021 ( .A1(n1336), .A2(n1293), .ZN(n1111) );
XOR2_X1 U1022 ( .A(n1337), .B(n1175), .Z(n1336) );
XOR2_X1 U1023 ( .A(n1338), .B(n1274), .Z(n1175) );
NAND2_X1 U1024 ( .A1(G210), .A2(n1306), .ZN(n1338) );
NOR2_X1 U1025 ( .A1(G953), .A2(G237), .ZN(n1306) );
NOR2_X1 U1026 ( .A1(KEYINPUT12), .A2(n1171), .ZN(n1337) );
XOR2_X1 U1027 ( .A(n1339), .B(n1340), .Z(n1171) );
XOR2_X1 U1028 ( .A(KEYINPUT42), .B(n1341), .Z(n1340) );
NOR2_X1 U1029 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
XOR2_X1 U1030 ( .A(n1344), .B(KEYINPUT57), .Z(n1343) );
NAND2_X1 U1031 ( .A1(n1345), .A2(n1286), .ZN(n1344) );
INV_X1 U1032 ( .A(G113), .ZN(n1286) );
NOR2_X1 U1033 ( .A1(n1345), .A2(n1346), .ZN(n1342) );
XOR2_X1 U1034 ( .A(KEYINPUT62), .B(G113), .Z(n1346) );
XOR2_X1 U1035 ( .A(G116), .B(n1347), .Z(n1345) );
XOR2_X1 U1036 ( .A(KEYINPUT3), .B(G119), .Z(n1347) );
XOR2_X1 U1037 ( .A(n1195), .B(n1348), .Z(n1339) );
NAND2_X1 U1038 ( .A1(KEYINPUT7), .A2(n1112), .ZN(n1335) );
XOR2_X1 U1039 ( .A(G472), .B(KEYINPUT30), .Z(n1112) );
AND2_X1 U1040 ( .A1(n1096), .A2(n1097), .ZN(n1264) );
NAND2_X1 U1041 ( .A1(G221), .A2(n1324), .ZN(n1097) );
NAND2_X1 U1042 ( .A1(G234), .A2(n1293), .ZN(n1324) );
NAND2_X1 U1043 ( .A1(n1349), .A2(n1350), .ZN(n1096) );
OR2_X1 U1044 ( .A1(n1109), .A2(G469), .ZN(n1350) );
XOR2_X1 U1045 ( .A(n1351), .B(KEYINPUT21), .Z(n1349) );
NAND2_X1 U1046 ( .A1(G469), .A2(n1109), .ZN(n1351) );
NAND2_X1 U1047 ( .A1(n1352), .A2(n1293), .ZN(n1109) );
XOR2_X1 U1048 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1049 ( .A(n1355), .B(n1188), .Z(n1354) );
NAND2_X1 U1050 ( .A1(G227), .A2(n1356), .ZN(n1188) );
XOR2_X1 U1051 ( .A(KEYINPUT9), .B(G953), .Z(n1356) );
NAND3_X1 U1052 ( .A1(n1357), .A2(n1358), .A3(n1359), .ZN(n1355) );
INV_X1 U1053 ( .A(n1190), .ZN(n1359) );
NOR3_X1 U1054 ( .A1(n1135), .A2(n1360), .A3(n1348), .ZN(n1190) );
NAND2_X1 U1055 ( .A1(n1361), .A2(n1362), .ZN(n1358) );
INV_X1 U1056 ( .A(KEYINPUT55), .ZN(n1362) );
XOR2_X1 U1057 ( .A(n1363), .B(n1348), .Z(n1361) );
NAND2_X1 U1058 ( .A1(n1360), .A2(n1135), .ZN(n1363) );
NAND2_X1 U1059 ( .A1(KEYINPUT55), .A2(n1191), .ZN(n1357) );
NAND2_X1 U1060 ( .A1(n1364), .A2(n1365), .ZN(n1191) );
NAND2_X1 U1061 ( .A1(n1348), .A2(n1366), .ZN(n1365) );
XOR2_X1 U1062 ( .A(n1360), .B(n1135), .Z(n1366) );
INV_X1 U1063 ( .A(n1367), .ZN(n1348) );
NAND3_X1 U1064 ( .A1(n1135), .A2(n1360), .A3(n1367), .ZN(n1364) );
XOR2_X1 U1065 ( .A(n1138), .B(n1137), .Z(n1367) );
XOR2_X1 U1066 ( .A(G134), .B(G137), .Z(n1137) );
INV_X1 U1067 ( .A(G131), .ZN(n1138) );
XNOR2_X1 U1068 ( .A(n1368), .B(n1274), .ZN(n1360) );
INV_X1 U1069 ( .A(G101), .ZN(n1274) );
NAND2_X1 U1070 ( .A1(KEYINPUT27), .A2(n1369), .ZN(n1368) );
XOR2_X1 U1071 ( .A(G104), .B(n1370), .Z(n1369) );
NOR2_X1 U1072 ( .A1(G107), .A2(KEYINPUT17), .ZN(n1370) );
XOR2_X1 U1073 ( .A(n1371), .B(n1372), .Z(n1135) );
NOR2_X1 U1074 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
NOR3_X1 U1075 ( .A1(KEYINPUT15), .A2(G146), .A3(n1248), .ZN(n1374) );
INV_X1 U1076 ( .A(G143), .ZN(n1248) );
NOR2_X1 U1077 ( .A1(n1375), .A2(n1376), .ZN(n1373) );
INV_X1 U1078 ( .A(KEYINPUT15), .ZN(n1376) );
XOR2_X1 U1079 ( .A(n1269), .B(KEYINPUT11), .Z(n1371) );
INV_X1 U1080 ( .A(G128), .ZN(n1269) );
NOR2_X1 U1081 ( .A1(KEYINPUT50), .A2(n1186), .ZN(n1353) );
XOR2_X1 U1082 ( .A(G140), .B(n1327), .Z(n1186) );
NAND2_X1 U1083 ( .A1(n1071), .A2(n1377), .ZN(n1275) );
NAND4_X1 U1084 ( .A1(G902), .A2(G953), .A3(n1280), .A4(n1378), .ZN(n1377) );
INV_X1 U1085 ( .A(G898), .ZN(n1378) );
NAND3_X1 U1086 ( .A1(n1280), .A2(n1122), .A3(G952), .ZN(n1071) );
NAND2_X1 U1087 ( .A1(G237), .A2(G234), .ZN(n1280) );
XOR2_X1 U1088 ( .A(KEYINPUT60), .B(n1276), .Z(n1288) );
INV_X1 U1089 ( .A(n1285), .ZN(n1276) );
NAND2_X1 U1090 ( .A1(n1086), .A2(n1087), .ZN(n1285) );
NAND2_X1 U1091 ( .A1(G214), .A2(n1379), .ZN(n1087) );
XNOR2_X1 U1092 ( .A(n1380), .B(n1201), .ZN(n1086) );
AND2_X1 U1093 ( .A1(G210), .A2(n1379), .ZN(n1201) );
NAND2_X1 U1094 ( .A1(n1381), .A2(n1293), .ZN(n1379) );
INV_X1 U1095 ( .A(G237), .ZN(n1381) );
NAND3_X1 U1096 ( .A1(n1382), .A2(n1383), .A3(n1293), .ZN(n1380) );
INV_X1 U1097 ( .A(G902), .ZN(n1293) );
NAND2_X1 U1098 ( .A1(n1384), .A2(n1385), .ZN(n1383) );
NAND2_X1 U1099 ( .A1(n1386), .A2(n1387), .ZN(n1384) );
NAND2_X1 U1100 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
INV_X1 U1101 ( .A(KEYINPUT40), .ZN(n1389) );
NAND2_X1 U1102 ( .A1(KEYINPUT40), .A2(n1148), .ZN(n1386) );
OR2_X1 U1103 ( .A1(n1385), .A2(n1388), .ZN(n1382) );
NAND2_X1 U1104 ( .A1(KEYINPUT47), .A2(n1148), .ZN(n1388) );
XOR2_X1 U1105 ( .A(n1390), .B(n1391), .Z(n1148) );
XOR2_X1 U1106 ( .A(G104), .B(n1392), .Z(n1391) );
XOR2_X1 U1107 ( .A(G119), .B(G113), .Z(n1392) );
XOR2_X1 U1108 ( .A(n1393), .B(n1314), .Z(n1390) );
XOR2_X1 U1109 ( .A(G107), .B(G116), .Z(n1314) );
XOR2_X1 U1110 ( .A(n1394), .B(G101), .Z(n1393) );
NAND3_X1 U1111 ( .A1(n1395), .A2(n1396), .A3(n1397), .ZN(n1394) );
NAND2_X1 U1112 ( .A1(KEYINPUT16), .A2(n1327), .ZN(n1397) );
OR3_X1 U1113 ( .A1(n1327), .A2(KEYINPUT16), .A3(G122), .ZN(n1396) );
INV_X1 U1114 ( .A(n1398), .ZN(n1327) );
NAND2_X1 U1115 ( .A1(G122), .A2(n1399), .ZN(n1395) );
NAND2_X1 U1116 ( .A1(n1400), .A2(n1401), .ZN(n1399) );
INV_X1 U1117 ( .A(KEYINPUT16), .ZN(n1401) );
XOR2_X1 U1118 ( .A(n1398), .B(KEYINPUT34), .Z(n1400) );
XNOR2_X1 U1119 ( .A(G110), .B(KEYINPUT14), .ZN(n1398) );
XOR2_X1 U1120 ( .A(n1195), .B(n1402), .Z(n1385) );
XOR2_X1 U1121 ( .A(n1200), .B(n1198), .Z(n1402) );
NAND2_X1 U1122 ( .A1(n1403), .A2(G224), .ZN(n1198) );
XOR2_X1 U1123 ( .A(n1122), .B(KEYINPUT38), .Z(n1403) );
INV_X1 U1124 ( .A(G953), .ZN(n1122) );
INV_X1 U1125 ( .A(G125), .ZN(n1200) );
XOR2_X1 U1126 ( .A(n1404), .B(G128), .Z(n1195) );
NAND2_X1 U1127 ( .A1(KEYINPUT4), .A2(n1375), .ZN(n1404) );
XOR2_X1 U1128 ( .A(G143), .B(G146), .Z(n1375) );
endmodule


