//Key = 1100101101010001011001101000000011100011111011100011110010111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401;

XNOR2_X1 U777 ( .A(G107), .B(n1064), .ZN(G9) );
NAND4_X1 U778 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1064) );
AND2_X1 U779 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XOR2_X1 U780 ( .A(KEYINPUT61), .B(n1071), .Z(n1065) );
NOR2_X1 U781 ( .A1(n1072), .A2(n1073), .ZN(G75) );
NOR4_X1 U782 ( .A1(G953), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1073) );
NOR3_X1 U783 ( .A1(n1077), .A2(KEYINPUT47), .A3(n1078), .ZN(n1075) );
INV_X1 U784 ( .A(n1079), .ZN(n1078) );
NOR2_X1 U785 ( .A1(n1080), .A2(n1081), .ZN(n1077) );
NOR4_X1 U786 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1081) );
NOR3_X1 U787 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1083) );
XOR2_X1 U788 ( .A(n1089), .B(KEYINPUT44), .Z(n1088) );
NOR2_X1 U789 ( .A1(n1090), .A2(n1091), .ZN(n1087) );
NOR2_X1 U790 ( .A1(n1069), .A2(n1092), .ZN(n1082) );
NOR2_X1 U791 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR3_X1 U792 ( .A1(n1094), .A2(n1095), .A3(n1086), .ZN(n1080) );
NOR2_X1 U793 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U794 ( .A1(n1098), .A2(n1084), .ZN(n1097) );
INV_X1 U795 ( .A(n1099), .ZN(n1084) );
NOR2_X1 U796 ( .A1(n1100), .A2(n1071), .ZN(n1098) );
AND2_X1 U797 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U798 ( .A1(n1103), .A2(n1085), .ZN(n1096) );
NOR2_X1 U799 ( .A1(n1070), .A2(n1104), .ZN(n1103) );
NOR3_X1 U800 ( .A1(n1074), .A2(G953), .A3(G952), .ZN(n1072) );
AND4_X1 U801 ( .A1(n1105), .A2(n1091), .A3(n1106), .A4(n1107), .ZN(n1074) );
NOR4_X1 U802 ( .A1(n1108), .A2(n1109), .A3(n1110), .A4(n1111), .ZN(n1107) );
XOR2_X1 U803 ( .A(KEYINPUT36), .B(n1112), .Z(n1109) );
NAND4_X1 U804 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1108) );
NAND2_X1 U805 ( .A1(KEYINPUT30), .A2(n1117), .ZN(n1116) );
NAND3_X1 U806 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1115) );
INV_X1 U807 ( .A(KEYINPUT30), .ZN(n1119) );
OR2_X1 U808 ( .A1(G478), .A2(KEYINPUT34), .ZN(n1114) );
NAND3_X1 U809 ( .A1(G478), .A2(n1121), .A3(KEYINPUT34), .ZN(n1113) );
NOR3_X1 U810 ( .A1(n1102), .A2(n1122), .A3(n1123), .ZN(n1106) );
XOR2_X1 U811 ( .A(n1124), .B(n1125), .Z(n1105) );
NOR2_X1 U812 ( .A1(n1126), .A2(KEYINPUT37), .ZN(n1125) );
INV_X1 U813 ( .A(n1127), .ZN(n1126) );
XOR2_X1 U814 ( .A(n1128), .B(n1129), .Z(G72) );
NOR2_X1 U815 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U816 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XNOR2_X1 U817 ( .A(n1134), .B(KEYINPUT31), .ZN(n1133) );
INV_X1 U818 ( .A(n1135), .ZN(n1132) );
NOR2_X1 U819 ( .A1(n1134), .A2(n1135), .ZN(n1130) );
NAND2_X1 U820 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U821 ( .A1(n1138), .A2(G953), .ZN(n1137) );
XOR2_X1 U822 ( .A(n1139), .B(n1140), .Z(n1136) );
XOR2_X1 U823 ( .A(n1141), .B(n1142), .Z(n1140) );
XNOR2_X1 U824 ( .A(n1143), .B(n1144), .ZN(n1139) );
NOR2_X1 U825 ( .A1(KEYINPUT23), .A2(n1145), .ZN(n1144) );
NOR2_X1 U826 ( .A1(G953), .A2(n1146), .ZN(n1134) );
NAND2_X1 U827 ( .A1(G953), .A2(n1147), .ZN(n1128) );
NAND2_X1 U828 ( .A1(G900), .A2(G227), .ZN(n1147) );
XOR2_X1 U829 ( .A(n1148), .B(n1149), .Z(G69) );
XOR2_X1 U830 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U831 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U832 ( .A1(n1154), .A2(n1155), .ZN(n1150) );
NAND3_X1 U833 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1155) );
XNOR2_X1 U834 ( .A(KEYINPUT33), .B(n1159), .ZN(n1156) );
XOR2_X1 U835 ( .A(KEYINPUT38), .B(G953), .Z(n1154) );
NAND2_X1 U836 ( .A1(G953), .A2(n1160), .ZN(n1148) );
NAND2_X1 U837 ( .A1(G898), .A2(G224), .ZN(n1160) );
NOR2_X1 U838 ( .A1(n1161), .A2(n1162), .ZN(G66) );
NOR3_X1 U839 ( .A1(n1163), .A2(n1124), .A3(n1164), .ZN(n1162) );
NOR2_X1 U840 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
AND2_X1 U841 ( .A1(n1076), .A2(G217), .ZN(n1165) );
XOR2_X1 U842 ( .A(n1167), .B(KEYINPUT62), .Z(n1163) );
NAND3_X1 U843 ( .A1(G217), .A2(n1166), .A3(n1168), .ZN(n1167) );
NOR2_X1 U844 ( .A1(n1161), .A2(n1169), .ZN(G63) );
XOR2_X1 U845 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U846 ( .A1(n1168), .A2(G478), .ZN(n1171) );
NOR2_X1 U847 ( .A1(n1172), .A2(n1173), .ZN(G60) );
XOR2_X1 U848 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND2_X1 U849 ( .A1(n1168), .A2(G475), .ZN(n1174) );
NOR2_X1 U850 ( .A1(n1176), .A2(n1177), .ZN(n1172) );
XOR2_X1 U851 ( .A(KEYINPUT43), .B(G952), .Z(n1177) );
XOR2_X1 U852 ( .A(KEYINPUT16), .B(n1178), .Z(n1176) );
XOR2_X1 U853 ( .A(G104), .B(n1179), .Z(G6) );
NOR2_X1 U854 ( .A1(n1161), .A2(n1180), .ZN(G57) );
NOR2_X1 U855 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U856 ( .A(KEYINPUT20), .B(n1183), .Z(n1182) );
NOR2_X1 U857 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
XOR2_X1 U858 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U859 ( .A1(n1188), .A2(n1189), .ZN(n1181) );
XOR2_X1 U860 ( .A(n1190), .B(n1187), .Z(n1189) );
XOR2_X1 U861 ( .A(n1191), .B(n1192), .Z(n1187) );
NAND2_X1 U862 ( .A1(n1168), .A2(G472), .ZN(n1191) );
INV_X1 U863 ( .A(n1186), .ZN(n1190) );
INV_X1 U864 ( .A(n1184), .ZN(n1188) );
XNOR2_X1 U865 ( .A(G101), .B(n1193), .ZN(n1184) );
NOR2_X1 U866 ( .A1(KEYINPUT48), .A2(n1194), .ZN(n1193) );
NOR2_X1 U867 ( .A1(n1195), .A2(n1196), .ZN(G54) );
XNOR2_X1 U868 ( .A(n1161), .B(KEYINPUT17), .ZN(n1196) );
XOR2_X1 U869 ( .A(n1197), .B(n1198), .Z(n1195) );
XOR2_X1 U870 ( .A(n1199), .B(n1200), .Z(n1198) );
NAND2_X1 U871 ( .A1(n1201), .A2(KEYINPUT22), .ZN(n1199) );
XOR2_X1 U872 ( .A(n1202), .B(n1203), .Z(n1201) );
NAND2_X1 U873 ( .A1(G227), .A2(n1178), .ZN(n1202) );
XOR2_X1 U874 ( .A(n1204), .B(n1205), .Z(n1197) );
NOR3_X1 U875 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1205) );
NOR2_X1 U876 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
INV_X1 U877 ( .A(KEYINPUT1), .ZN(n1210) );
NOR2_X1 U878 ( .A1(n1211), .A2(n1212), .ZN(n1209) );
NOR3_X1 U879 ( .A1(n1213), .A2(n1214), .A3(n1141), .ZN(n1212) );
NOR2_X1 U880 ( .A1(KEYINPUT40), .A2(n1215), .ZN(n1211) );
NOR2_X1 U881 ( .A1(KEYINPUT1), .A2(n1216), .ZN(n1207) );
NOR2_X1 U882 ( .A1(n1217), .A2(n1214), .ZN(n1216) );
XOR2_X1 U883 ( .A(n1213), .B(n1141), .Z(n1217) );
INV_X1 U884 ( .A(KEYINPUT40), .ZN(n1213) );
NAND2_X1 U885 ( .A1(KEYINPUT59), .A2(n1218), .ZN(n1204) );
NAND2_X1 U886 ( .A1(n1168), .A2(G469), .ZN(n1218) );
NOR3_X1 U887 ( .A1(n1161), .A2(n1219), .A3(n1220), .ZN(G51) );
NOR2_X1 U888 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NOR2_X1 U889 ( .A1(n1223), .A2(n1224), .ZN(n1221) );
NOR2_X1 U890 ( .A1(n1153), .A2(n1225), .ZN(n1224) );
NOR2_X1 U891 ( .A1(n1226), .A2(n1227), .ZN(n1223) );
NOR2_X1 U892 ( .A1(n1228), .A2(n1229), .ZN(n1219) );
NOR2_X1 U893 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NOR2_X1 U894 ( .A1(n1225), .A2(n1227), .ZN(n1231) );
XOR2_X1 U895 ( .A(n1226), .B(n1232), .Z(n1225) );
XOR2_X1 U896 ( .A(KEYINPUT3), .B(KEYINPUT0), .Z(n1232) );
NOR2_X1 U897 ( .A1(n1226), .A2(n1153), .ZN(n1230) );
AND2_X1 U898 ( .A1(n1168), .A2(n1120), .ZN(n1226) );
AND2_X1 U899 ( .A1(G902), .A2(n1076), .ZN(n1168) );
NAND4_X1 U900 ( .A1(n1233), .A2(n1146), .A3(n1158), .A4(n1159), .ZN(n1076) );
AND4_X1 U901 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1158) );
NOR4_X1 U902 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1179), .ZN(n1237) );
AND3_X1 U903 ( .A1(n1241), .A2(n1069), .A3(n1104), .ZN(n1179) );
NOR3_X1 U904 ( .A1(n1242), .A2(n1243), .A3(n1089), .ZN(n1239) );
NOR3_X1 U905 ( .A1(n1244), .A2(n1085), .A3(n1245), .ZN(n1243) );
NAND3_X1 U906 ( .A1(n1246), .A2(n1066), .A3(n1069), .ZN(n1244) );
INV_X1 U907 ( .A(KEYINPUT25), .ZN(n1242) );
NOR2_X1 U908 ( .A1(KEYINPUT25), .A2(n1247), .ZN(n1238) );
AND4_X1 U909 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1146) );
NOR4_X1 U910 ( .A1(n1252), .A2(n1253), .A3(n1254), .A4(n1255), .ZN(n1251) );
INV_X1 U911 ( .A(n1256), .ZN(n1255) );
NAND2_X1 U912 ( .A1(n1067), .A2(n1257), .ZN(n1250) );
NAND2_X1 U913 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NAND2_X1 U914 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XOR2_X1 U915 ( .A(KEYINPUT56), .B(n1262), .Z(n1258) );
XOR2_X1 U916 ( .A(n1157), .B(KEYINPUT12), .Z(n1233) );
NAND3_X1 U917 ( .A1(n1070), .A2(n1069), .A3(n1241), .ZN(n1157) );
INV_X1 U918 ( .A(n1222), .ZN(n1228) );
NAND2_X1 U919 ( .A1(KEYINPUT39), .A2(n1263), .ZN(n1222) );
XOR2_X1 U920 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U921 ( .A(n1266), .B(n1267), .Z(n1265) );
NOR2_X1 U922 ( .A1(KEYINPUT26), .A2(n1268), .ZN(n1267) );
INV_X1 U923 ( .A(G125), .ZN(n1268) );
NOR2_X1 U924 ( .A1(n1269), .A2(G952), .ZN(n1161) );
XNOR2_X1 U925 ( .A(KEYINPUT16), .B(G953), .ZN(n1269) );
XOR2_X1 U926 ( .A(n1270), .B(n1271), .Z(G48) );
NAND2_X1 U927 ( .A1(n1262), .A2(n1067), .ZN(n1271) );
AND2_X1 U928 ( .A1(n1272), .A2(n1104), .ZN(n1262) );
XNOR2_X1 U929 ( .A(G143), .B(n1248), .ZN(G45) );
NAND2_X1 U930 ( .A1(n1273), .A2(n1274), .ZN(n1248) );
XNOR2_X1 U931 ( .A(G140), .B(n1249), .ZN(G42) );
NAND3_X1 U932 ( .A1(n1275), .A2(n1071), .A3(n1261), .ZN(n1249) );
INV_X1 U933 ( .A(n1276), .ZN(n1261) );
XOR2_X1 U934 ( .A(G137), .B(n1254), .Z(G39) );
AND3_X1 U935 ( .A1(n1275), .A2(n1099), .A3(n1272), .ZN(n1254) );
XOR2_X1 U936 ( .A(G134), .B(n1253), .Z(G36) );
AND3_X1 U937 ( .A1(n1275), .A2(n1070), .A3(n1274), .ZN(n1253) );
XOR2_X1 U938 ( .A(G131), .B(n1252), .Z(G33) );
AND3_X1 U939 ( .A1(n1274), .A2(n1275), .A3(n1104), .ZN(n1252) );
INV_X1 U940 ( .A(n1094), .ZN(n1275) );
NAND2_X1 U941 ( .A1(n1277), .A2(n1091), .ZN(n1094) );
AND4_X1 U942 ( .A1(n1071), .A2(n1278), .A3(n1112), .A4(n1279), .ZN(n1274) );
NAND2_X1 U943 ( .A1(n1280), .A2(n1281), .ZN(G30) );
NAND2_X1 U944 ( .A1(n1282), .A2(n1256), .ZN(n1281) );
XOR2_X1 U945 ( .A(KEYINPUT11), .B(n1283), .Z(n1280) );
NOR2_X1 U946 ( .A1(n1282), .A2(n1256), .ZN(n1283) );
NAND3_X1 U947 ( .A1(n1070), .A2(n1067), .A3(n1272), .ZN(n1256) );
AND3_X1 U948 ( .A1(n1071), .A2(n1279), .A3(n1093), .ZN(n1272) );
NOR2_X1 U949 ( .A1(n1278), .A2(n1284), .ZN(n1093) );
XNOR2_X1 U950 ( .A(KEYINPUT7), .B(G128), .ZN(n1282) );
XNOR2_X1 U951 ( .A(G101), .B(n1159), .ZN(G3) );
NAND4_X1 U952 ( .A1(n1099), .A2(n1241), .A3(n1278), .A4(n1112), .ZN(n1159) );
XOR2_X1 U953 ( .A(G125), .B(n1285), .Z(G27) );
NOR3_X1 U954 ( .A1(n1276), .A2(n1286), .A3(n1089), .ZN(n1285) );
XOR2_X1 U955 ( .A(n1085), .B(KEYINPUT2), .Z(n1286) );
NAND4_X1 U956 ( .A1(n1287), .A2(n1104), .A3(n1284), .A4(n1279), .ZN(n1276) );
NAND2_X1 U957 ( .A1(n1288), .A2(n1289), .ZN(n1279) );
NAND4_X1 U958 ( .A1(n1138), .A2(G902), .A3(G953), .A4(n1079), .ZN(n1289) );
XNOR2_X1 U959 ( .A(G900), .B(KEYINPUT29), .ZN(n1138) );
NAND2_X1 U960 ( .A1(n1290), .A2(n1291), .ZN(G24) );
NAND2_X1 U961 ( .A1(G122), .A2(n1247), .ZN(n1291) );
XOR2_X1 U962 ( .A(KEYINPUT24), .B(n1292), .Z(n1290) );
NOR2_X1 U963 ( .A1(G122), .A2(n1247), .ZN(n1292) );
NAND4_X1 U964 ( .A1(n1260), .A2(n1273), .A3(n1069), .A4(n1066), .ZN(n1247) );
INV_X1 U965 ( .A(n1086), .ZN(n1069) );
NAND2_X1 U966 ( .A1(n1284), .A2(n1278), .ZN(n1086) );
NOR3_X1 U967 ( .A1(n1089), .A2(n1293), .A3(n1245), .ZN(n1273) );
NAND3_X1 U968 ( .A1(n1294), .A2(n1295), .A3(n1296), .ZN(G21) );
NAND2_X1 U969 ( .A1(n1240), .A2(n1297), .ZN(n1296) );
NAND2_X1 U970 ( .A1(n1298), .A2(n1299), .ZN(n1295) );
INV_X1 U971 ( .A(KEYINPUT21), .ZN(n1299) );
NAND2_X1 U972 ( .A1(G119), .A2(n1300), .ZN(n1298) );
XOR2_X1 U973 ( .A(KEYINPUT53), .B(n1240), .Z(n1300) );
INV_X1 U974 ( .A(n1301), .ZN(n1240) );
NAND2_X1 U975 ( .A1(KEYINPUT21), .A2(n1302), .ZN(n1294) );
NAND2_X1 U976 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
OR2_X1 U977 ( .A1(n1301), .A2(KEYINPUT53), .ZN(n1304) );
NAND3_X1 U978 ( .A1(G119), .A2(n1301), .A3(KEYINPUT53), .ZN(n1303) );
NAND3_X1 U979 ( .A1(n1287), .A2(n1099), .A3(n1305), .ZN(n1301) );
XNOR2_X1 U980 ( .A(G116), .B(n1236), .ZN(G18) );
NAND3_X1 U981 ( .A1(n1070), .A2(n1278), .A3(n1305), .ZN(n1236) );
NOR2_X1 U982 ( .A1(n1111), .A2(n1293), .ZN(n1070) );
XNOR2_X1 U983 ( .A(G113), .B(n1234), .ZN(G15) );
NAND3_X1 U984 ( .A1(n1104), .A2(n1278), .A3(n1305), .ZN(n1234) );
AND4_X1 U985 ( .A1(n1260), .A2(n1067), .A3(n1112), .A4(n1066), .ZN(n1305) );
INV_X1 U986 ( .A(n1284), .ZN(n1112) );
INV_X1 U987 ( .A(n1085), .ZN(n1260) );
NAND2_X1 U988 ( .A1(n1101), .A2(n1306), .ZN(n1085) );
INV_X1 U989 ( .A(n1287), .ZN(n1278) );
AND2_X1 U990 ( .A1(n1293), .A2(n1307), .ZN(n1104) );
XOR2_X1 U991 ( .A(KEYINPUT46), .B(n1245), .Z(n1307) );
XOR2_X1 U992 ( .A(n1111), .B(KEYINPUT58), .Z(n1245) );
XOR2_X1 U993 ( .A(n1235), .B(n1308), .Z(G12) );
NAND2_X1 U994 ( .A1(KEYINPUT42), .A2(G110), .ZN(n1308) );
NAND4_X1 U995 ( .A1(n1287), .A2(n1099), .A3(n1284), .A4(n1241), .ZN(n1235) );
AND3_X1 U996 ( .A1(n1071), .A2(n1066), .A3(n1067), .ZN(n1241) );
INV_X1 U997 ( .A(n1089), .ZN(n1067) );
NAND2_X1 U998 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U999 ( .A1(n1309), .A2(G214), .ZN(n1091) );
XOR2_X1 U1000 ( .A(n1310), .B(KEYINPUT14), .Z(n1309) );
INV_X1 U1001 ( .A(n1277), .ZN(n1090) );
NOR2_X1 U1002 ( .A1(n1123), .A2(n1311), .ZN(n1277) );
AND2_X1 U1003 ( .A1(n1120), .A2(n1118), .ZN(n1311) );
NOR2_X1 U1004 ( .A1(n1118), .A2(n1120), .ZN(n1123) );
INV_X1 U1005 ( .A(n1117), .ZN(n1120) );
NAND2_X1 U1006 ( .A1(G210), .A2(n1310), .ZN(n1117) );
NAND2_X1 U1007 ( .A1(n1312), .A2(n1313), .ZN(n1310) );
NAND2_X1 U1008 ( .A1(n1314), .A2(n1312), .ZN(n1118) );
XOR2_X1 U1009 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1010 ( .A(n1153), .B(n1264), .Z(n1316) );
INV_X1 U1011 ( .A(n1227), .ZN(n1153) );
XOR2_X1 U1012 ( .A(n1317), .B(n1318), .Z(n1227) );
XOR2_X1 U1013 ( .A(n1319), .B(n1320), .Z(n1318) );
XOR2_X1 U1014 ( .A(n1321), .B(n1322), .Z(n1317) );
XOR2_X1 U1015 ( .A(G113), .B(G101), .Z(n1322) );
NAND2_X1 U1016 ( .A1(n1323), .A2(KEYINPUT50), .ZN(n1321) );
XNOR2_X1 U1017 ( .A(n1324), .B(KEYINPUT54), .ZN(n1323) );
XOR2_X1 U1018 ( .A(G125), .B(n1266), .Z(n1315) );
AND2_X1 U1019 ( .A1(G224), .A2(n1178), .ZN(n1266) );
NAND2_X1 U1020 ( .A1(n1288), .A2(n1325), .ZN(n1066) );
NAND3_X1 U1021 ( .A1(n1152), .A2(n1079), .A3(G902), .ZN(n1325) );
NOR2_X1 U1022 ( .A1(n1178), .A2(G898), .ZN(n1152) );
NAND3_X1 U1023 ( .A1(n1079), .A2(n1178), .A3(G952), .ZN(n1288) );
NAND2_X1 U1024 ( .A1(G237), .A2(G234), .ZN(n1079) );
NOR2_X1 U1025 ( .A1(n1101), .A2(n1102), .ZN(n1071) );
INV_X1 U1026 ( .A(n1306), .ZN(n1102) );
NAND2_X1 U1027 ( .A1(G221), .A2(n1326), .ZN(n1306) );
NAND2_X1 U1028 ( .A1(G234), .A2(n1312), .ZN(n1326) );
XNOR2_X1 U1029 ( .A(n1110), .B(KEYINPUT13), .ZN(n1101) );
XNOR2_X1 U1030 ( .A(n1327), .B(G469), .ZN(n1110) );
NAND2_X1 U1031 ( .A1(n1328), .A2(n1312), .ZN(n1327) );
XOR2_X1 U1032 ( .A(n1329), .B(n1330), .Z(n1328) );
XNOR2_X1 U1033 ( .A(n1331), .B(n1203), .ZN(n1330) );
XOR2_X1 U1034 ( .A(G110), .B(G140), .Z(n1203) );
NAND3_X1 U1035 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1331) );
NAND2_X1 U1036 ( .A1(n1206), .A2(n1200), .ZN(n1334) );
AND2_X1 U1037 ( .A1(n1214), .A2(n1141), .ZN(n1206) );
OR3_X1 U1038 ( .A1(n1200), .A2(n1214), .A3(n1215), .ZN(n1333) );
NAND2_X1 U1039 ( .A1(n1335), .A2(n1215), .ZN(n1332) );
XOR2_X1 U1040 ( .A(n1200), .B(n1214), .Z(n1335) );
XOR2_X1 U1041 ( .A(G101), .B(n1324), .Z(n1214) );
XOR2_X1 U1042 ( .A(G104), .B(G107), .Z(n1324) );
XOR2_X1 U1043 ( .A(n1192), .B(KEYINPUT57), .Z(n1200) );
XOR2_X1 U1044 ( .A(n1336), .B(n1337), .Z(n1329) );
XOR2_X1 U1045 ( .A(KEYINPUT28), .B(KEYINPUT19), .Z(n1337) );
NOR2_X1 U1046 ( .A1(KEYINPUT10), .A2(n1338), .ZN(n1336) );
INV_X1 U1047 ( .A(G227), .ZN(n1338) );
XOR2_X1 U1048 ( .A(n1339), .B(G472), .Z(n1284) );
NAND2_X1 U1049 ( .A1(n1340), .A2(n1312), .ZN(n1339) );
XOR2_X1 U1050 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1051 ( .A(n1343), .B(n1186), .Z(n1342) );
XOR2_X1 U1052 ( .A(n1344), .B(n1264), .Z(n1186) );
XOR2_X1 U1053 ( .A(n1141), .B(KEYINPUT49), .Z(n1264) );
INV_X1 U1054 ( .A(n1215), .ZN(n1141) );
XOR2_X1 U1055 ( .A(n1270), .B(n1345), .Z(n1215) );
NAND3_X1 U1056 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1344) );
NAND2_X1 U1057 ( .A1(KEYINPUT5), .A2(n1349), .ZN(n1348) );
INV_X1 U1058 ( .A(n1350), .ZN(n1349) );
OR3_X1 U1059 ( .A1(n1351), .A2(KEYINPUT5), .A3(G113), .ZN(n1347) );
NAND2_X1 U1060 ( .A1(G113), .A2(n1351), .ZN(n1346) );
NAND2_X1 U1061 ( .A1(KEYINPUT41), .A2(n1350), .ZN(n1351) );
NAND2_X1 U1062 ( .A1(n1352), .A2(n1353), .ZN(n1350) );
NAND2_X1 U1063 ( .A1(G119), .A2(n1354), .ZN(n1353) );
NAND2_X1 U1064 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
NAND2_X1 U1065 ( .A1(KEYINPUT51), .A2(n1357), .ZN(n1356) );
INV_X1 U1066 ( .A(KEYINPUT9), .ZN(n1357) );
NAND3_X1 U1067 ( .A1(n1358), .A2(n1359), .A3(KEYINPUT9), .ZN(n1352) );
NAND2_X1 U1068 ( .A1(KEYINPUT51), .A2(n1360), .ZN(n1359) );
NAND2_X1 U1069 ( .A1(n1355), .A2(n1297), .ZN(n1360) );
OR2_X1 U1070 ( .A1(n1361), .A2(KEYINPUT51), .ZN(n1358) );
NAND2_X1 U1071 ( .A1(KEYINPUT18), .A2(n1192), .ZN(n1343) );
XNOR2_X1 U1072 ( .A(G131), .B(n1143), .ZN(n1192) );
XOR2_X1 U1073 ( .A(G134), .B(G137), .Z(n1143) );
XOR2_X1 U1074 ( .A(G101), .B(n1362), .Z(n1341) );
NOR2_X1 U1075 ( .A1(KEYINPUT55), .A2(n1194), .ZN(n1362) );
NAND3_X1 U1076 ( .A1(n1313), .A2(n1178), .A3(G210), .ZN(n1194) );
NOR2_X1 U1077 ( .A1(n1246), .A2(n1111), .ZN(n1099) );
XNOR2_X1 U1078 ( .A(n1363), .B(G475), .ZN(n1111) );
NAND2_X1 U1079 ( .A1(n1175), .A2(n1312), .ZN(n1363) );
XOR2_X1 U1080 ( .A(n1364), .B(n1365), .Z(n1175) );
XOR2_X1 U1081 ( .A(n1366), .B(n1367), .Z(n1365) );
NAND2_X1 U1082 ( .A1(KEYINPUT52), .A2(n1368), .ZN(n1367) );
NAND2_X1 U1083 ( .A1(n1369), .A2(n1370), .ZN(n1366) );
NAND2_X1 U1084 ( .A1(G146), .A2(n1142), .ZN(n1370) );
XOR2_X1 U1085 ( .A(KEYINPUT32), .B(n1371), .Z(n1369) );
NOR2_X1 U1086 ( .A1(G146), .A2(n1142), .ZN(n1371) );
XOR2_X1 U1087 ( .A(n1372), .B(n1373), .Z(n1364) );
XOR2_X1 U1088 ( .A(G113), .B(G104), .Z(n1373) );
NAND2_X1 U1089 ( .A1(KEYINPUT4), .A2(n1374), .ZN(n1372) );
XOR2_X1 U1090 ( .A(n1375), .B(n1376), .Z(n1374) );
XOR2_X1 U1091 ( .A(G143), .B(n1145), .Z(n1376) );
INV_X1 U1092 ( .A(G131), .ZN(n1145) );
NAND3_X1 U1093 ( .A1(n1313), .A2(n1178), .A3(n1377), .ZN(n1375) );
XNOR2_X1 U1094 ( .A(G214), .B(KEYINPUT15), .ZN(n1377) );
INV_X1 U1095 ( .A(G237), .ZN(n1313) );
INV_X1 U1096 ( .A(n1293), .ZN(n1246) );
NOR2_X1 U1097 ( .A1(n1122), .A2(n1378), .ZN(n1293) );
AND2_X1 U1098 ( .A1(G478), .A2(n1121), .ZN(n1378) );
NOR2_X1 U1099 ( .A1(n1121), .A2(G478), .ZN(n1122) );
NAND2_X1 U1100 ( .A1(n1312), .A2(n1170), .ZN(n1121) );
NAND2_X1 U1101 ( .A1(n1379), .A2(n1380), .ZN(n1170) );
NAND2_X1 U1102 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
XOR2_X1 U1103 ( .A(n1383), .B(KEYINPUT27), .Z(n1379) );
NAND2_X1 U1104 ( .A1(n1384), .A2(n1385), .ZN(n1383) );
XOR2_X1 U1105 ( .A(KEYINPUT6), .B(n1381), .Z(n1385) );
XNOR2_X1 U1106 ( .A(n1386), .B(n1387), .ZN(n1381) );
XOR2_X1 U1107 ( .A(G107), .B(n1388), .Z(n1387) );
NOR2_X1 U1108 ( .A1(G134), .A2(KEYINPUT8), .ZN(n1388) );
XNOR2_X1 U1109 ( .A(n1319), .B(n1345), .ZN(n1386) );
XOR2_X1 U1110 ( .A(G143), .B(G128), .Z(n1345) );
XNOR2_X1 U1111 ( .A(n1368), .B(n1361), .ZN(n1319) );
INV_X1 U1112 ( .A(n1355), .ZN(n1361) );
XNOR2_X1 U1113 ( .A(G116), .B(KEYINPUT45), .ZN(n1355) );
INV_X1 U1114 ( .A(G122), .ZN(n1368) );
INV_X1 U1115 ( .A(n1382), .ZN(n1384) );
NAND3_X1 U1116 ( .A1(G217), .A2(n1178), .A3(G234), .ZN(n1382) );
XOR2_X1 U1117 ( .A(n1389), .B(n1124), .Z(n1287) );
NOR2_X1 U1118 ( .A1(n1166), .A2(G902), .ZN(n1124) );
XNOR2_X1 U1119 ( .A(n1390), .B(n1391), .ZN(n1166) );
XOR2_X1 U1120 ( .A(G137), .B(n1392), .Z(n1391) );
AND3_X1 U1121 ( .A1(G221), .A2(n1178), .A3(G234), .ZN(n1392) );
INV_X1 U1122 ( .A(G953), .ZN(n1178) );
NAND2_X1 U1123 ( .A1(n1393), .A2(n1394), .ZN(n1390) );
NAND2_X1 U1124 ( .A1(n1395), .A2(n1396), .ZN(n1394) );
XOR2_X1 U1125 ( .A(G128), .B(n1320), .Z(n1396) );
XOR2_X1 U1126 ( .A(n1270), .B(n1142), .Z(n1395) );
INV_X1 U1127 ( .A(G146), .ZN(n1270) );
XOR2_X1 U1128 ( .A(n1397), .B(KEYINPUT35), .Z(n1393) );
NAND2_X1 U1129 ( .A1(n1398), .A2(n1399), .ZN(n1397) );
XOR2_X1 U1130 ( .A(G146), .B(n1142), .Z(n1399) );
XOR2_X1 U1131 ( .A(G140), .B(G125), .Z(n1142) );
XNOR2_X1 U1132 ( .A(G128), .B(n1320), .ZN(n1398) );
XNOR2_X1 U1133 ( .A(G110), .B(n1297), .ZN(n1320) );
INV_X1 U1134 ( .A(G119), .ZN(n1297) );
NAND2_X1 U1135 ( .A1(KEYINPUT60), .A2(n1127), .ZN(n1389) );
NAND2_X1 U1136 ( .A1(G217), .A2(n1400), .ZN(n1127) );
XOR2_X1 U1137 ( .A(KEYINPUT63), .B(n1401), .Z(n1400) );
AND2_X1 U1138 ( .A1(n1312), .A2(G234), .ZN(n1401) );
INV_X1 U1139 ( .A(G902), .ZN(n1312) );
endmodule


