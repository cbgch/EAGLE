//Key = 0100011001101001011110011101010110110101000011011100111001000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401;

NAND2_X1 U756 ( .A1(n1050), .A2(n1051), .ZN(G9) );
NAND2_X1 U757 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XNOR2_X1 U758 ( .A(n1054), .B(KEYINPUT35), .ZN(n1052) );
NAND2_X1 U759 ( .A1(G107), .A2(n1055), .ZN(n1050) );
XNOR2_X1 U760 ( .A(n1054), .B(KEYINPUT4), .ZN(n1055) );
NOR2_X1 U761 ( .A1(n1056), .A2(n1057), .ZN(G75) );
NOR4_X1 U762 ( .A1(G953), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1057) );
NOR2_X1 U763 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR2_X1 U764 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR3_X1 U765 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NOR2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR3_X1 U768 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1068) );
NOR3_X1 U769 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1074) );
NOR2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1073) );
NOR3_X1 U771 ( .A1(n1080), .A2(n1081), .A3(n1071), .ZN(n1063) );
INV_X1 U772 ( .A(n1078), .ZN(n1071) );
NOR3_X1 U773 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NOR2_X1 U774 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XNOR2_X1 U775 ( .A(KEYINPUT25), .B(n1065), .ZN(n1086) );
NOR3_X1 U776 ( .A1(n1087), .A2(n1088), .A3(n1065), .ZN(n1083) );
NOR2_X1 U777 ( .A1(n1089), .A2(n1067), .ZN(n1082) );
NOR2_X1 U778 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XNOR2_X1 U779 ( .A(n1092), .B(KEYINPUT27), .ZN(n1091) );
NOR3_X1 U780 ( .A1(n1058), .A2(G953), .A3(G952), .ZN(n1056) );
AND4_X1 U781 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1058) );
NOR4_X1 U782 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
XOR2_X1 U783 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U784 ( .A1(G472), .A2(KEYINPUT13), .ZN(n1102) );
XOR2_X1 U785 ( .A(n1103), .B(n1104), .Z(n1099) );
XNOR2_X1 U786 ( .A(KEYINPUT52), .B(n1105), .ZN(n1104) );
INV_X1 U787 ( .A(G469), .ZN(n1105) );
XNOR2_X1 U788 ( .A(n1106), .B(KEYINPUT1), .ZN(n1098) );
XNOR2_X1 U789 ( .A(G478), .B(n1107), .ZN(n1095) );
XOR2_X1 U790 ( .A(n1108), .B(n1109), .Z(G72) );
XOR2_X1 U791 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XOR2_X1 U793 ( .A(n1114), .B(n1115), .Z(n1113) );
XNOR2_X1 U794 ( .A(n1116), .B(n1117), .ZN(n1115) );
XOR2_X1 U795 ( .A(n1118), .B(n1119), .Z(n1114) );
XNOR2_X1 U796 ( .A(G131), .B(KEYINPUT63), .ZN(n1119) );
NAND2_X1 U797 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
NAND2_X1 U798 ( .A1(G134), .A2(n1122), .ZN(n1121) );
XOR2_X1 U799 ( .A(KEYINPUT24), .B(n1123), .Z(n1120) );
NOR2_X1 U800 ( .A1(G134), .A2(n1122), .ZN(n1123) );
NOR2_X1 U801 ( .A1(G900), .A2(n1124), .ZN(n1112) );
NOR2_X1 U802 ( .A1(n1125), .A2(G953), .ZN(n1110) );
NOR2_X1 U803 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XNOR2_X1 U804 ( .A(KEYINPUT41), .B(n1128), .ZN(n1127) );
NOR2_X1 U805 ( .A1(n1129), .A2(n1130), .ZN(n1108) );
AND2_X1 U806 ( .A1(G227), .A2(G900), .ZN(n1129) );
XOR2_X1 U807 ( .A(n1131), .B(n1132), .Z(G69) );
XOR2_X1 U808 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U809 ( .A1(n1135), .A2(G953), .ZN(n1134) );
NOR3_X1 U810 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1133) );
NOR2_X1 U811 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U812 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U813 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
INV_X1 U814 ( .A(KEYINPUT8), .ZN(n1139) );
NOR2_X1 U815 ( .A1(KEYINPUT8), .A2(n1145), .ZN(n1137) );
NOR2_X1 U816 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NOR2_X1 U817 ( .A1(n1142), .A2(n1144), .ZN(n1146) );
NOR2_X1 U818 ( .A1(G898), .A2(n1124), .ZN(n1136) );
NOR2_X1 U819 ( .A1(n1148), .A2(n1130), .ZN(n1131) );
NOR2_X1 U820 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U821 ( .A1(n1151), .A2(n1152), .ZN(G66) );
XNOR2_X1 U822 ( .A(n1153), .B(n1154), .ZN(n1152) );
NOR2_X1 U823 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U824 ( .A1(n1151), .A2(n1157), .ZN(G63) );
NOR3_X1 U825 ( .A1(n1107), .A2(n1158), .A3(n1159), .ZN(n1157) );
NOR3_X1 U826 ( .A1(n1160), .A2(n1161), .A3(n1156), .ZN(n1159) );
NOR2_X1 U827 ( .A1(n1162), .A2(n1163), .ZN(n1158) );
AND2_X1 U828 ( .A1(n1060), .A2(G478), .ZN(n1162) );
NOR3_X1 U829 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(G60) );
AND3_X1 U830 ( .A1(KEYINPUT59), .A2(G953), .A3(G952), .ZN(n1166) );
NOR2_X1 U831 ( .A1(KEYINPUT59), .A2(n1167), .ZN(n1165) );
INV_X1 U832 ( .A(n1151), .ZN(n1167) );
XOR2_X1 U833 ( .A(n1168), .B(n1169), .Z(n1164) );
NOR2_X1 U834 ( .A1(n1170), .A2(n1156), .ZN(n1169) );
NAND2_X1 U835 ( .A1(KEYINPUT23), .A2(n1171), .ZN(n1168) );
XOR2_X1 U836 ( .A(G104), .B(n1172), .Z(G6) );
NOR2_X1 U837 ( .A1(n1173), .A2(n1174), .ZN(G57) );
XOR2_X1 U838 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U839 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR2_X1 U840 ( .A1(KEYINPUT56), .A2(n1179), .ZN(n1175) );
XOR2_X1 U841 ( .A(n1180), .B(n1181), .Z(n1179) );
XNOR2_X1 U842 ( .A(n1182), .B(n1183), .ZN(n1181) );
XNOR2_X1 U843 ( .A(n1184), .B(n1185), .ZN(n1180) );
NOR2_X1 U844 ( .A1(n1186), .A2(n1156), .ZN(n1185) );
NOR2_X1 U845 ( .A1(G952), .A2(n1187), .ZN(n1173) );
XNOR2_X1 U846 ( .A(KEYINPUT12), .B(n1130), .ZN(n1187) );
NOR2_X1 U847 ( .A1(n1151), .A2(n1188), .ZN(G54) );
XOR2_X1 U848 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U849 ( .A(n1191), .B(n1192), .Z(n1189) );
NOR2_X1 U850 ( .A1(n1193), .A2(n1156), .ZN(n1192) );
XNOR2_X1 U851 ( .A(G469), .B(KEYINPUT3), .ZN(n1193) );
NAND3_X1 U852 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1191) );
NAND2_X1 U853 ( .A1(n1197), .A2(KEYINPUT40), .ZN(n1196) );
NAND3_X1 U854 ( .A1(n1198), .A2(n1199), .A3(n1116), .ZN(n1195) );
INV_X1 U855 ( .A(KEYINPUT40), .ZN(n1199) );
OR2_X1 U856 ( .A1(n1116), .A2(n1198), .ZN(n1194) );
NOR2_X1 U857 ( .A1(KEYINPUT51), .A2(n1197), .ZN(n1198) );
XNOR2_X1 U858 ( .A(n1200), .B(KEYINPUT34), .ZN(n1197) );
NOR2_X1 U859 ( .A1(n1151), .A2(n1201), .ZN(G51) );
XOR2_X1 U860 ( .A(n1202), .B(n1203), .Z(n1201) );
XNOR2_X1 U861 ( .A(n1204), .B(n1205), .ZN(n1203) );
NOR3_X1 U862 ( .A1(n1156), .A2(KEYINPUT22), .A3(n1206), .ZN(n1205) );
NAND2_X1 U863 ( .A1(G902), .A2(n1060), .ZN(n1156) );
NAND3_X1 U864 ( .A1(n1135), .A2(n1128), .A3(n1207), .ZN(n1060) );
INV_X1 U865 ( .A(n1126), .ZN(n1207) );
NAND4_X1 U866 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1126) );
NOR4_X1 U867 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1211) );
INV_X1 U868 ( .A(n1216), .ZN(n1213) );
INV_X1 U869 ( .A(n1217), .ZN(n1212) );
AND2_X1 U870 ( .A1(n1218), .A2(n1219), .ZN(n1135) );
NOR4_X1 U871 ( .A1(n1172), .A2(n1220), .A3(n1054), .A4(n1221), .ZN(n1219) );
AND3_X1 U872 ( .A1(n1078), .A2(n1222), .A3(n1090), .ZN(n1054) );
NOR3_X1 U873 ( .A1(n1065), .A2(n1223), .A3(n1224), .ZN(n1220) );
AND3_X1 U874 ( .A1(n1078), .A2(n1222), .A3(n1092), .ZN(n1172) );
NOR4_X1 U875 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1218) );
NOR2_X1 U876 ( .A1(n1070), .A2(n1229), .ZN(n1228) );
XOR2_X1 U877 ( .A(n1230), .B(KEYINPUT44), .Z(n1202) );
NOR2_X1 U878 ( .A1(n1130), .A2(G952), .ZN(n1151) );
NAND2_X1 U879 ( .A1(n1231), .A2(n1232), .ZN(G48) );
OR2_X1 U880 ( .A1(n1208), .A2(G146), .ZN(n1232) );
XOR2_X1 U881 ( .A(n1233), .B(KEYINPUT58), .Z(n1231) );
NAND2_X1 U882 ( .A1(G146), .A2(n1208), .ZN(n1233) );
NAND3_X1 U883 ( .A1(n1234), .A2(n1092), .A3(n1235), .ZN(n1208) );
XNOR2_X1 U884 ( .A(G143), .B(n1209), .ZN(G45) );
NAND4_X1 U885 ( .A1(n1235), .A2(n1077), .A3(n1236), .A4(n1237), .ZN(n1209) );
XNOR2_X1 U886 ( .A(n1238), .B(n1215), .ZN(G42) );
AND3_X1 U887 ( .A1(n1076), .A2(n1092), .A3(n1239), .ZN(n1215) );
XOR2_X1 U888 ( .A(n1214), .B(n1240), .Z(G39) );
NOR2_X1 U889 ( .A1(KEYINPUT21), .A2(n1122), .ZN(n1240) );
INV_X1 U890 ( .A(G137), .ZN(n1122) );
AND3_X1 U891 ( .A1(n1234), .A2(n1239), .A3(n1241), .ZN(n1214) );
XNOR2_X1 U892 ( .A(G134), .B(n1128), .ZN(G36) );
NAND3_X1 U893 ( .A1(n1239), .A2(n1090), .A3(n1077), .ZN(n1128) );
XNOR2_X1 U894 ( .A(G131), .B(n1216), .ZN(G33) );
NAND3_X1 U895 ( .A1(n1239), .A2(n1092), .A3(n1077), .ZN(n1216) );
NOR3_X1 U896 ( .A1(n1085), .A2(n1242), .A3(n1080), .ZN(n1239) );
INV_X1 U897 ( .A(n1094), .ZN(n1080) );
NOR2_X1 U898 ( .A1(n1072), .A2(n1075), .ZN(n1094) );
XOR2_X1 U899 ( .A(n1243), .B(n1244), .Z(G30) );
XNOR2_X1 U900 ( .A(KEYINPUT26), .B(n1245), .ZN(n1244) );
NAND2_X1 U901 ( .A1(n1246), .A2(n1247), .ZN(n1243) );
OR2_X1 U902 ( .A1(n1210), .A2(KEYINPUT38), .ZN(n1247) );
NAND3_X1 U903 ( .A1(n1234), .A2(n1090), .A3(n1235), .ZN(n1210) );
AND2_X1 U904 ( .A1(n1248), .A2(n1249), .ZN(n1235) );
NAND4_X1 U905 ( .A1(n1090), .A2(n1248), .A3(n1250), .A4(KEYINPUT38), .ZN(n1246) );
NOR2_X1 U906 ( .A1(n1251), .A2(n1249), .ZN(n1250) );
XOR2_X1 U907 ( .A(G101), .B(n1227), .Z(G3) );
AND3_X1 U908 ( .A1(n1077), .A2(n1222), .A3(n1241), .ZN(n1227) );
INV_X1 U909 ( .A(n1223), .ZN(n1222) );
NAND2_X1 U910 ( .A1(n1248), .A2(n1252), .ZN(n1223) );
NOR2_X1 U911 ( .A1(n1070), .A2(n1085), .ZN(n1248) );
XNOR2_X1 U912 ( .A(G125), .B(n1217), .ZN(G27) );
NAND4_X1 U913 ( .A1(n1076), .A2(n1253), .A3(n1254), .A4(n1092), .ZN(n1217) );
NOR2_X1 U914 ( .A1(n1242), .A2(n1070), .ZN(n1254) );
INV_X1 U915 ( .A(n1249), .ZN(n1242) );
NAND2_X1 U916 ( .A1(n1255), .A2(n1062), .ZN(n1249) );
NAND2_X1 U917 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
INV_X1 U918 ( .A(G900), .ZN(n1257) );
XNOR2_X1 U919 ( .A(G122), .B(n1258), .ZN(G24) );
NAND2_X1 U920 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
XOR2_X1 U921 ( .A(n1229), .B(KEYINPUT29), .Z(n1259) );
NAND3_X1 U922 ( .A1(n1253), .A2(n1078), .A3(n1261), .ZN(n1229) );
NOR3_X1 U923 ( .A1(n1262), .A2(n1263), .A3(n1093), .ZN(n1261) );
NOR2_X1 U924 ( .A1(n1264), .A2(n1106), .ZN(n1078) );
XNOR2_X1 U925 ( .A(n1226), .B(n1265), .ZN(G21) );
NAND2_X1 U926 ( .A1(KEYINPUT18), .A2(G119), .ZN(n1265) );
AND3_X1 U927 ( .A1(n1241), .A2(n1234), .A3(n1266), .ZN(n1226) );
INV_X1 U928 ( .A(n1251), .ZN(n1234) );
NAND2_X1 U929 ( .A1(n1106), .A2(n1264), .ZN(n1251) );
INV_X1 U930 ( .A(n1065), .ZN(n1241) );
XOR2_X1 U931 ( .A(G116), .B(n1225), .Z(G18) );
AND3_X1 U932 ( .A1(n1077), .A2(n1090), .A3(n1266), .ZN(n1225) );
NOR2_X1 U933 ( .A1(n1237), .A2(n1262), .ZN(n1090) );
XNOR2_X1 U934 ( .A(n1267), .B(n1221), .ZN(G15) );
AND3_X1 U935 ( .A1(n1077), .A2(n1092), .A3(n1266), .ZN(n1221) );
NOR3_X1 U936 ( .A1(n1070), .A2(n1263), .A3(n1067), .ZN(n1266) );
INV_X1 U937 ( .A(n1253), .ZN(n1067) );
NOR2_X1 U938 ( .A1(n1088), .A2(n1097), .ZN(n1253) );
INV_X1 U939 ( .A(n1087), .ZN(n1097) );
INV_X1 U940 ( .A(n1252), .ZN(n1263) );
NOR2_X1 U941 ( .A1(n1236), .A2(n1093), .ZN(n1092) );
INV_X1 U942 ( .A(n1262), .ZN(n1236) );
AND2_X1 U943 ( .A1(n1268), .A2(n1264), .ZN(n1077) );
XNOR2_X1 U944 ( .A(G110), .B(n1269), .ZN(G12) );
NAND4_X1 U945 ( .A1(n1270), .A2(n1252), .A3(n1271), .A4(n1272), .ZN(n1269) );
NOR2_X1 U946 ( .A1(n1224), .A2(n1065), .ZN(n1272) );
NAND2_X1 U947 ( .A1(n1273), .A2(n1262), .ZN(n1065) );
XNOR2_X1 U948 ( .A(n1274), .B(n1107), .ZN(n1262) );
NOR2_X1 U949 ( .A1(n1163), .A2(G902), .ZN(n1107) );
INV_X1 U950 ( .A(n1160), .ZN(n1163) );
XNOR2_X1 U951 ( .A(n1275), .B(n1276), .ZN(n1160) );
XOR2_X1 U952 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U953 ( .A(n1053), .B(n1279), .ZN(n1278) );
AND3_X1 U954 ( .A1(G234), .A2(n1130), .A3(G217), .ZN(n1279) );
INV_X1 U955 ( .A(G107), .ZN(n1053) );
XOR2_X1 U956 ( .A(n1280), .B(n1281), .Z(n1275) );
XNOR2_X1 U957 ( .A(n1282), .B(G134), .ZN(n1281) );
XNOR2_X1 U958 ( .A(G116), .B(G128), .ZN(n1280) );
NAND2_X1 U959 ( .A1(KEYINPUT6), .A2(n1161), .ZN(n1274) );
INV_X1 U960 ( .A(G478), .ZN(n1161) );
XNOR2_X1 U961 ( .A(KEYINPUT39), .B(n1093), .ZN(n1273) );
INV_X1 U962 ( .A(n1237), .ZN(n1093) );
XOR2_X1 U963 ( .A(n1283), .B(n1170), .Z(n1237) );
INV_X1 U964 ( .A(G475), .ZN(n1170) );
NAND2_X1 U965 ( .A1(n1171), .A2(n1284), .ZN(n1283) );
XNOR2_X1 U966 ( .A(n1285), .B(n1286), .ZN(n1171) );
XNOR2_X1 U967 ( .A(n1287), .B(n1288), .ZN(n1286) );
XOR2_X1 U968 ( .A(n1289), .B(n1290), .Z(n1288) );
NOR2_X1 U969 ( .A1(KEYINPUT11), .A2(n1277), .ZN(n1290) );
NAND3_X1 U970 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n1289) );
OR2_X1 U971 ( .A1(G140), .A2(KEYINPUT15), .ZN(n1293) );
NAND3_X1 U972 ( .A1(KEYINPUT15), .A2(G140), .A3(n1294), .ZN(n1292) );
NAND2_X1 U973 ( .A1(G125), .A2(n1295), .ZN(n1291) );
NAND2_X1 U974 ( .A1(n1296), .A2(KEYINPUT15), .ZN(n1295) );
XNOR2_X1 U975 ( .A(G140), .B(KEYINPUT19), .ZN(n1296) );
XOR2_X1 U976 ( .A(n1297), .B(n1298), .Z(n1285) );
XNOR2_X1 U977 ( .A(G146), .B(n1299), .ZN(n1298) );
XNOR2_X1 U978 ( .A(G113), .B(n1300), .ZN(n1297) );
NOR2_X1 U979 ( .A1(KEYINPUT60), .A2(n1301), .ZN(n1300) );
XNOR2_X1 U980 ( .A(n1282), .B(n1302), .ZN(n1301) );
NOR2_X1 U981 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
INV_X1 U982 ( .A(G214), .ZN(n1304) );
INV_X1 U983 ( .A(G143), .ZN(n1282) );
INV_X1 U984 ( .A(n1076), .ZN(n1224) );
NOR2_X1 U985 ( .A1(n1264), .A2(n1268), .ZN(n1076) );
INV_X1 U986 ( .A(n1106), .ZN(n1268) );
XOR2_X1 U987 ( .A(n1305), .B(n1155), .Z(n1106) );
NAND2_X1 U988 ( .A1(G217), .A2(n1306), .ZN(n1155) );
NAND2_X1 U989 ( .A1(n1153), .A2(n1284), .ZN(n1305) );
XNOR2_X1 U990 ( .A(n1307), .B(n1308), .ZN(n1153) );
NOR2_X1 U991 ( .A1(G137), .A2(KEYINPUT28), .ZN(n1308) );
XOR2_X1 U992 ( .A(n1309), .B(n1310), .Z(n1307) );
AND3_X1 U993 ( .A1(G221), .A2(n1130), .A3(G234), .ZN(n1310) );
NAND2_X1 U994 ( .A1(n1311), .A2(n1312), .ZN(n1309) );
NAND2_X1 U995 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U996 ( .A(G146), .B(n1117), .Z(n1314) );
XNOR2_X1 U997 ( .A(n1315), .B(n1316), .ZN(n1313) );
XOR2_X1 U998 ( .A(n1317), .B(KEYINPUT42), .Z(n1311) );
NAND2_X1 U999 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
XNOR2_X1 U1000 ( .A(G110), .B(n1315), .ZN(n1319) );
NAND2_X1 U1001 ( .A1(n1320), .A2(n1321), .ZN(n1315) );
NAND2_X1 U1002 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NAND2_X1 U1003 ( .A1(n1324), .A2(n1325), .ZN(n1322) );
NAND2_X1 U1004 ( .A1(n1245), .A2(n1326), .ZN(n1325) );
NAND2_X1 U1005 ( .A1(G128), .A2(n1327), .ZN(n1320) );
NAND2_X1 U1006 ( .A1(n1326), .A2(n1328), .ZN(n1327) );
NAND2_X1 U1007 ( .A1(G119), .A2(n1324), .ZN(n1328) );
INV_X1 U1008 ( .A(KEYINPUT2), .ZN(n1324) );
INV_X1 U1009 ( .A(KEYINPUT16), .ZN(n1326) );
XNOR2_X1 U1010 ( .A(G146), .B(n1117), .ZN(n1318) );
XNOR2_X1 U1011 ( .A(n1294), .B(G140), .ZN(n1117) );
XOR2_X1 U1012 ( .A(n1101), .B(n1186), .Z(n1264) );
INV_X1 U1013 ( .A(G472), .ZN(n1186) );
NAND2_X1 U1014 ( .A1(n1329), .A2(n1284), .ZN(n1101) );
XOR2_X1 U1015 ( .A(n1330), .B(n1331), .Z(n1329) );
NOR2_X1 U1016 ( .A1(n1178), .A2(n1332), .ZN(n1331) );
XOR2_X1 U1017 ( .A(KEYINPUT55), .B(n1177), .Z(n1332) );
AND2_X1 U1018 ( .A1(n1333), .A2(n1334), .ZN(n1177) );
OR2_X1 U1019 ( .A1(n1206), .A2(n1303), .ZN(n1334) );
NOR3_X1 U1020 ( .A1(n1333), .A2(n1303), .A3(n1206), .ZN(n1178) );
INV_X1 U1021 ( .A(G210), .ZN(n1206) );
NAND2_X1 U1022 ( .A1(n1335), .A2(n1130), .ZN(n1303) );
XNOR2_X1 U1023 ( .A(G237), .B(KEYINPUT36), .ZN(n1335) );
NAND2_X1 U1024 ( .A1(KEYINPUT31), .A2(n1336), .ZN(n1330) );
NAND2_X1 U1025 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
OR2_X1 U1026 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
XOR2_X1 U1027 ( .A(n1341), .B(KEYINPUT46), .Z(n1337) );
NAND2_X1 U1028 ( .A1(n1340), .A2(n1339), .ZN(n1341) );
XOR2_X1 U1029 ( .A(n1342), .B(n1343), .Z(n1339) );
INV_X1 U1030 ( .A(n1182), .ZN(n1343) );
XNOR2_X1 U1031 ( .A(n1344), .B(KEYINPUT9), .ZN(n1182) );
NAND2_X1 U1032 ( .A1(KEYINPUT54), .A2(n1345), .ZN(n1342) );
INV_X1 U1033 ( .A(n1085), .ZN(n1271) );
NAND2_X1 U1034 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NAND3_X1 U1035 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1088) );
OR2_X1 U1036 ( .A1(n1103), .A2(G469), .ZN(n1348) );
NAND2_X1 U1037 ( .A1(n1349), .A2(n1350), .ZN(n1347) );
INV_X1 U1038 ( .A(KEYINPUT57), .ZN(n1350) );
NAND2_X1 U1039 ( .A1(n1351), .A2(n1103), .ZN(n1349) );
XNOR2_X1 U1040 ( .A(KEYINPUT61), .B(G469), .ZN(n1351) );
NAND2_X1 U1041 ( .A1(KEYINPUT57), .A2(n1352), .ZN(n1346) );
NAND2_X1 U1042 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
OR2_X1 U1043 ( .A1(G469), .A2(KEYINPUT61), .ZN(n1354) );
NAND3_X1 U1044 ( .A1(G469), .A2(n1103), .A3(KEYINPUT61), .ZN(n1353) );
NAND2_X1 U1045 ( .A1(n1355), .A2(n1284), .ZN(n1103) );
XNOR2_X1 U1046 ( .A(n1116), .B(n1356), .ZN(n1355) );
XNOR2_X1 U1047 ( .A(n1190), .B(n1357), .ZN(n1356) );
XNOR2_X1 U1048 ( .A(n1358), .B(n1359), .ZN(n1190) );
XNOR2_X1 U1049 ( .A(n1316), .B(n1360), .ZN(n1359) );
XNOR2_X1 U1050 ( .A(KEYINPUT37), .B(n1238), .ZN(n1360) );
INV_X1 U1051 ( .A(G140), .ZN(n1238) );
INV_X1 U1052 ( .A(G110), .ZN(n1316) );
XNOR2_X1 U1053 ( .A(n1361), .B(n1345), .ZN(n1358) );
INV_X1 U1054 ( .A(n1184), .ZN(n1345) );
XNOR2_X1 U1055 ( .A(n1362), .B(n1363), .ZN(n1184) );
XNOR2_X1 U1056 ( .A(G137), .B(n1364), .ZN(n1363) );
NAND2_X1 U1057 ( .A1(KEYINPUT45), .A2(n1365), .ZN(n1364) );
INV_X1 U1058 ( .A(G134), .ZN(n1365) );
NAND2_X1 U1059 ( .A1(KEYINPUT10), .A2(n1299), .ZN(n1362) );
INV_X1 U1060 ( .A(G131), .ZN(n1299) );
NAND2_X1 U1061 ( .A1(G227), .A2(n1130), .ZN(n1361) );
XNOR2_X1 U1062 ( .A(n1366), .B(n1367), .ZN(n1116) );
NOR2_X1 U1063 ( .A1(G128), .A2(KEYINPUT30), .ZN(n1367) );
NAND2_X1 U1064 ( .A1(G221), .A2(n1306), .ZN(n1087) );
NAND2_X1 U1065 ( .A1(G234), .A2(n1284), .ZN(n1306) );
NAND2_X1 U1066 ( .A1(n1062), .A2(n1368), .ZN(n1252) );
NAND2_X1 U1067 ( .A1(n1256), .A2(n1150), .ZN(n1368) );
INV_X1 U1068 ( .A(G898), .ZN(n1150) );
NOR3_X1 U1069 ( .A1(n1124), .A2(n1369), .A3(n1284), .ZN(n1256) );
INV_X1 U1070 ( .A(G902), .ZN(n1284) );
AND2_X1 U1071 ( .A1(G234), .A2(G237), .ZN(n1369) );
XOR2_X1 U1072 ( .A(G953), .B(KEYINPUT20), .Z(n1124) );
NAND3_X1 U1073 ( .A1(n1370), .A2(n1130), .A3(n1371), .ZN(n1062) );
XOR2_X1 U1074 ( .A(KEYINPUT43), .B(G952), .Z(n1371) );
INV_X1 U1075 ( .A(G953), .ZN(n1130) );
NAND2_X1 U1076 ( .A1(G234), .A2(G237), .ZN(n1370) );
XNOR2_X1 U1077 ( .A(KEYINPUT14), .B(n1070), .ZN(n1270) );
INV_X1 U1078 ( .A(n1260), .ZN(n1070) );
NOR2_X1 U1079 ( .A1(n1372), .A2(n1075), .ZN(n1260) );
INV_X1 U1080 ( .A(n1079), .ZN(n1075) );
NAND2_X1 U1081 ( .A1(G214), .A2(n1373), .ZN(n1079) );
INV_X1 U1082 ( .A(n1072), .ZN(n1372) );
XNOR2_X1 U1083 ( .A(n1374), .B(n1375), .ZN(n1072) );
NOR2_X1 U1084 ( .A1(G902), .A2(n1376), .ZN(n1375) );
XOR2_X1 U1085 ( .A(n1377), .B(n1378), .Z(n1376) );
XOR2_X1 U1086 ( .A(n1230), .B(KEYINPUT49), .Z(n1378) );
NAND3_X1 U1087 ( .A1(n1379), .A2(n1380), .A3(n1381), .ZN(n1230) );
OR2_X1 U1088 ( .A1(n1144), .A2(n1142), .ZN(n1381) );
NAND2_X1 U1089 ( .A1(KEYINPUT62), .A2(n1382), .ZN(n1380) );
XOR2_X1 U1090 ( .A(n1143), .B(n1142), .Z(n1382) );
NAND2_X1 U1091 ( .A1(n1147), .A2(n1383), .ZN(n1379) );
INV_X1 U1092 ( .A(KEYINPUT62), .ZN(n1383) );
NAND2_X1 U1093 ( .A1(n1384), .A2(n1385), .ZN(n1147) );
NAND3_X1 U1094 ( .A1(n1142), .A2(n1144), .A3(n1143), .ZN(n1385) );
NAND3_X1 U1095 ( .A1(n1386), .A2(n1387), .A3(n1200), .ZN(n1144) );
NAND2_X1 U1096 ( .A1(KEYINPUT33), .A2(n1388), .ZN(n1387) );
NAND2_X1 U1097 ( .A1(G113), .A2(n1389), .ZN(n1388) );
NAND2_X1 U1098 ( .A1(n1340), .A2(n1390), .ZN(n1386) );
OR2_X1 U1099 ( .A1(n1143), .A2(n1142), .ZN(n1384) );
XNOR2_X1 U1100 ( .A(n1391), .B(n1277), .ZN(n1142) );
XOR2_X1 U1101 ( .A(G122), .B(KEYINPUT7), .Z(n1277) );
XNOR2_X1 U1102 ( .A(G110), .B(KEYINPUT47), .ZN(n1391) );
NAND3_X1 U1103 ( .A1(n1392), .A2(n1393), .A3(n1357), .ZN(n1143) );
INV_X1 U1104 ( .A(n1200), .ZN(n1357) );
XOR2_X1 U1105 ( .A(n1394), .B(n1395), .Z(n1200) );
INV_X1 U1106 ( .A(n1287), .ZN(n1395) );
XOR2_X1 U1107 ( .A(G104), .B(KEYINPUT48), .Z(n1287) );
XNOR2_X1 U1108 ( .A(G107), .B(n1333), .ZN(n1394) );
XOR2_X1 U1109 ( .A(G101), .B(KEYINPUT53), .Z(n1333) );
NAND2_X1 U1110 ( .A1(n1183), .A2(n1390), .ZN(n1393) );
INV_X1 U1111 ( .A(KEYINPUT33), .ZN(n1390) );
INV_X1 U1112 ( .A(n1340), .ZN(n1183) );
XOR2_X1 U1113 ( .A(n1389), .B(n1267), .Z(n1340) );
INV_X1 U1114 ( .A(G113), .ZN(n1267) );
NAND3_X1 U1115 ( .A1(G113), .A2(n1389), .A3(KEYINPUT33), .ZN(n1392) );
XOR2_X1 U1116 ( .A(G116), .B(n1396), .Z(n1389) );
XNOR2_X1 U1117 ( .A(KEYINPUT0), .B(n1323), .ZN(n1396) );
INV_X1 U1118 ( .A(G119), .ZN(n1323) );
NAND2_X1 U1119 ( .A1(KEYINPUT32), .A2(n1204), .ZN(n1377) );
XNOR2_X1 U1120 ( .A(n1397), .B(n1398), .ZN(n1204) );
XNOR2_X1 U1121 ( .A(KEYINPUT50), .B(n1294), .ZN(n1398) );
INV_X1 U1122 ( .A(G125), .ZN(n1294) );
XOR2_X1 U1123 ( .A(n1344), .B(n1399), .Z(n1397) );
NOR2_X1 U1124 ( .A1(n1400), .A2(n1149), .ZN(n1399) );
INV_X1 U1125 ( .A(G224), .ZN(n1149) );
XNOR2_X1 U1126 ( .A(G953), .B(KEYINPUT17), .ZN(n1400) );
XOR2_X1 U1127 ( .A(n1401), .B(n1366), .Z(n1344) );
XOR2_X1 U1128 ( .A(G143), .B(G146), .Z(n1366) );
NAND2_X1 U1129 ( .A1(KEYINPUT5), .A2(n1245), .ZN(n1401) );
INV_X1 U1130 ( .A(G128), .ZN(n1245) );
NAND2_X1 U1131 ( .A1(G210), .A2(n1373), .ZN(n1374) );
OR2_X1 U1132 ( .A1(G902), .A2(G237), .ZN(n1373) );
endmodule


