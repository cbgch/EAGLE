//Key = 1101101001101001000001010100101001000010111101011010101010011101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414, n1415, n1416;

XNOR2_X1 U782 ( .A(G107), .B(n1091), .ZN(G9) );
NOR2_X1 U783 ( .A1(n1092), .A2(n1093), .ZN(G75) );
NOR3_X1 U784 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
INV_X1 U785 ( .A(n1097), .ZN(n1096) );
NOR2_X1 U786 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
NOR3_X1 U787 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1098) );
AND2_X1 U788 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR3_X1 U789 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1101) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NOR2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NOR2_X1 U793 ( .A1(n1114), .A2(n1115), .ZN(n1108) );
NOR2_X1 U794 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NOR2_X1 U795 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
XOR2_X1 U796 ( .A(n1120), .B(KEYINPUT59), .Z(n1100) );
NAND2_X1 U797 ( .A1(n1104), .A2(n1121), .ZN(n1120) );
NAND3_X1 U798 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1094) );
NAND3_X1 U799 ( .A1(n1125), .A2(n1126), .A3(n1104), .ZN(n1124) );
NOR3_X1 U800 ( .A1(n1111), .A2(n1115), .A3(n1105), .ZN(n1104) );
NAND2_X1 U801 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U802 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR3_X1 U803 ( .A1(n1131), .A2(G953), .A3(G952), .ZN(n1092) );
INV_X1 U804 ( .A(n1122), .ZN(n1131) );
NAND4_X1 U805 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1122) );
XNOR2_X1 U806 ( .A(KEYINPUT25), .B(n1130), .ZN(n1134) );
XOR2_X1 U807 ( .A(n1136), .B(KEYINPUT12), .Z(n1133) );
NAND4_X1 U808 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1136) );
XOR2_X1 U809 ( .A(KEYINPUT61), .B(n1141), .Z(n1140) );
NOR2_X1 U810 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NOR2_X1 U811 ( .A1(n1144), .A2(n1145), .ZN(n1139) );
XNOR2_X1 U812 ( .A(n1146), .B(n1147), .ZN(n1145) );
XNOR2_X1 U813 ( .A(n1148), .B(KEYINPUT4), .ZN(n1146) );
AND2_X1 U814 ( .A1(n1143), .A2(n1142), .ZN(n1144) );
INV_X1 U815 ( .A(n1149), .ZN(n1138) );
NOR2_X1 U816 ( .A1(n1150), .A2(n1151), .ZN(n1132) );
AND2_X1 U817 ( .A1(n1111), .A2(KEYINPUT41), .ZN(n1151) );
INV_X1 U818 ( .A(n1152), .ZN(n1111) );
NOR2_X1 U819 ( .A1(KEYINPUT41), .A2(n1153), .ZN(n1150) );
NOR3_X1 U820 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1153) );
XOR2_X1 U821 ( .A(n1157), .B(n1158), .Z(G72) );
XOR2_X1 U822 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U823 ( .A1(n1161), .A2(n1123), .ZN(n1160) );
AND2_X1 U824 ( .A1(G227), .A2(G900), .ZN(n1161) );
NAND2_X1 U825 ( .A1(n1162), .A2(n1163), .ZN(n1159) );
NAND2_X1 U826 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XNOR2_X1 U827 ( .A(KEYINPUT19), .B(n1123), .ZN(n1164) );
XOR2_X1 U828 ( .A(n1166), .B(n1167), .Z(n1162) );
XNOR2_X1 U829 ( .A(n1168), .B(n1169), .ZN(n1167) );
XNOR2_X1 U830 ( .A(KEYINPUT3), .B(n1170), .ZN(n1169) );
NOR2_X1 U831 ( .A1(G131), .A2(KEYINPUT26), .ZN(n1170) );
XNOR2_X1 U832 ( .A(n1171), .B(n1172), .ZN(n1166) );
NAND2_X1 U833 ( .A1(n1123), .A2(n1173), .ZN(n1157) );
NAND2_X1 U834 ( .A1(n1174), .A2(n1175), .ZN(G69) );
NAND2_X1 U835 ( .A1(n1176), .A2(n1123), .ZN(n1175) );
XNOR2_X1 U836 ( .A(n1177), .B(n1178), .ZN(n1176) );
NAND2_X1 U837 ( .A1(n1179), .A2(G953), .ZN(n1174) );
NAND2_X1 U838 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NAND2_X1 U839 ( .A1(n1182), .A2(G224), .ZN(n1181) );
INV_X1 U840 ( .A(n1178), .ZN(n1182) );
NAND2_X1 U841 ( .A1(n1183), .A2(n1178), .ZN(n1180) );
NAND2_X1 U842 ( .A1(n1184), .A2(n1185), .ZN(n1178) );
NAND2_X1 U843 ( .A1(G953), .A2(n1186), .ZN(n1185) );
XNOR2_X1 U844 ( .A(n1187), .B(n1188), .ZN(n1184) );
NAND2_X1 U845 ( .A1(G898), .A2(G224), .ZN(n1183) );
NOR2_X1 U846 ( .A1(n1189), .A2(n1190), .ZN(G66) );
NOR3_X1 U847 ( .A1(n1191), .A2(n1148), .A3(n1192), .ZN(n1190) );
NOR2_X1 U848 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NOR2_X1 U849 ( .A1(n1097), .A2(n1147), .ZN(n1193) );
XOR2_X1 U850 ( .A(KEYINPUT55), .B(n1195), .Z(n1191) );
NOR3_X1 U851 ( .A1(n1196), .A2(n1147), .A3(n1197), .ZN(n1195) );
NOR2_X1 U852 ( .A1(n1189), .A2(n1198), .ZN(G63) );
XOR2_X1 U853 ( .A(n1199), .B(n1200), .Z(n1198) );
NAND3_X1 U854 ( .A1(n1201), .A2(n1202), .A3(G478), .ZN(n1199) );
OR2_X1 U855 ( .A1(n1203), .A2(KEYINPUT29), .ZN(n1202) );
NAND2_X1 U856 ( .A1(KEYINPUT29), .A2(n1204), .ZN(n1201) );
NAND2_X1 U857 ( .A1(n1097), .A2(G902), .ZN(n1204) );
NOR2_X1 U858 ( .A1(n1189), .A2(n1205), .ZN(G60) );
NOR3_X1 U859 ( .A1(n1142), .A2(n1206), .A3(n1207), .ZN(n1205) );
AND3_X1 U860 ( .A1(n1208), .A2(G475), .A3(n1203), .ZN(n1207) );
NOR2_X1 U861 ( .A1(n1209), .A2(n1208), .ZN(n1206) );
NOR2_X1 U862 ( .A1(n1097), .A2(n1143), .ZN(n1209) );
XOR2_X1 U863 ( .A(n1210), .B(n1211), .Z(G6) );
XNOR2_X1 U864 ( .A(G104), .B(KEYINPUT7), .ZN(n1211) );
NOR2_X1 U865 ( .A1(n1189), .A2(n1212), .ZN(G57) );
NOR2_X1 U866 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XOR2_X1 U867 ( .A(KEYINPUT44), .B(n1215), .Z(n1214) );
NOR2_X1 U868 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
AND2_X1 U869 ( .A1(n1217), .A2(n1216), .ZN(n1213) );
XNOR2_X1 U870 ( .A(n1218), .B(n1219), .ZN(n1216) );
XNOR2_X1 U871 ( .A(n1220), .B(n1221), .ZN(n1219) );
XOR2_X1 U872 ( .A(n1222), .B(KEYINPUT53), .Z(n1218) );
NAND2_X1 U873 ( .A1(n1203), .A2(G472), .ZN(n1222) );
XOR2_X1 U874 ( .A(G101), .B(n1223), .Z(n1217) );
NOR2_X1 U875 ( .A1(KEYINPUT39), .A2(n1224), .ZN(n1223) );
NOR2_X1 U876 ( .A1(n1189), .A2(n1225), .ZN(G54) );
XOR2_X1 U877 ( .A(n1226), .B(n1227), .Z(n1225) );
NOR2_X1 U878 ( .A1(n1154), .A2(n1196), .ZN(n1227) );
INV_X1 U879 ( .A(n1203), .ZN(n1196) );
NAND2_X1 U880 ( .A1(n1228), .A2(KEYINPUT50), .ZN(n1226) );
XOR2_X1 U881 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U882 ( .A(n1231), .B(n1232), .Z(n1229) );
NAND2_X1 U883 ( .A1(KEYINPUT21), .A2(n1172), .ZN(n1231) );
NOR2_X1 U884 ( .A1(n1189), .A2(n1233), .ZN(G51) );
XOR2_X1 U885 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U886 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U887 ( .A(n1238), .B(KEYINPUT1), .Z(n1234) );
NAND2_X1 U888 ( .A1(n1203), .A2(n1239), .ZN(n1238) );
NOR2_X1 U889 ( .A1(n1240), .A2(n1097), .ZN(n1203) );
NOR2_X1 U890 ( .A1(n1173), .A2(n1177), .ZN(n1097) );
NAND4_X1 U891 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1177) );
AND4_X1 U892 ( .A1(n1091), .A2(n1245), .A3(n1246), .A4(n1210), .ZN(n1244) );
NAND3_X1 U893 ( .A1(n1247), .A2(n1248), .A3(n1103), .ZN(n1210) );
NAND3_X1 U894 ( .A1(n1248), .A2(n1121), .A3(n1247), .ZN(n1091) );
NAND2_X1 U895 ( .A1(n1249), .A2(n1250), .ZN(n1243) );
NAND2_X1 U896 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U897 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
INV_X1 U898 ( .A(KEYINPUT6), .ZN(n1254) );
NAND4_X1 U899 ( .A1(n1125), .A2(n1117), .A3(n1113), .A4(n1255), .ZN(n1253) );
XNOR2_X1 U900 ( .A(KEYINPUT47), .B(n1256), .ZN(n1251) );
NAND3_X1 U901 ( .A1(n1257), .A2(n1258), .A3(n1152), .ZN(n1242) );
NAND2_X1 U902 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NAND3_X1 U903 ( .A1(n1261), .A2(n1149), .A3(n1248), .ZN(n1260) );
NAND2_X1 U904 ( .A1(n1125), .A2(n1262), .ZN(n1259) );
XOR2_X1 U905 ( .A(KEYINPUT17), .B(n1263), .Z(n1262) );
NAND2_X1 U906 ( .A1(KEYINPUT6), .A2(n1264), .ZN(n1241) );
NAND4_X1 U907 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1173) );
AND4_X1 U908 ( .A1(n1269), .A2(n1270), .A3(n1271), .A4(n1272), .ZN(n1268) );
NOR3_X1 U909 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1267) );
AND4_X1 U910 ( .A1(KEYINPUT27), .A2(n1276), .A3(n1099), .A4(n1103), .ZN(n1275) );
INV_X1 U911 ( .A(n1277), .ZN(n1099) );
NOR2_X1 U912 ( .A1(KEYINPUT27), .A2(n1278), .ZN(n1274) );
NOR2_X1 U913 ( .A1(n1123), .A2(G952), .ZN(n1189) );
XNOR2_X1 U914 ( .A(n1273), .B(n1279), .ZN(G48) );
NAND2_X1 U915 ( .A1(KEYINPUT48), .A2(G146), .ZN(n1279) );
AND2_X1 U916 ( .A1(n1280), .A2(n1103), .ZN(n1273) );
XNOR2_X1 U917 ( .A(G143), .B(n1265), .ZN(G45) );
NAND4_X1 U918 ( .A1(n1276), .A2(n1249), .A3(n1261), .A4(n1149), .ZN(n1265) );
XNOR2_X1 U919 ( .A(G140), .B(n1266), .ZN(G42) );
NAND4_X1 U920 ( .A1(n1103), .A2(n1112), .A3(n1281), .A4(n1277), .ZN(n1266) );
XNOR2_X1 U921 ( .A(G137), .B(n1269), .ZN(G39) );
NAND4_X1 U922 ( .A1(n1263), .A2(n1281), .A3(n1277), .A4(n1125), .ZN(n1269) );
XNOR2_X1 U923 ( .A(G134), .B(n1272), .ZN(G36) );
NAND3_X1 U924 ( .A1(n1277), .A2(n1121), .A3(n1276), .ZN(n1272) );
XNOR2_X1 U925 ( .A(G131), .B(n1278), .ZN(G33) );
NAND3_X1 U926 ( .A1(n1103), .A2(n1277), .A3(n1276), .ZN(n1278) );
AND2_X1 U927 ( .A1(n1281), .A2(n1113), .ZN(n1276) );
NOR2_X1 U928 ( .A1(n1282), .A2(n1129), .ZN(n1277) );
XNOR2_X1 U929 ( .A(n1271), .B(n1283), .ZN(G30) );
NOR2_X1 U930 ( .A1(KEYINPUT34), .A2(n1284), .ZN(n1283) );
NAND2_X1 U931 ( .A1(n1280), .A2(n1121), .ZN(n1271) );
AND3_X1 U932 ( .A1(n1281), .A2(n1249), .A3(n1263), .ZN(n1280) );
AND2_X1 U933 ( .A1(n1117), .A2(n1285), .ZN(n1281) );
NAND2_X1 U934 ( .A1(n1286), .A2(n1287), .ZN(G3) );
NAND2_X1 U935 ( .A1(n1264), .A2(n1288), .ZN(n1287) );
INV_X1 U936 ( .A(n1289), .ZN(n1264) );
XOR2_X1 U937 ( .A(n1290), .B(KEYINPUT13), .Z(n1286) );
NAND2_X1 U938 ( .A1(G101), .A2(n1289), .ZN(n1290) );
NAND3_X1 U939 ( .A1(n1125), .A2(n1113), .A3(n1247), .ZN(n1289) );
XNOR2_X1 U940 ( .A(G125), .B(n1270), .ZN(G27) );
NAND3_X1 U941 ( .A1(n1103), .A2(n1152), .A3(n1291), .ZN(n1270) );
AND3_X1 U942 ( .A1(n1112), .A2(n1285), .A3(n1249), .ZN(n1291) );
NAND2_X1 U943 ( .A1(n1105), .A2(n1292), .ZN(n1285) );
NAND4_X1 U944 ( .A1(G953), .A2(G902), .A3(n1165), .A4(n1293), .ZN(n1292) );
XOR2_X1 U945 ( .A(G900), .B(KEYINPUT40), .Z(n1165) );
XNOR2_X1 U946 ( .A(G122), .B(n1294), .ZN(G24) );
NAND4_X1 U947 ( .A1(n1295), .A2(n1296), .A3(n1152), .A4(n1297), .ZN(n1294) );
AND3_X1 U948 ( .A1(n1248), .A2(n1149), .A3(n1261), .ZN(n1297) );
XOR2_X1 U949 ( .A(n1298), .B(KEYINPUT33), .Z(n1261) );
INV_X1 U950 ( .A(n1115), .ZN(n1248) );
NAND2_X1 U951 ( .A1(n1299), .A2(n1300), .ZN(n1115) );
OR2_X1 U952 ( .A1(n1257), .A2(KEYINPUT16), .ZN(n1296) );
NAND2_X1 U953 ( .A1(KEYINPUT16), .A2(n1301), .ZN(n1295) );
NAND2_X1 U954 ( .A1(n1127), .A2(n1255), .ZN(n1301) );
XNOR2_X1 U955 ( .A(G119), .B(n1302), .ZN(G21) );
NAND4_X1 U956 ( .A1(n1152), .A2(n1125), .A3(n1257), .A4(n1303), .ZN(n1302) );
XOR2_X1 U957 ( .A(KEYINPUT49), .B(n1263), .Z(n1303) );
XOR2_X1 U958 ( .A(G116), .B(n1304), .Z(G18) );
NOR2_X1 U959 ( .A1(n1127), .A2(n1256), .ZN(n1304) );
NAND4_X1 U960 ( .A1(n1152), .A2(n1113), .A3(n1121), .A4(n1255), .ZN(n1256) );
NAND2_X1 U961 ( .A1(n1305), .A2(n1306), .ZN(n1121) );
OR2_X1 U962 ( .A1(n1107), .A2(KEYINPUT63), .ZN(n1306) );
INV_X1 U963 ( .A(n1125), .ZN(n1107) );
NAND3_X1 U964 ( .A1(n1149), .A2(n1298), .A3(KEYINPUT63), .ZN(n1305) );
INV_X1 U965 ( .A(n1249), .ZN(n1127) );
XOR2_X1 U966 ( .A(n1246), .B(n1307), .Z(G15) );
XNOR2_X1 U967 ( .A(G113), .B(KEYINPUT20), .ZN(n1307) );
NAND4_X1 U968 ( .A1(n1103), .A2(n1152), .A3(n1257), .A4(n1113), .ZN(n1246) );
NAND2_X1 U969 ( .A1(n1308), .A2(n1309), .ZN(n1113) );
OR3_X1 U970 ( .A1(n1310), .A2(n1299), .A3(KEYINPUT32), .ZN(n1309) );
NAND2_X1 U971 ( .A1(KEYINPUT32), .A2(n1263), .ZN(n1308) );
NOR2_X1 U972 ( .A1(n1300), .A2(n1299), .ZN(n1263) );
NOR2_X1 U973 ( .A1(n1118), .A2(n1156), .ZN(n1152) );
INV_X1 U974 ( .A(n1119), .ZN(n1156) );
NOR2_X1 U975 ( .A1(n1298), .A2(n1149), .ZN(n1103) );
XNOR2_X1 U976 ( .A(G110), .B(n1245), .ZN(G12) );
NAND3_X1 U977 ( .A1(n1247), .A2(n1125), .A3(n1112), .ZN(n1245) );
AND2_X1 U978 ( .A1(n1310), .A2(n1299), .ZN(n1112) );
NAND2_X1 U979 ( .A1(n1311), .A2(n1312), .ZN(n1299) );
NAND2_X1 U980 ( .A1(KEYINPUT9), .A2(n1137), .ZN(n1312) );
XOR2_X1 U981 ( .A(n1313), .B(G472), .Z(n1137) );
NAND3_X1 U982 ( .A1(G472), .A2(n1313), .A3(n1314), .ZN(n1311) );
INV_X1 U983 ( .A(KEYINPUT9), .ZN(n1314) );
NAND2_X1 U984 ( .A1(n1240), .A2(n1315), .ZN(n1313) );
NAND2_X1 U985 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
NAND2_X1 U986 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
XNOR2_X1 U987 ( .A(n1224), .B(n1288), .ZN(n1319) );
XNOR2_X1 U988 ( .A(n1220), .B(n1320), .ZN(n1318) );
XOR2_X1 U989 ( .A(n1321), .B(KEYINPUT18), .Z(n1316) );
NAND2_X1 U990 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XNOR2_X1 U991 ( .A(G101), .B(n1224), .ZN(n1323) );
NAND3_X1 U992 ( .A1(n1324), .A2(n1123), .A3(G210), .ZN(n1224) );
XNOR2_X1 U993 ( .A(n1320), .B(n1325), .ZN(n1322) );
INV_X1 U994 ( .A(n1220), .ZN(n1325) );
XOR2_X1 U995 ( .A(n1232), .B(n1326), .Z(n1220) );
NOR2_X1 U996 ( .A1(KEYINPUT46), .A2(n1221), .ZN(n1320) );
XOR2_X1 U997 ( .A(n1327), .B(KEYINPUT10), .Z(n1221) );
NAND2_X1 U998 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NAND2_X1 U999 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
XNOR2_X1 U1000 ( .A(KEYINPUT43), .B(n1332), .ZN(n1331) );
XNOR2_X1 U1001 ( .A(n1333), .B(n1334), .ZN(n1330) );
XOR2_X1 U1002 ( .A(n1335), .B(KEYINPUT22), .Z(n1328) );
NAND2_X1 U1003 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XNOR2_X1 U1004 ( .A(G119), .B(n1333), .ZN(n1337) );
NAND2_X1 U1005 ( .A1(KEYINPUT28), .A2(G116), .ZN(n1333) );
XNOR2_X1 U1006 ( .A(KEYINPUT43), .B(G113), .ZN(n1336) );
INV_X1 U1007 ( .A(n1300), .ZN(n1310) );
XOR2_X1 U1008 ( .A(n1338), .B(n1339), .Z(n1300) );
INV_X1 U1009 ( .A(n1148), .ZN(n1339) );
NOR2_X1 U1010 ( .A1(n1194), .A2(G902), .ZN(n1148) );
INV_X1 U1011 ( .A(n1197), .ZN(n1194) );
XNOR2_X1 U1012 ( .A(n1340), .B(n1341), .ZN(n1197) );
XNOR2_X1 U1013 ( .A(n1334), .B(n1342), .ZN(n1341) );
XNOR2_X1 U1014 ( .A(G137), .B(n1284), .ZN(n1342) );
INV_X1 U1015 ( .A(G119), .ZN(n1334) );
XOR2_X1 U1016 ( .A(n1343), .B(n1344), .Z(n1340) );
XNOR2_X1 U1017 ( .A(G110), .B(n1345), .ZN(n1344) );
NAND2_X1 U1018 ( .A1(n1346), .A2(KEYINPUT23), .ZN(n1345) );
XOR2_X1 U1019 ( .A(n1347), .B(G146), .Z(n1346) );
NAND2_X1 U1020 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
OR2_X1 U1021 ( .A1(n1350), .A2(G125), .ZN(n1349) );
XOR2_X1 U1022 ( .A(n1351), .B(KEYINPUT11), .Z(n1348) );
NAND2_X1 U1023 ( .A1(G125), .A2(n1350), .ZN(n1351) );
NAND3_X1 U1024 ( .A1(n1352), .A2(G221), .A3(KEYINPUT42), .ZN(n1343) );
NAND2_X1 U1025 ( .A1(KEYINPUT45), .A2(n1147), .ZN(n1338) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1353), .ZN(n1147) );
NOR2_X1 U1027 ( .A1(n1149), .A2(n1354), .ZN(n1125) );
INV_X1 U1028 ( .A(n1298), .ZN(n1354) );
XOR2_X1 U1029 ( .A(n1142), .B(n1355), .Z(n1298) );
XNOR2_X1 U1030 ( .A(KEYINPUT52), .B(n1143), .ZN(n1355) );
INV_X1 U1031 ( .A(G475), .ZN(n1143) );
NOR2_X1 U1032 ( .A1(n1208), .A2(G902), .ZN(n1142) );
XOR2_X1 U1033 ( .A(n1356), .B(KEYINPUT62), .Z(n1208) );
XOR2_X1 U1034 ( .A(n1357), .B(n1358), .Z(n1356) );
XOR2_X1 U1035 ( .A(n1359), .B(n1360), .Z(n1358) );
XNOR2_X1 U1036 ( .A(G131), .B(n1361), .ZN(n1360) );
XOR2_X1 U1037 ( .A(G146), .B(G143), .Z(n1359) );
XOR2_X1 U1038 ( .A(n1362), .B(n1363), .Z(n1357) );
XNOR2_X1 U1039 ( .A(n1332), .B(G104), .ZN(n1363) );
XOR2_X1 U1040 ( .A(n1364), .B(n1168), .Z(n1362) );
XNOR2_X1 U1041 ( .A(G125), .B(n1350), .ZN(n1168) );
NAND3_X1 U1042 ( .A1(n1324), .A2(n1123), .A3(n1365), .ZN(n1364) );
XOR2_X1 U1043 ( .A(KEYINPUT24), .B(G214), .Z(n1365) );
XNOR2_X1 U1044 ( .A(n1366), .B(G478), .ZN(n1149) );
NAND2_X1 U1045 ( .A1(n1200), .A2(n1367), .ZN(n1366) );
XNOR2_X1 U1046 ( .A(KEYINPUT56), .B(n1240), .ZN(n1367) );
XNOR2_X1 U1047 ( .A(n1368), .B(n1369), .ZN(n1200) );
XOR2_X1 U1048 ( .A(n1370), .B(n1371), .Z(n1369) );
NOR2_X1 U1049 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
NOR2_X1 U1050 ( .A1(KEYINPUT2), .A2(n1374), .ZN(n1373) );
AND2_X1 U1051 ( .A1(KEYINPUT58), .A2(n1374), .ZN(n1372) );
AND2_X1 U1052 ( .A1(n1352), .A2(G217), .ZN(n1370) );
AND2_X1 U1053 ( .A1(G234), .A2(n1123), .ZN(n1352) );
XOR2_X1 U1054 ( .A(n1375), .B(n1376), .Z(n1368) );
NOR2_X1 U1055 ( .A1(KEYINPUT51), .A2(n1377), .ZN(n1376) );
XNOR2_X1 U1056 ( .A(G116), .B(G122), .ZN(n1377) );
XNOR2_X1 U1057 ( .A(G107), .B(G134), .ZN(n1375) );
AND2_X1 U1058 ( .A1(n1117), .A2(n1257), .ZN(n1247) );
AND2_X1 U1059 ( .A1(n1249), .A2(n1255), .ZN(n1257) );
NAND2_X1 U1060 ( .A1(n1105), .A2(n1378), .ZN(n1255) );
NAND4_X1 U1061 ( .A1(G953), .A2(G902), .A3(n1293), .A4(n1186), .ZN(n1378) );
INV_X1 U1062 ( .A(G898), .ZN(n1186) );
NAND3_X1 U1063 ( .A1(n1293), .A2(n1123), .A3(G952), .ZN(n1105) );
NAND2_X1 U1064 ( .A1(G237), .A2(G234), .ZN(n1293) );
NOR2_X1 U1065 ( .A1(n1130), .A2(n1129), .ZN(n1249) );
INV_X1 U1066 ( .A(n1135), .ZN(n1129) );
NAND2_X1 U1067 ( .A1(G214), .A2(n1379), .ZN(n1135) );
INV_X1 U1068 ( .A(n1282), .ZN(n1130) );
XNOR2_X1 U1069 ( .A(n1380), .B(n1239), .ZN(n1282) );
AND2_X1 U1070 ( .A1(G210), .A2(n1379), .ZN(n1239) );
NAND2_X1 U1071 ( .A1(n1324), .A2(n1240), .ZN(n1379) );
INV_X1 U1072 ( .A(G237), .ZN(n1324) );
NAND3_X1 U1073 ( .A1(n1381), .A2(n1240), .A3(n1382), .ZN(n1380) );
XOR2_X1 U1074 ( .A(n1383), .B(KEYINPUT14), .Z(n1382) );
OR2_X1 U1075 ( .A1(n1384), .A2(n1237), .ZN(n1383) );
NAND2_X1 U1076 ( .A1(n1237), .A2(n1384), .ZN(n1381) );
XOR2_X1 U1077 ( .A(n1236), .B(KEYINPUT15), .Z(n1384) );
XNOR2_X1 U1078 ( .A(n1385), .B(n1326), .ZN(n1236) );
XNOR2_X1 U1079 ( .A(n1386), .B(G128), .ZN(n1326) );
NAND2_X1 U1080 ( .A1(KEYINPUT54), .A2(n1387), .ZN(n1386) );
XOR2_X1 U1081 ( .A(G143), .B(n1388), .Z(n1387) );
XOR2_X1 U1082 ( .A(KEYINPUT31), .B(G146), .Z(n1388) );
XNOR2_X1 U1083 ( .A(G125), .B(n1389), .ZN(n1385) );
AND2_X1 U1084 ( .A1(n1123), .A2(G224), .ZN(n1389) );
XOR2_X1 U1085 ( .A(n1390), .B(n1187), .Z(n1237) );
XOR2_X1 U1086 ( .A(n1391), .B(n1392), .Z(n1187) );
XNOR2_X1 U1087 ( .A(n1361), .B(G110), .ZN(n1392) );
INV_X1 U1088 ( .A(G122), .ZN(n1361) );
NAND2_X1 U1089 ( .A1(n1393), .A2(n1394), .ZN(n1391) );
NAND2_X1 U1090 ( .A1(n1395), .A2(n1396), .ZN(n1394) );
NAND2_X1 U1091 ( .A1(n1397), .A2(n1398), .ZN(n1396) );
NAND2_X1 U1092 ( .A1(KEYINPUT60), .A2(G113), .ZN(n1398) );
INV_X1 U1093 ( .A(KEYINPUT36), .ZN(n1397) );
NAND2_X1 U1094 ( .A1(n1399), .A2(n1332), .ZN(n1393) );
INV_X1 U1095 ( .A(G113), .ZN(n1332) );
NAND2_X1 U1096 ( .A1(KEYINPUT60), .A2(n1400), .ZN(n1399) );
OR2_X1 U1097 ( .A1(n1395), .A2(KEYINPUT36), .ZN(n1400) );
XOR2_X1 U1098 ( .A(G116), .B(n1401), .Z(n1395) );
NOR2_X1 U1099 ( .A1(G119), .A2(KEYINPUT35), .ZN(n1401) );
NAND2_X1 U1100 ( .A1(KEYINPUT38), .A2(n1188), .ZN(n1390) );
XOR2_X1 U1101 ( .A(n1402), .B(n1288), .Z(n1188) );
NAND2_X1 U1102 ( .A1(KEYINPUT0), .A2(n1403), .ZN(n1402) );
AND2_X1 U1103 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U1104 ( .A1(G221), .A2(n1353), .ZN(n1119) );
NAND2_X1 U1105 ( .A1(G234), .A2(n1240), .ZN(n1353) );
XNOR2_X1 U1106 ( .A(n1155), .B(n1154), .ZN(n1118) );
INV_X1 U1107 ( .A(G469), .ZN(n1154) );
AND2_X1 U1108 ( .A1(n1404), .A2(n1240), .ZN(n1155) );
INV_X1 U1109 ( .A(G902), .ZN(n1240) );
XOR2_X1 U1110 ( .A(n1230), .B(n1405), .Z(n1404) );
XNOR2_X1 U1111 ( .A(n1406), .B(n1407), .ZN(n1405) );
NOR2_X1 U1112 ( .A1(KEYINPUT57), .A2(n1172), .ZN(n1407) );
XOR2_X1 U1113 ( .A(n1408), .B(n1374), .Z(n1172) );
XNOR2_X1 U1114 ( .A(n1284), .B(G143), .ZN(n1374) );
INV_X1 U1115 ( .A(G128), .ZN(n1284) );
XNOR2_X1 U1116 ( .A(G146), .B(KEYINPUT37), .ZN(n1408) );
NAND2_X1 U1117 ( .A1(KEYINPUT30), .A2(n1232), .ZN(n1406) );
XNOR2_X1 U1118 ( .A(n1171), .B(G131), .ZN(n1232) );
XNOR2_X1 U1119 ( .A(G134), .B(n1409), .ZN(n1171) );
XOR2_X1 U1120 ( .A(KEYINPUT8), .B(G137), .Z(n1409) );
XNOR2_X1 U1121 ( .A(n1410), .B(n1411), .ZN(n1230) );
XNOR2_X1 U1122 ( .A(n1412), .B(n1413), .ZN(n1411) );
XNOR2_X1 U1123 ( .A(KEYINPUT5), .B(n1350), .ZN(n1413) );
INV_X1 U1124 ( .A(G140), .ZN(n1350) );
INV_X1 U1125 ( .A(G110), .ZN(n1412) );
XNOR2_X1 U1126 ( .A(n1403), .B(n1414), .ZN(n1410) );
XNOR2_X1 U1127 ( .A(n1288), .B(n1415), .ZN(n1414) );
AND2_X1 U1128 ( .A1(n1123), .A2(G227), .ZN(n1415) );
INV_X1 U1129 ( .A(G953), .ZN(n1123) );
INV_X1 U1130 ( .A(G101), .ZN(n1288) );
XNOR2_X1 U1131 ( .A(G104), .B(n1416), .ZN(n1403) );
INV_X1 U1132 ( .A(G107), .ZN(n1416) );
endmodule


