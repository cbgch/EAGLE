//Key = 0001011111100010001001011111000011010001000111110011111111010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351;

XOR2_X1 U749 ( .A(G107), .B(n1038), .Z(G9) );
NOR2_X1 U750 ( .A1(n1039), .A2(n1040), .ZN(G75) );
NOR3_X1 U751 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NOR2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U753 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR3_X1 U754 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
NOR2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U756 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR3_X1 U758 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1055) );
NOR2_X1 U759 ( .A1(n1060), .A2(n1061), .ZN(n1051) );
NOR2_X1 U760 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR3_X1 U761 ( .A1(n1061), .A2(n1064), .A3(n1054), .ZN(n1046) );
NOR3_X1 U762 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NOR2_X1 U763 ( .A1(n1068), .A2(n1048), .ZN(n1067) );
NOR2_X1 U764 ( .A1(n1069), .A2(n1050), .ZN(n1065) );
NAND3_X1 U765 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1041) );
NAND4_X1 U766 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1072) );
NOR3_X1 U767 ( .A1(n1077), .A2(n1045), .A3(n1078), .ZN(n1076) );
XOR2_X1 U768 ( .A(KEYINPUT25), .B(n1079), .Z(n1077) );
XNOR2_X1 U769 ( .A(KEYINPUT61), .B(n1080), .ZN(n1074) );
NOR3_X1 U770 ( .A1(n1081), .A2(G953), .A3(G952), .ZN(n1039) );
INV_X1 U771 ( .A(n1070), .ZN(n1081) );
NAND4_X1 U772 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1070) );
AND4_X1 U773 ( .A1(n1057), .A2(n1086), .A3(n1087), .A4(n1080), .ZN(n1085) );
NOR2_X1 U774 ( .A1(n1054), .A2(n1088), .ZN(n1084) );
XOR2_X1 U775 ( .A(n1089), .B(n1090), .Z(n1083) );
XNOR2_X1 U776 ( .A(KEYINPUT44), .B(n1091), .ZN(n1090) );
NOR2_X1 U777 ( .A1(KEYINPUT19), .A2(n1092), .ZN(n1089) );
XOR2_X1 U778 ( .A(n1093), .B(n1094), .Z(n1082) );
XNOR2_X1 U779 ( .A(G475), .B(KEYINPUT56), .ZN(n1094) );
XOR2_X1 U780 ( .A(n1095), .B(n1096), .Z(G72) );
XOR2_X1 U781 ( .A(n1097), .B(n1098), .Z(n1096) );
NAND2_X1 U782 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U783 ( .A1(G953), .A2(n1101), .ZN(n1100) );
XOR2_X1 U784 ( .A(n1102), .B(n1103), .Z(n1099) );
XNOR2_X1 U785 ( .A(n1104), .B(KEYINPUT21), .ZN(n1103) );
NAND2_X1 U786 ( .A1(n1105), .A2(KEYINPUT50), .ZN(n1104) );
XOR2_X1 U787 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U788 ( .A(G137), .B(G134), .Z(n1107) );
XOR2_X1 U789 ( .A(n1108), .B(G131), .Z(n1106) );
NOR2_X1 U790 ( .A1(n1109), .A2(n1110), .ZN(n1102) );
XOR2_X1 U791 ( .A(n1111), .B(KEYINPUT5), .Z(n1110) );
NAND2_X1 U792 ( .A1(G125), .A2(n1112), .ZN(n1111) );
NOR2_X1 U793 ( .A1(G125), .A2(n1112), .ZN(n1109) );
NAND3_X1 U794 ( .A1(G953), .A2(n1113), .A3(KEYINPUT23), .ZN(n1097) );
NAND2_X1 U795 ( .A1(G900), .A2(G227), .ZN(n1113) );
AND2_X1 U796 ( .A1(n1114), .A2(n1071), .ZN(n1095) );
XOR2_X1 U797 ( .A(n1115), .B(n1116), .Z(G69) );
XOR2_X1 U798 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
INV_X1 U800 ( .A(n1121), .ZN(n1120) );
XOR2_X1 U801 ( .A(n1122), .B(n1123), .Z(n1119) );
NAND2_X1 U802 ( .A1(KEYINPUT52), .A2(n1124), .ZN(n1122) );
NAND2_X1 U803 ( .A1(n1125), .A2(n1071), .ZN(n1117) );
NOR2_X1 U804 ( .A1(n1126), .A2(n1071), .ZN(n1115) );
AND2_X1 U805 ( .A1(G224), .A2(G898), .ZN(n1126) );
NOR2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XNOR2_X1 U807 ( .A(n1129), .B(n1130), .ZN(n1128) );
NOR2_X1 U808 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR3_X1 U809 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(G63) );
AND3_X1 U810 ( .A1(KEYINPUT60), .A2(n1136), .A3(G953), .ZN(n1135) );
NOR2_X1 U811 ( .A1(KEYINPUT60), .A2(n1137), .ZN(n1134) );
INV_X1 U812 ( .A(n1127), .ZN(n1137) );
NOR2_X1 U813 ( .A1(n1138), .A2(n1139), .ZN(n1133) );
XOR2_X1 U814 ( .A(KEYINPUT30), .B(n1140), .Z(n1139) );
NOR3_X1 U815 ( .A1(n1141), .A2(n1142), .A3(n1132), .ZN(n1140) );
XOR2_X1 U816 ( .A(KEYINPUT32), .B(n1143), .Z(n1141) );
NOR2_X1 U817 ( .A1(n1144), .A2(n1143), .ZN(n1138) );
NOR2_X1 U818 ( .A1(n1142), .A2(n1132), .ZN(n1144) );
INV_X1 U819 ( .A(G478), .ZN(n1142) );
NOR2_X1 U820 ( .A1(n1127), .A2(n1145), .ZN(G60) );
NOR3_X1 U821 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1145) );
AND3_X1 U822 ( .A1(n1149), .A2(G475), .A3(n1150), .ZN(n1148) );
INV_X1 U823 ( .A(n1132), .ZN(n1150) );
NOR2_X1 U824 ( .A1(n1151), .A2(n1149), .ZN(n1147) );
AND2_X1 U825 ( .A1(n1043), .A2(G475), .ZN(n1151) );
XOR2_X1 U826 ( .A(G104), .B(n1152), .Z(G6) );
NOR3_X1 U827 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(G57) );
NOR2_X1 U828 ( .A1(G101), .A2(n1156), .ZN(n1155) );
XOR2_X1 U829 ( .A(KEYINPUT36), .B(n1157), .Z(n1156) );
AND2_X1 U830 ( .A1(n1157), .A2(G101), .ZN(n1154) );
XNOR2_X1 U831 ( .A(n1158), .B(n1159), .ZN(n1157) );
NAND2_X1 U832 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
NAND2_X1 U833 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U834 ( .A(KEYINPUT26), .B(n1164), .Z(n1162) );
NOR2_X1 U835 ( .A1(n1165), .A2(n1132), .ZN(n1164) );
OR3_X1 U836 ( .A1(n1132), .A2(n1165), .A3(n1163), .ZN(n1160) );
XOR2_X1 U837 ( .A(n1166), .B(n1167), .Z(n1163) );
NAND2_X1 U838 ( .A1(KEYINPUT33), .A2(n1168), .ZN(n1166) );
INV_X1 U839 ( .A(G472), .ZN(n1165) );
NOR2_X1 U840 ( .A1(n1169), .A2(n1136), .ZN(n1153) );
XOR2_X1 U841 ( .A(n1071), .B(KEYINPUT37), .Z(n1169) );
NOR2_X1 U842 ( .A1(n1127), .A2(n1170), .ZN(G54) );
XOR2_X1 U843 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U844 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U845 ( .A1(n1092), .A2(n1132), .ZN(n1174) );
NOR2_X1 U846 ( .A1(n1175), .A2(n1176), .ZN(n1173) );
XOR2_X1 U847 ( .A(n1177), .B(KEYINPUT43), .Z(n1176) );
NAND2_X1 U848 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NOR2_X1 U849 ( .A1(n1179), .A2(n1180), .ZN(n1175) );
XNOR2_X1 U850 ( .A(KEYINPUT51), .B(n1178), .ZN(n1180) );
NAND2_X1 U851 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
NAND2_X1 U852 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
INV_X1 U853 ( .A(KEYINPUT16), .ZN(n1184) );
NAND3_X1 U854 ( .A1(n1108), .A2(n1185), .A3(KEYINPUT16), .ZN(n1181) );
XOR2_X1 U855 ( .A(n1186), .B(n1187), .Z(n1171) );
NAND2_X1 U856 ( .A1(KEYINPUT8), .A2(n1188), .ZN(n1186) );
NOR2_X1 U857 ( .A1(n1127), .A2(n1189), .ZN(G51) );
XOR2_X1 U858 ( .A(n1190), .B(n1191), .Z(n1189) );
XOR2_X1 U859 ( .A(n1192), .B(n1193), .Z(n1191) );
NOR2_X1 U860 ( .A1(n1194), .A2(n1132), .ZN(n1193) );
NAND2_X1 U861 ( .A1(G902), .A2(n1043), .ZN(n1132) );
OR2_X1 U862 ( .A1(n1114), .A2(n1125), .ZN(n1043) );
NAND4_X1 U863 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1125) );
NOR4_X1 U864 ( .A1(n1199), .A2(n1200), .A3(n1152), .A4(n1038), .ZN(n1198) );
AND3_X1 U865 ( .A1(n1073), .A2(n1201), .A3(n1202), .ZN(n1038) );
AND3_X1 U866 ( .A1(n1202), .A2(n1073), .A3(n1203), .ZN(n1152) );
NOR2_X1 U867 ( .A1(n1204), .A2(n1205), .ZN(n1197) );
NOR2_X1 U868 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
XOR2_X1 U869 ( .A(n1208), .B(KEYINPUT17), .Z(n1206) );
NAND3_X1 U870 ( .A1(n1066), .A2(n1062), .A3(n1209), .ZN(n1208) );
XOR2_X1 U871 ( .A(n1210), .B(KEYINPUT38), .Z(n1209) );
NOR3_X1 U872 ( .A1(n1211), .A2(n1068), .A3(n1212), .ZN(n1204) );
INV_X1 U873 ( .A(n1201), .ZN(n1068) );
NAND4_X1 U874 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1114) );
AND4_X1 U875 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1216) );
NOR2_X1 U876 ( .A1(n1221), .A2(n1222), .ZN(n1215) );
NOR2_X1 U877 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XOR2_X1 U878 ( .A(KEYINPUT35), .B(n1079), .Z(n1224) );
NAND4_X1 U879 ( .A1(n1225), .A2(n1226), .A3(n1066), .A4(n1063), .ZN(n1214) );
XOR2_X1 U880 ( .A(n1227), .B(KEYINPUT48), .Z(n1226) );
XOR2_X1 U881 ( .A(n1056), .B(KEYINPUT28), .Z(n1225) );
NAND3_X1 U882 ( .A1(n1228), .A2(n1203), .A3(n1229), .ZN(n1213) );
NOR3_X1 U883 ( .A1(n1212), .A2(n1230), .A3(n1069), .ZN(n1229) );
XOR2_X1 U884 ( .A(n1227), .B(KEYINPUT55), .Z(n1230) );
XOR2_X1 U885 ( .A(n1061), .B(KEYINPUT24), .Z(n1228) );
NOR3_X1 U886 ( .A1(n1231), .A2(KEYINPUT20), .A3(G953), .ZN(n1192) );
XOR2_X1 U887 ( .A(n1232), .B(n1233), .Z(n1190) );
NOR2_X1 U888 ( .A1(n1136), .A2(n1071), .ZN(n1127) );
XOR2_X1 U889 ( .A(G952), .B(KEYINPUT4), .Z(n1136) );
XOR2_X1 U890 ( .A(G146), .B(n1221), .Z(G48) );
AND3_X1 U891 ( .A1(n1056), .A2(n1234), .A3(n1203), .ZN(n1221) );
XNOR2_X1 U892 ( .A(G143), .B(n1220), .ZN(G45) );
NAND4_X1 U893 ( .A1(n1056), .A2(n1235), .A3(n1088), .A4(n1236), .ZN(n1220) );
XOR2_X1 U894 ( .A(G140), .B(n1237), .Z(G42) );
NOR2_X1 U895 ( .A1(n1238), .A2(n1219), .ZN(n1237) );
NAND4_X1 U896 ( .A1(n1063), .A2(n1203), .A3(n1239), .A4(n1075), .ZN(n1219) );
NOR2_X1 U897 ( .A1(n1240), .A2(n1069), .ZN(n1239) );
XNOR2_X1 U898 ( .A(KEYINPUT45), .B(KEYINPUT34), .ZN(n1238) );
XOR2_X1 U899 ( .A(n1241), .B(n1242), .Z(G39) );
OR2_X1 U900 ( .A1(n1223), .A2(n1050), .ZN(n1242) );
NAND2_X1 U901 ( .A1(n1075), .A2(n1234), .ZN(n1223) );
XNOR2_X1 U902 ( .A(G134), .B(n1218), .ZN(G36) );
NAND3_X1 U903 ( .A1(n1075), .A2(n1201), .A3(n1235), .ZN(n1218) );
XOR2_X1 U904 ( .A(n1243), .B(n1244), .Z(G33) );
NAND3_X1 U905 ( .A1(n1235), .A2(n1075), .A3(n1203), .ZN(n1244) );
INV_X1 U906 ( .A(n1061), .ZN(n1075) );
NAND3_X1 U907 ( .A1(n1087), .A2(n1057), .A3(n1245), .ZN(n1061) );
NOR3_X1 U908 ( .A1(n1069), .A2(n1240), .A3(n1212), .ZN(n1235) );
XOR2_X1 U909 ( .A(n1246), .B(n1217), .Z(G30) );
NAND3_X1 U910 ( .A1(n1056), .A2(n1201), .A3(n1234), .ZN(n1217) );
NOR4_X1 U911 ( .A1(n1069), .A2(n1247), .A3(n1248), .A4(n1240), .ZN(n1234) );
INV_X1 U912 ( .A(n1227), .ZN(n1240) );
XOR2_X1 U913 ( .A(G101), .B(n1200), .Z(G3) );
AND3_X1 U914 ( .A1(n1062), .A2(n1202), .A3(n1079), .ZN(n1200) );
XNOR2_X1 U915 ( .A(G125), .B(n1249), .ZN(G27) );
NAND4_X1 U916 ( .A1(n1066), .A2(n1063), .A3(n1056), .A4(n1227), .ZN(n1249) );
NAND2_X1 U917 ( .A1(n1045), .A2(n1250), .ZN(n1227) );
NAND4_X1 U918 ( .A1(G902), .A2(G953), .A3(n1251), .A4(n1101), .ZN(n1250) );
INV_X1 U919 ( .A(G900), .ZN(n1101) );
XOR2_X1 U920 ( .A(n1252), .B(n1195), .Z(G24) );
NAND4_X1 U921 ( .A1(n1253), .A2(n1073), .A3(n1088), .A4(n1236), .ZN(n1195) );
INV_X1 U922 ( .A(n1054), .ZN(n1073) );
NAND2_X1 U923 ( .A1(n1248), .A2(n1247), .ZN(n1054) );
XNOR2_X1 U924 ( .A(G119), .B(n1196), .ZN(G21) );
OR4_X1 U925 ( .A1(n1211), .A2(n1050), .A3(n1247), .A4(n1248), .ZN(n1196) );
INV_X1 U926 ( .A(n1079), .ZN(n1050) );
XNOR2_X1 U927 ( .A(G116), .B(n1254), .ZN(G18) );
NAND3_X1 U928 ( .A1(n1253), .A2(n1201), .A3(n1255), .ZN(n1254) );
XOR2_X1 U929 ( .A(n1212), .B(KEYINPUT27), .Z(n1255) );
NOR2_X1 U930 ( .A1(n1236), .A2(n1256), .ZN(n1201) );
INV_X1 U931 ( .A(n1211), .ZN(n1253) );
NAND3_X1 U932 ( .A1(n1056), .A2(n1210), .A3(n1257), .ZN(n1211) );
XOR2_X1 U933 ( .A(n1207), .B(KEYINPUT39), .Z(n1056) );
XNOR2_X1 U934 ( .A(G113), .B(n1258), .ZN(G15) );
NAND4_X1 U935 ( .A1(KEYINPUT7), .A2(n1066), .A3(n1259), .A4(n1062), .ZN(n1258) );
INV_X1 U936 ( .A(n1212), .ZN(n1062) );
NAND2_X1 U937 ( .A1(n1247), .A2(n1260), .ZN(n1212) );
NOR2_X1 U938 ( .A1(n1261), .A2(n1207), .ZN(n1259) );
AND2_X1 U939 ( .A1(n1257), .A2(n1203), .ZN(n1066) );
AND2_X1 U940 ( .A1(n1256), .A2(n1236), .ZN(n1203) );
INV_X1 U941 ( .A(n1048), .ZN(n1257) );
NAND2_X1 U942 ( .A1(n1262), .A2(n1263), .ZN(n1048) );
INV_X1 U943 ( .A(n1078), .ZN(n1262) );
XOR2_X1 U944 ( .A(G110), .B(n1199), .Z(G12) );
AND3_X1 U945 ( .A1(n1063), .A2(n1202), .A3(n1079), .ZN(n1199) );
NOR2_X1 U946 ( .A1(n1088), .A2(n1236), .ZN(n1079) );
XOR2_X1 U947 ( .A(G475), .B(n1264), .Z(n1236) );
NOR2_X1 U948 ( .A1(KEYINPUT11), .A2(n1093), .ZN(n1264) );
INV_X1 U949 ( .A(n1146), .ZN(n1093) );
NOR2_X1 U950 ( .A1(n1149), .A2(G902), .ZN(n1146) );
XNOR2_X1 U951 ( .A(n1265), .B(n1266), .ZN(n1149) );
XOR2_X1 U952 ( .A(n1267), .B(n1268), .Z(n1266) );
XNOR2_X1 U953 ( .A(n1269), .B(n1270), .ZN(n1268) );
NAND2_X1 U954 ( .A1(KEYINPUT47), .A2(G104), .ZN(n1269) );
XOR2_X1 U955 ( .A(n1271), .B(n1272), .Z(n1267) );
NAND2_X1 U956 ( .A1(KEYINPUT54), .A2(n1273), .ZN(n1272) );
NAND2_X1 U957 ( .A1(n1274), .A2(n1275), .ZN(n1271) );
NAND2_X1 U958 ( .A1(G113), .A2(n1252), .ZN(n1275) );
XOR2_X1 U959 ( .A(n1276), .B(KEYINPUT49), .Z(n1274) );
OR2_X1 U960 ( .A1(n1252), .A2(G113), .ZN(n1276) );
INV_X1 U961 ( .A(G122), .ZN(n1252) );
XOR2_X1 U962 ( .A(n1277), .B(n1278), .Z(n1265) );
XOR2_X1 U963 ( .A(G125), .B(n1279), .Z(n1278) );
AND3_X1 U964 ( .A1(G214), .A2(n1071), .A3(n1280), .ZN(n1279) );
XOR2_X1 U965 ( .A(n1243), .B(KEYINPUT9), .Z(n1277) );
INV_X1 U966 ( .A(G131), .ZN(n1243) );
INV_X1 U967 ( .A(n1256), .ZN(n1088) );
XOR2_X1 U968 ( .A(n1281), .B(G478), .Z(n1256) );
OR2_X1 U969 ( .A1(n1143), .A2(G902), .ZN(n1281) );
XNOR2_X1 U970 ( .A(n1282), .B(n1283), .ZN(n1143) );
XOR2_X1 U971 ( .A(G122), .B(n1284), .Z(n1283) );
NOR2_X1 U972 ( .A1(KEYINPUT41), .A2(n1285), .ZN(n1284) );
XOR2_X1 U973 ( .A(G134), .B(n1286), .Z(n1285) );
NOR2_X1 U974 ( .A1(KEYINPUT1), .A2(n1287), .ZN(n1286) );
XOR2_X1 U975 ( .A(G143), .B(n1246), .Z(n1287) );
XOR2_X1 U976 ( .A(n1288), .B(n1289), .Z(n1282) );
NAND2_X1 U977 ( .A1(n1290), .A2(G217), .ZN(n1288) );
NOR3_X1 U978 ( .A1(n1207), .A2(n1261), .A3(n1069), .ZN(n1202) );
NAND2_X1 U979 ( .A1(n1263), .A2(n1078), .ZN(n1069) );
XOR2_X1 U980 ( .A(n1091), .B(n1092), .Z(n1078) );
INV_X1 U981 ( .A(G469), .ZN(n1092) );
NAND2_X1 U982 ( .A1(n1291), .A2(n1292), .ZN(n1091) );
XNOR2_X1 U983 ( .A(n1293), .B(n1178), .ZN(n1291) );
XOR2_X1 U984 ( .A(n1294), .B(n1295), .Z(n1293) );
NOR2_X1 U985 ( .A1(KEYINPUT13), .A2(n1183), .ZN(n1295) );
XOR2_X1 U986 ( .A(n1108), .B(n1185), .Z(n1183) );
XOR2_X1 U987 ( .A(n1296), .B(n1297), .Z(n1185) );
INV_X1 U988 ( .A(G107), .ZN(n1296) );
XNOR2_X1 U989 ( .A(n1298), .B(KEYINPUT2), .ZN(n1108) );
NAND2_X1 U990 ( .A1(n1299), .A2(n1300), .ZN(n1294) );
OR2_X1 U991 ( .A1(n1301), .A2(KEYINPUT6), .ZN(n1300) );
XOR2_X1 U992 ( .A(n1302), .B(n1188), .Z(n1299) );
AND2_X1 U993 ( .A1(G227), .A2(n1071), .ZN(n1188) );
NAND2_X1 U994 ( .A1(KEYINPUT6), .A2(n1301), .ZN(n1302) );
XOR2_X1 U995 ( .A(n1187), .B(KEYINPUT12), .Z(n1301) );
XOR2_X1 U996 ( .A(n1303), .B(n1112), .Z(n1187) );
XOR2_X1 U997 ( .A(n1080), .B(KEYINPUT42), .Z(n1263) );
NAND2_X1 U998 ( .A1(G221), .A2(n1304), .ZN(n1080) );
INV_X1 U999 ( .A(n1210), .ZN(n1261) );
NAND2_X1 U1000 ( .A1(n1045), .A2(n1305), .ZN(n1210) );
NAND3_X1 U1001 ( .A1(n1121), .A2(n1251), .A3(G902), .ZN(n1305) );
NOR2_X1 U1002 ( .A1(n1071), .A2(G898), .ZN(n1121) );
NAND3_X1 U1003 ( .A1(n1251), .A2(n1071), .A3(G952), .ZN(n1045) );
NAND2_X1 U1004 ( .A1(G237), .A2(G234), .ZN(n1251) );
NAND2_X1 U1005 ( .A1(n1057), .A2(n1306), .ZN(n1207) );
NAND2_X1 U1006 ( .A1(n1245), .A2(n1087), .ZN(n1306) );
INV_X1 U1007 ( .A(n1058), .ZN(n1087) );
NOR2_X1 U1008 ( .A1(n1307), .A2(n1308), .ZN(n1058) );
NOR2_X1 U1009 ( .A1(n1280), .A2(n1194), .ZN(n1308) );
INV_X1 U1010 ( .A(n1059), .ZN(n1245) );
XOR2_X1 U1011 ( .A(n1086), .B(KEYINPUT46), .Z(n1059) );
NAND3_X1 U1012 ( .A1(n1309), .A2(n1307), .A3(G210), .ZN(n1086) );
NAND2_X1 U1013 ( .A1(n1310), .A2(n1292), .ZN(n1307) );
XOR2_X1 U1014 ( .A(n1232), .B(n1311), .Z(n1310) );
XNOR2_X1 U1015 ( .A(n1312), .B(KEYINPUT58), .ZN(n1311) );
NAND2_X1 U1016 ( .A1(n1313), .A2(KEYINPUT62), .ZN(n1312) );
XNOR2_X1 U1017 ( .A(n1233), .B(n1314), .ZN(n1313) );
NOR2_X1 U1018 ( .A1(G953), .A2(n1231), .ZN(n1314) );
INV_X1 U1019 ( .A(G224), .ZN(n1231) );
XOR2_X1 U1020 ( .A(n1298), .B(n1315), .Z(n1233) );
XOR2_X1 U1021 ( .A(KEYINPUT10), .B(G125), .Z(n1315) );
XOR2_X1 U1022 ( .A(n1124), .B(n1123), .Z(n1232) );
AND2_X1 U1023 ( .A1(n1316), .A2(n1317), .ZN(n1123) );
NAND2_X1 U1024 ( .A1(G122), .A2(n1303), .ZN(n1317) );
INV_X1 U1025 ( .A(G110), .ZN(n1303) );
XOR2_X1 U1026 ( .A(KEYINPUT3), .B(n1318), .Z(n1316) );
NOR2_X1 U1027 ( .A1(G122), .A2(n1319), .ZN(n1318) );
XOR2_X1 U1028 ( .A(KEYINPUT63), .B(G110), .Z(n1319) );
XNOR2_X1 U1029 ( .A(n1297), .B(n1320), .ZN(n1124) );
XOR2_X1 U1030 ( .A(n1289), .B(n1321), .Z(n1320) );
XOR2_X1 U1031 ( .A(G107), .B(G116), .Z(n1289) );
XOR2_X1 U1032 ( .A(G104), .B(G101), .Z(n1297) );
NAND2_X1 U1033 ( .A1(G214), .A2(n1309), .ZN(n1057) );
NAND2_X1 U1034 ( .A1(n1280), .A2(n1292), .ZN(n1309) );
INV_X1 U1035 ( .A(G237), .ZN(n1280) );
NOR2_X1 U1036 ( .A1(n1260), .A2(n1247), .ZN(n1063) );
XNOR2_X1 U1037 ( .A(n1322), .B(n1131), .ZN(n1247) );
NAND2_X1 U1038 ( .A1(G217), .A2(n1304), .ZN(n1131) );
NAND2_X1 U1039 ( .A1(G234), .A2(n1292), .ZN(n1304) );
NAND2_X1 U1040 ( .A1(n1129), .A2(n1292), .ZN(n1322) );
XNOR2_X1 U1041 ( .A(n1323), .B(n1324), .ZN(n1129) );
XOR2_X1 U1042 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1043 ( .A(G137), .B(G110), .Z(n1326) );
XOR2_X1 U1044 ( .A(KEYINPUT18), .B(KEYINPUT14), .Z(n1325) );
XOR2_X1 U1045 ( .A(n1327), .B(n1328), .Z(n1323) );
AND2_X1 U1046 ( .A1(G221), .A2(n1290), .ZN(n1328) );
AND2_X1 U1047 ( .A1(G234), .A2(n1071), .ZN(n1290) );
INV_X1 U1048 ( .A(G953), .ZN(n1071) );
XOR2_X1 U1049 ( .A(n1329), .B(n1330), .Z(n1327) );
NOR3_X1 U1050 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(n1330) );
NOR2_X1 U1051 ( .A1(G128), .A2(n1334), .ZN(n1333) );
NOR2_X1 U1052 ( .A1(KEYINPUT40), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1053 ( .A(KEYINPUT0), .B(G119), .Z(n1335) );
NOR3_X1 U1054 ( .A1(n1246), .A2(KEYINPUT40), .A3(G119), .ZN(n1332) );
INV_X1 U1055 ( .A(G128), .ZN(n1246) );
AND2_X1 U1056 ( .A1(G119), .A2(KEYINPUT40), .ZN(n1331) );
NAND3_X1 U1057 ( .A1(n1336), .A2(n1337), .A3(n1338), .ZN(n1329) );
NAND2_X1 U1058 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
INV_X1 U1059 ( .A(KEYINPUT57), .ZN(n1340) );
NAND3_X1 U1060 ( .A1(KEYINPUT57), .A2(n1341), .A3(n1342), .ZN(n1337) );
OR2_X1 U1061 ( .A1(n1342), .A2(n1341), .ZN(n1336) );
NOR2_X1 U1062 ( .A1(KEYINPUT29), .A2(n1339), .ZN(n1341) );
XOR2_X1 U1063 ( .A(G125), .B(n1273), .Z(n1339) );
XOR2_X1 U1064 ( .A(n1112), .B(KEYINPUT15), .Z(n1273) );
INV_X1 U1065 ( .A(G140), .ZN(n1112) );
INV_X1 U1066 ( .A(G146), .ZN(n1342) );
INV_X1 U1067 ( .A(n1248), .ZN(n1260) );
XOR2_X1 U1068 ( .A(n1343), .B(G472), .Z(n1248) );
NAND2_X1 U1069 ( .A1(n1344), .A2(n1292), .ZN(n1343) );
INV_X1 U1070 ( .A(G902), .ZN(n1292) );
XOR2_X1 U1071 ( .A(n1345), .B(n1346), .Z(n1344) );
XNOR2_X1 U1072 ( .A(n1159), .B(n1347), .ZN(n1346) );
XNOR2_X1 U1073 ( .A(G101), .B(KEYINPUT22), .ZN(n1347) );
NOR3_X1 U1074 ( .A1(G237), .A2(G953), .A3(n1194), .ZN(n1159) );
INV_X1 U1075 ( .A(G210), .ZN(n1194) );
XOR2_X1 U1076 ( .A(n1168), .B(n1167), .Z(n1345) );
XNOR2_X1 U1077 ( .A(n1348), .B(n1321), .ZN(n1167) );
XOR2_X1 U1078 ( .A(G113), .B(G119), .Z(n1321) );
XNOR2_X1 U1079 ( .A(G116), .B(KEYINPUT31), .ZN(n1348) );
XOR2_X1 U1080 ( .A(n1178), .B(n1298), .Z(n1168) );
XOR2_X1 U1081 ( .A(G128), .B(n1270), .Z(n1298) );
XOR2_X1 U1082 ( .A(G143), .B(G146), .Z(n1270) );
XOR2_X1 U1083 ( .A(n1349), .B(n1350), .Z(n1178) );
XOR2_X1 U1084 ( .A(G134), .B(G131), .Z(n1350) );
NAND2_X1 U1085 ( .A1(n1351), .A2(n1241), .ZN(n1349) );
INV_X1 U1086 ( .A(G137), .ZN(n1241) );
XNOR2_X1 U1087 ( .A(KEYINPUT59), .B(KEYINPUT53), .ZN(n1351) );
endmodule


