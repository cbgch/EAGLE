//Key = 1100111110110001111001110101010101111100010100011111011100010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372;

XOR2_X1 U756 ( .A(G107), .B(n1047), .Z(G9) );
AND2_X1 U757 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND3_X1 U758 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(G75) );
NAND2_X1 U759 ( .A1(G952), .A2(n1053), .ZN(n1052) );
NAND3_X1 U760 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NAND4_X1 U761 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1055) );
NOR3_X1 U762 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NOR2_X1 U763 ( .A1(KEYINPUT24), .A2(n1064), .ZN(n1063) );
NAND2_X1 U764 ( .A1(n1065), .A2(n1066), .ZN(n1058) );
NAND2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U766 ( .A1(KEYINPUT24), .A2(n1064), .ZN(n1068) );
NAND2_X1 U767 ( .A1(n1069), .A2(n1070), .ZN(n1057) );
NAND2_X1 U768 ( .A1(n1064), .A2(n1071), .ZN(n1070) );
OR2_X1 U769 ( .A1(n1049), .A2(n1072), .ZN(n1071) );
NAND4_X1 U770 ( .A1(n1073), .A2(n1074), .A3(n1067), .A4(n1075), .ZN(n1054) );
NOR2_X1 U771 ( .A1(n1076), .A2(n1065), .ZN(n1075) );
NAND2_X1 U772 ( .A1(n1062), .A2(n1077), .ZN(n1074) );
NAND2_X1 U773 ( .A1(n1059), .A2(n1078), .ZN(n1077) );
NAND3_X1 U774 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1073) );
NAND2_X1 U775 ( .A1(n1059), .A2(n1082), .ZN(n1080) );
NAND2_X1 U776 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U777 ( .A1(n1078), .A2(n1085), .ZN(n1079) );
NAND2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U779 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U780 ( .A1(n1090), .A2(n1091), .ZN(n1050) );
NOR4_X1 U781 ( .A1(n1088), .A2(n1062), .A3(n1061), .A4(n1092), .ZN(n1091) );
XOR2_X1 U782 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR4_X1 U783 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1090) );
XOR2_X1 U784 ( .A(KEYINPUT46), .B(n1099), .Z(n1098) );
XNOR2_X1 U785 ( .A(G475), .B(n1100), .ZN(n1097) );
NOR2_X1 U786 ( .A1(G469), .A2(n1101), .ZN(n1096) );
XNOR2_X1 U787 ( .A(KEYINPUT34), .B(n1102), .ZN(n1101) );
AND2_X1 U788 ( .A1(n1102), .A2(G469), .ZN(n1095) );
XOR2_X1 U789 ( .A(n1103), .B(n1104), .Z(G72) );
XOR2_X1 U790 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U791 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
AND2_X1 U792 ( .A1(G227), .A2(G900), .ZN(n1107) );
NAND2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1105) );
NAND2_X1 U794 ( .A1(G953), .A2(n1111), .ZN(n1110) );
XOR2_X1 U795 ( .A(n1112), .B(n1113), .Z(n1109) );
XOR2_X1 U796 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U797 ( .A1(KEYINPUT27), .A2(n1116), .ZN(n1114) );
XNOR2_X1 U798 ( .A(G131), .B(n1117), .ZN(n1116) );
NAND2_X1 U799 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U800 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U801 ( .A(KEYINPUT16), .B(n1122), .Z(n1118) );
NOR2_X1 U802 ( .A1(n1120), .A2(n1121), .ZN(n1122) );
XNOR2_X1 U803 ( .A(n1123), .B(n1124), .ZN(n1112) );
XOR2_X1 U804 ( .A(KEYINPUT57), .B(KEYINPUT22), .Z(n1124) );
NAND2_X1 U805 ( .A1(n1051), .A2(n1125), .ZN(n1103) );
XOR2_X1 U806 ( .A(n1126), .B(n1127), .Z(G69) );
XOR2_X1 U807 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U808 ( .A1(n1130), .A2(n1108), .ZN(n1129) );
XNOR2_X1 U809 ( .A(G953), .B(KEYINPUT3), .ZN(n1108) );
NOR2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U811 ( .A1(n1133), .A2(n1134), .ZN(n1128) );
NAND2_X1 U812 ( .A1(G953), .A2(n1132), .ZN(n1134) );
XOR2_X1 U813 ( .A(n1135), .B(n1136), .Z(n1133) );
NAND2_X1 U814 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
XNOR2_X1 U815 ( .A(KEYINPUT63), .B(KEYINPUT56), .ZN(n1137) );
NAND2_X1 U816 ( .A1(n1051), .A2(n1139), .ZN(n1126) );
NOR2_X1 U817 ( .A1(n1140), .A2(n1141), .ZN(G66) );
XOR2_X1 U818 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U819 ( .A1(n1144), .A2(n1145), .ZN(n1142) );
INV_X1 U820 ( .A(n1146), .ZN(n1145) );
NOR2_X1 U821 ( .A1(n1140), .A2(n1147), .ZN(G63) );
XOR2_X1 U822 ( .A(n1148), .B(n1149), .Z(n1147) );
AND2_X1 U823 ( .A1(G478), .A2(n1146), .ZN(n1148) );
NOR2_X1 U824 ( .A1(n1140), .A2(n1150), .ZN(G60) );
XOR2_X1 U825 ( .A(n1151), .B(n1152), .Z(n1150) );
AND2_X1 U826 ( .A1(G475), .A2(n1146), .ZN(n1151) );
XNOR2_X1 U827 ( .A(n1153), .B(n1154), .ZN(G6) );
NOR2_X1 U828 ( .A1(n1140), .A2(n1155), .ZN(G57) );
XOR2_X1 U829 ( .A(n1156), .B(n1157), .Z(n1155) );
XNOR2_X1 U830 ( .A(n1158), .B(n1159), .ZN(n1157) );
XNOR2_X1 U831 ( .A(n1160), .B(n1161), .ZN(n1156) );
XNOR2_X1 U832 ( .A(n1162), .B(KEYINPUT32), .ZN(n1161) );
NAND3_X1 U833 ( .A1(n1146), .A2(G472), .A3(KEYINPUT7), .ZN(n1162) );
NOR2_X1 U834 ( .A1(n1140), .A2(n1163), .ZN(G54) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(n1163) );
AND2_X1 U836 ( .A1(G469), .A2(n1146), .ZN(n1165) );
NOR3_X1 U837 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1164) );
NOR2_X1 U838 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
INV_X1 U839 ( .A(KEYINPUT31), .ZN(n1170) );
NOR2_X1 U840 ( .A1(n1171), .A2(n1172), .ZN(n1169) );
AND2_X1 U841 ( .A1(n1173), .A2(KEYINPUT39), .ZN(n1172) );
NOR3_X1 U842 ( .A1(KEYINPUT39), .A2(n1173), .A3(n1174), .ZN(n1171) );
NOR2_X1 U843 ( .A1(KEYINPUT31), .A2(n1175), .ZN(n1167) );
NOR2_X1 U844 ( .A1(n1174), .A2(n1176), .ZN(n1175) );
XNOR2_X1 U845 ( .A(n1177), .B(KEYINPUT39), .ZN(n1176) );
AND2_X1 U846 ( .A1(n1173), .A2(n1174), .ZN(n1166) );
XOR2_X1 U847 ( .A(n1178), .B(n1115), .Z(n1174) );
XNOR2_X1 U848 ( .A(n1179), .B(n1180), .ZN(n1178) );
NAND2_X1 U849 ( .A1(KEYINPUT25), .A2(n1181), .ZN(n1180) );
NAND2_X1 U850 ( .A1(KEYINPUT6), .A2(n1159), .ZN(n1179) );
NOR2_X1 U851 ( .A1(n1140), .A2(n1182), .ZN(G51) );
NOR2_X1 U852 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XOR2_X1 U853 ( .A(n1185), .B(KEYINPUT47), .Z(n1184) );
NAND2_X1 U854 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NOR2_X1 U855 ( .A1(n1186), .A2(n1187), .ZN(n1183) );
NAND3_X1 U856 ( .A1(G210), .A2(n1188), .A3(n1146), .ZN(n1187) );
NOR2_X1 U857 ( .A1(n1189), .A2(n1056), .ZN(n1146) );
NOR2_X1 U858 ( .A1(n1125), .A2(n1139), .ZN(n1056) );
NAND4_X1 U859 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1139) );
NOR4_X1 U860 ( .A1(n1194), .A2(n1154), .A3(n1195), .A4(n1196), .ZN(n1193) );
NOR2_X1 U861 ( .A1(n1084), .A2(n1197), .ZN(n1196) );
NOR4_X1 U862 ( .A1(n1061), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1195) );
XNOR2_X1 U863 ( .A(KEYINPUT38), .B(n1201), .ZN(n1200) );
AND2_X1 U864 ( .A1(n1072), .A2(n1048), .ZN(n1154) );
NOR3_X1 U865 ( .A1(n1061), .A2(n1202), .A3(n1198), .ZN(n1048) );
INV_X1 U866 ( .A(n1078), .ZN(n1061) );
NOR2_X1 U867 ( .A1(n1203), .A2(n1204), .ZN(n1192) );
NAND4_X1 U868 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1125) );
NOR4_X1 U869 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1208) );
INV_X1 U870 ( .A(n1213), .ZN(n1210) );
NOR2_X1 U871 ( .A1(n1214), .A2(n1215), .ZN(n1207) );
INV_X1 U872 ( .A(n1216), .ZN(n1215) );
XNOR2_X1 U873 ( .A(n1217), .B(KEYINPUT48), .ZN(n1189) );
XNOR2_X1 U874 ( .A(n1218), .B(n1219), .ZN(n1186) );
NAND2_X1 U875 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
NAND2_X1 U876 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
INV_X1 U877 ( .A(n1224), .ZN(n1223) );
NAND2_X1 U878 ( .A1(n1225), .A2(n1224), .ZN(n1220) );
NAND3_X1 U879 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1224) );
NAND2_X1 U880 ( .A1(KEYINPUT13), .A2(n1229), .ZN(n1228) );
NAND3_X1 U881 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1227) );
NAND2_X1 U882 ( .A1(G125), .A2(n1233), .ZN(n1226) );
NAND2_X1 U883 ( .A1(n1234), .A2(n1231), .ZN(n1233) );
INV_X1 U884 ( .A(KEYINPUT13), .ZN(n1231) );
XNOR2_X1 U885 ( .A(KEYINPUT45), .B(n1229), .ZN(n1234) );
XNOR2_X1 U886 ( .A(n1222), .B(KEYINPUT2), .ZN(n1225) );
NOR2_X1 U887 ( .A1(n1051), .A2(G952), .ZN(n1140) );
XNOR2_X1 U888 ( .A(G146), .B(n1205), .ZN(G48) );
NAND3_X1 U889 ( .A1(n1235), .A2(n1072), .A3(n1236), .ZN(n1205) );
XOR2_X1 U890 ( .A(n1206), .B(n1237), .Z(G45) );
NAND2_X1 U891 ( .A1(KEYINPUT49), .A2(G143), .ZN(n1237) );
NAND4_X1 U892 ( .A1(n1235), .A2(n1238), .A3(n1239), .A4(n1099), .ZN(n1206) );
XNOR2_X1 U893 ( .A(n1240), .B(n1214), .ZN(G42) );
AND3_X1 U894 ( .A1(n1059), .A2(n1065), .A3(n1241), .ZN(n1214) );
XOR2_X1 U895 ( .A(G137), .B(n1212), .Z(G39) );
AND3_X1 U896 ( .A1(n1059), .A2(n1067), .A3(n1236), .ZN(n1212) );
XNOR2_X1 U897 ( .A(G134), .B(n1242), .ZN(G36) );
NAND2_X1 U898 ( .A1(KEYINPUT11), .A2(n1211), .ZN(n1242) );
AND3_X1 U899 ( .A1(n1059), .A2(n1049), .A3(n1238), .ZN(n1211) );
XNOR2_X1 U900 ( .A(G131), .B(n1213), .ZN(G33) );
NAND3_X1 U901 ( .A1(n1072), .A2(n1059), .A3(n1238), .ZN(n1213) );
AND3_X1 U902 ( .A1(n1243), .A2(n1244), .A3(n1245), .ZN(n1238) );
NOR2_X1 U903 ( .A1(n1246), .A2(n1088), .ZN(n1059) );
XNOR2_X1 U904 ( .A(G128), .B(n1216), .ZN(G30) );
NAND3_X1 U905 ( .A1(n1235), .A2(n1049), .A3(n1236), .ZN(n1216) );
AND4_X1 U906 ( .A1(n1243), .A2(n1247), .A3(n1248), .A4(n1244), .ZN(n1236) );
XOR2_X1 U907 ( .A(G101), .B(n1194), .Z(G3) );
NOR2_X1 U908 ( .A1(n1197), .A2(n1083), .ZN(n1194) );
INV_X1 U909 ( .A(n1245), .ZN(n1083) );
NAND3_X1 U910 ( .A1(n1249), .A2(n1201), .A3(n1067), .ZN(n1197) );
XNOR2_X1 U911 ( .A(n1232), .B(n1209), .ZN(G27) );
AND3_X1 U912 ( .A1(n1235), .A2(n1069), .A3(n1241), .ZN(n1209) );
AND4_X1 U913 ( .A1(n1072), .A2(n1250), .A3(n1244), .A4(n1081), .ZN(n1241) );
NAND2_X1 U914 ( .A1(n1251), .A2(n1252), .ZN(n1244) );
NAND2_X1 U915 ( .A1(n1253), .A2(n1111), .ZN(n1252) );
INV_X1 U916 ( .A(G900), .ZN(n1111) );
XNOR2_X1 U917 ( .A(G122), .B(n1190), .ZN(G24) );
NAND4_X1 U918 ( .A1(n1239), .A2(n1254), .A3(n1078), .A4(n1099), .ZN(n1190) );
NOR2_X1 U919 ( .A1(n1248), .A2(n1247), .ZN(n1078) );
XNOR2_X1 U920 ( .A(G119), .B(n1255), .ZN(G21) );
NAND2_X1 U921 ( .A1(KEYINPUT43), .A2(n1256), .ZN(n1255) );
INV_X1 U922 ( .A(n1191), .ZN(n1256) );
NAND4_X1 U923 ( .A1(n1254), .A2(n1067), .A3(n1247), .A4(n1248), .ZN(n1191) );
XOR2_X1 U924 ( .A(G116), .B(n1204), .Z(G18) );
AND3_X1 U925 ( .A1(n1245), .A2(n1049), .A3(n1254), .ZN(n1204) );
AND2_X1 U926 ( .A1(n1257), .A2(n1235), .ZN(n1254) );
INV_X1 U927 ( .A(n1086), .ZN(n1235) );
XOR2_X1 U928 ( .A(n1258), .B(KEYINPUT53), .Z(n1086) );
INV_X1 U929 ( .A(n1199), .ZN(n1049) );
NAND2_X1 U930 ( .A1(n1099), .A2(n1259), .ZN(n1199) );
XOR2_X1 U931 ( .A(G113), .B(n1203), .Z(G15) );
AND4_X1 U932 ( .A1(n1257), .A2(n1245), .A3(n1072), .A4(n1258), .ZN(n1203) );
NOR2_X1 U933 ( .A1(n1259), .A2(n1099), .ZN(n1072) );
NOR2_X1 U934 ( .A1(n1247), .A2(n1260), .ZN(n1245) );
NOR3_X1 U935 ( .A1(n1202), .A2(n1062), .A3(n1065), .ZN(n1257) );
INV_X1 U936 ( .A(n1069), .ZN(n1065) );
INV_X1 U937 ( .A(n1201), .ZN(n1202) );
XNOR2_X1 U938 ( .A(G110), .B(n1261), .ZN(G12) );
NAND4_X1 U939 ( .A1(n1250), .A2(n1067), .A3(n1249), .A4(n1262), .ZN(n1261) );
XNOR2_X1 U940 ( .A(KEYINPUT4), .B(n1201), .ZN(n1262) );
NAND2_X1 U941 ( .A1(n1251), .A2(n1263), .ZN(n1201) );
NAND2_X1 U942 ( .A1(n1253), .A2(n1132), .ZN(n1263) );
INV_X1 U943 ( .A(G898), .ZN(n1132) );
NOR3_X1 U944 ( .A1(n1217), .A2(n1076), .A3(n1051), .ZN(n1253) );
NAND3_X1 U945 ( .A1(G952), .A2(n1051), .A3(n1264), .ZN(n1251) );
XNOR2_X1 U946 ( .A(n1076), .B(KEYINPUT30), .ZN(n1264) );
INV_X1 U947 ( .A(n1064), .ZN(n1076) );
NAND2_X1 U948 ( .A1(G237), .A2(G234), .ZN(n1064) );
INV_X1 U949 ( .A(n1198), .ZN(n1249) );
NAND2_X1 U950 ( .A1(n1243), .A2(n1258), .ZN(n1198) );
NOR2_X1 U951 ( .A1(n1089), .A2(n1088), .ZN(n1258) );
AND2_X1 U952 ( .A1(G214), .A2(n1188), .ZN(n1088) );
INV_X1 U953 ( .A(n1246), .ZN(n1089) );
NAND2_X1 U954 ( .A1(n1265), .A2(n1266), .ZN(n1246) );
NAND2_X1 U955 ( .A1(n1267), .A2(n1093), .ZN(n1266) );
XOR2_X1 U956 ( .A(KEYINPUT50), .B(n1268), .Z(n1265) );
NOR2_X1 U957 ( .A1(n1267), .A2(n1093), .ZN(n1268) );
NAND2_X1 U958 ( .A1(n1269), .A2(n1217), .ZN(n1093) );
XNOR2_X1 U959 ( .A(n1219), .B(n1270), .ZN(n1269) );
NOR2_X1 U960 ( .A1(KEYINPUT12), .A2(n1271), .ZN(n1270) );
XNOR2_X1 U961 ( .A(n1230), .B(n1272), .ZN(n1271) );
XNOR2_X1 U962 ( .A(n1232), .B(n1222), .ZN(n1272) );
NOR2_X1 U963 ( .A1(n1131), .A2(G953), .ZN(n1222) );
INV_X1 U964 ( .A(G224), .ZN(n1131) );
INV_X1 U965 ( .A(n1229), .ZN(n1230) );
XNOR2_X1 U966 ( .A(n1136), .B(n1138), .ZN(n1219) );
XNOR2_X1 U967 ( .A(n1273), .B(G110), .ZN(n1138) );
NAND2_X1 U968 ( .A1(KEYINPUT0), .A2(n1274), .ZN(n1273) );
XOR2_X1 U969 ( .A(n1275), .B(n1276), .Z(n1136) );
XOR2_X1 U970 ( .A(G113), .B(n1277), .Z(n1276) );
XNOR2_X1 U971 ( .A(KEYINPUT52), .B(n1278), .ZN(n1277) );
INV_X1 U972 ( .A(G119), .ZN(n1278) );
XOR2_X1 U973 ( .A(n1279), .B(n1280), .Z(n1275) );
XNOR2_X1 U974 ( .A(n1281), .B(n1282), .ZN(n1279) );
NAND2_X1 U975 ( .A1(KEYINPUT5), .A2(n1153), .ZN(n1281) );
XOR2_X1 U976 ( .A(n1094), .B(KEYINPUT35), .Z(n1267) );
NAND2_X1 U977 ( .A1(n1283), .A2(n1188), .ZN(n1094) );
NAND2_X1 U978 ( .A1(n1284), .A2(n1217), .ZN(n1188) );
XOR2_X1 U979 ( .A(KEYINPUT44), .B(G210), .Z(n1283) );
NOR2_X1 U980 ( .A1(n1069), .A2(n1062), .ZN(n1243) );
INV_X1 U981 ( .A(n1081), .ZN(n1062) );
NAND2_X1 U982 ( .A1(G221), .A2(n1285), .ZN(n1081) );
XOR2_X1 U983 ( .A(n1102), .B(G469), .Z(n1069) );
NAND2_X1 U984 ( .A1(n1286), .A2(n1217), .ZN(n1102) );
XOR2_X1 U985 ( .A(n1287), .B(n1288), .Z(n1286) );
XNOR2_X1 U986 ( .A(n1115), .B(n1173), .ZN(n1288) );
INV_X1 U987 ( .A(n1177), .ZN(n1173) );
XNOR2_X1 U988 ( .A(n1289), .B(n1290), .ZN(n1177) );
XNOR2_X1 U989 ( .A(n1240), .B(G110), .ZN(n1290) );
NAND2_X1 U990 ( .A1(G227), .A2(n1051), .ZN(n1289) );
XNOR2_X1 U991 ( .A(n1291), .B(n1292), .ZN(n1115) );
NOR2_X1 U992 ( .A1(KEYINPUT62), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U993 ( .A(n1159), .B(n1181), .ZN(n1287) );
XOR2_X1 U994 ( .A(n1280), .B(G104), .Z(n1181) );
XOR2_X1 U995 ( .A(G107), .B(n1294), .Z(n1280) );
NOR2_X1 U996 ( .A1(n1099), .A2(n1239), .ZN(n1067) );
INV_X1 U997 ( .A(n1259), .ZN(n1239) );
XNOR2_X1 U998 ( .A(n1100), .B(n1295), .ZN(n1259) );
NOR2_X1 U999 ( .A1(G475), .A2(KEYINPUT26), .ZN(n1295) );
OR2_X1 U1000 ( .A1(n1152), .A2(G902), .ZN(n1100) );
XNOR2_X1 U1001 ( .A(n1296), .B(n1297), .ZN(n1152) );
XNOR2_X1 U1002 ( .A(n1153), .B(n1298), .ZN(n1297) );
NOR2_X1 U1003 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XOR2_X1 U1004 ( .A(n1301), .B(KEYINPUT61), .Z(n1300) );
NAND2_X1 U1005 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NOR2_X1 U1006 ( .A1(n1302), .A2(n1303), .ZN(n1299) );
XOR2_X1 U1007 ( .A(n1304), .B(n1305), .Z(n1303) );
AND2_X1 U1008 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U1009 ( .A1(G143), .A2(n1308), .ZN(n1307) );
XOR2_X1 U1010 ( .A(KEYINPUT36), .B(n1309), .Z(n1306) );
NOR2_X1 U1011 ( .A1(n1308), .A2(G143), .ZN(n1309) );
AND3_X1 U1012 ( .A1(n1284), .A2(n1051), .A3(G214), .ZN(n1308) );
NOR2_X1 U1013 ( .A1(KEYINPUT20), .A2(n1310), .ZN(n1304) );
XNOR2_X1 U1014 ( .A(KEYINPUT23), .B(n1311), .ZN(n1310) );
INV_X1 U1015 ( .A(G131), .ZN(n1311) );
AND2_X1 U1016 ( .A1(n1312), .A2(n1313), .ZN(n1302) );
NAND2_X1 U1017 ( .A1(G146), .A2(n1314), .ZN(n1313) );
NAND2_X1 U1018 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XNOR2_X1 U1019 ( .A(KEYINPUT33), .B(n1317), .ZN(n1315) );
NAND2_X1 U1020 ( .A1(n1318), .A2(n1319), .ZN(n1312) );
NAND2_X1 U1021 ( .A1(n1320), .A2(n1321), .ZN(n1318) );
OR2_X1 U1022 ( .A1(n1317), .A2(KEYINPUT33), .ZN(n1321) );
NAND2_X1 U1023 ( .A1(n1123), .A2(KEYINPUT33), .ZN(n1320) );
INV_X1 U1024 ( .A(G104), .ZN(n1153) );
XNOR2_X1 U1025 ( .A(G113), .B(n1322), .ZN(n1296) );
XNOR2_X1 U1026 ( .A(KEYINPUT15), .B(n1274), .ZN(n1322) );
XNOR2_X1 U1027 ( .A(n1323), .B(G478), .ZN(n1099) );
OR2_X1 U1028 ( .A1(n1149), .A2(G902), .ZN(n1323) );
XNOR2_X1 U1029 ( .A(n1324), .B(n1325), .ZN(n1149) );
XOR2_X1 U1030 ( .A(n1326), .B(n1327), .Z(n1325) );
XNOR2_X1 U1031 ( .A(n1293), .B(G107), .ZN(n1327) );
XOR2_X1 U1032 ( .A(KEYINPUT21), .B(G143), .Z(n1326) );
XOR2_X1 U1033 ( .A(n1328), .B(n1329), .Z(n1324) );
XOR2_X1 U1034 ( .A(n1330), .B(n1331), .Z(n1329) );
NAND2_X1 U1035 ( .A1(G217), .A2(n1332), .ZN(n1331) );
NAND2_X1 U1036 ( .A1(n1333), .A2(n1334), .ZN(n1330) );
NAND2_X1 U1037 ( .A1(n1282), .A2(G122), .ZN(n1334) );
XOR2_X1 U1038 ( .A(n1335), .B(KEYINPUT19), .Z(n1333) );
NAND2_X1 U1039 ( .A1(n1336), .A2(n1274), .ZN(n1335) );
INV_X1 U1040 ( .A(G122), .ZN(n1274) );
INV_X1 U1041 ( .A(n1084), .ZN(n1250) );
NAND2_X1 U1042 ( .A1(n1260), .A2(n1247), .ZN(n1084) );
XOR2_X1 U1043 ( .A(n1337), .B(n1144), .Z(n1247) );
NAND2_X1 U1044 ( .A1(G217), .A2(n1285), .ZN(n1144) );
NAND2_X1 U1045 ( .A1(G234), .A2(n1217), .ZN(n1285) );
NAND2_X1 U1046 ( .A1(n1338), .A2(n1217), .ZN(n1337) );
XNOR2_X1 U1047 ( .A(n1143), .B(KEYINPUT58), .ZN(n1338) );
XNOR2_X1 U1048 ( .A(n1339), .B(n1340), .ZN(n1143) );
NOR2_X1 U1049 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
NOR2_X1 U1050 ( .A1(n1343), .A2(n1120), .ZN(n1342) );
NOR2_X1 U1051 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
INV_X1 U1052 ( .A(KEYINPUT37), .ZN(n1345) );
NOR2_X1 U1053 ( .A1(n1346), .A2(n1347), .ZN(n1341) );
XNOR2_X1 U1054 ( .A(KEYINPUT8), .B(n1348), .ZN(n1347) );
NOR2_X1 U1055 ( .A1(n1349), .A2(n1344), .ZN(n1346) );
XOR2_X1 U1056 ( .A(n1348), .B(KEYINPUT14), .Z(n1344) );
NAND2_X1 U1057 ( .A1(n1332), .A2(n1350), .ZN(n1348) );
XOR2_X1 U1058 ( .A(KEYINPUT42), .B(G221), .Z(n1350) );
AND2_X1 U1059 ( .A1(G234), .A2(n1051), .ZN(n1332) );
AND2_X1 U1060 ( .A1(n1120), .A2(KEYINPUT37), .ZN(n1349) );
NAND2_X1 U1061 ( .A1(KEYINPUT29), .A2(n1351), .ZN(n1339) );
XOR2_X1 U1062 ( .A(n1352), .B(n1353), .Z(n1351) );
XOR2_X1 U1063 ( .A(n1354), .B(n1355), .Z(n1353) );
XNOR2_X1 U1064 ( .A(n1123), .B(G119), .ZN(n1355) );
AND2_X1 U1065 ( .A1(n1317), .A2(n1316), .ZN(n1123) );
NAND2_X1 U1066 ( .A1(G125), .A2(n1240), .ZN(n1316) );
INV_X1 U1067 ( .A(G140), .ZN(n1240) );
NAND2_X1 U1068 ( .A1(G140), .A2(n1232), .ZN(n1317) );
INV_X1 U1069 ( .A(G125), .ZN(n1232) );
NAND2_X1 U1070 ( .A1(KEYINPUT18), .A2(n1356), .ZN(n1354) );
INV_X1 U1071 ( .A(G110), .ZN(n1356) );
XNOR2_X1 U1072 ( .A(n1293), .B(n1357), .ZN(n1352) );
XNOR2_X1 U1073 ( .A(KEYINPUT9), .B(n1319), .ZN(n1357) );
INV_X1 U1074 ( .A(G146), .ZN(n1319) );
INV_X1 U1075 ( .A(G128), .ZN(n1293) );
INV_X1 U1076 ( .A(n1248), .ZN(n1260) );
XNOR2_X1 U1077 ( .A(n1358), .B(G472), .ZN(n1248) );
NAND2_X1 U1078 ( .A1(n1359), .A2(n1217), .ZN(n1358) );
INV_X1 U1079 ( .A(G902), .ZN(n1217) );
XOR2_X1 U1080 ( .A(n1360), .B(n1361), .Z(n1359) );
NOR2_X1 U1081 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
NOR2_X1 U1082 ( .A1(KEYINPUT40), .A2(n1160), .ZN(n1363) );
NOR2_X1 U1083 ( .A1(KEYINPUT41), .A2(n1364), .ZN(n1362) );
INV_X1 U1084 ( .A(n1160), .ZN(n1364) );
XNOR2_X1 U1085 ( .A(n1365), .B(n1294), .ZN(n1160) );
XOR2_X1 U1086 ( .A(G101), .B(KEYINPUT10), .Z(n1294) );
NAND3_X1 U1087 ( .A1(n1284), .A2(n1051), .A3(G210), .ZN(n1365) );
INV_X1 U1088 ( .A(G953), .ZN(n1051) );
INV_X1 U1089 ( .A(G237), .ZN(n1284) );
XOR2_X1 U1090 ( .A(n1366), .B(n1158), .Z(n1360) );
XNOR2_X1 U1091 ( .A(n1229), .B(n1367), .ZN(n1158) );
XOR2_X1 U1092 ( .A(G113), .B(n1368), .Z(n1367) );
NOR2_X1 U1093 ( .A1(KEYINPUT60), .A2(n1369), .ZN(n1368) );
XNOR2_X1 U1094 ( .A(G119), .B(n1370), .ZN(n1369) );
NAND2_X1 U1095 ( .A1(KEYINPUT54), .A2(n1282), .ZN(n1370) );
INV_X1 U1096 ( .A(n1336), .ZN(n1282) );
XOR2_X1 U1097 ( .A(G116), .B(KEYINPUT28), .Z(n1336) );
XOR2_X1 U1098 ( .A(G128), .B(n1291), .Z(n1229) );
XNOR2_X1 U1099 ( .A(G143), .B(G146), .ZN(n1291) );
NAND2_X1 U1100 ( .A1(n1371), .A2(n1159), .ZN(n1366) );
XOR2_X1 U1101 ( .A(n1372), .B(n1121), .Z(n1159) );
XNOR2_X1 U1102 ( .A(n1328), .B(KEYINPUT51), .ZN(n1121) );
XNOR2_X1 U1103 ( .A(G134), .B(KEYINPUT17), .ZN(n1328) );
XNOR2_X1 U1104 ( .A(G131), .B(n1120), .ZN(n1372) );
XOR2_X1 U1105 ( .A(G137), .B(KEYINPUT59), .Z(n1120) );
XNOR2_X1 U1106 ( .A(KEYINPUT55), .B(KEYINPUT1), .ZN(n1371) );
endmodule


