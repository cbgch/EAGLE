//Key = 0001001010011001101011111001100111010110011110000111001111110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;

XOR2_X1 U742 ( .A(G107), .B(n1007), .Z(G9) );
NOR2_X1 U743 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
XOR2_X1 U744 ( .A(n1010), .B(KEYINPUT1), .Z(n1008) );
NOR2_X1 U745 ( .A1(n1011), .A2(n1012), .ZN(G75) );
NOR4_X1 U746 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
NAND2_X1 U747 ( .A1(n1017), .A2(n1018), .ZN(n1014) );
XOR2_X1 U748 ( .A(KEYINPUT54), .B(n1019), .Z(n1017) );
AND3_X1 U749 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1019) );
NAND4_X1 U750 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1013) );
NAND4_X1 U751 ( .A1(n1027), .A2(n1028), .A3(n1022), .A4(n1029), .ZN(n1024) );
NAND2_X1 U752 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U753 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U754 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U755 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
INV_X1 U756 ( .A(n1038), .ZN(n1034) );
NAND2_X1 U757 ( .A1(n1039), .A2(n1040), .ZN(n1030) );
NAND2_X1 U758 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
XOR2_X1 U759 ( .A(n1043), .B(KEYINPUT2), .Z(n1041) );
NAND2_X1 U760 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U761 ( .A1(n1020), .A2(n1046), .ZN(n1023) );
NAND2_X1 U762 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U763 ( .A1(n1028), .A2(n1049), .ZN(n1048) );
NAND2_X1 U764 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U765 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U766 ( .A1(n1054), .A2(n1022), .ZN(n1047) );
AND3_X1 U767 ( .A1(n1032), .A2(n1039), .A3(n1027), .ZN(n1020) );
INV_X1 U768 ( .A(n1055), .ZN(n1027) );
NOR3_X1 U769 ( .A1(n1056), .A2(G953), .A3(G952), .ZN(n1011) );
INV_X1 U770 ( .A(n1025), .ZN(n1056) );
NAND4_X1 U771 ( .A1(n1057), .A2(n1022), .A3(n1058), .A4(n1059), .ZN(n1025) );
NOR3_X1 U772 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
XOR2_X1 U773 ( .A(n1063), .B(n1064), .Z(n1061) );
XNOR2_X1 U774 ( .A(KEYINPUT36), .B(n1065), .ZN(n1064) );
NAND2_X1 U775 ( .A1(KEYINPUT38), .A2(n1066), .ZN(n1063) );
XOR2_X1 U776 ( .A(n1067), .B(n1068), .Z(n1058) );
NAND2_X1 U777 ( .A1(KEYINPUT37), .A2(G478), .ZN(n1067) );
XNOR2_X1 U778 ( .A(n1069), .B(G472), .ZN(n1057) );
XOR2_X1 U779 ( .A(n1070), .B(n1071), .Z(G72) );
XOR2_X1 U780 ( .A(n1072), .B(n1073), .Z(n1071) );
NOR2_X1 U781 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XOR2_X1 U782 ( .A(n1076), .B(n1077), .Z(n1075) );
XNOR2_X1 U783 ( .A(n1078), .B(n1079), .ZN(n1077) );
NAND3_X1 U784 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1078) );
NAND2_X1 U785 ( .A1(KEYINPUT48), .A2(n1083), .ZN(n1082) );
NAND2_X1 U786 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U787 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND4_X1 U788 ( .A1(n1084), .A2(n1088), .A3(KEYINPUT51), .A4(n1086), .ZN(n1081) );
NAND2_X1 U789 ( .A1(G131), .A2(n1089), .ZN(n1080) );
NAND3_X1 U790 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
NAND2_X1 U791 ( .A1(KEYINPUT51), .A2(KEYINPUT48), .ZN(n1092) );
NAND2_X1 U792 ( .A1(KEYINPUT20), .A2(n1093), .ZN(n1091) );
NAND2_X1 U793 ( .A1(n1084), .A2(n1094), .ZN(n1093) );
NAND2_X1 U794 ( .A1(n1088), .A2(n1087), .ZN(n1094) );
INV_X1 U795 ( .A(KEYINPUT51), .ZN(n1087) );
INV_X1 U796 ( .A(KEYINPUT48), .ZN(n1088) );
NAND2_X1 U797 ( .A1(n1084), .A2(n1095), .ZN(n1090) );
INV_X1 U798 ( .A(KEYINPUT20), .ZN(n1095) );
XOR2_X1 U799 ( .A(n1096), .B(n1097), .Z(n1084) );
NAND2_X1 U800 ( .A1(KEYINPUT32), .A2(n1098), .ZN(n1096) );
INV_X1 U801 ( .A(G137), .ZN(n1098) );
NOR2_X1 U802 ( .A1(G953), .A2(n1099), .ZN(n1072) );
NOR2_X1 U803 ( .A1(n1015), .A2(n1100), .ZN(n1099) );
XNOR2_X1 U804 ( .A(KEYINPUT6), .B(n1101), .ZN(n1100) );
NOR3_X1 U805 ( .A1(n1026), .A2(KEYINPUT46), .A3(n1102), .ZN(n1070) );
AND2_X1 U806 ( .A1(G227), .A2(G900), .ZN(n1102) );
XOR2_X1 U807 ( .A(n1103), .B(n1104), .Z(G69) );
XOR2_X1 U808 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U809 ( .A1(n1107), .A2(n1026), .ZN(n1106) );
AND2_X1 U810 ( .A1(G224), .A2(G898), .ZN(n1107) );
NOR2_X1 U811 ( .A1(KEYINPUT63), .A2(n1108), .ZN(n1105) );
NOR2_X1 U812 ( .A1(G953), .A2(n1109), .ZN(n1108) );
XOR2_X1 U813 ( .A(n1016), .B(KEYINPUT49), .Z(n1109) );
NAND2_X1 U814 ( .A1(n1110), .A2(n1111), .ZN(n1103) );
NAND2_X1 U815 ( .A1(n1112), .A2(G953), .ZN(n1111) );
XOR2_X1 U816 ( .A(n1113), .B(n1114), .Z(n1110) );
XNOR2_X1 U817 ( .A(KEYINPUT21), .B(n1115), .ZN(n1114) );
XNOR2_X1 U818 ( .A(n1116), .B(n1117), .ZN(n1113) );
NOR2_X1 U819 ( .A1(KEYINPUT29), .A2(n1118), .ZN(n1117) );
XOR2_X1 U820 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U821 ( .A1(KEYINPUT24), .A2(n1121), .ZN(n1119) );
XNOR2_X1 U822 ( .A(n1122), .B(n1123), .ZN(n1121) );
INV_X1 U823 ( .A(G113), .ZN(n1122) );
NOR2_X1 U824 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XOR2_X1 U825 ( .A(n1126), .B(n1127), .Z(n1125) );
OR2_X1 U826 ( .A1(n1128), .A2(n1065), .ZN(n1126) );
NOR2_X1 U827 ( .A1(n1124), .A2(n1129), .ZN(G63) );
NOR2_X1 U828 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U829 ( .A(n1132), .B(KEYINPUT58), .Z(n1131) );
NAND2_X1 U830 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U831 ( .A1(n1133), .A2(n1134), .ZN(n1130) );
AND2_X1 U832 ( .A1(n1135), .A2(G478), .ZN(n1133) );
NOR2_X1 U833 ( .A1(n1124), .A2(n1136), .ZN(G60) );
XOR2_X1 U834 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U835 ( .A1(n1135), .A2(G475), .ZN(n1137) );
XNOR2_X1 U836 ( .A(n1139), .B(n1140), .ZN(G6) );
NAND2_X1 U837 ( .A1(KEYINPUT12), .A2(n1141), .ZN(n1139) );
NOR2_X1 U838 ( .A1(n1124), .A2(n1142), .ZN(G57) );
XOR2_X1 U839 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U840 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND2_X1 U841 ( .A1(KEYINPUT16), .A2(n1147), .ZN(n1145) );
XOR2_X1 U842 ( .A(n1148), .B(n1149), .Z(n1143) );
XNOR2_X1 U843 ( .A(n1150), .B(n1151), .ZN(n1149) );
NAND2_X1 U844 ( .A1(n1135), .A2(G472), .ZN(n1148) );
INV_X1 U845 ( .A(n1128), .ZN(n1135) );
NOR2_X1 U846 ( .A1(n1124), .A2(n1152), .ZN(G54) );
XOR2_X1 U847 ( .A(n1153), .B(n1154), .Z(n1152) );
XNOR2_X1 U848 ( .A(n1155), .B(n1156), .ZN(n1154) );
NAND2_X1 U849 ( .A1(KEYINPUT41), .A2(n1115), .ZN(n1155) );
XOR2_X1 U850 ( .A(n1157), .B(n1158), .Z(n1153) );
NOR3_X1 U851 ( .A1(n1128), .A2(KEYINPUT47), .A3(n1159), .ZN(n1158) );
XNOR2_X1 U852 ( .A(G140), .B(KEYINPUT61), .ZN(n1157) );
NOR2_X1 U853 ( .A1(n1124), .A2(n1160), .ZN(G51) );
XOR2_X1 U854 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U855 ( .A(n1163), .B(n1164), .ZN(n1162) );
NOR3_X1 U856 ( .A1(n1128), .A2(KEYINPUT4), .A3(n1165), .ZN(n1164) );
NAND2_X1 U857 ( .A1(G902), .A2(n1166), .ZN(n1128) );
NAND3_X1 U858 ( .A1(n1167), .A2(n1018), .A3(n1168), .ZN(n1166) );
INV_X1 U859 ( .A(n1015), .ZN(n1168) );
NAND4_X1 U860 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1015) );
NAND2_X1 U861 ( .A1(n1173), .A2(n1032), .ZN(n1169) );
XNOR2_X1 U862 ( .A(n1174), .B(KEYINPUT57), .ZN(n1173) );
XNOR2_X1 U863 ( .A(n1101), .B(KEYINPUT34), .ZN(n1018) );
NAND3_X1 U864 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1101) );
NAND2_X1 U865 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND2_X1 U866 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NAND2_X1 U867 ( .A1(n1182), .A2(n1054), .ZN(n1181) );
XNOR2_X1 U868 ( .A(KEYINPUT39), .B(n1016), .ZN(n1167) );
NAND2_X1 U869 ( .A1(n1183), .A2(n1184), .ZN(n1016) );
AND4_X1 U870 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1184) );
NOR4_X1 U871 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1183) );
NOR2_X1 U872 ( .A1(n1010), .A2(n1009), .ZN(n1192) );
NAND4_X1 U873 ( .A1(n1193), .A2(n1021), .A3(n1039), .A4(n1194), .ZN(n1010) );
INV_X1 U874 ( .A(n1141), .ZN(n1191) );
NAND3_X1 U875 ( .A1(n1195), .A2(n1039), .A3(n1054), .ZN(n1141) );
NAND2_X1 U876 ( .A1(KEYINPUT22), .A2(n1196), .ZN(n1163) );
XNOR2_X1 U877 ( .A(n1197), .B(n1198), .ZN(n1196) );
XNOR2_X1 U878 ( .A(G125), .B(n1199), .ZN(n1198) );
NOR2_X1 U879 ( .A1(n1026), .A2(G952), .ZN(n1124) );
XNOR2_X1 U880 ( .A(G146), .B(n1200), .ZN(G48) );
NAND4_X1 U881 ( .A1(KEYINPUT15), .A2(n1182), .A3(n1054), .A4(n1178), .ZN(n1200) );
XOR2_X1 U882 ( .A(G143), .B(n1201), .Z(G45) );
NOR3_X1 U883 ( .A1(n1202), .A2(KEYINPUT30), .A3(n1042), .ZN(n1201) );
XOR2_X1 U884 ( .A(n1180), .B(KEYINPUT52), .Z(n1202) );
NAND3_X1 U885 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1180) );
XNOR2_X1 U886 ( .A(n1175), .B(n1206), .ZN(G42) );
XNOR2_X1 U887 ( .A(KEYINPUT19), .B(n1207), .ZN(n1206) );
NAND3_X1 U888 ( .A1(n1032), .A2(n1193), .A3(n1208), .ZN(n1175) );
XNOR2_X1 U889 ( .A(G137), .B(n1176), .ZN(G39) );
NAND3_X1 U890 ( .A1(n1028), .A2(n1032), .A3(n1182), .ZN(n1176) );
XNOR2_X1 U891 ( .A(G134), .B(n1209), .ZN(G36) );
NAND2_X1 U892 ( .A1(n1174), .A2(n1032), .ZN(n1209) );
AND2_X1 U893 ( .A1(n1205), .A2(n1021), .ZN(n1174) );
XOR2_X1 U894 ( .A(n1170), .B(n1210), .Z(G33) );
NAND2_X1 U895 ( .A1(KEYINPUT56), .A2(G131), .ZN(n1210) );
NAND3_X1 U896 ( .A1(n1054), .A2(n1032), .A3(n1205), .ZN(n1170) );
AND3_X1 U897 ( .A1(n1193), .A2(n1211), .A3(n1038), .ZN(n1205) );
INV_X1 U898 ( .A(n1060), .ZN(n1032) );
NAND2_X1 U899 ( .A1(n1045), .A2(n1212), .ZN(n1060) );
XNOR2_X1 U900 ( .A(G128), .B(n1171), .ZN(G30) );
NAND3_X1 U901 ( .A1(n1021), .A2(n1178), .A3(n1182), .ZN(n1171) );
AND4_X1 U902 ( .A1(n1036), .A2(n1193), .A3(n1213), .A4(n1211), .ZN(n1182) );
NAND2_X1 U903 ( .A1(n1214), .A2(n1215), .ZN(G3) );
NAND2_X1 U904 ( .A1(n1190), .A2(n1150), .ZN(n1215) );
XOR2_X1 U905 ( .A(KEYINPUT33), .B(n1216), .Z(n1214) );
NOR2_X1 U906 ( .A1(n1190), .A2(n1150), .ZN(n1216) );
INV_X1 U907 ( .A(G101), .ZN(n1150) );
AND3_X1 U908 ( .A1(n1028), .A2(n1195), .A3(n1038), .ZN(n1190) );
XNOR2_X1 U909 ( .A(G125), .B(n1172), .ZN(G27) );
NAND3_X1 U910 ( .A1(n1022), .A2(n1178), .A3(n1208), .ZN(n1172) );
AND4_X1 U911 ( .A1(n1036), .A2(n1054), .A3(n1037), .A4(n1211), .ZN(n1208) );
NAND2_X1 U912 ( .A1(n1055), .A2(n1217), .ZN(n1211) );
NAND3_X1 U913 ( .A1(G902), .A2(n1218), .A3(n1074), .ZN(n1217) );
NOR2_X1 U914 ( .A1(n1026), .A2(G900), .ZN(n1074) );
INV_X1 U915 ( .A(n1219), .ZN(n1022) );
XOR2_X1 U916 ( .A(G122), .B(n1189), .Z(G24) );
AND4_X1 U917 ( .A1(n1203), .A2(n1220), .A3(n1039), .A4(n1204), .ZN(n1189) );
NOR2_X1 U918 ( .A1(n1213), .A2(n1036), .ZN(n1039) );
XNOR2_X1 U919 ( .A(G119), .B(n1188), .ZN(G21) );
NAND4_X1 U920 ( .A1(n1220), .A2(n1028), .A3(n1213), .A4(n1036), .ZN(n1188) );
INV_X1 U921 ( .A(n1037), .ZN(n1213) );
XNOR2_X1 U922 ( .A(G116), .B(n1187), .ZN(G18) );
NAND3_X1 U923 ( .A1(n1038), .A2(n1021), .A3(n1220), .ZN(n1187) );
NOR3_X1 U924 ( .A1(n1042), .A2(n1221), .A3(n1219), .ZN(n1220) );
INV_X1 U925 ( .A(n1178), .ZN(n1042) );
XNOR2_X1 U926 ( .A(n1009), .B(KEYINPUT10), .ZN(n1178) );
NOR2_X1 U927 ( .A1(n1203), .A2(n1222), .ZN(n1021) );
XNOR2_X1 U928 ( .A(G113), .B(n1186), .ZN(G15) );
NAND3_X1 U929 ( .A1(n1038), .A2(n1054), .A3(n1223), .ZN(n1186) );
NOR3_X1 U930 ( .A1(n1219), .A2(n1221), .A3(n1009), .ZN(n1223) );
NAND2_X1 U931 ( .A1(n1053), .A2(n1224), .ZN(n1219) );
AND2_X1 U932 ( .A1(n1203), .A2(n1222), .ZN(n1054) );
INV_X1 U933 ( .A(n1204), .ZN(n1222) );
NOR2_X1 U934 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
XNOR2_X1 U935 ( .A(G110), .B(n1185), .ZN(G12) );
NAND4_X1 U936 ( .A1(n1028), .A2(n1195), .A3(n1037), .A4(n1036), .ZN(n1185) );
XNOR2_X1 U937 ( .A(n1225), .B(n1066), .ZN(n1036) );
NAND2_X1 U938 ( .A1(n1127), .A2(n1226), .ZN(n1066) );
XNOR2_X1 U939 ( .A(n1227), .B(n1228), .ZN(n1127) );
XNOR2_X1 U940 ( .A(G137), .B(n1229), .ZN(n1228) );
NAND3_X1 U941 ( .A1(n1230), .A2(n1026), .A3(G234), .ZN(n1229) );
XOR2_X1 U942 ( .A(KEYINPUT25), .B(G221), .Z(n1230) );
XNOR2_X1 U943 ( .A(n1231), .B(n1232), .ZN(n1227) );
NOR2_X1 U944 ( .A1(KEYINPUT53), .A2(n1233), .ZN(n1232) );
XNOR2_X1 U945 ( .A(G110), .B(n1234), .ZN(n1233) );
XNOR2_X1 U946 ( .A(n1235), .B(G119), .ZN(n1234) );
NAND2_X1 U947 ( .A1(KEYINPUT18), .A2(n1065), .ZN(n1225) );
NAND2_X1 U948 ( .A1(G217), .A2(n1236), .ZN(n1065) );
XOR2_X1 U949 ( .A(G472), .B(n1237), .Z(n1037) );
NOR2_X1 U950 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NOR2_X1 U951 ( .A1(KEYINPUT50), .A2(n1069), .ZN(n1239) );
AND2_X1 U952 ( .A1(KEYINPUT42), .A2(n1069), .ZN(n1238) );
AND2_X1 U953 ( .A1(n1226), .A2(n1240), .ZN(n1069) );
NAND2_X1 U954 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
NAND2_X1 U955 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XOR2_X1 U956 ( .A(n1245), .B(KEYINPUT26), .Z(n1241) );
OR2_X1 U957 ( .A1(n1244), .A2(n1243), .ZN(n1245) );
XOR2_X1 U958 ( .A(G101), .B(n1246), .Z(n1243) );
NOR2_X1 U959 ( .A1(n1151), .A2(KEYINPUT17), .ZN(n1246) );
AND3_X1 U960 ( .A1(G210), .A2(n1247), .A3(n1248), .ZN(n1151) );
XNOR2_X1 U961 ( .A(G953), .B(KEYINPUT7), .ZN(n1248) );
XOR2_X1 U962 ( .A(n1249), .B(n1197), .Z(n1244) );
XOR2_X1 U963 ( .A(n1146), .B(KEYINPUT5), .Z(n1249) );
XOR2_X1 U964 ( .A(n1250), .B(n1251), .Z(n1146) );
NOR2_X1 U965 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NOR3_X1 U966 ( .A1(KEYINPUT27), .A2(G119), .A3(n1254), .ZN(n1253) );
NOR2_X1 U967 ( .A1(n1123), .A2(n1255), .ZN(n1252) );
INV_X1 U968 ( .A(KEYINPUT27), .ZN(n1255) );
XNOR2_X1 U969 ( .A(G113), .B(n1256), .ZN(n1250) );
NOR3_X1 U970 ( .A1(n1050), .A2(n1221), .A3(n1009), .ZN(n1195) );
OR2_X1 U971 ( .A1(n1045), .A2(n1044), .ZN(n1009) );
INV_X1 U972 ( .A(n1212), .ZN(n1044) );
NAND2_X1 U973 ( .A1(G214), .A2(n1257), .ZN(n1212) );
XNOR2_X1 U974 ( .A(n1258), .B(n1165), .ZN(n1045) );
NAND2_X1 U975 ( .A1(G210), .A2(n1257), .ZN(n1165) );
NAND2_X1 U976 ( .A1(n1247), .A2(n1259), .ZN(n1257) );
NAND2_X1 U977 ( .A1(n1260), .A2(n1226), .ZN(n1258) );
XNOR2_X1 U978 ( .A(n1261), .B(n1161), .ZN(n1260) );
XNOR2_X1 U979 ( .A(n1262), .B(n1263), .ZN(n1161) );
XOR2_X1 U980 ( .A(n1123), .B(n1264), .Z(n1263) );
XNOR2_X1 U981 ( .A(n1254), .B(G119), .ZN(n1123) );
XNOR2_X1 U982 ( .A(n1265), .B(n1115), .ZN(n1262) );
INV_X1 U983 ( .A(G110), .ZN(n1115) );
NAND2_X1 U984 ( .A1(KEYINPUT11), .A2(n1120), .ZN(n1265) );
XNOR2_X1 U985 ( .A(G101), .B(n1266), .ZN(n1120) );
NAND3_X1 U986 ( .A1(KEYINPUT23), .A2(n1267), .A3(n1268), .ZN(n1261) );
XNOR2_X1 U987 ( .A(n1199), .B(n1269), .ZN(n1268) );
NOR2_X1 U988 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
AND2_X1 U989 ( .A1(G224), .A2(n1026), .ZN(n1199) );
NAND2_X1 U990 ( .A1(n1270), .A2(n1271), .ZN(n1267) );
INV_X1 U991 ( .A(KEYINPUT43), .ZN(n1271) );
NAND2_X1 U992 ( .A1(n1272), .A2(n1273), .ZN(n1270) );
NAND2_X1 U993 ( .A1(n1147), .A2(n1274), .ZN(n1273) );
INV_X1 U994 ( .A(G125), .ZN(n1274) );
NAND2_X1 U995 ( .A1(n1275), .A2(G125), .ZN(n1272) );
XNOR2_X1 U996 ( .A(KEYINPUT60), .B(n1147), .ZN(n1275) );
INV_X1 U997 ( .A(n1197), .ZN(n1147) );
XOR2_X1 U998 ( .A(n1276), .B(n1277), .Z(n1197) );
XNOR2_X1 U999 ( .A(n1278), .B(n1235), .ZN(n1276) );
NAND2_X1 U1000 ( .A1(KEYINPUT31), .A2(n1279), .ZN(n1278) );
INV_X1 U1001 ( .A(n1194), .ZN(n1221) );
NAND2_X1 U1002 ( .A1(n1055), .A2(n1280), .ZN(n1194) );
NAND4_X1 U1003 ( .A1(n1112), .A2(G953), .A3(G902), .A4(n1218), .ZN(n1280) );
XNOR2_X1 U1004 ( .A(G898), .B(KEYINPUT62), .ZN(n1112) );
NAND3_X1 U1005 ( .A1(n1218), .A2(n1026), .A3(G952), .ZN(n1055) );
NAND2_X1 U1006 ( .A1(G237), .A2(G234), .ZN(n1218) );
INV_X1 U1007 ( .A(n1193), .ZN(n1050) );
NOR2_X1 U1008 ( .A1(n1053), .A2(n1052), .ZN(n1193) );
INV_X1 U1009 ( .A(n1224), .ZN(n1052) );
NAND2_X1 U1010 ( .A1(G221), .A2(n1236), .ZN(n1224) );
NAND2_X1 U1011 ( .A1(G234), .A2(n1259), .ZN(n1236) );
XNOR2_X1 U1012 ( .A(n1281), .B(n1159), .ZN(n1053) );
INV_X1 U1013 ( .A(G469), .ZN(n1159) );
NAND2_X1 U1014 ( .A1(n1282), .A2(n1226), .ZN(n1281) );
XNOR2_X1 U1015 ( .A(n1283), .B(n1284), .ZN(n1282) );
XNOR2_X1 U1016 ( .A(n1207), .B(G110), .ZN(n1284) );
INV_X1 U1017 ( .A(G140), .ZN(n1207) );
INV_X1 U1018 ( .A(n1156), .ZN(n1283) );
XNOR2_X1 U1019 ( .A(n1285), .B(n1286), .ZN(n1156) );
XOR2_X1 U1020 ( .A(n1266), .B(n1076), .Z(n1286) );
XNOR2_X1 U1021 ( .A(n1287), .B(n1288), .ZN(n1076) );
NOR2_X1 U1022 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XOR2_X1 U1023 ( .A(KEYINPUT9), .B(n1291), .Z(n1290) );
NOR2_X1 U1024 ( .A1(n1277), .A2(n1279), .ZN(n1291) );
NOR2_X1 U1025 ( .A1(G146), .A2(n1292), .ZN(n1289) );
XNOR2_X1 U1026 ( .A(KEYINPUT0), .B(n1277), .ZN(n1292) );
XNOR2_X1 U1027 ( .A(G143), .B(KEYINPUT8), .ZN(n1277) );
NAND2_X1 U1028 ( .A1(KEYINPUT44), .A2(n1235), .ZN(n1287) );
XNOR2_X1 U1029 ( .A(n1140), .B(G107), .ZN(n1266) );
INV_X1 U1030 ( .A(G104), .ZN(n1140) );
XOR2_X1 U1031 ( .A(n1293), .B(n1256), .Z(n1285) );
XNOR2_X1 U1032 ( .A(n1294), .B(n1097), .ZN(n1256) );
XNOR2_X1 U1033 ( .A(G137), .B(G131), .ZN(n1294) );
XOR2_X1 U1034 ( .A(n1295), .B(n1296), .Z(n1293) );
NOR2_X1 U1035 ( .A1(G101), .A2(KEYINPUT45), .ZN(n1296) );
NAND2_X1 U1036 ( .A1(G227), .A2(n1026), .ZN(n1295) );
NOR2_X1 U1037 ( .A1(n1204), .A2(n1203), .ZN(n1028) );
XNOR2_X1 U1038 ( .A(n1062), .B(KEYINPUT55), .ZN(n1203) );
XNOR2_X1 U1039 ( .A(n1297), .B(G475), .ZN(n1062) );
NAND2_X1 U1040 ( .A1(n1138), .A2(n1226), .ZN(n1297) );
INV_X1 U1041 ( .A(n1298), .ZN(n1226) );
XOR2_X1 U1042 ( .A(n1264), .B(n1299), .Z(n1138) );
XNOR2_X1 U1043 ( .A(G104), .B(n1300), .ZN(n1299) );
NAND2_X1 U1044 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U1045 ( .A1(n1303), .A2(n1231), .ZN(n1302) );
XOR2_X1 U1046 ( .A(n1304), .B(KEYINPUT14), .Z(n1301) );
OR2_X1 U1047 ( .A1(n1231), .A2(n1303), .ZN(n1304) );
XNOR2_X1 U1048 ( .A(n1305), .B(n1306), .ZN(n1303) );
NOR2_X1 U1049 ( .A1(KEYINPUT40), .A2(n1086), .ZN(n1306) );
INV_X1 U1050 ( .A(G131), .ZN(n1086) );
XNOR2_X1 U1051 ( .A(G143), .B(n1307), .ZN(n1305) );
AND3_X1 U1052 ( .A1(G214), .A2(n1026), .A3(n1247), .ZN(n1307) );
INV_X1 U1053 ( .A(G237), .ZN(n1247) );
XNOR2_X1 U1054 ( .A(n1279), .B(n1079), .ZN(n1231) );
XOR2_X1 U1055 ( .A(G125), .B(G140), .Z(n1079) );
INV_X1 U1056 ( .A(G146), .ZN(n1279) );
XNOR2_X1 U1057 ( .A(G113), .B(n1308), .ZN(n1264) );
XOR2_X1 U1058 ( .A(n1068), .B(G478), .Z(n1204) );
NOR2_X1 U1059 ( .A1(n1134), .A2(n1298), .ZN(n1068) );
XOR2_X1 U1060 ( .A(n1259), .B(KEYINPUT28), .Z(n1298) );
INV_X1 U1061 ( .A(G902), .ZN(n1259) );
XNOR2_X1 U1062 ( .A(n1309), .B(n1310), .ZN(n1134) );
XOR2_X1 U1063 ( .A(n1311), .B(n1312), .Z(n1310) );
XNOR2_X1 U1064 ( .A(n1254), .B(G107), .ZN(n1312) );
INV_X1 U1065 ( .A(G116), .ZN(n1254) );
XNOR2_X1 U1066 ( .A(G143), .B(n1235), .ZN(n1311) );
INV_X1 U1067 ( .A(G128), .ZN(n1235) );
XNOR2_X1 U1068 ( .A(n1313), .B(n1308), .ZN(n1309) );
INV_X1 U1069 ( .A(n1116), .ZN(n1308) );
XOR2_X1 U1070 ( .A(G122), .B(KEYINPUT13), .Z(n1116) );
XOR2_X1 U1071 ( .A(n1314), .B(n1315), .Z(n1313) );
AND3_X1 U1072 ( .A1(G217), .A2(n1026), .A3(G234), .ZN(n1315) );
INV_X1 U1073 ( .A(G953), .ZN(n1026) );
NAND2_X1 U1074 ( .A1(n1316), .A2(n1097), .ZN(n1314) );
XOR2_X1 U1075 ( .A(G134), .B(KEYINPUT59), .Z(n1097) );
XNOR2_X1 U1076 ( .A(KEYINPUT35), .B(KEYINPUT3), .ZN(n1316) );
endmodule


