//Key = 1100000000100010000111010100011101110000000101010110001000101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361;

XOR2_X1 U748 ( .A(G107), .B(n1033), .Z(G9) );
NOR2_X1 U749 ( .A1(n1034), .A2(n1035), .ZN(G75) );
NOR4_X1 U750 ( .A1(G953), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1035) );
NOR2_X1 U751 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR2_X1 U752 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U753 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U754 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U756 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U760 ( .A1(n1057), .A2(n1058), .ZN(n1049) );
NOR2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR3_X1 U762 ( .A1(n1052), .A2(n1061), .A3(n1058), .ZN(n1045) );
NOR2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
XOR2_X1 U764 ( .A(n1064), .B(KEYINPUT10), .Z(n1063) );
NOR3_X1 U765 ( .A1(n1065), .A2(KEYINPUT27), .A3(n1066), .ZN(n1062) );
NOR4_X1 U766 ( .A1(n1066), .A2(n1058), .A3(n1048), .A4(n1052), .ZN(n1041) );
AND4_X1 U767 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
NAND2_X1 U768 ( .A1(KEYINPUT27), .A2(n1071), .ZN(n1067) );
NOR3_X1 U769 ( .A1(n1036), .A2(G953), .A3(G952), .ZN(n1034) );
AND4_X1 U770 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1036) );
NOR4_X1 U771 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1075) );
XOR2_X1 U772 ( .A(n1080), .B(KEYINPUT60), .Z(n1078) );
XOR2_X1 U773 ( .A(KEYINPUT61), .B(n1081), .Z(n1077) );
NOR2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U775 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XNOR2_X1 U776 ( .A(KEYINPUT43), .B(n1086), .ZN(n1085) );
NOR2_X1 U777 ( .A1(G472), .A2(n1087), .ZN(n1082) );
XOR2_X1 U778 ( .A(n1086), .B(KEYINPUT45), .Z(n1087) );
INV_X1 U779 ( .A(n1068), .ZN(n1076) );
XOR2_X1 U780 ( .A(n1088), .B(G478), .Z(n1074) );
XOR2_X1 U781 ( .A(n1089), .B(KEYINPUT39), .Z(n1072) );
NAND2_X1 U782 ( .A1(n1090), .A2(n1091), .ZN(G72) );
NAND3_X1 U783 ( .A1(n1092), .A2(n1093), .A3(G953), .ZN(n1091) );
XOR2_X1 U784 ( .A(n1094), .B(KEYINPUT52), .Z(n1090) );
NAND3_X1 U785 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1094) );
NAND2_X1 U786 ( .A1(n1098), .A2(n1093), .ZN(n1097) );
OR3_X1 U787 ( .A1(n1093), .A2(n1098), .A3(G953), .ZN(n1096) );
AND2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U789 ( .A(KEYINPUT58), .B(n1101), .ZN(n1100) );
NAND2_X1 U790 ( .A1(G953), .A2(n1102), .ZN(n1095) );
OR2_X1 U791 ( .A1(n1093), .A2(n1092), .ZN(n1102) );
NAND2_X1 U792 ( .A1(G900), .A2(G227), .ZN(n1092) );
NAND2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(n1093) );
NAND2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U795 ( .A(n1107), .B(KEYINPUT15), .Z(n1105) );
XOR2_X1 U796 ( .A(n1108), .B(n1109), .Z(n1103) );
XOR2_X1 U797 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U798 ( .A(G131), .B(n1112), .Z(n1108) );
NOR2_X1 U799 ( .A1(KEYINPUT6), .A2(n1113), .ZN(n1112) );
XOR2_X1 U800 ( .A(n1114), .B(n1115), .Z(G69) );
NAND2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND3_X1 U803 ( .A1(G898), .A2(G224), .A3(G953), .ZN(n1116) );
NAND2_X1 U804 ( .A1(n1120), .A2(n1121), .ZN(n1114) );
NAND2_X1 U805 ( .A1(n1106), .A2(n1122), .ZN(n1121) );
XOR2_X1 U806 ( .A(n1123), .B(n1124), .Z(n1120) );
XNOR2_X1 U807 ( .A(n1125), .B(KEYINPUT17), .ZN(n1123) );
NOR2_X1 U808 ( .A1(n1126), .A2(n1127), .ZN(G66) );
XOR2_X1 U809 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U810 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
NOR2_X1 U811 ( .A1(n1126), .A2(n1132), .ZN(G63) );
XOR2_X1 U812 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U813 ( .A1(n1135), .A2(n1131), .ZN(n1134) );
NAND2_X1 U814 ( .A1(KEYINPUT50), .A2(n1136), .ZN(n1133) );
NOR2_X1 U815 ( .A1(n1126), .A2(n1137), .ZN(G60) );
XNOR2_X1 U816 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR2_X1 U817 ( .A1(n1140), .A2(n1131), .ZN(n1139) );
INV_X1 U818 ( .A(G475), .ZN(n1140) );
XNOR2_X1 U819 ( .A(G104), .B(n1141), .ZN(G6) );
NAND2_X1 U820 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U821 ( .A1(KEYINPUT44), .A2(n1144), .ZN(n1143) );
OR2_X1 U822 ( .A1(KEYINPUT28), .A2(n1144), .ZN(n1142) );
INV_X1 U823 ( .A(n1145), .ZN(n1144) );
NOR2_X1 U824 ( .A1(n1126), .A2(n1146), .ZN(G57) );
XOR2_X1 U825 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U826 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U827 ( .A1(n1084), .A2(n1131), .ZN(n1149) );
INV_X1 U828 ( .A(G472), .ZN(n1084) );
XOR2_X1 U829 ( .A(n1151), .B(KEYINPUT48), .Z(n1147) );
NAND3_X1 U830 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
NAND2_X1 U831 ( .A1(KEYINPUT11), .A2(n1155), .ZN(n1154) );
NAND3_X1 U832 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1153) );
NAND2_X1 U833 ( .A1(n1159), .A2(n1160), .ZN(n1152) );
NAND2_X1 U834 ( .A1(n1161), .A2(n1157), .ZN(n1160) );
INV_X1 U835 ( .A(KEYINPUT11), .ZN(n1157) );
XOR2_X1 U836 ( .A(KEYINPUT3), .B(n1156), .Z(n1161) );
NOR2_X1 U837 ( .A1(n1126), .A2(n1162), .ZN(G54) );
XOR2_X1 U838 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U839 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U840 ( .A1(n1167), .A2(n1131), .ZN(n1166) );
INV_X1 U841 ( .A(G469), .ZN(n1167) );
NOR3_X1 U842 ( .A1(n1168), .A2(KEYINPUT59), .A3(n1169), .ZN(n1165) );
XOR2_X1 U843 ( .A(KEYINPUT7), .B(n1170), .Z(n1168) );
NOR2_X1 U844 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XNOR2_X1 U845 ( .A(n1173), .B(KEYINPUT31), .ZN(n1172) );
NOR2_X1 U846 ( .A1(n1126), .A2(n1174), .ZN(G51) );
XOR2_X1 U847 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U848 ( .A(n1177), .B(n1178), .Z(n1176) );
NOR2_X1 U849 ( .A1(n1179), .A2(n1131), .ZN(n1178) );
NAND2_X1 U850 ( .A1(G902), .A2(n1038), .ZN(n1131) );
NAND3_X1 U851 ( .A1(n1099), .A2(n1101), .A3(n1118), .ZN(n1038) );
AND4_X1 U852 ( .A1(n1145), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1118) );
NOR4_X1 U853 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1182) );
NOR3_X1 U854 ( .A1(n1070), .A2(n1187), .A3(n1052), .ZN(n1186) );
NOR2_X1 U855 ( .A1(n1033), .A2(n1188), .ZN(n1181) );
AND3_X1 U856 ( .A1(n1059), .A2(n1071), .A3(n1189), .ZN(n1033) );
NAND3_X1 U857 ( .A1(n1189), .A2(n1071), .A3(n1060), .ZN(n1145) );
AND4_X1 U858 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1099) );
NOR4_X1 U859 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
NOR2_X1 U860 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U861 ( .A(KEYINPUT21), .B(n1200), .Z(n1199) );
OR2_X1 U862 ( .A1(n1201), .A2(n1069), .ZN(n1192) );
NAND3_X1 U863 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1177) );
OR3_X1 U864 ( .A1(n1205), .A2(n1155), .A3(G125), .ZN(n1203) );
NAND2_X1 U865 ( .A1(n1206), .A2(G125), .ZN(n1202) );
XOR2_X1 U866 ( .A(n1205), .B(n1155), .Z(n1206) );
NOR2_X1 U867 ( .A1(n1119), .A2(G952), .ZN(n1126) );
XNOR2_X1 U868 ( .A(n1196), .B(n1207), .ZN(G48) );
NAND2_X1 U869 ( .A1(KEYINPUT1), .A2(G146), .ZN(n1207) );
AND3_X1 U870 ( .A1(n1060), .A2(n1054), .A3(n1208), .ZN(n1196) );
INV_X1 U871 ( .A(n1209), .ZN(n1054) );
XOR2_X1 U872 ( .A(G143), .B(n1210), .Z(G45) );
NOR2_X1 U873 ( .A1(n1211), .A2(n1201), .ZN(n1210) );
NAND3_X1 U874 ( .A1(n1200), .A2(n1212), .A3(n1213), .ZN(n1201) );
NOR3_X1 U875 ( .A1(n1209), .A2(n1214), .A3(n1215), .ZN(n1213) );
XOR2_X1 U876 ( .A(n1069), .B(KEYINPUT9), .Z(n1211) );
NAND2_X1 U877 ( .A1(n1216), .A2(n1217), .ZN(G42) );
NAND2_X1 U878 ( .A1(G140), .A2(n1190), .ZN(n1217) );
XOR2_X1 U879 ( .A(KEYINPUT0), .B(n1218), .Z(n1216) );
NOR2_X1 U880 ( .A1(G140), .A2(n1190), .ZN(n1218) );
NAND3_X1 U881 ( .A1(n1060), .A2(n1219), .A3(n1220), .ZN(n1190) );
XNOR2_X1 U882 ( .A(G137), .B(n1101), .ZN(G39) );
NAND2_X1 U883 ( .A1(n1219), .A2(n1221), .ZN(n1101) );
XOR2_X1 U884 ( .A(G134), .B(n1195), .Z(G36) );
AND3_X1 U885 ( .A1(n1219), .A2(n1059), .A3(n1222), .ZN(n1195) );
NAND2_X1 U886 ( .A1(n1223), .A2(n1224), .ZN(G33) );
NAND2_X1 U887 ( .A1(G131), .A2(n1191), .ZN(n1224) );
XOR2_X1 U888 ( .A(n1225), .B(KEYINPUT24), .Z(n1223) );
OR2_X1 U889 ( .A1(n1191), .A2(G131), .ZN(n1225) );
NAND3_X1 U890 ( .A1(n1060), .A2(n1219), .A3(n1222), .ZN(n1191) );
NOR3_X1 U891 ( .A1(n1209), .A2(n1214), .A3(n1048), .ZN(n1219) );
NAND2_X1 U892 ( .A1(n1080), .A2(n1068), .ZN(n1048) );
INV_X1 U893 ( .A(n1226), .ZN(n1214) );
XOR2_X1 U894 ( .A(n1227), .B(KEYINPUT38), .Z(n1209) );
XOR2_X1 U895 ( .A(G128), .B(n1194), .Z(G30) );
AND3_X1 U896 ( .A1(n1059), .A2(n1228), .A3(n1208), .ZN(n1194) );
AND4_X1 U897 ( .A1(n1229), .A2(n1200), .A3(n1230), .A4(n1226), .ZN(n1208) );
XOR2_X1 U898 ( .A(G101), .B(n1185), .Z(G3) );
NOR3_X1 U899 ( .A1(n1052), .A2(n1187), .A3(n1069), .ZN(n1185) );
INV_X1 U900 ( .A(n1189), .ZN(n1187) );
XOR2_X1 U901 ( .A(G125), .B(n1231), .Z(G27) );
NOR2_X1 U902 ( .A1(n1064), .A2(n1198), .ZN(n1231) );
NAND4_X1 U903 ( .A1(n1220), .A2(n1060), .A3(n1073), .A4(n1226), .ZN(n1198) );
NAND2_X1 U904 ( .A1(n1040), .A2(n1232), .ZN(n1226) );
NAND4_X1 U905 ( .A1(G902), .A2(n1106), .A3(n1233), .A4(n1107), .ZN(n1232) );
INV_X1 U906 ( .A(G900), .ZN(n1107) );
INV_X1 U907 ( .A(n1058), .ZN(n1073) );
XNOR2_X1 U908 ( .A(n1180), .B(n1234), .ZN(G24) );
NOR2_X1 U909 ( .A1(KEYINPUT53), .A2(n1235), .ZN(n1234) );
XNOR2_X1 U910 ( .A(G122), .B(KEYINPUT4), .ZN(n1235) );
NAND4_X1 U911 ( .A1(n1236), .A2(n1071), .A3(n1212), .A4(n1079), .ZN(n1180) );
XNOR2_X1 U912 ( .A(n1237), .B(KEYINPUT18), .ZN(n1212) );
INV_X1 U913 ( .A(n1044), .ZN(n1071) );
NAND2_X1 U914 ( .A1(n1238), .A2(n1239), .ZN(n1044) );
XOR2_X1 U915 ( .A(G119), .B(n1184), .Z(G21) );
AND2_X1 U916 ( .A1(n1236), .A2(n1221), .ZN(n1184) );
AND3_X1 U917 ( .A1(n1229), .A2(n1230), .A3(n1240), .ZN(n1221) );
XOR2_X1 U918 ( .A(G116), .B(n1183), .Z(G18) );
AND3_X1 U919 ( .A1(n1236), .A2(n1059), .A3(n1222), .ZN(n1183) );
NOR2_X1 U920 ( .A1(n1079), .A2(n1237), .ZN(n1059) );
XOR2_X1 U921 ( .A(G113), .B(n1188), .Z(G15) );
AND3_X1 U922 ( .A1(n1060), .A2(n1236), .A3(n1222), .ZN(n1188) );
INV_X1 U923 ( .A(n1069), .ZN(n1222) );
NAND2_X1 U924 ( .A1(n1239), .A2(n1230), .ZN(n1069) );
INV_X1 U925 ( .A(n1238), .ZN(n1230) );
XNOR2_X1 U926 ( .A(KEYINPUT42), .B(n1229), .ZN(n1239) );
NOR3_X1 U927 ( .A1(n1064), .A2(n1241), .A3(n1058), .ZN(n1236) );
NAND2_X1 U928 ( .A1(n1242), .A2(n1056), .ZN(n1058) );
INV_X1 U929 ( .A(n1055), .ZN(n1242) );
AND2_X1 U930 ( .A1(n1237), .A2(n1079), .ZN(n1060) );
INV_X1 U931 ( .A(n1215), .ZN(n1079) );
NAND2_X1 U932 ( .A1(n1243), .A2(n1244), .ZN(G12) );
NAND2_X1 U933 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
XOR2_X1 U934 ( .A(KEYINPUT20), .B(n1247), .Z(n1243) );
NOR2_X1 U935 ( .A1(n1246), .A2(n1245), .ZN(n1247) );
XNOR2_X1 U936 ( .A(KEYINPUT51), .B(G110), .ZN(n1245) );
AND4_X1 U937 ( .A1(n1220), .A2(n1240), .A3(n1248), .A4(n1249), .ZN(n1246) );
OR2_X1 U938 ( .A1(n1189), .A2(KEYINPUT2), .ZN(n1249) );
NOR3_X1 U939 ( .A1(n1064), .A2(n1241), .A3(n1227), .ZN(n1189) );
NAND2_X1 U940 ( .A1(KEYINPUT2), .A2(n1250), .ZN(n1248) );
NAND3_X1 U941 ( .A1(n1228), .A2(n1200), .A3(n1241), .ZN(n1250) );
AND2_X1 U942 ( .A1(n1251), .A2(n1040), .ZN(n1241) );
NAND3_X1 U943 ( .A1(n1233), .A2(n1119), .A3(G952), .ZN(n1040) );
XOR2_X1 U944 ( .A(n1252), .B(KEYINPUT12), .Z(n1251) );
NAND4_X1 U945 ( .A1(G902), .A2(n1106), .A3(n1233), .A4(n1122), .ZN(n1252) );
INV_X1 U946 ( .A(G898), .ZN(n1122) );
NAND2_X1 U947 ( .A1(G237), .A2(G234), .ZN(n1233) );
XOR2_X1 U948 ( .A(G953), .B(KEYINPUT56), .Z(n1106) );
INV_X1 U949 ( .A(n1064), .ZN(n1200) );
NAND2_X1 U950 ( .A1(n1065), .A2(n1068), .ZN(n1064) );
NAND2_X1 U951 ( .A1(G214), .A2(n1253), .ZN(n1068) );
INV_X1 U952 ( .A(n1080), .ZN(n1065) );
XNOR2_X1 U953 ( .A(n1254), .B(n1179), .ZN(n1080) );
NAND2_X1 U954 ( .A1(G210), .A2(n1253), .ZN(n1179) );
NAND2_X1 U955 ( .A1(n1255), .A2(n1256), .ZN(n1253) );
XOR2_X1 U956 ( .A(n1257), .B(KEYINPUT37), .Z(n1255) );
NAND2_X1 U957 ( .A1(n1258), .A2(n1256), .ZN(n1254) );
XOR2_X1 U958 ( .A(n1175), .B(n1259), .Z(n1258) );
NOR3_X1 U959 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1259) );
NOR3_X1 U960 ( .A1(n1205), .A2(n1263), .A3(n1264), .ZN(n1262) );
AND2_X1 U961 ( .A1(n1205), .A2(n1263), .ZN(n1261) );
AND2_X1 U962 ( .A1(n1265), .A2(n1156), .ZN(n1263) );
XNOR2_X1 U963 ( .A(G125), .B(KEYINPUT34), .ZN(n1265) );
INV_X1 U964 ( .A(n1204), .ZN(n1260) );
NAND2_X1 U965 ( .A1(n1264), .A2(n1205), .ZN(n1204) );
NAND2_X1 U966 ( .A1(G224), .A2(n1119), .ZN(n1205) );
NOR2_X1 U967 ( .A1(n1156), .A2(G125), .ZN(n1264) );
NAND2_X1 U968 ( .A1(n1266), .A2(n1267), .ZN(n1175) );
OR2_X1 U969 ( .A1(n1124), .A2(n1125), .ZN(n1267) );
NAND2_X1 U970 ( .A1(n1125), .A2(n1268), .ZN(n1266) );
XNOR2_X1 U971 ( .A(n1124), .B(KEYINPUT35), .ZN(n1268) );
XNOR2_X1 U972 ( .A(n1269), .B(n1270), .ZN(n1124) );
XOR2_X1 U973 ( .A(G113), .B(G110), .Z(n1270) );
XOR2_X1 U974 ( .A(n1271), .B(n1272), .Z(n1269) );
NOR2_X1 U975 ( .A1(KEYINPUT55), .A2(n1273), .ZN(n1272) );
XNOR2_X1 U976 ( .A(n1274), .B(n1275), .ZN(n1125) );
NOR2_X1 U977 ( .A1(KEYINPUT16), .A2(n1276), .ZN(n1275) );
INV_X1 U978 ( .A(G101), .ZN(n1274) );
INV_X1 U979 ( .A(n1227), .ZN(n1228) );
NAND2_X1 U980 ( .A1(n1055), .A2(n1056), .ZN(n1227) );
NAND2_X1 U981 ( .A1(G221), .A2(n1277), .ZN(n1056) );
XNOR2_X1 U982 ( .A(n1278), .B(G469), .ZN(n1055) );
NAND2_X1 U983 ( .A1(n1279), .A2(n1256), .ZN(n1278) );
XOR2_X1 U984 ( .A(n1280), .B(n1281), .Z(n1279) );
INV_X1 U985 ( .A(n1163), .ZN(n1281) );
XOR2_X1 U986 ( .A(n1282), .B(n1283), .Z(n1163) );
XOR2_X1 U987 ( .A(n1276), .B(n1111), .Z(n1283) );
NAND2_X1 U988 ( .A1(n1284), .A2(n1285), .ZN(n1111) );
NAND2_X1 U989 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U990 ( .A(n1288), .B(KEYINPUT57), .Z(n1286) );
NAND2_X1 U991 ( .A1(n1289), .A2(n1290), .ZN(n1284) );
XOR2_X1 U992 ( .A(n1288), .B(KEYINPUT23), .Z(n1290) );
XNOR2_X1 U993 ( .A(G104), .B(G107), .ZN(n1276) );
XOR2_X1 U994 ( .A(n1158), .B(G101), .Z(n1282) );
NOR2_X1 U995 ( .A1(n1291), .A2(n1169), .ZN(n1280) );
AND2_X1 U996 ( .A1(n1173), .A2(n1171), .ZN(n1169) );
NOR2_X1 U997 ( .A1(n1173), .A2(n1171), .ZN(n1291) );
XNOR2_X1 U998 ( .A(G140), .B(G110), .ZN(n1171) );
AND2_X1 U999 ( .A1(G227), .A2(n1119), .ZN(n1173) );
INV_X1 U1000 ( .A(n1052), .ZN(n1240) );
NAND2_X1 U1001 ( .A1(n1237), .A2(n1215), .ZN(n1052) );
XOR2_X1 U1002 ( .A(n1292), .B(G475), .Z(n1215) );
NAND2_X1 U1003 ( .A1(n1138), .A2(n1256), .ZN(n1292) );
XNOR2_X1 U1004 ( .A(n1293), .B(n1294), .ZN(n1138) );
XOR2_X1 U1005 ( .A(n1295), .B(n1271), .Z(n1294) );
NAND2_X1 U1006 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
NAND2_X1 U1007 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
XNOR2_X1 U1008 ( .A(n1300), .B(n1301), .ZN(n1299) );
XOR2_X1 U1009 ( .A(n1302), .B(G131), .Z(n1298) );
XOR2_X1 U1010 ( .A(n1303), .B(KEYINPUT8), .Z(n1296) );
NAND2_X1 U1011 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
XOR2_X1 U1012 ( .A(n1300), .B(n1301), .Z(n1305) );
NAND2_X1 U1013 ( .A1(KEYINPUT54), .A2(n1306), .ZN(n1300) );
XNOR2_X1 U1014 ( .A(G131), .B(n1302), .ZN(n1304) );
NAND2_X1 U1015 ( .A1(n1307), .A2(n1308), .ZN(n1302) );
NAND4_X1 U1016 ( .A1(G214), .A2(G143), .A3(n1257), .A4(n1119), .ZN(n1308) );
NAND2_X1 U1017 ( .A1(n1309), .A2(n1310), .ZN(n1307) );
NAND3_X1 U1018 ( .A1(n1257), .A2(n1119), .A3(G214), .ZN(n1310) );
XOR2_X1 U1019 ( .A(KEYINPUT19), .B(G143), .Z(n1309) );
XNOR2_X1 U1020 ( .A(G104), .B(G113), .ZN(n1293) );
XOR2_X1 U1021 ( .A(n1088), .B(n1311), .Z(n1237) );
NOR2_X1 U1022 ( .A1(KEYINPUT5), .A2(n1135), .ZN(n1311) );
INV_X1 U1023 ( .A(G478), .ZN(n1135) );
NAND2_X1 U1024 ( .A1(n1136), .A2(n1256), .ZN(n1088) );
XOR2_X1 U1025 ( .A(n1312), .B(n1313), .Z(n1136) );
XOR2_X1 U1026 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1027 ( .A(G116), .B(G107), .Z(n1315) );
XOR2_X1 U1028 ( .A(KEYINPUT62), .B(G134), .Z(n1314) );
XOR2_X1 U1029 ( .A(n1316), .B(n1317), .Z(n1312) );
INV_X1 U1030 ( .A(n1271), .ZN(n1317) );
XNOR2_X1 U1031 ( .A(G122), .B(KEYINPUT36), .ZN(n1271) );
XOR2_X1 U1032 ( .A(n1318), .B(n1319), .Z(n1316) );
AND2_X1 U1033 ( .A1(n1320), .A2(G217), .ZN(n1319) );
NAND2_X1 U1034 ( .A1(n1321), .A2(KEYINPUT14), .ZN(n1318) );
XOR2_X1 U1035 ( .A(n1322), .B(n1323), .Z(n1321) );
INV_X1 U1036 ( .A(G143), .ZN(n1322) );
INV_X1 U1037 ( .A(n1070), .ZN(n1220) );
NAND2_X1 U1038 ( .A1(n1238), .A2(n1229), .ZN(n1070) );
XOR2_X1 U1039 ( .A(n1089), .B(KEYINPUT47), .Z(n1229) );
XNOR2_X1 U1040 ( .A(n1324), .B(n1130), .ZN(n1089) );
NAND2_X1 U1041 ( .A1(G217), .A2(n1277), .ZN(n1130) );
NAND2_X1 U1042 ( .A1(G234), .A2(n1256), .ZN(n1277) );
OR2_X1 U1043 ( .A1(n1129), .A2(G902), .ZN(n1324) );
XNOR2_X1 U1044 ( .A(n1325), .B(n1326), .ZN(n1129) );
NOR2_X1 U1045 ( .A1(KEYINPUT41), .A2(n1327), .ZN(n1326) );
XOR2_X1 U1046 ( .A(n1328), .B(G137), .Z(n1327) );
NAND2_X1 U1047 ( .A1(n1320), .A2(G221), .ZN(n1328) );
AND2_X1 U1048 ( .A1(G234), .A2(n1119), .ZN(n1320) );
NAND2_X1 U1049 ( .A1(n1329), .A2(n1330), .ZN(n1325) );
NAND2_X1 U1050 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U1051 ( .A(KEYINPUT29), .B(n1333), .Z(n1329) );
NOR2_X1 U1052 ( .A1(n1332), .A2(n1331), .ZN(n1333) );
XNOR2_X1 U1053 ( .A(G110), .B(n1334), .ZN(n1331) );
NAND3_X1 U1054 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1334) );
NAND2_X1 U1055 ( .A1(n1323), .A2(n1338), .ZN(n1337) );
NAND3_X1 U1056 ( .A1(n1339), .A2(n1340), .A3(n1341), .ZN(n1338) );
NAND2_X1 U1057 ( .A1(KEYINPUT40), .A2(n1342), .ZN(n1341) );
NAND2_X1 U1058 ( .A1(KEYINPUT46), .A2(n1343), .ZN(n1340) );
NAND2_X1 U1059 ( .A1(n1344), .A2(n1345), .ZN(n1339) );
INV_X1 U1060 ( .A(KEYINPUT46), .ZN(n1345) );
NAND2_X1 U1061 ( .A1(n1343), .A2(n1346), .ZN(n1344) );
NAND2_X1 U1062 ( .A1(KEYINPUT26), .A2(n1347), .ZN(n1346) );
NAND4_X1 U1063 ( .A1(n1343), .A2(n1342), .A3(n1288), .A4(n1347), .ZN(n1336) );
INV_X1 U1064 ( .A(KEYINPUT40), .ZN(n1347) );
INV_X1 U1065 ( .A(KEYINPUT26), .ZN(n1342) );
NAND2_X1 U1066 ( .A1(KEYINPUT40), .A2(n1348), .ZN(n1335) );
NAND2_X1 U1067 ( .A1(n1343), .A2(n1349), .ZN(n1348) );
NAND2_X1 U1068 ( .A1(KEYINPUT26), .A2(n1288), .ZN(n1349) );
XNOR2_X1 U1069 ( .A(n1301), .B(n1306), .ZN(n1332) );
XNOR2_X1 U1070 ( .A(n1110), .B(KEYINPUT63), .ZN(n1306) );
XNOR2_X1 U1071 ( .A(G140), .B(G125), .ZN(n1110) );
XNOR2_X1 U1072 ( .A(G146), .B(KEYINPUT22), .ZN(n1301) );
XOR2_X1 U1073 ( .A(n1086), .B(G472), .Z(n1238) );
NAND3_X1 U1074 ( .A1(n1350), .A2(n1256), .A3(n1351), .ZN(n1086) );
NAND2_X1 U1075 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
XOR2_X1 U1076 ( .A(KEYINPUT30), .B(n1354), .Z(n1353) );
XOR2_X1 U1077 ( .A(KEYINPUT13), .B(n1156), .Z(n1352) );
INV_X1 U1078 ( .A(G902), .ZN(n1256) );
NAND2_X1 U1079 ( .A1(n1355), .A2(n1356), .ZN(n1350) );
XNOR2_X1 U1080 ( .A(n1354), .B(KEYINPUT33), .ZN(n1356) );
XOR2_X1 U1081 ( .A(n1150), .B(n1159), .Z(n1354) );
INV_X1 U1082 ( .A(n1158), .ZN(n1159) );
XNOR2_X1 U1083 ( .A(n1357), .B(n1113), .ZN(n1158) );
XNOR2_X1 U1084 ( .A(G134), .B(G137), .ZN(n1113) );
XNOR2_X1 U1085 ( .A(KEYINPUT25), .B(n1358), .ZN(n1357) );
NOR2_X1 U1086 ( .A1(G131), .A2(KEYINPUT32), .ZN(n1358) );
XNOR2_X1 U1087 ( .A(n1359), .B(n1360), .ZN(n1150) );
XOR2_X1 U1088 ( .A(G113), .B(G101), .Z(n1360) );
XNOR2_X1 U1089 ( .A(n1361), .B(n1273), .ZN(n1359) );
XOR2_X1 U1090 ( .A(G116), .B(n1343), .Z(n1273) );
INV_X1 U1091 ( .A(G119), .ZN(n1343) );
NAND3_X1 U1092 ( .A1(n1257), .A2(n1119), .A3(G210), .ZN(n1361) );
INV_X1 U1093 ( .A(G953), .ZN(n1119) );
INV_X1 U1094 ( .A(G237), .ZN(n1257) );
XOR2_X1 U1095 ( .A(KEYINPUT13), .B(n1155), .Z(n1355) );
INV_X1 U1096 ( .A(n1156), .ZN(n1155) );
XNOR2_X1 U1097 ( .A(n1287), .B(n1323), .ZN(n1156) );
INV_X1 U1098 ( .A(n1288), .ZN(n1323) );
XNOR2_X1 U1099 ( .A(G128), .B(KEYINPUT49), .ZN(n1288) );
INV_X1 U1100 ( .A(n1289), .ZN(n1287) );
XOR2_X1 U1101 ( .A(G146), .B(G143), .Z(n1289) );
endmodule


