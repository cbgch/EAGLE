//Key = 0100010100110011101001011101110010011101101011000000011111010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327;

XOR2_X1 U733 ( .A(G107), .B(n1012), .Z(G9) );
NOR2_X1 U734 ( .A1(n1013), .A2(n1014), .ZN(G75) );
NOR3_X1 U735 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NAND3_X1 U736 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1015) );
NAND2_X1 U737 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U738 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND3_X1 U739 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1024) );
NAND2_X1 U740 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
OR3_X1 U741 ( .A1(n1030), .A2(KEYINPUT21), .A3(n1031), .ZN(n1028) );
NAND3_X1 U742 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1025) );
NAND2_X1 U743 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NAND2_X1 U744 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND4_X1 U745 ( .A1(n1039), .A2(G221), .A3(n1040), .A4(n1041), .ZN(n1038) );
INV_X1 U746 ( .A(KEYINPUT30), .ZN(n1041) );
NAND2_X1 U747 ( .A1(KEYINPUT21), .A2(n1042), .ZN(n1037) );
NAND2_X1 U748 ( .A1(n1043), .A2(n1044), .ZN(n1032) );
NAND2_X1 U749 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND3_X1 U750 ( .A1(n1043), .A2(n1047), .A3(n1035), .ZN(n1023) );
NAND2_X1 U751 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U752 ( .A1(n1034), .A2(n1050), .ZN(n1049) );
NAND2_X1 U753 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U754 ( .A1(n1027), .A2(n1053), .ZN(n1048) );
NAND3_X1 U755 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NAND2_X1 U756 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U757 ( .A1(KEYINPUT30), .A2(n1034), .ZN(n1054) );
INV_X1 U758 ( .A(n1059), .ZN(n1021) );
NOR3_X1 U759 ( .A1(n1060), .A2(G953), .A3(G952), .ZN(n1013) );
INV_X1 U760 ( .A(n1018), .ZN(n1060) );
NAND4_X1 U761 ( .A1(n1057), .A2(n1027), .A3(n1043), .A4(n1061), .ZN(n1018) );
NOR3_X1 U762 ( .A1(n1062), .A2(n1058), .A3(n1063), .ZN(n1061) );
XOR2_X1 U763 ( .A(n1064), .B(n1065), .Z(n1063) );
NOR2_X1 U764 ( .A1(G478), .A2(KEYINPUT58), .ZN(n1065) );
XOR2_X1 U765 ( .A(n1066), .B(n1067), .Z(G72) );
NOR2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
XOR2_X1 U767 ( .A(KEYINPUT3), .B(n1019), .Z(n1069) );
NOR2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
XNOR2_X1 U769 ( .A(G227), .B(KEYINPUT9), .ZN(n1070) );
NAND2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1066) );
NAND2_X1 U771 ( .A1(n1074), .A2(n1019), .ZN(n1073) );
XOR2_X1 U772 ( .A(n1075), .B(n1076), .Z(n1074) );
NAND2_X1 U773 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NAND2_X1 U774 ( .A1(n1017), .A2(n1079), .ZN(n1078) );
INV_X1 U775 ( .A(KEYINPUT51), .ZN(n1079) );
NAND2_X1 U776 ( .A1(KEYINPUT51), .A2(n1080), .ZN(n1077) );
NAND2_X1 U777 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND3_X1 U778 ( .A1(n1083), .A2(n1076), .A3(G953), .ZN(n1072) );
XNOR2_X1 U779 ( .A(n1084), .B(n1085), .ZN(n1076) );
XNOR2_X1 U780 ( .A(G131), .B(n1086), .ZN(n1085) );
XNOR2_X1 U781 ( .A(n1087), .B(n1088), .ZN(n1084) );
XOR2_X1 U782 ( .A(KEYINPUT31), .B(G900), .Z(n1083) );
XOR2_X1 U783 ( .A(n1089), .B(n1090), .Z(G69) );
XOR2_X1 U784 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U785 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U786 ( .A(KEYINPUT20), .B(G953), .Z(n1094) );
NAND2_X1 U787 ( .A1(n1095), .A2(n1096), .ZN(n1091) );
NAND2_X1 U788 ( .A1(G898), .A2(G224), .ZN(n1096) );
XOR2_X1 U789 ( .A(KEYINPUT3), .B(G953), .Z(n1095) );
NAND2_X1 U790 ( .A1(n1097), .A2(n1098), .ZN(n1089) );
NAND2_X1 U791 ( .A1(G953), .A2(n1099), .ZN(n1098) );
XNOR2_X1 U792 ( .A(n1100), .B(n1101), .ZN(n1097) );
NOR2_X1 U793 ( .A1(n1102), .A2(n1103), .ZN(G66) );
XOR2_X1 U794 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U795 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NOR2_X1 U796 ( .A1(n1102), .A2(n1108), .ZN(G63) );
NOR3_X1 U797 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1108) );
NOR3_X1 U798 ( .A1(n1112), .A2(n1113), .A3(n1107), .ZN(n1111) );
NOR2_X1 U799 ( .A1(n1114), .A2(n1115), .ZN(n1110) );
NOR2_X1 U800 ( .A1(n1116), .A2(n1113), .ZN(n1114) );
NOR2_X1 U801 ( .A1(n1102), .A2(n1117), .ZN(G60) );
XNOR2_X1 U802 ( .A(n1118), .B(n1119), .ZN(n1117) );
NOR3_X1 U803 ( .A1(n1107), .A2(KEYINPUT4), .A3(n1120), .ZN(n1119) );
INV_X1 U804 ( .A(G475), .ZN(n1120) );
XNOR2_X1 U805 ( .A(n1121), .B(n1122), .ZN(G6) );
NOR2_X1 U806 ( .A1(KEYINPUT52), .A2(n1123), .ZN(n1122) );
NOR2_X1 U807 ( .A1(n1124), .A2(n1125), .ZN(G57) );
XOR2_X1 U808 ( .A(n1126), .B(n1127), .Z(n1125) );
XNOR2_X1 U809 ( .A(n1128), .B(n1129), .ZN(n1127) );
XOR2_X1 U810 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U811 ( .A1(KEYINPUT57), .A2(n1132), .ZN(n1130) );
XOR2_X1 U812 ( .A(n1133), .B(n1134), .Z(n1126) );
XOR2_X1 U813 ( .A(KEYINPUT2), .B(G101), .Z(n1134) );
AND2_X1 U814 ( .A1(G472), .A2(n1135), .ZN(n1133) );
NOR2_X1 U815 ( .A1(G952), .A2(n1136), .ZN(n1124) );
XOR2_X1 U816 ( .A(KEYINPUT5), .B(G953), .Z(n1136) );
NOR2_X1 U817 ( .A1(n1102), .A2(n1137), .ZN(G54) );
XOR2_X1 U818 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U819 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U820 ( .A1(KEYINPUT46), .A2(n1142), .ZN(n1141) );
XOR2_X1 U821 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U822 ( .A1(KEYINPUT35), .A2(n1145), .ZN(n1143) );
NAND2_X1 U823 ( .A1(n1135), .A2(G469), .ZN(n1140) );
NOR2_X1 U824 ( .A1(n1102), .A2(n1146), .ZN(G51) );
XOR2_X1 U825 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U826 ( .A1(n1149), .A2(n1107), .ZN(n1147) );
INV_X1 U827 ( .A(n1135), .ZN(n1107) );
NOR2_X1 U828 ( .A1(n1150), .A2(n1116), .ZN(n1135) );
AND2_X1 U829 ( .A1(n1151), .A2(n1093), .ZN(n1116) );
INV_X1 U830 ( .A(n1016), .ZN(n1093) );
NAND4_X1 U831 ( .A1(n1121), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1016) );
NOR4_X1 U832 ( .A1(n1012), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1154) );
NOR2_X1 U833 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NOR2_X1 U834 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
XOR2_X1 U835 ( .A(n1052), .B(KEYINPUT14), .Z(n1161) );
NOR2_X1 U836 ( .A1(n1051), .A2(n1162), .ZN(n1160) );
NOR3_X1 U837 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1156) );
NOR4_X1 U838 ( .A1(n1166), .A2(n1051), .A3(n1030), .A4(n1031), .ZN(n1155) );
INV_X1 U839 ( .A(n1035), .ZN(n1031) );
INV_X1 U840 ( .A(n1042), .ZN(n1030) );
NAND3_X1 U841 ( .A1(n1167), .A2(n1162), .A3(n1055), .ZN(n1166) );
INV_X1 U842 ( .A(KEYINPUT7), .ZN(n1162) );
AND2_X1 U843 ( .A1(n1168), .A2(n1169), .ZN(n1012) );
NOR2_X1 U844 ( .A1(n1170), .A2(n1171), .ZN(n1153) );
NAND2_X1 U845 ( .A1(n1172), .A2(n1169), .ZN(n1121) );
AND4_X1 U846 ( .A1(n1042), .A2(n1173), .A3(n1027), .A4(n1167), .ZN(n1169) );
XOR2_X1 U847 ( .A(n1017), .B(KEYINPUT29), .Z(n1151) );
NAND4_X1 U848 ( .A1(n1174), .A2(n1082), .A3(n1175), .A4(n1176), .ZN(n1017) );
NOR2_X1 U849 ( .A1(n1177), .A2(n1081), .ZN(n1176) );
NAND4_X1 U850 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1081) );
NAND4_X1 U851 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1042), .ZN(n1178) );
NOR2_X1 U852 ( .A1(n1185), .A2(n1055), .ZN(n1184) );
XOR2_X1 U853 ( .A(n1186), .B(KEYINPUT59), .Z(n1185) );
INV_X1 U854 ( .A(n1165), .ZN(n1183) );
NOR3_X1 U855 ( .A1(n1187), .A2(n1046), .A3(n1029), .ZN(n1177) );
OR3_X1 U856 ( .A1(n1045), .A2(n1029), .A3(n1187), .ZN(n1082) );
INV_X1 U857 ( .A(n1034), .ZN(n1029) );
NOR2_X1 U858 ( .A1(n1019), .A2(G952), .ZN(n1102) );
NAND2_X1 U859 ( .A1(n1188), .A2(n1189), .ZN(G48) );
NAND2_X1 U860 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
INV_X1 U861 ( .A(G146), .ZN(n1191) );
XNOR2_X1 U862 ( .A(KEYINPUT43), .B(n1179), .ZN(n1190) );
NAND2_X1 U863 ( .A1(G146), .A2(n1192), .ZN(n1188) );
XOR2_X1 U864 ( .A(n1179), .B(KEYINPUT47), .Z(n1192) );
NAND3_X1 U865 ( .A1(n1193), .A2(n1173), .A3(n1172), .ZN(n1179) );
XOR2_X1 U866 ( .A(G143), .B(n1194), .Z(G45) );
NOR4_X1 U867 ( .A1(KEYINPUT60), .A2(n1055), .A3(n1165), .A4(n1187), .ZN(n1194) );
INV_X1 U868 ( .A(n1173), .ZN(n1055) );
XNOR2_X1 U869 ( .A(G140), .B(n1180), .ZN(G42) );
NAND3_X1 U870 ( .A1(n1034), .A2(n1042), .A3(n1195), .ZN(n1180) );
XNOR2_X1 U871 ( .A(G137), .B(n1181), .ZN(G39) );
NAND3_X1 U872 ( .A1(n1193), .A2(n1034), .A3(n1035), .ZN(n1181) );
XNOR2_X1 U873 ( .A(G134), .B(n1196), .ZN(G36) );
NAND4_X1 U874 ( .A1(n1034), .A2(n1168), .A3(n1197), .A4(n1198), .ZN(n1196) );
NAND2_X1 U875 ( .A1(n1187), .A2(n1199), .ZN(n1198) );
INV_X1 U876 ( .A(KEYINPUT8), .ZN(n1199) );
NAND2_X1 U877 ( .A1(KEYINPUT8), .A2(n1200), .ZN(n1197) );
NAND3_X1 U878 ( .A1(n1186), .A2(n1052), .A3(n1042), .ZN(n1200) );
XOR2_X1 U879 ( .A(G131), .B(n1201), .Z(G33) );
NOR4_X1 U880 ( .A1(KEYINPUT38), .A2(n1045), .A3(n1187), .A4(n1202), .ZN(n1201) );
XOR2_X1 U881 ( .A(KEYINPUT56), .B(n1034), .Z(n1202) );
NOR2_X1 U882 ( .A1(n1203), .A2(n1204), .ZN(n1034) );
XOR2_X1 U883 ( .A(KEYINPUT37), .B(n1057), .Z(n1203) );
NAND3_X1 U884 ( .A1(n1042), .A2(n1186), .A3(n1182), .ZN(n1187) );
XNOR2_X1 U885 ( .A(G128), .B(n1175), .ZN(G30) );
NAND3_X1 U886 ( .A1(n1168), .A2(n1173), .A3(n1193), .ZN(n1175) );
AND4_X1 U887 ( .A1(n1042), .A2(n1205), .A3(n1206), .A4(n1186), .ZN(n1193) );
NAND3_X1 U888 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(G3) );
NAND2_X1 U889 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND3_X1 U890 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1211) );
NAND2_X1 U891 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND2_X1 U892 ( .A1(n1217), .A2(n1218), .ZN(n1213) );
INV_X1 U893 ( .A(KEYINPUT50), .ZN(n1218) );
NAND2_X1 U894 ( .A1(n1219), .A2(n1220), .ZN(n1217) );
NAND2_X1 U895 ( .A1(KEYINPUT44), .A2(KEYINPUT13), .ZN(n1220) );
NAND2_X1 U896 ( .A1(KEYINPUT50), .A2(n1219), .ZN(n1212) );
INV_X1 U897 ( .A(n1221), .ZN(n1210) );
NAND4_X1 U898 ( .A1(n1221), .A2(n1215), .A3(n1219), .A4(KEYINPUT44), .ZN(n1208) );
INV_X1 U899 ( .A(KEYINPUT13), .ZN(n1215) );
NAND2_X1 U900 ( .A1(n1222), .A2(n1216), .ZN(n1207) );
INV_X1 U901 ( .A(KEYINPUT44), .ZN(n1216) );
NAND2_X1 U902 ( .A1(n1219), .A2(n1223), .ZN(n1222) );
NAND2_X1 U903 ( .A1(KEYINPUT13), .A2(n1221), .ZN(n1223) );
NAND2_X1 U904 ( .A1(n1224), .A2(n1182), .ZN(n1221) );
INV_X1 U905 ( .A(n1052), .ZN(n1182) );
XOR2_X1 U906 ( .A(n1225), .B(KEYINPUT40), .Z(n1219) );
XOR2_X1 U907 ( .A(n1174), .B(n1226), .Z(G27) );
NAND2_X1 U908 ( .A1(KEYINPUT42), .A2(G125), .ZN(n1226) );
NAND3_X1 U909 ( .A1(n1043), .A2(n1173), .A3(n1195), .ZN(n1174) );
AND3_X1 U910 ( .A1(n1172), .A2(n1186), .A3(n1227), .ZN(n1195) );
NAND2_X1 U911 ( .A1(n1059), .A2(n1228), .ZN(n1186) );
NAND4_X1 U912 ( .A1(G953), .A2(G902), .A3(n1229), .A4(n1071), .ZN(n1228) );
INV_X1 U913 ( .A(G900), .ZN(n1071) );
INV_X1 U914 ( .A(n1045), .ZN(n1172) );
XNOR2_X1 U915 ( .A(G122), .B(n1230), .ZN(G24) );
NAND3_X1 U916 ( .A1(n1231), .A2(n1027), .A3(n1232), .ZN(n1230) );
XOR2_X1 U917 ( .A(n1165), .B(KEYINPUT32), .Z(n1232) );
NAND2_X1 U918 ( .A1(n1062), .A2(n1233), .ZN(n1165) );
INV_X1 U919 ( .A(n1164), .ZN(n1027) );
NAND2_X1 U920 ( .A1(n1234), .A2(n1235), .ZN(n1164) );
XOR2_X1 U921 ( .A(n1236), .B(n1237), .Z(G21) );
NAND2_X1 U922 ( .A1(KEYINPUT27), .A2(n1238), .ZN(n1237) );
INV_X1 U923 ( .A(n1152), .ZN(n1238) );
NAND4_X1 U924 ( .A1(n1231), .A2(n1035), .A3(n1205), .A4(n1206), .ZN(n1152) );
INV_X1 U925 ( .A(n1163), .ZN(n1231) );
XOR2_X1 U926 ( .A(G116), .B(n1171), .Z(G18) );
NOR3_X1 U927 ( .A1(n1052), .A2(n1046), .A3(n1163), .ZN(n1171) );
INV_X1 U928 ( .A(n1168), .ZN(n1046) );
NOR2_X1 U929 ( .A1(n1062), .A2(n1239), .ZN(n1168) );
XOR2_X1 U930 ( .A(G113), .B(n1170), .Z(G15) );
NOR3_X1 U931 ( .A1(n1052), .A2(n1045), .A3(n1163), .ZN(n1170) );
NAND3_X1 U932 ( .A1(n1173), .A2(n1167), .A3(n1043), .ZN(n1163) );
AND2_X1 U933 ( .A1(n1039), .A2(n1240), .ZN(n1043) );
NAND2_X1 U934 ( .A1(G221), .A2(n1040), .ZN(n1240) );
NAND2_X1 U935 ( .A1(n1239), .A2(n1062), .ZN(n1045) );
INV_X1 U936 ( .A(n1233), .ZN(n1239) );
NAND2_X1 U937 ( .A1(n1234), .A2(n1206), .ZN(n1052) );
INV_X1 U938 ( .A(n1235), .ZN(n1206) );
XNOR2_X1 U939 ( .A(G110), .B(n1241), .ZN(G12) );
NAND3_X1 U940 ( .A1(n1224), .A2(n1227), .A3(KEYINPUT10), .ZN(n1241) );
INV_X1 U941 ( .A(n1051), .ZN(n1227) );
NAND2_X1 U942 ( .A1(n1235), .A2(n1205), .ZN(n1051) );
XNOR2_X1 U943 ( .A(n1234), .B(KEYINPUT41), .ZN(n1205) );
XNOR2_X1 U944 ( .A(n1242), .B(n1106), .ZN(n1234) );
NAND2_X1 U945 ( .A1(G217), .A2(n1040), .ZN(n1106) );
OR2_X1 U946 ( .A1(n1105), .A2(G902), .ZN(n1242) );
XNOR2_X1 U947 ( .A(n1243), .B(n1244), .ZN(n1105) );
XOR2_X1 U948 ( .A(n1245), .B(n1246), .Z(n1243) );
XOR2_X1 U949 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U950 ( .A(KEYINPUT11), .B(G137), .Z(n1248) );
XOR2_X1 U951 ( .A(KEYINPUT49), .B(KEYINPUT12), .Z(n1247) );
XOR2_X1 U952 ( .A(n1249), .B(n1250), .Z(n1245) );
XOR2_X1 U953 ( .A(G128), .B(G119), .Z(n1250) );
XOR2_X1 U954 ( .A(n1251), .B(G110), .Z(n1249) );
NAND2_X1 U955 ( .A1(G221), .A2(n1252), .ZN(n1251) );
XOR2_X1 U956 ( .A(n1253), .B(G472), .Z(n1235) );
NAND2_X1 U957 ( .A1(n1254), .A2(n1150), .ZN(n1253) );
XOR2_X1 U958 ( .A(n1255), .B(n1256), .Z(n1254) );
XNOR2_X1 U959 ( .A(n1132), .B(n1128), .ZN(n1256) );
XNOR2_X1 U960 ( .A(n1236), .B(n1257), .ZN(n1128) );
XOR2_X1 U961 ( .A(n1258), .B(n1131), .Z(n1255) );
XNOR2_X1 U962 ( .A(n1259), .B(n1260), .ZN(n1131) );
AND3_X1 U963 ( .A1(G210), .A2(n1019), .A3(n1261), .ZN(n1260) );
NAND2_X1 U964 ( .A1(KEYINPUT23), .A2(n1225), .ZN(n1258) );
INV_X1 U965 ( .A(n1159), .ZN(n1224) );
NAND4_X1 U966 ( .A1(n1035), .A2(n1042), .A3(n1173), .A4(n1167), .ZN(n1159) );
NAND2_X1 U967 ( .A1(n1059), .A2(n1262), .ZN(n1167) );
NAND4_X1 U968 ( .A1(G953), .A2(G902), .A3(n1229), .A4(n1099), .ZN(n1262) );
INV_X1 U969 ( .A(G898), .ZN(n1099) );
NAND3_X1 U970 ( .A1(n1229), .A2(n1019), .A3(G952), .ZN(n1059) );
NAND2_X1 U971 ( .A1(G237), .A2(n1263), .ZN(n1229) );
NOR2_X1 U972 ( .A1(n1057), .A2(n1204), .ZN(n1173) );
XNOR2_X1 U973 ( .A(n1058), .B(KEYINPUT55), .ZN(n1204) );
AND2_X1 U974 ( .A1(G214), .A2(n1264), .ZN(n1058) );
XNOR2_X1 U975 ( .A(n1265), .B(n1149), .ZN(n1057) );
NAND2_X1 U976 ( .A1(G210), .A2(n1264), .ZN(n1149) );
NAND2_X1 U977 ( .A1(n1261), .A2(n1150), .ZN(n1264) );
OR2_X1 U978 ( .A1(n1148), .A2(G902), .ZN(n1265) );
XNOR2_X1 U979 ( .A(n1266), .B(n1267), .ZN(n1148) );
XOR2_X1 U980 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U981 ( .A(n1259), .B(G125), .Z(n1269) );
NAND2_X1 U982 ( .A1(n1270), .A2(n1271), .ZN(n1259) );
NAND2_X1 U983 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
XOR2_X1 U984 ( .A(KEYINPUT18), .B(n1274), .Z(n1270) );
NOR2_X1 U985 ( .A1(n1272), .A2(n1273), .ZN(n1274) );
NAND2_X1 U986 ( .A1(G224), .A2(n1019), .ZN(n1268) );
XOR2_X1 U987 ( .A(n1275), .B(n1101), .Z(n1266) );
XOR2_X1 U988 ( .A(G110), .B(G122), .Z(n1101) );
NAND2_X1 U989 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND3_X1 U990 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1277) );
INV_X1 U991 ( .A(KEYINPUT39), .ZN(n1280) );
NAND2_X1 U992 ( .A1(n1100), .A2(KEYINPUT39), .ZN(n1276) );
XOR2_X1 U993 ( .A(n1278), .B(n1279), .Z(n1100) );
XNOR2_X1 U994 ( .A(n1281), .B(n1257), .ZN(n1279) );
XNOR2_X1 U995 ( .A(n1282), .B(n1283), .ZN(n1257) );
XNOR2_X1 U996 ( .A(G116), .B(KEYINPUT15), .ZN(n1282) );
XOR2_X1 U997 ( .A(n1284), .B(KEYINPUT48), .Z(n1281) );
NAND2_X1 U998 ( .A1(KEYINPUT25), .A2(n1236), .ZN(n1284) );
INV_X1 U999 ( .A(G119), .ZN(n1236) );
XOR2_X1 U1000 ( .A(n1285), .B(n1286), .Z(n1278) );
NOR2_X1 U1001 ( .A1(KEYINPUT0), .A2(n1287), .ZN(n1286) );
XOR2_X1 U1002 ( .A(n1288), .B(G107), .Z(n1287) );
NAND2_X1 U1003 ( .A1(KEYINPUT1), .A2(G104), .ZN(n1288) );
NOR2_X1 U1004 ( .A1(n1039), .A2(n1289), .ZN(n1042) );
AND2_X1 U1005 ( .A1(G221), .A2(n1040), .ZN(n1289) );
NAND2_X1 U1006 ( .A1(n1263), .A2(n1150), .ZN(n1040) );
XNOR2_X1 U1007 ( .A(G234), .B(KEYINPUT53), .ZN(n1263) );
XOR2_X1 U1008 ( .A(n1290), .B(G469), .Z(n1039) );
NAND2_X1 U1009 ( .A1(n1291), .A2(n1150), .ZN(n1290) );
XOR2_X1 U1010 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U1011 ( .A(n1294), .B(n1145), .Z(n1293) );
XOR2_X1 U1012 ( .A(n1088), .B(KEYINPUT17), .Z(n1145) );
XOR2_X1 U1013 ( .A(n1272), .B(n1273), .Z(n1088) );
XOR2_X1 U1014 ( .A(G143), .B(G146), .Z(n1273) );
XOR2_X1 U1015 ( .A(G128), .B(KEYINPUT34), .Z(n1272) );
INV_X1 U1016 ( .A(n1138), .ZN(n1294) );
XOR2_X1 U1017 ( .A(n1295), .B(n1296), .Z(n1138) );
XOR2_X1 U1018 ( .A(G140), .B(G110), .Z(n1296) );
NAND2_X1 U1019 ( .A1(G227), .A2(n1019), .ZN(n1295) );
INV_X1 U1020 ( .A(n1144), .ZN(n1292) );
XOR2_X1 U1021 ( .A(n1297), .B(n1298), .Z(n1144) );
XOR2_X1 U1022 ( .A(G107), .B(G104), .Z(n1298) );
XNOR2_X1 U1023 ( .A(n1132), .B(n1285), .ZN(n1297) );
XNOR2_X1 U1024 ( .A(n1225), .B(KEYINPUT19), .ZN(n1285) );
INV_X1 U1025 ( .A(G101), .ZN(n1225) );
XNOR2_X1 U1026 ( .A(n1299), .B(G131), .ZN(n1132) );
NAND2_X1 U1027 ( .A1(KEYINPUT16), .A2(n1086), .ZN(n1299) );
XNOR2_X1 U1028 ( .A(G137), .B(n1300), .ZN(n1086) );
NOR2_X1 U1029 ( .A1(n1233), .A2(n1062), .ZN(n1035) );
XNOR2_X1 U1030 ( .A(n1301), .B(G475), .ZN(n1062) );
NAND2_X1 U1031 ( .A1(n1302), .A2(n1118), .ZN(n1301) );
XNOR2_X1 U1032 ( .A(n1303), .B(n1304), .ZN(n1118) );
XOR2_X1 U1033 ( .A(n1244), .B(n1305), .Z(n1304) );
XNOR2_X1 U1034 ( .A(n1306), .B(n1307), .ZN(n1305) );
NOR2_X1 U1035 ( .A1(KEYINPUT26), .A2(n1308), .ZN(n1307) );
XOR2_X1 U1036 ( .A(G122), .B(n1283), .Z(n1308) );
XOR2_X1 U1037 ( .A(G113), .B(KEYINPUT6), .Z(n1283) );
NAND3_X1 U1038 ( .A1(n1309), .A2(n1310), .A3(KEYINPUT61), .ZN(n1306) );
NAND2_X1 U1039 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NAND3_X1 U1040 ( .A1(n1261), .A2(n1019), .A3(G214), .ZN(n1312) );
XOR2_X1 U1041 ( .A(n1313), .B(KEYINPUT28), .Z(n1311) );
INV_X1 U1042 ( .A(G143), .ZN(n1313) );
NAND4_X1 U1043 ( .A1(G214), .A2(n1314), .A3(n1261), .A4(n1019), .ZN(n1309) );
INV_X1 U1044 ( .A(G237), .ZN(n1261) );
XOR2_X1 U1045 ( .A(KEYINPUT36), .B(G143), .Z(n1314) );
XOR2_X1 U1046 ( .A(G146), .B(n1087), .Z(n1244) );
XOR2_X1 U1047 ( .A(G125), .B(G140), .Z(n1087) );
XOR2_X1 U1048 ( .A(n1123), .B(n1315), .Z(n1303) );
XOR2_X1 U1049 ( .A(KEYINPUT22), .B(G131), .Z(n1315) );
INV_X1 U1050 ( .A(G104), .ZN(n1123) );
XOR2_X1 U1051 ( .A(KEYINPUT24), .B(G902), .Z(n1302) );
NAND2_X1 U1052 ( .A1(n1316), .A2(n1317), .ZN(n1233) );
NAND2_X1 U1053 ( .A1(G478), .A2(n1064), .ZN(n1317) );
XOR2_X1 U1054 ( .A(n1318), .B(KEYINPUT33), .Z(n1316) );
NAND2_X1 U1055 ( .A1(n1109), .A2(n1113), .ZN(n1318) );
INV_X1 U1056 ( .A(G478), .ZN(n1113) );
INV_X1 U1057 ( .A(n1064), .ZN(n1109) );
NAND2_X1 U1058 ( .A1(n1112), .A2(n1150), .ZN(n1064) );
INV_X1 U1059 ( .A(G902), .ZN(n1150) );
INV_X1 U1060 ( .A(n1115), .ZN(n1112) );
XOR2_X1 U1061 ( .A(n1319), .B(n1320), .Z(n1115) );
XNOR2_X1 U1062 ( .A(n1321), .B(n1300), .ZN(n1320) );
XOR2_X1 U1063 ( .A(G134), .B(KEYINPUT63), .Z(n1300) );
NAND2_X1 U1064 ( .A1(G217), .A2(n1252), .ZN(n1321) );
AND2_X1 U1065 ( .A1(G234), .A2(n1019), .ZN(n1252) );
INV_X1 U1066 ( .A(G953), .ZN(n1019) );
XOR2_X1 U1067 ( .A(n1322), .B(n1323), .Z(n1319) );
XOR2_X1 U1068 ( .A(G143), .B(G128), .Z(n1323) );
NAND2_X1 U1069 ( .A1(KEYINPUT54), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1070 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1071 ( .A(G122), .B(G107), .Z(n1326) );
NOR2_X1 U1072 ( .A1(KEYINPUT62), .A2(n1327), .ZN(n1325) );
XNOR2_X1 U1073 ( .A(G116), .B(KEYINPUT45), .ZN(n1327) );
endmodule


