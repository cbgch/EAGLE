//Key = 1000101111111011000100100101010111111010000010000000100000010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297;

XNOR2_X1 U722 ( .A(G107), .B(n984), .ZN(G9) );
NOR2_X1 U723 ( .A1(n985), .A2(KEYINPUT50), .ZN(n984) );
NAND4_X1 U724 ( .A1(n986), .A2(n987), .A3(n988), .A4(n989), .ZN(G75) );
NAND4_X1 U725 ( .A1(n990), .A2(n991), .A3(n992), .A4(n993), .ZN(n988) );
NOR4_X1 U726 ( .A1(n994), .A2(n995), .A3(n996), .A4(n997), .ZN(n993) );
XNOR2_X1 U727 ( .A(n998), .B(KEYINPUT52), .ZN(n995) );
XNOR2_X1 U728 ( .A(G469), .B(n999), .ZN(n994) );
NOR2_X1 U729 ( .A1(n1000), .A2(KEYINPUT54), .ZN(n999) );
NOR3_X1 U730 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n992) );
NAND2_X1 U731 ( .A1(n1004), .A2(n1005), .ZN(n987) );
NAND2_X1 U732 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NAND3_X1 U733 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1007) );
NAND2_X1 U734 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NAND2_X1 U735 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U736 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U737 ( .A1(n1017), .A2(n1018), .ZN(n1011) );
NAND2_X1 U738 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
XNOR2_X1 U739 ( .A(n1021), .B(KEYINPUT62), .ZN(n1019) );
NAND3_X1 U740 ( .A1(n1017), .A2(n1022), .A3(n1013), .ZN(n1006) );
NAND3_X1 U741 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NAND2_X1 U742 ( .A1(n1008), .A2(n1026), .ZN(n1025) );
NAND2_X1 U743 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U744 ( .A1(n1029), .A2(n1003), .ZN(n1028) );
NAND3_X1 U745 ( .A1(n1030), .A2(n1010), .A3(n1031), .ZN(n1023) );
INV_X1 U746 ( .A(n1032), .ZN(n1004) );
XOR2_X1 U747 ( .A(n1033), .B(n1034), .Z(G72) );
XOR2_X1 U748 ( .A(n1035), .B(n1036), .Z(n1034) );
NOR3_X1 U749 ( .A1(n1037), .A2(KEYINPUT61), .A3(G953), .ZN(n1036) );
NOR2_X1 U750 ( .A1(n1038), .A2(n1039), .ZN(n1035) );
XNOR2_X1 U751 ( .A(n1040), .B(n1041), .ZN(n1039) );
XNOR2_X1 U752 ( .A(n1042), .B(n1043), .ZN(n1041) );
NOR2_X1 U753 ( .A1(KEYINPUT24), .A2(n1044), .ZN(n1043) );
XOR2_X1 U754 ( .A(n1045), .B(n1046), .Z(n1044) );
XOR2_X1 U755 ( .A(n1047), .B(G134), .Z(n1045) );
NAND2_X1 U756 ( .A1(KEYINPUT14), .A2(n1048), .ZN(n1047) );
NAND2_X1 U757 ( .A1(n1049), .A2(KEYINPUT9), .ZN(n1042) );
XNOR2_X1 U758 ( .A(G125), .B(G140), .ZN(n1049) );
NOR2_X1 U759 ( .A1(G900), .A2(n989), .ZN(n1038) );
NOR3_X1 U760 ( .A1(n989), .A2(KEYINPUT20), .A3(n1050), .ZN(n1033) );
NOR2_X1 U761 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U762 ( .A(n1053), .B(n1054), .Z(G69) );
NOR2_X1 U763 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XNOR2_X1 U764 ( .A(n1057), .B(n1058), .ZN(n1056) );
XOR2_X1 U765 ( .A(n1059), .B(n1060), .Z(n1058) );
NOR2_X1 U766 ( .A1(KEYINPUT5), .A2(n1061), .ZN(n1059) );
NOR2_X1 U767 ( .A1(n1062), .A2(n989), .ZN(n1055) );
XNOR2_X1 U768 ( .A(G898), .B(KEYINPUT34), .ZN(n1062) );
XOR2_X1 U769 ( .A(n1063), .B(n1064), .Z(n1053) );
NOR2_X1 U770 ( .A1(KEYINPUT21), .A2(n1065), .ZN(n1064) );
NOR2_X1 U771 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
XNOR2_X1 U772 ( .A(G953), .B(KEYINPUT4), .ZN(n1067) );
NAND2_X1 U773 ( .A1(G953), .A2(n1068), .ZN(n1063) );
NAND2_X1 U774 ( .A1(G224), .A2(G898), .ZN(n1068) );
NOR2_X1 U775 ( .A1(n1069), .A2(n1070), .ZN(G66) );
XOR2_X1 U776 ( .A(n1071), .B(n1072), .Z(n1070) );
NAND2_X1 U777 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U778 ( .A1(n1069), .A2(n1075), .ZN(G63) );
XNOR2_X1 U779 ( .A(n1076), .B(n1077), .ZN(n1075) );
NAND2_X1 U780 ( .A1(n1073), .A2(G478), .ZN(n1076) );
NOR2_X1 U781 ( .A1(n1069), .A2(n1078), .ZN(G60) );
XOR2_X1 U782 ( .A(n1079), .B(n1080), .Z(n1078) );
XOR2_X1 U783 ( .A(n1081), .B(KEYINPUT53), .Z(n1080) );
NAND2_X1 U784 ( .A1(n1073), .A2(G475), .ZN(n1081) );
XNOR2_X1 U785 ( .A(n1082), .B(n1083), .ZN(G6) );
NOR2_X1 U786 ( .A1(n1069), .A2(n1084), .ZN(G57) );
XOR2_X1 U787 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR3_X1 U788 ( .A1(KEYINPUT17), .A2(n1087), .A3(n1088), .ZN(n1086) );
NOR2_X1 U789 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XOR2_X1 U790 ( .A(KEYINPUT49), .B(n1091), .Z(n1090) );
AND2_X1 U791 ( .A1(n1089), .A2(n1091), .ZN(n1087) );
AND2_X1 U792 ( .A1(n1073), .A2(G472), .ZN(n1089) );
XNOR2_X1 U793 ( .A(n1092), .B(G101), .ZN(n1085) );
NOR2_X1 U794 ( .A1(n1069), .A2(n1093), .ZN(G54) );
XOR2_X1 U795 ( .A(n1094), .B(n1095), .Z(n1093) );
XOR2_X1 U796 ( .A(n1096), .B(n1097), .Z(n1095) );
XOR2_X1 U797 ( .A(n1098), .B(n1099), .Z(n1096) );
XOR2_X1 U798 ( .A(n1100), .B(n1101), .Z(n1094) );
XNOR2_X1 U799 ( .A(n1102), .B(G110), .ZN(n1101) );
XOR2_X1 U800 ( .A(n1103), .B(n1104), .Z(n1100) );
NAND2_X1 U801 ( .A1(n1073), .A2(G469), .ZN(n1103) );
NOR2_X1 U802 ( .A1(n1069), .A2(n1105), .ZN(G51) );
XOR2_X1 U803 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR3_X1 U804 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1107) );
NOR2_X1 U805 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
INV_X1 U806 ( .A(KEYINPUT16), .ZN(n1112) );
NOR2_X1 U807 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
XNOR2_X1 U808 ( .A(KEYINPUT43), .B(n1115), .ZN(n1114) );
INV_X1 U809 ( .A(n1116), .ZN(n1113) );
NOR3_X1 U810 ( .A1(KEYINPUT16), .A2(n1117), .A3(n1118), .ZN(n1109) );
AND2_X1 U811 ( .A1(n1118), .A2(n1117), .ZN(n1108) );
XNOR2_X1 U812 ( .A(n1119), .B(n1061), .ZN(n1117) );
XNOR2_X1 U813 ( .A(n1120), .B(G110), .ZN(n1061) );
NAND3_X1 U814 ( .A1(KEYINPUT32), .A2(n1116), .A3(n1121), .ZN(n1118) );
XOR2_X1 U815 ( .A(n1115), .B(KEYINPUT43), .Z(n1121) );
NAND2_X1 U816 ( .A1(n1122), .A2(n1123), .ZN(n1115) );
XNOR2_X1 U817 ( .A(G125), .B(n1124), .ZN(n1123) );
NAND2_X1 U818 ( .A1(n1125), .A2(n1126), .ZN(n1116) );
XNOR2_X1 U819 ( .A(n1124), .B(n1127), .ZN(n1125) );
NAND2_X1 U820 ( .A1(n1073), .A2(n1128), .ZN(n1106) );
NOR2_X1 U821 ( .A1(n1129), .A2(n986), .ZN(n1073) );
AND2_X1 U822 ( .A1(n1037), .A2(n1066), .ZN(n986) );
AND2_X1 U823 ( .A1(n1130), .A2(n1131), .ZN(n1066) );
NOR4_X1 U824 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1131) );
NOR4_X1 U825 ( .A1(n1136), .A2(n985), .A3(n1137), .A4(n1083), .ZN(n1130) );
AND3_X1 U826 ( .A1(n1138), .A2(n1017), .A3(n1021), .ZN(n1083) );
AND3_X1 U827 ( .A1(n1139), .A2(n1017), .A3(n1138), .ZN(n985) );
NOR2_X1 U828 ( .A1(n1140), .A2(n1141), .ZN(n1136) );
AND4_X1 U829 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1037) );
AND4_X1 U830 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1145) );
NAND2_X1 U831 ( .A1(n1021), .A2(n1150), .ZN(n1144) );
NAND2_X1 U832 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NAND3_X1 U833 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1142) );
NOR2_X1 U834 ( .A1(n989), .A2(G952), .ZN(n1069) );
XNOR2_X1 U835 ( .A(G146), .B(n1143), .ZN(G48) );
NAND4_X1 U836 ( .A1(n1021), .A2(n1153), .A3(n1156), .A4(n1154), .ZN(n1143) );
XNOR2_X1 U837 ( .A(G143), .B(n1157), .ZN(G45) );
NAND3_X1 U838 ( .A1(n1155), .A2(n1153), .A3(n1158), .ZN(n1157) );
XNOR2_X1 U839 ( .A(n1154), .B(KEYINPUT38), .ZN(n1158) );
AND3_X1 U840 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1155) );
XNOR2_X1 U841 ( .A(G140), .B(n1149), .ZN(G42) );
NAND3_X1 U842 ( .A1(n1162), .A2(n1163), .A3(n1021), .ZN(n1149) );
XNOR2_X1 U843 ( .A(G137), .B(n1148), .ZN(G39) );
NAND3_X1 U844 ( .A1(n1163), .A2(n1156), .A3(n1013), .ZN(n1148) );
XOR2_X1 U845 ( .A(n1147), .B(n1164), .Z(G36) );
NAND2_X1 U846 ( .A1(KEYINPUT59), .A2(G134), .ZN(n1164) );
OR2_X1 U847 ( .A1(n1152), .A2(n1020), .ZN(n1147) );
XNOR2_X1 U848 ( .A(n1048), .B(n1165), .ZN(G33) );
NOR2_X1 U849 ( .A1(n1152), .A2(n1166), .ZN(n1165) );
XOR2_X1 U850 ( .A(KEYINPUT12), .B(n1021), .Z(n1166) );
NAND2_X1 U851 ( .A1(n1161), .A2(n1163), .ZN(n1152) );
AND2_X1 U852 ( .A1(n1008), .A2(n1153), .ZN(n1163) );
NOR2_X1 U853 ( .A1(n1027), .A2(n1167), .ZN(n1153) );
INV_X1 U854 ( .A(n1168), .ZN(n1167) );
XOR2_X1 U855 ( .A(n1169), .B(KEYINPUT22), .Z(n1027) );
INV_X1 U856 ( .A(n996), .ZN(n1008) );
NAND2_X1 U857 ( .A1(n1030), .A2(n1170), .ZN(n996) );
XOR2_X1 U858 ( .A(n1146), .B(n1171), .Z(G30) );
NAND2_X1 U859 ( .A1(KEYINPUT36), .A2(G128), .ZN(n1171) );
NAND4_X1 U860 ( .A1(n1156), .A2(n1139), .A3(n1172), .A4(n1169), .ZN(n1146) );
AND2_X1 U861 ( .A1(n1168), .A2(n1154), .ZN(n1172) );
INV_X1 U862 ( .A(n1020), .ZN(n1139) );
XNOR2_X1 U863 ( .A(n1173), .B(n1135), .ZN(G3) );
AND3_X1 U864 ( .A1(n1161), .A2(n1138), .A3(n1013), .ZN(n1135) );
XNOR2_X1 U865 ( .A(n1127), .B(n1174), .ZN(G27) );
NOR2_X1 U866 ( .A1(n1151), .A2(n1175), .ZN(n1174) );
XOR2_X1 U867 ( .A(KEYINPUT35), .B(n1021), .Z(n1175) );
NAND3_X1 U868 ( .A1(n1162), .A2(n1168), .A3(n1176), .ZN(n1151) );
NAND2_X1 U869 ( .A1(n1032), .A2(n1177), .ZN(n1168) );
NAND4_X1 U870 ( .A1(G953), .A2(G902), .A3(n1178), .A4(n1052), .ZN(n1177) );
INV_X1 U871 ( .A(G900), .ZN(n1052) );
XNOR2_X1 U872 ( .A(n1120), .B(n1179), .ZN(G24) );
NOR2_X1 U873 ( .A1(n1141), .A2(n1180), .ZN(n1179) );
XNOR2_X1 U874 ( .A(KEYINPUT40), .B(n1181), .ZN(n1180) );
NAND4_X1 U875 ( .A1(n1176), .A2(n1017), .A3(n1159), .A4(n1160), .ZN(n1141) );
AND2_X1 U876 ( .A1(n1182), .A2(n1183), .ZN(n1017) );
XNOR2_X1 U877 ( .A(n1134), .B(n1184), .ZN(G21) );
NAND2_X1 U878 ( .A1(KEYINPUT33), .A2(G119), .ZN(n1184) );
AND4_X1 U879 ( .A1(n1176), .A2(n1013), .A3(n1156), .A4(n1181), .ZN(n1134) );
NOR2_X1 U880 ( .A1(n1183), .A2(n1185), .ZN(n1156) );
INV_X1 U881 ( .A(n997), .ZN(n1183) );
INV_X1 U882 ( .A(n1024), .ZN(n1176) );
NAND3_X1 U883 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(G18) );
NAND2_X1 U884 ( .A1(n1137), .A2(n1189), .ZN(n1188) );
NAND2_X1 U885 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
INV_X1 U886 ( .A(KEYINPUT48), .ZN(n1191) );
XNOR2_X1 U887 ( .A(G116), .B(KEYINPUT25), .ZN(n1190) );
OR3_X1 U888 ( .A1(n1192), .A2(n1137), .A3(KEYINPUT48), .ZN(n1187) );
NOR4_X1 U889 ( .A1(n1024), .A2(n1016), .A3(n1020), .A4(n1140), .ZN(n1137) );
INV_X1 U890 ( .A(n1181), .ZN(n1140) );
NAND2_X1 U891 ( .A1(n1193), .A2(n1160), .ZN(n1020) );
INV_X1 U892 ( .A(n1161), .ZN(n1016) );
NAND2_X1 U893 ( .A1(n1010), .A2(n1154), .ZN(n1024) );
NAND2_X1 U894 ( .A1(KEYINPUT48), .A2(n1192), .ZN(n1186) );
XNOR2_X1 U895 ( .A(n1133), .B(n1194), .ZN(G15) );
NAND2_X1 U896 ( .A1(KEYINPUT27), .A2(G113), .ZN(n1194) );
AND4_X1 U897 ( .A1(n1195), .A2(n1181), .A3(n1161), .A4(n1196), .ZN(n1133) );
AND2_X1 U898 ( .A1(n1021), .A2(n1010), .ZN(n1196) );
NOR2_X1 U899 ( .A1(n1197), .A2(n1198), .ZN(n1010) );
NOR2_X1 U900 ( .A1(n1160), .A2(n1193), .ZN(n1021) );
INV_X1 U901 ( .A(n1159), .ZN(n1193) );
NOR2_X1 U902 ( .A1(n997), .A2(n1185), .ZN(n1161) );
INV_X1 U903 ( .A(n998), .ZN(n1185) );
XOR2_X1 U904 ( .A(n1132), .B(n1199), .Z(G12) );
NOR2_X1 U905 ( .A1(KEYINPUT45), .A2(n1200), .ZN(n1199) );
XNOR2_X1 U906 ( .A(G110), .B(KEYINPUT37), .ZN(n1200) );
AND3_X1 U907 ( .A1(n1013), .A2(n1138), .A3(n1162), .ZN(n1132) );
INV_X1 U908 ( .A(n1015), .ZN(n1162) );
NAND2_X1 U909 ( .A1(n1182), .A2(n997), .ZN(n1015) );
XNOR2_X1 U910 ( .A(n1201), .B(n1074), .ZN(n997) );
AND2_X1 U911 ( .A1(G217), .A2(n1202), .ZN(n1074) );
NAND2_X1 U912 ( .A1(n1072), .A2(n1129), .ZN(n1201) );
XNOR2_X1 U913 ( .A(n1203), .B(n1204), .ZN(n1072) );
XOR2_X1 U914 ( .A(n1205), .B(n1206), .Z(n1204) );
XNOR2_X1 U915 ( .A(n1207), .B(G140), .ZN(n1206) );
XOR2_X1 U916 ( .A(KEYINPUT47), .B(KEYINPUT10), .Z(n1205) );
XOR2_X1 U917 ( .A(n1208), .B(n1209), .Z(n1203) );
XOR2_X1 U918 ( .A(n1210), .B(n1211), .Z(n1209) );
NOR2_X1 U919 ( .A1(G119), .A2(KEYINPUT1), .ZN(n1211) );
AND3_X1 U920 ( .A1(G221), .A2(n989), .A3(G234), .ZN(n1210) );
XOR2_X1 U921 ( .A(n1212), .B(n1213), .Z(n1208) );
XNOR2_X1 U922 ( .A(n998), .B(KEYINPUT58), .ZN(n1182) );
XNOR2_X1 U923 ( .A(n1214), .B(G472), .ZN(n998) );
NAND2_X1 U924 ( .A1(n1215), .A2(n1129), .ZN(n1214) );
XOR2_X1 U925 ( .A(n1216), .B(n1217), .Z(n1215) );
XNOR2_X1 U926 ( .A(n1218), .B(n1091), .ZN(n1217) );
XNOR2_X1 U927 ( .A(n1219), .B(n1220), .ZN(n1091) );
XOR2_X1 U928 ( .A(G113), .B(n1221), .Z(n1220) );
NOR4_X1 U929 ( .A1(n1222), .A2(n1223), .A3(KEYINPUT39), .A4(n1224), .ZN(n1221) );
AND2_X1 U930 ( .A1(n1225), .A2(KEYINPUT56), .ZN(n1224) );
NOR2_X1 U931 ( .A1(n1226), .A2(n1192), .ZN(n1223) );
NOR2_X1 U932 ( .A1(KEYINPUT56), .A2(n1227), .ZN(n1226) );
XNOR2_X1 U933 ( .A(KEYINPUT0), .B(n1225), .ZN(n1227) );
NOR3_X1 U934 ( .A1(G116), .A2(KEYINPUT56), .A3(n1225), .ZN(n1222) );
INV_X1 U935 ( .A(G119), .ZN(n1225) );
XNOR2_X1 U936 ( .A(n1098), .B(n1228), .ZN(n1219) );
XOR2_X1 U937 ( .A(n1212), .B(n1229), .Z(n1098) );
XNOR2_X1 U938 ( .A(G128), .B(n1046), .ZN(n1212) );
NAND2_X1 U939 ( .A1(KEYINPUT63), .A2(n1092), .ZN(n1218) );
AND3_X1 U940 ( .A1(n1230), .A2(n989), .A3(G210), .ZN(n1092) );
XNOR2_X1 U941 ( .A(KEYINPUT42), .B(n1173), .ZN(n1216) );
INV_X1 U942 ( .A(G101), .ZN(n1173) );
AND3_X1 U943 ( .A1(n1195), .A2(n1181), .A3(n1169), .ZN(n1138) );
NOR2_X1 U944 ( .A1(n1198), .A2(n1029), .ZN(n1169) );
INV_X1 U945 ( .A(n1197), .ZN(n1029) );
XOR2_X1 U946 ( .A(n1000), .B(G469), .Z(n1197) );
AND2_X1 U947 ( .A1(n1231), .A2(n1129), .ZN(n1000) );
XOR2_X1 U948 ( .A(n1232), .B(n1233), .Z(n1231) );
XNOR2_X1 U949 ( .A(n1099), .B(n1234), .ZN(n1233) );
XNOR2_X1 U950 ( .A(n1046), .B(n1229), .ZN(n1234) );
XNOR2_X1 U951 ( .A(n1048), .B(G134), .ZN(n1229) );
XOR2_X1 U952 ( .A(G137), .B(KEYINPUT28), .Z(n1046) );
XOR2_X1 U953 ( .A(n1235), .B(n1236), .Z(n1232) );
XOR2_X1 U954 ( .A(n1237), .B(n1238), .Z(n1236) );
NOR2_X1 U955 ( .A1(KEYINPUT2), .A2(n1040), .ZN(n1238) );
XOR2_X1 U956 ( .A(G128), .B(n1097), .Z(n1040) );
XNOR2_X1 U957 ( .A(n1207), .B(n1239), .ZN(n1097) );
NOR2_X1 U958 ( .A1(G143), .A2(KEYINPUT3), .ZN(n1239) );
INV_X1 U959 ( .A(G146), .ZN(n1207) );
NOR2_X1 U960 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
XOR2_X1 U961 ( .A(KEYINPUT18), .B(n1242), .Z(n1241) );
NOR2_X1 U962 ( .A1(G140), .A2(n1243), .ZN(n1242) );
INV_X1 U963 ( .A(G110), .ZN(n1243) );
NOR2_X1 U964 ( .A1(G110), .A2(n1102), .ZN(n1240) );
NAND2_X1 U965 ( .A1(KEYINPUT44), .A2(n1104), .ZN(n1235) );
NOR2_X1 U966 ( .A1(n1051), .A2(G953), .ZN(n1104) );
INV_X1 U967 ( .A(G227), .ZN(n1051) );
XOR2_X1 U968 ( .A(n1003), .B(KEYINPUT26), .Z(n1198) );
AND2_X1 U969 ( .A1(G221), .A2(n1202), .ZN(n1003) );
NAND2_X1 U970 ( .A1(G234), .A2(n1129), .ZN(n1202) );
NAND2_X1 U971 ( .A1(n1032), .A2(n1244), .ZN(n1181) );
NAND4_X1 U972 ( .A1(G953), .A2(G902), .A3(n1245), .A4(n1178), .ZN(n1244) );
XOR2_X1 U973 ( .A(KEYINPUT34), .B(G898), .Z(n1245) );
NAND3_X1 U974 ( .A1(n1178), .A2(n989), .A3(G952), .ZN(n1032) );
NAND2_X1 U975 ( .A1(G237), .A2(G234), .ZN(n1178) );
XOR2_X1 U976 ( .A(n1154), .B(KEYINPUT13), .Z(n1195) );
NOR2_X1 U977 ( .A1(n1030), .A2(n1031), .ZN(n1154) );
INV_X1 U978 ( .A(n1170), .ZN(n1031) );
NAND2_X1 U979 ( .A1(G214), .A2(n1246), .ZN(n1170) );
XOR2_X1 U980 ( .A(n1247), .B(n1128), .Z(n1030) );
AND2_X1 U981 ( .A1(G210), .A2(n1246), .ZN(n1128) );
NAND2_X1 U982 ( .A1(n1129), .A2(n1230), .ZN(n1246) );
NAND2_X1 U983 ( .A1(n1248), .A2(n1129), .ZN(n1247) );
INV_X1 U984 ( .A(G902), .ZN(n1129) );
XOR2_X1 U985 ( .A(n1249), .B(n1250), .Z(n1248) );
XNOR2_X1 U986 ( .A(n1119), .B(n1213), .ZN(n1250) );
XOR2_X1 U987 ( .A(G110), .B(G125), .Z(n1213) );
NAND3_X1 U988 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1119) );
NAND2_X1 U989 ( .A1(n1057), .A2(n1060), .ZN(n1253) );
NAND2_X1 U990 ( .A1(KEYINPUT60), .A2(n1254), .ZN(n1252) );
NAND2_X1 U991 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
INV_X1 U992 ( .A(n1057), .ZN(n1256) );
XNOR2_X1 U993 ( .A(KEYINPUT23), .B(n1060), .ZN(n1255) );
NAND2_X1 U994 ( .A1(n1257), .A2(n1258), .ZN(n1251) );
INV_X1 U995 ( .A(KEYINPUT60), .ZN(n1258) );
NAND2_X1 U996 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
OR3_X1 U997 ( .A1(n1057), .A2(n1060), .A3(KEYINPUT23), .ZN(n1260) );
XOR2_X1 U998 ( .A(n1099), .B(KEYINPUT29), .Z(n1057) );
XOR2_X1 U999 ( .A(G101), .B(n1261), .Z(n1099) );
XNOR2_X1 U1000 ( .A(n1262), .B(G104), .ZN(n1261) );
INV_X1 U1001 ( .A(G107), .ZN(n1262) );
NAND2_X1 U1002 ( .A1(KEYINPUT23), .A2(n1060), .ZN(n1259) );
XNOR2_X1 U1003 ( .A(n1263), .B(n1264), .ZN(n1060) );
NOR2_X1 U1004 ( .A1(KEYINPUT57), .A2(n1192), .ZN(n1264) );
INV_X1 U1005 ( .A(G116), .ZN(n1192) );
XNOR2_X1 U1006 ( .A(G119), .B(n1265), .ZN(n1263) );
NOR2_X1 U1007 ( .A1(G113), .A2(KEYINPUT55), .ZN(n1265) );
XOR2_X1 U1008 ( .A(n1266), .B(n1267), .Z(n1249) );
XNOR2_X1 U1009 ( .A(G122), .B(n1122), .ZN(n1267) );
INV_X1 U1010 ( .A(n1126), .ZN(n1122) );
NAND2_X1 U1011 ( .A1(G224), .A2(n989), .ZN(n1126) );
NAND2_X1 U1012 ( .A1(KEYINPUT8), .A2(n1124), .ZN(n1266) );
XNOR2_X1 U1013 ( .A(n1228), .B(n1268), .ZN(n1124) );
INV_X1 U1014 ( .A(G128), .ZN(n1268) );
NAND2_X1 U1015 ( .A1(n1269), .A2(KEYINPUT15), .ZN(n1228) );
XNOR2_X1 U1016 ( .A(G143), .B(G146), .ZN(n1269) );
NOR2_X1 U1017 ( .A1(n1160), .A2(n1159), .ZN(n1013) );
NAND2_X1 U1018 ( .A1(n1270), .A2(n990), .ZN(n1159) );
NAND2_X1 U1019 ( .A1(G475), .A2(n1271), .ZN(n990) );
NAND2_X1 U1020 ( .A1(n1079), .A2(n1272), .ZN(n1271) );
XNOR2_X1 U1021 ( .A(n1002), .B(KEYINPUT41), .ZN(n1270) );
AND3_X1 U1022 ( .A1(n1272), .A2(n1273), .A3(n1079), .ZN(n1002) );
XOR2_X1 U1023 ( .A(n1274), .B(n1275), .Z(n1079) );
XNOR2_X1 U1024 ( .A(G113), .B(n1276), .ZN(n1275) );
NAND2_X1 U1025 ( .A1(KEYINPUT19), .A2(n1127), .ZN(n1276) );
INV_X1 U1026 ( .A(G125), .ZN(n1127) );
XOR2_X1 U1027 ( .A(n1277), .B(n1278), .Z(n1274) );
NOR2_X1 U1028 ( .A1(G146), .A2(KEYINPUT46), .ZN(n1278) );
XOR2_X1 U1029 ( .A(n1279), .B(n1280), .Z(n1277) );
XNOR2_X1 U1030 ( .A(n1048), .B(n1281), .ZN(n1280) );
XNOR2_X1 U1031 ( .A(G143), .B(n1102), .ZN(n1281) );
INV_X1 U1032 ( .A(G140), .ZN(n1102) );
INV_X1 U1033 ( .A(G131), .ZN(n1048) );
XOR2_X1 U1034 ( .A(n1282), .B(n1283), .Z(n1279) );
AND3_X1 U1035 ( .A1(G214), .A2(n989), .A3(n1230), .ZN(n1283) );
INV_X1 U1036 ( .A(G237), .ZN(n1230) );
XNOR2_X1 U1037 ( .A(n1284), .B(n1120), .ZN(n1282) );
NAND2_X1 U1038 ( .A1(KEYINPUT11), .A2(n1082), .ZN(n1284) );
INV_X1 U1039 ( .A(G104), .ZN(n1082) );
INV_X1 U1040 ( .A(G475), .ZN(n1273) );
XNOR2_X1 U1041 ( .A(G902), .B(KEYINPUT30), .ZN(n1272) );
NAND2_X1 U1042 ( .A1(n1285), .A2(n991), .ZN(n1160) );
NAND2_X1 U1043 ( .A1(G478), .A2(n1286), .ZN(n991) );
OR2_X1 U1044 ( .A1(n1077), .A2(G902), .ZN(n1286) );
XNOR2_X1 U1045 ( .A(n1001), .B(KEYINPUT51), .ZN(n1285) );
NOR3_X1 U1046 ( .A1(G478), .A2(G902), .A3(n1077), .ZN(n1001) );
XNOR2_X1 U1047 ( .A(n1287), .B(n1288), .ZN(n1077) );
AND3_X1 U1048 ( .A1(G217), .A2(n989), .A3(G234), .ZN(n1288) );
INV_X1 U1049 ( .A(G953), .ZN(n989) );
NAND2_X1 U1050 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
NAND2_X1 U1051 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XOR2_X1 U1052 ( .A(KEYINPUT31), .B(n1293), .Z(n1289) );
NOR2_X1 U1053 ( .A1(n1291), .A2(n1292), .ZN(n1293) );
XOR2_X1 U1054 ( .A(n1294), .B(n1295), .Z(n1292) );
XNOR2_X1 U1055 ( .A(KEYINPUT6), .B(n1120), .ZN(n1295) );
INV_X1 U1056 ( .A(G122), .ZN(n1120) );
XNOR2_X1 U1057 ( .A(G107), .B(G116), .ZN(n1294) );
XOR2_X1 U1058 ( .A(n1296), .B(n1297), .Z(n1291) );
XOR2_X1 U1059 ( .A(G143), .B(G134), .Z(n1297) );
NAND2_X1 U1060 ( .A1(KEYINPUT7), .A2(G128), .ZN(n1296) );
endmodule


