//Key = 0101111010111101001000001100100001011111101110100010100110100000


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159;

XOR2_X2 U1213 ( .A(RESTART), .B(KEYINPUT46), .Z(n1914) );
INV_X2 U1214 ( .A(n1837), .ZN(n1762) );
INV_X2 U1215 ( .A(U280), .ZN(n1763) );
NAND2_X1 U1216 ( .A1(n1620), .A2(n1621), .ZN(U344) );
NAND2_X1 U1217 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1622), .ZN(n1621) );
NAND2_X1 U1218 ( .A1(n1623), .A2(DATA_IN_7_), .ZN(n1620) );
NAND2_X1 U1219 ( .A1(n1624), .A2(n1625), .ZN(U343) );
NAND2_X1 U1220 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1622), .ZN(n1625) );
XOR2_X1 U1221 ( .A(KEYINPUT15), .B(n1626), .Z(n1624) );
NOR2_X1 U1222 ( .A1(n1627), .A2(n1622), .ZN(n1626) );
NAND2_X1 U1223 ( .A1(n1628), .A2(n1629), .ZN(U342) );
NAND2_X1 U1224 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1622), .ZN(n1629) );
NAND2_X1 U1225 ( .A1(n1623), .A2(DATA_IN_5_), .ZN(n1628) );
NAND2_X1 U1226 ( .A1(n1630), .A2(n1631), .ZN(U341) );
NAND2_X1 U1227 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1622), .ZN(n1631) );
NAND2_X1 U1228 ( .A1(n1623), .A2(DATA_IN_4_), .ZN(n1630) );
NAND2_X1 U1229 ( .A1(n1632), .A2(n1633), .ZN(U340) );
NAND2_X1 U1230 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1622), .ZN(n1633) );
NAND2_X1 U1231 ( .A1(n1623), .A2(DATA_IN_3_), .ZN(n1632) );
NAND2_X1 U1232 ( .A1(n1634), .A2(n1635), .ZN(U339) );
NAND2_X1 U1233 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1622), .ZN(n1635) );
NAND2_X1 U1234 ( .A1(n1623), .A2(DATA_IN_2_), .ZN(n1634) );
NAND2_X1 U1235 ( .A1(n1636), .A2(n1637), .ZN(U338) );
NAND2_X1 U1236 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1622), .ZN(n1637) );
NAND2_X1 U1237 ( .A1(n1623), .A2(DATA_IN_1_), .ZN(n1636) );
NAND2_X1 U1238 ( .A1(n1638), .A2(n1639), .ZN(U337) );
NAND2_X1 U1239 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1622), .ZN(n1639) );
NAND2_X1 U1240 ( .A1(n1623), .A2(DATA_IN_0_), .ZN(n1638) );
INV_X1 U1241 ( .A(n1622), .ZN(n1623) );
NAND2_X1 U1242 ( .A1(n1640), .A2(n1641), .ZN(n1622) );
NAND3_X1 U1243 ( .A1(n1642), .A2(n1643), .A3(n1644), .ZN(n1641) );
NAND2_X1 U1244 ( .A1(n1645), .A2(n1646), .ZN(U336) );
NAND2_X1 U1245 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1647), .ZN(n1646) );
NAND2_X1 U1246 ( .A1(n1648), .A2(DATA_IN_7_), .ZN(n1645) );
NAND2_X1 U1247 ( .A1(n1649), .A2(n1650), .ZN(U335) );
NAND2_X1 U1248 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1647), .ZN(n1650) );
NAND2_X1 U1249 ( .A1(n1648), .A2(DATA_IN_6_), .ZN(n1649) );
NAND2_X1 U1250 ( .A1(n1651), .A2(n1652), .ZN(U334) );
NAND2_X1 U1251 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1647), .ZN(n1652) );
NAND2_X1 U1252 ( .A1(n1653), .A2(n1648), .ZN(n1651) );
XNOR2_X1 U1253 ( .A(KEYINPUT23), .B(n1654), .ZN(n1653) );
NAND2_X1 U1254 ( .A1(n1655), .A2(n1656), .ZN(U333) );
NAND2_X1 U1255 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1647), .ZN(n1656) );
NAND2_X1 U1256 ( .A1(n1657), .A2(n1648), .ZN(n1655) );
XOR2_X1 U1257 ( .A(KEYINPUT2), .B(DATA_IN_4_), .Z(n1657) );
NAND2_X1 U1258 ( .A1(n1658), .A2(n1659), .ZN(U332) );
NAND2_X1 U1259 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1647), .ZN(n1659) );
XOR2_X1 U1260 ( .A(n1660), .B(KEYINPUT57), .Z(n1658) );
NAND2_X1 U1261 ( .A1(n1648), .A2(DATA_IN_3_), .ZN(n1660) );
NAND2_X1 U1262 ( .A1(n1661), .A2(n1662), .ZN(U331) );
NAND2_X1 U1263 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1647), .ZN(n1662) );
NAND2_X1 U1264 ( .A1(n1648), .A2(DATA_IN_2_), .ZN(n1661) );
NAND2_X1 U1265 ( .A1(n1663), .A2(n1664), .ZN(U330) );
NAND2_X1 U1266 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1647), .ZN(n1664) );
NAND2_X1 U1267 ( .A1(n1648), .A2(DATA_IN_1_), .ZN(n1663) );
NAND2_X1 U1268 ( .A1(n1665), .A2(n1666), .ZN(U329) );
NAND2_X1 U1269 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1647), .ZN(n1666) );
NAND2_X1 U1270 ( .A1(n1648), .A2(DATA_IN_0_), .ZN(n1665) );
INV_X1 U1271 ( .A(n1647), .ZN(n1648) );
NAND2_X1 U1272 ( .A1(n1640), .A2(n1667), .ZN(n1647) );
NAND2_X1 U1273 ( .A1(n1668), .A2(n1643), .ZN(n1667) );
NAND3_X1 U1274 ( .A1(n1644), .A2(n1642), .A3(n1669), .ZN(n1668) );
NAND2_X1 U1275 ( .A1(n1670), .A2(n1671), .ZN(n1669) );
NAND3_X1 U1276 ( .A1(n1672), .A2(n1673), .A3(n1674), .ZN(n1671) );
NAND2_X1 U1277 ( .A1(DATA_IN_6_), .A2(n1675), .ZN(n1674) );
NAND3_X1 U1278 ( .A1(n1676), .A2(n1677), .A3(n1678), .ZN(n1673) );
NAND2_X1 U1279 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1627), .ZN(n1678) );
NAND3_X1 U1280 ( .A1(n1679), .A2(n1680), .A3(n1681), .ZN(n1677) );
NAND2_X1 U1281 ( .A1(DATA_IN_4_), .A2(n1682), .ZN(n1681) );
NAND3_X1 U1282 ( .A1(n1683), .A2(n1684), .A3(n1685), .ZN(n1680) );
OR2_X1 U1283 ( .A1(n1682), .A2(DATA_IN_4_), .ZN(n1685) );
INV_X1 U1284 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1682) );
NAND3_X1 U1285 ( .A1(n1686), .A2(n1687), .A3(n1688), .ZN(n1684) );
NAND2_X1 U1286 ( .A1(DATA_IN_3_), .A2(n1689), .ZN(n1688) );
NAND3_X1 U1287 ( .A1(n1690), .A2(n1691), .A3(n1692), .ZN(n1687) );
NAND2_X1 U1288 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1693), .ZN(n1692) );
NAND3_X1 U1289 ( .A1(n1694), .A2(n1695), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1691) );
INV_X1 U1290 ( .A(DATA_IN_0_), .ZN(n1695) );
NAND2_X1 U1291 ( .A1(DATA_IN_1_), .A2(n1696), .ZN(n1694) );
NAND2_X1 U1292 ( .A1(n1697), .A2(n1698), .ZN(n1690) );
XNOR2_X1 U1293 ( .A(n1699), .B(KEYINPUT16), .ZN(n1697) );
NAND2_X1 U1294 ( .A1(DATA_IN_2_), .A2(n1699), .ZN(n1686) );
NAND2_X1 U1295 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1700), .ZN(n1683) );
NAND2_X1 U1296 ( .A1(DATA_IN_5_), .A2(n1701), .ZN(n1679) );
XOR2_X1 U1297 ( .A(RMIN_REG_5__SCAN_IN), .B(KEYINPUT4), .Z(n1701) );
NAND2_X1 U1298 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1654), .ZN(n1676) );
NAND2_X1 U1299 ( .A1(n1702), .A2(RMIN_REG_7__SCAN_IN), .ZN(n1672) );
XNOR2_X1 U1300 ( .A(DATA_IN_7_), .B(KEYINPUT45), .ZN(n1702) );
NAND2_X1 U1301 ( .A1(DATA_IN_7_), .A2(n1703), .ZN(n1670) );
NAND2_X1 U1302 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1704), .ZN(n1642) );
XNOR2_X1 U1303 ( .A(KEYINPUT55), .B(n1705), .ZN(n1704) );
NAND3_X1 U1304 ( .A1(n1706), .A2(n1707), .A3(n1708), .ZN(n1644) );
NAND2_X1 U1305 ( .A1(DATA_IN_7_), .A2(n1709), .ZN(n1708) );
NAND3_X1 U1306 ( .A1(n1710), .A2(n1711), .A3(n1712), .ZN(n1707) );
XOR2_X1 U1307 ( .A(KEYINPUT50), .B(n1713), .Z(n1712) );
NOR2_X1 U1308 ( .A1(n1714), .A2(n1715), .ZN(n1713) );
NOR2_X1 U1309 ( .A1(n1716), .A2(n1717), .ZN(n1715) );
AND2_X1 U1310 ( .A1(n1718), .A2(DATA_IN_4_), .ZN(n1717) );
NOR2_X1 U1311 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1719), .ZN(n1716) );
NOR2_X1 U1312 ( .A1(DATA_IN_4_), .A2(n1718), .ZN(n1719) );
NAND2_X1 U1313 ( .A1(n1720), .A2(n1721), .ZN(n1718) );
NAND2_X1 U1314 ( .A1(DATA_IN_3_), .A2(n1722), .ZN(n1721) );
XOR2_X1 U1315 ( .A(KEYINPUT39), .B(n1723), .Z(n1720) );
NOR3_X1 U1316 ( .A1(n1724), .A2(n1725), .A3(n1726), .ZN(n1723) );
NOR2_X1 U1317 ( .A1(DATA_IN_2_), .A2(n1727), .ZN(n1726) );
NOR3_X1 U1318 ( .A1(n1728), .A2(n1729), .A3(n1730), .ZN(n1725) );
NOR2_X1 U1319 ( .A1(n1698), .A2(n1731), .ZN(n1730) );
XNOR2_X1 U1320 ( .A(n1727), .B(KEYINPUT32), .ZN(n1731) );
INV_X1 U1321 ( .A(DATA_IN_2_), .ZN(n1698) );
NOR3_X1 U1322 ( .A1(n1732), .A2(RMAX_REG_0__SCAN_IN), .A3(n1733), .ZN(n1729));
NOR2_X1 U1323 ( .A1(DATA_IN_1_), .A2(n1734), .ZN(n1733) );
XNOR2_X1 U1324 ( .A(DATA_IN_0_), .B(KEYINPUT0), .ZN(n1732) );
NOR2_X1 U1325 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1693), .ZN(n1728) );
NOR2_X1 U1326 ( .A1(DATA_IN_3_), .A2(n1722), .ZN(n1724) );
NOR2_X1 U1327 ( .A1(DATA_IN_5_), .A2(n1735), .ZN(n1714) );
NAND2_X1 U1328 ( .A1(DATA_IN_5_), .A2(n1735), .ZN(n1711) );
INV_X1 U1329 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1735) );
NAND2_X1 U1330 ( .A1(DATA_IN_6_), .A2(n1736), .ZN(n1710) );
NAND2_X1 U1331 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1627), .ZN(n1706) );
INV_X1 U1332 ( .A(DATA_IN_6_), .ZN(n1627) );
NAND2_X1 U1333 ( .A1(n1737), .A2(n1738), .ZN(U328) );
NAND2_X1 U1334 ( .A1(n1739), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1738) );
XOR2_X1 U1335 ( .A(n1740), .B(KEYINPUT7), .Z(n1739) );
NAND2_X1 U1336 ( .A1(n1741), .A2(DATA_IN_7_), .ZN(n1737) );
NAND2_X1 U1337 ( .A1(n1742), .A2(n1743), .ZN(U327) );
NAND2_X1 U1338 ( .A1(n1741), .A2(DATA_IN_6_), .ZN(n1743) );
NAND2_X1 U1339 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1740), .ZN(n1742) );
NAND2_X1 U1340 ( .A1(n1744), .A2(n1745), .ZN(U326) );
NAND2_X1 U1341 ( .A1(n1746), .A2(n1741), .ZN(n1745) );
XNOR2_X1 U1342 ( .A(DATA_IN_5_), .B(KEYINPUT1), .ZN(n1746) );
NAND2_X1 U1343 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1740), .ZN(n1744) );
NAND2_X1 U1344 ( .A1(n1747), .A2(n1748), .ZN(U325) );
NAND2_X1 U1345 ( .A1(n1741), .A2(DATA_IN_4_), .ZN(n1748) );
NAND2_X1 U1346 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1740), .ZN(n1747) );
NAND2_X1 U1347 ( .A1(n1749), .A2(n1750), .ZN(U324) );
NAND2_X1 U1348 ( .A1(n1741), .A2(DATA_IN_3_), .ZN(n1750) );
NAND2_X1 U1349 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1740), .ZN(n1749) );
NAND2_X1 U1350 ( .A1(n1751), .A2(n1752), .ZN(U323) );
NAND2_X1 U1351 ( .A1(n1753), .A2(n1740), .ZN(n1752) );
XOR2_X1 U1352 ( .A(RLAST_REG_2__SCAN_IN), .B(KEYINPUT59), .Z(n1753) );
NAND2_X1 U1353 ( .A1(n1741), .A2(DATA_IN_2_), .ZN(n1751) );
NAND2_X1 U1354 ( .A1(n1754), .A2(n1755), .ZN(U322) );
NAND2_X1 U1355 ( .A1(n1741), .A2(DATA_IN_1_), .ZN(n1755) );
NAND2_X1 U1356 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1740), .ZN(n1754) );
NAND2_X1 U1357 ( .A1(n1756), .A2(n1757), .ZN(U321) );
NAND2_X1 U1358 ( .A1(n1741), .A2(DATA_IN_0_), .ZN(n1757) );
AND2_X1 U1359 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1758), .ZN(n1741) );
NAND2_X1 U1360 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1740), .ZN(n1756) );
NAND2_X1 U1361 ( .A1(n1640), .A2(n1758), .ZN(n1740) );
NAND2_X1 U1362 ( .A1(n1759), .A2(n1643), .ZN(n1758) );
INV_X1 U1363 ( .A(U375), .ZN(n1640) );
NOR2_X1 U1364 ( .A1(STATO_REG_0__SCAN_IN), .A2(STATO_REG_1__SCAN_IN), .ZN(U375) );
NAND2_X1 U1365 ( .A1(n1760), .A2(n1761), .ZN(U320) );
NAND2_X1 U1366 ( .A1(n1762), .A2(DATA_IN_7_), .ZN(n1761) );
NAND2_X1 U1367 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1763), .ZN(n1760) );
NAND2_X1 U1368 ( .A1(n1764), .A2(n1765), .ZN(U319) );
NAND2_X1 U1369 ( .A1(n1762), .A2(DATA_IN_6_), .ZN(n1765) );
NAND2_X1 U1370 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1763), .ZN(n1764) );
NAND2_X1 U1371 ( .A1(n1766), .A2(n1767), .ZN(U318) );
NAND2_X1 U1372 ( .A1(n1762), .A2(n1768), .ZN(n1767) );
XNOR2_X1 U1373 ( .A(KEYINPUT30), .B(n1654), .ZN(n1768) );
NAND2_X1 U1374 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1763), .ZN(n1766) );
NAND2_X1 U1375 ( .A1(n1769), .A2(n1770), .ZN(U317) );
NAND2_X1 U1376 ( .A1(n1762), .A2(DATA_IN_4_), .ZN(n1770) );
NAND2_X1 U1377 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1763), .ZN(n1769) );
NAND2_X1 U1378 ( .A1(n1771), .A2(n1772), .ZN(U316) );
NAND2_X1 U1379 ( .A1(n1762), .A2(DATA_IN_3_), .ZN(n1772) );
NAND2_X1 U1380 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1763), .ZN(n1771) );
NAND2_X1 U1381 ( .A1(n1773), .A2(n1774), .ZN(U315) );
NAND2_X1 U1382 ( .A1(n1762), .A2(DATA_IN_2_), .ZN(n1774) );
NAND2_X1 U1383 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1763), .ZN(n1773) );
NAND2_X1 U1384 ( .A1(n1775), .A2(n1776), .ZN(U314) );
NAND2_X1 U1385 ( .A1(n1762), .A2(DATA_IN_1_), .ZN(n1776) );
NAND2_X1 U1386 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1763), .ZN(n1775) );
NAND2_X1 U1387 ( .A1(n1777), .A2(n1778), .ZN(U313) );
NAND2_X1 U1388 ( .A1(n1762), .A2(DATA_IN_0_), .ZN(n1778) );
NAND2_X1 U1389 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1763), .ZN(n1777) );
NAND2_X1 U1390 ( .A1(n1779), .A2(n1780), .ZN(U312) );
NAND2_X1 U1391 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1762), .ZN(n1780) );
NAND2_X1 U1392 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1763), .ZN(n1779) );
NAND2_X1 U1393 ( .A1(n1781), .A2(n1782), .ZN(U311) );
NAND2_X1 U1394 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1763), .ZN(n1782) );
XOR2_X1 U1395 ( .A(KEYINPUT38), .B(n1783), .Z(n1781) );
AND2_X1 U1396 ( .A1(n1762), .A2(REG1_REG_6__SCAN_IN), .ZN(n1783) );
NAND2_X1 U1397 ( .A1(n1784), .A2(n1785), .ZN(U310) );
NAND2_X1 U1398 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1762), .ZN(n1785) );
NAND2_X1 U1399 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1763), .ZN(n1784) );
NAND2_X1 U1400 ( .A1(n1786), .A2(n1787), .ZN(U309) );
NAND2_X1 U1401 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1762), .ZN(n1787) );
NAND2_X1 U1402 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1763), .ZN(n1786) );
NAND2_X1 U1403 ( .A1(n1788), .A2(n1789), .ZN(U308) );
NAND2_X1 U1404 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1762), .ZN(n1789) );
NAND2_X1 U1405 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1763), .ZN(n1788) );
NAND2_X1 U1406 ( .A1(n1790), .A2(n1791), .ZN(U307) );
NAND2_X1 U1407 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1762), .ZN(n1791) );
XOR2_X1 U1408 ( .A(KEYINPUT12), .B(n1792), .Z(n1790) );
AND2_X1 U1409 ( .A1(n1763), .A2(REG2_REG_2__SCAN_IN), .ZN(n1792) );
NAND2_X1 U1410 ( .A1(n1793), .A2(n1794), .ZN(U306) );
NAND2_X1 U1411 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1762), .ZN(n1794) );
NAND2_X1 U1412 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1763), .ZN(n1793) );
NAND2_X1 U1413 ( .A1(n1795), .A2(n1796), .ZN(U305) );
NAND2_X1 U1414 ( .A1(n1797), .A2(n1763), .ZN(n1796) );
XNOR2_X1 U1415 ( .A(REG2_REG_0__SCAN_IN), .B(KEYINPUT42), .ZN(n1797) );
NAND2_X1 U1416 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1762), .ZN(n1795) );
NAND2_X1 U1417 ( .A1(n1798), .A2(n1799), .ZN(U304) );
NAND2_X1 U1418 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1762), .ZN(n1799) );
NAND2_X1 U1419 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1763), .ZN(n1798) );
NAND2_X1 U1420 ( .A1(n1800), .A2(n1801), .ZN(U303) );
NAND2_X1 U1421 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1762), .ZN(n1801) );
NAND2_X1 U1422 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1763), .ZN(n1800) );
NAND2_X1 U1423 ( .A1(n1802), .A2(n1803), .ZN(U302) );
NAND2_X1 U1424 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1762), .ZN(n1803) );
NAND2_X1 U1425 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1763), .ZN(n1802) );
NAND2_X1 U1426 ( .A1(n1804), .A2(n1805), .ZN(U301) );
NAND2_X1 U1427 ( .A1(n1762), .A2(n1806), .ZN(n1805) );
XOR2_X1 U1428 ( .A(REG2_REG_4__SCAN_IN), .B(KEYINPUT49), .Z(n1806) );
NAND2_X1 U1429 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1763), .ZN(n1804) );
NAND2_X1 U1430 ( .A1(n1807), .A2(n1808), .ZN(U300) );
NAND2_X1 U1431 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1762), .ZN(n1808) );
XOR2_X1 U1432 ( .A(KEYINPUT3), .B(n1809), .Z(n1807) );
AND2_X1 U1433 ( .A1(n1763), .A2(REG3_REG_3__SCAN_IN), .ZN(n1809) );
NAND2_X1 U1434 ( .A1(n1810), .A2(n1811), .ZN(U299) );
NAND2_X1 U1435 ( .A1(n1812), .A2(n1763), .ZN(n1811) );
XNOR2_X1 U1436 ( .A(REG3_REG_2__SCAN_IN), .B(KEYINPUT33), .ZN(n1812) );
NAND2_X1 U1437 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1762), .ZN(n1810) );
NAND2_X1 U1438 ( .A1(n1813), .A2(n1814), .ZN(U298) );
NAND2_X1 U1439 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1762), .ZN(n1814) );
NAND2_X1 U1440 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1763), .ZN(n1813) );
NAND2_X1 U1441 ( .A1(n1815), .A2(n1816), .ZN(U297) );
NAND2_X1 U1442 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1762), .ZN(n1816) );
NAND2_X1 U1443 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1763), .ZN(n1815) );
NAND2_X1 U1444 ( .A1(n1817), .A2(n1818), .ZN(U296) );
NAND2_X1 U1445 ( .A1(n1819), .A2(REG3_REG_7__SCAN_IN), .ZN(n1818) );
XNOR2_X1 U1446 ( .A(n1762), .B(KEYINPUT24), .ZN(n1819) );
NAND2_X1 U1447 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1763), .ZN(n1817) );
NAND2_X1 U1448 ( .A1(n1820), .A2(n1821), .ZN(U295) );
NAND2_X1 U1449 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1762), .ZN(n1821) );
NAND2_X1 U1450 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1763), .ZN(n1820) );
NAND2_X1 U1451 ( .A1(n1822), .A2(n1823), .ZN(U294) );
NAND2_X1 U1452 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1762), .ZN(n1823) );
NAND2_X1 U1453 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1763), .ZN(n1822) );
NAND2_X1 U1454 ( .A1(n1824), .A2(n1825), .ZN(U293) );
NAND2_X1 U1455 ( .A1(n1826), .A2(n1762), .ZN(n1825) );
XNOR2_X1 U1456 ( .A(REG3_REG_4__SCAN_IN), .B(KEYINPUT28), .ZN(n1826) );
NAND2_X1 U1457 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1763), .ZN(n1824) );
NAND2_X1 U1458 ( .A1(n1827), .A2(n1828), .ZN(U292) );
NAND2_X1 U1459 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1762), .ZN(n1828) );
XOR2_X1 U1460 ( .A(KEYINPUT36), .B(n1829), .Z(n1827) );
NOR2_X1 U1461 ( .A1(U280), .A2(n1830), .ZN(n1829) );
NAND2_X1 U1462 ( .A1(n1831), .A2(n1832), .ZN(U291) );
NAND2_X1 U1463 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1762), .ZN(n1832) );
NAND2_X1 U1464 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1763), .ZN(n1831) );
NAND2_X1 U1465 ( .A1(n1833), .A2(n1834), .ZN(U290) );
NAND2_X1 U1466 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1762), .ZN(n1834) );
NAND2_X1 U1467 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1763), .ZN(n1833) );
NAND2_X1 U1468 ( .A1(n1835), .A2(n1836), .ZN(U289) );
NAND2_X1 U1469 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1762), .ZN(n1836) );
NAND2_X1 U1470 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1763), .ZN(n1835) );
NAND4_X1 U1471 ( .A1(n1838), .A2(n1839), .A3(n1840), .A4(n1841), .ZN(U288));
OR2_X1 U1472 ( .A1(n1842), .A2(n1843), .ZN(n1841) );
NOR2_X1 U1473 ( .A1(n1844), .A2(n1845), .ZN(n1840) );
NOR2_X1 U1474 ( .A1(n1846), .A2(n1847), .ZN(n1845) );
XNOR2_X1 U1475 ( .A(n1848), .B(KEYINPUT51), .ZN(n1846) );
NAND2_X1 U1476 ( .A1(n1849), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1839) );
NAND2_X1 U1477 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1763), .ZN(n1838) );
NAND4_X1 U1478 ( .A1(n1850), .A2(n1851), .A3(n1852), .A4(n1853), .ZN(U287));
NOR4_X1 U1479 ( .A1(n1844), .A2(n1854), .A3(n1855), .A4(n1856), .ZN(n1853));
NOR2_X1 U1480 ( .A1(n1857), .A2(n1858), .ZN(n1856) );
INV_X1 U1481 ( .A(RLAST_REG_6__SCAN_IN), .ZN(n1858) );
XNOR2_X1 U1482 ( .A(n1849), .B(KEYINPUT47), .ZN(n1857) );
NOR2_X1 U1483 ( .A1(n1859), .A2(n1860), .ZN(n1855) );
XNOR2_X1 U1484 ( .A(REG4_REG_6__SCAN_IN), .B(KEYINPUT9), .ZN(n1859) );
NOR3_X1 U1485 ( .A1(n1861), .A2(n1862), .A3(n1863), .ZN(n1854) );
AND3_X1 U1486 ( .A1(n1862), .A2(n1861), .A3(n1864), .ZN(n1844) );
OR2_X1 U1487 ( .A1(n1865), .A2(n1866), .ZN(n1861) );
NOR2_X1 U1488 ( .A1(n1867), .A2(n1868), .ZN(n1852) );
NOR3_X1 U1489 ( .A1(n1869), .A2(n1870), .A3(n1871), .ZN(n1868) );
INV_X1 U1490 ( .A(n1843), .ZN(n1869) );
NOR3_X1 U1491 ( .A1(n1843), .A2(KEYINPUT14), .A3(n1842), .ZN(n1867) );
NAND2_X1 U1492 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1763), .ZN(n1851) );
NAND2_X1 U1493 ( .A1(KEYINPUT14), .A2(n1872), .ZN(n1850) );
NAND2_X1 U1494 ( .A1(n1871), .A2(n1873), .ZN(n1872) );
NAND2_X1 U1495 ( .A1(n1874), .A2(n1843), .ZN(n1873) );
NAND4_X1 U1496 ( .A1(n1875), .A2(n1876), .A3(n1877), .A4(n1878), .ZN(U286));
NOR4_X1 U1497 ( .A1(n1879), .A2(n1880), .A3(n1881), .A4(n1882), .ZN(n1878));
AND2_X1 U1498 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1763), .ZN(n1882) );
NOR2_X1 U1499 ( .A1(n1883), .A2(n1860), .ZN(n1881) );
INV_X1 U1500 ( .A(n1848), .ZN(n1860) );
NOR2_X1 U1501 ( .A1(n1871), .A2(n1884), .ZN(n1880) );
NAND3_X1 U1502 ( .A1(n1885), .A2(n1886), .A3(n1874), .ZN(n1871) );
NOR2_X1 U1503 ( .A1(n1870), .A2(n1842), .ZN(n1879) );
INV_X1 U1504 ( .A(n1884), .ZN(n1870) );
NAND2_X1 U1505 ( .A1(n1843), .A2(n1887), .ZN(n1884) );
NAND2_X1 U1506 ( .A1(n1888), .A2(n1889), .ZN(n1887) );
NAND2_X1 U1507 ( .A1(n1890), .A2(n1891), .ZN(n1843) );
XNOR2_X1 U1508 ( .A(n1888), .B(KEYINPUT22), .ZN(n1890) );
NAND2_X1 U1509 ( .A1(n1849), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1877) );
NAND2_X1 U1510 ( .A1(n1892), .A2(n1864), .ZN(n1876) );
XNOR2_X1 U1511 ( .A(n1893), .B(n1866), .ZN(n1892) );
NOR2_X1 U1512 ( .A1(n1862), .A2(n1894), .ZN(n1866) );
AND2_X1 U1513 ( .A1(n1888), .A2(n1895), .ZN(n1894) );
NOR2_X1 U1514 ( .A1(n1895), .A2(n1888), .ZN(n1862) );
NAND2_X1 U1515 ( .A1(n1896), .A2(n1888), .ZN(n1875) );
AND2_X1 U1516 ( .A1(n1897), .A2(n1898), .ZN(n1888) );
NAND3_X1 U1517 ( .A1(n1899), .A2(n1900), .A3(n1901), .ZN(n1898) );
XOR2_X1 U1518 ( .A(n1902), .B(n1903), .Z(n1901) );
XOR2_X1 U1519 ( .A(KEYINPUT8), .B(n1904), .Z(n1899) );
NOR2_X1 U1520 ( .A1(n1905), .A2(n1906), .ZN(n1904) );
NAND3_X1 U1521 ( .A1(n1907), .A2(n1908), .A3(n1909), .ZN(n1897) );
XOR2_X1 U1522 ( .A(n1910), .B(n1903), .Z(n1909) );
AND2_X1 U1523 ( .A1(n1911), .A2(n1912), .ZN(n1903) );
NAND2_X1 U1524 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1913), .ZN(n1912) );
XOR2_X1 U1525 ( .A(RESTART), .B(KEYINPUT29), .Z(n1913) );
NAND2_X1 U1526 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1914), .ZN(n1911) );
NAND2_X1 U1527 ( .A1(KEYINPUT43), .A2(n1902), .ZN(n1910) );
NAND2_X1 U1528 ( .A1(n1915), .A2(n1916), .ZN(n1902) );
NAND2_X1 U1529 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1917), .ZN(n1916) );
XOR2_X1 U1530 ( .A(RESTART), .B(KEYINPUT48), .Z(n1917) );
NAND2_X1 U1531 ( .A1(DATA_IN_6_), .A2(n1914), .ZN(n1915) );
NAND2_X1 U1532 ( .A1(n1900), .A2(n1906), .ZN(n1907) );
NAND4_X1 U1533 ( .A1(n1918), .A2(n1919), .A3(n1920), .A4(n1921), .ZN(U285));
NOR3_X1 U1534 ( .A1(n1922), .A2(n1923), .A3(n1924), .ZN(n1921) );
NOR2_X1 U1535 ( .A1(n1925), .A2(n1842), .ZN(n1924) );
NAND2_X1 U1536 ( .A1(n1874), .A2(n1926), .ZN(n1842) );
NAND2_X1 U1537 ( .A1(n1885), .A2(n1886), .ZN(n1926) );
NOR2_X1 U1538 ( .A1(n1885), .A2(n1927), .ZN(n1925) );
XOR2_X1 U1539 ( .A(n1886), .B(KEYINPUT27), .Z(n1927) );
NAND2_X1 U1540 ( .A1(n1889), .A2(n1928), .ZN(n1886) );
NAND2_X1 U1541 ( .A1(n1929), .A2(n1930), .ZN(n1928) );
INV_X1 U1542 ( .A(n1891), .ZN(n1889) );
NOR2_X1 U1543 ( .A1(n1930), .A2(n1929), .ZN(n1891) );
NOR3_X1 U1544 ( .A1(n1863), .A2(n1893), .A3(n1931), .ZN(n1923) );
XOR2_X1 U1545 ( .A(n1932), .B(KEYINPUT35), .Z(n1931) );
NAND2_X1 U1546 ( .A1(n1933), .A2(n1934), .ZN(n1932) );
NAND2_X1 U1547 ( .A1(n1935), .A2(n1936), .ZN(n1934) );
INV_X1 U1548 ( .A(n1937), .ZN(n1933) );
INV_X1 U1549 ( .A(n1865), .ZN(n1893) );
NAND3_X1 U1550 ( .A1(n1937), .A2(n1936), .A3(n1935), .ZN(n1865) );
NAND2_X1 U1551 ( .A1(n1895), .A2(n1938), .ZN(n1937) );
NAND2_X1 U1552 ( .A1(n1930), .A2(n1939), .ZN(n1938) );
NAND2_X1 U1553 ( .A1(n1940), .A2(n1941), .ZN(n1895) );
XNOR2_X1 U1554 ( .A(KEYINPUT19), .B(n1939), .ZN(n1941) );
NOR2_X1 U1555 ( .A1(n1940), .A2(n1942), .ZN(n1922) );
INV_X1 U1556 ( .A(n1930), .ZN(n1940) );
NAND2_X1 U1557 ( .A1(n1943), .A2(n1944), .ZN(n1930) );
NAND2_X1 U1558 ( .A1(n1945), .A2(n1946), .ZN(n1944) );
NAND2_X1 U1559 ( .A1(n1908), .A2(n1900), .ZN(n1946) );
NAND2_X1 U1560 ( .A1(n1947), .A2(n1948), .ZN(n1900) );
INV_X1 U1561 ( .A(n1905), .ZN(n1908) );
NOR2_X1 U1562 ( .A1(n1948), .A2(n1947), .ZN(n1905) );
INV_X1 U1563 ( .A(n1906), .ZN(n1945) );
NAND2_X1 U1564 ( .A1(n1949), .A2(n1906), .ZN(n1943) );
NAND2_X1 U1565 ( .A1(n1950), .A2(n1951), .ZN(n1906) );
NAND2_X1 U1566 ( .A1(n1952), .A2(n1953), .ZN(n1951) );
NAND2_X1 U1567 ( .A1(n1954), .A2(n1955), .ZN(n1953) );
OR2_X1 U1568 ( .A1(n1955), .A2(n1954), .ZN(n1950) );
XOR2_X1 U1569 ( .A(n1948), .B(n1947), .Z(n1949) );
NAND2_X1 U1570 ( .A1(n1956), .A2(n1957), .ZN(n1947) );
NAND2_X1 U1571 ( .A1(DATA_IN_5_), .A2(n1914), .ZN(n1957) );
NAND2_X1 U1572 ( .A1(RESTART), .A2(RMAX_REG_5__SCAN_IN), .ZN(n1956) );
NAND2_X1 U1573 ( .A1(n1958), .A2(n1959), .ZN(n1948) );
NAND2_X1 U1574 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1914), .ZN(n1959) );
NAND2_X1 U1575 ( .A1(RESTART), .A2(RMIN_REG_5__SCAN_IN), .ZN(n1958) );
XOR2_X1 U1576 ( .A(n1960), .B(KEYINPUT20), .Z(n1920) );
NAND2_X1 U1577 ( .A1(n1848), .A2(REG4_REG_4__SCAN_IN), .ZN(n1960) );
NAND2_X1 U1578 ( .A1(n1849), .A2(RLAST_REG_4__SCAN_IN), .ZN(n1919) );
NAND2_X1 U1579 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1763), .ZN(n1918) );
NAND4_X1 U1580 ( .A1(n1961), .A2(n1962), .A3(n1963), .A4(n1964), .ZN(U284));
NOR3_X1 U1581 ( .A1(n1965), .A2(n1966), .A3(n1967), .ZN(n1964) );
NOR2_X1 U1582 ( .A1(n1863), .A2(n1968), .ZN(n1967) );
XNOR2_X1 U1583 ( .A(n1935), .B(n1936), .ZN(n1968) );
NAND2_X1 U1584 ( .A1(n1939), .A2(n1969), .ZN(n1936) );
NAND2_X1 U1585 ( .A1(n1970), .A2(n1971), .ZN(n1969) );
NAND2_X1 U1586 ( .A1(n1972), .A2(n1973), .ZN(n1971) );
XNOR2_X1 U1587 ( .A(n1974), .B(KEYINPUT52), .ZN(n1972) );
INV_X1 U1588 ( .A(n1975), .ZN(n1939) );
NOR3_X1 U1589 ( .A1(n1976), .A2(n1885), .A3(n1977), .ZN(n1966) );
NOR2_X1 U1590 ( .A1(n1978), .A2(n1979), .ZN(n1977) );
AND2_X1 U1591 ( .A1(n1978), .A2(n1979), .ZN(n1885) );
NAND2_X1 U1592 ( .A1(n1929), .A2(n1980), .ZN(n1979) );
NAND2_X1 U1593 ( .A1(n1970), .A2(n1981), .ZN(n1980) );
NAND2_X1 U1594 ( .A1(n1973), .A2(n1974), .ZN(n1981) );
AND2_X1 U1595 ( .A1(n1982), .A2(n1983), .ZN(n1929) );
OR4_X1 U1596 ( .A1(n1970), .A2(n1974), .A3(n1984), .A4(KEYINPUT56), .ZN(n1983) );
NAND2_X1 U1597 ( .A1(n1975), .A2(KEYINPUT56), .ZN(n1982) );
NOR3_X1 U1598 ( .A1(n1985), .A2(n1970), .A3(n1984), .ZN(n1975) );
NOR2_X1 U1599 ( .A1(n1986), .A2(n1987), .ZN(n1965) );
INV_X1 U1600 ( .A(RLAST_REG_3__SCAN_IN), .ZN(n1987) );
XNOR2_X1 U1601 ( .A(n1849), .B(KEYINPUT53), .ZN(n1986) );
NAND2_X1 U1602 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1763), .ZN(n1963) );
NAND2_X1 U1603 ( .A1(n1896), .A2(n1970), .ZN(n1962) );
XOR2_X1 U1604 ( .A(n1955), .B(n1988), .Z(n1970) );
XOR2_X1 U1605 ( .A(n1952), .B(n1989), .Z(n1988) );
NOR2_X1 U1606 ( .A1(KEYINPUT63), .A2(n1954), .ZN(n1989) );
AND2_X1 U1607 ( .A1(n1990), .A2(n1991), .ZN(n1954) );
NAND2_X1 U1608 ( .A1(n1992), .A2(n1993), .ZN(n1991) );
XOR2_X1 U1609 ( .A(n1994), .B(KEYINPUT44), .Z(n1992) );
NAND2_X1 U1610 ( .A1(n1995), .A2(n1996), .ZN(n1990) );
NAND2_X1 U1611 ( .A1(n1997), .A2(n1998), .ZN(n1996) );
XNOR2_X1 U1612 ( .A(KEYINPUT44), .B(n1994), .ZN(n1998) );
XNOR2_X1 U1613 ( .A(n1993), .B(KEYINPUT31), .ZN(n1997) );
INV_X1 U1614 ( .A(n1999), .ZN(n1993) );
AND2_X1 U1615 ( .A1(n2000), .A2(n2001), .ZN(n1952) );
NAND2_X1 U1616 ( .A1(RESTART), .A2(RMIN_REG_4__SCAN_IN), .ZN(n2001) );
XOR2_X1 U1617 ( .A(n2002), .B(KEYINPUT62), .Z(n2000) );
NAND2_X1 U1618 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1914), .ZN(n2002) );
NAND2_X1 U1619 ( .A1(n2003), .A2(n2004), .ZN(n1955) );
NAND2_X1 U1620 ( .A1(DATA_IN_4_), .A2(n1914), .ZN(n2004) );
NAND2_X1 U1621 ( .A1(RESTART), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2003) );
NAND2_X1 U1622 ( .A1(n1848), .A2(REG4_REG_3__SCAN_IN), .ZN(n1961) );
NAND4_X1 U1623 ( .A1(n2005), .A2(n2006), .A3(n2007), .A4(n2008), .ZN(U283));
NOR3_X1 U1624 ( .A1(n2009), .A2(n2010), .A3(n2011), .ZN(n2008) );
NOR2_X1 U1625 ( .A1(n2012), .A2(n1976), .ZN(n2011) );
INV_X1 U1626 ( .A(n1874), .ZN(n1976) );
XOR2_X1 U1627 ( .A(n2013), .B(KEYINPUT41), .Z(n2012) );
OR2_X1 U1628 ( .A1(n1978), .A2(n2014), .ZN(n2013) );
AND2_X1 U1629 ( .A1(n2015), .A2(n2016), .ZN(n1978) );
XNOR2_X1 U1630 ( .A(n1974), .B(n1973), .ZN(n2015) );
NOR3_X1 U1631 ( .A1(n2017), .A2(n1935), .A3(n1863), .ZN(n2010) );
INV_X1 U1632 ( .A(n1864), .ZN(n1863) );
AND2_X1 U1633 ( .A1(n2016), .A2(n2018), .ZN(n1935) );
XNOR2_X1 U1634 ( .A(n1974), .B(n2019), .ZN(n2018) );
NAND2_X1 U1635 ( .A1(KEYINPUT13), .A2(n1984), .ZN(n2019) );
XOR2_X1 U1636 ( .A(n2020), .B(KEYINPUT34), .Z(n2017) );
NAND2_X1 U1637 ( .A1(n2021), .A2(n2022), .ZN(n2020) );
OR3_X1 U1638 ( .A1(n1974), .A2(n2016), .A3(KEYINPUT13), .ZN(n2022) );
NAND2_X1 U1639 ( .A1(n2014), .A2(KEYINPUT13), .ZN(n2021) );
NOR2_X1 U1640 ( .A1(n1985), .A2(n2016), .ZN(n2014) );
NOR2_X1 U1641 ( .A1(n1974), .A2(n1942), .ZN(n2009) );
INV_X1 U1642 ( .A(n1985), .ZN(n1974) );
NAND2_X1 U1643 ( .A1(n2023), .A2(n2024), .ZN(n1985) );
OR2_X1 U1644 ( .A1(n2025), .A2(n1994), .ZN(n2024) );
XOR2_X1 U1645 ( .A(n2026), .B(KEYINPUT26), .Z(n2023) );
NAND2_X1 U1646 ( .A1(n2025), .A2(n1994), .ZN(n2026) );
NAND2_X1 U1647 ( .A1(n2027), .A2(n2028), .ZN(n1994) );
NAND2_X1 U1648 ( .A1(n2029), .A2(n2030), .ZN(n2028) );
XOR2_X1 U1649 ( .A(KEYINPUT40), .B(n2031), .Z(n2027) );
NOR2_X1 U1650 ( .A1(n2032), .A2(n2033), .ZN(n2031) );
XNOR2_X1 U1651 ( .A(n2034), .B(n1995), .ZN(n2025) );
AND2_X1 U1652 ( .A1(n2035), .A2(n2036), .ZN(n1995) );
NAND2_X1 U1653 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1914), .ZN(n2036) );
XOR2_X1 U1654 ( .A(n2037), .B(KEYINPUT54), .Z(n2035) );
NAND2_X1 U1655 ( .A1(RESTART), .A2(RMIN_REG_3__SCAN_IN), .ZN(n2037) );
NAND2_X1 U1656 ( .A1(KEYINPUT5), .A2(n1999), .ZN(n2034) );
NAND2_X1 U1657 ( .A1(n2038), .A2(n2039), .ZN(n1999) );
NAND2_X1 U1658 ( .A1(DATA_IN_3_), .A2(n1914), .ZN(n2039) );
NAND2_X1 U1659 ( .A1(RESTART), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2038) );
NAND2_X1 U1660 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1763), .ZN(n2007) );
NAND2_X1 U1661 ( .A1(n1849), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2006) );
NAND2_X1 U1662 ( .A1(n1848), .A2(REG4_REG_2__SCAN_IN), .ZN(n2005) );
NAND4_X1 U1663 ( .A1(n2040), .A2(n2041), .A3(n2042), .A4(n2043), .ZN(U282));
NAND2_X1 U1664 ( .A1(n1849), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2043) );
NOR2_X1 U1665 ( .A1(n2044), .A2(n2045), .ZN(n2042) );
AND2_X1 U1666 ( .A1(n2046), .A2(n1896), .ZN(n2045) );
INV_X1 U1667 ( .A(n1942), .ZN(n1896) );
NOR3_X1 U1668 ( .A1(n2047), .A2(n2016), .A3(n2048), .ZN(n2044) );
AND2_X1 U1669 ( .A1(n2049), .A2(n2050), .ZN(n2016) );
NAND2_X1 U1670 ( .A1(n2051), .A2(n1984), .ZN(n2050) );
INV_X1 U1671 ( .A(n1973), .ZN(n1984) );
NOR2_X1 U1672 ( .A1(n2052), .A2(n2046), .ZN(n1973) );
NAND2_X1 U1673 ( .A1(n2046), .A2(n2052), .ZN(n2051) );
NOR2_X1 U1674 ( .A1(n2046), .A2(n2049), .ZN(n2047) );
XOR2_X1 U1675 ( .A(n2053), .B(n2033), .Z(n2046) );
NAND2_X1 U1676 ( .A1(n2054), .A2(n2055), .ZN(n2033) );
NAND2_X1 U1677 ( .A1(n2056), .A2(n2057), .ZN(n2055) );
NAND2_X1 U1678 ( .A1(n2058), .A2(n2059), .ZN(n2056) );
OR2_X1 U1679 ( .A1(n2058), .A2(n2059), .ZN(n2054) );
NAND4_X1 U1680 ( .A1(KEYINPUT6), .A2(n2060), .A3(n2061), .A4(n2062), .ZN(n2053) );
NAND3_X1 U1681 ( .A1(n2029), .A2(n2030), .A3(n2063), .ZN(n2062) );
OR2_X1 U1682 ( .A1(n2063), .A2(n2030), .ZN(n2061) );
INV_X1 U1683 ( .A(KEYINPUT21), .ZN(n2063) );
INV_X1 U1684 ( .A(n2032), .ZN(n2060) );
NOR2_X1 U1685 ( .A1(n2030), .A2(n2029), .ZN(n2032) );
NAND2_X1 U1686 ( .A1(n2064), .A2(n2065), .ZN(n2029) );
NAND2_X1 U1687 ( .A1(DATA_IN_2_), .A2(n1914), .ZN(n2065) );
NAND2_X1 U1688 ( .A1(RESTART), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2064) );
NAND2_X1 U1689 ( .A1(n2066), .A2(n2067), .ZN(n2030) );
NAND2_X1 U1690 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1914), .ZN(n2067) );
NAND2_X1 U1691 ( .A1(RESTART), .A2(RMIN_REG_2__SCAN_IN), .ZN(n2066) );
NAND2_X1 U1692 ( .A1(n1848), .A2(REG4_REG_1__SCAN_IN), .ZN(n2041) );
NAND2_X1 U1693 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1763), .ZN(n2040) );
NAND3_X1 U1694 ( .A1(n2068), .A2(n2069), .A3(n2070), .ZN(U281) );
NOR3_X1 U1695 ( .A1(n2071), .A2(n2072), .A3(n2073), .ZN(n2070) );
AND2_X1 U1696 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1849), .ZN(n2073) );
AND3_X1 U1697 ( .A1(n2074), .A2(n1914), .A3(n2075), .ZN(n1849) );
XNOR2_X1 U1698 ( .A(KEYINPUT58), .B(n1759), .ZN(n2074) );
INV_X1 U1699 ( .A(ENABLE), .ZN(n1759) );
NOR2_X1 U1700 ( .A1(n2048), .A2(n2049), .ZN(n2072) );
NAND2_X1 U1701 ( .A1(n2052), .A2(n2076), .ZN(n2049) );
NAND3_X1 U1702 ( .A1(n2077), .A2(n2057), .A3(n2078), .ZN(n2076) );
INV_X1 U1703 ( .A(n2079), .ZN(n2078) );
NAND2_X1 U1704 ( .A1(n2079), .A2(n2080), .ZN(n2052) );
NAND2_X1 U1705 ( .A1(n2077), .A2(n2057), .ZN(n2080) );
OR2_X1 U1706 ( .A1(n2081), .A2(n2082), .ZN(n2077) );
NOR2_X1 U1707 ( .A1(n1864), .A2(n1874), .ZN(n2048) );
NOR2_X1 U1708 ( .A1(n2083), .A2(n2084), .ZN(n1874) );
NOR3_X1 U1709 ( .A1(n2085), .A2(AVERAGE), .A3(n2086), .ZN(n1864) );
NOR2_X1 U1710 ( .A1(n2079), .A2(n1942), .ZN(n2071) );
NAND3_X1 U1711 ( .A1(n2087), .A2(n2083), .A3(n2075), .ZN(n1942) );
NAND3_X1 U1712 ( .A1(n2088), .A2(n2089), .A3(RESTART), .ZN(n2083) );
NAND3_X1 U1713 ( .A1(n2090), .A2(n2091), .A3(n2092), .ZN(n2089) );
XOR2_X1 U1714 ( .A(n2093), .B(KEYINPUT61), .Z(n2092) );
NAND2_X1 U1715 ( .A1(n1675), .A2(n2094), .ZN(n2093) );
NAND2_X1 U1716 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n2095), .ZN(n2094) );
INV_X1 U1717 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1675) );
NAND2_X1 U1718 ( .A1(n2096), .A2(n1736), .ZN(n2091) );
INV_X1 U1719 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1736) );
XNOR2_X1 U1720 ( .A(KEYINPUT17), .B(n2095), .ZN(n2096) );
NAND2_X1 U1721 ( .A1(n2097), .A2(n2098), .ZN(n2095) );
NAND2_X1 U1722 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n2099), .ZN(n2098) );
OR2_X1 U1723 ( .A1(n2100), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2099) );
NAND2_X1 U1724 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n2100), .ZN(n2097) );
XNOR2_X1 U1725 ( .A(n2101), .B(KEYINPUT18), .ZN(n2100) );
NAND2_X1 U1726 ( .A1(n2102), .A2(n2103), .ZN(n2101) );
NAND2_X1 U1727 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2103) );
NAND3_X1 U1728 ( .A1(n2104), .A2(n2105), .A3(n2106), .ZN(n2102) );
OR2_X1 U1729 ( .A1(RMAX_REG_4__SCAN_IN), .A2(RMIN_REG_4__SCAN_IN), .ZN(n2106) );
NAND3_X1 U1730 ( .A1(n2107), .A2(n2108), .A3(n2109), .ZN(n2105) );
NAND2_X1 U1731 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2109) );
NAND4_X1 U1732 ( .A1(n2110), .A2(n2111), .A3(n2112), .A4(n2113), .ZN(n2108));
NAND2_X1 U1733 ( .A1(KEYINPUT60), .A2(n2114), .ZN(n2113) );
NAND2_X1 U1734 ( .A1(n1696), .A2(n1734), .ZN(n2114) );
NAND2_X1 U1735 ( .A1(n2115), .A2(n1696), .ZN(n2112) );
INV_X1 U1736 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1696) );
NAND2_X1 U1737 ( .A1(n2116), .A2(n2117), .ZN(n2115) );
OR2_X1 U1738 ( .A1(KEYINPUT60), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2117) );
INV_X1 U1739 ( .A(n2118), .ZN(n2116) );
NAND2_X1 U1740 ( .A1(n2118), .A2(n1734), .ZN(n2111) );
INV_X1 U1741 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1734) );
NAND2_X1 U1742 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2118) );
NAND2_X1 U1743 ( .A1(n1727), .A2(n1699), .ZN(n2110) );
INV_X1 U1744 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1699) );
INV_X1 U1745 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1727) );
NAND2_X1 U1746 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2107) );
NAND2_X1 U1747 ( .A1(n1722), .A2(n1689), .ZN(n2104) );
INV_X1 U1748 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1689) );
INV_X1 U1749 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1722) );
NAND2_X1 U1750 ( .A1(n2119), .A2(RMIN_REG_7__SCAN_IN), .ZN(n2090) );
XNOR2_X1 U1751 ( .A(RMAX_REG_7__SCAN_IN), .B(KEYINPUT10), .ZN(n2119) );
NAND2_X1 U1752 ( .A1(n1709), .A2(n1703), .ZN(n2088) );
INV_X1 U1753 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1703) );
INV_X1 U1754 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1709) );
NAND2_X1 U1755 ( .A1(n1914), .A2(n2120), .ZN(n2087) );
NAND3_X1 U1756 ( .A1(n2085), .A2(n2121), .A3(ENABLE), .ZN(n2120) );
NAND2_X1 U1757 ( .A1(n2122), .A2(n2123), .ZN(n2085) );
NAND2_X1 U1758 ( .A1(n2124), .A2(n2125), .ZN(n2123) );
NAND2_X1 U1759 ( .A1(REG4_REG_7__SCAN_IN), .A2(DATA_IN_7_), .ZN(n2125) );
NAND2_X1 U1760 ( .A1(n2126), .A2(n2127), .ZN(n2124) );
NAND2_X1 U1761 ( .A1(REG4_REG_6__SCAN_IN), .A2(DATA_IN_6_), .ZN(n2127) );
NAND3_X1 U1762 ( .A1(n2128), .A2(n2129), .A3(n2130), .ZN(n2126) );
OR2_X1 U1763 ( .A1(DATA_IN_6_), .A2(REG4_REG_6__SCAN_IN), .ZN(n2130) );
NAND3_X1 U1764 ( .A1(n2131), .A2(n2132), .A3(n2133), .ZN(n2129) );
NAND2_X1 U1765 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2133) );
NAND3_X1 U1766 ( .A1(n2134), .A2(n2135), .A3(n2136), .ZN(n2132) );
NAND2_X1 U1767 ( .A1(n1700), .A2(n1830), .ZN(n2136) );
INV_X1 U1768 ( .A(REG4_REG_3__SCAN_IN), .ZN(n1830) );
INV_X1 U1769 ( .A(DATA_IN_3_), .ZN(n1700) );
NAND3_X1 U1770 ( .A1(n2137), .A2(n2138), .A3(n2139), .ZN(n2135) );
NAND2_X1 U1771 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2139) );
NAND3_X1 U1772 ( .A1(n2140), .A2(n2141), .A3(n2142), .ZN(n2138) );
OR2_X1 U1773 ( .A1(DATA_IN_2_), .A2(REG4_REG_2__SCAN_IN), .ZN(n2142) );
NAND2_X1 U1774 ( .A1(n2143), .A2(n2144), .ZN(n2141) );
INV_X1 U1775 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2144) );
OR2_X1 U1776 ( .A1(n2145), .A2(n1693), .ZN(n2143) );
NAND2_X1 U1777 ( .A1(n2145), .A2(n1693), .ZN(n2140) );
INV_X1 U1778 ( .A(DATA_IN_1_), .ZN(n1693) );
NAND2_X1 U1779 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2145) );
NAND2_X1 U1780 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2137) );
NAND2_X1 U1781 ( .A1(n2146), .A2(n2147), .ZN(n2134) );
INV_X1 U1782 ( .A(REG4_REG_4__SCAN_IN), .ZN(n2147) );
XOR2_X1 U1783 ( .A(KEYINPUT25), .B(DATA_IN_4_), .Z(n2146) );
NAND2_X1 U1784 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2131) );
NAND2_X1 U1785 ( .A1(n1654), .A2(n1883), .ZN(n2128) );
INV_X1 U1786 ( .A(REG4_REG_5__SCAN_IN), .ZN(n1883) );
INV_X1 U1787 ( .A(DATA_IN_5_), .ZN(n1654) );
NAND2_X1 U1788 ( .A1(n1705), .A2(n1847), .ZN(n2122) );
INV_X1 U1789 ( .A(REG4_REG_7__SCAN_IN), .ZN(n1847) );
INV_X1 U1790 ( .A(DATA_IN_7_), .ZN(n1705) );
XOR2_X1 U1791 ( .A(n2148), .B(n2059), .Z(n2079) );
NAND2_X1 U1792 ( .A1(n2149), .A2(n2150), .ZN(n2059) );
NAND2_X1 U1793 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1914), .ZN(n2150) );
NAND2_X1 U1794 ( .A1(RESTART), .A2(RMIN_REG_1__SCAN_IN), .ZN(n2149) );
NAND2_X1 U1795 ( .A1(n2151), .A2(KEYINPUT37), .ZN(n2148) );
XNOR2_X1 U1796 ( .A(n2057), .B(n2058), .ZN(n2151) );
NAND2_X1 U1797 ( .A1(n2152), .A2(n2153), .ZN(n2058) );
NAND2_X1 U1798 ( .A1(DATA_IN_1_), .A2(n1914), .ZN(n2153) );
NAND2_X1 U1799 ( .A1(RESTART), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2152) );
NAND2_X1 U1800 ( .A1(n2081), .A2(n2082), .ZN(n2057) );
NAND2_X1 U1801 ( .A1(n2154), .A2(n2155), .ZN(n2082) );
NAND2_X1 U1802 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1914), .ZN(n2155) );
NAND2_X1 U1803 ( .A1(RESTART), .A2(RMIN_REG_0__SCAN_IN), .ZN(n2154) );
NAND2_X1 U1804 ( .A1(n2156), .A2(n2157), .ZN(n2081) );
NAND2_X1 U1805 ( .A1(DATA_IN_0_), .A2(n1914), .ZN(n2157) );
NAND2_X1 U1806 ( .A1(RESTART), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2156) );
NAND2_X1 U1807 ( .A1(n1848), .A2(REG4_REG_0__SCAN_IN), .ZN(n2069) );
NOR2_X1 U1808 ( .A1(n2121), .A2(n2086), .ZN(n1848) );
NAND3_X1 U1809 ( .A1(n2075), .A2(n1914), .A3(ENABLE), .ZN(n2086) );
INV_X1 U1810 ( .A(n2084), .ZN(n2075) );
NAND2_X1 U1811 ( .A1(STATO_REG_1__SCAN_IN), .A2(U280), .ZN(n2084) );
INV_X1 U1812 ( .A(AVERAGE), .ZN(n2121) );
NAND2_X1 U1813 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1763), .ZN(n2068) );
NAND2_X1 U1814 ( .A1(n1837), .A2(n2158), .ZN(U280) );
OR2_X1 U1815 ( .A1(n1643), .A2(STATO_REG_1__SCAN_IN), .ZN(n2158) );
NAND2_X1 U1816 ( .A1(STATO_REG_1__SCAN_IN), .A2(n2159), .ZN(n1837) );
XNOR2_X1 U1817 ( .A(n1643), .B(KEYINPUT11), .ZN(n2159) );
INV_X1 U1818 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1643) );
endmodule


