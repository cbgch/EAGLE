//Key = 1111111101010010110000110101110110101100001101001000011011010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373;

XNOR2_X1 U742 ( .A(n1039), .B(n1040), .ZN(G9) );
XNOR2_X1 U743 ( .A(G107), .B(KEYINPUT38), .ZN(n1040) );
NOR2_X1 U744 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR3_X1 U745 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
NOR2_X1 U746 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U747 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U748 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
INV_X1 U749 ( .A(KEYINPUT40), .ZN(n1051) );
NOR4_X1 U750 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1050) );
NOR2_X1 U751 ( .A1(n1056), .A2(n1055), .ZN(n1048) );
NOR2_X1 U752 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U753 ( .A1(n1059), .A2(n1054), .ZN(n1058) );
NOR2_X1 U754 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR3_X1 U755 ( .A1(n1053), .A2(KEYINPUT40), .A3(n1052), .ZN(n1061) );
NOR3_X1 U756 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1060) );
XNOR2_X1 U757 ( .A(n1065), .B(KEYINPUT33), .ZN(n1062) );
NOR3_X1 U758 ( .A1(n1052), .A2(n1066), .A3(n1067), .ZN(n1057) );
NOR2_X1 U759 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NAND3_X1 U760 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1043) );
NAND3_X1 U761 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
INV_X1 U762 ( .A(n1055), .ZN(n1075) );
NAND2_X1 U763 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NAND4_X1 U764 ( .A1(n1063), .A2(n1078), .A3(n1064), .A4(n1065), .ZN(n1077) );
NAND2_X1 U765 ( .A1(n1079), .A2(n1080), .ZN(n1076) );
NAND2_X1 U766 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U767 ( .A1(n1065), .A2(n1083), .ZN(n1082) );
NAND3_X1 U768 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1083) );
NAND2_X1 U769 ( .A1(n1078), .A2(n1087), .ZN(n1085) );
OR3_X1 U770 ( .A1(n1088), .A2(n1089), .A3(n1087), .ZN(n1084) );
INV_X1 U771 ( .A(KEYINPUT16), .ZN(n1087) );
NAND2_X1 U772 ( .A1(n1090), .A2(n1078), .ZN(n1081) );
AND3_X1 U773 ( .A1(n1070), .A2(n1071), .A3(n1091), .ZN(n1041) );
NAND4_X1 U774 ( .A1(n1079), .A2(n1078), .A3(n1092), .A4(n1093), .ZN(n1070) );
NOR4_X1 U775 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1093) );
NOR2_X1 U776 ( .A1(n1098), .A2(n1099), .ZN(n1094) );
XOR2_X1 U777 ( .A(n1100), .B(KEYINPUT10), .Z(n1092) );
XOR2_X1 U778 ( .A(n1101), .B(n1102), .Z(G72) );
NOR2_X1 U779 ( .A1(n1103), .A2(n1071), .ZN(n1102) );
NOR2_X1 U780 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U781 ( .A1(n1106), .A2(n1107), .ZN(n1101) );
NAND2_X1 U782 ( .A1(n1108), .A2(n1071), .ZN(n1107) );
XNOR2_X1 U783 ( .A(n1109), .B(n1110), .ZN(n1108) );
NOR2_X1 U784 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
INV_X1 U785 ( .A(n1113), .ZN(n1112) );
XOR2_X1 U786 ( .A(n1114), .B(KEYINPUT23), .Z(n1111) );
NAND3_X1 U787 ( .A1(G900), .A2(n1109), .A3(G953), .ZN(n1106) );
XNOR2_X1 U788 ( .A(n1115), .B(n1116), .ZN(n1109) );
XNOR2_X1 U789 ( .A(n1117), .B(n1118), .ZN(n1116) );
NAND2_X1 U790 ( .A1(KEYINPUT32), .A2(n1119), .ZN(n1117) );
XOR2_X1 U791 ( .A(n1120), .B(n1121), .Z(n1115) );
NOR2_X1 U792 ( .A1(KEYINPUT51), .A2(n1122), .ZN(n1121) );
XNOR2_X1 U793 ( .A(G125), .B(G146), .ZN(n1120) );
XOR2_X1 U794 ( .A(n1123), .B(n1124), .Z(G69) );
NAND2_X1 U795 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
OR3_X1 U796 ( .A1(n1071), .A2(G224), .A3(n1127), .ZN(n1126) );
NAND2_X1 U797 ( .A1(n1128), .A2(n1127), .ZN(n1125) );
OR2_X1 U798 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
XNOR2_X1 U799 ( .A(n1131), .B(n1132), .ZN(n1129) );
XNOR2_X1 U800 ( .A(n1133), .B(n1134), .ZN(n1131) );
NAND2_X1 U801 ( .A1(KEYINPUT54), .A2(n1135), .ZN(n1133) );
INV_X1 U802 ( .A(n1136), .ZN(n1135) );
NAND2_X1 U803 ( .A1(G953), .A2(n1137), .ZN(n1128) );
NAND2_X1 U804 ( .A1(G898), .A2(G224), .ZN(n1137) );
NAND2_X1 U805 ( .A1(n1071), .A2(n1138), .ZN(n1123) );
NAND2_X1 U806 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XNOR2_X1 U807 ( .A(KEYINPUT9), .B(n1141), .ZN(n1140) );
NOR3_X1 U808 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(G66) );
AND2_X1 U809 ( .A1(KEYINPUT7), .A2(n1145), .ZN(n1144) );
NOR3_X1 U810 ( .A1(KEYINPUT7), .A2(n1071), .A3(n1091), .ZN(n1143) );
INV_X1 U811 ( .A(G952), .ZN(n1091) );
XOR2_X1 U812 ( .A(n1146), .B(n1147), .Z(n1142) );
NOR2_X1 U813 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
NOR2_X1 U814 ( .A1(n1145), .A2(n1150), .ZN(G63) );
XOR2_X1 U815 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U816 ( .A1(n1099), .A2(n1149), .ZN(n1151) );
NOR2_X1 U817 ( .A1(n1145), .A2(n1153), .ZN(G60) );
XNOR2_X1 U818 ( .A(n1154), .B(n1155), .ZN(n1153) );
AND2_X1 U819 ( .A1(G475), .A2(n1156), .ZN(n1155) );
XNOR2_X1 U820 ( .A(G104), .B(n1157), .ZN(G6) );
NAND2_X1 U821 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XNOR2_X1 U822 ( .A(KEYINPUT26), .B(n1160), .ZN(n1159) );
NOR2_X1 U823 ( .A1(n1145), .A2(n1161), .ZN(G57) );
XOR2_X1 U824 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U825 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
NOR2_X1 U826 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
INV_X1 U827 ( .A(n1168), .ZN(n1167) );
NOR2_X1 U828 ( .A1(n1169), .A2(n1168), .ZN(n1164) );
XOR2_X1 U829 ( .A(n1170), .B(n1171), .Z(n1168) );
XNOR2_X1 U830 ( .A(n1172), .B(n1173), .ZN(n1170) );
NAND2_X1 U831 ( .A1(KEYINPUT1), .A2(n1174), .ZN(n1172) );
XOR2_X1 U832 ( .A(KEYINPUT27), .B(n1166), .Z(n1169) );
AND2_X1 U833 ( .A1(n1156), .A2(G472), .ZN(n1166) );
NOR2_X1 U834 ( .A1(n1145), .A2(n1175), .ZN(G54) );
XOR2_X1 U835 ( .A(n1176), .B(n1177), .Z(n1175) );
AND2_X1 U836 ( .A1(G469), .A2(n1156), .ZN(n1176) );
NOR2_X1 U837 ( .A1(n1145), .A2(n1178), .ZN(G51) );
NOR2_X1 U838 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XOR2_X1 U839 ( .A(n1181), .B(KEYINPUT6), .Z(n1180) );
NAND2_X1 U840 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NOR2_X1 U841 ( .A1(n1182), .A2(n1183), .ZN(n1179) );
AND2_X1 U842 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NAND2_X1 U843 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
XNOR2_X1 U844 ( .A(n1188), .B(n1189), .ZN(n1186) );
XOR2_X1 U845 ( .A(n1190), .B(KEYINPUT21), .Z(n1184) );
NAND2_X1 U846 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XNOR2_X1 U847 ( .A(n1193), .B(n1188), .ZN(n1191) );
INV_X1 U848 ( .A(n1189), .ZN(n1193) );
AND2_X1 U849 ( .A1(n1156), .A2(n1194), .ZN(n1182) );
INV_X1 U850 ( .A(n1149), .ZN(n1156) );
NAND2_X1 U851 ( .A1(G902), .A2(n1045), .ZN(n1149) );
NAND4_X1 U852 ( .A1(n1113), .A2(n1139), .A3(n1114), .A4(n1141), .ZN(n1045) );
AND4_X1 U853 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1139) );
NOR4_X1 U854 ( .A1(n1199), .A2(n1200), .A3(n1039), .A4(n1201), .ZN(n1198) );
AND3_X1 U855 ( .A1(n1202), .A2(n1068), .A3(n1203), .ZN(n1201) );
AND2_X1 U856 ( .A1(n1068), .A2(n1158), .ZN(n1039) );
OR2_X1 U857 ( .A1(n1204), .A2(n1205), .ZN(n1197) );
NAND3_X1 U858 ( .A1(n1206), .A2(n1207), .A3(n1079), .ZN(n1196) );
NAND2_X1 U859 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U860 ( .A1(n1210), .A2(n1211), .ZN(n1206) );
NAND4_X1 U861 ( .A1(n1097), .A2(n1204), .A3(n1096), .A4(n1212), .ZN(n1211) );
NOR2_X1 U862 ( .A1(n1086), .A2(n1054), .ZN(n1212) );
INV_X1 U863 ( .A(KEYINPUT5), .ZN(n1204) );
NAND2_X1 U864 ( .A1(n1069), .A2(n1158), .ZN(n1195) );
AND2_X1 U865 ( .A1(n1213), .A2(n1065), .ZN(n1158) );
NOR4_X1 U866 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1113) );
OR3_X1 U867 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1217) );
NOR3_X1 U868 ( .A1(n1221), .A2(n1222), .A3(n1047), .ZN(n1220) );
INV_X1 U869 ( .A(KEYINPUT63), .ZN(n1221) );
NOR2_X1 U870 ( .A1(KEYINPUT63), .A2(n1223), .ZN(n1219) );
NOR2_X1 U871 ( .A1(n1224), .A2(n1086), .ZN(n1218) );
NOR2_X1 U872 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
NOR2_X1 U873 ( .A1(n1227), .A2(n1228), .ZN(n1225) );
AND3_X1 U874 ( .A1(n1069), .A2(n1229), .A3(n1090), .ZN(n1216) );
NAND2_X1 U875 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND3_X1 U876 ( .A1(n1232), .A2(n1233), .A3(n1079), .ZN(n1231) );
NAND2_X1 U877 ( .A1(n1234), .A2(n1078), .ZN(n1230) );
NOR2_X1 U878 ( .A1(n1071), .A2(G952), .ZN(n1145) );
XOR2_X1 U879 ( .A(G146), .B(n1215), .Z(G48) );
NOR3_X1 U880 ( .A1(n1160), .A2(n1086), .A3(n1228), .ZN(n1215) );
XNOR2_X1 U881 ( .A(n1235), .B(n1236), .ZN(G45) );
NOR2_X1 U882 ( .A1(n1086), .A2(n1237), .ZN(n1236) );
XNOR2_X1 U883 ( .A(n1226), .B(KEYINPUT60), .ZN(n1237) );
AND3_X1 U884 ( .A1(n1095), .A2(n1238), .A3(n1239), .ZN(n1226) );
XNOR2_X1 U885 ( .A(G140), .B(n1240), .ZN(G42) );
NAND4_X1 U886 ( .A1(n1241), .A2(n1090), .A3(n1069), .A4(n1234), .ZN(n1240) );
XNOR2_X1 U887 ( .A(n1078), .B(KEYINPUT36), .ZN(n1241) );
XOR2_X1 U888 ( .A(G137), .B(n1214), .Z(G39) );
NOR3_X1 U889 ( .A1(n1228), .A2(n1047), .A3(n1054), .ZN(n1214) );
INV_X1 U890 ( .A(n1073), .ZN(n1054) );
XNOR2_X1 U891 ( .A(n1242), .B(n1223), .ZN(G36) );
NAND2_X1 U892 ( .A1(n1222), .A2(n1078), .ZN(n1223) );
AND2_X1 U893 ( .A1(n1239), .A2(n1068), .ZN(n1222) );
NAND2_X1 U894 ( .A1(KEYINPUT4), .A2(n1243), .ZN(n1242) );
XNOR2_X1 U895 ( .A(G131), .B(n1114), .ZN(G33) );
NAND3_X1 U896 ( .A1(n1239), .A2(n1078), .A3(n1069), .ZN(n1114) );
INV_X1 U897 ( .A(n1047), .ZN(n1078) );
NAND2_X1 U898 ( .A1(n1244), .A2(n1088), .ZN(n1047) );
INV_X1 U899 ( .A(n1089), .ZN(n1244) );
AND2_X1 U900 ( .A1(n1202), .A2(n1234), .ZN(n1239) );
XOR2_X1 U901 ( .A(G128), .B(n1245), .Z(G30) );
NOR3_X1 U902 ( .A1(n1228), .A2(n1246), .A3(n1227), .ZN(n1245) );
XNOR2_X1 U903 ( .A(n1232), .B(KEYINPUT52), .ZN(n1246) );
NAND3_X1 U904 ( .A1(n1096), .A2(n1097), .A3(n1234), .ZN(n1228) );
NOR3_X1 U905 ( .A1(n1247), .A2(n1063), .A3(n1064), .ZN(n1234) );
INV_X1 U906 ( .A(n1248), .ZN(n1064) );
XOR2_X1 U907 ( .A(G101), .B(n1200), .Z(G3) );
AND3_X1 U908 ( .A1(n1202), .A2(n1213), .A3(n1073), .ZN(n1200) );
XNOR2_X1 U909 ( .A(n1249), .B(n1250), .ZN(G27) );
NOR4_X1 U910 ( .A1(n1251), .A2(n1086), .A3(KEYINPUT55), .A4(n1247), .ZN(n1250) );
INV_X1 U911 ( .A(n1233), .ZN(n1247) );
NAND2_X1 U912 ( .A1(n1055), .A2(n1252), .ZN(n1233) );
NAND4_X1 U913 ( .A1(G953), .A2(G902), .A3(n1253), .A4(n1105), .ZN(n1252) );
INV_X1 U914 ( .A(G900), .ZN(n1105) );
NAND3_X1 U915 ( .A1(n1069), .A2(n1079), .A3(n1090), .ZN(n1251) );
XOR2_X1 U916 ( .A(n1141), .B(n1254), .Z(G24) );
NAND2_X1 U917 ( .A1(KEYINPUT45), .A2(G122), .ZN(n1254) );
NAND4_X1 U918 ( .A1(n1203), .A2(n1065), .A3(n1095), .A4(n1238), .ZN(n1141) );
INV_X1 U919 ( .A(n1067), .ZN(n1065) );
NAND2_X1 U920 ( .A1(n1255), .A2(n1256), .ZN(n1067) );
XNOR2_X1 U921 ( .A(n1096), .B(KEYINPUT18), .ZN(n1255) );
NAND3_X1 U922 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(G21) );
NAND2_X1 U923 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND2_X1 U924 ( .A1(n1262), .A2(KEYINPUT2), .ZN(n1260) );
XOR2_X1 U925 ( .A(n1205), .B(KEYINPUT35), .Z(n1262) );
NAND3_X1 U926 ( .A1(KEYINPUT2), .A2(G119), .A3(n1205), .ZN(n1258) );
OR2_X1 U927 ( .A1(n1205), .A2(KEYINPUT2), .ZN(n1257) );
NAND4_X1 U928 ( .A1(n1073), .A2(n1203), .A3(n1096), .A4(n1097), .ZN(n1205) );
XNOR2_X1 U929 ( .A(G116), .B(n1263), .ZN(G18) );
NAND3_X1 U930 ( .A1(n1203), .A2(n1264), .A3(n1202), .ZN(n1263) );
XNOR2_X1 U931 ( .A(KEYINPUT50), .B(n1227), .ZN(n1264) );
INV_X1 U932 ( .A(n1068), .ZN(n1227) );
NOR2_X1 U933 ( .A1(n1095), .A2(n1265), .ZN(n1068) );
NOR3_X1 U934 ( .A1(n1086), .A2(n1210), .A3(n1052), .ZN(n1203) );
INV_X1 U935 ( .A(n1079), .ZN(n1052) );
INV_X1 U936 ( .A(n1232), .ZN(n1086) );
XNOR2_X1 U937 ( .A(n1266), .B(KEYINPUT46), .ZN(n1232) );
XOR2_X1 U938 ( .A(n1267), .B(n1268), .Z(G15) );
NOR3_X1 U939 ( .A1(n1208), .A2(n1210), .A3(n1269), .ZN(n1268) );
XNOR2_X1 U940 ( .A(n1079), .B(KEYINPUT49), .ZN(n1269) );
NOR2_X1 U941 ( .A1(n1248), .A2(n1063), .ZN(n1079) );
INV_X1 U942 ( .A(n1270), .ZN(n1063) );
INV_X1 U943 ( .A(n1209), .ZN(n1210) );
NAND3_X1 U944 ( .A1(n1271), .A2(n1202), .A3(n1069), .ZN(n1208) );
INV_X1 U945 ( .A(n1160), .ZN(n1069) );
NAND2_X1 U946 ( .A1(n1265), .A2(n1095), .ZN(n1160) );
INV_X1 U947 ( .A(n1238), .ZN(n1265) );
INV_X1 U948 ( .A(n1053), .ZN(n1202) );
NAND2_X1 U949 ( .A1(n1256), .A2(n1096), .ZN(n1053) );
XNOR2_X1 U950 ( .A(G113), .B(KEYINPUT3), .ZN(n1267) );
NAND3_X1 U951 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(G12) );
NAND2_X1 U952 ( .A1(n1199), .A2(n1275), .ZN(n1274) );
NAND2_X1 U953 ( .A1(KEYINPUT28), .A2(n1276), .ZN(n1275) );
XOR2_X1 U954 ( .A(KEYINPUT39), .B(G110), .Z(n1276) );
INV_X1 U955 ( .A(n1277), .ZN(n1199) );
NAND3_X1 U956 ( .A1(KEYINPUT28), .A2(n1277), .A3(G110), .ZN(n1273) );
NAND3_X1 U957 ( .A1(n1073), .A2(n1213), .A3(n1090), .ZN(n1277) );
NOR2_X1 U958 ( .A1(n1096), .A2(n1256), .ZN(n1090) );
INV_X1 U959 ( .A(n1097), .ZN(n1256) );
XOR2_X1 U960 ( .A(n1278), .B(n1148), .Z(n1097) );
NAND2_X1 U961 ( .A1(G217), .A2(n1279), .ZN(n1148) );
OR2_X1 U962 ( .A1(n1147), .A2(n1280), .ZN(n1278) );
XNOR2_X1 U963 ( .A(n1281), .B(n1282), .ZN(n1147) );
XOR2_X1 U964 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U965 ( .A(KEYINPUT25), .B(n1285), .Z(n1284) );
NOR2_X1 U966 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U967 ( .A(n1288), .B(KEYINPUT34), .Z(n1287) );
NAND2_X1 U968 ( .A1(G110), .A2(n1289), .ZN(n1288) );
NOR2_X1 U969 ( .A1(G110), .A2(n1289), .ZN(n1286) );
XNOR2_X1 U970 ( .A(G128), .B(n1261), .ZN(n1289) );
AND2_X1 U971 ( .A1(n1290), .A2(G221), .ZN(n1283) );
XNOR2_X1 U972 ( .A(n1291), .B(n1292), .ZN(n1281) );
XNOR2_X1 U973 ( .A(n1293), .B(G472), .ZN(n1096) );
NAND2_X1 U974 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
XOR2_X1 U975 ( .A(n1296), .B(n1297), .Z(n1294) );
XNOR2_X1 U976 ( .A(n1174), .B(n1163), .ZN(n1297) );
XNOR2_X1 U977 ( .A(n1298), .B(n1299), .ZN(n1163) );
NAND2_X1 U978 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
XOR2_X1 U979 ( .A(KEYINPUT24), .B(G210), .Z(n1301) );
INV_X1 U980 ( .A(n1119), .ZN(n1174) );
XOR2_X1 U981 ( .A(n1302), .B(n1303), .Z(n1296) );
NOR2_X1 U982 ( .A1(KEYINPUT62), .A2(n1171), .ZN(n1303) );
XOR2_X1 U983 ( .A(n1304), .B(n1305), .Z(n1171) );
XNOR2_X1 U984 ( .A(G113), .B(G119), .ZN(n1304) );
XNOR2_X1 U985 ( .A(KEYINPUT12), .B(n1306), .ZN(n1302) );
NOR2_X1 U986 ( .A1(KEYINPUT44), .A2(n1173), .ZN(n1306) );
AND4_X1 U987 ( .A1(n1271), .A2(n1248), .A3(n1209), .A4(n1270), .ZN(n1213) );
NAND2_X1 U988 ( .A1(G221), .A2(n1279), .ZN(n1270) );
NAND2_X1 U989 ( .A1(G234), .A2(n1307), .ZN(n1279) );
NAND2_X1 U990 ( .A1(n1055), .A2(n1308), .ZN(n1209) );
NAND3_X1 U991 ( .A1(G902), .A2(n1253), .A3(n1130), .ZN(n1308) );
NOR2_X1 U992 ( .A1(n1071), .A2(G898), .ZN(n1130) );
NAND3_X1 U993 ( .A1(n1253), .A2(n1071), .A3(G952), .ZN(n1055) );
NAND2_X1 U994 ( .A1(G237), .A2(G234), .ZN(n1253) );
XNOR2_X1 U995 ( .A(n1309), .B(G469), .ZN(n1248) );
OR2_X1 U996 ( .A1(n1177), .A2(n1280), .ZN(n1309) );
XNOR2_X1 U997 ( .A(n1310), .B(n1311), .ZN(n1177) );
XOR2_X1 U998 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U999 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1000 ( .A(n1316), .B(n1317), .Z(n1310) );
XOR2_X1 U1001 ( .A(KEYINPUT56), .B(G110), .Z(n1317) );
XNOR2_X1 U1002 ( .A(n1119), .B(n1318), .ZN(n1316) );
NOR2_X1 U1003 ( .A1(G953), .A2(n1104), .ZN(n1318) );
INV_X1 U1004 ( .A(G227), .ZN(n1104) );
XNOR2_X1 U1005 ( .A(n1319), .B(n1320), .ZN(n1119) );
XNOR2_X1 U1006 ( .A(KEYINPUT17), .B(n1243), .ZN(n1320) );
INV_X1 U1007 ( .A(G134), .ZN(n1243) );
XNOR2_X1 U1008 ( .A(G131), .B(n1292), .ZN(n1319) );
XOR2_X1 U1009 ( .A(G137), .B(KEYINPUT15), .Z(n1292) );
XOR2_X1 U1010 ( .A(n1266), .B(KEYINPUT22), .Z(n1271) );
NAND2_X1 U1011 ( .A1(n1089), .A2(n1088), .ZN(n1266) );
NAND2_X1 U1012 ( .A1(G214), .A2(n1321), .ZN(n1088) );
XNOR2_X1 U1013 ( .A(n1322), .B(n1194), .ZN(n1089) );
AND2_X1 U1014 ( .A1(G210), .A2(n1321), .ZN(n1194) );
NAND2_X1 U1015 ( .A1(n1323), .A2(n1307), .ZN(n1321) );
INV_X1 U1016 ( .A(G902), .ZN(n1307) );
INV_X1 U1017 ( .A(G237), .ZN(n1323) );
NAND2_X1 U1018 ( .A1(n1324), .A2(n1295), .ZN(n1322) );
XOR2_X1 U1019 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1020 ( .A(n1327), .B(n1328), .Z(n1326) );
NOR2_X1 U1021 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
AND2_X1 U1022 ( .A1(KEYINPUT43), .A2(n1188), .ZN(n1330) );
XOR2_X1 U1023 ( .A(n1173), .B(G125), .Z(n1188) );
INV_X1 U1024 ( .A(n1331), .ZN(n1173) );
NOR3_X1 U1025 ( .A1(KEYINPUT43), .A2(n1331), .A3(n1249), .ZN(n1329) );
INV_X1 U1026 ( .A(G125), .ZN(n1249) );
XOR2_X1 U1027 ( .A(G128), .B(n1332), .Z(n1331) );
NOR2_X1 U1028 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
NOR2_X1 U1029 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
INV_X1 U1030 ( .A(n1337), .ZN(n1336) );
XOR2_X1 U1031 ( .A(KEYINPUT42), .B(n1338), .Z(n1335) );
NOR2_X1 U1032 ( .A1(n1337), .A2(n1338), .ZN(n1333) );
XNOR2_X1 U1033 ( .A(n1235), .B(KEYINPUT11), .ZN(n1338) );
XOR2_X1 U1034 ( .A(G146), .B(KEYINPUT57), .Z(n1337) );
NOR2_X1 U1035 ( .A1(KEYINPUT19), .A2(n1339), .ZN(n1327) );
XNOR2_X1 U1036 ( .A(n1192), .B(KEYINPUT14), .ZN(n1339) );
INV_X1 U1037 ( .A(n1187), .ZN(n1192) );
NAND2_X1 U1038 ( .A1(n1340), .A2(n1341), .ZN(n1187) );
NAND2_X1 U1039 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
INV_X1 U1040 ( .A(n1134), .ZN(n1343) );
XNOR2_X1 U1041 ( .A(n1132), .B(n1344), .ZN(n1342) );
XOR2_X1 U1042 ( .A(n1345), .B(KEYINPUT41), .Z(n1340) );
NAND2_X1 U1043 ( .A1(n1346), .A2(n1134), .ZN(n1345) );
XNOR2_X1 U1044 ( .A(G122), .B(G110), .ZN(n1134) );
XNOR2_X1 U1045 ( .A(n1344), .B(n1347), .ZN(n1346) );
INV_X1 U1046 ( .A(n1132), .ZN(n1347) );
XOR2_X1 U1047 ( .A(G113), .B(n1348), .Z(n1132) );
NOR2_X1 U1048 ( .A1(KEYINPUT8), .A2(n1349), .ZN(n1348) );
XOR2_X1 U1049 ( .A(n1350), .B(n1305), .Z(n1349) );
NAND2_X1 U1050 ( .A1(KEYINPUT29), .A2(n1261), .ZN(n1350) );
INV_X1 U1051 ( .A(G119), .ZN(n1261) );
XNOR2_X1 U1052 ( .A(KEYINPUT53), .B(n1351), .ZN(n1344) );
NOR2_X1 U1053 ( .A1(KEYINPUT58), .A2(n1136), .ZN(n1351) );
XNOR2_X1 U1054 ( .A(n1312), .B(n1352), .ZN(n1136) );
XNOR2_X1 U1055 ( .A(KEYINPUT13), .B(n1353), .ZN(n1352) );
INV_X1 U1056 ( .A(G107), .ZN(n1353) );
XNOR2_X1 U1057 ( .A(G104), .B(n1299), .ZN(n1312) );
XOR2_X1 U1058 ( .A(G101), .B(KEYINPUT31), .Z(n1299) );
XNOR2_X1 U1059 ( .A(KEYINPUT47), .B(n1189), .ZN(n1325) );
NAND2_X1 U1060 ( .A1(G224), .A2(n1071), .ZN(n1189) );
NOR2_X1 U1061 ( .A1(n1238), .A2(n1095), .ZN(n1073) );
XNOR2_X1 U1062 ( .A(n1354), .B(G475), .ZN(n1095) );
NAND2_X1 U1063 ( .A1(n1295), .A2(n1154), .ZN(n1354) );
NAND2_X1 U1064 ( .A1(n1355), .A2(n1356), .ZN(n1154) );
NAND2_X1 U1065 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
XOR2_X1 U1066 ( .A(n1359), .B(KEYINPUT30), .Z(n1355) );
OR2_X1 U1067 ( .A1(n1358), .A2(n1357), .ZN(n1359) );
XOR2_X1 U1068 ( .A(n1360), .B(n1361), .Z(n1357) );
XOR2_X1 U1069 ( .A(n1362), .B(n1363), .Z(n1361) );
NAND2_X1 U1070 ( .A1(KEYINPUT59), .A2(n1364), .ZN(n1363) );
XNOR2_X1 U1071 ( .A(KEYINPUT61), .B(n1365), .ZN(n1364) );
INV_X1 U1072 ( .A(n1291), .ZN(n1365) );
XOR2_X1 U1073 ( .A(G125), .B(n1315), .Z(n1291) );
XNOR2_X1 U1074 ( .A(n1122), .B(G146), .ZN(n1315) );
INV_X1 U1075 ( .A(G140), .ZN(n1122) );
NAND2_X1 U1076 ( .A1(G214), .A2(n1300), .ZN(n1362) );
NOR2_X1 U1077 ( .A1(G953), .A2(G237), .ZN(n1300) );
XNOR2_X1 U1078 ( .A(n1366), .B(n1367), .ZN(n1360) );
NAND2_X1 U1079 ( .A1(KEYINPUT37), .A2(G131), .ZN(n1367) );
NAND2_X1 U1080 ( .A1(KEYINPUT0), .A2(n1235), .ZN(n1366) );
XOR2_X1 U1081 ( .A(G104), .B(n1368), .Z(n1358) );
XOR2_X1 U1082 ( .A(G122), .B(G113), .Z(n1368) );
INV_X1 U1083 ( .A(n1280), .ZN(n1295) );
NAND2_X1 U1084 ( .A1(n1100), .A2(n1369), .ZN(n1238) );
OR2_X1 U1085 ( .A1(n1099), .A2(n1098), .ZN(n1369) );
NAND2_X1 U1086 ( .A1(n1098), .A2(n1099), .ZN(n1100) );
INV_X1 U1087 ( .A(G478), .ZN(n1099) );
NOR2_X1 U1088 ( .A1(n1280), .A2(n1152), .ZN(n1098) );
XNOR2_X1 U1089 ( .A(n1370), .B(n1371), .ZN(n1152) );
XOR2_X1 U1090 ( .A(n1372), .B(n1373), .Z(n1371) );
XNOR2_X1 U1091 ( .A(G134), .B(G122), .ZN(n1373) );
NAND2_X1 U1092 ( .A1(G217), .A2(n1290), .ZN(n1372) );
AND2_X1 U1093 ( .A1(G234), .A2(n1071), .ZN(n1290) );
INV_X1 U1094 ( .A(G953), .ZN(n1071) );
XOR2_X1 U1095 ( .A(n1314), .B(n1305), .Z(n1370) );
XOR2_X1 U1096 ( .A(G116), .B(KEYINPUT48), .Z(n1305) );
XNOR2_X1 U1097 ( .A(G107), .B(n1118), .ZN(n1314) );
XNOR2_X1 U1098 ( .A(G128), .B(n1235), .ZN(n1118) );
INV_X1 U1099 ( .A(G143), .ZN(n1235) );
XOR2_X1 U1100 ( .A(G902), .B(KEYINPUT20), .Z(n1280) );
OR2_X1 U1101 ( .A1(G110), .A2(KEYINPUT28), .ZN(n1272) );
endmodule


