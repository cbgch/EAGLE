//Key = 1100010001100101101010011001100111101001011011011011100100101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370;

XNOR2_X1 U741 ( .A(G107), .B(n1024), .ZN(G9) );
NAND2_X1 U742 ( .A1(KEYINPUT31), .A2(n1025), .ZN(n1024) );
NOR2_X1 U743 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR4_X1 U744 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1027) );
NOR2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR2_X1 U746 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U747 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR2_X1 U748 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U749 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR3_X1 U750 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1040) );
NOR2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U752 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U753 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR3_X1 U754 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1043) );
XOR2_X1 U755 ( .A(n1054), .B(KEYINPUT11), .Z(n1053) );
NOR2_X1 U756 ( .A1(n1054), .A2(n1055), .ZN(n1042) );
NOR3_X1 U757 ( .A1(n1054), .A2(n1056), .A3(n1046), .ZN(n1038) );
NOR2_X1 U758 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR4_X1 U760 ( .A1(n1061), .A2(n1046), .A3(n1041), .A4(n1054), .ZN(n1034) );
NOR2_X1 U761 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND3_X1 U762 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1028) );
NOR3_X1 U763 ( .A1(n1067), .A2(G953), .A3(G952), .ZN(n1026) );
INV_X1 U764 ( .A(n1064), .ZN(n1067) );
NAND4_X1 U765 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1064) );
NOR3_X1 U766 ( .A1(n1054), .A2(n1072), .A3(n1073), .ZN(n1071) );
NOR3_X1 U767 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1070) );
NOR2_X1 U768 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XNOR2_X1 U769 ( .A(G469), .B(KEYINPUT12), .ZN(n1078) );
INV_X1 U770 ( .A(n1079), .ZN(n1077) );
NOR2_X1 U771 ( .A1(G469), .A2(n1079), .ZN(n1075) );
XOR2_X1 U772 ( .A(n1080), .B(n1081), .Z(n1074) );
XNOR2_X1 U773 ( .A(KEYINPUT60), .B(n1082), .ZN(n1081) );
NOR2_X1 U774 ( .A1(n1083), .A2(KEYINPUT38), .ZN(n1080) );
NAND2_X1 U775 ( .A1(KEYINPUT20), .A2(n1037), .ZN(n1069) );
NAND2_X1 U776 ( .A1(n1084), .A2(n1085), .ZN(n1068) );
INV_X1 U777 ( .A(KEYINPUT20), .ZN(n1085) );
NAND2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
XOR2_X1 U779 ( .A(n1088), .B(n1089), .Z(G72) );
XOR2_X1 U780 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND3_X1 U781 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
NAND2_X1 U782 ( .A1(G953), .A2(n1095), .ZN(n1094) );
XNOR2_X1 U783 ( .A(KEYINPUT15), .B(n1096), .ZN(n1095) );
NAND2_X1 U784 ( .A1(n1097), .A2(n1098), .ZN(n1093) );
NAND3_X1 U785 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
NAND2_X1 U786 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NAND2_X1 U787 ( .A1(n1104), .A2(G125), .ZN(n1099) );
NAND2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(n1092) );
INV_X1 U789 ( .A(n1097), .ZN(n1106) );
XNOR2_X1 U790 ( .A(n1102), .B(n1104), .ZN(n1105) );
NOR2_X1 U791 ( .A1(n1103), .A2(n1107), .ZN(n1104) );
INV_X1 U792 ( .A(KEYINPUT52), .ZN(n1103) );
INV_X1 U793 ( .A(G125), .ZN(n1102) );
NAND3_X1 U794 ( .A1(G953), .A2(n1108), .A3(KEYINPUT42), .ZN(n1090) );
XOR2_X1 U795 ( .A(KEYINPUT58), .B(n1109), .Z(n1108) );
AND2_X1 U796 ( .A1(G227), .A2(G900), .ZN(n1109) );
NOR2_X1 U797 ( .A1(n1110), .A2(G953), .ZN(n1088) );
XOR2_X1 U798 ( .A(n1111), .B(n1112), .Z(G69) );
NOR3_X1 U799 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1112) );
NOR2_X1 U800 ( .A1(G953), .A2(n1116), .ZN(n1115) );
NOR2_X1 U801 ( .A1(n1031), .A2(n1117), .ZN(n1116) );
XNOR2_X1 U802 ( .A(KEYINPUT35), .B(n1066), .ZN(n1117) );
NOR2_X1 U803 ( .A1(G224), .A2(n1065), .ZN(n1114) );
OR2_X1 U804 ( .A1(n1118), .A2(n1113), .ZN(n1111) );
NOR2_X1 U805 ( .A1(n1119), .A2(n1120), .ZN(G66) );
XOR2_X1 U806 ( .A(n1121), .B(n1122), .Z(n1120) );
NAND2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
NOR2_X1 U808 ( .A1(n1119), .A2(n1125), .ZN(G63) );
XOR2_X1 U809 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U810 ( .A1(n1123), .A2(G478), .ZN(n1126) );
NOR2_X1 U811 ( .A1(n1119), .A2(n1128), .ZN(G60) );
XOR2_X1 U812 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND3_X1 U813 ( .A1(KEYINPUT24), .A2(n1123), .A3(n1131), .ZN(n1129) );
XNOR2_X1 U814 ( .A(G475), .B(KEYINPUT32), .ZN(n1131) );
XNOR2_X1 U815 ( .A(G104), .B(n1132), .ZN(G6) );
NOR2_X1 U816 ( .A1(n1133), .A2(KEYINPUT40), .ZN(n1132) );
INV_X1 U817 ( .A(n1134), .ZN(n1133) );
NOR2_X1 U818 ( .A1(n1119), .A2(n1135), .ZN(G57) );
XOR2_X1 U819 ( .A(n1136), .B(n1137), .Z(n1135) );
NOR2_X1 U820 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
XOR2_X1 U821 ( .A(KEYINPUT53), .B(n1140), .Z(n1139) );
NOR2_X1 U822 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
AND2_X1 U823 ( .A1(n1142), .A2(n1141), .ZN(n1138) );
NAND2_X1 U824 ( .A1(n1123), .A2(G472), .ZN(n1142) );
NAND2_X1 U825 ( .A1(n1143), .A2(n1144), .ZN(n1136) );
XOR2_X1 U826 ( .A(n1145), .B(KEYINPUT30), .Z(n1143) );
OR2_X1 U827 ( .A1(G101), .A2(n1146), .ZN(n1145) );
NOR2_X1 U828 ( .A1(n1119), .A2(n1147), .ZN(G54) );
XOR2_X1 U829 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U830 ( .A(n1150), .B(n1151), .ZN(n1149) );
NOR2_X1 U831 ( .A1(KEYINPUT46), .A2(n1152), .ZN(n1150) );
XNOR2_X1 U832 ( .A(n1097), .B(n1153), .ZN(n1152) );
XOR2_X1 U833 ( .A(n1154), .B(KEYINPUT45), .Z(n1153) );
XOR2_X1 U834 ( .A(n1155), .B(n1156), .Z(n1097) );
XOR2_X1 U835 ( .A(n1157), .B(n1158), .Z(n1148) );
NAND2_X1 U836 ( .A1(n1123), .A2(G469), .ZN(n1157) );
INV_X1 U837 ( .A(n1159), .ZN(n1123) );
NOR2_X1 U838 ( .A1(n1160), .A2(n1161), .ZN(G51) );
XNOR2_X1 U839 ( .A(n1119), .B(KEYINPUT51), .ZN(n1161) );
NOR2_X1 U840 ( .A1(n1065), .A2(G952), .ZN(n1119) );
NOR3_X1 U841 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1160) );
AND2_X1 U842 ( .A1(n1165), .A2(KEYINPUT21), .ZN(n1164) );
NOR3_X1 U843 ( .A1(n1165), .A2(KEYINPUT21), .A3(n1166), .ZN(n1163) );
NOR3_X1 U844 ( .A1(n1159), .A2(KEYINPUT7), .A3(n1167), .ZN(n1166) );
NOR3_X1 U845 ( .A1(n1159), .A2(n1168), .A3(n1167), .ZN(n1162) );
NOR2_X1 U846 ( .A1(n1169), .A2(KEYINPUT21), .ZN(n1168) );
NOR2_X1 U847 ( .A1(KEYINPUT7), .A2(n1170), .ZN(n1169) );
INV_X1 U848 ( .A(n1165), .ZN(n1170) );
XOR2_X1 U849 ( .A(n1118), .B(n1171), .Z(n1165) );
NOR2_X1 U850 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NOR2_X1 U851 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XNOR2_X1 U852 ( .A(n1176), .B(KEYINPUT18), .ZN(n1175) );
INV_X1 U853 ( .A(n1177), .ZN(n1174) );
NOR2_X1 U854 ( .A1(n1177), .A2(n1178), .ZN(n1172) );
NAND2_X1 U855 ( .A1(G902), .A2(n1179), .ZN(n1159) );
NAND3_X1 U856 ( .A1(n1180), .A2(n1066), .A3(n1110), .ZN(n1179) );
INV_X1 U857 ( .A(n1029), .ZN(n1110) );
NAND4_X1 U858 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1029) );
NOR4_X1 U859 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1184) );
NOR3_X1 U860 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1188) );
INV_X1 U861 ( .A(n1192), .ZN(n1187) );
NOR2_X1 U862 ( .A1(n1193), .A2(n1194), .ZN(n1183) );
NAND4_X1 U863 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1182) );
XNOR2_X1 U864 ( .A(n1190), .B(KEYINPUT43), .ZN(n1198) );
XNOR2_X1 U865 ( .A(n1048), .B(KEYINPUT55), .ZN(n1195) );
INV_X1 U866 ( .A(n1031), .ZN(n1180) );
NAND4_X1 U867 ( .A1(n1134), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1031) );
NOR4_X1 U868 ( .A1(n1202), .A2(n1203), .A3(n1025), .A4(n1204), .ZN(n1201) );
AND2_X1 U869 ( .A1(n1205), .A2(n1063), .ZN(n1025) );
NAND2_X1 U870 ( .A1(n1206), .A2(n1058), .ZN(n1200) );
XOR2_X1 U871 ( .A(n1207), .B(KEYINPUT33), .Z(n1206) );
NAND2_X1 U872 ( .A1(n1208), .A2(n1048), .ZN(n1207) );
NAND2_X1 U873 ( .A1(n1062), .A2(n1205), .ZN(n1134) );
NOR4_X1 U874 ( .A1(n1055), .A2(n1054), .A3(n1190), .A4(n1209), .ZN(n1205) );
XNOR2_X1 U875 ( .A(n1156), .B(n1210), .ZN(G48) );
NOR3_X1 U876 ( .A1(n1211), .A2(n1191), .A3(n1189), .ZN(n1210) );
INV_X1 U877 ( .A(n1062), .ZN(n1191) );
XNOR2_X1 U878 ( .A(n1190), .B(KEYINPUT50), .ZN(n1211) );
NAND2_X1 U879 ( .A1(n1212), .A2(n1213), .ZN(G45) );
NAND2_X1 U880 ( .A1(G143), .A2(n1214), .ZN(n1213) );
XOR2_X1 U881 ( .A(KEYINPUT27), .B(n1215), .Z(n1212) );
NOR2_X1 U882 ( .A1(G143), .A2(n1214), .ZN(n1215) );
NAND4_X1 U883 ( .A1(n1216), .A2(n1048), .A3(n1197), .A4(n1196), .ZN(n1214) );
NOR2_X1 U884 ( .A1(n1086), .A2(n1217), .ZN(n1197) );
XNOR2_X1 U885 ( .A(KEYINPUT16), .B(n1058), .ZN(n1216) );
XNOR2_X1 U886 ( .A(n1107), .B(n1218), .ZN(G42) );
NOR2_X1 U887 ( .A1(KEYINPUT37), .A2(n1192), .ZN(n1218) );
NAND3_X1 U888 ( .A1(n1062), .A2(n1196), .A3(n1219), .ZN(n1192) );
NOR3_X1 U889 ( .A1(n1041), .A2(n1049), .A3(n1050), .ZN(n1219) );
XOR2_X1 U890 ( .A(n1186), .B(n1220), .Z(G39) );
NOR2_X1 U891 ( .A1(KEYINPUT25), .A2(n1221), .ZN(n1220) );
NOR3_X1 U892 ( .A1(n1037), .A2(n1041), .A3(n1189), .ZN(n1186) );
XOR2_X1 U893 ( .A(G134), .B(n1194), .Z(G36) );
AND2_X1 U894 ( .A1(n1222), .A2(n1063), .ZN(n1194) );
XOR2_X1 U895 ( .A(G131), .B(n1193), .Z(G33) );
AND2_X1 U896 ( .A1(n1222), .A2(n1062), .ZN(n1193) );
AND3_X1 U897 ( .A1(n1196), .A2(n1223), .A3(n1048), .ZN(n1222) );
XOR2_X1 U898 ( .A(G128), .B(n1185), .Z(G30) );
NOR3_X1 U899 ( .A1(n1224), .A2(n1190), .A3(n1189), .ZN(n1185) );
NAND3_X1 U900 ( .A1(n1050), .A2(n1225), .A3(n1196), .ZN(n1189) );
AND2_X1 U901 ( .A1(n1226), .A2(n1227), .ZN(n1196) );
INV_X1 U902 ( .A(n1063), .ZN(n1224) );
XOR2_X1 U903 ( .A(n1228), .B(n1229), .Z(G3) );
XNOR2_X1 U904 ( .A(G101), .B(KEYINPUT14), .ZN(n1229) );
NAND4_X1 U905 ( .A1(n1230), .A2(n1048), .A3(n1231), .A4(n1232), .ZN(n1228) );
NOR2_X1 U906 ( .A1(n1209), .A2(n1190), .ZN(n1231) );
XNOR2_X1 U907 ( .A(n1226), .B(KEYINPUT10), .ZN(n1230) );
XNOR2_X1 U908 ( .A(G125), .B(n1181), .ZN(G27) );
NAND4_X1 U909 ( .A1(n1233), .A2(n1062), .A3(n1234), .A4(n1227), .ZN(n1181) );
NAND2_X1 U910 ( .A1(n1033), .A2(n1235), .ZN(n1227) );
NAND4_X1 U911 ( .A1(G902), .A2(G953), .A3(n1236), .A4(n1096), .ZN(n1235) );
INV_X1 U912 ( .A(G900), .ZN(n1096) );
NAND2_X1 U913 ( .A1(n1237), .A2(n1238), .ZN(G24) );
OR2_X1 U914 ( .A1(n1199), .A2(G122), .ZN(n1238) );
XOR2_X1 U915 ( .A(n1239), .B(KEYINPUT8), .Z(n1237) );
NAND2_X1 U916 ( .A1(G122), .A2(n1199), .ZN(n1239) );
OR4_X1 U917 ( .A1(n1240), .A2(n1054), .A3(n1217), .A4(n1086), .ZN(n1199) );
XNOR2_X1 U918 ( .A(KEYINPUT29), .B(n1087), .ZN(n1217) );
NAND2_X1 U919 ( .A1(n1049), .A2(n1241), .ZN(n1054) );
NAND2_X1 U920 ( .A1(n1242), .A2(n1243), .ZN(G21) );
NAND2_X1 U921 ( .A1(n1203), .A2(n1244), .ZN(n1243) );
XOR2_X1 U922 ( .A(KEYINPUT47), .B(n1245), .Z(n1242) );
NOR2_X1 U923 ( .A1(n1203), .A2(n1244), .ZN(n1245) );
NOR4_X1 U924 ( .A1(n1240), .A2(n1037), .A3(n1241), .A4(n1049), .ZN(n1203) );
INV_X1 U925 ( .A(n1246), .ZN(n1240) );
XNOR2_X1 U926 ( .A(G116), .B(n1066), .ZN(G18) );
NAND3_X1 U927 ( .A1(n1048), .A2(n1063), .A3(n1246), .ZN(n1066) );
NAND2_X1 U928 ( .A1(n1247), .A2(n1248), .ZN(n1063) );
NAND3_X1 U929 ( .A1(n1087), .A2(n1086), .A3(n1249), .ZN(n1248) );
INV_X1 U930 ( .A(KEYINPUT29), .ZN(n1249) );
NAND2_X1 U931 ( .A1(KEYINPUT29), .A2(n1232), .ZN(n1247) );
XOR2_X1 U932 ( .A(G113), .B(n1202), .Z(G15) );
AND3_X1 U933 ( .A1(n1062), .A2(n1048), .A3(n1246), .ZN(n1202) );
NOR3_X1 U934 ( .A1(n1190), .A2(n1209), .A3(n1046), .ZN(n1246) );
INV_X1 U935 ( .A(n1234), .ZN(n1046) );
NAND2_X1 U936 ( .A1(n1250), .A2(n1251), .ZN(n1234) );
OR3_X1 U937 ( .A1(n1052), .A2(n1073), .A3(KEYINPUT4), .ZN(n1251) );
INV_X1 U938 ( .A(n1051), .ZN(n1073) );
NAND2_X1 U939 ( .A1(KEYINPUT4), .A2(n1226), .ZN(n1250) );
INV_X1 U940 ( .A(n1055), .ZN(n1226) );
NOR2_X1 U941 ( .A1(n1225), .A2(n1241), .ZN(n1048) );
INV_X1 U942 ( .A(n1050), .ZN(n1241) );
NOR2_X1 U943 ( .A1(n1087), .A2(n1086), .ZN(n1062) );
INV_X1 U944 ( .A(n1252), .ZN(n1086) );
XOR2_X1 U945 ( .A(G110), .B(n1204), .Z(G12) );
AND2_X1 U946 ( .A1(n1208), .A2(n1233), .ZN(n1204) );
NOR3_X1 U947 ( .A1(n1190), .A2(n1049), .A3(n1050), .ZN(n1233) );
XNOR2_X1 U948 ( .A(n1253), .B(G472), .ZN(n1050) );
NAND2_X1 U949 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
XOR2_X1 U950 ( .A(n1256), .B(n1141), .Z(n1254) );
XOR2_X1 U951 ( .A(n1257), .B(n1258), .Z(n1141) );
XNOR2_X1 U952 ( .A(G113), .B(n1259), .ZN(n1258) );
XOR2_X1 U953 ( .A(n1155), .B(n1260), .Z(n1257) );
NOR2_X1 U954 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
NOR3_X1 U955 ( .A1(KEYINPUT34), .A2(G119), .A3(n1263), .ZN(n1262) );
NOR2_X1 U956 ( .A1(n1264), .A2(n1265), .ZN(n1261) );
INV_X1 U957 ( .A(KEYINPUT34), .ZN(n1265) );
XNOR2_X1 U958 ( .A(n1244), .B(G116), .ZN(n1264) );
XNOR2_X1 U959 ( .A(n1266), .B(n1267), .ZN(n1155) );
NAND3_X1 U960 ( .A1(n1268), .A2(n1269), .A3(n1144), .ZN(n1256) );
NAND2_X1 U961 ( .A1(n1146), .A2(G101), .ZN(n1144) );
OR3_X1 U962 ( .A1(n1146), .A2(G101), .A3(KEYINPUT22), .ZN(n1269) );
NAND2_X1 U963 ( .A1(KEYINPUT22), .A2(n1146), .ZN(n1268) );
AND2_X1 U964 ( .A1(G210), .A2(n1270), .ZN(n1146) );
INV_X1 U965 ( .A(n1225), .ZN(n1049) );
XNOR2_X1 U966 ( .A(n1271), .B(n1124), .ZN(n1225) );
AND2_X1 U967 ( .A1(G217), .A2(n1272), .ZN(n1124) );
NAND2_X1 U968 ( .A1(n1122), .A2(n1255), .ZN(n1271) );
XNOR2_X1 U969 ( .A(n1273), .B(n1274), .ZN(n1122) );
XNOR2_X1 U970 ( .A(n1275), .B(n1276), .ZN(n1274) );
NAND2_X1 U971 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND2_X1 U972 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
INV_X1 U973 ( .A(KEYINPUT49), .ZN(n1280) );
NAND2_X1 U974 ( .A1(n1281), .A2(n1282), .ZN(n1279) );
NAND2_X1 U975 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NAND2_X1 U976 ( .A1(n1285), .A2(n1286), .ZN(n1281) );
NAND2_X1 U977 ( .A1(KEYINPUT49), .A2(n1287), .ZN(n1277) );
NAND2_X1 U978 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U979 ( .A1(n1286), .A2(n1284), .ZN(n1289) );
NAND2_X1 U980 ( .A1(n1101), .A2(n1290), .ZN(n1284) );
NAND2_X1 U981 ( .A1(G125), .A2(G140), .ZN(n1290) );
INV_X1 U982 ( .A(n1291), .ZN(n1101) );
INV_X1 U983 ( .A(n1283), .ZN(n1286) );
NAND2_X1 U984 ( .A1(n1285), .A2(n1283), .ZN(n1288) );
XNOR2_X1 U985 ( .A(n1292), .B(n1293), .ZN(n1283) );
NOR2_X1 U986 ( .A1(KEYINPUT57), .A2(G137), .ZN(n1293) );
NAND2_X1 U987 ( .A1(n1294), .A2(G221), .ZN(n1292) );
XNOR2_X1 U988 ( .A(n1107), .B(G125), .ZN(n1285) );
XNOR2_X1 U989 ( .A(G128), .B(n1295), .ZN(n1273) );
INV_X1 U990 ( .A(n1058), .ZN(n1190) );
NAND2_X1 U991 ( .A1(n1296), .A2(n1297), .ZN(n1058) );
OR2_X1 U992 ( .A1(n1041), .A2(KEYINPUT39), .ZN(n1297) );
INV_X1 U993 ( .A(n1223), .ZN(n1041) );
NOR2_X1 U994 ( .A1(n1059), .A2(n1072), .ZN(n1223) );
INV_X1 U995 ( .A(n1060), .ZN(n1072) );
NAND3_X1 U996 ( .A1(n1059), .A2(n1060), .A3(KEYINPUT39), .ZN(n1296) );
NAND2_X1 U997 ( .A1(G214), .A2(n1298), .ZN(n1060) );
XNOR2_X1 U998 ( .A(n1082), .B(n1083), .ZN(n1059) );
INV_X1 U999 ( .A(n1167), .ZN(n1083) );
NAND2_X1 U1000 ( .A1(G210), .A2(n1298), .ZN(n1167) );
NAND2_X1 U1001 ( .A1(n1299), .A2(n1255), .ZN(n1298) );
INV_X1 U1002 ( .A(G237), .ZN(n1299) );
NAND3_X1 U1003 ( .A1(n1300), .A2(n1255), .A3(n1301), .ZN(n1082) );
NAND2_X1 U1004 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NAND2_X1 U1005 ( .A1(n1118), .A2(n1304), .ZN(n1303) );
NAND2_X1 U1006 ( .A1(KEYINPUT54), .A2(KEYINPUT28), .ZN(n1304) );
XNOR2_X1 U1007 ( .A(n1305), .B(n1178), .ZN(n1302) );
NAND3_X1 U1008 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1300) );
XNOR2_X1 U1009 ( .A(n1118), .B(KEYINPUT28), .ZN(n1308) );
XNOR2_X1 U1010 ( .A(n1309), .B(n1310), .ZN(n1118) );
XNOR2_X1 U1011 ( .A(n1263), .B(n1311), .ZN(n1310) );
XNOR2_X1 U1012 ( .A(KEYINPUT63), .B(n1312), .ZN(n1311) );
INV_X1 U1013 ( .A(G116), .ZN(n1263) );
XNOR2_X1 U1014 ( .A(n1313), .B(n1314), .ZN(n1309) );
XNOR2_X1 U1015 ( .A(n1315), .B(n1275), .ZN(n1314) );
XNOR2_X1 U1016 ( .A(G110), .B(n1244), .ZN(n1275) );
INV_X1 U1017 ( .A(G119), .ZN(n1244) );
INV_X1 U1018 ( .A(n1316), .ZN(n1315) );
INV_X1 U1019 ( .A(KEYINPUT54), .ZN(n1307) );
XNOR2_X1 U1020 ( .A(n1176), .B(n1305), .ZN(n1306) );
NAND2_X1 U1021 ( .A1(KEYINPUT48), .A2(n1177), .ZN(n1305) );
XOR2_X1 U1022 ( .A(n1267), .B(n1317), .Z(n1177) );
XNOR2_X1 U1023 ( .A(G125), .B(n1259), .ZN(n1317) );
XNOR2_X1 U1024 ( .A(KEYINPUT59), .B(n1318), .ZN(n1259) );
NOR2_X1 U1025 ( .A1(KEYINPUT17), .A2(n1156), .ZN(n1318) );
INV_X1 U1026 ( .A(n1178), .ZN(n1176) );
NAND2_X1 U1027 ( .A1(G224), .A2(n1065), .ZN(n1178) );
NOR3_X1 U1028 ( .A1(n1055), .A2(n1209), .A3(n1037), .ZN(n1208) );
INV_X1 U1029 ( .A(n1232), .ZN(n1037) );
NOR2_X1 U1030 ( .A1(n1252), .A2(n1087), .ZN(n1232) );
XNOR2_X1 U1031 ( .A(n1319), .B(G478), .ZN(n1087) );
NAND2_X1 U1032 ( .A1(n1127), .A2(n1255), .ZN(n1319) );
XOR2_X1 U1033 ( .A(n1320), .B(n1321), .Z(n1127) );
XOR2_X1 U1034 ( .A(n1322), .B(n1323), .Z(n1321) );
NAND2_X1 U1035 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
NAND2_X1 U1036 ( .A1(G128), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1037 ( .A(n1327), .B(KEYINPUT26), .Z(n1324) );
OR2_X1 U1038 ( .A1(n1326), .A2(G128), .ZN(n1327) );
NAND2_X1 U1039 ( .A1(n1294), .A2(G217), .ZN(n1322) );
AND2_X1 U1040 ( .A1(G234), .A2(n1065), .ZN(n1294) );
XOR2_X1 U1041 ( .A(n1328), .B(G134), .Z(n1320) );
NAND3_X1 U1042 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1328) );
OR2_X1 U1043 ( .A1(n1332), .A2(G107), .ZN(n1331) );
NAND2_X1 U1044 ( .A1(n1333), .A2(n1334), .ZN(n1330) );
INV_X1 U1045 ( .A(KEYINPUT13), .ZN(n1334) );
NAND2_X1 U1046 ( .A1(G107), .A2(n1335), .ZN(n1333) );
XNOR2_X1 U1047 ( .A(KEYINPUT36), .B(n1332), .ZN(n1335) );
NAND2_X1 U1048 ( .A1(KEYINPUT13), .A2(n1336), .ZN(n1329) );
NAND2_X1 U1049 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
NAND3_X1 U1050 ( .A1(KEYINPUT36), .A2(G107), .A3(n1332), .ZN(n1338) );
OR2_X1 U1051 ( .A1(n1332), .A2(KEYINPUT36), .ZN(n1337) );
NAND2_X1 U1052 ( .A1(n1339), .A2(n1340), .ZN(n1332) );
NAND2_X1 U1053 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
XNOR2_X1 U1054 ( .A(n1343), .B(KEYINPUT44), .ZN(n1342) );
XNOR2_X1 U1055 ( .A(G122), .B(KEYINPUT19), .ZN(n1341) );
XOR2_X1 U1056 ( .A(KEYINPUT0), .B(n1344), .Z(n1339) );
NOR2_X1 U1057 ( .A1(n1312), .A2(n1343), .ZN(n1344) );
XOR2_X1 U1058 ( .A(G116), .B(KEYINPUT61), .Z(n1343) );
XNOR2_X1 U1059 ( .A(n1345), .B(G475), .ZN(n1252) );
NAND2_X1 U1060 ( .A1(n1130), .A2(n1255), .ZN(n1345) );
XNOR2_X1 U1061 ( .A(n1346), .B(n1347), .ZN(n1130) );
XOR2_X1 U1062 ( .A(n1348), .B(n1349), .Z(n1347) );
XNOR2_X1 U1063 ( .A(n1350), .B(n1351), .ZN(n1349) );
NOR2_X1 U1064 ( .A1(KEYINPUT3), .A2(n1352), .ZN(n1351) );
XOR2_X1 U1065 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1066 ( .A(n1355), .B(G131), .Z(n1354) );
NAND2_X1 U1067 ( .A1(G214), .A2(n1270), .ZN(n1355) );
NOR2_X1 U1068 ( .A1(G953), .A2(G237), .ZN(n1270) );
XNOR2_X1 U1069 ( .A(G143), .B(KEYINPUT6), .ZN(n1353) );
NAND2_X1 U1070 ( .A1(KEYINPUT23), .A2(n1312), .ZN(n1350) );
INV_X1 U1071 ( .A(G122), .ZN(n1312) );
NOR3_X1 U1072 ( .A1(n1291), .A2(n1356), .A3(n1357), .ZN(n1348) );
AND3_X1 U1073 ( .A1(KEYINPUT5), .A2(G140), .A3(G125), .ZN(n1357) );
NOR2_X1 U1074 ( .A1(KEYINPUT5), .A2(G125), .ZN(n1356) );
NOR2_X1 U1075 ( .A1(G125), .A2(G140), .ZN(n1291) );
XNOR2_X1 U1076 ( .A(n1316), .B(n1295), .ZN(n1346) );
XNOR2_X1 U1077 ( .A(n1156), .B(KEYINPUT56), .ZN(n1295) );
INV_X1 U1078 ( .A(G146), .ZN(n1156) );
XOR2_X1 U1079 ( .A(G104), .B(G113), .Z(n1316) );
AND2_X1 U1080 ( .A1(n1033), .A2(n1358), .ZN(n1209) );
NAND3_X1 U1081 ( .A1(n1113), .A2(n1236), .A3(G902), .ZN(n1358) );
NOR2_X1 U1082 ( .A1(G898), .A2(n1065), .ZN(n1113) );
NAND3_X1 U1083 ( .A1(n1236), .A2(n1065), .A3(G952), .ZN(n1033) );
NAND2_X1 U1084 ( .A1(G237), .A2(G234), .ZN(n1236) );
NAND2_X1 U1085 ( .A1(n1052), .A2(n1051), .ZN(n1055) );
NAND2_X1 U1086 ( .A1(G221), .A2(n1272), .ZN(n1051) );
NAND2_X1 U1087 ( .A1(G234), .A2(n1255), .ZN(n1272) );
XOR2_X1 U1088 ( .A(n1359), .B(G469), .Z(n1052) );
NAND2_X1 U1089 ( .A1(KEYINPUT9), .A2(n1079), .ZN(n1359) );
NAND2_X1 U1090 ( .A1(n1360), .A2(n1255), .ZN(n1079) );
INV_X1 U1091 ( .A(G902), .ZN(n1255) );
XOR2_X1 U1092 ( .A(n1361), .B(n1362), .Z(n1360) );
XNOR2_X1 U1093 ( .A(n1154), .B(n1363), .ZN(n1362) );
INV_X1 U1094 ( .A(n1266), .ZN(n1363) );
XOR2_X1 U1095 ( .A(G131), .B(n1364), .Z(n1266) );
XNOR2_X1 U1096 ( .A(n1221), .B(G134), .ZN(n1364) );
INV_X1 U1097 ( .A(G137), .ZN(n1221) );
XNOR2_X1 U1098 ( .A(G104), .B(n1313), .ZN(n1154) );
XOR2_X1 U1099 ( .A(G101), .B(G107), .Z(n1313) );
XOR2_X1 U1100 ( .A(n1365), .B(n1366), .Z(n1361) );
NOR2_X1 U1101 ( .A1(KEYINPUT2), .A2(n1367), .ZN(n1366) );
XNOR2_X1 U1102 ( .A(G146), .B(n1267), .ZN(n1367) );
XNOR2_X1 U1103 ( .A(G128), .B(n1326), .ZN(n1267) );
INV_X1 U1104 ( .A(G143), .ZN(n1326) );
NAND2_X1 U1105 ( .A1(n1368), .A2(n1369), .ZN(n1365) );
XOR2_X1 U1106 ( .A(KEYINPUT62), .B(KEYINPUT41), .Z(n1369) );
XOR2_X1 U1107 ( .A(n1370), .B(n1158), .Z(n1368) );
XNOR2_X1 U1108 ( .A(G110), .B(n1107), .ZN(n1158) );
INV_X1 U1109 ( .A(G140), .ZN(n1107) );
NAND2_X1 U1110 ( .A1(KEYINPUT1), .A2(n1151), .ZN(n1370) );
NAND2_X1 U1111 ( .A1(G227), .A2(n1065), .ZN(n1151) );
INV_X1 U1112 ( .A(G953), .ZN(n1065) );
endmodule


