//Key = 0110010111110011000011100000110110100111011101111111000101110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342;

XNOR2_X1 U734 ( .A(G107), .B(n1018), .ZN(G9) );
NOR2_X1 U735 ( .A1(n1019), .A2(n1020), .ZN(G75) );
NOR4_X1 U736 ( .A1(n1021), .A2(n1022), .A3(G953), .A4(n1023), .ZN(n1020) );
NOR2_X1 U737 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U738 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U739 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR2_X1 U740 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR2_X1 U741 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U742 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U743 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR2_X1 U744 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U745 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U746 ( .A1(n1042), .A2(n1043), .ZN(n1034) );
NOR2_X1 U747 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
AND4_X1 U748 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1030) );
NOR3_X1 U749 ( .A1(n1037), .A2(n1050), .A3(n1043), .ZN(n1026) );
INV_X1 U750 ( .A(n1048), .ZN(n1043) );
NOR2_X1 U751 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U752 ( .A1(n1053), .A2(n1033), .ZN(n1052) );
NOR3_X1 U753 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NOR2_X1 U754 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
INV_X1 U755 ( .A(KEYINPUT35), .ZN(n1058) );
NOR2_X1 U756 ( .A1(n1059), .A2(n1060), .ZN(n1054) );
NOR4_X1 U757 ( .A1(KEYINPUT35), .A2(n1047), .A3(n1057), .A4(n1046), .ZN(n1051) );
XNOR2_X1 U758 ( .A(n1061), .B(KEYINPUT52), .ZN(n1057) );
NAND3_X1 U759 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1021) );
XNOR2_X1 U760 ( .A(n1065), .B(KEYINPUT41), .ZN(n1064) );
NOR3_X1 U761 ( .A1(n1023), .A2(G953), .A3(G952), .ZN(n1019) );
AND4_X1 U762 ( .A1(n1061), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1023) );
NOR4_X1 U763 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1068) );
INV_X1 U764 ( .A(n1073), .ZN(n1070) );
XNOR2_X1 U765 ( .A(n1074), .B(n1075), .ZN(n1067) );
NAND2_X1 U766 ( .A1(KEYINPUT45), .A2(n1076), .ZN(n1074) );
NAND2_X1 U767 ( .A1(n1077), .A2(n1078), .ZN(G72) );
NAND2_X1 U768 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U769 ( .A1(G953), .A2(n1081), .ZN(n1080) );
NAND3_X1 U770 ( .A1(G953), .A2(n1082), .A3(n1083), .ZN(n1077) );
INV_X1 U771 ( .A(n1079), .ZN(n1083) );
NOR2_X1 U772 ( .A1(KEYINPUT56), .A2(n1084), .ZN(n1079) );
XOR2_X1 U773 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U774 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U775 ( .A(n1089), .B(n1090), .Z(n1088) );
XNOR2_X1 U776 ( .A(n1091), .B(n1092), .ZN(n1090) );
XOR2_X1 U777 ( .A(n1093), .B(n1094), .Z(n1091) );
NAND2_X1 U778 ( .A1(KEYINPUT11), .A2(G125), .ZN(n1093) );
XOR2_X1 U779 ( .A(n1095), .B(n1096), .Z(n1089) );
XNOR2_X1 U780 ( .A(KEYINPUT7), .B(n1097), .ZN(n1096) );
NAND2_X1 U781 ( .A1(KEYINPUT1), .A2(G131), .ZN(n1095) );
NOR2_X1 U782 ( .A1(G900), .A2(n1098), .ZN(n1087) );
NAND2_X1 U783 ( .A1(n1098), .A2(n1099), .ZN(n1085) );
NAND3_X1 U784 ( .A1(n1063), .A2(n1100), .A3(n1101), .ZN(n1099) );
XOR2_X1 U785 ( .A(n1102), .B(KEYINPUT39), .Z(n1101) );
NAND2_X1 U786 ( .A1(G900), .A2(G227), .ZN(n1082) );
XOR2_X1 U787 ( .A(n1103), .B(n1104), .Z(G69) );
XOR2_X1 U788 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U789 ( .A1(n1107), .A2(n1098), .ZN(n1106) );
AND2_X1 U790 ( .A1(G224), .A2(G898), .ZN(n1107) );
NAND2_X1 U791 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
NAND2_X1 U792 ( .A1(G953), .A2(n1110), .ZN(n1109) );
XNOR2_X1 U793 ( .A(n1111), .B(n1112), .ZN(n1108) );
NAND2_X1 U794 ( .A1(n1098), .A2(n1113), .ZN(n1103) );
NOR2_X1 U795 ( .A1(n1114), .A2(n1115), .ZN(G66) );
XOR2_X1 U796 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U797 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U798 ( .A1(n1114), .A2(n1120), .ZN(G63) );
NOR2_X1 U799 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U800 ( .A(KEYINPUT3), .B(n1123), .Z(n1122) );
AND2_X1 U801 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NOR2_X1 U802 ( .A1(n1125), .A2(n1124), .ZN(n1121) );
NOR2_X1 U803 ( .A1(n1119), .A2(n1126), .ZN(n1125) );
INV_X1 U804 ( .A(G478), .ZN(n1126) );
NOR2_X1 U805 ( .A1(n1114), .A2(n1127), .ZN(G60) );
XOR2_X1 U806 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U807 ( .A1(n1130), .A2(n1119), .ZN(n1128) );
XOR2_X1 U808 ( .A(G104), .B(n1131), .Z(G6) );
NOR2_X1 U809 ( .A1(n1132), .A2(n1133), .ZN(G57) );
XOR2_X1 U810 ( .A(KEYINPUT24), .B(n1114), .Z(n1133) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(n1132) );
XNOR2_X1 U812 ( .A(n1136), .B(n1137), .ZN(n1135) );
NAND2_X1 U813 ( .A1(KEYINPUT38), .A2(n1138), .ZN(n1136) );
XOR2_X1 U814 ( .A(n1139), .B(n1140), .Z(n1134) );
NOR2_X1 U815 ( .A1(n1075), .A2(n1119), .ZN(n1140) );
NAND2_X1 U816 ( .A1(KEYINPUT50), .A2(n1141), .ZN(n1139) );
NOR2_X1 U817 ( .A1(n1114), .A2(n1142), .ZN(G54) );
XOR2_X1 U818 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U819 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR2_X1 U820 ( .A1(n1147), .A2(n1119), .ZN(n1146) );
NOR2_X1 U821 ( .A1(KEYINPUT40), .A2(n1148), .ZN(n1145) );
XOR2_X1 U822 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U823 ( .A1(KEYINPUT23), .A2(n1151), .ZN(n1150) );
NAND3_X1 U824 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1149) );
NAND2_X1 U825 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
OR3_X1 U826 ( .A1(n1156), .A2(n1155), .A3(n1157), .ZN(n1153) );
XOR2_X1 U827 ( .A(n1158), .B(KEYINPUT49), .Z(n1155) );
OR2_X1 U828 ( .A1(KEYINPUT36), .A2(n1159), .ZN(n1156) );
NAND2_X1 U829 ( .A1(n1159), .A2(n1157), .ZN(n1152) );
INV_X1 U830 ( .A(KEYINPUT58), .ZN(n1157) );
NAND3_X1 U831 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1143) );
NAND2_X1 U832 ( .A1(n1163), .A2(KEYINPUT47), .ZN(n1161) );
NAND2_X1 U833 ( .A1(n1164), .A2(n1165), .ZN(n1160) );
INV_X1 U834 ( .A(KEYINPUT47), .ZN(n1165) );
NOR2_X1 U835 ( .A1(n1114), .A2(n1166), .ZN(G51) );
XNOR2_X1 U836 ( .A(n1167), .B(n1168), .ZN(n1166) );
XOR2_X1 U837 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U838 ( .A1(n1171), .A2(n1119), .ZN(n1170) );
NAND2_X1 U839 ( .A1(G902), .A2(n1172), .ZN(n1119) );
NAND3_X1 U840 ( .A1(n1063), .A2(n1065), .A3(n1062), .ZN(n1172) );
AND2_X1 U841 ( .A1(n1173), .A2(n1100), .ZN(n1062) );
NAND2_X1 U842 ( .A1(n1174), .A2(n1061), .ZN(n1100) );
XNOR2_X1 U843 ( .A(KEYINPUT63), .B(n1102), .ZN(n1173) );
NAND4_X1 U844 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1102) );
NAND3_X1 U845 ( .A1(n1179), .A2(n1044), .A3(n1039), .ZN(n1175) );
INV_X1 U846 ( .A(n1113), .ZN(n1065) );
NAND4_X1 U847 ( .A1(n1180), .A2(n1018), .A3(n1181), .A4(n1182), .ZN(n1113) );
NOR4_X1 U848 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1131), .ZN(n1182) );
AND3_X1 U849 ( .A1(n1186), .A2(n1045), .A3(n1048), .ZN(n1131) );
NAND2_X1 U850 ( .A1(n1187), .A2(n1188), .ZN(n1181) );
NAND2_X1 U851 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U852 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XNOR2_X1 U853 ( .A(KEYINPUT16), .B(n1037), .ZN(n1192) );
NAND2_X1 U854 ( .A1(n1039), .A2(n1044), .ZN(n1189) );
NAND3_X1 U855 ( .A1(n1048), .A2(n1186), .A3(n1044), .ZN(n1018) );
AND3_X1 U856 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1063) );
NOR2_X1 U857 ( .A1(n1196), .A2(n1197), .ZN(n1169) );
XNOR2_X1 U858 ( .A(n1198), .B(KEYINPUT10), .ZN(n1197) );
NOR2_X1 U859 ( .A1(n1199), .A2(n1200), .ZN(n1196) );
NOR2_X1 U860 ( .A1(n1201), .A2(G952), .ZN(n1114) );
XNOR2_X1 U861 ( .A(n1098), .B(KEYINPUT22), .ZN(n1201) );
NAND2_X1 U862 ( .A1(n1202), .A2(n1203), .ZN(G48) );
OR2_X1 U863 ( .A1(n1195), .A2(G146), .ZN(n1203) );
XOR2_X1 U864 ( .A(n1204), .B(KEYINPUT30), .Z(n1202) );
NAND2_X1 U865 ( .A1(G146), .A2(n1195), .ZN(n1204) );
NAND3_X1 U866 ( .A1(n1191), .A2(n1045), .A3(n1205), .ZN(n1195) );
XNOR2_X1 U867 ( .A(G143), .B(n1193), .ZN(G45) );
NAND3_X1 U868 ( .A1(n1039), .A2(n1205), .A3(n1206), .ZN(n1193) );
XNOR2_X1 U869 ( .A(G140), .B(n1194), .ZN(G42) );
NAND2_X1 U870 ( .A1(n1179), .A2(n1207), .ZN(n1194) );
XOR2_X1 U871 ( .A(n1208), .B(n1209), .Z(G39) );
NAND2_X1 U872 ( .A1(KEYINPUT21), .A2(G137), .ZN(n1209) );
NAND2_X1 U873 ( .A1(n1061), .A2(n1210), .ZN(n1208) );
XOR2_X1 U874 ( .A(KEYINPUT18), .B(n1174), .Z(n1210) );
AND3_X1 U875 ( .A1(n1211), .A2(n1191), .A3(n1049), .ZN(n1174) );
XNOR2_X1 U876 ( .A(G134), .B(n1212), .ZN(G36) );
NAND3_X1 U877 ( .A1(n1179), .A2(n1044), .A3(n1213), .ZN(n1212) );
XNOR2_X1 U878 ( .A(n1039), .B(KEYINPUT29), .ZN(n1213) );
XNOR2_X1 U879 ( .A(G131), .B(n1176), .ZN(G33) );
NAND3_X1 U880 ( .A1(n1179), .A2(n1045), .A3(n1039), .ZN(n1176) );
AND2_X1 U881 ( .A1(n1211), .A2(n1061), .ZN(n1179) );
INV_X1 U882 ( .A(n1029), .ZN(n1061) );
NAND2_X1 U883 ( .A1(n1214), .A2(n1060), .ZN(n1029) );
INV_X1 U884 ( .A(n1059), .ZN(n1214) );
XOR2_X1 U885 ( .A(n1177), .B(n1215), .Z(G30) );
XOR2_X1 U886 ( .A(KEYINPUT32), .B(G128), .Z(n1215) );
NAND3_X1 U887 ( .A1(n1191), .A2(n1044), .A3(n1205), .ZN(n1177) );
AND2_X1 U888 ( .A1(n1211), .A2(n1055), .ZN(n1205) );
AND3_X1 U889 ( .A1(n1216), .A2(n1046), .A3(n1047), .ZN(n1211) );
XOR2_X1 U890 ( .A(G101), .B(n1185), .Z(G3) );
AND3_X1 U891 ( .A1(n1049), .A2(n1186), .A3(n1039), .ZN(n1185) );
XNOR2_X1 U892 ( .A(G125), .B(n1178), .ZN(G27) );
NAND4_X1 U893 ( .A1(n1207), .A2(n1066), .A3(n1055), .A4(n1216), .ZN(n1178) );
NAND2_X1 U894 ( .A1(n1025), .A2(n1217), .ZN(n1216) );
NAND4_X1 U895 ( .A1(G953), .A2(G902), .A3(n1218), .A4(n1219), .ZN(n1217) );
INV_X1 U896 ( .A(G900), .ZN(n1219) );
AND3_X1 U897 ( .A1(n1045), .A2(n1071), .A3(n1220), .ZN(n1207) );
XNOR2_X1 U898 ( .A(G122), .B(n1221), .ZN(G24) );
NOR2_X1 U899 ( .A1(n1222), .A2(KEYINPUT6), .ZN(n1221) );
INV_X1 U900 ( .A(n1180), .ZN(n1222) );
NAND3_X1 U901 ( .A1(n1206), .A2(n1048), .A3(n1187), .ZN(n1180) );
NOR2_X1 U902 ( .A1(n1071), .A2(n1041), .ZN(n1048) );
INV_X1 U903 ( .A(n1220), .ZN(n1041) );
AND2_X1 U904 ( .A1(n1223), .A2(n1072), .ZN(n1206) );
XNOR2_X1 U905 ( .A(n1224), .B(KEYINPUT26), .ZN(n1223) );
XNOR2_X1 U906 ( .A(n1225), .B(n1226), .ZN(G21) );
AND3_X1 U907 ( .A1(n1187), .A2(n1191), .A3(n1049), .ZN(n1226) );
NOR2_X1 U908 ( .A1(n1220), .A2(n1040), .ZN(n1191) );
INV_X1 U909 ( .A(n1071), .ZN(n1040) );
XNOR2_X1 U910 ( .A(G116), .B(n1227), .ZN(G18) );
NAND4_X1 U911 ( .A1(n1228), .A2(n1229), .A3(n1044), .A4(n1230), .ZN(n1227) );
AND2_X1 U912 ( .A1(n1066), .A2(n1039), .ZN(n1230) );
NOR2_X1 U913 ( .A1(n1072), .A2(n1224), .ZN(n1044) );
XOR2_X1 U914 ( .A(KEYINPUT19), .B(n1055), .Z(n1228) );
XOR2_X1 U915 ( .A(G113), .B(n1184), .Z(G15) );
AND3_X1 U916 ( .A1(n1039), .A2(n1045), .A3(n1187), .ZN(n1184) );
AND3_X1 U917 ( .A1(n1055), .A2(n1229), .A3(n1066), .ZN(n1187) );
INV_X1 U918 ( .A(n1033), .ZN(n1066) );
NAND2_X1 U919 ( .A1(n1231), .A2(n1046), .ZN(n1033) );
INV_X1 U920 ( .A(n1047), .ZN(n1231) );
NAND2_X1 U921 ( .A1(n1232), .A2(n1233), .ZN(n1045) );
OR2_X1 U922 ( .A1(n1037), .A2(KEYINPUT51), .ZN(n1233) );
INV_X1 U923 ( .A(n1049), .ZN(n1037) );
NAND3_X1 U924 ( .A1(n1224), .A2(n1072), .A3(KEYINPUT51), .ZN(n1232) );
INV_X1 U925 ( .A(n1234), .ZN(n1224) );
NOR2_X1 U926 ( .A1(n1071), .A2(n1220), .ZN(n1039) );
XOR2_X1 U927 ( .A(G110), .B(n1183), .Z(G12) );
AND4_X1 U928 ( .A1(n1049), .A2(n1186), .A3(n1220), .A4(n1071), .ZN(n1183) );
NAND3_X1 U929 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1071) );
NAND2_X1 U930 ( .A1(n1238), .A2(n1116), .ZN(n1237) );
OR3_X1 U931 ( .A1(n1116), .A2(n1238), .A3(G902), .ZN(n1236) );
NOR2_X1 U932 ( .A1(n1118), .A2(G234), .ZN(n1238) );
INV_X1 U933 ( .A(G217), .ZN(n1118) );
XOR2_X1 U934 ( .A(n1239), .B(n1240), .Z(n1116) );
XNOR2_X1 U935 ( .A(n1241), .B(n1242), .ZN(n1240) );
NAND2_X1 U936 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
OR2_X1 U937 ( .A1(n1245), .A2(KEYINPUT17), .ZN(n1244) );
NAND3_X1 U938 ( .A1(G140), .A2(n1246), .A3(KEYINPUT17), .ZN(n1243) );
XOR2_X1 U939 ( .A(n1247), .B(n1248), .Z(n1239) );
XNOR2_X1 U940 ( .A(n1225), .B(G110), .ZN(n1248) );
NAND2_X1 U941 ( .A1(n1249), .A2(n1250), .ZN(n1247) );
NAND4_X1 U942 ( .A1(n1251), .A2(G221), .A3(G234), .A4(n1098), .ZN(n1250) );
XOR2_X1 U943 ( .A(n1252), .B(KEYINPUT0), .Z(n1249) );
NAND2_X1 U944 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NAND3_X1 U945 ( .A1(G234), .A2(n1098), .A3(G221), .ZN(n1254) );
NAND2_X1 U946 ( .A1(G902), .A2(G217), .ZN(n1235) );
XOR2_X1 U947 ( .A(n1076), .B(n1075), .Z(n1220) );
INV_X1 U948 ( .A(G472), .ZN(n1075) );
AND3_X1 U949 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1076) );
NAND2_X1 U950 ( .A1(n1258), .A2(n1141), .ZN(n1257) );
XNOR2_X1 U951 ( .A(n1259), .B(n1260), .ZN(n1258) );
INV_X1 U952 ( .A(n1137), .ZN(n1260) );
NAND2_X1 U953 ( .A1(n1261), .A2(n1262), .ZN(n1255) );
XOR2_X1 U954 ( .A(n1141), .B(n1263), .Z(n1262) );
XNOR2_X1 U955 ( .A(KEYINPUT5), .B(KEYINPUT37), .ZN(n1263) );
XNOR2_X1 U956 ( .A(G101), .B(n1264), .ZN(n1141) );
AND3_X1 U957 ( .A1(G210), .A2(n1098), .A3(n1265), .ZN(n1264) );
XNOR2_X1 U958 ( .A(n1259), .B(n1137), .ZN(n1261) );
XNOR2_X1 U959 ( .A(n1266), .B(n1267), .ZN(n1137) );
XNOR2_X1 U960 ( .A(KEYINPUT9), .B(n1225), .ZN(n1267) );
XNOR2_X1 U961 ( .A(G113), .B(G116), .ZN(n1266) );
NAND2_X1 U962 ( .A1(KEYINPUT15), .A2(n1268), .ZN(n1259) );
XOR2_X1 U963 ( .A(KEYINPUT57), .B(n1138), .Z(n1268) );
XOR2_X1 U964 ( .A(n1151), .B(n1269), .Z(n1138) );
AND4_X1 U965 ( .A1(n1047), .A2(n1055), .A3(n1229), .A4(n1046), .ZN(n1186) );
NAND2_X1 U966 ( .A1(n1270), .A2(G221), .ZN(n1046) );
XOR2_X1 U967 ( .A(n1271), .B(KEYINPUT54), .Z(n1270) );
NAND2_X1 U968 ( .A1(G234), .A2(n1256), .ZN(n1271) );
NAND2_X1 U969 ( .A1(n1025), .A2(n1272), .ZN(n1229) );
NAND4_X1 U970 ( .A1(G953), .A2(G902), .A3(n1273), .A4(n1110), .ZN(n1272) );
INV_X1 U971 ( .A(G898), .ZN(n1110) );
XNOR2_X1 U972 ( .A(KEYINPUT48), .B(n1218), .ZN(n1273) );
NAND3_X1 U973 ( .A1(n1218), .A2(n1098), .A3(G952), .ZN(n1025) );
NAND2_X1 U974 ( .A1(G237), .A2(G234), .ZN(n1218) );
AND2_X1 U975 ( .A1(n1059), .A2(n1060), .ZN(n1055) );
NAND2_X1 U976 ( .A1(G214), .A2(n1274), .ZN(n1060) );
XOR2_X1 U977 ( .A(n1275), .B(n1171), .Z(n1059) );
NAND2_X1 U978 ( .A1(G210), .A2(n1274), .ZN(n1171) );
NAND2_X1 U979 ( .A1(n1265), .A2(n1256), .ZN(n1274) );
NAND2_X1 U980 ( .A1(n1276), .A2(n1256), .ZN(n1275) );
XNOR2_X1 U981 ( .A(n1277), .B(n1278), .ZN(n1276) );
INV_X1 U982 ( .A(n1167), .ZN(n1278) );
XNOR2_X1 U983 ( .A(n1111), .B(n1279), .ZN(n1167) );
XNOR2_X1 U984 ( .A(n1280), .B(KEYINPUT60), .ZN(n1279) );
NAND2_X1 U985 ( .A1(KEYINPUT46), .A2(n1112), .ZN(n1280) );
XNOR2_X1 U986 ( .A(G110), .B(n1281), .ZN(n1112) );
XNOR2_X1 U987 ( .A(KEYINPUT2), .B(n1282), .ZN(n1281) );
XOR2_X1 U988 ( .A(n1283), .B(n1284), .Z(n1111) );
XOR2_X1 U989 ( .A(n1285), .B(n1286), .Z(n1284) );
NOR2_X1 U990 ( .A1(KEYINPUT27), .A2(n1225), .ZN(n1286) );
INV_X1 U991 ( .A(G119), .ZN(n1225) );
NOR2_X1 U992 ( .A1(G113), .A2(KEYINPUT53), .ZN(n1285) );
XNOR2_X1 U993 ( .A(n1287), .B(n1288), .ZN(n1283) );
NAND2_X1 U994 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
NAND3_X1 U995 ( .A1(n1291), .A2(n1292), .A3(G101), .ZN(n1290) );
XOR2_X1 U996 ( .A(KEYINPUT14), .B(n1293), .Z(n1289) );
NOR2_X1 U997 ( .A1(G101), .A2(n1294), .ZN(n1293) );
AND2_X1 U998 ( .A1(n1291), .A2(n1292), .ZN(n1294) );
NAND3_X1 U999 ( .A1(n1295), .A2(n1296), .A3(G104), .ZN(n1292) );
OR2_X1 U1000 ( .A1(n1296), .A2(n1297), .ZN(n1291) );
INV_X1 U1001 ( .A(KEYINPUT31), .ZN(n1296) );
NOR2_X1 U1002 ( .A1(n1198), .A2(n1298), .ZN(n1277) );
NOR2_X1 U1003 ( .A1(n1200), .A2(n1299), .ZN(n1298) );
XNOR2_X1 U1004 ( .A(KEYINPUT55), .B(n1199), .ZN(n1299) );
AND2_X1 U1005 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND2_X1 U1006 ( .A1(G224), .A2(n1098), .ZN(n1200) );
XOR2_X1 U1007 ( .A(n1246), .B(n1269), .Z(n1199) );
XNOR2_X1 U1008 ( .A(n1092), .B(KEYINPUT62), .ZN(n1269) );
INV_X1 U1009 ( .A(G125), .ZN(n1246) );
XOR2_X1 U1010 ( .A(n1300), .B(n1301), .Z(n1047) );
XNOR2_X1 U1011 ( .A(KEYINPUT61), .B(n1147), .ZN(n1301) );
INV_X1 U1012 ( .A(G469), .ZN(n1147) );
NAND2_X1 U1013 ( .A1(n1302), .A2(n1256), .ZN(n1300) );
INV_X1 U1014 ( .A(G902), .ZN(n1256) );
XOR2_X1 U1015 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U1016 ( .A(n1092), .B(n1159), .ZN(n1304) );
XOR2_X1 U1017 ( .A(G101), .B(n1297), .Z(n1159) );
XNOR2_X1 U1018 ( .A(G104), .B(n1295), .ZN(n1297) );
INV_X1 U1019 ( .A(G107), .ZN(n1295) );
INV_X1 U1020 ( .A(n1158), .ZN(n1092) );
XOR2_X1 U1021 ( .A(G143), .B(n1241), .Z(n1158) );
XOR2_X1 U1022 ( .A(G128), .B(G146), .Z(n1241) );
XOR2_X1 U1023 ( .A(n1305), .B(n1306), .Z(n1303) );
NOR2_X1 U1024 ( .A1(KEYINPUT12), .A2(n1151), .ZN(n1306) );
XOR2_X1 U1025 ( .A(n1094), .B(G131), .Z(n1151) );
XNOR2_X1 U1026 ( .A(G134), .B(n1251), .ZN(n1094) );
INV_X1 U1027 ( .A(n1253), .ZN(n1251) );
XOR2_X1 U1028 ( .A(G137), .B(KEYINPUT43), .Z(n1253) );
NAND2_X1 U1029 ( .A1(n1307), .A2(n1162), .ZN(n1305) );
NAND2_X1 U1030 ( .A1(n1308), .A2(n1164), .ZN(n1162) );
INV_X1 U1031 ( .A(n1163), .ZN(n1307) );
NOR2_X1 U1032 ( .A1(n1164), .A2(n1308), .ZN(n1163) );
NOR2_X1 U1033 ( .A1(n1081), .A2(G953), .ZN(n1308) );
INV_X1 U1034 ( .A(G227), .ZN(n1081) );
XOR2_X1 U1035 ( .A(G110), .B(n1097), .Z(n1164) );
NOR2_X1 U1036 ( .A1(n1234), .A2(n1072), .ZN(n1049) );
XOR2_X1 U1037 ( .A(n1309), .B(n1130), .Z(n1072) );
INV_X1 U1038 ( .A(G475), .ZN(n1130) );
OR2_X1 U1039 ( .A1(n1129), .A2(G902), .ZN(n1309) );
XNOR2_X1 U1040 ( .A(n1310), .B(n1311), .ZN(n1129) );
XOR2_X1 U1041 ( .A(n1312), .B(n1245), .Z(n1311) );
XNOR2_X1 U1042 ( .A(G125), .B(n1097), .ZN(n1245) );
INV_X1 U1043 ( .A(G140), .ZN(n1097) );
NOR2_X1 U1044 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U1045 ( .A(KEYINPUT25), .B(n1315), .Z(n1314) );
NOR2_X1 U1046 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
AND2_X1 U1047 ( .A1(n1316), .A2(n1317), .ZN(n1313) );
NAND3_X1 U1048 ( .A1(n1265), .A2(n1098), .A3(n1318), .ZN(n1317) );
XNOR2_X1 U1049 ( .A(G214), .B(KEYINPUT34), .ZN(n1318) );
INV_X1 U1050 ( .A(G237), .ZN(n1265) );
XOR2_X1 U1051 ( .A(n1319), .B(n1320), .Z(n1310) );
XOR2_X1 U1052 ( .A(G146), .B(G131), .Z(n1320) );
NAND2_X1 U1053 ( .A1(n1321), .A2(KEYINPUT42), .ZN(n1319) );
XOR2_X1 U1054 ( .A(n1322), .B(G104), .Z(n1321) );
NAND2_X1 U1055 ( .A1(KEYINPUT28), .A2(n1323), .ZN(n1322) );
XOR2_X1 U1056 ( .A(G113), .B(n1324), .Z(n1323) );
XNOR2_X1 U1057 ( .A(KEYINPUT44), .B(n1282), .ZN(n1324) );
NAND2_X1 U1058 ( .A1(n1325), .A2(n1073), .ZN(n1234) );
NAND2_X1 U1059 ( .A1(G478), .A2(n1326), .ZN(n1073) );
OR2_X1 U1060 ( .A1(n1124), .A2(G902), .ZN(n1326) );
XNOR2_X1 U1061 ( .A(n1069), .B(KEYINPUT13), .ZN(n1325) );
NOR3_X1 U1062 ( .A1(G478), .A2(G902), .A3(n1124), .ZN(n1069) );
XNOR2_X1 U1063 ( .A(n1327), .B(n1328), .ZN(n1124) );
XNOR2_X1 U1064 ( .A(G107), .B(n1329), .ZN(n1328) );
NAND3_X1 U1065 ( .A1(G217), .A2(n1098), .A3(n1330), .ZN(n1329) );
XNOR2_X1 U1066 ( .A(G234), .B(KEYINPUT59), .ZN(n1330) );
INV_X1 U1067 ( .A(G953), .ZN(n1098) );
XOR2_X1 U1068 ( .A(n1331), .B(n1332), .Z(n1327) );
NOR3_X1 U1069 ( .A1(n1333), .A2(n1334), .A3(n1335), .ZN(n1332) );
NOR2_X1 U1070 ( .A1(n1336), .A2(n1288), .ZN(n1335) );
INV_X1 U1071 ( .A(G116), .ZN(n1288) );
AND3_X1 U1072 ( .A1(n1336), .A2(n1282), .A3(n1337), .ZN(n1334) );
INV_X1 U1073 ( .A(KEYINPUT33), .ZN(n1336) );
NOR2_X1 U1074 ( .A1(n1337), .A2(n1282), .ZN(n1333) );
INV_X1 U1075 ( .A(G122), .ZN(n1282) );
NOR2_X1 U1076 ( .A1(G116), .A2(KEYINPUT4), .ZN(n1337) );
NAND3_X1 U1077 ( .A1(n1338), .A2(n1339), .A3(KEYINPUT20), .ZN(n1331) );
OR3_X1 U1078 ( .A1(n1340), .A2(G134), .A3(KEYINPUT8), .ZN(n1339) );
NAND2_X1 U1079 ( .A1(n1341), .A2(KEYINPUT8), .ZN(n1338) );
XNOR2_X1 U1080 ( .A(n1342), .B(n1340), .ZN(n1341) );
XNOR2_X1 U1081 ( .A(G128), .B(n1316), .ZN(n1340) );
INV_X1 U1082 ( .A(G143), .ZN(n1316) );
INV_X1 U1083 ( .A(G134), .ZN(n1342) );
endmodule


