//Key = 1010111001101001011001110100010000010001100101110111010011110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276;

XOR2_X1 U702 ( .A(n969), .B(n970), .Z(G9) );
NOR2_X1 U703 ( .A1(KEYINPUT30), .A2(n971), .ZN(n970) );
NOR2_X1 U704 ( .A1(n972), .A2(n973), .ZN(n969) );
NOR2_X1 U705 ( .A1(n974), .A2(n975), .ZN(G75) );
NOR4_X1 U706 ( .A1(n976), .A2(n977), .A3(G953), .A4(n978), .ZN(n975) );
AND3_X1 U707 ( .A1(n979), .A2(n980), .A3(n981), .ZN(n977) );
NAND3_X1 U708 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n976) );
XOR2_X1 U709 ( .A(n985), .B(KEYINPUT4), .Z(n984) );
NAND2_X1 U710 ( .A1(n986), .A2(n987), .ZN(n985) );
NAND3_X1 U711 ( .A1(n988), .A2(n980), .A3(n979), .ZN(n987) );
NAND3_X1 U712 ( .A1(n989), .A2(n990), .A3(n991), .ZN(n986) );
NAND2_X1 U713 ( .A1(n992), .A2(n993), .ZN(n990) );
NAND2_X1 U714 ( .A1(n994), .A2(n980), .ZN(n993) );
NAND2_X1 U715 ( .A1(n995), .A2(n996), .ZN(n992) );
NAND2_X1 U716 ( .A1(n997), .A2(n998), .ZN(n996) );
NAND2_X1 U717 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND2_X1 U718 ( .A1(n1001), .A2(n980), .ZN(n997) );
NAND2_X1 U719 ( .A1(n989), .A2(n1002), .ZN(n983) );
NAND2_X1 U720 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND3_X1 U721 ( .A1(n1005), .A2(n1006), .A3(n979), .ZN(n1004) );
AND3_X1 U722 ( .A1(n1000), .A2(n995), .A3(n991), .ZN(n979) );
NAND3_X1 U723 ( .A1(n1007), .A2(n1008), .A3(n980), .ZN(n1003) );
NAND2_X1 U724 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND4_X1 U725 ( .A1(n1011), .A2(n1012), .A3(n995), .A4(n1013), .ZN(n1009) );
INV_X1 U726 ( .A(KEYINPUT5), .ZN(n1013) );
NAND3_X1 U727 ( .A1(n1014), .A2(n1015), .A3(n991), .ZN(n1007) );
INV_X1 U728 ( .A(n1010), .ZN(n991) );
NAND4_X1 U729 ( .A1(KEYINPUT5), .A2(n1012), .A3(n1011), .A4(n995), .ZN(n1015) );
NAND3_X1 U730 ( .A1(n1016), .A2(n1000), .A3(n1017), .ZN(n1014) );
XOR2_X1 U731 ( .A(n1018), .B(KEYINPUT41), .Z(n1017) );
NOR3_X1 U732 ( .A1(n978), .A2(G953), .A3(G952), .ZN(n974) );
AND4_X1 U733 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n978) );
NOR4_X1 U734 ( .A1(n1012), .A2(n1023), .A3(n1006), .A4(n1024), .ZN(n1022) );
XOR2_X1 U735 ( .A(n1025), .B(KEYINPUT58), .Z(n1023) );
XOR2_X1 U736 ( .A(n1026), .B(n1027), .Z(n1021) );
NOR2_X1 U737 ( .A1(KEYINPUT1), .A2(n1028), .ZN(n1027) );
XOR2_X1 U738 ( .A(n1029), .B(G478), .Z(n1020) );
XOR2_X1 U739 ( .A(n1030), .B(G472), .Z(n1019) );
XOR2_X1 U740 ( .A(n1031), .B(n1032), .Z(G72) );
XOR2_X1 U741 ( .A(n1033), .B(n1034), .Z(n1032) );
NAND2_X1 U742 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U743 ( .A1(G953), .A2(n1037), .ZN(n1036) );
XOR2_X1 U744 ( .A(n1038), .B(n1039), .Z(n1035) );
XNOR2_X1 U745 ( .A(G140), .B(n1040), .ZN(n1039) );
NAND2_X1 U746 ( .A1(n1041), .A2(KEYINPUT35), .ZN(n1040) );
XNOR2_X1 U747 ( .A(n1042), .B(n1043), .ZN(n1041) );
XOR2_X1 U748 ( .A(n1044), .B(KEYINPUT18), .Z(n1042) );
NAND2_X1 U749 ( .A1(n1045), .A2(n1046), .ZN(n1033) );
NAND2_X1 U750 ( .A1(G900), .A2(G227), .ZN(n1046) );
AND2_X1 U751 ( .A1(n1047), .A2(n1048), .ZN(n1031) );
XOR2_X1 U752 ( .A(n1049), .B(n1050), .Z(G69) );
NOR2_X1 U753 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U754 ( .A(KEYINPUT20), .B(n1053), .Z(n1052) );
NOR2_X1 U755 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
AND2_X1 U756 ( .A1(n1055), .A2(n1054), .ZN(n1051) );
AND2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NAND2_X1 U758 ( .A1(G953), .A2(n1058), .ZN(n1057) );
XOR2_X1 U759 ( .A(n1059), .B(n1060), .Z(n1056) );
NOR2_X1 U760 ( .A1(KEYINPUT54), .A2(n1061), .ZN(n1059) );
NAND2_X1 U761 ( .A1(n1062), .A2(n1063), .ZN(n1055) );
XOR2_X1 U762 ( .A(n1048), .B(KEYINPUT37), .Z(n1062) );
NAND2_X1 U763 ( .A1(n1045), .A2(n1064), .ZN(n1049) );
NAND2_X1 U764 ( .A1(G898), .A2(G224), .ZN(n1064) );
XOR2_X1 U765 ( .A(G953), .B(KEYINPUT55), .Z(n1045) );
NOR2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(G66) );
XNOR2_X1 U767 ( .A(n1067), .B(n1068), .ZN(n1066) );
NOR2_X1 U768 ( .A1(KEYINPUT33), .A2(n1069), .ZN(n1068) );
NAND3_X1 U769 ( .A1(n1070), .A2(G217), .A3(KEYINPUT53), .ZN(n1067) );
NOR2_X1 U770 ( .A1(n1065), .A2(n1071), .ZN(G63) );
XOR2_X1 U771 ( .A(n1072), .B(n1073), .Z(n1071) );
NAND2_X1 U772 ( .A1(n1070), .A2(G478), .ZN(n1072) );
NOR2_X1 U773 ( .A1(n1065), .A2(n1074), .ZN(G60) );
XOR2_X1 U774 ( .A(n1075), .B(n1076), .Z(n1074) );
AND2_X1 U775 ( .A1(G475), .A2(n1070), .ZN(n1076) );
NAND2_X1 U776 ( .A1(KEYINPUT22), .A2(n1077), .ZN(n1075) );
XOR2_X1 U777 ( .A(G104), .B(n1078), .Z(G6) );
NOR2_X1 U778 ( .A1(n973), .A2(n1079), .ZN(n1078) );
NOR2_X1 U779 ( .A1(n1065), .A2(n1080), .ZN(G57) );
XOR2_X1 U780 ( .A(n1081), .B(n1082), .Z(n1080) );
XOR2_X1 U781 ( .A(n1083), .B(n1084), .Z(n1082) );
XOR2_X1 U782 ( .A(n1085), .B(n1086), .Z(n1081) );
NOR2_X1 U783 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U784 ( .A(KEYINPUT44), .B(n1089), .Z(n1088) );
NOR2_X1 U785 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
AND2_X1 U786 ( .A1(n1090), .A2(n1091), .ZN(n1087) );
NAND2_X1 U787 ( .A1(n1070), .A2(G472), .ZN(n1085) );
NOR2_X1 U788 ( .A1(n1065), .A2(n1092), .ZN(G54) );
XOR2_X1 U789 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND2_X1 U790 ( .A1(n1070), .A2(G469), .ZN(n1094) );
NAND3_X1 U791 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1093) );
OR2_X1 U792 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U793 ( .A1(KEYINPUT36), .A2(n1100), .ZN(n1096) );
NAND2_X1 U794 ( .A1(n1101), .A2(n1099), .ZN(n1100) );
XNOR2_X1 U795 ( .A(n1098), .B(KEYINPUT39), .ZN(n1101) );
NAND2_X1 U796 ( .A1(n1102), .A2(n1103), .ZN(n1095) );
INV_X1 U797 ( .A(KEYINPUT36), .ZN(n1103) );
NAND2_X1 U798 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
OR2_X1 U799 ( .A1(n1098), .A2(KEYINPUT39), .ZN(n1105) );
NAND3_X1 U800 ( .A1(n1098), .A2(n1099), .A3(KEYINPUT39), .ZN(n1104) );
XNOR2_X1 U801 ( .A(n1106), .B(n1107), .ZN(n1098) );
XOR2_X1 U802 ( .A(n1108), .B(n1109), .Z(n1106) );
NAND2_X1 U803 ( .A1(KEYINPUT57), .A2(n1110), .ZN(n1108) );
NOR2_X1 U804 ( .A1(n1111), .A2(n1112), .ZN(G51) );
XNOR2_X1 U805 ( .A(n1065), .B(KEYINPUT9), .ZN(n1112) );
NOR2_X1 U806 ( .A1(n1048), .A2(G952), .ZN(n1065) );
XOR2_X1 U807 ( .A(n1113), .B(n1114), .Z(n1111) );
NOR3_X1 U808 ( .A1(n1115), .A2(KEYINPUT3), .A3(n1116), .ZN(n1114) );
NAND2_X1 U809 ( .A1(n1070), .A2(n1117), .ZN(n1113) );
NOR2_X1 U810 ( .A1(n1118), .A2(n982), .ZN(n1070) );
NOR2_X1 U811 ( .A1(n1047), .A2(n1063), .ZN(n982) );
NAND4_X1 U812 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1063) );
NOR4_X1 U813 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n1122) );
INV_X1 U814 ( .A(n1127), .ZN(n1126) );
NAND2_X1 U815 ( .A1(n1001), .A2(n1128), .ZN(n1121) );
NAND2_X1 U816 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XNOR2_X1 U817 ( .A(KEYINPUT10), .B(n972), .ZN(n1130) );
NAND2_X1 U818 ( .A1(n1131), .A2(n981), .ZN(n972) );
XOR2_X1 U819 ( .A(n1079), .B(KEYINPUT32), .Z(n1129) );
NAND2_X1 U820 ( .A1(n988), .A2(n1131), .ZN(n1079) );
AND3_X1 U821 ( .A1(n1132), .A2(n1133), .A3(n980), .ZN(n1131) );
NAND4_X1 U822 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1047) );
NOR4_X1 U823 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1137) );
INV_X1 U824 ( .A(n1142), .ZN(n1140) );
NOR3_X1 U825 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1136) );
NOR3_X1 U826 ( .A1(n973), .A2(n1146), .A3(n1147), .ZN(n1145) );
XOR2_X1 U827 ( .A(KEYINPUT17), .B(n995), .Z(n1146) );
AND4_X1 U828 ( .A1(n973), .A2(n988), .A3(n1148), .A4(n1149), .ZN(n1144) );
NOR2_X1 U829 ( .A1(n1150), .A2(n1148), .ZN(n1143) );
INV_X1 U830 ( .A(KEYINPUT47), .ZN(n1148) );
NAND3_X1 U831 ( .A1(n1025), .A2(n994), .A3(n1151), .ZN(n1134) );
XOR2_X1 U832 ( .A(n1150), .B(n1152), .Z(G48) );
NAND2_X1 U833 ( .A1(KEYINPUT43), .A2(G146), .ZN(n1152) );
NAND3_X1 U834 ( .A1(n1149), .A2(n1001), .A3(n988), .ZN(n1150) );
XNOR2_X1 U835 ( .A(G143), .B(n1135), .ZN(G45) );
NAND4_X1 U836 ( .A1(n1151), .A2(n1001), .A3(n1132), .A4(n1153), .ZN(n1135) );
XOR2_X1 U837 ( .A(G140), .B(n1141), .Z(G42) );
NOR2_X1 U838 ( .A1(n1147), .A2(n1154), .ZN(n1141) );
NAND3_X1 U839 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(G39) );
OR2_X1 U840 ( .A1(n1142), .A2(KEYINPUT46), .ZN(n1157) );
NAND3_X1 U841 ( .A1(KEYINPUT46), .A2(n1142), .A3(G137), .ZN(n1156) );
NAND2_X1 U842 ( .A1(n1158), .A2(n1044), .ZN(n1155) );
NAND2_X1 U843 ( .A1(n1159), .A2(KEYINPUT46), .ZN(n1158) );
XOR2_X1 U844 ( .A(n1142), .B(KEYINPUT48), .Z(n1159) );
NAND3_X1 U845 ( .A1(n1000), .A2(n1149), .A3(n989), .ZN(n1142) );
INV_X1 U846 ( .A(n1160), .ZN(n1149) );
XOR2_X1 U847 ( .A(n1161), .B(n1162), .Z(G36) );
NAND4_X1 U848 ( .A1(n1151), .A2(n1000), .A3(n1025), .A4(n1163), .ZN(n1162) );
XOR2_X1 U849 ( .A(KEYINPUT28), .B(n1132), .Z(n1163) );
AND3_X1 U850 ( .A1(n1164), .A2(n1165), .A3(n999), .ZN(n1151) );
XNOR2_X1 U851 ( .A(n1139), .B(n1166), .ZN(G33) );
XOR2_X1 U852 ( .A(KEYINPUT49), .B(G131), .Z(n1166) );
AND4_X1 U853 ( .A1(n999), .A2(n988), .A3(n994), .A4(n1165), .ZN(n1139) );
INV_X1 U854 ( .A(n1154), .ZN(n994) );
NAND2_X1 U855 ( .A1(n1000), .A2(n1132), .ZN(n1154) );
AND2_X1 U856 ( .A1(n1011), .A2(n1167), .ZN(n1000) );
XOR2_X1 U857 ( .A(G128), .B(n1138), .Z(G30) );
NOR3_X1 U858 ( .A1(n973), .A2(n1168), .A3(n1160), .ZN(n1138) );
NAND4_X1 U859 ( .A1(n1132), .A2(n1169), .A3(n1165), .A4(n1006), .ZN(n1160) );
XOR2_X1 U860 ( .A(G101), .B(n1125), .Z(G3) );
AND2_X1 U861 ( .A1(n1170), .A2(n999), .ZN(n1125) );
XOR2_X1 U862 ( .A(G125), .B(n1171), .Z(G27) );
NOR3_X1 U863 ( .A1(n1147), .A2(n973), .A3(n1024), .ZN(n1171) );
INV_X1 U864 ( .A(n995), .ZN(n1024) );
INV_X1 U865 ( .A(n1001), .ZN(n973) );
NAND4_X1 U866 ( .A1(n1005), .A2(n988), .A3(n1165), .A4(n1006), .ZN(n1147) );
NAND2_X1 U867 ( .A1(n1010), .A2(n1172), .ZN(n1165) );
NAND4_X1 U868 ( .A1(G902), .A2(G953), .A3(n1173), .A4(n1037), .ZN(n1172) );
INV_X1 U869 ( .A(G900), .ZN(n1037) );
XNOR2_X1 U870 ( .A(G122), .B(n1119), .ZN(G24) );
NAND4_X1 U871 ( .A1(n1164), .A2(n1174), .A3(n980), .A4(n1153), .ZN(n1119) );
NOR2_X1 U872 ( .A1(n1006), .A2(n1169), .ZN(n980) );
XOR2_X1 U873 ( .A(n1175), .B(n1120), .Z(G21) );
NAND4_X1 U874 ( .A1(n1174), .A2(n989), .A3(n1169), .A4(n1006), .ZN(n1120) );
INV_X1 U875 ( .A(n1005), .ZN(n1169) );
XOR2_X1 U876 ( .A(G116), .B(n1124), .Z(G18) );
AND3_X1 U877 ( .A1(n999), .A2(n981), .A3(n1174), .ZN(n1124) );
INV_X1 U878 ( .A(n1168), .ZN(n981) );
NAND2_X1 U879 ( .A1(n1164), .A2(n1025), .ZN(n1168) );
NAND2_X1 U880 ( .A1(n1176), .A2(n1177), .ZN(G15) );
NAND2_X1 U881 ( .A1(G113), .A2(n1127), .ZN(n1177) );
XOR2_X1 U882 ( .A(KEYINPUT25), .B(n1178), .Z(n1176) );
NOR2_X1 U883 ( .A1(G113), .A2(n1127), .ZN(n1178) );
NAND3_X1 U884 ( .A1(n999), .A2(n988), .A3(n1174), .ZN(n1127) );
AND3_X1 U885 ( .A1(n1001), .A2(n1133), .A3(n995), .ZN(n1174) );
NOR2_X1 U886 ( .A1(n1179), .A2(n1016), .ZN(n995) );
INV_X1 U887 ( .A(n1018), .ZN(n1179) );
NOR2_X1 U888 ( .A1(n1025), .A2(n1164), .ZN(n988) );
NOR2_X1 U889 ( .A1(n1006), .A2(n1005), .ZN(n999) );
XOR2_X1 U890 ( .A(n1123), .B(n1180), .Z(G12) );
XOR2_X1 U891 ( .A(KEYINPUT19), .B(G110), .Z(n1180) );
AND3_X1 U892 ( .A1(n1005), .A2(n1006), .A3(n1170), .ZN(n1123) );
AND4_X1 U893 ( .A1(n989), .A2(n1001), .A3(n1132), .A4(n1133), .ZN(n1170) );
NAND2_X1 U894 ( .A1(n1010), .A2(n1181), .ZN(n1133) );
NAND4_X1 U895 ( .A1(G902), .A2(G953), .A3(n1173), .A4(n1058), .ZN(n1181) );
INV_X1 U896 ( .A(G898), .ZN(n1058) );
NAND3_X1 U897 ( .A1(n1173), .A2(n1048), .A3(G952), .ZN(n1010) );
NAND2_X1 U898 ( .A1(G234), .A2(G237), .ZN(n1173) );
NOR2_X1 U899 ( .A1(n1018), .A2(n1016), .ZN(n1132) );
AND2_X1 U900 ( .A1(G221), .A2(n1182), .ZN(n1016) );
NAND2_X1 U901 ( .A1(G234), .A2(n1118), .ZN(n1182) );
XOR2_X1 U902 ( .A(n1183), .B(G469), .Z(n1018) );
NAND2_X1 U903 ( .A1(n1184), .A2(n1118), .ZN(n1183) );
XNOR2_X1 U904 ( .A(n1185), .B(n1099), .ZN(n1184) );
XNOR2_X1 U905 ( .A(n1186), .B(n1187), .ZN(n1099) );
NAND2_X1 U906 ( .A1(G227), .A2(n1048), .ZN(n1186) );
NAND2_X1 U907 ( .A1(KEYINPUT51), .A2(n1188), .ZN(n1185) );
XOR2_X1 U908 ( .A(n1189), .B(n1107), .Z(n1188) );
NAND2_X1 U909 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND2_X1 U910 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U911 ( .A(KEYINPUT14), .B(n1194), .Z(n1192) );
NAND2_X1 U912 ( .A1(n1109), .A2(n1195), .ZN(n1190) );
XNOR2_X1 U913 ( .A(n1194), .B(KEYINPUT34), .ZN(n1195) );
NOR2_X1 U914 ( .A1(KEYINPUT42), .A2(n1110), .ZN(n1194) );
INV_X1 U915 ( .A(n1193), .ZN(n1109) );
XOR2_X1 U916 ( .A(n1083), .B(n1196), .Z(n1193) );
NOR2_X1 U917 ( .A1(n1011), .A2(n1012), .ZN(n1001) );
INV_X1 U918 ( .A(n1167), .ZN(n1012) );
NAND2_X1 U919 ( .A1(G214), .A2(n1197), .ZN(n1167) );
XNOR2_X1 U920 ( .A(n1198), .B(n1117), .ZN(n1011) );
INV_X1 U921 ( .A(n1026), .ZN(n1117) );
NAND2_X1 U922 ( .A1(G210), .A2(n1197), .ZN(n1026) );
NAND2_X1 U923 ( .A1(n1199), .A2(n1118), .ZN(n1197) );
XOR2_X1 U924 ( .A(KEYINPUT63), .B(G237), .Z(n1199) );
NAND2_X1 U925 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
NAND2_X1 U926 ( .A1(KEYINPUT38), .A2(n1028), .ZN(n1201) );
INV_X1 U927 ( .A(n1202), .ZN(n1028) );
NAND2_X1 U928 ( .A1(KEYINPUT45), .A2(n1202), .ZN(n1200) );
NOR3_X1 U929 ( .A1(n1116), .A2(G902), .A3(n1203), .ZN(n1202) );
XNOR2_X1 U930 ( .A(KEYINPUT2), .B(n1115), .ZN(n1203) );
AND2_X1 U931 ( .A1(n1204), .A2(n1205), .ZN(n1115) );
NOR2_X1 U932 ( .A1(n1205), .A2(n1204), .ZN(n1116) );
XOR2_X1 U933 ( .A(n1060), .B(n1061), .Z(n1204) );
XNOR2_X1 U934 ( .A(n1206), .B(n1207), .ZN(n1061) );
XOR2_X1 U935 ( .A(n1208), .B(KEYINPUT13), .Z(n1206) );
INV_X1 U936 ( .A(G110), .ZN(n1208) );
XNOR2_X1 U937 ( .A(n1209), .B(n1210), .ZN(n1060) );
XOR2_X1 U938 ( .A(G113), .B(n1211), .Z(n1210) );
XOR2_X1 U939 ( .A(G119), .B(G116), .Z(n1211) );
XOR2_X1 U940 ( .A(n1083), .B(n1212), .Z(n1209) );
NOR2_X1 U941 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
AND3_X1 U942 ( .A1(KEYINPUT31), .A2(n971), .A3(G104), .ZN(n1214) );
NOR2_X1 U943 ( .A1(KEYINPUT31), .A2(n1196), .ZN(n1213) );
XOR2_X1 U944 ( .A(G104), .B(G107), .Z(n1196) );
XNOR2_X1 U945 ( .A(n1215), .B(n1216), .ZN(n1205) );
INV_X1 U946 ( .A(n1038), .ZN(n1216) );
XOR2_X1 U947 ( .A(n1217), .B(G125), .Z(n1038) );
NAND2_X1 U948 ( .A1(G224), .A2(n1048), .ZN(n1215) );
NOR2_X1 U949 ( .A1(n1153), .A2(n1164), .ZN(n989) );
XNOR2_X1 U950 ( .A(n1218), .B(n1029), .ZN(n1164) );
NAND2_X1 U951 ( .A1(n1073), .A2(n1219), .ZN(n1029) );
XOR2_X1 U952 ( .A(KEYINPUT29), .B(G902), .Z(n1219) );
XOR2_X1 U953 ( .A(n1220), .B(n1221), .Z(n1073) );
NOR3_X1 U954 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1221) );
XOR2_X1 U955 ( .A(n1048), .B(KEYINPUT21), .Z(n1224) );
NAND2_X1 U956 ( .A1(n1225), .A2(KEYINPUT23), .ZN(n1220) );
XOR2_X1 U957 ( .A(n1226), .B(n1227), .Z(n1225) );
XOR2_X1 U958 ( .A(n1207), .B(n1228), .Z(n1227) );
XOR2_X1 U959 ( .A(n971), .B(n1229), .Z(n1226) );
XOR2_X1 U960 ( .A(G134), .B(G116), .Z(n1229) );
INV_X1 U961 ( .A(G107), .ZN(n971) );
NAND2_X1 U962 ( .A1(KEYINPUT0), .A2(n1230), .ZN(n1218) );
INV_X1 U963 ( .A(G478), .ZN(n1230) );
INV_X1 U964 ( .A(n1025), .ZN(n1153) );
XOR2_X1 U965 ( .A(n1231), .B(G475), .Z(n1025) );
NAND2_X1 U966 ( .A1(n1077), .A2(n1118), .ZN(n1231) );
XNOR2_X1 U967 ( .A(n1232), .B(n1233), .ZN(n1077) );
XOR2_X1 U968 ( .A(n1234), .B(n1235), .Z(n1233) );
XNOR2_X1 U969 ( .A(n1236), .B(n1237), .ZN(n1235) );
NAND2_X1 U970 ( .A1(KEYINPUT59), .A2(n1238), .ZN(n1237) );
XOR2_X1 U971 ( .A(G113), .B(n1207), .Z(n1238) );
XOR2_X1 U972 ( .A(G122), .B(KEYINPUT8), .Z(n1207) );
NAND2_X1 U973 ( .A1(KEYINPUT56), .A2(G140), .ZN(n1236) );
XOR2_X1 U974 ( .A(n1239), .B(n1240), .Z(n1232) );
XOR2_X1 U975 ( .A(G104), .B(n1241), .Z(n1240) );
AND3_X1 U976 ( .A1(G214), .A2(n1048), .A3(n1242), .ZN(n1241) );
XNOR2_X1 U977 ( .A(G131), .B(G143), .ZN(n1239) );
NAND3_X1 U978 ( .A1(n1243), .A2(n1244), .A3(n1245), .ZN(n1006) );
NAND2_X1 U979 ( .A1(G902), .A2(G217), .ZN(n1245) );
OR3_X1 U980 ( .A1(n1246), .A2(G902), .A3(n1247), .ZN(n1244) );
NAND2_X1 U981 ( .A1(n1247), .A2(n1246), .ZN(n1243) );
INV_X1 U982 ( .A(n1069), .ZN(n1246) );
XOR2_X1 U983 ( .A(n1248), .B(n1249), .Z(n1069) );
XOR2_X1 U984 ( .A(n1250), .B(n1251), .Z(n1249) );
XOR2_X1 U985 ( .A(n1252), .B(n1187), .Z(n1251) );
XOR2_X1 U986 ( .A(G110), .B(G140), .Z(n1187) );
INV_X1 U987 ( .A(n1234), .ZN(n1252) );
XNOR2_X1 U988 ( .A(G125), .B(G146), .ZN(n1234) );
XOR2_X1 U989 ( .A(n1253), .B(n1254), .Z(n1250) );
NAND2_X1 U990 ( .A1(KEYINPUT6), .A2(G137), .ZN(n1254) );
NAND3_X1 U991 ( .A1(G221), .A2(n1255), .A3(n1256), .ZN(n1253) );
XOR2_X1 U992 ( .A(n1048), .B(KEYINPUT26), .Z(n1256) );
INV_X1 U993 ( .A(n1223), .ZN(n1255) );
XNOR2_X1 U994 ( .A(G234), .B(KEYINPUT61), .ZN(n1223) );
XOR2_X1 U995 ( .A(n1257), .B(n1258), .Z(n1248) );
XOR2_X1 U996 ( .A(G128), .B(G119), .Z(n1258) );
XNOR2_X1 U997 ( .A(KEYINPUT15), .B(KEYINPUT11), .ZN(n1257) );
NOR2_X1 U998 ( .A1(n1222), .A2(G234), .ZN(n1247) );
INV_X1 U999 ( .A(G217), .ZN(n1222) );
XOR2_X1 U1000 ( .A(n1030), .B(n1259), .Z(n1005) );
XOR2_X1 U1001 ( .A(KEYINPUT40), .B(n1260), .Z(n1259) );
NOR2_X1 U1002 ( .A1(KEYINPUT27), .A2(G472), .ZN(n1260) );
NAND2_X1 U1003 ( .A1(n1261), .A2(n1118), .ZN(n1030) );
INV_X1 U1004 ( .A(G902), .ZN(n1118) );
XOR2_X1 U1005 ( .A(n1262), .B(n1263), .Z(n1261) );
XNOR2_X1 U1006 ( .A(n1084), .B(n1091), .ZN(n1263) );
XNOR2_X1 U1007 ( .A(n1264), .B(n1265), .ZN(n1091) );
NOR2_X1 U1008 ( .A1(G113), .A2(KEYINPUT16), .ZN(n1265) );
NAND2_X1 U1009 ( .A1(n1266), .A2(n1267), .ZN(n1264) );
NAND2_X1 U1010 ( .A1(G116), .A2(n1175), .ZN(n1267) );
XOR2_X1 U1011 ( .A(KEYINPUT50), .B(n1268), .Z(n1266) );
NOR2_X1 U1012 ( .A1(G116), .A2(n1175), .ZN(n1268) );
INV_X1 U1013 ( .A(G119), .ZN(n1175) );
NAND3_X1 U1014 ( .A1(n1242), .A2(n1048), .A3(G210), .ZN(n1084) );
INV_X1 U1015 ( .A(G953), .ZN(n1048) );
INV_X1 U1016 ( .A(G237), .ZN(n1242) );
XOR2_X1 U1017 ( .A(n1269), .B(n1270), .Z(n1262) );
XNOR2_X1 U1018 ( .A(KEYINPUT60), .B(n1271), .ZN(n1270) );
NOR2_X1 U1019 ( .A1(KEYINPUT62), .A2(n1090), .ZN(n1271) );
XNOR2_X1 U1020 ( .A(n1107), .B(n1110), .ZN(n1090) );
AND2_X1 U1021 ( .A1(n1272), .A2(n1273), .ZN(n1110) );
NAND2_X1 U1022 ( .A1(n1043), .A2(G137), .ZN(n1273) );
NAND2_X1 U1023 ( .A1(n1274), .A2(n1044), .ZN(n1272) );
INV_X1 U1024 ( .A(G137), .ZN(n1044) );
XNOR2_X1 U1025 ( .A(KEYINPUT52), .B(n1043), .ZN(n1274) );
XOR2_X1 U1026 ( .A(G131), .B(n1161), .Z(n1043) );
INV_X1 U1027 ( .A(G134), .ZN(n1161) );
INV_X1 U1028 ( .A(n1217), .ZN(n1107) );
XOR2_X1 U1029 ( .A(n1275), .B(n1276), .Z(n1217) );
XOR2_X1 U1030 ( .A(KEYINPUT7), .B(KEYINPUT24), .Z(n1276) );
XNOR2_X1 U1031 ( .A(G146), .B(n1228), .ZN(n1275) );
XOR2_X1 U1032 ( .A(G128), .B(G143), .Z(n1228) );
NAND2_X1 U1033 ( .A1(KEYINPUT12), .A2(n1083), .ZN(n1269) );
INV_X1 U1034 ( .A(G101), .ZN(n1083) );
endmodule


