//Key = 0110010110111001010100000001100001100000000001100110111100110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319;

XNOR2_X1 U731 ( .A(G107), .B(n1005), .ZN(G9) );
NAND2_X1 U732 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
XNOR2_X1 U733 ( .A(KEYINPUT36), .B(n1008), .ZN(n1007) );
NOR2_X1 U734 ( .A1(n1009), .A2(n1010), .ZN(G75) );
NOR4_X1 U735 ( .A1(G953), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1010) );
XOR2_X1 U736 ( .A(KEYINPUT2), .B(n1014), .Z(n1013) );
NOR2_X1 U737 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NOR4_X1 U738 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
XOR2_X1 U739 ( .A(n1021), .B(KEYINPUT48), .Z(n1017) );
NOR3_X1 U740 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1015) );
NOR2_X1 U741 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR3_X1 U742 ( .A1(n1019), .A2(n1026), .A3(n1027), .ZN(n1025) );
NOR3_X1 U743 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
NOR2_X1 U744 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U745 ( .A1(n1033), .A2(n1006), .ZN(n1031) );
NOR2_X1 U746 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR2_X1 U747 ( .A1(n1036), .A2(n1020), .ZN(n1029) );
NOR2_X1 U748 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
AND2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR2_X1 U750 ( .A1(n1041), .A2(n1042), .ZN(n1026) );
NOR2_X1 U751 ( .A1(n1043), .A2(n1032), .ZN(n1041) );
XNOR2_X1 U752 ( .A(n1044), .B(KEYINPUT61), .ZN(n1043) );
NOR4_X1 U753 ( .A1(n1028), .A2(n1045), .A3(n1032), .A4(n1020), .ZN(n1024) );
INV_X1 U754 ( .A(n1046), .ZN(n1032) );
NOR2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR3_X1 U756 ( .A1(n1011), .A2(G953), .A3(G952), .ZN(n1009) );
AND4_X1 U757 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1011) );
NOR4_X1 U758 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
INV_X1 U759 ( .A(n1057), .ZN(n1054) );
NAND2_X1 U760 ( .A1(n1058), .A2(n1059), .ZN(n1053) );
NAND2_X1 U761 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
XNOR2_X1 U762 ( .A(G472), .B(KEYINPUT8), .ZN(n1060) );
NOR3_X1 U763 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1051) );
XOR2_X1 U764 ( .A(n1065), .B(n1066), .Z(n1064) );
XNOR2_X1 U765 ( .A(KEYINPUT11), .B(n1067), .ZN(n1066) );
XNOR2_X1 U766 ( .A(n1028), .B(KEYINPUT27), .ZN(n1063) );
XOR2_X1 U767 ( .A(n1068), .B(KEYINPUT19), .Z(n1050) );
NAND3_X1 U768 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1068) );
NAND2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U770 ( .A1(KEYINPUT30), .A2(n1074), .ZN(n1070) );
NAND2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
XNOR2_X1 U772 ( .A(n1072), .B(KEYINPUT25), .ZN(n1075) );
NAND2_X1 U773 ( .A1(n1077), .A2(n1078), .ZN(n1069) );
INV_X1 U774 ( .A(KEYINPUT30), .ZN(n1078) );
NAND2_X1 U775 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
OR3_X1 U776 ( .A1(n1073), .A2(n1072), .A3(KEYINPUT25), .ZN(n1080) );
INV_X1 U777 ( .A(n1076), .ZN(n1073) );
NAND2_X1 U778 ( .A1(KEYINPUT25), .A2(n1072), .ZN(n1079) );
XNOR2_X1 U779 ( .A(n1023), .B(KEYINPUT4), .ZN(n1049) );
XOR2_X1 U780 ( .A(n1081), .B(n1082), .Z(G72) );
NOR2_X1 U781 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U782 ( .A(n1085), .B(KEYINPUT50), .Z(n1083) );
NAND2_X1 U783 ( .A1(G900), .A2(G227), .ZN(n1085) );
NAND2_X1 U784 ( .A1(n1086), .A2(n1087), .ZN(n1081) );
NAND3_X1 U785 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1087) );
INV_X1 U786 ( .A(n1091), .ZN(n1089) );
OR2_X1 U787 ( .A1(n1088), .A2(n1090), .ZN(n1086) );
NAND2_X1 U788 ( .A1(n1084), .A2(n1092), .ZN(n1090) );
NAND2_X1 U789 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U790 ( .A(n1095), .B(n1096), .Z(n1088) );
XNOR2_X1 U791 ( .A(n1097), .B(n1098), .ZN(n1096) );
XNOR2_X1 U792 ( .A(G131), .B(n1099), .ZN(n1095) );
NOR2_X1 U793 ( .A1(KEYINPUT35), .A2(n1100), .ZN(n1099) );
XNOR2_X1 U794 ( .A(G137), .B(n1101), .ZN(n1100) );
NAND2_X1 U795 ( .A1(KEYINPUT7), .A2(n1102), .ZN(n1101) );
XOR2_X1 U796 ( .A(n1103), .B(n1104), .Z(G69) );
NOR2_X1 U797 ( .A1(n1105), .A2(n1084), .ZN(n1104) );
AND2_X1 U798 ( .A1(G224), .A2(G898), .ZN(n1105) );
NAND2_X1 U799 ( .A1(n1106), .A2(n1107), .ZN(n1103) );
NAND2_X1 U800 ( .A1(n1108), .A2(n1084), .ZN(n1107) );
XNOR2_X1 U801 ( .A(n1109), .B(n1110), .ZN(n1108) );
OR3_X1 U802 ( .A1(n1111), .A2(n1112), .A3(n1084), .ZN(n1106) );
INV_X1 U803 ( .A(n1109), .ZN(n1111) );
NOR2_X1 U804 ( .A1(n1113), .A2(n1114), .ZN(G66) );
NOR3_X1 U805 ( .A1(n1076), .A2(n1115), .A3(n1116), .ZN(n1114) );
NOR3_X1 U806 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1116) );
NOR2_X1 U807 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
AND2_X1 U808 ( .A1(n1012), .A2(n1072), .ZN(n1120) );
INV_X1 U809 ( .A(n1118), .ZN(n1072) );
NOR2_X1 U810 ( .A1(n1113), .A2(n1122), .ZN(G63) );
XOR2_X1 U811 ( .A(n1123), .B(n1124), .Z(n1122) );
AND2_X1 U812 ( .A1(G478), .A2(n1125), .ZN(n1123) );
NOR2_X1 U813 ( .A1(n1113), .A2(n1126), .ZN(G60) );
XNOR2_X1 U814 ( .A(n1127), .B(n1128), .ZN(n1126) );
AND2_X1 U815 ( .A1(G475), .A2(n1125), .ZN(n1128) );
XNOR2_X1 U816 ( .A(G104), .B(n1129), .ZN(G6) );
NOR2_X1 U817 ( .A1(n1113), .A2(n1130), .ZN(G57) );
XNOR2_X1 U818 ( .A(n1131), .B(n1132), .ZN(n1130) );
NAND2_X1 U819 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
XOR2_X1 U820 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U821 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U822 ( .A1(KEYINPUT44), .A2(n1139), .ZN(n1138) );
AND2_X1 U823 ( .A1(G472), .A2(n1125), .ZN(n1137) );
XNOR2_X1 U824 ( .A(KEYINPUT56), .B(KEYINPUT40), .ZN(n1133) );
NOR2_X1 U825 ( .A1(n1113), .A2(n1140), .ZN(G54) );
XOR2_X1 U826 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U827 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U828 ( .A1(KEYINPUT34), .A2(n1145), .ZN(n1144) );
NAND3_X1 U829 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1143) );
OR3_X1 U830 ( .A1(n1149), .A2(n1150), .A3(KEYINPUT3), .ZN(n1147) );
NAND2_X1 U831 ( .A1(KEYINPUT3), .A2(n1150), .ZN(n1146) );
XOR2_X1 U832 ( .A(n1151), .B(n1152), .Z(n1141) );
NAND2_X1 U833 ( .A1(n1125), .A2(G469), .ZN(n1151) );
INV_X1 U834 ( .A(n1119), .ZN(n1125) );
NOR2_X1 U835 ( .A1(n1153), .A2(n1154), .ZN(G51) );
XOR2_X1 U836 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U837 ( .A1(n1067), .A2(n1119), .ZN(n1156) );
NAND2_X1 U838 ( .A1(G902), .A2(n1012), .ZN(n1119) );
NAND3_X1 U839 ( .A1(n1093), .A2(n1157), .A3(n1110), .ZN(n1012) );
AND2_X1 U840 ( .A1(n1158), .A2(n1159), .ZN(n1110) );
NOR4_X1 U841 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1159) );
INV_X1 U842 ( .A(n1164), .ZN(n1160) );
AND4_X1 U843 ( .A1(n1165), .A2(n1166), .A3(n1129), .A4(n1167), .ZN(n1158) );
OR2_X1 U844 ( .A1(n1008), .A2(n1168), .ZN(n1167) );
NAND3_X1 U845 ( .A1(n1169), .A2(n1170), .A3(n1047), .ZN(n1008) );
INV_X1 U846 ( .A(n1018), .ZN(n1169) );
NAND2_X1 U847 ( .A1(n1046), .A2(n1171), .ZN(n1018) );
NAND3_X1 U848 ( .A1(n1172), .A2(n1046), .A3(n1048), .ZN(n1129) );
XOR2_X1 U849 ( .A(KEYINPUT32), .B(n1094), .Z(n1157) );
AND4_X1 U850 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1094) );
NAND3_X1 U851 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1173) );
XNOR2_X1 U852 ( .A(n1044), .B(KEYINPUT58), .ZN(n1179) );
AND4_X1 U853 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1093) );
NOR2_X1 U854 ( .A1(KEYINPUT62), .A2(n1184), .ZN(n1155) );
XOR2_X1 U855 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U856 ( .A1(KEYINPUT31), .A2(n1109), .ZN(n1186) );
NAND2_X1 U857 ( .A1(n1187), .A2(n1188), .ZN(n1185) );
NAND2_X1 U858 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U859 ( .A(n1191), .B(KEYINPUT16), .Z(n1187) );
OR2_X1 U860 ( .A1(n1189), .A2(n1190), .ZN(n1191) );
XNOR2_X1 U861 ( .A(n1113), .B(KEYINPUT1), .ZN(n1153) );
NOR2_X1 U862 ( .A1(n1084), .A2(G952), .ZN(n1113) );
XNOR2_X1 U863 ( .A(G146), .B(n1174), .ZN(G48) );
NAND3_X1 U864 ( .A1(n1048), .A2(n1006), .A3(n1177), .ZN(n1174) );
XNOR2_X1 U865 ( .A(G143), .B(n1175), .ZN(G45) );
NAND3_X1 U866 ( .A1(n1192), .A2(n1038), .A3(n1193), .ZN(n1175) );
NOR3_X1 U867 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1193) );
XNOR2_X1 U868 ( .A(G140), .B(n1176), .ZN(G42) );
NAND2_X1 U869 ( .A1(n1197), .A2(n1198), .ZN(n1176) );
XNOR2_X1 U870 ( .A(n1199), .B(n1200), .ZN(G39) );
NOR3_X1 U871 ( .A1(n1020), .A2(n1019), .A3(n1201), .ZN(n1200) );
INV_X1 U872 ( .A(n1178), .ZN(n1019) );
INV_X1 U873 ( .A(n1044), .ZN(n1020) );
XNOR2_X1 U874 ( .A(n1102), .B(n1202), .ZN(G36) );
NOR2_X1 U875 ( .A1(KEYINPUT29), .A2(n1180), .ZN(n1202) );
NAND3_X1 U876 ( .A1(n1038), .A2(n1047), .A3(n1197), .ZN(n1180) );
XOR2_X1 U877 ( .A(n1181), .B(n1203), .Z(G33) );
XNOR2_X1 U878 ( .A(KEYINPUT10), .B(n1204), .ZN(n1203) );
NAND3_X1 U879 ( .A1(n1048), .A2(n1038), .A3(n1197), .ZN(n1181) );
AND3_X1 U880 ( .A1(n1171), .A2(n1205), .A3(n1044), .ZN(n1197) );
NOR2_X1 U881 ( .A1(n1034), .A2(n1055), .ZN(n1044) );
INV_X1 U882 ( .A(n1035), .ZN(n1055) );
XOR2_X1 U883 ( .A(n1182), .B(n1206), .Z(G30) );
NAND2_X1 U884 ( .A1(KEYINPUT52), .A2(G128), .ZN(n1206) );
NAND3_X1 U885 ( .A1(n1006), .A2(n1047), .A3(n1177), .ZN(n1182) );
INV_X1 U886 ( .A(n1201), .ZN(n1177) );
NAND4_X1 U887 ( .A1(n1171), .A2(n1039), .A3(n1205), .A4(n1207), .ZN(n1201) );
XNOR2_X1 U888 ( .A(G101), .B(n1166), .ZN(G3) );
NAND3_X1 U889 ( .A1(n1172), .A2(n1178), .A3(n1038), .ZN(n1166) );
XOR2_X1 U890 ( .A(n1183), .B(n1208), .Z(G27) );
NOR2_X1 U891 ( .A1(G125), .A2(KEYINPUT41), .ZN(n1208) );
NAND3_X1 U892 ( .A1(n1194), .A2(n1198), .A3(n1192), .ZN(n1183) );
AND3_X1 U893 ( .A1(n1205), .A2(n1042), .A3(n1006), .ZN(n1192) );
NAND2_X1 U894 ( .A1(n1021), .A2(n1209), .ZN(n1205) );
NAND3_X1 U895 ( .A1(G902), .A2(n1210), .A3(n1091), .ZN(n1209) );
NOR2_X1 U896 ( .A1(n1084), .A2(G900), .ZN(n1091) );
AND3_X1 U897 ( .A1(n1040), .A2(n1039), .A3(n1048), .ZN(n1198) );
XNOR2_X1 U898 ( .A(G122), .B(n1165), .ZN(G24) );
NAND4_X1 U899 ( .A1(n1211), .A2(n1046), .A3(n1062), .A4(n1212), .ZN(n1165) );
NOR2_X1 U900 ( .A1(n1207), .A2(n1039), .ZN(n1046) );
XOR2_X1 U901 ( .A(G119), .B(n1163), .Z(G21) );
AND4_X1 U902 ( .A1(n1211), .A2(n1178), .A3(n1039), .A4(n1207), .ZN(n1163) );
XNOR2_X1 U903 ( .A(n1213), .B(n1162), .ZN(G18) );
AND3_X1 U904 ( .A1(n1038), .A2(n1047), .A3(n1211), .ZN(n1162) );
NOR2_X1 U905 ( .A1(n1062), .A2(n1195), .ZN(n1047) );
INV_X1 U906 ( .A(n1212), .ZN(n1195) );
XOR2_X1 U907 ( .A(G113), .B(n1161), .Z(G15) );
AND3_X1 U908 ( .A1(n1048), .A2(n1038), .A3(n1211), .ZN(n1161) );
AND4_X1 U909 ( .A1(n1194), .A2(n1006), .A3(n1042), .A4(n1170), .ZN(n1211) );
NOR2_X1 U910 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U911 ( .A1(n1212), .A2(n1196), .ZN(n1048) );
INV_X1 U912 ( .A(n1062), .ZN(n1196) );
XNOR2_X1 U913 ( .A(G110), .B(n1164), .ZN(G12) );
NAND4_X1 U914 ( .A1(n1172), .A2(n1178), .A3(n1040), .A4(n1039), .ZN(n1164) );
XOR2_X1 U915 ( .A(n1214), .B(n1118), .Z(n1039) );
NAND2_X1 U916 ( .A1(G217), .A2(n1215), .ZN(n1118) );
XNOR2_X1 U917 ( .A(n1076), .B(KEYINPUT39), .ZN(n1214) );
NOR2_X1 U918 ( .A1(n1121), .A2(G902), .ZN(n1076) );
INV_X1 U919 ( .A(n1117), .ZN(n1121) );
XNOR2_X1 U920 ( .A(n1216), .B(n1217), .ZN(n1117) );
XOR2_X1 U921 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U922 ( .A(G128), .B(G119), .Z(n1219) );
XNOR2_X1 U923 ( .A(KEYINPUT0), .B(n1199), .ZN(n1218) );
INV_X1 U924 ( .A(G137), .ZN(n1199) );
XOR2_X1 U925 ( .A(n1220), .B(n1221), .Z(n1216) );
XNOR2_X1 U926 ( .A(G110), .B(n1222), .ZN(n1221) );
NAND3_X1 U927 ( .A1(n1223), .A2(n1084), .A3(G221), .ZN(n1222) );
NAND2_X1 U928 ( .A1(n1224), .A2(KEYINPUT33), .ZN(n1220) );
XOR2_X1 U929 ( .A(n1225), .B(n1098), .Z(n1224) );
INV_X1 U930 ( .A(n1207), .ZN(n1040) );
NAND2_X1 U931 ( .A1(n1059), .A2(n1226), .ZN(n1207) );
NAND2_X1 U932 ( .A1(G472), .A2(n1061), .ZN(n1226) );
OR2_X1 U933 ( .A1(n1061), .A2(G472), .ZN(n1059) );
NAND2_X1 U934 ( .A1(n1227), .A2(n1228), .ZN(n1061) );
XOR2_X1 U935 ( .A(n1229), .B(n1230), .Z(n1227) );
XOR2_X1 U936 ( .A(n1139), .B(n1135), .Z(n1230) );
AND2_X1 U937 ( .A1(n1231), .A2(n1232), .ZN(n1135) );
NAND2_X1 U938 ( .A1(n1233), .A2(n1213), .ZN(n1232) );
XOR2_X1 U939 ( .A(KEYINPUT23), .B(n1234), .Z(n1233) );
NAND2_X1 U940 ( .A1(G116), .A2(n1235), .ZN(n1231) );
XNOR2_X1 U941 ( .A(n1234), .B(KEYINPUT43), .ZN(n1235) );
XOR2_X1 U942 ( .A(G119), .B(n1236), .Z(n1234) );
NOR2_X1 U943 ( .A1(KEYINPUT9), .A2(n1237), .ZN(n1236) );
XNOR2_X1 U944 ( .A(n1238), .B(n1239), .ZN(n1139) );
XNOR2_X1 U945 ( .A(KEYINPUT51), .B(n1240), .ZN(n1229) );
INV_X1 U946 ( .A(n1132), .ZN(n1240) );
XNOR2_X1 U947 ( .A(n1241), .B(G101), .ZN(n1132) );
NAND2_X1 U948 ( .A1(n1242), .A2(G210), .ZN(n1241) );
NOR2_X1 U949 ( .A1(n1212), .A2(n1062), .ZN(n1178) );
XNOR2_X1 U950 ( .A(n1243), .B(G475), .ZN(n1062) );
NAND2_X1 U951 ( .A1(n1228), .A2(n1127), .ZN(n1243) );
NAND2_X1 U952 ( .A1(n1244), .A2(n1245), .ZN(n1127) );
OR2_X1 U953 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XOR2_X1 U954 ( .A(n1248), .B(KEYINPUT13), .Z(n1244) );
NAND2_X1 U955 ( .A1(n1247), .A2(n1246), .ZN(n1248) );
NAND2_X1 U956 ( .A1(n1249), .A2(n1250), .ZN(n1246) );
NAND2_X1 U957 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XOR2_X1 U958 ( .A(n1253), .B(n1254), .Z(n1252) );
XNOR2_X1 U959 ( .A(n1255), .B(n1098), .ZN(n1251) );
XOR2_X1 U960 ( .A(n1256), .B(KEYINPUT37), .Z(n1249) );
NAND2_X1 U961 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XNOR2_X1 U962 ( .A(n1254), .B(n1253), .ZN(n1258) );
NAND2_X1 U963 ( .A1(KEYINPUT45), .A2(G131), .ZN(n1253) );
XOR2_X1 U964 ( .A(n1259), .B(G143), .Z(n1254) );
NAND3_X1 U965 ( .A1(n1242), .A2(G214), .A3(KEYINPUT46), .ZN(n1259) );
NOR2_X1 U966 ( .A1(G953), .A2(G237), .ZN(n1242) );
XOR2_X1 U967 ( .A(n1255), .B(n1098), .Z(n1257) );
XOR2_X1 U968 ( .A(G125), .B(G140), .Z(n1098) );
NAND2_X1 U969 ( .A1(n1260), .A2(KEYINPUT55), .ZN(n1255) );
XOR2_X1 U970 ( .A(n1225), .B(KEYINPUT42), .Z(n1260) );
XNOR2_X1 U971 ( .A(G146), .B(KEYINPUT17), .ZN(n1225) );
XNOR2_X1 U972 ( .A(n1261), .B(n1262), .ZN(n1247) );
NOR2_X1 U973 ( .A1(KEYINPUT38), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U974 ( .A(G113), .B(G122), .ZN(n1261) );
NAND3_X1 U975 ( .A1(n1264), .A2(n1265), .A3(n1057), .ZN(n1212) );
NAND2_X1 U976 ( .A1(G478), .A2(n1266), .ZN(n1057) );
OR2_X1 U977 ( .A1(n1124), .A2(G902), .ZN(n1266) );
NAND2_X1 U978 ( .A1(n1056), .A2(n1267), .ZN(n1265) );
INV_X1 U979 ( .A(KEYINPUT21), .ZN(n1267) );
NOR3_X1 U980 ( .A1(G478), .A2(G902), .A3(n1124), .ZN(n1056) );
XNOR2_X1 U981 ( .A(n1268), .B(n1269), .ZN(n1124) );
XNOR2_X1 U982 ( .A(n1102), .B(n1270), .ZN(n1269) );
NOR2_X1 U983 ( .A1(KEYINPUT18), .A2(n1271), .ZN(n1270) );
XNOR2_X1 U984 ( .A(G128), .B(n1272), .ZN(n1271) );
XOR2_X1 U985 ( .A(KEYINPUT59), .B(G143), .Z(n1272) );
INV_X1 U986 ( .A(G134), .ZN(n1102) );
XOR2_X1 U987 ( .A(n1273), .B(n1274), .Z(n1268) );
AND3_X1 U988 ( .A1(G217), .A2(n1084), .A3(n1223), .ZN(n1274) );
XOR2_X1 U989 ( .A(G234), .B(KEYINPUT22), .Z(n1223) );
NAND2_X1 U990 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
OR2_X1 U991 ( .A1(n1277), .A2(G107), .ZN(n1276) );
XOR2_X1 U992 ( .A(n1278), .B(KEYINPUT60), .Z(n1275) );
NAND2_X1 U993 ( .A1(G107), .A2(n1277), .ZN(n1278) );
XNOR2_X1 U994 ( .A(G116), .B(n1279), .ZN(n1277) );
NAND2_X1 U995 ( .A1(KEYINPUT21), .A2(G478), .ZN(n1264) );
AND3_X1 U996 ( .A1(n1171), .A2(n1170), .A3(n1006), .ZN(n1172) );
INV_X1 U997 ( .A(n1168), .ZN(n1006) );
NAND2_X1 U998 ( .A1(n1034), .A2(n1035), .ZN(n1168) );
NAND2_X1 U999 ( .A1(G214), .A2(n1280), .ZN(n1035) );
XNOR2_X1 U1000 ( .A(n1281), .B(n1067), .ZN(n1034) );
NAND2_X1 U1001 ( .A1(G210), .A2(n1280), .ZN(n1067) );
NAND2_X1 U1002 ( .A1(n1282), .A2(n1228), .ZN(n1280) );
INV_X1 U1003 ( .A(G237), .ZN(n1282) );
NAND2_X1 U1004 ( .A1(KEYINPUT49), .A2(n1065), .ZN(n1281) );
NAND2_X1 U1005 ( .A1(n1283), .A2(n1228), .ZN(n1065) );
XOR2_X1 U1006 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U1007 ( .A(KEYINPUT6), .B(n1190), .ZN(n1285) );
NAND2_X1 U1008 ( .A1(G224), .A2(n1084), .ZN(n1190) );
XNOR2_X1 U1009 ( .A(n1109), .B(n1189), .ZN(n1284) );
XNOR2_X1 U1010 ( .A(G125), .B(n1238), .ZN(n1189) );
XNOR2_X1 U1011 ( .A(n1286), .B(n1287), .ZN(n1238) );
XNOR2_X1 U1012 ( .A(n1288), .B(n1289), .ZN(n1109) );
XOR2_X1 U1013 ( .A(G101), .B(n1290), .Z(n1289) );
XNOR2_X1 U1014 ( .A(n1279), .B(G110), .ZN(n1290) );
INV_X1 U1015 ( .A(G122), .ZN(n1279) );
XOR2_X1 U1016 ( .A(n1291), .B(n1292), .Z(n1288) );
NOR2_X1 U1017 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U1018 ( .A(KEYINPUT47), .B(n1295), .Z(n1294) );
NOR2_X1 U1019 ( .A1(n1237), .A2(n1296), .ZN(n1295) );
AND2_X1 U1020 ( .A1(n1296), .A2(n1237), .ZN(n1293) );
XOR2_X1 U1021 ( .A(G113), .B(KEYINPUT57), .Z(n1237) );
XNOR2_X1 U1022 ( .A(n1213), .B(G119), .ZN(n1296) );
INV_X1 U1023 ( .A(G116), .ZN(n1213) );
NAND3_X1 U1024 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1291) );
NAND2_X1 U1025 ( .A1(KEYINPUT20), .A2(n1300), .ZN(n1299) );
OR3_X1 U1026 ( .A1(n1300), .A2(KEYINPUT20), .A3(G107), .ZN(n1298) );
NAND2_X1 U1027 ( .A1(G107), .A2(n1301), .ZN(n1297) );
NAND2_X1 U1028 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
INV_X1 U1029 ( .A(KEYINPUT20), .ZN(n1303) );
XOR2_X1 U1030 ( .A(KEYINPUT15), .B(n1300), .Z(n1302) );
NAND2_X1 U1031 ( .A1(n1021), .A2(n1304), .ZN(n1170) );
NAND4_X1 U1032 ( .A1(G953), .A2(G902), .A3(n1112), .A4(n1210), .ZN(n1304) );
XOR2_X1 U1033 ( .A(G898), .B(KEYINPUT54), .Z(n1112) );
NAND3_X1 U1034 ( .A1(n1210), .A2(n1084), .A3(G952), .ZN(n1021) );
NAND2_X1 U1035 ( .A1(G237), .A2(G234), .ZN(n1210) );
NOR2_X1 U1036 ( .A1(n1194), .A2(n1028), .ZN(n1171) );
INV_X1 U1037 ( .A(n1042), .ZN(n1028) );
NAND2_X1 U1038 ( .A1(G221), .A2(n1215), .ZN(n1042) );
NAND2_X1 U1039 ( .A1(G234), .A2(n1228), .ZN(n1215) );
INV_X1 U1040 ( .A(n1023), .ZN(n1194) );
XNOR2_X1 U1041 ( .A(n1305), .B(G469), .ZN(n1023) );
NAND2_X1 U1042 ( .A1(n1306), .A2(n1228), .ZN(n1305) );
INV_X1 U1043 ( .A(G902), .ZN(n1228) );
XOR2_X1 U1044 ( .A(n1307), .B(n1152), .Z(n1306) );
XNOR2_X1 U1045 ( .A(n1097), .B(n1239), .ZN(n1152) );
XNOR2_X1 U1046 ( .A(n1308), .B(n1309), .ZN(n1239) );
XNOR2_X1 U1047 ( .A(G137), .B(n1310), .ZN(n1309) );
NAND2_X1 U1048 ( .A1(n1311), .A2(KEYINPUT12), .ZN(n1310) );
XNOR2_X1 U1049 ( .A(G134), .B(KEYINPUT14), .ZN(n1311) );
NAND2_X1 U1050 ( .A1(KEYINPUT53), .A2(n1204), .ZN(n1308) );
INV_X1 U1051 ( .A(G131), .ZN(n1204) );
XOR2_X1 U1052 ( .A(n1312), .B(n1287), .Z(n1097) );
XOR2_X1 U1053 ( .A(G128), .B(KEYINPUT24), .Z(n1287) );
NAND2_X1 U1054 ( .A1(KEYINPUT28), .A2(n1286), .ZN(n1312) );
XOR2_X1 U1055 ( .A(G146), .B(G143), .Z(n1286) );
XOR2_X1 U1056 ( .A(n1145), .B(n1313), .Z(n1307) );
NOR2_X1 U1057 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
INV_X1 U1058 ( .A(n1148), .ZN(n1315) );
NAND2_X1 U1059 ( .A1(n1150), .A2(n1149), .ZN(n1148) );
NOR2_X1 U1060 ( .A1(n1150), .A2(n1149), .ZN(n1314) );
NAND2_X1 U1061 ( .A1(G227), .A2(n1084), .ZN(n1149) );
INV_X1 U1062 ( .A(G953), .ZN(n1084) );
XNOR2_X1 U1063 ( .A(G140), .B(n1316), .ZN(n1150) );
INV_X1 U1064 ( .A(G110), .ZN(n1316) );
XOR2_X1 U1065 ( .A(n1317), .B(G101), .Z(n1145) );
NAND2_X1 U1066 ( .A1(KEYINPUT63), .A2(n1318), .ZN(n1317) );
XOR2_X1 U1067 ( .A(n1319), .B(n1300), .Z(n1318) );
XNOR2_X1 U1068 ( .A(n1263), .B(KEYINPUT5), .ZN(n1300) );
INV_X1 U1069 ( .A(G104), .ZN(n1263) );
NOR2_X1 U1070 ( .A1(G107), .A2(KEYINPUT26), .ZN(n1319) );
endmodule


