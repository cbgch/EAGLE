//Key = 1101010000100000110111111001001100010100100010001100011111111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;

XNOR2_X1 U726 ( .A(G107), .B(n1020), .ZN(G9) );
NOR2_X1 U727 ( .A1(n1021), .A2(n1022), .ZN(G75) );
NOR4_X1 U728 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1022) );
XOR2_X1 U729 ( .A(n1027), .B(KEYINPUT30), .Z(n1026) );
NAND4_X1 U730 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1027) );
XNOR2_X1 U731 ( .A(KEYINPUT2), .B(n1032), .ZN(n1031) );
NOR3_X1 U732 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1025) );
NOR3_X1 U733 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NOR2_X1 U734 ( .A1(n1039), .A2(n1032), .ZN(n1038) );
NOR3_X1 U735 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
NOR3_X1 U736 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
NOR2_X1 U737 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U738 ( .A1(n1048), .A2(n1049), .ZN(n1044) );
NOR3_X1 U739 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1041) );
NOR2_X1 U740 ( .A1(KEYINPUT51), .A2(n1053), .ZN(n1040) );
NOR2_X1 U741 ( .A1(n1054), .A2(n1055), .ZN(n1037) );
INV_X1 U742 ( .A(n1029), .ZN(n1055) );
NOR2_X1 U743 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U744 ( .A1(KEYINPUT6), .A2(n1058), .ZN(n1056) );
NOR2_X1 U745 ( .A1(n1028), .A2(n1059), .ZN(n1034) );
AND3_X1 U746 ( .A1(KEYINPUT6), .A2(n1060), .A3(n1029), .ZN(n1059) );
NAND3_X1 U747 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1023) );
NAND3_X1 U748 ( .A1(n1064), .A2(n1065), .A3(n1028), .ZN(n1063) );
INV_X1 U749 ( .A(n1036), .ZN(n1028) );
NAND2_X1 U750 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND3_X1 U751 ( .A1(n1068), .A2(n1033), .A3(KEYINPUT51), .ZN(n1067) );
NAND2_X1 U752 ( .A1(n1029), .A2(n1069), .ZN(n1066) );
NOR2_X1 U753 ( .A1(n1043), .A2(n1051), .ZN(n1029) );
NOR3_X1 U754 ( .A1(n1070), .A2(G953), .A3(G952), .ZN(n1021) );
INV_X1 U755 ( .A(n1061), .ZN(n1070) );
NAND4_X1 U756 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1061) );
NOR4_X1 U757 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
XOR2_X1 U758 ( .A(n1079), .B(n1080), .Z(n1077) );
NAND2_X1 U759 ( .A1(n1081), .A2(KEYINPUT17), .ZN(n1079) );
XNOR2_X1 U760 ( .A(G475), .B(KEYINPUT33), .ZN(n1081) );
XOR2_X1 U761 ( .A(n1082), .B(n1083), .Z(n1076) );
NAND2_X1 U762 ( .A1(KEYINPUT35), .A2(n1084), .ZN(n1082) );
XNOR2_X1 U763 ( .A(n1085), .B(n1086), .ZN(n1073) );
XNOR2_X1 U764 ( .A(n1052), .B(KEYINPUT45), .ZN(n1071) );
XOR2_X1 U765 ( .A(n1087), .B(n1088), .Z(G72) );
NOR2_X1 U766 ( .A1(n1089), .A2(n1062), .ZN(n1088) );
AND2_X1 U767 ( .A1(G227), .A2(G900), .ZN(n1089) );
NAND2_X1 U768 ( .A1(n1090), .A2(n1091), .ZN(n1087) );
NAND3_X1 U769 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
NAND2_X1 U770 ( .A1(n1095), .A2(G953), .ZN(n1093) );
OR2_X1 U771 ( .A1(n1092), .A2(n1094), .ZN(n1090) );
NAND2_X1 U772 ( .A1(n1062), .A2(n1096), .ZN(n1094) );
NAND3_X1 U773 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
NOR3_X1 U774 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
XOR2_X1 U775 ( .A(n1103), .B(KEYINPUT24), .Z(n1098) );
INV_X1 U776 ( .A(n1104), .ZN(n1097) );
XOR2_X1 U777 ( .A(n1105), .B(n1106), .Z(n1092) );
XNOR2_X1 U778 ( .A(n1107), .B(n1108), .ZN(n1105) );
NAND2_X1 U779 ( .A1(n1109), .A2(n1110), .ZN(G69) );
NAND2_X1 U780 ( .A1(G953), .A2(n1111), .ZN(n1110) );
NAND2_X1 U781 ( .A1(G898), .A2(n1112), .ZN(n1111) );
XNOR2_X1 U782 ( .A(G224), .B(n1113), .ZN(n1112) );
NAND2_X1 U783 ( .A1(n1114), .A2(n1062), .ZN(n1109) );
XOR2_X1 U784 ( .A(n1115), .B(n1113), .Z(n1114) );
XNOR2_X1 U785 ( .A(n1116), .B(KEYINPUT7), .ZN(n1113) );
NAND2_X1 U786 ( .A1(KEYINPUT19), .A2(n1117), .ZN(n1115) );
NOR2_X1 U787 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XOR2_X1 U788 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR3_X1 U789 ( .A1(n1122), .A2(KEYINPUT12), .A3(n1123), .ZN(n1120) );
NOR2_X1 U790 ( .A1(n1118), .A2(n1124), .ZN(G63) );
NOR3_X1 U791 ( .A1(n1083), .A2(n1125), .A3(n1126), .ZN(n1124) );
NOR3_X1 U792 ( .A1(n1127), .A2(n1084), .A3(n1122), .ZN(n1126) );
NOR2_X1 U793 ( .A1(n1128), .A2(n1129), .ZN(n1125) );
NOR2_X1 U794 ( .A1(n1130), .A2(n1084), .ZN(n1128) );
INV_X1 U795 ( .A(G478), .ZN(n1084) );
NOR2_X1 U796 ( .A1(n1118), .A2(n1131), .ZN(G60) );
NOR3_X1 U797 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
NOR2_X1 U798 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
AND3_X1 U799 ( .A1(n1136), .A2(n1135), .A3(n1137), .ZN(n1133) );
INV_X1 U800 ( .A(KEYINPUT50), .ZN(n1136) );
NOR2_X1 U801 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
NOR2_X1 U802 ( .A1(KEYINPUT50), .A2(n1139), .ZN(n1138) );
XOR2_X1 U803 ( .A(KEYINPUT53), .B(n1135), .Z(n1139) );
NOR2_X1 U804 ( .A1(n1122), .A2(n1140), .ZN(n1137) );
XNOR2_X1 U805 ( .A(G104), .B(n1141), .ZN(G6) );
NOR2_X1 U806 ( .A1(n1118), .A2(n1142), .ZN(G57) );
XOR2_X1 U807 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U808 ( .A1(KEYINPUT39), .A2(n1145), .ZN(n1143) );
XOR2_X1 U809 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U810 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U811 ( .A1(n1086), .A2(n1122), .ZN(n1148) );
INV_X1 U812 ( .A(G472), .ZN(n1086) );
NOR2_X1 U813 ( .A1(n1118), .A2(n1150), .ZN(G54) );
XOR2_X1 U814 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U815 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U816 ( .A(n1155), .B(n1156), .Z(n1153) );
XNOR2_X1 U817 ( .A(G110), .B(n1157), .ZN(n1156) );
XNOR2_X1 U818 ( .A(KEYINPUT26), .B(KEYINPUT14), .ZN(n1157) );
XNOR2_X1 U819 ( .A(n1158), .B(n1159), .ZN(n1155) );
XOR2_X1 U820 ( .A(n1160), .B(n1108), .Z(n1159) );
NOR2_X1 U821 ( .A1(n1161), .A2(n1122), .ZN(n1160) );
XNOR2_X1 U822 ( .A(n1162), .B(n1163), .ZN(n1151) );
NAND2_X1 U823 ( .A1(KEYINPUT55), .A2(n1107), .ZN(n1162) );
NOR2_X1 U824 ( .A1(n1118), .A2(n1164), .ZN(G51) );
XOR2_X1 U825 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U826 ( .A(KEYINPUT5), .B(n1167), .Z(n1166) );
NOR2_X1 U827 ( .A1(n1168), .A2(n1122), .ZN(n1167) );
NAND2_X1 U828 ( .A1(G902), .A2(n1024), .ZN(n1122) );
INV_X1 U829 ( .A(n1130), .ZN(n1024) );
NOR4_X1 U830 ( .A1(n1104), .A2(n1103), .A3(n1117), .A4(n1169), .ZN(n1130) );
OR3_X1 U831 ( .A1(n1170), .A2(n1101), .A3(n1102), .ZN(n1169) );
AND4_X1 U832 ( .A1(n1171), .A2(n1060), .A3(n1069), .A4(n1172), .ZN(n1101) );
XNOR2_X1 U833 ( .A(KEYINPUT46), .B(n1043), .ZN(n1172) );
INV_X1 U834 ( .A(n1173), .ZN(n1043) );
XNOR2_X1 U835 ( .A(n1100), .B(KEYINPUT23), .ZN(n1170) );
INV_X1 U836 ( .A(n1174), .ZN(n1100) );
NAND4_X1 U837 ( .A1(n1020), .A2(n1141), .A3(n1175), .A4(n1176), .ZN(n1117) );
NOR4_X1 U838 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
NOR3_X1 U839 ( .A1(n1053), .A2(n1181), .A3(n1182), .ZN(n1180) );
NOR2_X1 U840 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NOR2_X1 U841 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NOR2_X1 U842 ( .A1(n1030), .A2(n1187), .ZN(n1185) );
XOR2_X1 U843 ( .A(KEYINPUT8), .B(n1069), .Z(n1187) );
NOR3_X1 U844 ( .A1(n1033), .A2(n1188), .A3(n1189), .ZN(n1183) );
INV_X1 U845 ( .A(n1068), .ZN(n1053) );
NOR3_X1 U846 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1178) );
INV_X1 U847 ( .A(KEYINPUT43), .ZN(n1190) );
NOR2_X1 U848 ( .A1(KEYINPUT43), .A2(n1193), .ZN(n1177) );
NAND3_X1 U849 ( .A1(n1064), .A2(n1194), .A3(n1069), .ZN(n1141) );
NAND3_X1 U850 ( .A1(n1030), .A2(n1194), .A3(n1064), .ZN(n1020) );
NAND4_X1 U851 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1103) );
NAND2_X1 U852 ( .A1(n1199), .A2(n1200), .ZN(n1104) );
NAND4_X1 U853 ( .A1(n1186), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1200) );
OR2_X1 U854 ( .A1(n1204), .A2(n1203), .ZN(n1199) );
INV_X1 U855 ( .A(KEYINPUT20), .ZN(n1203) );
XNOR2_X1 U856 ( .A(n1116), .B(n1205), .ZN(n1165) );
AND2_X1 U857 ( .A1(n1206), .A2(G953), .ZN(n1118) );
XNOR2_X1 U858 ( .A(G952), .B(KEYINPUT25), .ZN(n1206) );
XNOR2_X1 U859 ( .A(G146), .B(n1174), .ZN(G48) );
NAND3_X1 U860 ( .A1(n1069), .A2(n1207), .A3(n1208), .ZN(n1174) );
XNOR2_X1 U861 ( .A(G143), .B(n1204), .ZN(G45) );
NAND3_X1 U862 ( .A1(n1057), .A2(n1201), .A3(n1202), .ZN(n1204) );
NOR3_X1 U863 ( .A1(n1192), .A2(n1209), .A3(n1210), .ZN(n1202) );
XNOR2_X1 U864 ( .A(G140), .B(n1211), .ZN(G42) );
NAND2_X1 U865 ( .A1(n1212), .A2(n1060), .ZN(n1211) );
NAND3_X1 U866 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(G39) );
NAND2_X1 U867 ( .A1(G137), .A2(n1216), .ZN(n1215) );
NAND2_X1 U868 ( .A1(n1217), .A2(n1218), .ZN(n1214) );
INV_X1 U869 ( .A(KEYINPUT27), .ZN(n1218) );
NAND2_X1 U870 ( .A1(n1102), .A2(n1219), .ZN(n1217) );
XNOR2_X1 U871 ( .A(KEYINPUT49), .B(n1220), .ZN(n1219) );
NAND2_X1 U872 ( .A1(KEYINPUT27), .A2(n1221), .ZN(n1213) );
NAND2_X1 U873 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NAND3_X1 U874 ( .A1(KEYINPUT49), .A2(n1102), .A3(n1220), .ZN(n1223) );
INV_X1 U875 ( .A(n1216), .ZN(n1102) );
NAND3_X1 U876 ( .A1(n1208), .A2(n1173), .A3(n1224), .ZN(n1216) );
OR2_X1 U877 ( .A1(n1220), .A2(KEYINPUT49), .ZN(n1222) );
XOR2_X1 U878 ( .A(n1195), .B(n1225), .Z(G36) );
XNOR2_X1 U879 ( .A(G134), .B(KEYINPUT29), .ZN(n1225) );
NAND4_X1 U880 ( .A1(n1171), .A2(n1173), .A3(n1030), .A4(n1057), .ZN(n1195) );
XNOR2_X1 U881 ( .A(G131), .B(n1196), .ZN(G33) );
NAND2_X1 U882 ( .A1(n1212), .A2(n1057), .ZN(n1196) );
AND3_X1 U883 ( .A1(n1069), .A2(n1173), .A3(n1171), .ZN(n1212) );
INV_X1 U884 ( .A(n1210), .ZN(n1171) );
NOR2_X1 U885 ( .A1(n1052), .A2(n1075), .ZN(n1173) );
INV_X1 U886 ( .A(n1050), .ZN(n1075) );
XOR2_X1 U887 ( .A(n1197), .B(n1226), .Z(G30) );
NAND2_X1 U888 ( .A1(KEYINPUT44), .A2(G128), .ZN(n1226) );
NAND3_X1 U889 ( .A1(n1030), .A2(n1207), .A3(n1208), .ZN(n1197) );
NOR3_X1 U890 ( .A1(n1210), .A2(n1188), .A3(n1189), .ZN(n1208) );
NAND3_X1 U891 ( .A1(n1227), .A2(n1046), .A3(n1049), .ZN(n1210) );
XOR2_X1 U892 ( .A(n1228), .B(n1179), .Z(G3) );
AND3_X1 U893 ( .A1(n1194), .A2(n1057), .A3(n1224), .ZN(n1179) );
AND4_X1 U894 ( .A1(n1049), .A2(n1207), .A3(n1229), .A4(n1046), .ZN(n1194) );
XNOR2_X1 U895 ( .A(G101), .B(KEYINPUT56), .ZN(n1228) );
XNOR2_X1 U896 ( .A(G125), .B(n1198), .ZN(G27) );
NAND4_X1 U897 ( .A1(n1068), .A2(n1060), .A3(n1069), .A4(n1227), .ZN(n1198) );
NAND2_X1 U898 ( .A1(n1230), .A2(n1036), .ZN(n1227) );
NAND4_X1 U899 ( .A1(n1231), .A2(n1095), .A3(G902), .A4(n1232), .ZN(n1230) );
XNOR2_X1 U900 ( .A(G900), .B(KEYINPUT34), .ZN(n1095) );
XNOR2_X1 U901 ( .A(G953), .B(KEYINPUT48), .ZN(n1231) );
XNOR2_X1 U902 ( .A(G122), .B(n1175), .ZN(G24) );
NAND3_X1 U903 ( .A1(n1068), .A2(n1064), .A3(n1233), .ZN(n1175) );
NOR3_X1 U904 ( .A1(n1234), .A2(n1181), .A3(n1209), .ZN(n1233) );
XNOR2_X1 U905 ( .A(G119), .B(n1235), .ZN(G21) );
NAND3_X1 U906 ( .A1(n1068), .A2(n1224), .A3(n1236), .ZN(n1235) );
NOR3_X1 U907 ( .A1(n1189), .A2(n1188), .A3(n1237), .ZN(n1236) );
XNOR2_X1 U908 ( .A(n1181), .B(KEYINPUT21), .ZN(n1237) );
XNOR2_X1 U909 ( .A(G116), .B(n1238), .ZN(G18) );
NAND4_X1 U910 ( .A1(n1239), .A2(n1068), .A3(n1030), .A4(n1229), .ZN(n1238) );
NOR2_X1 U911 ( .A1(n1201), .A2(n1209), .ZN(n1030) );
XOR2_X1 U912 ( .A(n1240), .B(KEYINPUT4), .Z(n1209) );
NOR2_X1 U913 ( .A1(n1051), .A2(n1192), .ZN(n1068) );
XNOR2_X1 U914 ( .A(KEYINPUT10), .B(n1057), .ZN(n1239) );
XNOR2_X1 U915 ( .A(G113), .B(n1241), .ZN(G15) );
NAND4_X1 U916 ( .A1(n1069), .A2(n1072), .A3(n1242), .A4(n1243), .ZN(n1241) );
XNOR2_X1 U917 ( .A(KEYINPUT9), .B(n1192), .ZN(n1243) );
NOR2_X1 U918 ( .A1(n1181), .A2(n1186), .ZN(n1242) );
INV_X1 U919 ( .A(n1057), .ZN(n1186) );
NAND2_X1 U920 ( .A1(n1244), .A2(n1245), .ZN(n1057) );
OR3_X1 U921 ( .A1(n1078), .A2(n1189), .A3(KEYINPUT62), .ZN(n1245) );
NAND2_X1 U922 ( .A1(KEYINPUT62), .A2(n1064), .ZN(n1244) );
INV_X1 U923 ( .A(n1032), .ZN(n1064) );
NAND2_X1 U924 ( .A1(n1188), .A2(n1189), .ZN(n1032) );
INV_X1 U925 ( .A(n1078), .ZN(n1188) );
INV_X1 U926 ( .A(n1051), .ZN(n1072) );
NAND2_X1 U927 ( .A1(n1047), .A2(n1046), .ZN(n1051) );
AND2_X1 U928 ( .A1(n1240), .A2(n1201), .ZN(n1069) );
INV_X1 U929 ( .A(n1234), .ZN(n1201) );
XNOR2_X1 U930 ( .A(G110), .B(n1246), .ZN(G12) );
NOR2_X1 U931 ( .A1(n1247), .A2(KEYINPUT52), .ZN(n1246) );
INV_X1 U932 ( .A(n1193), .ZN(n1247) );
NAND2_X1 U933 ( .A1(n1191), .A2(n1207), .ZN(n1193) );
INV_X1 U934 ( .A(n1192), .ZN(n1207) );
NAND2_X1 U935 ( .A1(n1248), .A2(n1050), .ZN(n1192) );
NAND2_X1 U936 ( .A1(G214), .A2(n1249), .ZN(n1050) );
XNOR2_X1 U937 ( .A(n1052), .B(KEYINPUT63), .ZN(n1248) );
XOR2_X1 U938 ( .A(n1250), .B(n1168), .Z(n1052) );
NAND2_X1 U939 ( .A1(G210), .A2(n1249), .ZN(n1168) );
NAND2_X1 U940 ( .A1(n1251), .A2(n1252), .ZN(n1249) );
INV_X1 U941 ( .A(G237), .ZN(n1251) );
NAND2_X1 U942 ( .A1(n1253), .A2(n1252), .ZN(n1250) );
XNOR2_X1 U943 ( .A(n1254), .B(n1255), .ZN(n1253) );
INV_X1 U944 ( .A(n1116), .ZN(n1255) );
XNOR2_X1 U945 ( .A(n1256), .B(n1257), .ZN(n1116) );
XNOR2_X1 U946 ( .A(G110), .B(n1258), .ZN(n1257) );
XNOR2_X1 U947 ( .A(KEYINPUT3), .B(KEYINPUT13), .ZN(n1258) );
XOR2_X1 U948 ( .A(n1259), .B(n1260), .Z(n1256) );
XOR2_X1 U949 ( .A(n1261), .B(n1262), .Z(n1259) );
NOR2_X1 U950 ( .A1(KEYINPUT42), .A2(n1205), .ZN(n1254) );
XNOR2_X1 U951 ( .A(n1263), .B(n1264), .ZN(n1205) );
XNOR2_X1 U952 ( .A(G125), .B(n1265), .ZN(n1263) );
AND2_X1 U953 ( .A1(n1062), .A2(G224), .ZN(n1265) );
AND4_X1 U954 ( .A1(n1224), .A2(n1060), .A3(n1266), .A4(n1049), .ZN(n1191) );
XOR2_X1 U955 ( .A(n1047), .B(KEYINPUT0), .Z(n1049) );
XNOR2_X1 U956 ( .A(n1267), .B(n1161), .ZN(n1047) );
INV_X1 U957 ( .A(G469), .ZN(n1161) );
NAND2_X1 U958 ( .A1(n1268), .A2(n1252), .ZN(n1267) );
XOR2_X1 U959 ( .A(n1269), .B(n1270), .Z(n1268) );
NOR2_X1 U960 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XOR2_X1 U961 ( .A(n1273), .B(KEYINPUT16), .Z(n1272) );
NAND2_X1 U962 ( .A1(n1274), .A2(n1163), .ZN(n1273) );
NOR2_X1 U963 ( .A1(n1274), .A2(n1163), .ZN(n1271) );
NAND2_X1 U964 ( .A1(G227), .A2(n1062), .ZN(n1163) );
XOR2_X1 U965 ( .A(n1154), .B(n1275), .Z(n1274) );
NOR2_X1 U966 ( .A1(KEYINPUT38), .A2(n1276), .ZN(n1275) );
INV_X1 U967 ( .A(G110), .ZN(n1276) );
XOR2_X1 U968 ( .A(G140), .B(KEYINPUT41), .Z(n1154) );
NAND2_X1 U969 ( .A1(n1277), .A2(n1278), .ZN(n1269) );
NAND2_X1 U970 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
XNOR2_X1 U971 ( .A(KEYINPUT31), .B(n1281), .ZN(n1280) );
INV_X1 U972 ( .A(n1107), .ZN(n1281) );
XOR2_X1 U973 ( .A(n1282), .B(n1283), .Z(n1279) );
XOR2_X1 U974 ( .A(n1284), .B(KEYINPUT36), .Z(n1277) );
NAND2_X1 U975 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
XNOR2_X1 U976 ( .A(n1282), .B(n1283), .ZN(n1286) );
XOR2_X1 U977 ( .A(n1108), .B(KEYINPUT61), .Z(n1283) );
XOR2_X1 U978 ( .A(n1287), .B(n1288), .Z(n1108) );
XNOR2_X1 U979 ( .A(G128), .B(KEYINPUT28), .ZN(n1287) );
NAND2_X1 U980 ( .A1(KEYINPUT1), .A2(n1158), .ZN(n1282) );
XOR2_X1 U981 ( .A(n1262), .B(KEYINPUT58), .Z(n1158) );
XOR2_X1 U982 ( .A(G101), .B(n1289), .Z(n1262) );
XOR2_X1 U983 ( .A(G107), .B(G104), .Z(n1289) );
XNOR2_X1 U984 ( .A(n1107), .B(KEYINPUT31), .ZN(n1285) );
NOR2_X1 U985 ( .A1(n1048), .A2(n1181), .ZN(n1266) );
INV_X1 U986 ( .A(n1229), .ZN(n1181) );
NAND2_X1 U987 ( .A1(n1036), .A2(n1290), .ZN(n1229) );
NAND4_X1 U988 ( .A1(G953), .A2(G902), .A3(n1232), .A4(n1291), .ZN(n1290) );
INV_X1 U989 ( .A(G898), .ZN(n1291) );
NAND3_X1 U990 ( .A1(n1232), .A2(n1062), .A3(G952), .ZN(n1036) );
NAND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1232) );
INV_X1 U992 ( .A(n1046), .ZN(n1048) );
NAND2_X1 U993 ( .A1(G221), .A2(n1292), .ZN(n1046) );
NAND2_X1 U994 ( .A1(G234), .A2(n1252), .ZN(n1292) );
INV_X1 U995 ( .A(n1058), .ZN(n1060) );
NAND2_X1 U996 ( .A1(n1189), .A2(n1078), .ZN(n1058) );
NAND3_X1 U997 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(n1078) );
NAND2_X1 U998 ( .A1(n1296), .A2(n1121), .ZN(n1295) );
OR3_X1 U999 ( .A1(n1121), .A2(n1296), .A3(G902), .ZN(n1294) );
NOR2_X1 U1000 ( .A1(n1123), .A2(G234), .ZN(n1296) );
INV_X1 U1001 ( .A(G217), .ZN(n1123) );
XNOR2_X1 U1002 ( .A(n1297), .B(n1298), .ZN(n1121) );
XOR2_X1 U1003 ( .A(n1299), .B(n1300), .Z(n1298) );
XNOR2_X1 U1004 ( .A(n1301), .B(G110), .ZN(n1300) );
INV_X1 U1005 ( .A(G119), .ZN(n1301) );
XNOR2_X1 U1006 ( .A(KEYINPUT22), .B(n1302), .ZN(n1299) );
XNOR2_X1 U1007 ( .A(n1303), .B(n1304), .ZN(n1297) );
XOR2_X1 U1008 ( .A(n1305), .B(n1306), .Z(n1304) );
NAND2_X1 U1009 ( .A1(KEYINPUT57), .A2(n1307), .ZN(n1306) );
INV_X1 U1010 ( .A(G146), .ZN(n1307) );
NAND2_X1 U1011 ( .A1(n1308), .A2(n1309), .ZN(n1305) );
NAND4_X1 U1012 ( .A1(G234), .A2(G221), .A3(G137), .A4(n1062), .ZN(n1309) );
NAND2_X1 U1013 ( .A1(n1310), .A2(n1311), .ZN(n1308) );
NAND3_X1 U1014 ( .A1(G221), .A2(n1062), .A3(G234), .ZN(n1311) );
XNOR2_X1 U1015 ( .A(G137), .B(KEYINPUT32), .ZN(n1310) );
NAND2_X1 U1016 ( .A1(G902), .A2(G217), .ZN(n1293) );
XNOR2_X1 U1017 ( .A(n1312), .B(G472), .ZN(n1189) );
NAND2_X1 U1018 ( .A1(KEYINPUT54), .A2(n1085), .ZN(n1312) );
NAND2_X1 U1019 ( .A1(n1313), .A2(n1252), .ZN(n1085) );
INV_X1 U1020 ( .A(G902), .ZN(n1252) );
XNOR2_X1 U1021 ( .A(n1144), .B(n1314), .ZN(n1313) );
XNOR2_X1 U1022 ( .A(n1315), .B(KEYINPUT59), .ZN(n1314) );
NAND2_X1 U1023 ( .A1(KEYINPUT37), .A2(n1316), .ZN(n1315) );
XNOR2_X1 U1024 ( .A(n1317), .B(n1149), .ZN(n1316) );
XOR2_X1 U1025 ( .A(n1107), .B(n1264), .Z(n1149) );
XNOR2_X1 U1026 ( .A(n1288), .B(n1318), .ZN(n1264) );
NOR2_X1 U1027 ( .A1(KEYINPUT15), .A2(n1302), .ZN(n1318) );
XOR2_X1 U1028 ( .A(G131), .B(n1319), .Z(n1107) );
XNOR2_X1 U1029 ( .A(n1220), .B(G134), .ZN(n1319) );
INV_X1 U1030 ( .A(G137), .ZN(n1220) );
NAND2_X1 U1031 ( .A1(KEYINPUT60), .A2(n1146), .ZN(n1317) );
XNOR2_X1 U1032 ( .A(n1261), .B(n1320), .ZN(n1146) );
XNOR2_X1 U1033 ( .A(G119), .B(n1321), .ZN(n1261) );
XOR2_X1 U1034 ( .A(n1322), .B(n1323), .Z(n1144) );
INV_X1 U1035 ( .A(G101), .ZN(n1323) );
NAND2_X1 U1036 ( .A1(G210), .A2(n1324), .ZN(n1322) );
INV_X1 U1037 ( .A(n1033), .ZN(n1224) );
NAND2_X1 U1038 ( .A1(n1234), .A2(n1240), .ZN(n1033) );
XNOR2_X1 U1039 ( .A(n1083), .B(G478), .ZN(n1240) );
NOR2_X1 U1040 ( .A1(n1129), .A2(G902), .ZN(n1083) );
INV_X1 U1041 ( .A(n1127), .ZN(n1129) );
XNOR2_X1 U1042 ( .A(n1325), .B(n1326), .ZN(n1127) );
XNOR2_X1 U1043 ( .A(n1302), .B(n1327), .ZN(n1326) );
XOR2_X1 U1044 ( .A(G143), .B(G134), .Z(n1327) );
INV_X1 U1045 ( .A(G128), .ZN(n1302) );
XOR2_X1 U1046 ( .A(n1328), .B(n1329), .Z(n1325) );
AND3_X1 U1047 ( .A1(G234), .A2(n1062), .A3(G217), .ZN(n1329) );
INV_X1 U1048 ( .A(G953), .ZN(n1062) );
NAND2_X1 U1049 ( .A1(n1330), .A2(n1331), .ZN(n1328) );
NAND2_X1 U1050 ( .A1(G107), .A2(n1260), .ZN(n1331) );
XOR2_X1 U1051 ( .A(n1332), .B(KEYINPUT11), .Z(n1330) );
OR2_X1 U1052 ( .A1(n1260), .A2(G107), .ZN(n1332) );
XOR2_X1 U1053 ( .A(G122), .B(n1320), .Z(n1260) );
XOR2_X1 U1054 ( .A(G116), .B(KEYINPUT18), .Z(n1320) );
XOR2_X1 U1055 ( .A(n1080), .B(n1140), .Z(n1234) );
INV_X1 U1056 ( .A(G475), .ZN(n1140) );
NOR2_X1 U1057 ( .A1(n1135), .A2(G902), .ZN(n1080) );
XNOR2_X1 U1058 ( .A(n1333), .B(n1334), .ZN(n1135) );
XNOR2_X1 U1059 ( .A(n1335), .B(n1336), .ZN(n1334) );
XNOR2_X1 U1060 ( .A(n1288), .B(n1321), .ZN(n1336) );
XOR2_X1 U1061 ( .A(G113), .B(KEYINPUT47), .Z(n1321) );
XNOR2_X1 U1062 ( .A(G143), .B(G146), .ZN(n1288) );
INV_X1 U1063 ( .A(n1303), .ZN(n1335) );
XOR2_X1 U1064 ( .A(n1106), .B(KEYINPUT40), .Z(n1303) );
XOR2_X1 U1065 ( .A(G125), .B(G140), .Z(n1106) );
XOR2_X1 U1066 ( .A(n1337), .B(n1338), .Z(n1333) );
XOR2_X1 U1067 ( .A(G131), .B(G122), .Z(n1338) );
XOR2_X1 U1068 ( .A(n1339), .B(G104), .Z(n1337) );
NAND2_X1 U1069 ( .A1(G214), .A2(n1324), .ZN(n1339) );
NOR2_X1 U1070 ( .A1(G953), .A2(G237), .ZN(n1324) );
endmodule


