//Key = 0011111101111110000101011110011000000111001101110110001001001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355;

XNOR2_X1 U738 ( .A(G107), .B(n1021), .ZN(G9) );
NOR2_X1 U739 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR4_X1 U740 ( .A1(n1024), .A2(n1025), .A3(G953), .A4(n1026), .ZN(n1023) );
NOR3_X1 U741 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1025) );
NOR2_X1 U742 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR2_X1 U743 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U744 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U745 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR2_X1 U746 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U747 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR3_X1 U748 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1034) );
NOR3_X1 U749 ( .A1(n1037), .A2(n1045), .A3(n1043), .ZN(n1030) );
NAND3_X1 U750 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1024) );
NAND2_X1 U751 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NAND2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U754 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND3_X1 U755 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
NAND2_X1 U756 ( .A1(n1060), .A2(n1061), .ZN(n1055) );
NAND2_X1 U757 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND3_X1 U758 ( .A1(n1058), .A2(n1064), .A3(KEYINPUT37), .ZN(n1063) );
NAND2_X1 U759 ( .A1(n1057), .A2(n1065), .ZN(n1062) );
OR2_X1 U760 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(n1051) );
INV_X1 U762 ( .A(KEYINPUT37), .ZN(n1069) );
NAND4_X1 U763 ( .A1(n1053), .A2(n1060), .A3(n1058), .A4(n1064), .ZN(n1068) );
INV_X1 U764 ( .A(n1027), .ZN(n1053) );
NOR3_X1 U765 ( .A1(n1026), .A2(G953), .A3(G952), .ZN(n1022) );
AND4_X1 U766 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1026) );
NOR4_X1 U767 ( .A1(n1074), .A2(n1075), .A3(n1043), .A4(n1076), .ZN(n1073) );
XOR2_X1 U768 ( .A(n1077), .B(n1078), .Z(n1076) );
NOR2_X1 U769 ( .A1(KEYINPUT40), .A2(n1079), .ZN(n1078) );
XOR2_X1 U770 ( .A(n1080), .B(KEYINPUT11), .Z(n1075) );
XNOR2_X1 U771 ( .A(n1081), .B(KEYINPUT26), .ZN(n1074) );
NOR3_X1 U772 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1072) );
INV_X1 U773 ( .A(n1085), .ZN(n1084) );
AND2_X1 U774 ( .A1(n1079), .A2(KEYINPUT40), .ZN(n1082) );
XOR2_X1 U775 ( .A(n1086), .B(n1087), .Z(n1071) );
NAND2_X1 U776 ( .A1(KEYINPUT54), .A2(n1088), .ZN(n1087) );
INV_X1 U777 ( .A(G478), .ZN(n1088) );
XNOR2_X1 U778 ( .A(n1089), .B(n1090), .ZN(n1070) );
NAND2_X1 U779 ( .A1(KEYINPUT9), .A2(n1091), .ZN(n1090) );
XOR2_X1 U780 ( .A(n1092), .B(n1093), .Z(G72) );
XOR2_X1 U781 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND3_X1 U782 ( .A1(n1096), .A2(n1097), .A3(KEYINPUT4), .ZN(n1095) );
NAND2_X1 U783 ( .A1(G900), .A2(G227), .ZN(n1097) );
INV_X1 U784 ( .A(n1098), .ZN(n1096) );
NAND2_X1 U785 ( .A1(n1099), .A2(n1100), .ZN(n1094) );
INV_X1 U786 ( .A(n1101), .ZN(n1100) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(n1099) );
XOR2_X1 U788 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U789 ( .A1(KEYINPUT50), .A2(n1106), .ZN(n1105) );
NOR2_X1 U790 ( .A1(n1107), .A2(G953), .ZN(n1092) );
NOR3_X1 U791 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1107) );
XOR2_X1 U792 ( .A(n1111), .B(KEYINPUT61), .Z(n1110) );
XOR2_X1 U793 ( .A(n1112), .B(n1113), .Z(G69) );
XOR2_X1 U794 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U795 ( .A1(n1116), .A2(n1098), .ZN(n1115) );
XOR2_X1 U796 ( .A(n1117), .B(KEYINPUT56), .Z(n1098) );
NOR2_X1 U797 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NAND2_X1 U798 ( .A1(n1120), .A2(n1121), .ZN(n1114) );
NAND2_X1 U799 ( .A1(G953), .A2(n1119), .ZN(n1121) );
XNOR2_X1 U800 ( .A(n1122), .B(n1123), .ZN(n1120) );
NAND2_X1 U801 ( .A1(n1124), .A2(n1117), .ZN(n1112) );
XOR2_X1 U802 ( .A(KEYINPUT43), .B(n1048), .Z(n1124) );
NOR2_X1 U803 ( .A1(n1125), .A2(n1126), .ZN(G66) );
NOR3_X1 U804 ( .A1(n1089), .A2(n1127), .A3(n1128), .ZN(n1126) );
NOR3_X1 U805 ( .A1(n1129), .A2(n1091), .A3(n1130), .ZN(n1128) );
INV_X1 U806 ( .A(n1131), .ZN(n1129) );
NOR2_X1 U807 ( .A1(n1132), .A2(n1131), .ZN(n1127) );
NOR2_X1 U808 ( .A1(n1133), .A2(n1091), .ZN(n1132) );
NOR3_X1 U809 ( .A1(n1125), .A2(n1134), .A3(n1135), .ZN(G63) );
NOR2_X1 U810 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NOR2_X1 U811 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
AND2_X1 U812 ( .A1(n1140), .A2(KEYINPUT53), .ZN(n1139) );
NOR3_X1 U813 ( .A1(KEYINPUT53), .A2(n1140), .A3(n1141), .ZN(n1138) );
INV_X1 U814 ( .A(n1142), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1143), .A2(n1142), .ZN(n1134) );
XNOR2_X1 U816 ( .A(n1144), .B(KEYINPUT25), .ZN(n1142) );
NOR2_X1 U817 ( .A1(n1140), .A2(n1141), .ZN(n1143) );
INV_X1 U818 ( .A(KEYINPUT38), .ZN(n1141) );
NAND2_X1 U819 ( .A1(n1145), .A2(G478), .ZN(n1140) );
NOR2_X1 U820 ( .A1(n1125), .A2(n1146), .ZN(G60) );
XOR2_X1 U821 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U822 ( .A1(KEYINPUT27), .A2(n1149), .ZN(n1148) );
NAND2_X1 U823 ( .A1(n1145), .A2(G475), .ZN(n1147) );
XOR2_X1 U824 ( .A(n1150), .B(n1151), .Z(G6) );
NOR2_X1 U825 ( .A1(n1125), .A2(n1152), .ZN(G57) );
XOR2_X1 U826 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U827 ( .A(n1155), .B(n1156), .Z(n1154) );
AND2_X1 U828 ( .A1(G472), .A2(n1145), .ZN(n1155) );
XNOR2_X1 U829 ( .A(n1157), .B(n1158), .ZN(n1153) );
NOR2_X1 U830 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U831 ( .A(KEYINPUT36), .B(n1161), .Z(n1160) );
NOR2_X1 U832 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
AND2_X1 U833 ( .A1(n1163), .A2(n1162), .ZN(n1159) );
NOR2_X1 U834 ( .A1(n1125), .A2(n1164), .ZN(G54) );
XOR2_X1 U835 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U836 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U837 ( .A1(n1169), .A2(n1130), .ZN(n1167) );
INV_X1 U838 ( .A(n1145), .ZN(n1130) );
XOR2_X1 U839 ( .A(n1170), .B(KEYINPUT62), .Z(n1165) );
NAND2_X1 U840 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
INV_X1 U841 ( .A(n1173), .ZN(n1171) );
NOR2_X1 U842 ( .A1(n1125), .A2(n1174), .ZN(G51) );
XOR2_X1 U843 ( .A(n1175), .B(n1176), .Z(n1174) );
AND2_X1 U844 ( .A1(G210), .A2(n1145), .ZN(n1176) );
NOR2_X1 U845 ( .A1(n1177), .A2(n1133), .ZN(n1145) );
AND2_X1 U846 ( .A1(n1048), .A2(n1178), .ZN(n1133) );
XOR2_X1 U847 ( .A(KEYINPUT58), .B(n1046), .Z(n1178) );
AND3_X1 U848 ( .A1(n1179), .A2(n1111), .A3(n1180), .ZN(n1046) );
INV_X1 U849 ( .A(n1108), .ZN(n1180) );
NAND4_X1 U850 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1108) );
AND3_X1 U851 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
NAND2_X1 U852 ( .A1(n1039), .A2(n1188), .ZN(n1183) );
NAND2_X1 U853 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U854 ( .A1(n1191), .A2(n1059), .ZN(n1190) );
XOR2_X1 U855 ( .A(KEYINPUT5), .B(n1192), .Z(n1189) );
OR4_X1 U856 ( .A1(n1043), .A2(n1064), .A3(n1193), .A4(KEYINPUT21), .ZN(n1182) );
NAND2_X1 U857 ( .A1(n1194), .A2(KEYINPUT21), .ZN(n1181) );
XOR2_X1 U858 ( .A(KEYINPUT47), .B(n1109), .Z(n1179) );
INV_X1 U859 ( .A(n1195), .ZN(n1109) );
AND4_X1 U860 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1048) );
AND4_X1 U861 ( .A1(n1200), .A2(n1021), .A3(n1201), .A4(n1202), .ZN(n1199) );
NAND3_X1 U862 ( .A1(n1203), .A2(n1204), .A3(n1058), .ZN(n1021) );
NOR3_X1 U863 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1198) );
NOR2_X1 U864 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NOR4_X1 U865 ( .A1(n1039), .A2(n1210), .A3(n1029), .A4(n1211), .ZN(n1206) );
INV_X1 U866 ( .A(n1058), .ZN(n1029) );
NAND3_X1 U867 ( .A1(n1212), .A2(n1213), .A3(n1064), .ZN(n1210) );
NOR2_X1 U868 ( .A1(n1151), .A2(n1213), .ZN(n1205) );
INV_X1 U869 ( .A(KEYINPUT57), .ZN(n1213) );
NAND3_X1 U870 ( .A1(n1058), .A2(n1204), .A3(n1059), .ZN(n1151) );
NAND3_X1 U871 ( .A1(n1214), .A2(n1203), .A3(n1067), .ZN(n1196) );
NAND3_X1 U872 ( .A1(n1215), .A2(n1216), .A3(KEYINPUT12), .ZN(n1175) );
NAND2_X1 U873 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
INV_X1 U874 ( .A(KEYINPUT35), .ZN(n1218) );
XOR2_X1 U875 ( .A(n1219), .B(n1220), .Z(n1217) );
NAND2_X1 U876 ( .A1(KEYINPUT35), .A2(n1221), .ZN(n1215) );
NAND2_X1 U877 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NAND3_X1 U878 ( .A1(KEYINPUT51), .A2(n1224), .A3(n1225), .ZN(n1223) );
INV_X1 U879 ( .A(n1226), .ZN(n1224) );
NAND2_X1 U880 ( .A1(n1219), .A2(n1220), .ZN(n1222) );
INV_X1 U881 ( .A(n1225), .ZN(n1220) );
NOR2_X1 U882 ( .A1(n1226), .A2(KEYINPUT51), .ZN(n1219) );
XOR2_X1 U883 ( .A(n1227), .B(KEYINPUT3), .Z(n1226) );
NOR2_X1 U884 ( .A1(n1117), .A2(G952), .ZN(n1125) );
NAND3_X1 U885 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(G48) );
NAND4_X1 U886 ( .A1(n1191), .A2(n1059), .A3(n1039), .A4(n1231), .ZN(n1230) );
NAND2_X1 U887 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NAND2_X1 U888 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND3_X1 U889 ( .A1(G146), .A2(n1236), .A3(n1232), .ZN(n1229) );
INV_X1 U890 ( .A(KEYINPUT33), .ZN(n1232) );
NAND4_X1 U891 ( .A1(n1191), .A2(n1059), .A3(n1039), .A4(n1235), .ZN(n1236) );
INV_X1 U892 ( .A(KEYINPUT17), .ZN(n1235) );
NAND2_X1 U893 ( .A1(KEYINPUT33), .A2(n1234), .ZN(n1228) );
INV_X1 U894 ( .A(G146), .ZN(n1234) );
XOR2_X1 U895 ( .A(n1237), .B(n1185), .Z(G45) );
NAND4_X1 U896 ( .A1(n1238), .A2(n1239), .A3(n1039), .A4(n1240), .ZN(n1185) );
XOR2_X1 U897 ( .A(G140), .B(n1194), .Z(G42) );
NOR3_X1 U898 ( .A1(n1043), .A2(n1241), .A3(n1193), .ZN(n1194) );
XOR2_X1 U899 ( .A(G137), .B(n1242), .Z(G39) );
NOR2_X1 U900 ( .A1(KEYINPUT15), .A2(n1195), .ZN(n1242) );
NAND3_X1 U901 ( .A1(n1060), .A2(n1049), .A3(n1191), .ZN(n1195) );
XOR2_X1 U902 ( .A(n1243), .B(G134), .Z(G36) );
NAND2_X1 U903 ( .A1(KEYINPUT24), .A2(n1187), .ZN(n1243) );
NAND3_X1 U904 ( .A1(n1049), .A2(n1203), .A3(n1239), .ZN(n1187) );
XOR2_X1 U905 ( .A(n1186), .B(n1244), .Z(G33) );
NAND2_X1 U906 ( .A1(KEYINPUT49), .A2(G131), .ZN(n1244) );
NAND3_X1 U907 ( .A1(n1059), .A2(n1049), .A3(n1239), .ZN(n1186) );
AND3_X1 U908 ( .A1(n1064), .A2(n1245), .A3(n1067), .ZN(n1239) );
INV_X1 U909 ( .A(n1043), .ZN(n1049) );
NAND2_X1 U910 ( .A1(n1246), .A2(n1041), .ZN(n1043) );
INV_X1 U911 ( .A(n1040), .ZN(n1246) );
XOR2_X1 U912 ( .A(n1247), .B(n1111), .Z(G30) );
NAND3_X1 U913 ( .A1(n1203), .A2(n1039), .A3(n1191), .ZN(n1111) );
AND4_X1 U914 ( .A1(n1064), .A2(n1081), .A3(n1248), .A4(n1245), .ZN(n1191) );
INV_X1 U915 ( .A(n1045), .ZN(n1203) );
XOR2_X1 U916 ( .A(G101), .B(n1249), .Z(G3) );
NOR2_X1 U917 ( .A1(n1208), .A2(n1250), .ZN(n1249) );
XNOR2_X1 U918 ( .A(KEYINPUT19), .B(n1209), .ZN(n1250) );
NAND4_X1 U919 ( .A1(n1067), .A2(n1060), .A3(n1064), .A4(n1212), .ZN(n1209) );
XOR2_X1 U920 ( .A(n1251), .B(n1252), .Z(G27) );
NAND2_X1 U921 ( .A1(n1192), .A2(n1039), .ZN(n1252) );
NOR2_X1 U922 ( .A1(n1193), .A2(n1037), .ZN(n1192) );
INV_X1 U923 ( .A(n1057), .ZN(n1037) );
NAND3_X1 U924 ( .A1(n1066), .A2(n1245), .A3(n1059), .ZN(n1193) );
NAND2_X1 U925 ( .A1(n1027), .A2(n1253), .ZN(n1245) );
NAND3_X1 U926 ( .A1(G902), .A2(n1254), .A3(n1101), .ZN(n1253) );
NOR2_X1 U927 ( .A1(n1117), .A2(G900), .ZN(n1101) );
XOR2_X1 U928 ( .A(n1200), .B(n1255), .Z(G24) );
XOR2_X1 U929 ( .A(n1256), .B(KEYINPUT31), .Z(n1255) );
NAND4_X1 U930 ( .A1(n1238), .A2(n1214), .A3(n1058), .A4(n1240), .ZN(n1200) );
NAND2_X1 U931 ( .A1(n1257), .A2(n1258), .ZN(G21) );
NAND2_X1 U932 ( .A1(G119), .A2(n1197), .ZN(n1258) );
XOR2_X1 U933 ( .A(KEYINPUT29), .B(n1259), .Z(n1257) );
NOR2_X1 U934 ( .A1(G119), .A2(n1197), .ZN(n1259) );
NAND4_X1 U935 ( .A1(n1060), .A2(n1214), .A3(n1081), .A4(n1248), .ZN(n1197) );
XOR2_X1 U936 ( .A(n1260), .B(n1261), .Z(G18) );
XNOR2_X1 U937 ( .A(G116), .B(KEYINPUT41), .ZN(n1261) );
NAND4_X1 U938 ( .A1(n1262), .A2(n1067), .A3(n1263), .A4(n1057), .ZN(n1260) );
NOR2_X1 U939 ( .A1(n1208), .A2(n1045), .ZN(n1263) );
NAND2_X1 U940 ( .A1(n1240), .A2(n1264), .ZN(n1045) );
INV_X1 U941 ( .A(n1265), .ZN(n1240) );
XOR2_X1 U942 ( .A(n1212), .B(KEYINPUT59), .Z(n1262) );
XOR2_X1 U943 ( .A(n1266), .B(n1202), .Z(G15) );
NAND3_X1 U944 ( .A1(n1067), .A2(n1214), .A3(n1059), .ZN(n1202) );
INV_X1 U945 ( .A(n1211), .ZN(n1059) );
NAND2_X1 U946 ( .A1(n1265), .A2(n1238), .ZN(n1211) );
AND3_X1 U947 ( .A1(n1039), .A2(n1212), .A3(n1057), .ZN(n1214) );
NOR2_X1 U948 ( .A1(n1044), .A2(n1083), .ZN(n1057) );
INV_X1 U949 ( .A(n1042), .ZN(n1083) );
AND2_X1 U950 ( .A1(n1267), .A2(n1081), .ZN(n1067) );
XOR2_X1 U951 ( .A(KEYINPUT2), .B(n1248), .Z(n1267) );
XNOR2_X1 U952 ( .A(G110), .B(n1201), .ZN(G12) );
NAND3_X1 U953 ( .A1(n1204), .A2(n1066), .A3(n1060), .ZN(n1201) );
INV_X1 U954 ( .A(n1033), .ZN(n1060) );
NAND2_X1 U955 ( .A1(n1265), .A2(n1264), .ZN(n1033) );
INV_X1 U956 ( .A(n1238), .ZN(n1264) );
XOR2_X1 U957 ( .A(n1268), .B(n1077), .Z(n1238) );
NOR2_X1 U958 ( .A1(n1149), .A2(G902), .ZN(n1077) );
XNOR2_X1 U959 ( .A(n1269), .B(n1270), .ZN(n1149) );
XOR2_X1 U960 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR4_X1 U961 ( .A1(n1273), .A2(n1274), .A3(KEYINPUT32), .A4(n1275), .ZN(n1272) );
NOR2_X1 U962 ( .A1(G104), .A2(n1276), .ZN(n1275) );
NOR2_X1 U963 ( .A1(KEYINPUT22), .A2(n1277), .ZN(n1276) );
AND2_X1 U964 ( .A1(KEYINPUT52), .A2(n1277), .ZN(n1274) );
NOR4_X1 U965 ( .A1(KEYINPUT52), .A2(n1150), .A3(KEYINPUT22), .A4(n1277), .ZN(n1273) );
XOR2_X1 U966 ( .A(n1266), .B(n1256), .Z(n1277) );
INV_X1 U967 ( .A(G122), .ZN(n1256) );
NOR3_X1 U968 ( .A1(n1278), .A2(G953), .A3(G237), .ZN(n1271) );
XNOR2_X1 U969 ( .A(G214), .B(KEYINPUT0), .ZN(n1278) );
XNOR2_X1 U970 ( .A(n1102), .B(n1279), .ZN(n1269) );
XOR2_X1 U971 ( .A(G131), .B(n1280), .Z(n1102) );
NAND2_X1 U972 ( .A1(KEYINPUT45), .A2(n1079), .ZN(n1268) );
INV_X1 U973 ( .A(G475), .ZN(n1079) );
XOR2_X1 U974 ( .A(n1086), .B(G478), .Z(n1265) );
NAND2_X1 U975 ( .A1(n1144), .A2(n1177), .ZN(n1086) );
XNOR2_X1 U976 ( .A(n1281), .B(n1282), .ZN(n1144) );
XOR2_X1 U977 ( .A(G116), .B(n1283), .Z(n1282) );
XOR2_X1 U978 ( .A(G134), .B(G122), .Z(n1283) );
XOR2_X1 U979 ( .A(n1284), .B(n1285), .Z(n1281) );
XOR2_X1 U980 ( .A(G107), .B(n1286), .Z(n1285) );
AND3_X1 U981 ( .A1(G217), .A2(n1117), .A3(G234), .ZN(n1286) );
NAND2_X1 U982 ( .A1(KEYINPUT30), .A2(n1287), .ZN(n1284) );
XOR2_X1 U983 ( .A(G143), .B(G128), .Z(n1287) );
NAND2_X1 U984 ( .A1(n1288), .A2(n1289), .ZN(n1066) );
OR3_X1 U985 ( .A1(n1290), .A2(n1081), .A3(KEYINPUT48), .ZN(n1289) );
NAND2_X1 U986 ( .A1(KEYINPUT48), .A2(n1058), .ZN(n1288) );
NOR2_X1 U987 ( .A1(n1248), .A2(n1081), .ZN(n1058) );
XNOR2_X1 U988 ( .A(n1291), .B(G472), .ZN(n1081) );
NAND2_X1 U989 ( .A1(n1292), .A2(n1177), .ZN(n1291) );
XOR2_X1 U990 ( .A(n1293), .B(n1294), .Z(n1292) );
XNOR2_X1 U991 ( .A(KEYINPUT63), .B(n1162), .ZN(n1294) );
NAND3_X1 U992 ( .A1(n1295), .A2(n1117), .A3(G210), .ZN(n1162) );
XOR2_X1 U993 ( .A(KEYINPUT7), .B(G237), .Z(n1295) );
XNOR2_X1 U994 ( .A(n1156), .B(n1296), .ZN(n1293) );
XNOR2_X1 U995 ( .A(n1297), .B(n1298), .ZN(n1156) );
XOR2_X1 U996 ( .A(n1299), .B(G113), .Z(n1297) );
INV_X1 U997 ( .A(n1290), .ZN(n1248) );
XOR2_X1 U998 ( .A(n1089), .B(n1091), .Z(n1290) );
NAND2_X1 U999 ( .A1(G217), .A2(n1300), .ZN(n1091) );
NOR2_X1 U1000 ( .A1(n1131), .A2(G902), .ZN(n1089) );
XOR2_X1 U1001 ( .A(n1301), .B(n1302), .Z(n1131) );
XOR2_X1 U1002 ( .A(G137), .B(n1303), .Z(n1302) );
AND3_X1 U1003 ( .A1(G234), .A2(n1117), .A3(G221), .ZN(n1303) );
NAND2_X1 U1004 ( .A1(KEYINPUT13), .A2(n1304), .ZN(n1301) );
XOR2_X1 U1005 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1006 ( .A(n1280), .B(n1307), .ZN(n1306) );
XNOR2_X1 U1007 ( .A(n1251), .B(G140), .ZN(n1280) );
INV_X1 U1008 ( .A(G125), .ZN(n1251) );
XNOR2_X1 U1009 ( .A(G110), .B(n1308), .ZN(n1305) );
XOR2_X1 U1010 ( .A(G146), .B(G128), .Z(n1308) );
AND3_X1 U1011 ( .A1(n1039), .A2(n1212), .A3(n1064), .ZN(n1204) );
INV_X1 U1012 ( .A(n1241), .ZN(n1064) );
NAND2_X1 U1013 ( .A1(n1042), .A2(n1044), .ZN(n1241) );
NAND2_X1 U1014 ( .A1(n1085), .A2(n1080), .ZN(n1044) );
NAND2_X1 U1015 ( .A1(G469), .A2(n1309), .ZN(n1080) );
NAND2_X1 U1016 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NAND3_X1 U1017 ( .A1(n1311), .A2(n1169), .A3(n1310), .ZN(n1085) );
XOR2_X1 U1018 ( .A(KEYINPUT20), .B(n1177), .Z(n1310) );
INV_X1 U1019 ( .A(G469), .ZN(n1169) );
XNOR2_X1 U1020 ( .A(n1168), .B(n1312), .ZN(n1311) );
XOR2_X1 U1021 ( .A(KEYINPUT16), .B(n1313), .Z(n1312) );
NOR2_X1 U1022 ( .A1(n1173), .A2(n1314), .ZN(n1313) );
XNOR2_X1 U1023 ( .A(KEYINPUT18), .B(n1172), .ZN(n1314) );
NAND3_X1 U1024 ( .A1(G227), .A2(n1117), .A3(n1315), .ZN(n1172) );
NOR2_X1 U1025 ( .A1(n1315), .A2(n1316), .ZN(n1173) );
AND2_X1 U1026 ( .A1(G227), .A2(n1117), .ZN(n1316) );
XNOR2_X1 U1027 ( .A(G140), .B(G110), .ZN(n1315) );
XNOR2_X1 U1028 ( .A(n1317), .B(n1318), .ZN(n1168) );
XOR2_X1 U1029 ( .A(G104), .B(n1319), .Z(n1318) );
XOR2_X1 U1030 ( .A(KEYINPUT34), .B(G107), .Z(n1319) );
XOR2_X1 U1031 ( .A(n1296), .B(n1104), .Z(n1317) );
NAND2_X1 U1032 ( .A1(n1320), .A2(n1321), .ZN(n1104) );
NAND2_X1 U1033 ( .A1(n1322), .A2(n1247), .ZN(n1321) );
XOR2_X1 U1034 ( .A(n1323), .B(KEYINPUT44), .Z(n1320) );
OR2_X1 U1035 ( .A1(n1322), .A2(n1247), .ZN(n1323) );
XNOR2_X1 U1036 ( .A(n1324), .B(G146), .ZN(n1322) );
NAND2_X1 U1037 ( .A1(KEYINPUT39), .A2(n1237), .ZN(n1324) );
INV_X1 U1038 ( .A(G143), .ZN(n1237) );
XOR2_X1 U1039 ( .A(n1157), .B(n1163), .Z(n1296) );
NAND2_X1 U1040 ( .A1(n1325), .A2(n1326), .ZN(n1157) );
NAND2_X1 U1041 ( .A1(G131), .A2(n1327), .ZN(n1326) );
XOR2_X1 U1042 ( .A(KEYINPUT14), .B(n1328), .Z(n1325) );
NOR2_X1 U1043 ( .A1(G131), .A2(n1327), .ZN(n1328) );
INV_X1 U1044 ( .A(n1106), .ZN(n1327) );
XOR2_X1 U1045 ( .A(n1329), .B(G137), .Z(n1106) );
INV_X1 U1046 ( .A(G134), .ZN(n1329) );
NAND2_X1 U1047 ( .A1(G221), .A2(n1300), .ZN(n1042) );
NAND2_X1 U1048 ( .A1(G234), .A2(n1330), .ZN(n1300) );
XOR2_X1 U1049 ( .A(KEYINPUT42), .B(G902), .Z(n1330) );
NAND2_X1 U1050 ( .A1(n1027), .A2(n1331), .ZN(n1212) );
NAND4_X1 U1051 ( .A1(G953), .A2(G902), .A3(n1254), .A4(n1119), .ZN(n1331) );
INV_X1 U1052 ( .A(G898), .ZN(n1119) );
NAND3_X1 U1053 ( .A1(n1254), .A2(n1117), .A3(G952), .ZN(n1027) );
INV_X1 U1054 ( .A(G953), .ZN(n1117) );
NAND2_X1 U1055 ( .A1(G237), .A2(G234), .ZN(n1254) );
INV_X1 U1056 ( .A(n1208), .ZN(n1039) );
NAND2_X1 U1057 ( .A1(n1040), .A2(n1041), .ZN(n1208) );
NAND2_X1 U1058 ( .A1(G214), .A2(n1332), .ZN(n1041) );
NAND2_X1 U1059 ( .A1(n1333), .A2(n1177), .ZN(n1332) );
NAND2_X1 U1060 ( .A1(n1334), .A2(n1335), .ZN(n1040) );
NAND2_X1 U1061 ( .A1(G210), .A2(n1336), .ZN(n1335) );
NAND2_X1 U1062 ( .A1(n1177), .A2(n1337), .ZN(n1336) );
OR2_X1 U1063 ( .A1(n1338), .A2(n1333), .ZN(n1337) );
INV_X1 U1064 ( .A(G237), .ZN(n1333) );
NAND3_X1 U1065 ( .A1(n1339), .A2(n1177), .A3(n1338), .ZN(n1334) );
XOR2_X1 U1066 ( .A(n1225), .B(n1227), .Z(n1338) );
XOR2_X1 U1067 ( .A(n1340), .B(n1123), .Z(n1227) );
XNOR2_X1 U1068 ( .A(n1341), .B(n1342), .ZN(n1123) );
XNOR2_X1 U1069 ( .A(G110), .B(n1343), .ZN(n1342) );
NAND2_X1 U1070 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
OR2_X1 U1071 ( .A1(n1346), .A2(n1163), .ZN(n1345) );
XOR2_X1 U1072 ( .A(n1347), .B(KEYINPUT55), .Z(n1344) );
NAND2_X1 U1073 ( .A1(n1346), .A2(n1163), .ZN(n1347) );
INV_X1 U1074 ( .A(G101), .ZN(n1163) );
XNOR2_X1 U1075 ( .A(n1150), .B(n1348), .ZN(n1346) );
NOR2_X1 U1076 ( .A1(G107), .A2(KEYINPUT8), .ZN(n1348) );
INV_X1 U1077 ( .A(G104), .ZN(n1150) );
XOR2_X1 U1078 ( .A(n1349), .B(G122), .Z(n1341) );
XNOR2_X1 U1079 ( .A(KEYINPUT10), .B(KEYINPUT1), .ZN(n1349) );
XOR2_X1 U1080 ( .A(n1350), .B(KEYINPUT23), .Z(n1340) );
NAND2_X1 U1081 ( .A1(KEYINPUT6), .A2(n1122), .ZN(n1350) );
XNOR2_X1 U1082 ( .A(n1351), .B(n1352), .ZN(n1122) );
INV_X1 U1083 ( .A(n1299), .ZN(n1352) );
XNOR2_X1 U1084 ( .A(G116), .B(n1307), .ZN(n1299) );
XOR2_X1 U1085 ( .A(G119), .B(KEYINPUT28), .Z(n1307) );
NAND2_X1 U1086 ( .A1(KEYINPUT60), .A2(n1266), .ZN(n1351) );
INV_X1 U1087 ( .A(G113), .ZN(n1266) );
XNOR2_X1 U1088 ( .A(n1298), .B(n1353), .ZN(n1225) );
XOR2_X1 U1089 ( .A(G125), .B(n1354), .Z(n1353) );
NOR2_X1 U1090 ( .A1(G953), .A2(n1118), .ZN(n1354) );
INV_X1 U1091 ( .A(G224), .ZN(n1118) );
XNOR2_X1 U1092 ( .A(n1355), .B(n1279), .ZN(n1298) );
XOR2_X1 U1093 ( .A(G143), .B(G146), .Z(n1279) );
NAND2_X1 U1094 ( .A1(KEYINPUT46), .A2(n1247), .ZN(n1355) );
INV_X1 U1095 ( .A(G128), .ZN(n1247) );
INV_X1 U1096 ( .A(G902), .ZN(n1177) );
NAND2_X1 U1097 ( .A1(G210), .A2(G237), .ZN(n1339) );
endmodule


