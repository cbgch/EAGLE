//Key = 1110001100100010011101001110011111010010011110100010001001110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;

XOR2_X1 U760 ( .A(G107), .B(n1051), .Z(G9) );
NAND3_X1 U761 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(G75) );
NAND2_X1 U762 ( .A1(G952), .A2(n1055), .ZN(n1054) );
NAND3_X1 U763 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NAND4_X1 U764 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1057) );
NAND2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NAND2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U767 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
OR2_X1 U768 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U769 ( .A1(n1071), .A2(n1072), .ZN(n1063) );
NAND2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1056) );
NAND2_X1 U771 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND3_X1 U772 ( .A1(n1076), .A2(n1062), .A3(n1065), .ZN(n1075) );
NAND2_X1 U773 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U774 ( .A1(n1060), .A2(n1079), .ZN(n1078) );
NAND2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U776 ( .A1(n1059), .A2(n1082), .ZN(n1077) );
NAND2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U779 ( .A(n1087), .B(KEYINPUT28), .Z(n1074) );
NAND4_X1 U780 ( .A1(n1059), .A2(n1060), .A3(n1088), .A4(n1062), .ZN(n1087) );
NAND3_X1 U781 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1052) );
NOR4_X1 U782 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1091) );
NOR3_X1 U783 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
INV_X1 U784 ( .A(KEYINPUT0), .ZN(n1096) );
NOR2_X1 U785 ( .A1(KEYINPUT0), .A2(G478), .ZN(n1094) );
NAND3_X1 U786 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1092) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U788 ( .A1(KEYINPUT3), .A2(n1104), .ZN(n1103) );
XNOR2_X1 U789 ( .A(G472), .B(KEYINPUT19), .ZN(n1104) );
NAND2_X1 U790 ( .A1(n1105), .A2(n1106), .ZN(n1100) );
XNOR2_X1 U791 ( .A(n1107), .B(n1108), .ZN(n1099) );
XNOR2_X1 U792 ( .A(KEYINPUT17), .B(KEYINPUT12), .ZN(n1108) );
NOR3_X1 U793 ( .A1(n1109), .A2(n1110), .A3(n1085), .ZN(n1090) );
INV_X1 U794 ( .A(n1111), .ZN(n1110) );
AND3_X1 U795 ( .A1(n1112), .A2(n1069), .A3(n1113), .ZN(n1089) );
XOR2_X1 U796 ( .A(n1114), .B(n1115), .Z(G72) );
NAND2_X1 U797 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
OR3_X1 U798 ( .A1(n1053), .A2(G227), .A3(n1118), .ZN(n1117) );
NAND2_X1 U799 ( .A1(n1119), .A2(n1118), .ZN(n1116) );
OR2_X1 U800 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
XNOR2_X1 U801 ( .A(n1122), .B(n1123), .ZN(n1120) );
NOR3_X1 U802 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
AND2_X1 U803 ( .A1(G125), .A2(KEYINPUT8), .ZN(n1126) );
NOR2_X1 U804 ( .A1(KEYINPUT8), .A2(n1127), .ZN(n1125) );
NOR2_X1 U805 ( .A1(KEYINPUT20), .A2(n1128), .ZN(n1122) );
XOR2_X1 U806 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U807 ( .A1(KEYINPUT32), .A2(n1131), .ZN(n1129) );
NAND2_X1 U808 ( .A1(G953), .A2(n1132), .ZN(n1119) );
NAND2_X1 U809 ( .A1(G900), .A2(G227), .ZN(n1132) );
NAND2_X1 U810 ( .A1(n1053), .A2(n1133), .ZN(n1114) );
XOR2_X1 U811 ( .A(n1134), .B(n1135), .Z(G69) );
XOR2_X1 U812 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND3_X1 U813 ( .A1(n1138), .A2(n1053), .A3(KEYINPUT58), .ZN(n1137) );
NAND2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
NAND2_X1 U815 ( .A1(G953), .A2(n1141), .ZN(n1140) );
XNOR2_X1 U816 ( .A(n1142), .B(n1143), .ZN(n1139) );
XOR2_X1 U817 ( .A(n1144), .B(KEYINPUT6), .Z(n1143) );
NOR3_X1 U818 ( .A1(n1053), .A2(KEYINPUT5), .A3(n1145), .ZN(n1134) );
AND2_X1 U819 ( .A1(G224), .A2(G898), .ZN(n1145) );
NOR2_X1 U820 ( .A1(n1146), .A2(n1147), .ZN(G66) );
XOR2_X1 U821 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U822 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
AND2_X1 U823 ( .A1(KEYINPUT60), .A2(n1152), .ZN(n1151) );
NOR2_X1 U824 ( .A1(KEYINPUT51), .A2(n1152), .ZN(n1150) );
NAND2_X1 U825 ( .A1(n1153), .A2(n1105), .ZN(n1152) );
NOR2_X1 U826 ( .A1(n1146), .A2(n1154), .ZN(G63) );
XOR2_X1 U827 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U828 ( .A1(n1098), .A2(n1157), .ZN(n1156) );
NOR2_X1 U829 ( .A1(n1146), .A2(n1158), .ZN(G60) );
XOR2_X1 U830 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND3_X1 U831 ( .A1(n1161), .A2(n1162), .A3(G475), .ZN(n1159) );
NAND2_X1 U832 ( .A1(KEYINPUT35), .A2(n1157), .ZN(n1162) );
NAND2_X1 U833 ( .A1(n1163), .A2(n1164), .ZN(n1161) );
INV_X1 U834 ( .A(KEYINPUT35), .ZN(n1164) );
NAND2_X1 U835 ( .A1(n1058), .A2(G902), .ZN(n1163) );
XNOR2_X1 U836 ( .A(G104), .B(n1165), .ZN(G6) );
NOR2_X1 U837 ( .A1(n1146), .A2(n1166), .ZN(G57) );
XNOR2_X1 U838 ( .A(n1167), .B(n1168), .ZN(n1166) );
NAND2_X1 U839 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
NAND2_X1 U840 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XOR2_X1 U841 ( .A(n1173), .B(n1174), .Z(n1169) );
AND2_X1 U842 ( .A1(G472), .A2(n1153), .ZN(n1174) );
OR2_X1 U843 ( .A1(n1172), .A2(n1171), .ZN(n1173) );
NAND3_X1 U844 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1171) );
NAND2_X1 U845 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND3_X1 U846 ( .A1(n1180), .A2(n1181), .A3(KEYINPUT41), .ZN(n1176) );
INV_X1 U847 ( .A(n1179), .ZN(n1180) );
NAND2_X1 U848 ( .A1(n1182), .A2(n1183), .ZN(n1179) );
XOR2_X1 U849 ( .A(KEYINPUT37), .B(KEYINPUT25), .Z(n1182) );
OR2_X1 U850 ( .A1(n1183), .A2(KEYINPUT41), .ZN(n1175) );
INV_X1 U851 ( .A(KEYINPUT14), .ZN(n1172) );
NOR2_X1 U852 ( .A1(n1146), .A2(n1184), .ZN(G54) );
XOR2_X1 U853 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U854 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U855 ( .A(G110), .B(n1189), .Z(n1188) );
NOR2_X1 U856 ( .A1(KEYINPUT53), .A2(n1190), .ZN(n1189) );
AND2_X1 U857 ( .A1(G469), .A2(n1153), .ZN(n1187) );
XNOR2_X1 U858 ( .A(n1191), .B(n1192), .ZN(n1185) );
XNOR2_X1 U859 ( .A(n1193), .B(n1131), .ZN(n1192) );
NAND2_X1 U860 ( .A1(KEYINPUT43), .A2(n1194), .ZN(n1193) );
NOR2_X1 U861 ( .A1(n1146), .A2(n1195), .ZN(G51) );
XOR2_X1 U862 ( .A(n1196), .B(n1197), .Z(n1195) );
NOR2_X1 U863 ( .A1(n1198), .A2(n1157), .ZN(n1197) );
INV_X1 U864 ( .A(n1153), .ZN(n1157) );
NOR2_X1 U865 ( .A1(n1199), .A2(n1058), .ZN(n1153) );
NOR2_X1 U866 ( .A1(n1133), .A2(n1138), .ZN(n1058) );
NAND4_X1 U867 ( .A1(n1165), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1138) );
NOR4_X1 U868 ( .A1(n1051), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1202) );
INV_X1 U869 ( .A(n1206), .ZN(n1205) );
AND3_X1 U870 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1051) );
NAND2_X1 U871 ( .A1(n1210), .A2(n1211), .ZN(n1201) );
NAND2_X1 U872 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XOR2_X1 U873 ( .A(KEYINPUT29), .B(n1214), .Z(n1213) );
XOR2_X1 U874 ( .A(KEYINPUT24), .B(n1215), .Z(n1212) );
NAND3_X1 U875 ( .A1(n1209), .A2(n1208), .A3(n1216), .ZN(n1165) );
NAND4_X1 U876 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1133) );
NOR4_X1 U877 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1220) );
NAND2_X1 U878 ( .A1(n1225), .A2(n1226), .ZN(n1219) );
NAND2_X1 U879 ( .A1(n1227), .A2(n1081), .ZN(n1226) );
XNOR2_X1 U880 ( .A(KEYINPUT30), .B(n1080), .ZN(n1227) );
INV_X1 U881 ( .A(n1228), .ZN(n1225) );
NOR2_X1 U882 ( .A1(KEYINPUT36), .A2(n1229), .ZN(n1196) );
XOR2_X1 U883 ( .A(n1230), .B(n1231), .Z(n1229) );
XNOR2_X1 U884 ( .A(n1232), .B(n1233), .ZN(n1231) );
XNOR2_X1 U885 ( .A(KEYINPUT38), .B(n1234), .ZN(n1233) );
XNOR2_X1 U886 ( .A(n1235), .B(n1236), .ZN(n1230) );
AND2_X1 U887 ( .A1(G953), .A2(n1237), .ZN(n1146) );
XOR2_X1 U888 ( .A(KEYINPUT46), .B(G952), .Z(n1237) );
XOR2_X1 U889 ( .A(n1238), .B(n1239), .Z(G48) );
NOR2_X1 U890 ( .A1(KEYINPUT39), .A2(n1240), .ZN(n1239) );
NOR2_X1 U891 ( .A1(n1080), .A2(n1228), .ZN(n1238) );
XOR2_X1 U892 ( .A(G143), .B(n1223), .Z(G45) );
AND4_X1 U893 ( .A1(n1241), .A2(n1242), .A3(n1093), .A4(n1243), .ZN(n1223) );
AND3_X1 U894 ( .A1(n1088), .A2(n1210), .A3(n1209), .ZN(n1243) );
NAND2_X1 U895 ( .A1(n1244), .A2(n1245), .ZN(G42) );
NAND2_X1 U896 ( .A1(n1224), .A2(n1194), .ZN(n1245) );
INV_X1 U897 ( .A(n1246), .ZN(n1224) );
XOR2_X1 U898 ( .A(n1247), .B(KEYINPUT49), .Z(n1244) );
NAND2_X1 U899 ( .A1(G140), .A2(n1246), .ZN(n1247) );
NAND3_X1 U900 ( .A1(n1216), .A2(n1248), .A3(n1071), .ZN(n1246) );
XNOR2_X1 U901 ( .A(n1217), .B(n1249), .ZN(G39) );
XOR2_X1 U902 ( .A(KEYINPUT27), .B(G137), .Z(n1249) );
NAND2_X1 U903 ( .A1(n1250), .A2(n1248), .ZN(n1217) );
XNOR2_X1 U904 ( .A(n1251), .B(n1222), .ZN(G36) );
AND3_X1 U905 ( .A1(n1248), .A2(n1207), .A3(n1088), .ZN(n1222) );
XOR2_X1 U906 ( .A(G131), .B(n1221), .Z(G33) );
AND3_X1 U907 ( .A1(n1088), .A2(n1248), .A3(n1216), .ZN(n1221) );
AND3_X1 U908 ( .A1(n1209), .A2(n1241), .A3(n1072), .ZN(n1248) );
NOR2_X1 U909 ( .A1(n1070), .A2(n1252), .ZN(n1072) );
INV_X1 U910 ( .A(n1069), .ZN(n1252) );
XNOR2_X1 U911 ( .A(G128), .B(n1253), .ZN(G30) );
NOR2_X1 U912 ( .A1(n1254), .A2(KEYINPUT23), .ZN(n1253) );
NOR2_X1 U913 ( .A1(n1081), .A2(n1228), .ZN(n1254) );
NAND4_X1 U914 ( .A1(n1241), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1228) );
NOR2_X1 U915 ( .A1(n1067), .A2(n1083), .ZN(n1257) );
INV_X1 U916 ( .A(n1209), .ZN(n1083) );
INV_X1 U917 ( .A(n1207), .ZN(n1081) );
XOR2_X1 U918 ( .A(n1200), .B(n1258), .Z(G3) );
XNOR2_X1 U919 ( .A(KEYINPUT44), .B(n1259), .ZN(n1258) );
NAND4_X1 U920 ( .A1(n1059), .A2(n1088), .A3(n1209), .A4(n1260), .ZN(n1200) );
XNOR2_X1 U921 ( .A(G125), .B(n1218), .ZN(G27) );
NAND4_X1 U922 ( .A1(n1060), .A2(n1071), .A3(n1261), .A4(n1216), .ZN(n1218) );
AND2_X1 U923 ( .A1(n1241), .A2(n1210), .ZN(n1261) );
NAND2_X1 U924 ( .A1(n1262), .A2(n1263), .ZN(n1241) );
NAND3_X1 U925 ( .A1(G902), .A2(n1062), .A3(n1121), .ZN(n1263) );
NOR2_X1 U926 ( .A1(n1053), .A2(G900), .ZN(n1121) );
XNOR2_X1 U927 ( .A(G122), .B(n1206), .ZN(G24) );
NAND4_X1 U928 ( .A1(n1060), .A2(n1208), .A3(n1093), .A4(n1242), .ZN(n1206) );
AND2_X1 U929 ( .A1(n1065), .A2(n1260), .ZN(n1208) );
NOR2_X1 U930 ( .A1(n1255), .A2(n1256), .ZN(n1065) );
XOR2_X1 U931 ( .A(G119), .B(n1204), .Z(G21) );
AND3_X1 U932 ( .A1(n1060), .A2(n1260), .A3(n1250), .ZN(n1204) );
AND3_X1 U933 ( .A1(n1256), .A2(n1255), .A3(n1059), .ZN(n1250) );
XNOR2_X1 U934 ( .A(G116), .B(n1264), .ZN(G18) );
NOR2_X1 U935 ( .A1(n1203), .A2(KEYINPUT16), .ZN(n1264) );
AND4_X1 U936 ( .A1(n1060), .A2(n1088), .A3(n1207), .A4(n1260), .ZN(n1203) );
AND2_X1 U937 ( .A1(n1210), .A2(n1265), .ZN(n1260) );
NOR2_X1 U938 ( .A1(n1093), .A2(n1266), .ZN(n1207) );
NAND3_X1 U939 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(G15) );
NAND3_X1 U940 ( .A1(n1210), .A2(n1270), .A3(n1214), .ZN(n1269) );
NAND2_X1 U941 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND2_X1 U942 ( .A1(KEYINPUT50), .A2(n1273), .ZN(n1272) );
NAND3_X1 U943 ( .A1(G113), .A2(n1274), .A3(n1271), .ZN(n1268) );
INV_X1 U944 ( .A(KEYINPUT56), .ZN(n1271) );
NAND3_X1 U945 ( .A1(n1214), .A2(n1210), .A3(KEYINPUT50), .ZN(n1274) );
AND4_X1 U946 ( .A1(n1060), .A2(n1216), .A3(n1088), .A4(n1265), .ZN(n1214) );
NOR2_X1 U947 ( .A1(n1255), .A2(n1275), .ZN(n1088) );
INV_X1 U948 ( .A(n1256), .ZN(n1275) );
INV_X1 U949 ( .A(n1080), .ZN(n1216) );
NAND2_X1 U950 ( .A1(n1266), .A2(n1093), .ZN(n1080) );
INV_X1 U951 ( .A(n1242), .ZN(n1266) );
NOR2_X1 U952 ( .A1(n1107), .A2(n1085), .ZN(n1060) );
NAND2_X1 U953 ( .A1(KEYINPUT56), .A2(n1273), .ZN(n1267) );
XOR2_X1 U954 ( .A(n1276), .B(n1277), .Z(G12) );
NOR2_X1 U955 ( .A1(G110), .A2(KEYINPUT13), .ZN(n1277) );
NAND2_X1 U956 ( .A1(n1215), .A2(n1210), .ZN(n1276) );
INV_X1 U957 ( .A(n1067), .ZN(n1210) );
NAND2_X1 U958 ( .A1(n1070), .A2(n1069), .ZN(n1067) );
NAND2_X1 U959 ( .A1(G214), .A2(n1278), .ZN(n1069) );
NAND2_X1 U960 ( .A1(n1279), .A2(n1112), .ZN(n1070) );
NAND2_X1 U961 ( .A1(n1280), .A2(n1198), .ZN(n1112) );
XOR2_X1 U962 ( .A(KEYINPUT59), .B(n1109), .Z(n1279) );
NOR2_X1 U963 ( .A1(n1198), .A2(n1280), .ZN(n1109) );
AND2_X1 U964 ( .A1(n1281), .A2(n1199), .ZN(n1280) );
XOR2_X1 U965 ( .A(n1282), .B(KEYINPUT7), .Z(n1281) );
NAND2_X1 U966 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NAND2_X1 U967 ( .A1(n1235), .A2(n1285), .ZN(n1284) );
XOR2_X1 U968 ( .A(n1286), .B(KEYINPUT40), .Z(n1283) );
OR2_X1 U969 ( .A1(n1285), .A2(n1235), .ZN(n1286) );
XNOR2_X1 U970 ( .A(n1144), .B(n1287), .ZN(n1235) );
NOR2_X1 U971 ( .A1(KEYINPUT52), .A2(n1288), .ZN(n1287) );
XOR2_X1 U972 ( .A(n1289), .B(n1290), .Z(n1144) );
XNOR2_X1 U973 ( .A(KEYINPUT45), .B(n1291), .ZN(n1290) );
XNOR2_X1 U974 ( .A(n1183), .B(G110), .ZN(n1289) );
NAND3_X1 U975 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n1285) );
NAND2_X1 U976 ( .A1(n1232), .A2(n1295), .ZN(n1294) );
NAND2_X1 U977 ( .A1(n1296), .A2(n1297), .ZN(n1293) );
INV_X1 U978 ( .A(KEYINPUT33), .ZN(n1297) );
NAND2_X1 U979 ( .A1(n1298), .A2(n1299), .ZN(n1296) );
INV_X1 U980 ( .A(n1232), .ZN(n1299) );
XNOR2_X1 U981 ( .A(n1295), .B(n1300), .ZN(n1298) );
NAND2_X1 U982 ( .A1(KEYINPUT33), .A2(n1301), .ZN(n1292) );
NAND2_X1 U983 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NAND2_X1 U984 ( .A1(n1295), .A2(n1300), .ZN(n1303) );
OR3_X1 U985 ( .A1(n1295), .A2(n1232), .A3(n1300), .ZN(n1302) );
INV_X1 U986 ( .A(KEYINPUT31), .ZN(n1300) );
NAND2_X1 U987 ( .A1(G224), .A2(n1053), .ZN(n1232) );
NAND2_X1 U988 ( .A1(n1304), .A2(n1305), .ZN(n1295) );
NAND2_X1 U989 ( .A1(n1306), .A2(G125), .ZN(n1305) );
XOR2_X1 U990 ( .A(n1307), .B(KEYINPUT11), .Z(n1304) );
NAND2_X1 U991 ( .A1(n1236), .A2(n1234), .ZN(n1307) );
NAND2_X1 U992 ( .A1(G210), .A2(n1278), .ZN(n1198) );
NAND2_X1 U993 ( .A1(n1199), .A2(n1308), .ZN(n1278) );
INV_X1 U994 ( .A(G237), .ZN(n1308) );
AND4_X1 U995 ( .A1(n1059), .A2(n1071), .A3(n1209), .A4(n1265), .ZN(n1215) );
NAND2_X1 U996 ( .A1(n1262), .A2(n1309), .ZN(n1265) );
NAND4_X1 U997 ( .A1(G953), .A2(G902), .A3(n1062), .A4(n1141), .ZN(n1309) );
INV_X1 U998 ( .A(G898), .ZN(n1141) );
NAND3_X1 U999 ( .A1(G952), .A2(n1053), .A3(n1310), .ZN(n1262) );
XOR2_X1 U1000 ( .A(n1062), .B(KEYINPUT15), .Z(n1310) );
NAND2_X1 U1001 ( .A1(G237), .A2(G234), .ZN(n1062) );
NOR2_X1 U1002 ( .A1(n1086), .A2(n1085), .ZN(n1209) );
AND2_X1 U1003 ( .A1(G221), .A2(n1311), .ZN(n1085) );
INV_X1 U1004 ( .A(n1107), .ZN(n1086) );
XNOR2_X1 U1005 ( .A(n1312), .B(G469), .ZN(n1107) );
NAND2_X1 U1006 ( .A1(n1313), .A2(n1199), .ZN(n1312) );
XOR2_X1 U1007 ( .A(n1314), .B(n1315), .Z(n1313) );
XNOR2_X1 U1008 ( .A(n1316), .B(n1317), .ZN(n1315) );
INV_X1 U1009 ( .A(n1131), .ZN(n1317) );
NAND2_X1 U1010 ( .A1(KEYINPUT1), .A2(n1318), .ZN(n1316) );
INV_X1 U1011 ( .A(n1190), .ZN(n1318) );
NAND2_X1 U1012 ( .A1(G227), .A2(n1053), .ZN(n1190) );
XOR2_X1 U1013 ( .A(n1319), .B(n1320), .Z(n1314) );
NOR2_X1 U1014 ( .A1(KEYINPUT34), .A2(n1191), .ZN(n1320) );
XNOR2_X1 U1015 ( .A(n1130), .B(n1288), .ZN(n1191) );
INV_X1 U1016 ( .A(n1142), .ZN(n1288) );
XOR2_X1 U1017 ( .A(G101), .B(n1321), .Z(n1142) );
XOR2_X1 U1018 ( .A(G107), .B(G104), .Z(n1321) );
XOR2_X1 U1019 ( .A(G128), .B(n1322), .Z(n1130) );
XNOR2_X1 U1020 ( .A(G110), .B(G140), .ZN(n1319) );
AND2_X1 U1021 ( .A1(n1323), .A2(n1255), .ZN(n1071) );
NAND3_X1 U1022 ( .A1(n1324), .A2(n1325), .A3(n1113), .ZN(n1255) );
OR2_X1 U1023 ( .A1(n1106), .A2(n1105), .ZN(n1113) );
NAND3_X1 U1024 ( .A1(n1105), .A2(n1106), .A3(n1326), .ZN(n1325) );
INV_X1 U1025 ( .A(KEYINPUT22), .ZN(n1326) );
NAND2_X1 U1026 ( .A1(n1149), .A2(n1199), .ZN(n1106) );
XNOR2_X1 U1027 ( .A(n1327), .B(n1328), .ZN(n1149) );
XOR2_X1 U1028 ( .A(G137), .B(n1329), .Z(n1328) );
XNOR2_X1 U1029 ( .A(KEYINPUT48), .B(n1240), .ZN(n1329) );
XOR2_X1 U1030 ( .A(n1330), .B(n1331), .Z(n1327) );
XOR2_X1 U1031 ( .A(n1332), .B(n1333), .Z(n1331) );
NAND3_X1 U1032 ( .A1(n1127), .A2(n1334), .A3(KEYINPUT42), .ZN(n1333) );
NAND2_X1 U1033 ( .A1(n1335), .A2(n1336), .ZN(n1332) );
NAND2_X1 U1034 ( .A1(G110), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1035 ( .A(KEYINPUT10), .B(n1338), .Z(n1335) );
NOR2_X1 U1036 ( .A1(G110), .A2(n1337), .ZN(n1338) );
XNOR2_X1 U1037 ( .A(n1339), .B(G119), .ZN(n1337) );
NAND2_X1 U1038 ( .A1(n1340), .A2(G221), .ZN(n1330) );
INV_X1 U1039 ( .A(n1341), .ZN(n1105) );
NAND2_X1 U1040 ( .A1(KEYINPUT22), .A2(n1341), .ZN(n1324) );
NAND2_X1 U1041 ( .A1(G217), .A2(n1311), .ZN(n1341) );
NAND2_X1 U1042 ( .A1(G234), .A2(n1199), .ZN(n1311) );
XNOR2_X1 U1043 ( .A(n1256), .B(KEYINPUT47), .ZN(n1323) );
XOR2_X1 U1044 ( .A(G472), .B(n1102), .Z(n1256) );
AND2_X1 U1045 ( .A1(n1342), .A2(n1199), .ZN(n1102) );
NAND2_X1 U1046 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
OR3_X1 U1047 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1344) );
XOR2_X1 U1048 ( .A(KEYINPUT18), .B(n1348), .Z(n1343) );
NOR2_X1 U1049 ( .A1(n1349), .A2(n1168), .ZN(n1348) );
INV_X1 U1050 ( .A(n1345), .ZN(n1168) );
XOR2_X1 U1051 ( .A(n1350), .B(n1259), .Z(n1345) );
INV_X1 U1052 ( .A(G101), .ZN(n1259) );
NAND2_X1 U1053 ( .A1(G210), .A2(n1351), .ZN(n1350) );
NOR2_X1 U1054 ( .A1(n1346), .A2(n1347), .ZN(n1349) );
XNOR2_X1 U1055 ( .A(n1352), .B(KEYINPUT62), .ZN(n1347) );
NAND2_X1 U1056 ( .A1(n1178), .A2(n1183), .ZN(n1352) );
NOR2_X1 U1057 ( .A1(n1183), .A2(n1178), .ZN(n1346) );
INV_X1 U1058 ( .A(n1181), .ZN(n1178) );
XNOR2_X1 U1059 ( .A(n1131), .B(n1306), .ZN(n1181) );
INV_X1 U1060 ( .A(n1236), .ZN(n1306) );
XOR2_X1 U1061 ( .A(n1353), .B(n1339), .Z(n1236) );
INV_X1 U1062 ( .A(G128), .ZN(n1339) );
NAND2_X1 U1063 ( .A1(KEYINPUT2), .A2(n1322), .ZN(n1353) );
XNOR2_X1 U1064 ( .A(n1354), .B(n1355), .ZN(n1131) );
XOR2_X1 U1065 ( .A(KEYINPUT21), .B(G137), .Z(n1355) );
XNOR2_X1 U1066 ( .A(G131), .B(G134), .ZN(n1354) );
XOR2_X1 U1067 ( .A(G113), .B(n1356), .Z(n1183) );
XOR2_X1 U1068 ( .A(G119), .B(G116), .Z(n1356) );
NOR2_X1 U1069 ( .A1(n1242), .A2(n1093), .ZN(n1059) );
XOR2_X1 U1070 ( .A(G475), .B(n1357), .Z(n1093) );
AND2_X1 U1071 ( .A1(n1160), .A2(n1199), .ZN(n1357) );
INV_X1 U1072 ( .A(G902), .ZN(n1199) );
NAND2_X1 U1073 ( .A1(n1358), .A2(n1359), .ZN(n1160) );
NAND2_X1 U1074 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
XOR2_X1 U1075 ( .A(KEYINPUT54), .B(n1362), .Z(n1358) );
NOR2_X1 U1076 ( .A1(n1360), .A2(n1361), .ZN(n1362) );
XNOR2_X1 U1077 ( .A(n1363), .B(n1364), .ZN(n1361) );
XNOR2_X1 U1078 ( .A(G131), .B(n1365), .ZN(n1364) );
NAND3_X1 U1079 ( .A1(n1366), .A2(n1367), .A3(n1334), .ZN(n1365) );
INV_X1 U1080 ( .A(n1124), .ZN(n1334) );
NOR2_X1 U1081 ( .A1(n1234), .A2(n1194), .ZN(n1124) );
OR2_X1 U1082 ( .A1(n1127), .A2(KEYINPUT61), .ZN(n1367) );
NAND2_X1 U1083 ( .A1(n1234), .A2(n1194), .ZN(n1127) );
INV_X1 U1084 ( .A(G140), .ZN(n1194) );
INV_X1 U1085 ( .A(G125), .ZN(n1234) );
NAND2_X1 U1086 ( .A1(KEYINPUT61), .A2(G125), .ZN(n1366) );
XOR2_X1 U1087 ( .A(n1368), .B(n1322), .Z(n1363) );
XNOR2_X1 U1088 ( .A(G143), .B(n1240), .ZN(n1322) );
INV_X1 U1089 ( .A(G146), .ZN(n1240) );
NAND2_X1 U1090 ( .A1(G214), .A2(n1351), .ZN(n1368) );
NOR2_X1 U1091 ( .A1(G953), .A2(G237), .ZN(n1351) );
XOR2_X1 U1092 ( .A(n1369), .B(n1370), .Z(n1360) );
NOR2_X1 U1093 ( .A1(n1371), .A2(G104), .ZN(n1370) );
INV_X1 U1094 ( .A(KEYINPUT63), .ZN(n1371) );
NAND2_X1 U1095 ( .A1(n1372), .A2(n1373), .ZN(n1369) );
NAND2_X1 U1096 ( .A1(G113), .A2(n1291), .ZN(n1373) );
XOR2_X1 U1097 ( .A(n1374), .B(KEYINPUT9), .Z(n1372) );
NAND2_X1 U1098 ( .A1(G122), .A2(n1273), .ZN(n1374) );
INV_X1 U1099 ( .A(G113), .ZN(n1273) );
NAND2_X1 U1100 ( .A1(n1375), .A2(n1111), .ZN(n1242) );
NAND2_X1 U1101 ( .A1(n1097), .A2(n1098), .ZN(n1111) );
OR2_X1 U1102 ( .A1(n1098), .A2(n1097), .ZN(n1375) );
NOR2_X1 U1103 ( .A1(n1155), .A2(G902), .ZN(n1097) );
XOR2_X1 U1104 ( .A(n1376), .B(n1377), .Z(n1155) );
AND2_X1 U1105 ( .A1(n1340), .A2(G217), .ZN(n1377) );
AND2_X1 U1106 ( .A1(G234), .A2(n1053), .ZN(n1340) );
INV_X1 U1107 ( .A(G953), .ZN(n1053) );
NAND3_X1 U1108 ( .A1(n1378), .A2(n1379), .A3(n1380), .ZN(n1376) );
NAND2_X1 U1109 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
OR3_X1 U1110 ( .A1(n1382), .A2(n1381), .A3(n1383), .ZN(n1379) );
XNOR2_X1 U1111 ( .A(n1384), .B(n1385), .ZN(n1381) );
NOR2_X1 U1112 ( .A1(KEYINPUT4), .A2(n1251), .ZN(n1385) );
INV_X1 U1113 ( .A(G134), .ZN(n1251) );
XNOR2_X1 U1114 ( .A(G143), .B(G128), .ZN(n1384) );
OR2_X1 U1115 ( .A1(KEYINPUT55), .A2(n1386), .ZN(n1382) );
NAND2_X1 U1116 ( .A1(n1386), .A2(n1383), .ZN(n1378) );
INV_X1 U1117 ( .A(KEYINPUT26), .ZN(n1383) );
XOR2_X1 U1118 ( .A(n1387), .B(G107), .Z(n1386) );
NAND2_X1 U1119 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
NAND2_X1 U1120 ( .A1(G116), .A2(n1291), .ZN(n1389) );
XOR2_X1 U1121 ( .A(KEYINPUT57), .B(n1390), .Z(n1388) );
NOR2_X1 U1122 ( .A1(G116), .A2(n1291), .ZN(n1390) );
INV_X1 U1123 ( .A(G122), .ZN(n1291) );
INV_X1 U1124 ( .A(G478), .ZN(n1098) );
endmodule


