//Key = 0110001101011100100111111100000000011001110001001101001101000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394;

XNOR2_X1 U759 ( .A(G107), .B(n1055), .ZN(G9) );
NOR2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(G75) );
XOR2_X1 U761 ( .A(KEYINPUT8), .B(n1058), .Z(n1057) );
NOR3_X1 U762 ( .A1(n1059), .A2(G953), .A3(n1060), .ZN(n1058) );
XOR2_X1 U763 ( .A(KEYINPUT33), .B(G952), .Z(n1059) );
NOR4_X1 U764 ( .A1(n1061), .A2(n1062), .A3(G953), .A4(n1060), .ZN(n1056) );
AND4_X1 U765 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1060) );
NOR4_X1 U766 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
XNOR2_X1 U767 ( .A(n1071), .B(n1072), .ZN(n1070) );
NOR2_X1 U768 ( .A1(n1073), .A2(KEYINPUT3), .ZN(n1072) );
XNOR2_X1 U769 ( .A(n1074), .B(KEYINPUT23), .ZN(n1069) );
NAND3_X1 U770 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1067) );
XOR2_X1 U771 ( .A(n1078), .B(G475), .Z(n1077) );
OR2_X1 U772 ( .A1(G478), .A2(KEYINPUT16), .ZN(n1076) );
NAND3_X1 U773 ( .A1(G478), .A2(n1079), .A3(KEYINPUT16), .ZN(n1075) );
NOR3_X1 U774 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1065) );
NAND2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(n1063) );
NOR2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1062) );
NOR2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR3_X1 U778 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
NOR3_X1 U779 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1090) );
NOR2_X1 U780 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XNOR2_X1 U781 ( .A(KEYINPUT41), .B(n1097), .ZN(n1096) );
NOR4_X1 U782 ( .A1(KEYINPUT50), .A2(n1098), .A3(n1097), .A4(n1064), .ZN(n1093) );
NOR2_X1 U783 ( .A1(n1099), .A2(n1100), .ZN(n1092) );
NOR3_X1 U784 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1099) );
NOR2_X1 U785 ( .A1(n1097), .A2(n1104), .ZN(n1102) );
INV_X1 U786 ( .A(KEYINPUT50), .ZN(n1104) );
XOR2_X1 U787 ( .A(KEYINPUT53), .B(n1105), .Z(n1101) );
NOR2_X1 U788 ( .A1(n1074), .A2(n1106), .ZN(n1105) );
NOR3_X1 U789 ( .A1(n1097), .A2(n1107), .A3(n1100), .ZN(n1087) );
INV_X1 U790 ( .A(n1108), .ZN(n1100) );
NOR3_X1 U791 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1107) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1091), .ZN(n1111) );
NOR2_X1 U793 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR3_X1 U794 ( .A1(n1115), .A2(n1116), .A3(n1068), .ZN(n1110) );
XNOR2_X1 U795 ( .A(KEYINPUT7), .B(n1089), .ZN(n1115) );
AND2_X1 U796 ( .A1(n1117), .A2(n1118), .ZN(n1109) );
NAND3_X1 U797 ( .A1(n1119), .A2(G952), .A3(n1120), .ZN(n1061) );
XOR2_X1 U798 ( .A(n1121), .B(n1122), .Z(G72) );
NAND2_X1 U799 ( .A1(G953), .A2(n1123), .ZN(n1122) );
NAND2_X1 U800 ( .A1(G900), .A2(G227), .ZN(n1123) );
NAND2_X1 U801 ( .A1(KEYINPUT35), .A2(n1124), .ZN(n1121) );
XOR2_X1 U802 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U803 ( .A1(n1119), .A2(G953), .ZN(n1126) );
NOR2_X1 U804 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
XOR2_X1 U805 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U806 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U807 ( .A(n1133), .B(n1134), .ZN(n1132) );
NOR2_X1 U808 ( .A1(KEYINPUT43), .A2(n1135), .ZN(n1134) );
NAND2_X1 U809 ( .A1(KEYINPUT39), .A2(n1136), .ZN(n1133) );
XNOR2_X1 U810 ( .A(n1137), .B(n1138), .ZN(n1129) );
XOR2_X1 U811 ( .A(G134), .B(G131), .Z(n1138) );
XOR2_X1 U812 ( .A(n1139), .B(n1140), .Z(G69) );
NOR2_X1 U813 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
AND2_X1 U814 ( .A1(G224), .A2(G898), .ZN(n1141) );
NAND2_X1 U815 ( .A1(n1143), .A2(n1144), .ZN(n1139) );
NAND2_X1 U816 ( .A1(KEYINPUT60), .A2(n1145), .ZN(n1144) );
XOR2_X1 U817 ( .A(n1146), .B(n1147), .Z(n1143) );
NOR2_X1 U818 ( .A1(n1120), .A2(G953), .ZN(n1147) );
OR2_X1 U819 ( .A1(n1145), .A2(KEYINPUT60), .ZN(n1146) );
NAND2_X1 U820 ( .A1(n1148), .A2(n1149), .ZN(n1145) );
NAND2_X1 U821 ( .A1(G953), .A2(n1150), .ZN(n1149) );
XNOR2_X1 U822 ( .A(n1151), .B(n1152), .ZN(n1148) );
XNOR2_X1 U823 ( .A(n1153), .B(n1154), .ZN(n1151) );
NAND2_X1 U824 ( .A1(KEYINPUT49), .A2(n1155), .ZN(n1154) );
NAND2_X1 U825 ( .A1(KEYINPUT22), .A2(n1156), .ZN(n1153) );
INV_X1 U826 ( .A(n1157), .ZN(n1156) );
NOR2_X1 U827 ( .A1(n1158), .A2(n1159), .ZN(G66) );
NOR3_X1 U828 ( .A1(n1071), .A2(n1160), .A3(n1161), .ZN(n1159) );
NOR2_X1 U829 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NOR2_X1 U830 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
NOR2_X1 U831 ( .A1(n1166), .A2(n1167), .ZN(n1164) );
AND3_X1 U832 ( .A1(n1163), .A2(n1073), .A3(n1168), .ZN(n1160) );
INV_X1 U833 ( .A(n1165), .ZN(n1073) );
NOR2_X1 U834 ( .A1(n1158), .A2(n1169), .ZN(G63) );
XNOR2_X1 U835 ( .A(n1170), .B(n1171), .ZN(n1169) );
AND2_X1 U836 ( .A1(G478), .A2(n1168), .ZN(n1171) );
NOR2_X1 U837 ( .A1(n1158), .A2(n1172), .ZN(G60) );
XOR2_X1 U838 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U839 ( .A(KEYINPUT13), .B(n1175), .Z(n1174) );
AND2_X1 U840 ( .A1(G475), .A2(n1168), .ZN(n1175) );
NAND2_X1 U841 ( .A1(n1176), .A2(n1177), .ZN(G6) );
NAND2_X1 U842 ( .A1(G104), .A2(n1178), .ZN(n1177) );
XOR2_X1 U843 ( .A(n1179), .B(KEYINPUT10), .Z(n1176) );
OR2_X1 U844 ( .A1(n1178), .A2(G104), .ZN(n1179) );
NOR2_X1 U845 ( .A1(n1180), .A2(n1181), .ZN(G57) );
XOR2_X1 U846 ( .A(n1182), .B(n1183), .Z(n1181) );
NOR2_X1 U847 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U848 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NOR2_X1 U849 ( .A1(n1188), .A2(KEYINPUT18), .ZN(n1186) );
AND2_X1 U850 ( .A1(n1189), .A2(KEYINPUT63), .ZN(n1188) );
NOR2_X1 U851 ( .A1(n1190), .A2(n1189), .ZN(n1184) );
NAND2_X1 U852 ( .A1(n1168), .A2(G472), .ZN(n1189) );
INV_X1 U853 ( .A(n1191), .ZN(n1168) );
NOR2_X1 U854 ( .A1(n1192), .A2(n1193), .ZN(n1190) );
INV_X1 U855 ( .A(KEYINPUT63), .ZN(n1193) );
NOR2_X1 U856 ( .A1(KEYINPUT18), .A2(n1194), .ZN(n1192) );
XOR2_X1 U857 ( .A(n1195), .B(n1196), .Z(n1182) );
NOR2_X1 U858 ( .A1(KEYINPUT32), .A2(G101), .ZN(n1196) );
NOR2_X1 U859 ( .A1(n1197), .A2(n1142), .ZN(n1180) );
XNOR2_X1 U860 ( .A(G952), .B(KEYINPUT36), .ZN(n1197) );
NOR2_X1 U861 ( .A1(n1158), .A2(n1198), .ZN(G54) );
XOR2_X1 U862 ( .A(n1199), .B(n1200), .Z(n1198) );
XNOR2_X1 U863 ( .A(n1201), .B(n1202), .ZN(n1200) );
XNOR2_X1 U864 ( .A(n1203), .B(n1204), .ZN(n1201) );
NOR2_X1 U865 ( .A1(n1084), .A2(n1191), .ZN(n1204) );
XOR2_X1 U866 ( .A(n1205), .B(n1206), .Z(n1199) );
XNOR2_X1 U867 ( .A(KEYINPUT34), .B(n1207), .ZN(n1206) );
NAND2_X1 U868 ( .A1(KEYINPUT19), .A2(n1208), .ZN(n1205) );
XOR2_X1 U869 ( .A(KEYINPUT62), .B(n1209), .Z(n1208) );
NOR2_X1 U870 ( .A1(n1158), .A2(n1210), .ZN(G51) );
XOR2_X1 U871 ( .A(KEYINPUT28), .B(n1211), .Z(n1210) );
NOR2_X1 U872 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XOR2_X1 U873 ( .A(KEYINPUT52), .B(n1214), .Z(n1213) );
NOR3_X1 U874 ( .A1(n1215), .A2(n1216), .A3(n1191), .ZN(n1214) );
INV_X1 U875 ( .A(n1217), .ZN(n1215) );
NOR2_X1 U876 ( .A1(n1218), .A2(n1217), .ZN(n1212) );
XNOR2_X1 U877 ( .A(n1219), .B(n1220), .ZN(n1217) );
XOR2_X1 U878 ( .A(KEYINPUT57), .B(n1221), .Z(n1220) );
XOR2_X1 U879 ( .A(n1222), .B(n1223), .Z(n1219) );
NAND2_X1 U880 ( .A1(KEYINPUT25), .A2(n1224), .ZN(n1222) );
NOR2_X1 U881 ( .A1(n1216), .A2(n1191), .ZN(n1218) );
NAND2_X1 U882 ( .A1(G902), .A2(n1225), .ZN(n1191) );
NAND2_X1 U883 ( .A1(n1120), .A2(n1119), .ZN(n1225) );
INV_X1 U884 ( .A(n1166), .ZN(n1119) );
NAND2_X1 U885 ( .A1(n1226), .A2(n1227), .ZN(n1166) );
NOR4_X1 U886 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1227) );
INV_X1 U887 ( .A(n1232), .ZN(n1231) );
AND4_X1 U888 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1226) );
INV_X1 U889 ( .A(n1167), .ZN(n1120) );
NAND2_X1 U890 ( .A1(n1237), .A2(n1238), .ZN(n1167) );
AND4_X1 U891 ( .A1(n1055), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1238) );
NAND3_X1 U892 ( .A1(n1113), .A2(n1242), .A3(n1243), .ZN(n1055) );
AND4_X1 U893 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1178), .ZN(n1237) );
NAND3_X1 U894 ( .A1(n1243), .A2(n1242), .A3(n1114), .ZN(n1178) );
NOR2_X1 U895 ( .A1(n1142), .A2(G952), .ZN(n1158) );
XNOR2_X1 U896 ( .A(G146), .B(n1236), .ZN(G48) );
NAND4_X1 U897 ( .A1(n1247), .A2(n1248), .A3(n1114), .A4(n1068), .ZN(n1236) );
XOR2_X1 U898 ( .A(n1235), .B(n1249), .Z(G45) );
XNOR2_X1 U899 ( .A(G143), .B(KEYINPUT26), .ZN(n1249) );
NAND4_X1 U900 ( .A1(n1250), .A2(n1118), .A3(n1247), .A4(n1251), .ZN(n1235) );
NOR3_X1 U901 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1251) );
INV_X1 U902 ( .A(n1095), .ZN(n1247) );
XOR2_X1 U903 ( .A(n1234), .B(n1255), .Z(G42) );
XNOR2_X1 U904 ( .A(G140), .B(KEYINPUT47), .ZN(n1255) );
NAND4_X1 U905 ( .A1(n1256), .A2(n1114), .A3(n1257), .A4(n1258), .ZN(n1234) );
XOR2_X1 U906 ( .A(G137), .B(n1230), .Z(G39) );
AND4_X1 U907 ( .A1(n1256), .A2(n1117), .A3(n1258), .A4(n1068), .ZN(n1230) );
XOR2_X1 U908 ( .A(G134), .B(n1229), .Z(G36) );
AND3_X1 U909 ( .A1(n1118), .A2(n1113), .A3(n1256), .ZN(n1229) );
XOR2_X1 U910 ( .A(G131), .B(n1228), .Z(G33) );
AND3_X1 U911 ( .A1(n1114), .A2(n1118), .A3(n1256), .ZN(n1228) );
NOR3_X1 U912 ( .A1(n1095), .A2(n1253), .A3(n1097), .ZN(n1256) );
NAND2_X1 U913 ( .A1(n1259), .A2(n1106), .ZN(n1097) );
XOR2_X1 U914 ( .A(n1260), .B(KEYINPUT55), .Z(n1095) );
XNOR2_X1 U915 ( .A(G128), .B(n1233), .ZN(G30) );
NAND4_X1 U916 ( .A1(n1248), .A2(n1113), .A3(n1260), .A4(n1068), .ZN(n1233) );
XNOR2_X1 U917 ( .A(G101), .B(n1246), .ZN(G3) );
NAND3_X1 U918 ( .A1(n1117), .A2(n1243), .A3(n1118), .ZN(n1246) );
XNOR2_X1 U919 ( .A(G125), .B(n1232), .ZN(G27) );
NAND4_X1 U920 ( .A1(n1248), .A2(n1114), .A3(n1257), .A4(n1108), .ZN(n1232) );
NOR3_X1 U921 ( .A1(n1116), .A2(n1253), .A3(n1254), .ZN(n1248) );
INV_X1 U922 ( .A(n1103), .ZN(n1254) );
AND2_X1 U923 ( .A1(n1261), .A2(n1086), .ZN(n1253) );
NAND3_X1 U924 ( .A1(G902), .A2(n1262), .A3(n1127), .ZN(n1261) );
NOR2_X1 U925 ( .A1(n1142), .A2(G900), .ZN(n1127) );
XNOR2_X1 U926 ( .A(G122), .B(n1245), .ZN(G24) );
OR4_X1 U927 ( .A1(n1263), .A2(n1264), .A3(n1252), .A4(n1091), .ZN(n1245) );
INV_X1 U928 ( .A(n1242), .ZN(n1091) );
NOR2_X1 U929 ( .A1(n1068), .A2(n1258), .ZN(n1242) );
XNOR2_X1 U930 ( .A(G119), .B(n1244), .ZN(G21) );
NAND4_X1 U931 ( .A1(n1265), .A2(n1117), .A3(n1258), .A4(n1068), .ZN(n1244) );
XOR2_X1 U932 ( .A(n1241), .B(n1266), .Z(G18) );
XNOR2_X1 U933 ( .A(KEYINPUT2), .B(n1267), .ZN(n1266) );
NAND3_X1 U934 ( .A1(n1265), .A2(n1113), .A3(n1118), .ZN(n1241) );
NOR2_X1 U935 ( .A1(n1252), .A2(n1250), .ZN(n1113) );
XOR2_X1 U936 ( .A(n1268), .B(KEYINPUT5), .Z(n1252) );
XNOR2_X1 U937 ( .A(G113), .B(n1240), .ZN(G15) );
NAND3_X1 U938 ( .A1(n1118), .A2(n1265), .A3(n1114), .ZN(n1240) );
AND2_X1 U939 ( .A1(n1250), .A2(n1268), .ZN(n1114) );
INV_X1 U940 ( .A(n1263), .ZN(n1250) );
INV_X1 U941 ( .A(n1264), .ZN(n1265) );
NAND2_X1 U942 ( .A1(n1108), .A2(n1269), .ZN(n1264) );
NOR2_X1 U943 ( .A1(n1098), .A2(n1270), .ZN(n1108) );
INV_X1 U944 ( .A(n1064), .ZN(n1270) );
NOR2_X1 U945 ( .A1(n1258), .A2(n1257), .ZN(n1118) );
XOR2_X1 U946 ( .A(n1239), .B(n1271), .Z(G12) );
XNOR2_X1 U947 ( .A(KEYINPUT40), .B(n1272), .ZN(n1271) );
NAND4_X1 U948 ( .A1(n1117), .A2(n1243), .A3(n1257), .A4(n1258), .ZN(n1239) );
INV_X1 U949 ( .A(n1116), .ZN(n1258) );
XOR2_X1 U950 ( .A(n1071), .B(n1165), .Z(n1116) );
NAND2_X1 U951 ( .A1(G217), .A2(n1273), .ZN(n1165) );
NOR2_X1 U952 ( .A1(n1163), .A2(G902), .ZN(n1071) );
XOR2_X1 U953 ( .A(n1274), .B(n1275), .Z(n1163) );
XNOR2_X1 U954 ( .A(n1276), .B(n1277), .ZN(n1275) );
NAND2_X1 U955 ( .A1(n1278), .A2(G221), .ZN(n1276) );
NAND2_X1 U956 ( .A1(n1279), .A2(n1280), .ZN(n1274) );
NAND2_X1 U957 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND2_X1 U958 ( .A1(n1283), .A2(n1284), .ZN(n1281) );
NAND2_X1 U959 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND2_X1 U960 ( .A1(n1287), .A2(n1288), .ZN(n1283) );
NAND2_X1 U961 ( .A1(n1289), .A2(n1290), .ZN(n1279) );
NAND2_X1 U962 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
NAND2_X1 U963 ( .A1(n1288), .A2(n1286), .ZN(n1292) );
INV_X1 U964 ( .A(n1285), .ZN(n1288) );
NAND2_X1 U965 ( .A1(n1285), .A2(n1287), .ZN(n1291) );
XOR2_X1 U966 ( .A(n1286), .B(KEYINPUT20), .Z(n1287) );
NAND2_X1 U967 ( .A1(n1293), .A2(n1294), .ZN(n1286) );
NAND2_X1 U968 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
XNOR2_X1 U969 ( .A(KEYINPUT1), .B(n1272), .ZN(n1296) );
XNOR2_X1 U970 ( .A(n1297), .B(G119), .ZN(n1295) );
INV_X1 U971 ( .A(G128), .ZN(n1297) );
NAND2_X1 U972 ( .A1(n1298), .A2(n1299), .ZN(n1293) );
XNOR2_X1 U973 ( .A(KEYINPUT46), .B(n1272), .ZN(n1299) );
XNOR2_X1 U974 ( .A(G119), .B(G128), .ZN(n1298) );
NOR2_X1 U975 ( .A1(G146), .A2(KEYINPUT37), .ZN(n1285) );
INV_X1 U976 ( .A(n1068), .ZN(n1257) );
XNOR2_X1 U977 ( .A(n1300), .B(G472), .ZN(n1068) );
NAND2_X1 U978 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
XNOR2_X1 U979 ( .A(n1187), .B(n1303), .ZN(n1301) );
XNOR2_X1 U980 ( .A(G101), .B(n1195), .ZN(n1303) );
NAND3_X1 U981 ( .A1(n1304), .A2(n1142), .A3(G210), .ZN(n1195) );
INV_X1 U982 ( .A(n1194), .ZN(n1187) );
XNOR2_X1 U983 ( .A(n1305), .B(n1306), .ZN(n1194) );
XNOR2_X1 U984 ( .A(n1203), .B(n1307), .ZN(n1306) );
XOR2_X1 U985 ( .A(n1152), .B(KEYINPUT59), .Z(n1305) );
AND2_X1 U986 ( .A1(n1269), .A2(n1260), .ZN(n1243) );
AND2_X1 U987 ( .A1(n1064), .A2(n1098), .ZN(n1260) );
NAND2_X1 U988 ( .A1(n1308), .A2(n1309), .ZN(n1098) );
NAND2_X1 U989 ( .A1(n1310), .A2(n1084), .ZN(n1309) );
NAND2_X1 U990 ( .A1(KEYINPUT11), .A2(n1311), .ZN(n1310) );
NAND2_X1 U991 ( .A1(n1081), .A2(KEYINPUT11), .ZN(n1308) );
NOR2_X1 U992 ( .A1(n1084), .A2(n1083), .ZN(n1081) );
INV_X1 U993 ( .A(n1311), .ZN(n1083) );
NAND2_X1 U994 ( .A1(n1312), .A2(n1302), .ZN(n1311) );
XOR2_X1 U995 ( .A(n1209), .B(n1313), .Z(n1312) );
XNOR2_X1 U996 ( .A(n1314), .B(n1315), .ZN(n1313) );
NOR2_X1 U997 ( .A1(KEYINPUT30), .A2(n1207), .ZN(n1315) );
NAND2_X1 U998 ( .A1(G227), .A2(n1142), .ZN(n1207) );
NAND4_X1 U999 ( .A1(KEYINPUT6), .A2(n1316), .A3(n1317), .A4(n1318), .ZN(n1314) );
NAND2_X1 U1000 ( .A1(KEYINPUT14), .A2(n1319), .ZN(n1318) );
NAND2_X1 U1001 ( .A1(n1320), .A2(n1203), .ZN(n1319) );
XNOR2_X1 U1002 ( .A(KEYINPUT9), .B(n1202), .ZN(n1320) );
NAND2_X1 U1003 ( .A1(n1321), .A2(n1322), .ZN(n1317) );
INV_X1 U1004 ( .A(KEYINPUT14), .ZN(n1322) );
NAND2_X1 U1005 ( .A1(n1323), .A2(n1324), .ZN(n1321) );
NAND3_X1 U1006 ( .A1(KEYINPUT9), .A2(n1203), .A3(n1202), .ZN(n1324) );
OR2_X1 U1007 ( .A1(n1202), .A2(KEYINPUT9), .ZN(n1323) );
OR2_X1 U1008 ( .A1(n1203), .A2(n1202), .ZN(n1316) );
XOR2_X1 U1009 ( .A(n1325), .B(n1131), .Z(n1202) );
XNOR2_X1 U1010 ( .A(n1326), .B(n1327), .ZN(n1131) );
NAND2_X1 U1011 ( .A1(n1328), .A2(n1329), .ZN(n1326) );
XOR2_X1 U1012 ( .A(KEYINPUT51), .B(KEYINPUT38), .Z(n1328) );
NAND3_X1 U1013 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n1325) );
OR2_X1 U1014 ( .A1(n1333), .A2(KEYINPUT31), .ZN(n1331) );
NAND2_X1 U1015 ( .A1(n1334), .A2(KEYINPUT31), .ZN(n1330) );
XNOR2_X1 U1016 ( .A(n1335), .B(n1336), .ZN(n1334) );
NOR2_X1 U1017 ( .A1(G104), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1018 ( .A(G131), .B(n1338), .Z(n1203) );
NOR2_X1 U1019 ( .A1(KEYINPUT56), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1020 ( .A(n1340), .B(G134), .Z(n1339) );
NAND2_X1 U1021 ( .A1(KEYINPUT45), .A2(n1341), .ZN(n1340) );
XNOR2_X1 U1022 ( .A(KEYINPUT42), .B(n1135), .ZN(n1341) );
INV_X1 U1023 ( .A(n1277), .ZN(n1135) );
XOR2_X1 U1024 ( .A(G137), .B(KEYINPUT48), .Z(n1277) );
XNOR2_X1 U1025 ( .A(n1272), .B(G140), .ZN(n1209) );
INV_X1 U1026 ( .A(G110), .ZN(n1272) );
INV_X1 U1027 ( .A(G469), .ZN(n1084) );
NAND2_X1 U1028 ( .A1(G221), .A2(n1273), .ZN(n1064) );
NAND2_X1 U1029 ( .A1(G234), .A2(n1302), .ZN(n1273) );
AND2_X1 U1030 ( .A1(n1103), .A2(n1342), .ZN(n1269) );
NAND2_X1 U1031 ( .A1(n1086), .A2(n1343), .ZN(n1342) );
NAND4_X1 U1032 ( .A1(G902), .A2(G953), .A3(n1262), .A4(n1150), .ZN(n1343) );
INV_X1 U1033 ( .A(G898), .ZN(n1150) );
NAND3_X1 U1034 ( .A1(n1262), .A2(n1142), .A3(G952), .ZN(n1086) );
NAND2_X1 U1035 ( .A1(G237), .A2(G234), .ZN(n1262) );
NOR2_X1 U1036 ( .A1(n1259), .A2(n1080), .ZN(n1103) );
INV_X1 U1037 ( .A(n1106), .ZN(n1080) );
NAND2_X1 U1038 ( .A1(G214), .A2(n1344), .ZN(n1106) );
INV_X1 U1039 ( .A(n1074), .ZN(n1259) );
XOR2_X1 U1040 ( .A(n1345), .B(n1216), .Z(n1074) );
NAND2_X1 U1041 ( .A1(G210), .A2(n1344), .ZN(n1216) );
NAND2_X1 U1042 ( .A1(n1304), .A2(n1302), .ZN(n1344) );
NAND2_X1 U1043 ( .A1(n1346), .A2(n1302), .ZN(n1345) );
XNOR2_X1 U1044 ( .A(n1223), .B(n1347), .ZN(n1346) );
XNOR2_X1 U1045 ( .A(n1224), .B(n1221), .ZN(n1347) );
AND2_X1 U1046 ( .A1(n1348), .A2(n1349), .ZN(n1221) );
NAND2_X1 U1047 ( .A1(n1157), .A2(n1350), .ZN(n1349) );
XOR2_X1 U1048 ( .A(n1351), .B(KEYINPUT17), .Z(n1348) );
OR2_X1 U1049 ( .A1(n1350), .A2(n1157), .ZN(n1351) );
XOR2_X1 U1050 ( .A(G110), .B(G122), .Z(n1157) );
NAND3_X1 U1051 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1350) );
NAND2_X1 U1052 ( .A1(n1152), .A2(n1155), .ZN(n1354) );
NAND2_X1 U1053 ( .A1(KEYINPUT27), .A2(n1355), .ZN(n1353) );
NAND2_X1 U1054 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
XNOR2_X1 U1055 ( .A(KEYINPUT58), .B(n1152), .ZN(n1357) );
INV_X1 U1056 ( .A(n1155), .ZN(n1356) );
NAND2_X1 U1057 ( .A1(n1358), .A2(n1359), .ZN(n1352) );
INV_X1 U1058 ( .A(KEYINPUT27), .ZN(n1359) );
NAND2_X1 U1059 ( .A1(n1360), .A2(n1361), .ZN(n1358) );
OR3_X1 U1060 ( .A1(n1155), .A2(n1152), .A3(KEYINPUT58), .ZN(n1361) );
NAND2_X1 U1061 ( .A1(n1333), .A2(n1332), .ZN(n1155) );
NAND3_X1 U1062 ( .A1(G101), .A2(n1337), .A3(G104), .ZN(n1332) );
INV_X1 U1063 ( .A(G107), .ZN(n1337) );
AND2_X1 U1064 ( .A1(n1362), .A2(n1363), .ZN(n1333) );
OR3_X1 U1065 ( .A1(G101), .A2(G104), .A3(G107), .ZN(n1363) );
NAND2_X1 U1066 ( .A1(n1364), .A2(G107), .ZN(n1362) );
XNOR2_X1 U1067 ( .A(G104), .B(n1335), .ZN(n1364) );
INV_X1 U1068 ( .A(G101), .ZN(n1335) );
NAND2_X1 U1069 ( .A1(KEYINPUT58), .A2(n1152), .ZN(n1360) );
XNOR2_X1 U1070 ( .A(G113), .B(n1365), .ZN(n1152) );
XNOR2_X1 U1071 ( .A(G119), .B(n1267), .ZN(n1365) );
AND2_X1 U1072 ( .A1(n1366), .A2(G224), .ZN(n1224) );
XNOR2_X1 U1073 ( .A(G953), .B(KEYINPUT29), .ZN(n1366) );
XOR2_X1 U1074 ( .A(n1307), .B(n1137), .Z(n1223) );
INV_X1 U1075 ( .A(G125), .ZN(n1137) );
NAND2_X1 U1076 ( .A1(n1367), .A2(n1368), .ZN(n1307) );
NAND2_X1 U1077 ( .A1(n1369), .A2(n1329), .ZN(n1368) );
XOR2_X1 U1078 ( .A(KEYINPUT24), .B(n1327), .Z(n1369) );
NAND2_X1 U1079 ( .A1(G146), .A2(n1370), .ZN(n1367) );
XNOR2_X1 U1080 ( .A(n1327), .B(KEYINPUT21), .ZN(n1370) );
INV_X1 U1081 ( .A(n1089), .ZN(n1117) );
NAND2_X1 U1082 ( .A1(n1268), .A2(n1263), .ZN(n1089) );
XNOR2_X1 U1083 ( .A(n1078), .B(n1371), .ZN(n1263) );
XOR2_X1 U1084 ( .A(KEYINPUT4), .B(n1372), .Z(n1371) );
NOR2_X1 U1085 ( .A1(KEYINPUT44), .A2(G475), .ZN(n1372) );
NAND2_X1 U1086 ( .A1(n1173), .A2(n1302), .ZN(n1078) );
XOR2_X1 U1087 ( .A(n1373), .B(n1374), .Z(n1173) );
XOR2_X1 U1088 ( .A(G113), .B(n1375), .Z(n1374) );
XNOR2_X1 U1089 ( .A(n1329), .B(G122), .ZN(n1375) );
INV_X1 U1090 ( .A(G146), .ZN(n1329) );
XNOR2_X1 U1091 ( .A(n1376), .B(n1282), .ZN(n1373) );
INV_X1 U1092 ( .A(n1289), .ZN(n1282) );
XNOR2_X1 U1093 ( .A(G125), .B(n1136), .ZN(n1289) );
INV_X1 U1094 ( .A(G140), .ZN(n1136) );
XOR2_X1 U1095 ( .A(n1377), .B(G104), .Z(n1376) );
NAND2_X1 U1096 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
OR2_X1 U1097 ( .A1(n1380), .A2(G131), .ZN(n1379) );
XOR2_X1 U1098 ( .A(n1381), .B(KEYINPUT15), .Z(n1378) );
NAND2_X1 U1099 ( .A1(G131), .A2(n1380), .ZN(n1381) );
XNOR2_X1 U1100 ( .A(n1382), .B(n1383), .ZN(n1380) );
XOR2_X1 U1101 ( .A(n1384), .B(KEYINPUT0), .Z(n1382) );
NAND3_X1 U1102 ( .A1(n1385), .A2(n1304), .A3(G214), .ZN(n1384) );
INV_X1 U1103 ( .A(G237), .ZN(n1304) );
XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1142), .ZN(n1385) );
NOR2_X1 U1105 ( .A1(n1082), .A2(n1386), .ZN(n1268) );
AND2_X1 U1106 ( .A1(G478), .A2(n1079), .ZN(n1386) );
NOR2_X1 U1107 ( .A1(n1079), .A2(G478), .ZN(n1082) );
NAND2_X1 U1108 ( .A1(n1170), .A2(n1302), .ZN(n1079) );
INV_X1 U1109 ( .A(G902), .ZN(n1302) );
XNOR2_X1 U1110 ( .A(n1387), .B(n1388), .ZN(n1170) );
XOR2_X1 U1111 ( .A(n1389), .B(n1390), .Z(n1388) );
XNOR2_X1 U1112 ( .A(G134), .B(G107), .ZN(n1390) );
NAND2_X1 U1113 ( .A1(n1391), .A2(n1392), .ZN(n1389) );
NAND2_X1 U1114 ( .A1(G122), .A2(n1267), .ZN(n1392) );
XOR2_X1 U1115 ( .A(KEYINPUT12), .B(n1393), .Z(n1391) );
NOR2_X1 U1116 ( .A1(G122), .A2(n1267), .ZN(n1393) );
INV_X1 U1117 ( .A(G116), .ZN(n1267) );
XNOR2_X1 U1118 ( .A(n1327), .B(n1394), .ZN(n1387) );
AND2_X1 U1119 ( .A1(n1278), .A2(G217), .ZN(n1394) );
AND2_X1 U1120 ( .A1(G234), .A2(n1142), .ZN(n1278) );
INV_X1 U1121 ( .A(G953), .ZN(n1142) );
XOR2_X1 U1122 ( .A(G128), .B(n1383), .Z(n1327) );
XOR2_X1 U1123 ( .A(G143), .B(KEYINPUT54), .Z(n1383) );
endmodule


