//Key = 1101001001110101100011001001000001101110100111010110110001110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321;

XNOR2_X1 U730 ( .A(G107), .B(n1001), .ZN(G9) );
NOR2_X1 U731 ( .A1(n1002), .A2(n1003), .ZN(G75) );
NOR3_X1 U732 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1003) );
NAND3_X1 U733 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1004) );
NAND2_X1 U734 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND2_X1 U735 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND4_X1 U736 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1013) );
NAND2_X1 U737 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NAND2_X1 U738 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
OR2_X1 U739 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U740 ( .A1(n1024), .A2(n1025), .ZN(n1018) );
NAND2_X1 U741 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U742 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND3_X1 U743 ( .A1(n1020), .A2(n1030), .A3(n1024), .ZN(n1012) );
NAND2_X1 U744 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND3_X1 U745 ( .A1(n1033), .A2(n1034), .A3(n1014), .ZN(n1032) );
OR2_X1 U746 ( .A1(n1017), .A2(n1015), .ZN(n1034) );
NAND3_X1 U747 ( .A1(n1035), .A2(n1036), .A3(n1017), .ZN(n1033) );
NAND2_X1 U748 ( .A1(n1015), .A2(n1037), .ZN(n1031) );
INV_X1 U749 ( .A(n1038), .ZN(n1010) );
NOR3_X1 U750 ( .A1(n1039), .A2(G953), .A3(n1040), .ZN(n1002) );
INV_X1 U751 ( .A(n1007), .ZN(n1040) );
NAND4_X1 U752 ( .A1(n1041), .A2(n1024), .A3(n1042), .A4(n1043), .ZN(n1007) );
NOR3_X1 U753 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
XOR2_X1 U754 ( .A(n1047), .B(n1048), .Z(n1046) );
XNOR2_X1 U755 ( .A(KEYINPUT8), .B(n1049), .ZN(n1048) );
NAND2_X1 U756 ( .A1(KEYINPUT16), .A2(n1050), .ZN(n1047) );
XNOR2_X1 U757 ( .A(n1051), .B(n1052), .ZN(n1042) );
XNOR2_X1 U758 ( .A(n1053), .B(KEYINPUT46), .ZN(n1051) );
XNOR2_X1 U759 ( .A(n1054), .B(KEYINPUT17), .ZN(n1041) );
XNOR2_X1 U760 ( .A(KEYINPUT54), .B(n1005), .ZN(n1039) );
INV_X1 U761 ( .A(G952), .ZN(n1005) );
XOR2_X1 U762 ( .A(n1055), .B(n1056), .Z(G72) );
XOR2_X1 U763 ( .A(n1057), .B(n1058), .Z(n1056) );
NOR2_X1 U764 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XNOR2_X1 U765 ( .A(G953), .B(KEYINPUT40), .ZN(n1060) );
INV_X1 U766 ( .A(n1061), .ZN(n1059) );
NAND2_X1 U767 ( .A1(n1062), .A2(n1063), .ZN(n1057) );
OR2_X1 U768 ( .A1(n1008), .A2(G900), .ZN(n1063) );
XOR2_X1 U769 ( .A(n1064), .B(n1065), .Z(n1062) );
XOR2_X1 U770 ( .A(n1066), .B(n1067), .Z(n1065) );
XNOR2_X1 U771 ( .A(G125), .B(n1068), .ZN(n1067) );
NAND2_X1 U772 ( .A1(KEYINPUT58), .A2(G140), .ZN(n1068) );
XOR2_X1 U773 ( .A(n1069), .B(n1070), .Z(n1064) );
XOR2_X1 U774 ( .A(G134), .B(G131), .Z(n1070) );
XNOR2_X1 U775 ( .A(KEYINPUT30), .B(n1071), .ZN(n1069) );
NAND2_X1 U776 ( .A1(G953), .A2(n1072), .ZN(n1055) );
NAND2_X1 U777 ( .A1(G900), .A2(G227), .ZN(n1072) );
XOR2_X1 U778 ( .A(n1073), .B(n1074), .Z(G69) );
NOR2_X1 U779 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
XOR2_X1 U780 ( .A(n1077), .B(n1078), .Z(n1076) );
NOR2_X1 U781 ( .A1(KEYINPUT7), .A2(n1079), .ZN(n1078) );
XOR2_X1 U782 ( .A(n1080), .B(n1081), .Z(n1079) );
NAND2_X1 U783 ( .A1(KEYINPUT44), .A2(n1082), .ZN(n1080) );
NOR2_X1 U784 ( .A1(G898), .A2(n1008), .ZN(n1075) );
NAND3_X1 U785 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1073) );
NAND2_X1 U786 ( .A1(n1086), .A2(n1008), .ZN(n1085) );
OR3_X1 U787 ( .A1(n1087), .A2(n1008), .A3(KEYINPUT27), .ZN(n1084) );
NAND3_X1 U788 ( .A1(G953), .A2(n1087), .A3(KEYINPUT27), .ZN(n1083) );
NAND2_X1 U789 ( .A1(G898), .A2(G224), .ZN(n1087) );
NOR2_X1 U790 ( .A1(n1088), .A2(n1089), .ZN(G66) );
NOR3_X1 U791 ( .A1(n1053), .A2(n1090), .A3(n1091), .ZN(n1089) );
NOR3_X1 U792 ( .A1(n1092), .A2(n1052), .A3(n1093), .ZN(n1091) );
NOR2_X1 U793 ( .A1(n1094), .A2(n1095), .ZN(n1090) );
NOR2_X1 U794 ( .A1(n1096), .A2(n1052), .ZN(n1094) );
NOR2_X1 U795 ( .A1(n1088), .A2(n1097), .ZN(G63) );
XNOR2_X1 U796 ( .A(n1098), .B(n1099), .ZN(n1097) );
NOR2_X1 U797 ( .A1(n1100), .A2(n1093), .ZN(n1098) );
XNOR2_X1 U798 ( .A(G478), .B(KEYINPUT19), .ZN(n1100) );
NOR2_X1 U799 ( .A1(n1088), .A2(n1101), .ZN(G60) );
XOR2_X1 U800 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U801 ( .A1(n1104), .A2(n1093), .ZN(n1102) );
XNOR2_X1 U802 ( .A(G104), .B(n1105), .ZN(G6) );
NOR2_X1 U803 ( .A1(n1088), .A2(n1106), .ZN(G57) );
XOR2_X1 U804 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U805 ( .A(n1109), .B(n1110), .Z(n1107) );
NOR2_X1 U806 ( .A1(n1050), .A2(n1093), .ZN(n1110) );
INV_X1 U807 ( .A(G472), .ZN(n1050) );
NOR2_X1 U808 ( .A1(n1088), .A2(n1111), .ZN(G54) );
XOR2_X1 U809 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U810 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U811 ( .A(n1116), .B(n1117), .Z(n1112) );
NOR2_X1 U812 ( .A1(n1118), .A2(n1093), .ZN(n1117) );
NAND2_X1 U813 ( .A1(G902), .A2(n1006), .ZN(n1093) );
INV_X1 U814 ( .A(n1096), .ZN(n1006) );
XOR2_X1 U815 ( .A(n1119), .B(KEYINPUT59), .Z(n1116) );
NAND2_X1 U816 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U817 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
OR2_X1 U818 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U819 ( .A(KEYINPUT11), .B(n1126), .Z(n1120) );
NOR3_X1 U820 ( .A1(n1124), .A2(n1122), .A3(n1125), .ZN(n1126) );
AND3_X1 U821 ( .A1(G140), .A2(n1127), .A3(KEYINPUT25), .ZN(n1125) );
NOR2_X1 U822 ( .A1(n1128), .A2(KEYINPUT25), .ZN(n1124) );
NOR2_X1 U823 ( .A1(n1088), .A2(n1129), .ZN(G51) );
XOR2_X1 U824 ( .A(n1130), .B(n1131), .Z(n1129) );
XNOR2_X1 U825 ( .A(n1132), .B(n1133), .ZN(n1131) );
NAND2_X1 U826 ( .A1(KEYINPUT33), .A2(n1134), .ZN(n1132) );
XOR2_X1 U827 ( .A(n1135), .B(n1136), .Z(n1130) );
XNOR2_X1 U828 ( .A(G125), .B(n1137), .ZN(n1136) );
NAND3_X1 U829 ( .A1(G902), .A2(G210), .A3(n1138), .ZN(n1135) );
XNOR2_X1 U830 ( .A(n1096), .B(KEYINPUT31), .ZN(n1138) );
NOR2_X1 U831 ( .A1(n1086), .A2(n1061), .ZN(n1096) );
NAND4_X1 U832 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1061) );
NOR4_X1 U833 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1142) );
NOR2_X1 U834 ( .A1(n1147), .A2(n1148), .ZN(n1141) );
NOR3_X1 U835 ( .A1(n1149), .A2(n1035), .A3(n1044), .ZN(n1148) );
INV_X1 U836 ( .A(n1150), .ZN(n1147) );
NAND2_X1 U837 ( .A1(n1151), .A2(n1152), .ZN(n1140) );
NAND2_X1 U838 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND4_X1 U839 ( .A1(n1037), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1154) );
NOR2_X1 U840 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
OR2_X1 U841 ( .A1(n1149), .A2(n1160), .ZN(n1153) );
OR2_X1 U842 ( .A1(n1155), .A2(n1161), .ZN(n1139) );
INV_X1 U843 ( .A(KEYINPUT50), .ZN(n1155) );
NAND2_X1 U844 ( .A1(n1162), .A2(n1163), .ZN(n1086) );
AND4_X1 U845 ( .A1(n1001), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1163) );
NAND3_X1 U846 ( .A1(n1015), .A2(n1023), .A3(n1167), .ZN(n1001) );
AND4_X1 U847 ( .A1(n1168), .A2(n1169), .A3(n1105), .A4(n1170), .ZN(n1162) );
NAND3_X1 U848 ( .A1(n1171), .A2(n1015), .A3(n1172), .ZN(n1170) );
NAND3_X1 U849 ( .A1(n1167), .A2(n1015), .A3(n1022), .ZN(n1105) );
NOR2_X1 U850 ( .A1(n1008), .A2(G952), .ZN(n1088) );
XOR2_X1 U851 ( .A(G146), .B(n1173), .Z(G48) );
NOR4_X1 U852 ( .A1(KEYINPUT42), .A2(n1160), .A3(n1026), .A4(n1149), .ZN(n1173) );
INV_X1 U853 ( .A(n1151), .ZN(n1026) );
INV_X1 U854 ( .A(n1174), .ZN(n1160) );
XOR2_X1 U855 ( .A(n1161), .B(n1175), .Z(G45) );
NAND2_X1 U856 ( .A1(KEYINPUT49), .A2(G143), .ZN(n1175) );
NAND3_X1 U857 ( .A1(n1171), .A2(n1156), .A3(n1176), .ZN(n1161) );
XOR2_X1 U858 ( .A(G140), .B(n1146), .Z(G42) );
AND3_X1 U859 ( .A1(n1022), .A2(n1177), .A3(n1178), .ZN(n1146) );
XOR2_X1 U860 ( .A(n1145), .B(n1179), .Z(G39) );
XNOR2_X1 U861 ( .A(KEYINPUT14), .B(n1071), .ZN(n1179) );
AND3_X1 U862 ( .A1(n1024), .A2(n1174), .A3(n1178), .ZN(n1145) );
XOR2_X1 U863 ( .A(G134), .B(n1144), .Z(G36) );
AND3_X1 U864 ( .A1(n1156), .A2(n1023), .A3(n1178), .ZN(n1144) );
XOR2_X1 U865 ( .A(G131), .B(n1143), .Z(G33) );
AND3_X1 U866 ( .A1(n1022), .A2(n1156), .A3(n1178), .ZN(n1143) );
AND4_X1 U867 ( .A1(n1014), .A2(n1151), .A3(n1159), .A4(n1017), .ZN(n1178) );
XNOR2_X1 U868 ( .A(G128), .B(n1150), .ZN(G30) );
NAND3_X1 U869 ( .A1(n1023), .A2(n1174), .A3(n1176), .ZN(n1150) );
AND3_X1 U870 ( .A1(n1151), .A2(n1159), .A3(n1037), .ZN(n1176) );
XNOR2_X1 U871 ( .A(G101), .B(n1169), .ZN(G3) );
NAND3_X1 U872 ( .A1(n1024), .A2(n1167), .A3(n1156), .ZN(n1169) );
XOR2_X1 U873 ( .A(n1180), .B(n1181), .Z(G27) );
NOR3_X1 U874 ( .A1(n1149), .A2(n1035), .A3(n1182), .ZN(n1181) );
XNOR2_X1 U875 ( .A(n1020), .B(KEYINPUT12), .ZN(n1182) );
INV_X1 U876 ( .A(n1177), .ZN(n1035) );
NAND3_X1 U877 ( .A1(n1037), .A2(n1159), .A3(n1022), .ZN(n1149) );
NAND2_X1 U878 ( .A1(n1038), .A2(n1183), .ZN(n1159) );
NAND4_X1 U879 ( .A1(G953), .A2(G902), .A3(n1184), .A4(n1185), .ZN(n1183) );
XOR2_X1 U880 ( .A(KEYINPUT0), .B(G900), .Z(n1184) );
XNOR2_X1 U881 ( .A(G125), .B(KEYINPUT10), .ZN(n1180) );
XOR2_X1 U882 ( .A(n1186), .B(n1187), .Z(G24) );
XNOR2_X1 U883 ( .A(KEYINPUT37), .B(n1188), .ZN(n1187) );
NAND4_X1 U884 ( .A1(n1171), .A2(n1020), .A3(n1189), .A4(n1015), .ZN(n1186) );
NOR2_X1 U885 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
INV_X1 U886 ( .A(n1037), .ZN(n1191) );
XOR2_X1 U887 ( .A(n1192), .B(KEYINPUT36), .Z(n1190) );
INV_X1 U888 ( .A(n1158), .ZN(n1171) );
NAND2_X1 U889 ( .A1(n1193), .A2(n1194), .ZN(n1158) );
XOR2_X1 U890 ( .A(n1168), .B(n1195), .Z(G21) );
NAND2_X1 U891 ( .A1(KEYINPUT15), .A2(G119), .ZN(n1195) );
NAND3_X1 U892 ( .A1(n1024), .A2(n1174), .A3(n1172), .ZN(n1168) );
NAND2_X1 U893 ( .A1(n1196), .A2(n1197), .ZN(n1174) );
NAND3_X1 U894 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1197) );
INV_X1 U895 ( .A(KEYINPUT32), .ZN(n1200) );
NAND2_X1 U896 ( .A1(KEYINPUT32), .A2(n1156), .ZN(n1196) );
XNOR2_X1 U897 ( .A(G116), .B(n1166), .ZN(G18) );
NAND3_X1 U898 ( .A1(n1156), .A2(n1023), .A3(n1172), .ZN(n1166) );
NOR2_X1 U899 ( .A1(n1194), .A2(n1201), .ZN(n1023) );
XNOR2_X1 U900 ( .A(G113), .B(n1165), .ZN(G15) );
NAND3_X1 U901 ( .A1(n1022), .A2(n1156), .A3(n1172), .ZN(n1165) );
AND3_X1 U902 ( .A1(n1037), .A2(n1192), .A3(n1020), .ZN(n1172) );
INV_X1 U903 ( .A(n1044), .ZN(n1020) );
NAND2_X1 U904 ( .A1(n1029), .A2(n1202), .ZN(n1044) );
INV_X1 U905 ( .A(n1036), .ZN(n1156) );
NAND2_X1 U906 ( .A1(n1203), .A2(n1198), .ZN(n1036) );
AND2_X1 U907 ( .A1(n1201), .A2(n1194), .ZN(n1022) );
INV_X1 U908 ( .A(n1193), .ZN(n1201) );
XNOR2_X1 U909 ( .A(G110), .B(n1164), .ZN(G12) );
NAND3_X1 U910 ( .A1(n1167), .A2(n1177), .A3(n1024), .ZN(n1164) );
NOR2_X1 U911 ( .A1(n1193), .A2(n1194), .ZN(n1024) );
XOR2_X1 U912 ( .A(n1204), .B(n1104), .Z(n1194) );
INV_X1 U913 ( .A(G475), .ZN(n1104) );
OR2_X1 U914 ( .A1(n1103), .A2(G902), .ZN(n1204) );
XNOR2_X1 U915 ( .A(n1205), .B(n1206), .ZN(n1103) );
XOR2_X1 U916 ( .A(n1207), .B(n1208), .Z(n1206) );
XNOR2_X1 U917 ( .A(n1209), .B(G104), .ZN(n1208) );
INV_X1 U918 ( .A(G113), .ZN(n1209) );
XOR2_X1 U919 ( .A(n1210), .B(n1211), .Z(n1205) );
XOR2_X1 U920 ( .A(n1212), .B(n1213), .Z(n1211) );
NAND3_X1 U921 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1213) );
NAND2_X1 U922 ( .A1(KEYINPUT22), .A2(n1217), .ZN(n1216) );
OR3_X1 U923 ( .A1(n1217), .A2(KEYINPUT22), .A3(n1218), .ZN(n1215) );
NAND2_X1 U924 ( .A1(n1218), .A2(n1219), .ZN(n1214) );
NAND2_X1 U925 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
INV_X1 U926 ( .A(KEYINPUT22), .ZN(n1221) );
XNOR2_X1 U927 ( .A(KEYINPUT18), .B(n1217), .ZN(n1220) );
XOR2_X1 U928 ( .A(G140), .B(KEYINPUT61), .Z(n1218) );
NAND2_X1 U929 ( .A1(n1222), .A2(G214), .ZN(n1212) );
XOR2_X1 U930 ( .A(n1223), .B(n1224), .Z(n1210) );
NOR2_X1 U931 ( .A1(G131), .A2(KEYINPUT41), .ZN(n1224) );
NAND2_X1 U932 ( .A1(KEYINPUT43), .A2(n1188), .ZN(n1223) );
XNOR2_X1 U933 ( .A(n1225), .B(G478), .ZN(n1193) );
NAND2_X1 U934 ( .A1(n1099), .A2(n1226), .ZN(n1225) );
XNOR2_X1 U935 ( .A(KEYINPUT57), .B(n1227), .ZN(n1226) );
XOR2_X1 U936 ( .A(n1228), .B(n1229), .Z(n1099) );
XNOR2_X1 U937 ( .A(n1230), .B(n1231), .ZN(n1229) );
XOR2_X1 U938 ( .A(n1232), .B(n1233), .Z(n1231) );
AND3_X1 U939 ( .A1(G217), .A2(n1008), .A3(G234), .ZN(n1233) );
NAND2_X1 U940 ( .A1(KEYINPUT52), .A2(G116), .ZN(n1232) );
XOR2_X1 U941 ( .A(n1234), .B(n1235), .Z(n1228) );
XOR2_X1 U942 ( .A(G143), .B(G134), .Z(n1235) );
XNOR2_X1 U943 ( .A(G122), .B(G128), .ZN(n1234) );
NAND2_X1 U944 ( .A1(n1236), .A2(n1237), .ZN(n1177) );
OR3_X1 U945 ( .A1(n1198), .A2(n1203), .A3(KEYINPUT32), .ZN(n1237) );
NAND2_X1 U946 ( .A1(KEYINPUT32), .A2(n1015), .ZN(n1236) );
NOR2_X1 U947 ( .A1(n1198), .A2(n1199), .ZN(n1015) );
INV_X1 U948 ( .A(n1203), .ZN(n1199) );
XOR2_X1 U949 ( .A(n1238), .B(n1239), .Z(n1203) );
INV_X1 U950 ( .A(n1053), .ZN(n1239) );
NOR2_X1 U951 ( .A1(n1095), .A2(G902), .ZN(n1053) );
INV_X1 U952 ( .A(n1092), .ZN(n1095) );
XNOR2_X1 U953 ( .A(n1240), .B(n1241), .ZN(n1092) );
XOR2_X1 U954 ( .A(n1242), .B(n1243), .Z(n1241) );
XNOR2_X1 U955 ( .A(G146), .B(n1244), .ZN(n1243) );
XOR2_X1 U956 ( .A(KEYINPUT60), .B(KEYINPUT2), .Z(n1242) );
XOR2_X1 U957 ( .A(n1245), .B(n1246), .Z(n1240) );
XNOR2_X1 U958 ( .A(n1217), .B(G119), .ZN(n1246) );
XOR2_X1 U959 ( .A(n1247), .B(n1128), .Z(n1245) );
XOR2_X1 U960 ( .A(G110), .B(G140), .Z(n1128) );
NAND2_X1 U961 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND4_X1 U962 ( .A1(G221), .A2(G234), .A3(n1250), .A4(n1008), .ZN(n1249) );
NAND2_X1 U963 ( .A1(n1251), .A2(n1252), .ZN(n1248) );
NAND3_X1 U964 ( .A1(G234), .A2(n1008), .A3(G221), .ZN(n1252) );
XOR2_X1 U965 ( .A(KEYINPUT47), .B(n1250), .Z(n1251) );
XNOR2_X1 U966 ( .A(n1071), .B(KEYINPUT4), .ZN(n1250) );
NAND2_X1 U967 ( .A1(KEYINPUT13), .A2(n1052), .ZN(n1238) );
NAND2_X1 U968 ( .A1(G217), .A2(n1253), .ZN(n1052) );
XNOR2_X1 U969 ( .A(n1049), .B(G472), .ZN(n1198) );
NAND3_X1 U970 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1049) );
XNOR2_X1 U971 ( .A(G902), .B(KEYINPUT5), .ZN(n1256) );
NAND3_X1 U972 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1255) );
INV_X1 U973 ( .A(KEYINPUT21), .ZN(n1259) );
XNOR2_X1 U974 ( .A(G101), .B(n1260), .ZN(n1258) );
XOR2_X1 U975 ( .A(n1261), .B(n1262), .Z(n1257) );
NAND2_X1 U976 ( .A1(n1263), .A2(KEYINPUT21), .ZN(n1254) );
XNOR2_X1 U977 ( .A(n1261), .B(n1108), .ZN(n1263) );
XNOR2_X1 U978 ( .A(n1114), .B(n1260), .ZN(n1108) );
NAND2_X1 U979 ( .A1(n1222), .A2(G210), .ZN(n1260) );
NOR2_X1 U980 ( .A1(G953), .A2(G237), .ZN(n1222) );
XOR2_X1 U981 ( .A(n1262), .B(n1264), .Z(n1114) );
XOR2_X1 U982 ( .A(n1109), .B(KEYINPUT38), .Z(n1261) );
XNOR2_X1 U983 ( .A(n1133), .B(n1265), .ZN(n1109) );
XNOR2_X1 U984 ( .A(G113), .B(n1266), .ZN(n1265) );
NAND2_X1 U985 ( .A1(KEYINPUT24), .A2(n1267), .ZN(n1266) );
XNOR2_X1 U986 ( .A(n1268), .B(G116), .ZN(n1267) );
AND3_X1 U987 ( .A1(n1151), .A2(n1192), .A3(n1037), .ZN(n1167) );
NOR2_X1 U988 ( .A1(n1014), .A2(n1045), .ZN(n1037) );
INV_X1 U989 ( .A(n1017), .ZN(n1045) );
NAND2_X1 U990 ( .A1(G214), .A2(n1269), .ZN(n1017) );
INV_X1 U991 ( .A(n1054), .ZN(n1014) );
XNOR2_X1 U992 ( .A(n1270), .B(n1271), .ZN(n1054) );
NOR2_X1 U993 ( .A1(G902), .A2(n1272), .ZN(n1271) );
XNOR2_X1 U994 ( .A(n1134), .B(n1273), .ZN(n1272) );
XOR2_X1 U995 ( .A(n1274), .B(n1275), .Z(n1273) );
NOR2_X1 U996 ( .A1(KEYINPUT48), .A2(n1137), .ZN(n1275) );
NAND2_X1 U997 ( .A1(G224), .A2(n1008), .ZN(n1137) );
NAND2_X1 U998 ( .A1(n1276), .A2(n1277), .ZN(n1274) );
NAND2_X1 U999 ( .A1(G125), .A2(n1278), .ZN(n1277) );
INV_X1 U1000 ( .A(n1133), .ZN(n1278) );
XOR2_X1 U1001 ( .A(n1279), .B(KEYINPUT26), .Z(n1276) );
NAND2_X1 U1002 ( .A1(n1133), .A2(n1217), .ZN(n1279) );
INV_X1 U1003 ( .A(G125), .ZN(n1217) );
XOR2_X1 U1004 ( .A(G128), .B(n1207), .Z(n1133) );
XNOR2_X1 U1005 ( .A(n1077), .B(n1280), .ZN(n1134) );
NOR2_X1 U1006 ( .A1(KEYINPUT23), .A2(n1281), .ZN(n1280) );
XOR2_X1 U1007 ( .A(n1082), .B(n1081), .Z(n1281) );
XOR2_X1 U1008 ( .A(n1282), .B(G101), .Z(n1081) );
XOR2_X1 U1009 ( .A(n1283), .B(n1284), .Z(n1082) );
NOR2_X1 U1010 ( .A1(G113), .A2(KEYINPUT28), .ZN(n1284) );
NAND3_X1 U1011 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(n1283) );
NAND2_X1 U1012 ( .A1(G116), .A2(n1268), .ZN(n1287) );
INV_X1 U1013 ( .A(G119), .ZN(n1268) );
NAND2_X1 U1014 ( .A1(n1288), .A2(n1289), .ZN(n1286) );
INV_X1 U1015 ( .A(KEYINPUT6), .ZN(n1289) );
NAND2_X1 U1016 ( .A1(n1290), .A2(n1291), .ZN(n1288) );
XNOR2_X1 U1017 ( .A(KEYINPUT53), .B(G119), .ZN(n1290) );
NAND2_X1 U1018 ( .A1(KEYINPUT6), .A2(n1292), .ZN(n1285) );
NAND2_X1 U1019 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
OR2_X1 U1020 ( .A1(G119), .A2(KEYINPUT53), .ZN(n1294) );
NAND3_X1 U1021 ( .A1(G119), .A2(n1291), .A3(KEYINPUT53), .ZN(n1293) );
INV_X1 U1022 ( .A(G116), .ZN(n1291) );
XNOR2_X1 U1023 ( .A(n1295), .B(n1188), .ZN(n1077) );
INV_X1 U1024 ( .A(G122), .ZN(n1188) );
NAND2_X1 U1025 ( .A1(KEYINPUT34), .A2(n1127), .ZN(n1295) );
INV_X1 U1026 ( .A(G110), .ZN(n1127) );
NAND2_X1 U1027 ( .A1(n1296), .A2(n1269), .ZN(n1270) );
NAND2_X1 U1028 ( .A1(n1297), .A2(n1227), .ZN(n1269) );
INV_X1 U1029 ( .A(G237), .ZN(n1297) );
XNOR2_X1 U1030 ( .A(G210), .B(KEYINPUT63), .ZN(n1296) );
NAND2_X1 U1031 ( .A1(n1038), .A2(n1298), .ZN(n1192) );
NAND4_X1 U1032 ( .A1(G953), .A2(G902), .A3(n1185), .A4(n1299), .ZN(n1298) );
INV_X1 U1033 ( .A(G898), .ZN(n1299) );
NAND3_X1 U1034 ( .A1(n1185), .A2(n1008), .A3(G952), .ZN(n1038) );
NAND2_X1 U1035 ( .A1(G237), .A2(G234), .ZN(n1185) );
NOR2_X1 U1036 ( .A1(n1029), .A2(n1028), .ZN(n1151) );
INV_X1 U1037 ( .A(n1202), .ZN(n1028) );
NAND2_X1 U1038 ( .A1(G221), .A2(n1253), .ZN(n1202) );
NAND2_X1 U1039 ( .A1(G234), .A2(n1227), .ZN(n1253) );
XNOR2_X1 U1040 ( .A(n1300), .B(n1118), .ZN(n1029) );
INV_X1 U1041 ( .A(G469), .ZN(n1118) );
NAND2_X1 U1042 ( .A1(n1301), .A2(n1227), .ZN(n1300) );
INV_X1 U1043 ( .A(G902), .ZN(n1227) );
XOR2_X1 U1044 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U1045 ( .A(n1122), .B(n1115), .Z(n1303) );
XNOR2_X1 U1046 ( .A(n1304), .B(n1066), .ZN(n1115) );
XNOR2_X1 U1047 ( .A(n1305), .B(n1207), .ZN(n1066) );
XOR2_X1 U1048 ( .A(G146), .B(G143), .Z(n1207) );
NAND2_X1 U1049 ( .A1(n1306), .A2(n1244), .ZN(n1305) );
INV_X1 U1050 ( .A(G128), .ZN(n1244) );
XOR2_X1 U1051 ( .A(KEYINPUT39), .B(KEYINPUT3), .Z(n1306) );
XNOR2_X1 U1052 ( .A(KEYINPUT9), .B(n1307), .ZN(n1304) );
NOR2_X1 U1053 ( .A1(KEYINPUT35), .A2(n1282), .ZN(n1307) );
XOR2_X1 U1054 ( .A(G104), .B(n1230), .Z(n1282) );
XOR2_X1 U1055 ( .A(G107), .B(KEYINPUT1), .Z(n1230) );
AND2_X1 U1056 ( .A1(G227), .A2(n1008), .ZN(n1122) );
INV_X1 U1057 ( .A(G953), .ZN(n1008) );
XOR2_X1 U1058 ( .A(n1308), .B(n1309), .Z(n1302) );
XNOR2_X1 U1059 ( .A(n1264), .B(n1310), .ZN(n1309) );
NOR2_X1 U1060 ( .A1(KEYINPUT56), .A2(n1311), .ZN(n1310) );
XOR2_X1 U1061 ( .A(n1312), .B(n1313), .Z(n1311) );
NOR2_X1 U1062 ( .A1(G110), .A2(KEYINPUT51), .ZN(n1313) );
XNOR2_X1 U1063 ( .A(G140), .B(KEYINPUT20), .ZN(n1312) );
INV_X1 U1064 ( .A(G101), .ZN(n1264) );
NOR2_X1 U1065 ( .A1(KEYINPUT29), .A2(n1262), .ZN(n1308) );
XOR2_X1 U1066 ( .A(n1314), .B(n1315), .Z(n1262) );
XOR2_X1 U1067 ( .A(KEYINPUT45), .B(G131), .Z(n1315) );
NAND3_X1 U1068 ( .A1(n1316), .A2(n1317), .A3(n1318), .ZN(n1314) );
NAND2_X1 U1069 ( .A1(KEYINPUT55), .A2(G134), .ZN(n1318) );
OR3_X1 U1070 ( .A1(G134), .A2(KEYINPUT55), .A3(n1071), .ZN(n1317) );
NAND2_X1 U1071 ( .A1(n1319), .A2(n1071), .ZN(n1316) );
INV_X1 U1072 ( .A(G137), .ZN(n1071) );
NAND2_X1 U1073 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
INV_X1 U1074 ( .A(KEYINPUT55), .ZN(n1321) );
XNOR2_X1 U1075 ( .A(G134), .B(KEYINPUT62), .ZN(n1320) );
endmodule


