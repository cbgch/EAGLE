//Key = 1101101011010110010011111010110010111010100000010000100110001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;

XOR2_X1 U731 ( .A(G107), .B(n1006), .Z(G9) );
NOR2_X1 U732 ( .A1(n1007), .A2(n1008), .ZN(G75) );
NOR4_X1 U733 ( .A1(n1009), .A2(n1010), .A3(n1011), .A4(n1012), .ZN(n1008) );
INV_X1 U734 ( .A(G952), .ZN(n1012) );
NOR3_X1 U735 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1011) );
INV_X1 U736 ( .A(n1016), .ZN(n1014) );
NAND3_X1 U737 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1013) );
NAND2_X1 U738 ( .A1(n1020), .A2(n1021), .ZN(n1017) );
INV_X1 U739 ( .A(n1022), .ZN(n1021) );
NAND3_X1 U740 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1020) );
NAND2_X1 U741 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NAND3_X1 U742 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1023) );
NAND3_X1 U743 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1009) );
NAND4_X1 U744 ( .A1(n1034), .A2(n1030), .A3(n1016), .A4(n1035), .ZN(n1033) );
NOR2_X1 U745 ( .A1(n1027), .A2(n1036), .ZN(n1035) );
XNOR2_X1 U746 ( .A(n1037), .B(KEYINPUT52), .ZN(n1016) );
NAND2_X1 U747 ( .A1(n1038), .A2(n1039), .ZN(n1034) );
NAND3_X1 U748 ( .A1(n1040), .A2(n1041), .A3(n1019), .ZN(n1039) );
NAND2_X1 U749 ( .A1(n1042), .A2(n1015), .ZN(n1041) );
NAND3_X1 U750 ( .A1(n1043), .A2(n1044), .A3(n1018), .ZN(n1040) );
NAND2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1038) );
NOR3_X1 U752 ( .A1(n1047), .A2(G953), .A3(n1048), .ZN(n1007) );
INV_X1 U753 ( .A(n1031), .ZN(n1048) );
NAND4_X1 U754 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1031) );
NOR4_X1 U755 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
XNOR2_X1 U756 ( .A(KEYINPUT18), .B(n1057), .ZN(n1056) );
XNOR2_X1 U757 ( .A(n1036), .B(KEYINPUT3), .ZN(n1053) );
NOR3_X1 U758 ( .A1(n1042), .A2(n1058), .A3(n1026), .ZN(n1051) );
NAND2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1050) );
XNOR2_X1 U760 ( .A(KEYINPUT46), .B(n1061), .ZN(n1059) );
XNOR2_X1 U761 ( .A(n1062), .B(n1063), .ZN(n1049) );
NOR2_X1 U762 ( .A1(KEYINPUT44), .A2(n1064), .ZN(n1063) );
XNOR2_X1 U763 ( .A(G952), .B(KEYINPUT32), .ZN(n1047) );
XOR2_X1 U764 ( .A(n1065), .B(n1066), .Z(G72) );
XOR2_X1 U765 ( .A(n1067), .B(n1068), .Z(n1066) );
NOR2_X1 U766 ( .A1(n1069), .A2(n1032), .ZN(n1068) );
AND2_X1 U767 ( .A1(G227), .A2(G900), .ZN(n1069) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1067) );
NAND2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U770 ( .A(n1074), .B(n1075), .Z(n1070) );
NAND2_X1 U771 ( .A1(KEYINPUT29), .A2(n1076), .ZN(n1075) );
NAND3_X1 U772 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1074) );
OR2_X1 U773 ( .A1(n1080), .A2(KEYINPUT39), .ZN(n1078) );
NAND2_X1 U774 ( .A1(KEYINPUT39), .A2(G140), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1032), .A2(n1081), .ZN(n1065) );
XOR2_X1 U776 ( .A(n1082), .B(n1083), .Z(G69) );
NOR2_X1 U777 ( .A1(n1084), .A2(n1032), .ZN(n1083) );
NOR2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U779 ( .A1(KEYINPUT31), .A2(n1087), .ZN(n1082) );
XOR2_X1 U780 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR3_X1 U781 ( .A1(n1090), .A2(KEYINPUT43), .A3(n1091), .ZN(n1089) );
NOR2_X1 U782 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U783 ( .A(KEYINPUT12), .B(n1032), .ZN(n1090) );
NAND2_X1 U784 ( .A1(n1094), .A2(n1095), .ZN(n1088) );
NAND2_X1 U785 ( .A1(n1072), .A2(n1086), .ZN(n1095) );
XNOR2_X1 U786 ( .A(n1096), .B(n1097), .ZN(n1094) );
NAND2_X1 U787 ( .A1(KEYINPUT38), .A2(n1098), .ZN(n1096) );
NOR2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(G66) );
XNOR2_X1 U789 ( .A(n1101), .B(n1102), .ZN(n1100) );
NOR2_X1 U790 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U791 ( .A1(n1099), .A2(n1105), .ZN(G63) );
XOR2_X1 U792 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U793 ( .A1(n1108), .A2(n1104), .ZN(n1106) );
NOR2_X1 U794 ( .A1(n1099), .A2(n1109), .ZN(G60) );
XOR2_X1 U795 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U796 ( .A1(n1061), .A2(n1104), .ZN(n1110) );
INV_X1 U797 ( .A(G475), .ZN(n1061) );
XNOR2_X1 U798 ( .A(G104), .B(n1112), .ZN(G6) );
NOR2_X1 U799 ( .A1(n1113), .A2(n1114), .ZN(G57) );
XOR2_X1 U800 ( .A(KEYINPUT51), .B(n1099), .Z(n1114) );
XOR2_X1 U801 ( .A(n1115), .B(n1116), .Z(n1113) );
XOR2_X1 U802 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U803 ( .A1(KEYINPUT35), .A2(n1119), .ZN(n1117) );
XOR2_X1 U804 ( .A(G101), .B(n1120), .Z(n1115) );
NOR2_X1 U805 ( .A1(n1121), .A2(n1104), .ZN(n1120) );
NOR2_X1 U806 ( .A1(n1099), .A2(n1122), .ZN(G54) );
XOR2_X1 U807 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U808 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND2_X1 U809 ( .A1(n1127), .A2(KEYINPUT56), .ZN(n1126) );
XNOR2_X1 U810 ( .A(n1128), .B(n1076), .ZN(n1127) );
NAND2_X1 U811 ( .A1(KEYINPUT26), .A2(n1129), .ZN(n1128) );
NAND2_X1 U812 ( .A1(n1130), .A2(n1131), .ZN(n1125) );
NAND2_X1 U813 ( .A1(G110), .A2(n1132), .ZN(n1131) );
NAND2_X1 U814 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U815 ( .A1(G140), .A2(n1135), .ZN(n1134) );
NAND2_X1 U816 ( .A1(n1136), .A2(n1137), .ZN(n1130) );
NAND2_X1 U817 ( .A1(n1135), .A2(n1138), .ZN(n1136) );
NAND2_X1 U818 ( .A1(n1139), .A2(n1133), .ZN(n1138) );
INV_X1 U819 ( .A(KEYINPUT10), .ZN(n1133) );
INV_X1 U820 ( .A(KEYINPUT16), .ZN(n1135) );
XOR2_X1 U821 ( .A(n1140), .B(n1141), .Z(n1123) );
NOR2_X1 U822 ( .A1(n1142), .A2(n1104), .ZN(n1141) );
NOR2_X1 U823 ( .A1(n1099), .A2(n1143), .ZN(G51) );
XOR2_X1 U824 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U825 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U826 ( .A1(n1148), .A2(n1104), .ZN(n1146) );
NAND2_X1 U827 ( .A1(G902), .A2(n1010), .ZN(n1104) );
OR3_X1 U828 ( .A1(n1093), .A2(n1149), .A3(n1081), .ZN(n1010) );
NAND4_X1 U829 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1081) );
NOR4_X1 U830 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1153) );
NAND2_X1 U831 ( .A1(n1158), .A2(n1046), .ZN(n1152) );
XOR2_X1 U832 ( .A(n1159), .B(KEYINPUT40), .Z(n1158) );
OR2_X1 U833 ( .A1(n1160), .A2(n1044), .ZN(n1159) );
NAND2_X1 U834 ( .A1(n1161), .A2(n1162), .ZN(n1150) );
NAND2_X1 U835 ( .A1(n1028), .A2(n1029), .ZN(n1162) );
INV_X1 U836 ( .A(n1163), .ZN(n1161) );
XNOR2_X1 U837 ( .A(KEYINPUT6), .B(n1092), .ZN(n1149) );
NAND4_X1 U838 ( .A1(n1164), .A2(n1112), .A3(n1165), .A4(n1166), .ZN(n1093) );
NOR4_X1 U839 ( .A1(n1006), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1166) );
NOR2_X1 U840 ( .A1(n1029), .A2(n1170), .ZN(n1006) );
OR3_X1 U841 ( .A1(n1043), .A2(n1028), .A3(n1171), .ZN(n1165) );
OR2_X1 U842 ( .A1(n1028), .A2(n1170), .ZN(n1112) );
NAND3_X1 U843 ( .A1(n1172), .A2(n1173), .A3(n1045), .ZN(n1170) );
NAND4_X1 U844 ( .A1(n1022), .A2(n1174), .A3(n1175), .A4(n1173), .ZN(n1164) );
XNOR2_X1 U845 ( .A(KEYINPUT42), .B(n1176), .ZN(n1175) );
INV_X1 U846 ( .A(n1044), .ZN(n1174) );
XOR2_X1 U847 ( .A(n1177), .B(KEYINPUT9), .Z(n1144) );
NAND2_X1 U848 ( .A1(n1178), .A2(KEYINPUT60), .ZN(n1177) );
XNOR2_X1 U849 ( .A(n1179), .B(n1180), .ZN(n1178) );
XOR2_X1 U850 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U851 ( .A1(G125), .A2(KEYINPUT2), .ZN(n1182) );
NOR2_X1 U852 ( .A1(n1032), .A2(G952), .ZN(n1099) );
XNOR2_X1 U853 ( .A(n1183), .B(n1184), .ZN(G48) );
NOR2_X1 U854 ( .A1(n1028), .A2(n1163), .ZN(n1184) );
XNOR2_X1 U855 ( .A(G143), .B(n1151), .ZN(G45) );
NAND3_X1 U856 ( .A1(n1185), .A2(n1172), .A3(n1186), .ZN(n1151) );
NOR3_X1 U857 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1186) );
NAND3_X1 U858 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(G42) );
NAND2_X1 U859 ( .A1(n1157), .A2(n1137), .ZN(n1192) );
NAND2_X1 U860 ( .A1(n1193), .A2(n1194), .ZN(n1191) );
INV_X1 U861 ( .A(KEYINPUT4), .ZN(n1194) );
NAND2_X1 U862 ( .A1(n1195), .A2(n1196), .ZN(n1193) );
XNOR2_X1 U863 ( .A(KEYINPUT36), .B(G140), .ZN(n1195) );
NAND2_X1 U864 ( .A1(KEYINPUT4), .A2(n1197), .ZN(n1190) );
NAND2_X1 U865 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
OR2_X1 U866 ( .A1(G140), .A2(KEYINPUT36), .ZN(n1199) );
NAND3_X1 U867 ( .A1(G140), .A2(n1196), .A3(KEYINPUT36), .ZN(n1198) );
INV_X1 U868 ( .A(n1157), .ZN(n1196) );
NOR3_X1 U869 ( .A1(n1200), .A2(n1028), .A3(n1044), .ZN(n1157) );
XOR2_X1 U870 ( .A(G137), .B(n1155), .Z(G39) );
NOR3_X1 U871 ( .A1(n1201), .A2(n1200), .A3(n1027), .ZN(n1155) );
XNOR2_X1 U872 ( .A(G134), .B(n1202), .ZN(G36) );
NAND2_X1 U873 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NAND2_X1 U874 ( .A1(KEYINPUT20), .A2(n1205), .ZN(n1204) );
INV_X1 U875 ( .A(n1156), .ZN(n1205) );
NAND2_X1 U876 ( .A1(KEYINPUT48), .A2(n1156), .ZN(n1203) );
NOR3_X1 U877 ( .A1(n1043), .A2(n1029), .A3(n1200), .ZN(n1156) );
XOR2_X1 U878 ( .A(G131), .B(n1154), .Z(G33) );
NOR3_X1 U879 ( .A1(n1043), .A2(n1028), .A3(n1200), .ZN(n1154) );
NAND3_X1 U880 ( .A1(n1036), .A2(n1019), .A3(n1206), .ZN(n1200) );
NOR3_X1 U881 ( .A1(n1189), .A2(n1026), .A3(n1042), .ZN(n1206) );
INV_X1 U882 ( .A(n1207), .ZN(n1189) );
XNOR2_X1 U883 ( .A(n1208), .B(n1209), .ZN(G30) );
NOR3_X1 U884 ( .A1(n1163), .A2(KEYINPUT54), .A3(n1029), .ZN(n1209) );
NAND3_X1 U885 ( .A1(n1172), .A2(n1207), .A3(n1210), .ZN(n1163) );
NOR3_X1 U886 ( .A1(n1025), .A2(n1026), .A3(n1176), .ZN(n1172) );
XOR2_X1 U887 ( .A(G101), .B(n1169), .Z(G3) );
NOR2_X1 U888 ( .A1(n1211), .A2(n1043), .ZN(n1169) );
XNOR2_X1 U889 ( .A(n1212), .B(n1213), .ZN(G27) );
NOR3_X1 U890 ( .A1(n1214), .A2(n1176), .A3(n1160), .ZN(n1213) );
NAND4_X1 U891 ( .A1(n1025), .A2(n1215), .A3(n1207), .A4(n1030), .ZN(n1160) );
NAND2_X1 U892 ( .A1(n1216), .A2(n1217), .ZN(n1207) );
NAND2_X1 U893 ( .A1(n1218), .A2(n1073), .ZN(n1217) );
INV_X1 U894 ( .A(G900), .ZN(n1073) );
INV_X1 U895 ( .A(n1046), .ZN(n1176) );
XNOR2_X1 U896 ( .A(KEYINPUT61), .B(n1044), .ZN(n1214) );
XOR2_X1 U897 ( .A(G122), .B(n1168), .Z(G24) );
NOR4_X1 U898 ( .A1(n1171), .A2(n1015), .A3(n1187), .A4(n1188), .ZN(n1168) );
INV_X1 U899 ( .A(n1045), .ZN(n1015) );
NOR2_X1 U900 ( .A1(n1219), .A2(n1054), .ZN(n1045) );
XNOR2_X1 U901 ( .A(n1220), .B(n1221), .ZN(G21) );
NAND2_X1 U902 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
OR4_X1 U903 ( .A1(n1027), .A2(n1210), .A3(n1171), .A4(KEYINPUT21), .ZN(n1223) );
INV_X1 U904 ( .A(n1201), .ZN(n1210) );
NAND2_X1 U905 ( .A1(n1092), .A2(KEYINPUT21), .ZN(n1222) );
NOR3_X1 U906 ( .A1(n1027), .A2(n1201), .A3(n1171), .ZN(n1092) );
NAND2_X1 U907 ( .A1(n1054), .A2(n1219), .ZN(n1201) );
XNOR2_X1 U908 ( .A(n1224), .B(n1167), .ZN(G18) );
NOR3_X1 U909 ( .A1(n1043), .A2(n1029), .A3(n1171), .ZN(n1167) );
NAND2_X1 U910 ( .A1(n1188), .A2(n1225), .ZN(n1029) );
XNOR2_X1 U911 ( .A(n1226), .B(n1227), .ZN(G15) );
NOR4_X1 U912 ( .A1(KEYINPUT30), .A2(n1028), .A3(n1043), .A4(n1171), .ZN(n1227) );
NAND4_X1 U913 ( .A1(n1025), .A2(n1046), .A3(n1030), .A4(n1173), .ZN(n1171) );
INV_X1 U914 ( .A(n1185), .ZN(n1043) );
NOR2_X1 U915 ( .A1(n1054), .A2(n1057), .ZN(n1185) );
INV_X1 U916 ( .A(n1215), .ZN(n1028) );
NOR2_X1 U917 ( .A1(n1225), .A2(n1188), .ZN(n1215) );
XNOR2_X1 U918 ( .A(n1139), .B(n1228), .ZN(G12) );
NOR3_X1 U919 ( .A1(n1211), .A2(KEYINPUT53), .A3(n1044), .ZN(n1228) );
NAND2_X1 U920 ( .A1(n1057), .A2(n1054), .ZN(n1044) );
XOR2_X1 U921 ( .A(n1229), .B(n1103), .Z(n1054) );
NAND2_X1 U922 ( .A1(G217), .A2(n1230), .ZN(n1103) );
NAND2_X1 U923 ( .A1(n1101), .A2(n1231), .ZN(n1229) );
XNOR2_X1 U924 ( .A(n1232), .B(n1233), .ZN(n1101) );
XOR2_X1 U925 ( .A(n1234), .B(n1235), .Z(n1233) );
XNOR2_X1 U926 ( .A(n1139), .B(n1236), .ZN(n1235) );
NOR2_X1 U927 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XOR2_X1 U928 ( .A(KEYINPUT33), .B(n1239), .Z(n1238) );
NOR2_X1 U929 ( .A1(n1183), .A2(n1240), .ZN(n1239) );
AND2_X1 U930 ( .A1(n1183), .A2(n1240), .ZN(n1237) );
NAND3_X1 U931 ( .A1(n1241), .A2(n1242), .A3(n1080), .ZN(n1240) );
INV_X1 U932 ( .A(n1243), .ZN(n1080) );
OR2_X1 U933 ( .A1(G140), .A2(KEYINPUT0), .ZN(n1242) );
NAND2_X1 U934 ( .A1(n1244), .A2(KEYINPUT0), .ZN(n1241) );
AND2_X1 U935 ( .A1(n1245), .A2(G221), .ZN(n1234) );
XOR2_X1 U936 ( .A(n1246), .B(n1247), .Z(n1232) );
XNOR2_X1 U937 ( .A(n1208), .B(G119), .ZN(n1247) );
XNOR2_X1 U938 ( .A(G137), .B(KEYINPUT49), .ZN(n1246) );
INV_X1 U939 ( .A(n1219), .ZN(n1057) );
XOR2_X1 U940 ( .A(n1248), .B(n1121), .Z(n1219) );
INV_X1 U941 ( .A(G472), .ZN(n1121) );
NAND2_X1 U942 ( .A1(n1249), .A2(n1231), .ZN(n1248) );
XOR2_X1 U943 ( .A(n1250), .B(n1251), .Z(n1249) );
XOR2_X1 U944 ( .A(n1118), .B(n1252), .Z(n1251) );
NOR2_X1 U945 ( .A1(G101), .A2(KEYINPUT19), .ZN(n1252) );
XOR2_X1 U946 ( .A(n1253), .B(n1254), .Z(n1118) );
XNOR2_X1 U947 ( .A(G128), .B(n1255), .ZN(n1254) );
NAND2_X1 U948 ( .A1(G210), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U949 ( .A(n1119), .B(KEYINPUT50), .ZN(n1250) );
AND2_X1 U950 ( .A1(n1257), .A2(n1258), .ZN(n1119) );
OR2_X1 U951 ( .A1(n1259), .A2(n1226), .ZN(n1258) );
XOR2_X1 U952 ( .A(n1260), .B(KEYINPUT5), .Z(n1257) );
NAND2_X1 U953 ( .A1(n1259), .A2(n1226), .ZN(n1260) );
XOR2_X1 U954 ( .A(G116), .B(n1261), .Z(n1259) );
XNOR2_X1 U955 ( .A(KEYINPUT11), .B(n1221), .ZN(n1261) );
NAND3_X1 U956 ( .A1(n1046), .A2(n1173), .A3(n1022), .ZN(n1211) );
NOR3_X1 U957 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1022) );
NAND2_X1 U958 ( .A1(n1187), .A2(n1188), .ZN(n1027) );
NOR2_X1 U959 ( .A1(n1262), .A2(n1058), .ZN(n1188) );
NOR2_X1 U960 ( .A1(n1060), .A2(G475), .ZN(n1058) );
AND2_X1 U961 ( .A1(G475), .A2(n1060), .ZN(n1262) );
OR2_X1 U962 ( .A1(n1111), .A2(G902), .ZN(n1060) );
XNOR2_X1 U963 ( .A(n1263), .B(n1264), .ZN(n1111) );
XOR2_X1 U964 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U965 ( .A(n1267), .B(n1268), .Z(n1266) );
NOR2_X1 U966 ( .A1(G131), .A2(KEYINPUT7), .ZN(n1268) );
NAND3_X1 U967 ( .A1(n1269), .A2(n1270), .A3(n1079), .ZN(n1267) );
INV_X1 U968 ( .A(n1244), .ZN(n1079) );
NOR2_X1 U969 ( .A1(n1137), .A2(n1212), .ZN(n1244) );
INV_X1 U970 ( .A(G140), .ZN(n1137) );
OR2_X1 U971 ( .A1(n1212), .A2(KEYINPUT22), .ZN(n1270) );
NAND2_X1 U972 ( .A1(n1243), .A2(KEYINPUT22), .ZN(n1269) );
NOR2_X1 U973 ( .A1(G125), .A2(G140), .ZN(n1243) );
NAND2_X1 U974 ( .A1(G214), .A2(n1256), .ZN(n1265) );
NOR2_X1 U975 ( .A1(G953), .A2(G237), .ZN(n1256) );
XOR2_X1 U976 ( .A(n1271), .B(n1272), .Z(n1263) );
NAND2_X1 U977 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
NAND2_X1 U978 ( .A1(G104), .A2(n1275), .ZN(n1274) );
XOR2_X1 U979 ( .A(KEYINPUT24), .B(n1276), .Z(n1273) );
NOR2_X1 U980 ( .A1(G104), .A2(n1275), .ZN(n1276) );
XNOR2_X1 U981 ( .A(G122), .B(n1226), .ZN(n1275) );
INV_X1 U982 ( .A(G113), .ZN(n1226) );
INV_X1 U983 ( .A(n1225), .ZN(n1187) );
XOR2_X1 U984 ( .A(n1277), .B(n1064), .Z(n1225) );
XOR2_X1 U985 ( .A(n1108), .B(KEYINPUT47), .Z(n1064) );
INV_X1 U986 ( .A(G478), .ZN(n1108) );
NAND2_X1 U987 ( .A1(KEYINPUT17), .A2(n1062), .ZN(n1277) );
OR2_X1 U988 ( .A1(n1278), .A2(n1107), .ZN(n1062) );
XNOR2_X1 U989 ( .A(n1279), .B(n1280), .ZN(n1107) );
XOR2_X1 U990 ( .A(n1281), .B(n1282), .Z(n1280) );
XNOR2_X1 U991 ( .A(KEYINPUT14), .B(n1283), .ZN(n1282) );
NOR2_X1 U992 ( .A1(G128), .A2(KEYINPUT37), .ZN(n1283) );
NAND2_X1 U993 ( .A1(G217), .A2(n1245), .ZN(n1281) );
AND2_X1 U994 ( .A1(G234), .A2(n1032), .ZN(n1245) );
XOR2_X1 U995 ( .A(n1284), .B(n1285), .Z(n1279) );
XOR2_X1 U996 ( .A(n1286), .B(n1287), .Z(n1284) );
XNOR2_X1 U997 ( .A(n1231), .B(KEYINPUT59), .ZN(n1278) );
INV_X1 U998 ( .A(n1030), .ZN(n1026) );
NAND2_X1 U999 ( .A1(G221), .A2(n1230), .ZN(n1030) );
NAND2_X1 U1000 ( .A1(G234), .A2(n1231), .ZN(n1230) );
INV_X1 U1001 ( .A(n1036), .ZN(n1025) );
XOR2_X1 U1002 ( .A(n1288), .B(n1142), .Z(n1036) );
INV_X1 U1003 ( .A(G469), .ZN(n1142) );
NAND2_X1 U1004 ( .A1(n1289), .A2(n1231), .ZN(n1288) );
XOR2_X1 U1005 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U1006 ( .A(n1140), .B(n1292), .Z(n1291) );
NAND2_X1 U1007 ( .A1(KEYINPUT63), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U1008 ( .A(n1076), .B(n1294), .ZN(n1293) );
XOR2_X1 U1009 ( .A(KEYINPUT58), .B(n1129), .Z(n1294) );
XNOR2_X1 U1010 ( .A(n1295), .B(G101), .ZN(n1129) );
NAND4_X1 U1011 ( .A1(KEYINPUT55), .A2(n1296), .A3(n1297), .A4(n1298), .ZN(n1295) );
OR3_X1 U1012 ( .A1(n1299), .A2(n1287), .A3(KEYINPUT45), .ZN(n1298) );
NAND2_X1 U1013 ( .A1(KEYINPUT45), .A2(n1299), .ZN(n1297) );
XNOR2_X1 U1014 ( .A(n1300), .B(n1253), .ZN(n1076) );
XOR2_X1 U1015 ( .A(n1301), .B(n1302), .Z(n1253) );
XNOR2_X1 U1016 ( .A(n1183), .B(G137), .ZN(n1302) );
XOR2_X1 U1017 ( .A(n1286), .B(G131), .Z(n1301) );
XNOR2_X1 U1018 ( .A(G134), .B(n1303), .ZN(n1286) );
XOR2_X1 U1019 ( .A(KEYINPUT23), .B(G143), .Z(n1303) );
NAND2_X1 U1020 ( .A1(KEYINPUT62), .A2(n1208), .ZN(n1300) );
INV_X1 U1021 ( .A(G128), .ZN(n1208) );
NAND2_X1 U1022 ( .A1(n1304), .A2(n1032), .ZN(n1140) );
XNOR2_X1 U1023 ( .A(G227), .B(KEYINPUT13), .ZN(n1304) );
XNOR2_X1 U1024 ( .A(G110), .B(G140), .ZN(n1290) );
NAND2_X1 U1025 ( .A1(n1216), .A2(n1305), .ZN(n1173) );
NAND2_X1 U1026 ( .A1(n1218), .A2(n1086), .ZN(n1305) );
INV_X1 U1027 ( .A(G898), .ZN(n1086) );
AND3_X1 U1028 ( .A1(G902), .A2(n1037), .A3(n1072), .ZN(n1218) );
XNOR2_X1 U1029 ( .A(G953), .B(KEYINPUT28), .ZN(n1072) );
NAND3_X1 U1030 ( .A1(n1037), .A2(n1032), .A3(G952), .ZN(n1216) );
INV_X1 U1031 ( .A(G953), .ZN(n1032) );
NAND2_X1 U1032 ( .A1(G237), .A2(G234), .ZN(n1037) );
NOR2_X1 U1033 ( .A1(n1019), .A2(n1042), .ZN(n1046) );
INV_X1 U1034 ( .A(n1018), .ZN(n1042) );
NAND2_X1 U1035 ( .A1(G214), .A2(n1306), .ZN(n1018) );
XOR2_X1 U1036 ( .A(n1055), .B(KEYINPUT8), .Z(n1019) );
XOR2_X1 U1037 ( .A(n1307), .B(n1148), .Z(n1055) );
NAND2_X1 U1038 ( .A1(G210), .A2(n1306), .ZN(n1148) );
NAND2_X1 U1039 ( .A1(n1308), .A2(n1231), .ZN(n1306) );
INV_X1 U1040 ( .A(G237), .ZN(n1308) );
NAND2_X1 U1041 ( .A1(n1309), .A2(n1231), .ZN(n1307) );
INV_X1 U1042 ( .A(G902), .ZN(n1231) );
XOR2_X1 U1043 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U1044 ( .A(n1181), .B(n1312), .ZN(n1311) );
NAND3_X1 U1045 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1312) );
OR2_X1 U1046 ( .A1(n1316), .A2(KEYINPUT34), .ZN(n1315) );
INV_X1 U1047 ( .A(n1179), .ZN(n1316) );
NAND3_X1 U1048 ( .A1(KEYINPUT34), .A2(n1317), .A3(n1212), .ZN(n1314) );
OR2_X1 U1049 ( .A1(n1212), .A2(n1317), .ZN(n1313) );
NOR2_X1 U1050 ( .A1(KEYINPUT15), .A2(n1179), .ZN(n1317) );
XOR2_X1 U1051 ( .A(G128), .B(n1272), .Z(n1179) );
XNOR2_X1 U1052 ( .A(n1183), .B(G143), .ZN(n1272) );
INV_X1 U1053 ( .A(G146), .ZN(n1183) );
INV_X1 U1054 ( .A(G125), .ZN(n1212) );
NOR2_X1 U1055 ( .A1(n1085), .A2(G953), .ZN(n1181) );
INV_X1 U1056 ( .A(G224), .ZN(n1085) );
NOR2_X1 U1057 ( .A1(KEYINPUT25), .A2(n1147), .ZN(n1310) );
XOR2_X1 U1058 ( .A(n1098), .B(n1097), .Z(n1147) );
XNOR2_X1 U1059 ( .A(n1318), .B(n1319), .ZN(n1097) );
XOR2_X1 U1060 ( .A(n1320), .B(n1285), .Z(n1319) );
XNOR2_X1 U1061 ( .A(n1224), .B(G122), .ZN(n1285) );
INV_X1 U1062 ( .A(G116), .ZN(n1224) );
NOR2_X1 U1063 ( .A1(KEYINPUT41), .A2(n1221), .ZN(n1320) );
INV_X1 U1064 ( .A(G119), .ZN(n1221) );
XNOR2_X1 U1065 ( .A(G110), .B(G113), .ZN(n1318) );
XOR2_X1 U1066 ( .A(G101), .B(n1321), .Z(n1098) );
NOR2_X1 U1067 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NOR2_X1 U1068 ( .A1(n1287), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1069 ( .A(KEYINPUT57), .B(n1299), .Z(n1324) );
INV_X1 U1070 ( .A(n1296), .ZN(n1322) );
NAND2_X1 U1071 ( .A1(n1299), .A2(n1287), .ZN(n1296) );
XOR2_X1 U1072 ( .A(G107), .B(KEYINPUT27), .Z(n1287) );
XOR2_X1 U1073 ( .A(G104), .B(KEYINPUT1), .Z(n1299) );
INV_X1 U1074 ( .A(G110), .ZN(n1139) );
endmodule


