//Key = 1011011000110000010001000111111101111010110110010110010011001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352;

XOR2_X1 U723 ( .A(G107), .B(n1015), .Z(G9) );
NAND3_X1 U724 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(G75) );
NAND2_X1 U725 ( .A1(G952), .A2(n1019), .ZN(n1018) );
NAND4_X1 U726 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1019) );
NOR2_X1 U727 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
XOR2_X1 U728 ( .A(KEYINPUT29), .B(n1026), .Z(n1025) );
NOR2_X1 U729 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NOR3_X1 U730 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NOR2_X1 U731 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR2_X1 U732 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR2_X1 U733 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U734 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
AND2_X1 U735 ( .A1(n1040), .A2(KEYINPUT58), .ZN(n1036) );
NOR3_X1 U736 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1032) );
NOR3_X1 U737 ( .A1(n1043), .A2(n1044), .A3(n1035), .ZN(n1027) );
NOR2_X1 U738 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
AND3_X1 U739 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NOR4_X1 U740 ( .A1(KEYINPUT58), .A2(n1031), .A3(n1050), .A4(n1051), .ZN(n1045) );
INV_X1 U741 ( .A(n1052), .ZN(n1031) );
NAND2_X1 U742 ( .A1(n1053), .A2(n1054), .ZN(n1022) );
NAND4_X1 U743 ( .A1(n1040), .A2(n1052), .A3(n1055), .A4(n1056), .ZN(n1021) );
XNOR2_X1 U744 ( .A(KEYINPUT18), .B(n1035), .ZN(n1056) );
NAND2_X1 U745 ( .A1(n1047), .A2(n1057), .ZN(n1020) );
NAND2_X1 U746 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U747 ( .A1(n1052), .A2(n1060), .ZN(n1059) );
NAND2_X1 U748 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND3_X1 U749 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
NAND2_X1 U750 ( .A1(n1040), .A2(n1066), .ZN(n1061) );
XOR2_X1 U751 ( .A(KEYINPUT60), .B(n1067), .Z(n1058) );
AND2_X1 U752 ( .A1(n1068), .A2(n1040), .ZN(n1067) );
INV_X1 U753 ( .A(n1043), .ZN(n1040) );
NAND2_X1 U754 ( .A1(n1065), .A2(n1069), .ZN(n1043) );
INV_X1 U755 ( .A(n1039), .ZN(n1065) );
NAND2_X1 U756 ( .A1(n1070), .A2(n1071), .ZN(n1016) );
NAND2_X1 U757 ( .A1(G952), .A2(n1054), .ZN(n1071) );
INV_X1 U758 ( .A(KEYINPUT47), .ZN(n1054) );
INV_X1 U759 ( .A(n1053), .ZN(n1070) );
NAND4_X1 U760 ( .A1(n1072), .A2(n1052), .A3(n1073), .A4(n1074), .ZN(n1053) );
XOR2_X1 U761 ( .A(KEYINPUT14), .B(n1075), .Z(n1074) );
NOR3_X1 U762 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
XOR2_X1 U763 ( .A(KEYINPUT37), .B(n1079), .Z(n1078) );
NOR2_X1 U764 ( .A1(G469), .A2(n1080), .ZN(n1079) );
XOR2_X1 U765 ( .A(n1081), .B(n1082), .Z(n1077) );
XOR2_X1 U766 ( .A(n1083), .B(n1084), .Z(n1082) );
NAND2_X1 U767 ( .A1(KEYINPUT10), .A2(n1085), .ZN(n1084) );
XOR2_X1 U768 ( .A(KEYINPUT32), .B(KEYINPUT17), .Z(n1081) );
NAND3_X1 U769 ( .A1(n1050), .A2(n1041), .A3(n1086), .ZN(n1076) );
NAND2_X1 U770 ( .A1(G469), .A2(n1080), .ZN(n1086) );
NOR2_X1 U771 ( .A1(n1087), .A2(n1088), .ZN(n1073) );
XOR2_X1 U772 ( .A(n1089), .B(KEYINPUT2), .Z(n1088) );
XNOR2_X1 U773 ( .A(n1090), .B(KEYINPUT19), .ZN(n1072) );
NAND2_X1 U774 ( .A1(n1091), .A2(n1092), .ZN(G72) );
NAND3_X1 U775 ( .A1(G953), .A2(n1093), .A3(n1094), .ZN(n1092) );
XOR2_X1 U776 ( .A(KEYINPUT43), .B(n1095), .Z(n1091) );
NOR2_X1 U777 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XNOR2_X1 U778 ( .A(n1094), .B(KEYINPUT61), .ZN(n1097) );
AND2_X1 U779 ( .A1(n1098), .A2(n1099), .ZN(n1094) );
NAND3_X1 U780 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
XOR2_X1 U781 ( .A(KEYINPUT28), .B(n1103), .Z(n1102) );
NAND2_X1 U782 ( .A1(G953), .A2(n1104), .ZN(n1101) );
XOR2_X1 U783 ( .A(n1105), .B(n1106), .Z(n1100) );
NAND2_X1 U784 ( .A1(n1107), .A2(n1103), .ZN(n1098) );
AND2_X1 U785 ( .A1(n1017), .A2(n1108), .ZN(n1103) );
XNOR2_X1 U786 ( .A(n1106), .B(n1105), .ZN(n1107) );
NOR2_X1 U787 ( .A1(KEYINPUT8), .A2(n1109), .ZN(n1105) );
XOR2_X1 U788 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U789 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U790 ( .A1(KEYINPUT22), .A2(n1114), .ZN(n1112) );
XNOR2_X1 U791 ( .A(G128), .B(n1115), .ZN(n1110) );
XNOR2_X1 U792 ( .A(KEYINPUT38), .B(n1116), .ZN(n1115) );
AND2_X1 U793 ( .A1(n1093), .A2(G953), .ZN(n1096) );
NAND2_X1 U794 ( .A1(G900), .A2(G227), .ZN(n1093) );
XOR2_X1 U795 ( .A(n1117), .B(n1118), .Z(G69) );
XOR2_X1 U796 ( .A(n1119), .B(n1120), .Z(n1118) );
NOR2_X1 U797 ( .A1(n1121), .A2(n1017), .ZN(n1120) );
NOR2_X1 U798 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U799 ( .A1(n1124), .A2(n1125), .ZN(n1119) );
XOR2_X1 U800 ( .A(n1126), .B(n1127), .Z(n1125) );
XNOR2_X1 U801 ( .A(n1128), .B(n1129), .ZN(n1127) );
NOR2_X1 U802 ( .A1(G898), .A2(n1017), .ZN(n1124) );
AND2_X1 U803 ( .A1(n1130), .A2(n1017), .ZN(n1117) );
NOR2_X1 U804 ( .A1(n1131), .A2(n1132), .ZN(G66) );
XOR2_X1 U805 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U806 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NOR2_X1 U807 ( .A1(n1131), .A2(n1137), .ZN(G63) );
XNOR2_X1 U808 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR2_X1 U809 ( .A1(n1140), .A2(n1136), .ZN(n1139) );
NOR2_X1 U810 ( .A1(n1131), .A2(n1141), .ZN(G60) );
XNOR2_X1 U811 ( .A(n1142), .B(n1143), .ZN(n1141) );
NOR2_X1 U812 ( .A1(n1144), .A2(n1136), .ZN(n1143) );
XOR2_X1 U813 ( .A(G104), .B(n1145), .Z(G6) );
NOR2_X1 U814 ( .A1(n1131), .A2(n1146), .ZN(G57) );
XOR2_X1 U815 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U816 ( .A(G101), .B(n1149), .ZN(n1148) );
NAND3_X1 U817 ( .A1(n1150), .A2(n1151), .A3(KEYINPUT53), .ZN(n1149) );
NAND2_X1 U818 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND3_X1 U819 ( .A1(G902), .A2(n1154), .A3(G472), .ZN(n1153) );
XNOR2_X1 U820 ( .A(KEYINPUT34), .B(n1024), .ZN(n1154) );
NAND4_X1 U821 ( .A1(n1155), .A2(n1156), .A3(G472), .A4(n1157), .ZN(n1150) );
INV_X1 U822 ( .A(n1152), .ZN(n1157) );
XNOR2_X1 U823 ( .A(n1158), .B(n1159), .ZN(n1152) );
XOR2_X1 U824 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U825 ( .A(n1162), .B(n1163), .Z(n1158) );
XOR2_X1 U826 ( .A(n1164), .B(KEYINPUT15), .Z(n1162) );
NAND2_X1 U827 ( .A1(KEYINPUT34), .A2(n1136), .ZN(n1156) );
NAND2_X1 U828 ( .A1(n1165), .A2(n1166), .ZN(n1155) );
INV_X1 U829 ( .A(KEYINPUT34), .ZN(n1166) );
NAND2_X1 U830 ( .A1(n1167), .A2(G902), .ZN(n1165) );
NOR2_X1 U831 ( .A1(KEYINPUT63), .A2(n1168), .ZN(n1147) );
NOR2_X1 U832 ( .A1(n1131), .A2(n1169), .ZN(G54) );
XOR2_X1 U833 ( .A(n1170), .B(n1171), .Z(n1169) );
XNOR2_X1 U834 ( .A(n1172), .B(n1173), .ZN(n1171) );
XOR2_X1 U835 ( .A(n1174), .B(n1175), .Z(n1170) );
XOR2_X1 U836 ( .A(KEYINPUT24), .B(n1176), .Z(n1175) );
NOR2_X1 U837 ( .A1(n1177), .A2(n1136), .ZN(n1176) );
NOR2_X1 U838 ( .A1(n1131), .A2(n1178), .ZN(G51) );
XOR2_X1 U839 ( .A(n1179), .B(n1180), .Z(n1178) );
XNOR2_X1 U840 ( .A(n1181), .B(n1182), .ZN(n1180) );
NOR2_X1 U841 ( .A1(n1085), .A2(n1136), .ZN(n1181) );
NAND2_X1 U842 ( .A1(G902), .A2(n1024), .ZN(n1136) );
INV_X1 U843 ( .A(n1167), .ZN(n1024) );
NOR2_X1 U844 ( .A1(n1130), .A2(n1108), .ZN(n1167) );
NAND4_X1 U845 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1108) );
AND4_X1 U846 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1186) );
NOR2_X1 U847 ( .A1(n1191), .A2(n1192), .ZN(n1185) );
NOR2_X1 U848 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NOR2_X1 U849 ( .A1(n1064), .A2(n1195), .ZN(n1193) );
XNOR2_X1 U850 ( .A(KEYINPUT12), .B(n1038), .ZN(n1195) );
NOR3_X1 U851 ( .A1(n1196), .A2(n1055), .A3(n1197), .ZN(n1191) );
NOR2_X1 U852 ( .A1(n1198), .A2(n1199), .ZN(n1196) );
NOR4_X1 U853 ( .A1(KEYINPUT27), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1199) );
NOR2_X1 U854 ( .A1(n1203), .A2(n1204), .ZN(n1198) );
NAND2_X1 U855 ( .A1(KEYINPUT27), .A2(n1205), .ZN(n1184) );
NAND2_X1 U856 ( .A1(n1206), .A2(n1204), .ZN(n1183) );
INV_X1 U857 ( .A(KEYINPUT54), .ZN(n1204) );
NAND4_X1 U858 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1130) );
NOR4_X1 U859 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1145), .ZN(n1210) );
AND3_X1 U860 ( .A1(n1052), .A2(n1064), .A3(n1214), .ZN(n1145) );
NOR2_X1 U861 ( .A1(n1015), .A2(n1215), .ZN(n1209) );
AND3_X1 U862 ( .A1(n1216), .A2(n1052), .A3(n1214), .ZN(n1015) );
XOR2_X1 U863 ( .A(n1217), .B(n1218), .Z(n1179) );
NOR2_X1 U864 ( .A1(n1017), .A2(G952), .ZN(n1131) );
XNOR2_X1 U865 ( .A(G146), .B(n1190), .ZN(G48) );
NAND4_X1 U866 ( .A1(n1219), .A2(n1066), .A3(n1055), .A4(n1220), .ZN(n1190) );
XOR2_X1 U867 ( .A(G143), .B(n1205), .Z(G45) );
AND4_X1 U868 ( .A1(n1055), .A2(n1221), .A3(n1066), .A4(n1222), .ZN(n1205) );
NOR2_X1 U869 ( .A1(n1201), .A2(n1202), .ZN(n1222) );
XNOR2_X1 U870 ( .A(G140), .B(n1189), .ZN(G42) );
NAND4_X1 U871 ( .A1(n1047), .A2(n1219), .A3(n1049), .A4(n1066), .ZN(n1189) );
INV_X1 U872 ( .A(n1029), .ZN(n1047) );
XNOR2_X1 U873 ( .A(G137), .B(n1188), .ZN(G39) );
NAND3_X1 U874 ( .A1(n1223), .A2(n1220), .A3(n1224), .ZN(n1188) );
XOR2_X1 U875 ( .A(G134), .B(n1225), .Z(G36) );
NOR2_X1 U876 ( .A1(n1038), .A2(n1194), .ZN(n1225) );
INV_X1 U877 ( .A(n1216), .ZN(n1038) );
XOR2_X1 U878 ( .A(n1226), .B(n1227), .Z(G33) );
NAND2_X1 U879 ( .A1(n1228), .A2(n1064), .ZN(n1227) );
INV_X1 U880 ( .A(n1194), .ZN(n1228) );
NAND2_X1 U881 ( .A1(n1224), .A2(n1229), .ZN(n1194) );
NOR3_X1 U882 ( .A1(n1200), .A2(n1197), .A3(n1029), .ZN(n1224) );
NAND2_X1 U883 ( .A1(n1230), .A2(n1050), .ZN(n1029) );
INV_X1 U884 ( .A(n1051), .ZN(n1230) );
NAND2_X1 U885 ( .A1(n1231), .A2(KEYINPUT25), .ZN(n1226) );
XNOR2_X1 U886 ( .A(G131), .B(KEYINPUT3), .ZN(n1231) );
NAND2_X1 U887 ( .A1(n1232), .A2(n1233), .ZN(G30) );
NAND2_X1 U888 ( .A1(n1206), .A2(n1234), .ZN(n1233) );
XOR2_X1 U889 ( .A(n1235), .B(KEYINPUT16), .Z(n1232) );
OR2_X1 U890 ( .A1(n1234), .A2(n1206), .ZN(n1235) );
NOR3_X1 U891 ( .A1(n1236), .A2(n1197), .A3(n1203), .ZN(n1206) );
NAND4_X1 U892 ( .A1(n1237), .A2(n1216), .A3(n1048), .A4(n1220), .ZN(n1203) );
INV_X1 U893 ( .A(n1221), .ZN(n1197) );
XOR2_X1 U894 ( .A(G101), .B(n1213), .Z(G3) );
AND3_X1 U895 ( .A1(n1214), .A2(n1069), .A3(n1229), .ZN(n1213) );
XNOR2_X1 U896 ( .A(G125), .B(n1187), .ZN(G27) );
NAND4_X1 U897 ( .A1(n1219), .A2(n1063), .A3(n1049), .A4(n1055), .ZN(n1187) );
AND3_X1 U898 ( .A1(n1048), .A2(n1221), .A3(n1064), .ZN(n1219) );
NAND2_X1 U899 ( .A1(n1039), .A2(n1238), .ZN(n1221) );
NAND4_X1 U900 ( .A1(G953), .A2(G902), .A3(n1239), .A4(n1104), .ZN(n1238) );
INV_X1 U901 ( .A(G900), .ZN(n1104) );
XOR2_X1 U902 ( .A(G122), .B(n1212), .Z(G24) );
AND3_X1 U903 ( .A1(n1240), .A2(n1052), .A3(n1241), .ZN(n1212) );
NOR2_X1 U904 ( .A1(n1220), .A2(n1048), .ZN(n1052) );
XNOR2_X1 U905 ( .A(n1211), .B(n1242), .ZN(G21) );
XNOR2_X1 U906 ( .A(G119), .B(KEYINPUT9), .ZN(n1242) );
AND3_X1 U907 ( .A1(n1223), .A2(n1220), .A3(n1241), .ZN(n1211) );
XNOR2_X1 U908 ( .A(G116), .B(n1207), .ZN(G18) );
NAND3_X1 U909 ( .A1(n1229), .A2(n1216), .A3(n1241), .ZN(n1207) );
AND3_X1 U910 ( .A1(n1055), .A2(n1243), .A3(n1063), .ZN(n1241) );
XNOR2_X1 U911 ( .A(n1244), .B(n1208), .ZN(G15) );
NAND4_X1 U912 ( .A1(n1245), .A2(n1068), .A3(n1064), .A4(n1243), .ZN(n1208) );
NAND2_X1 U913 ( .A1(n1246), .A2(n1247), .ZN(n1064) );
NAND3_X1 U914 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1247) );
INV_X1 U915 ( .A(KEYINPUT52), .ZN(n1250) );
NAND2_X1 U916 ( .A1(KEYINPUT52), .A2(n1240), .ZN(n1246) );
INV_X1 U917 ( .A(n1202), .ZN(n1240) );
NAND2_X1 U918 ( .A1(n1248), .A2(n1090), .ZN(n1202) );
NOR2_X1 U919 ( .A1(n1201), .A2(n1035), .ZN(n1068) );
INV_X1 U920 ( .A(n1063), .ZN(n1035) );
NOR2_X1 U921 ( .A1(n1042), .A2(n1251), .ZN(n1063) );
INV_X1 U922 ( .A(n1041), .ZN(n1251) );
XNOR2_X1 U923 ( .A(n1252), .B(KEYINPUT31), .ZN(n1042) );
INV_X1 U924 ( .A(n1229), .ZN(n1201) );
NOR2_X1 U925 ( .A1(n1048), .A2(n1049), .ZN(n1229) );
NAND2_X1 U926 ( .A1(KEYINPUT26), .A2(n1253), .ZN(n1244) );
XOR2_X1 U927 ( .A(G110), .B(n1215), .Z(G12) );
AND3_X1 U928 ( .A1(n1049), .A2(n1214), .A3(n1223), .ZN(n1215) );
AND2_X1 U929 ( .A1(n1069), .A2(n1048), .ZN(n1223) );
XOR2_X1 U930 ( .A(n1254), .B(n1135), .Z(n1048) );
NAND2_X1 U931 ( .A1(G217), .A2(n1255), .ZN(n1135) );
NAND2_X1 U932 ( .A1(n1256), .A2(n1257), .ZN(n1254) );
XNOR2_X1 U933 ( .A(n1134), .B(KEYINPUT4), .ZN(n1256) );
XNOR2_X1 U934 ( .A(n1258), .B(n1259), .ZN(n1134) );
XNOR2_X1 U935 ( .A(G119), .B(n1260), .ZN(n1259) );
NAND2_X1 U936 ( .A1(n1261), .A2(G221), .ZN(n1260) );
XNOR2_X1 U937 ( .A(n1174), .B(n1262), .ZN(n1258) );
NOR2_X1 U938 ( .A1(G125), .A2(KEYINPUT39), .ZN(n1262) );
XOR2_X1 U939 ( .A(n1263), .B(n1264), .Z(n1174) );
NAND2_X1 U940 ( .A1(n1265), .A2(n1266), .ZN(n1069) );
OR3_X1 U941 ( .A1(n1248), .A2(n1090), .A3(KEYINPUT52), .ZN(n1266) );
NAND2_X1 U942 ( .A1(KEYINPUT52), .A2(n1216), .ZN(n1265) );
NOR2_X1 U943 ( .A1(n1248), .A2(n1249), .ZN(n1216) );
INV_X1 U944 ( .A(n1090), .ZN(n1249) );
XOR2_X1 U945 ( .A(n1267), .B(n1140), .Z(n1090) );
INV_X1 U946 ( .A(G478), .ZN(n1140) );
NAND2_X1 U947 ( .A1(n1138), .A2(n1257), .ZN(n1267) );
XNOR2_X1 U948 ( .A(n1268), .B(n1269), .ZN(n1138) );
XOR2_X1 U949 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U950 ( .A(G107), .B(n1272), .Z(n1271) );
NOR2_X1 U951 ( .A1(KEYINPUT7), .A2(n1273), .ZN(n1272) );
XNOR2_X1 U952 ( .A(n1234), .B(n1274), .ZN(n1273) );
XOR2_X1 U953 ( .A(G143), .B(G134), .Z(n1274) );
INV_X1 U954 ( .A(G128), .ZN(n1234) );
AND2_X1 U955 ( .A1(n1261), .A2(G217), .ZN(n1270) );
AND2_X1 U956 ( .A1(G234), .A2(n1017), .ZN(n1261) );
XNOR2_X1 U957 ( .A(G116), .B(n1275), .ZN(n1268) );
XOR2_X1 U958 ( .A(KEYINPUT49), .B(G122), .Z(n1275) );
NAND2_X1 U959 ( .A1(n1276), .A2(n1277), .ZN(n1248) );
NAND2_X1 U960 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
INV_X1 U961 ( .A(KEYINPUT45), .ZN(n1279) );
NAND2_X1 U962 ( .A1(n1280), .A2(n1089), .ZN(n1278) );
NAND2_X1 U963 ( .A1(n1281), .A2(n1144), .ZN(n1089) );
INV_X1 U964 ( .A(n1087), .ZN(n1280) );
NOR2_X1 U965 ( .A1(n1144), .A2(n1281), .ZN(n1087) );
INV_X1 U966 ( .A(G475), .ZN(n1144) );
NAND2_X1 U967 ( .A1(KEYINPUT45), .A2(n1282), .ZN(n1276) );
XNOR2_X1 U968 ( .A(n1281), .B(G475), .ZN(n1282) );
AND2_X1 U969 ( .A1(n1283), .A2(n1257), .ZN(n1281) );
XNOR2_X1 U970 ( .A(KEYINPUT62), .B(n1284), .ZN(n1283) );
INV_X1 U971 ( .A(n1142), .ZN(n1284) );
XNOR2_X1 U972 ( .A(n1285), .B(n1286), .ZN(n1142) );
XOR2_X1 U973 ( .A(G104), .B(n1287), .Z(n1286) );
XNOR2_X1 U974 ( .A(G122), .B(n1253), .ZN(n1287) );
INV_X1 U975 ( .A(G113), .ZN(n1253) );
XOR2_X1 U976 ( .A(n1288), .B(n1289), .Z(n1285) );
XOR2_X1 U977 ( .A(n1290), .B(n1291), .Z(n1289) );
NAND3_X1 U978 ( .A1(n1292), .A2(n1017), .A3(G214), .ZN(n1291) );
NAND2_X1 U979 ( .A1(n1293), .A2(n1294), .ZN(n1290) );
OR2_X1 U980 ( .A1(n1106), .A2(n1295), .ZN(n1294) );
XOR2_X1 U981 ( .A(n1296), .B(KEYINPUT59), .Z(n1293) );
NAND2_X1 U982 ( .A1(n1295), .A2(n1106), .ZN(n1296) );
XNOR2_X1 U983 ( .A(G140), .B(n1297), .ZN(n1106) );
XOR2_X1 U984 ( .A(G146), .B(KEYINPUT55), .Z(n1295) );
AND3_X1 U985 ( .A1(n1237), .A2(n1243), .A3(n1245), .ZN(n1214) );
XNOR2_X1 U986 ( .A(n1055), .B(KEYINPUT40), .ZN(n1245) );
INV_X1 U987 ( .A(n1236), .ZN(n1055) );
NAND2_X1 U988 ( .A1(n1051), .A2(n1050), .ZN(n1236) );
NAND2_X1 U989 ( .A1(G214), .A2(n1298), .ZN(n1050) );
XOR2_X1 U990 ( .A(n1083), .B(n1085), .Z(n1051) );
NAND2_X1 U991 ( .A1(G210), .A2(n1298), .ZN(n1085) );
NAND2_X1 U992 ( .A1(n1292), .A2(n1257), .ZN(n1298) );
NAND2_X1 U993 ( .A1(n1299), .A2(n1257), .ZN(n1083) );
XOR2_X1 U994 ( .A(n1300), .B(n1301), .Z(n1299) );
XNOR2_X1 U995 ( .A(KEYINPUT13), .B(n1302), .ZN(n1301) );
NOR2_X1 U996 ( .A1(n1217), .A2(KEYINPUT46), .ZN(n1302) );
AND2_X1 U997 ( .A1(n1303), .A2(n1304), .ZN(n1217) );
NAND2_X1 U998 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND2_X1 U999 ( .A1(KEYINPUT57), .A2(n1307), .ZN(n1306) );
NAND2_X1 U1000 ( .A1(KEYINPUT35), .A2(n1128), .ZN(n1307) );
NAND2_X1 U1001 ( .A1(n1308), .A2(n1309), .ZN(n1303) );
NAND2_X1 U1002 ( .A1(KEYINPUT35), .A2(n1310), .ZN(n1309) );
NAND2_X1 U1003 ( .A1(n1311), .A2(KEYINPUT57), .ZN(n1310) );
INV_X1 U1004 ( .A(n1305), .ZN(n1311) );
NAND2_X1 U1005 ( .A1(n1312), .A2(n1313), .ZN(n1305) );
OR2_X1 U1006 ( .A1(n1126), .A2(n1129), .ZN(n1313) );
XOR2_X1 U1007 ( .A(n1314), .B(KEYINPUT42), .Z(n1312) );
NAND2_X1 U1008 ( .A1(n1129), .A2(n1126), .ZN(n1314) );
XOR2_X1 U1009 ( .A(n1160), .B(KEYINPUT36), .Z(n1126) );
XOR2_X1 U1010 ( .A(G101), .B(n1315), .Z(n1129) );
NOR2_X1 U1011 ( .A1(KEYINPUT51), .A2(n1316), .ZN(n1315) );
XOR2_X1 U1012 ( .A(n1317), .B(n1318), .Z(n1316) );
XOR2_X1 U1013 ( .A(KEYINPUT30), .B(G104), .Z(n1318) );
NOR2_X1 U1014 ( .A1(G107), .A2(KEYINPUT20), .ZN(n1317) );
INV_X1 U1015 ( .A(n1128), .ZN(n1308) );
XNOR2_X1 U1016 ( .A(G110), .B(G122), .ZN(n1128) );
NAND2_X1 U1017 ( .A1(n1319), .A2(n1320), .ZN(n1300) );
NAND2_X1 U1018 ( .A1(n1182), .A2(n1321), .ZN(n1320) );
NAND2_X1 U1019 ( .A1(KEYINPUT41), .A2(G224), .ZN(n1321) );
INV_X1 U1020 ( .A(n1322), .ZN(n1182) );
NAND3_X1 U1021 ( .A1(KEYINPUT41), .A2(n1218), .A3(n1322), .ZN(n1319) );
XOR2_X1 U1022 ( .A(n1323), .B(n1297), .Z(n1322) );
INV_X1 U1023 ( .A(G125), .ZN(n1297) );
NOR2_X1 U1024 ( .A1(n1122), .A2(G953), .ZN(n1218) );
INV_X1 U1025 ( .A(G224), .ZN(n1122) );
NAND2_X1 U1026 ( .A1(n1039), .A2(n1324), .ZN(n1243) );
NAND4_X1 U1027 ( .A1(G953), .A2(G902), .A3(n1325), .A4(n1123), .ZN(n1324) );
INV_X1 U1028 ( .A(G898), .ZN(n1123) );
XNOR2_X1 U1029 ( .A(KEYINPUT56), .B(n1239), .ZN(n1325) );
NAND3_X1 U1030 ( .A1(n1239), .A2(n1017), .A3(G952), .ZN(n1039) );
NAND2_X1 U1031 ( .A1(G237), .A2(G234), .ZN(n1239) );
XNOR2_X1 U1032 ( .A(n1066), .B(KEYINPUT21), .ZN(n1237) );
INV_X1 U1033 ( .A(n1200), .ZN(n1066) );
NAND2_X1 U1034 ( .A1(n1252), .A2(n1041), .ZN(n1200) );
NAND2_X1 U1035 ( .A1(G221), .A2(n1255), .ZN(n1041) );
NAND2_X1 U1036 ( .A1(G234), .A2(n1257), .ZN(n1255) );
XOR2_X1 U1037 ( .A(n1080), .B(n1177), .Z(n1252) );
INV_X1 U1038 ( .A(G469), .ZN(n1177) );
NAND2_X1 U1039 ( .A1(n1326), .A2(n1257), .ZN(n1080) );
XNOR2_X1 U1040 ( .A(n1327), .B(n1328), .ZN(n1326) );
INV_X1 U1041 ( .A(n1172), .ZN(n1328) );
XNOR2_X1 U1042 ( .A(n1329), .B(KEYINPUT0), .ZN(n1172) );
NAND2_X1 U1043 ( .A1(G227), .A2(n1017), .ZN(n1329) );
XNOR2_X1 U1044 ( .A(n1264), .B(n1330), .ZN(n1327) );
NOR2_X1 U1045 ( .A1(KEYINPUT1), .A2(n1331), .ZN(n1330) );
XOR2_X1 U1046 ( .A(n1173), .B(n1263), .Z(n1331) );
XOR2_X1 U1047 ( .A(G128), .B(n1163), .Z(n1263) );
XNOR2_X1 U1048 ( .A(n1114), .B(G146), .ZN(n1163) );
INV_X1 U1049 ( .A(G137), .ZN(n1114) );
XOR2_X1 U1050 ( .A(n1332), .B(n1333), .Z(n1173) );
XOR2_X1 U1051 ( .A(G107), .B(G104), .Z(n1333) );
XOR2_X1 U1052 ( .A(n1334), .B(n1113), .Z(n1332) );
XOR2_X1 U1053 ( .A(n1161), .B(KEYINPUT5), .Z(n1113) );
XNOR2_X1 U1054 ( .A(n1288), .B(n1335), .ZN(n1161) );
XNOR2_X1 U1055 ( .A(G131), .B(G143), .ZN(n1288) );
XNOR2_X1 U1056 ( .A(G110), .B(n1336), .ZN(n1264) );
INV_X1 U1057 ( .A(G140), .ZN(n1336) );
INV_X1 U1058 ( .A(n1220), .ZN(n1049) );
XNOR2_X1 U1059 ( .A(n1337), .B(G472), .ZN(n1220) );
NAND2_X1 U1060 ( .A1(n1338), .A2(n1257), .ZN(n1337) );
INV_X1 U1061 ( .A(G902), .ZN(n1257) );
XOR2_X1 U1062 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1063 ( .A(n1341), .B(n1342), .Z(n1340) );
XNOR2_X1 U1064 ( .A(n1343), .B(n1344), .ZN(n1342) );
INV_X1 U1065 ( .A(G131), .ZN(n1344) );
NAND2_X1 U1066 ( .A1(KEYINPUT50), .A2(n1345), .ZN(n1343) );
INV_X1 U1067 ( .A(n1168), .ZN(n1345) );
NAND3_X1 U1068 ( .A1(n1292), .A2(n1017), .A3(G210), .ZN(n1168) );
INV_X1 U1069 ( .A(G953), .ZN(n1017) );
INV_X1 U1070 ( .A(G237), .ZN(n1292) );
XNOR2_X1 U1071 ( .A(G137), .B(KEYINPUT11), .ZN(n1341) );
XOR2_X1 U1072 ( .A(n1346), .B(n1347), .Z(n1339) );
XNOR2_X1 U1073 ( .A(n1348), .B(n1349), .ZN(n1347) );
NOR2_X1 U1074 ( .A1(KEYINPUT48), .A2(n1323), .ZN(n1349) );
XOR2_X1 U1075 ( .A(n1164), .B(n1350), .Z(n1323) );
XNOR2_X1 U1076 ( .A(n1116), .B(G143), .ZN(n1350) );
INV_X1 U1077 ( .A(G146), .ZN(n1116) );
NAND2_X1 U1078 ( .A1(n1351), .A2(KEYINPUT44), .ZN(n1164) );
XNOR2_X1 U1079 ( .A(G128), .B(KEYINPUT23), .ZN(n1351) );
NAND2_X1 U1080 ( .A1(KEYINPUT6), .A2(n1160), .ZN(n1348) );
XOR2_X1 U1081 ( .A(G113), .B(n1352), .Z(n1160) );
XOR2_X1 U1082 ( .A(G119), .B(G116), .Z(n1352) );
XOR2_X1 U1083 ( .A(n1334), .B(n1335), .Z(n1346) );
XOR2_X1 U1084 ( .A(G134), .B(KEYINPUT33), .Z(n1335) );
XNOR2_X1 U1085 ( .A(KEYINPUT15), .B(G101), .ZN(n1334) );
endmodule


