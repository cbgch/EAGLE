//Key = 0010011111001001101110010100011111111001000111101110110010011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380;

XNOR2_X1 U751 ( .A(G107), .B(n1048), .ZN(G9) );
NAND4_X1 U752 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(G75) );
NAND4_X1 U753 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1051) );
NOR4_X1 U754 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
NOR3_X1 U755 ( .A1(n1061), .A2(KEYINPUT41), .A3(n1062), .ZN(n1060) );
AND2_X1 U756 ( .A1(n1061), .A2(KEYINPUT41), .ZN(n1059) );
NAND3_X1 U757 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1057) );
XNOR2_X1 U758 ( .A(KEYINPUT8), .B(n1066), .ZN(n1065) );
XOR2_X1 U759 ( .A(n1067), .B(n1068), .Z(n1064) );
XOR2_X1 U760 ( .A(KEYINPUT57), .B(KEYINPUT2), .Z(n1068) );
XNOR2_X1 U761 ( .A(n1069), .B(n1070), .ZN(n1063) );
NAND2_X1 U762 ( .A1(KEYINPUT9), .A2(n1071), .ZN(n1070) );
NOR3_X1 U763 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1055) );
NAND2_X1 U764 ( .A1(n1075), .A2(n1076), .ZN(n1050) );
NAND2_X1 U765 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND4_X1 U766 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1053), .ZN(n1078) );
NAND2_X1 U767 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U768 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
OR2_X1 U769 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U770 ( .A1(n1088), .A2(n1089), .ZN(n1082) );
NAND2_X1 U771 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND3_X1 U772 ( .A1(n1092), .A2(n1054), .A3(n1074), .ZN(n1091) );
INV_X1 U773 ( .A(n1093), .ZN(n1074) );
NAND3_X1 U774 ( .A1(n1088), .A2(n1094), .A3(n1084), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND3_X1 U776 ( .A1(n1097), .A2(n1098), .A3(n1080), .ZN(n1096) );
OR2_X1 U777 ( .A1(n1053), .A2(n1079), .ZN(n1098) );
OR3_X1 U778 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1097) );
NAND2_X1 U779 ( .A1(n1102), .A2(n1079), .ZN(n1095) );
INV_X1 U780 ( .A(n1103), .ZN(n1075) );
XOR2_X1 U781 ( .A(n1104), .B(n1105), .Z(G72) );
NAND2_X1 U782 ( .A1(G953), .A2(n1106), .ZN(n1105) );
NAND2_X1 U783 ( .A1(G900), .A2(G227), .ZN(n1106) );
NAND2_X1 U784 ( .A1(KEYINPUT5), .A2(n1107), .ZN(n1104) );
XOR2_X1 U785 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U786 ( .A1(n1052), .A2(n1110), .ZN(n1109) );
NAND2_X1 U787 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
NAND2_X1 U788 ( .A1(G953), .A2(n1113), .ZN(n1112) );
XOR2_X1 U789 ( .A(n1114), .B(n1115), .Z(n1111) );
XNOR2_X1 U790 ( .A(n1116), .B(n1117), .ZN(n1115) );
NAND2_X1 U791 ( .A1(KEYINPUT49), .A2(n1118), .ZN(n1116) );
XNOR2_X1 U792 ( .A(KEYINPUT34), .B(n1119), .ZN(n1114) );
NOR2_X1 U793 ( .A1(KEYINPUT4), .A2(n1120), .ZN(n1119) );
XOR2_X1 U794 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U795 ( .A1(KEYINPUT21), .A2(n1123), .ZN(n1121) );
XOR2_X1 U796 ( .A(n1124), .B(n1125), .Z(G69) );
NOR2_X1 U797 ( .A1(n1052), .A2(n1126), .ZN(n1125) );
XOR2_X1 U798 ( .A(KEYINPUT58), .B(n1127), .Z(n1126) );
NOR2_X1 U799 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U800 ( .A1(n1130), .A2(n1131), .ZN(n1124) );
NAND2_X1 U801 ( .A1(n1132), .A2(n1052), .ZN(n1131) );
XOR2_X1 U802 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND3_X1 U803 ( .A1(G898), .A2(n1133), .A3(G953), .ZN(n1130) );
XOR2_X1 U804 ( .A(n1135), .B(KEYINPUT55), .Z(n1133) );
NOR2_X1 U805 ( .A1(n1136), .A2(n1137), .ZN(G66) );
XOR2_X1 U806 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND3_X1 U807 ( .A1(n1140), .A2(n1141), .A3(KEYINPUT56), .ZN(n1138) );
NOR2_X1 U808 ( .A1(n1136), .A2(n1142), .ZN(G63) );
XOR2_X1 U809 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U810 ( .A(n1145), .B(n1146), .ZN(n1144) );
AND2_X1 U811 ( .A1(G478), .A2(n1140), .ZN(n1146) );
XOR2_X1 U812 ( .A(KEYINPUT60), .B(KEYINPUT38), .Z(n1143) );
NOR2_X1 U813 ( .A1(n1136), .A2(n1147), .ZN(G60) );
NOR3_X1 U814 ( .A1(n1069), .A2(n1148), .A3(n1149), .ZN(n1147) );
AND4_X1 U815 ( .A1(n1150), .A2(KEYINPUT15), .A3(G475), .A4(n1140), .ZN(n1149) );
NOR2_X1 U816 ( .A1(n1151), .A2(n1150), .ZN(n1148) );
NOR3_X1 U817 ( .A1(n1152), .A2(n1049), .A3(n1071), .ZN(n1151) );
INV_X1 U818 ( .A(KEYINPUT15), .ZN(n1152) );
XNOR2_X1 U819 ( .A(G104), .B(n1153), .ZN(G6) );
NOR2_X1 U820 ( .A1(n1154), .A2(n1155), .ZN(G57) );
XOR2_X1 U821 ( .A(n1156), .B(n1157), .Z(n1155) );
XNOR2_X1 U822 ( .A(n1158), .B(n1159), .ZN(n1157) );
NAND2_X1 U823 ( .A1(KEYINPUT63), .A2(n1160), .ZN(n1158) );
XOR2_X1 U824 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U825 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U826 ( .A1(KEYINPUT62), .A2(n1165), .ZN(n1164) );
AND2_X1 U827 ( .A1(G472), .A2(n1140), .ZN(n1163) );
NAND2_X1 U828 ( .A1(KEYINPUT44), .A2(G101), .ZN(n1156) );
XNOR2_X1 U829 ( .A(n1136), .B(KEYINPUT36), .ZN(n1154) );
NOR2_X1 U830 ( .A1(n1136), .A2(n1166), .ZN(G54) );
XOR2_X1 U831 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U832 ( .A(KEYINPUT1), .B(n1169), .Z(n1168) );
NOR2_X1 U833 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NOR2_X1 U834 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NOR2_X1 U835 ( .A1(n1174), .A2(n1175), .ZN(n1172) );
INV_X1 U836 ( .A(KEYINPUT16), .ZN(n1175) );
NOR2_X1 U837 ( .A1(n1176), .A2(n1177), .ZN(n1174) );
NOR2_X1 U838 ( .A1(n1178), .A2(n1179), .ZN(n1170) );
NOR2_X1 U839 ( .A1(n1180), .A2(n1177), .ZN(n1179) );
INV_X1 U840 ( .A(KEYINPUT31), .ZN(n1177) );
AND2_X1 U841 ( .A1(n1173), .A2(KEYINPUT16), .ZN(n1180) );
NAND2_X1 U842 ( .A1(n1181), .A2(n1182), .ZN(n1173) );
NAND2_X1 U843 ( .A1(KEYINPUT10), .A2(n1183), .ZN(n1182) );
NAND2_X1 U844 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
INV_X1 U845 ( .A(n1186), .ZN(n1184) );
NAND2_X1 U846 ( .A1(n1187), .A2(n1188), .ZN(n1181) );
INV_X1 U847 ( .A(KEYINPUT10), .ZN(n1188) );
XNOR2_X1 U848 ( .A(G110), .B(n1189), .ZN(n1187) );
INV_X1 U849 ( .A(n1176), .ZN(n1178) );
XOR2_X1 U850 ( .A(n1190), .B(n1191), .Z(n1167) );
NOR2_X1 U851 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NOR2_X1 U852 ( .A1(n1136), .A2(n1194), .ZN(G51) );
XOR2_X1 U853 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U854 ( .A(n1197), .B(n1198), .Z(n1196) );
XNOR2_X1 U855 ( .A(n1135), .B(n1199), .ZN(n1195) );
NOR2_X1 U856 ( .A1(n1200), .A2(n1193), .ZN(n1199) );
INV_X1 U857 ( .A(n1140), .ZN(n1193) );
NOR2_X1 U858 ( .A1(n1201), .A2(n1049), .ZN(n1140) );
NOR2_X1 U859 ( .A1(n1110), .A2(n1134), .ZN(n1049) );
NAND4_X1 U860 ( .A1(n1202), .A2(n1153), .A3(n1203), .A4(n1204), .ZN(n1134) );
AND4_X1 U861 ( .A1(n1048), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1204) );
NAND3_X1 U862 ( .A1(n1087), .A2(n1079), .A3(n1208), .ZN(n1048) );
NAND2_X1 U863 ( .A1(n1209), .A2(n1210), .ZN(n1203) );
INV_X1 U864 ( .A(KEYINPUT40), .ZN(n1210) );
NAND3_X1 U865 ( .A1(n1208), .A2(n1079), .A3(n1086), .ZN(n1153) );
NAND2_X1 U866 ( .A1(n1102), .A2(n1211), .ZN(n1202) );
NAND3_X1 U867 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1211) );
NAND2_X1 U868 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND4_X1 U869 ( .A1(KEYINPUT40), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1212) );
NAND4_X1 U870 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1110) );
NOR4_X1 U871 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1223) );
INV_X1 U872 ( .A(n1228), .ZN(n1224) );
NOR2_X1 U873 ( .A1(n1229), .A2(n1230), .ZN(n1222) );
INV_X1 U874 ( .A(n1231), .ZN(n1230) );
OR2_X1 U875 ( .A1(n1218), .A2(n1232), .ZN(n1220) );
NOR2_X1 U876 ( .A1(n1052), .A2(G952), .ZN(n1136) );
XNOR2_X1 U877 ( .A(G146), .B(n1231), .ZN(G48) );
NAND2_X1 U878 ( .A1(n1086), .A2(n1233), .ZN(n1231) );
XNOR2_X1 U879 ( .A(G143), .B(n1221), .ZN(G45) );
NAND4_X1 U880 ( .A1(n1234), .A2(n1100), .A3(n1235), .A4(n1236), .ZN(n1221) );
XOR2_X1 U881 ( .A(G140), .B(n1229), .Z(G42) );
AND3_X1 U882 ( .A1(n1237), .A2(n1086), .A3(n1099), .ZN(n1229) );
XNOR2_X1 U883 ( .A(n1227), .B(n1238), .ZN(G39) );
NOR2_X1 U884 ( .A1(G137), .A2(KEYINPUT47), .ZN(n1238) );
AND2_X1 U885 ( .A1(n1217), .A2(n1237), .ZN(n1227) );
XOR2_X1 U886 ( .A(G134), .B(n1226), .Z(G36) );
AND3_X1 U887 ( .A1(n1087), .A2(n1100), .A3(n1237), .ZN(n1226) );
XOR2_X1 U888 ( .A(G131), .B(n1225), .Z(G33) );
AND2_X1 U889 ( .A1(n1237), .A2(n1216), .ZN(n1225) );
INV_X1 U890 ( .A(n1239), .ZN(n1216) );
AND4_X1 U891 ( .A1(n1235), .A2(n1080), .A3(n1236), .A4(n1053), .ZN(n1237) );
XNOR2_X1 U892 ( .A(G128), .B(n1228), .ZN(G30) );
NAND2_X1 U893 ( .A1(n1233), .A2(n1087), .ZN(n1228) );
AND4_X1 U894 ( .A1(n1236), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1233) );
AND2_X1 U895 ( .A1(n1235), .A2(n1102), .ZN(n1242) );
XNOR2_X1 U896 ( .A(G101), .B(n1207), .ZN(G3) );
NAND3_X1 U897 ( .A1(n1208), .A2(n1100), .A3(n1088), .ZN(n1207) );
XOR2_X1 U898 ( .A(G125), .B(n1243), .Z(G27) );
NOR2_X1 U899 ( .A1(n1244), .A2(n1232), .ZN(n1243) );
NAND4_X1 U900 ( .A1(n1099), .A2(n1086), .A3(n1102), .A4(n1236), .ZN(n1232) );
NAND2_X1 U901 ( .A1(n1103), .A2(n1245), .ZN(n1236) );
NAND2_X1 U902 ( .A1(n1246), .A2(n1113), .ZN(n1245) );
INV_X1 U903 ( .A(G900), .ZN(n1113) );
XNOR2_X1 U904 ( .A(n1084), .B(KEYINPUT3), .ZN(n1244) );
XOR2_X1 U905 ( .A(n1206), .B(n1247), .Z(G24) );
NAND2_X1 U906 ( .A1(KEYINPUT39), .A2(G122), .ZN(n1247) );
NAND3_X1 U907 ( .A1(n1234), .A2(n1079), .A3(n1215), .ZN(n1206) );
NAND2_X1 U908 ( .A1(n1248), .A2(n1249), .ZN(n1079) );
OR3_X1 U909 ( .A1(n1240), .A2(n1241), .A3(KEYINPUT54), .ZN(n1249) );
NAND2_X1 U910 ( .A1(KEYINPUT54), .A2(n1100), .ZN(n1248) );
AND3_X1 U911 ( .A1(n1250), .A2(n1058), .A3(n1102), .ZN(n1234) );
XNOR2_X1 U912 ( .A(n1251), .B(n1209), .ZN(G21) );
AND3_X1 U913 ( .A1(n1217), .A2(n1102), .A3(n1215), .ZN(n1209) );
AND3_X1 U914 ( .A1(n1241), .A2(n1240), .A3(n1088), .ZN(n1217) );
XOR2_X1 U915 ( .A(n1252), .B(n1253), .Z(G18) );
XNOR2_X1 U916 ( .A(G116), .B(KEYINPUT11), .ZN(n1253) );
NAND2_X1 U917 ( .A1(n1254), .A2(n1102), .ZN(n1252) );
XOR2_X1 U918 ( .A(n1213), .B(KEYINPUT48), .Z(n1254) );
NAND3_X1 U919 ( .A1(n1087), .A2(n1100), .A3(n1215), .ZN(n1213) );
INV_X1 U920 ( .A(n1255), .ZN(n1215) );
NOR2_X1 U921 ( .A1(n1250), .A2(n1256), .ZN(n1087) );
XOR2_X1 U922 ( .A(G113), .B(n1257), .Z(G15) );
NOR3_X1 U923 ( .A1(n1255), .A2(n1258), .A3(n1239), .ZN(n1257) );
NAND2_X1 U924 ( .A1(n1086), .A2(n1100), .ZN(n1239) );
NOR2_X1 U925 ( .A1(n1240), .A2(n1066), .ZN(n1100) );
INV_X1 U926 ( .A(n1241), .ZN(n1066) );
AND2_X1 U927 ( .A1(n1256), .A2(n1250), .ZN(n1086) );
INV_X1 U928 ( .A(n1058), .ZN(n1256) );
XNOR2_X1 U929 ( .A(n1102), .B(KEYINPUT0), .ZN(n1258) );
NAND2_X1 U930 ( .A1(n1084), .A2(n1219), .ZN(n1255) );
INV_X1 U931 ( .A(n1218), .ZN(n1084) );
NAND3_X1 U932 ( .A1(n1054), .A2(n1093), .A3(n1092), .ZN(n1218) );
XNOR2_X1 U933 ( .A(G110), .B(n1205), .ZN(G12) );
NAND3_X1 U934 ( .A1(n1088), .A2(n1208), .A3(n1099), .ZN(n1205) );
AND2_X1 U935 ( .A1(n1259), .A2(n1240), .ZN(n1099) );
OR2_X1 U936 ( .A1(n1073), .A2(n1260), .ZN(n1240) );
NOR2_X1 U937 ( .A1(n1061), .A2(n1062), .ZN(n1260) );
INV_X1 U938 ( .A(n1261), .ZN(n1062) );
NOR2_X1 U939 ( .A1(n1261), .A2(n1141), .ZN(n1073) );
INV_X1 U940 ( .A(n1061), .ZN(n1141) );
NAND2_X1 U941 ( .A1(G217), .A2(n1262), .ZN(n1061) );
NAND2_X1 U942 ( .A1(n1139), .A2(n1201), .ZN(n1261) );
XOR2_X1 U943 ( .A(n1263), .B(n1264), .Z(n1139) );
XOR2_X1 U944 ( .A(n1265), .B(n1266), .Z(n1264) );
XNOR2_X1 U945 ( .A(n1267), .B(n1268), .ZN(n1266) );
NOR2_X1 U946 ( .A1(KEYINPUT42), .A2(n1269), .ZN(n1268) );
XNOR2_X1 U947 ( .A(G146), .B(KEYINPUT50), .ZN(n1269) );
XNOR2_X1 U948 ( .A(KEYINPUT53), .B(n1123), .ZN(n1265) );
XOR2_X1 U949 ( .A(n1270), .B(n1118), .Z(n1263) );
XOR2_X1 U950 ( .A(n1271), .B(n1272), .Z(n1270) );
AND3_X1 U951 ( .A1(G221), .A2(n1052), .A3(G234), .ZN(n1272) );
NAND2_X1 U952 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
NAND2_X1 U953 ( .A1(G119), .A2(n1275), .ZN(n1274) );
XOR2_X1 U954 ( .A(KEYINPUT6), .B(n1276), .Z(n1273) );
NOR2_X1 U955 ( .A1(G119), .A2(n1275), .ZN(n1276) );
XNOR2_X1 U956 ( .A(KEYINPUT54), .B(n1241), .ZN(n1259) );
XNOR2_X1 U957 ( .A(n1277), .B(G472), .ZN(n1241) );
NAND2_X1 U958 ( .A1(n1278), .A2(n1201), .ZN(n1277) );
XOR2_X1 U959 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U960 ( .A(n1165), .B(n1161), .Z(n1280) );
XNOR2_X1 U961 ( .A(n1281), .B(n1282), .ZN(n1161) );
XNOR2_X1 U962 ( .A(n1283), .B(n1284), .ZN(n1165) );
NOR2_X1 U963 ( .A1(G119), .A2(KEYINPUT51), .ZN(n1284) );
XOR2_X1 U964 ( .A(n1159), .B(n1285), .Z(n1279) );
XOR2_X1 U965 ( .A(KEYINPUT46), .B(G101), .Z(n1285) );
NAND2_X1 U966 ( .A1(n1286), .A2(G210), .ZN(n1159) );
AND3_X1 U967 ( .A1(n1235), .A2(n1219), .A3(n1102), .ZN(n1208) );
NOR2_X1 U968 ( .A1(n1080), .A2(n1101), .ZN(n1102) );
INV_X1 U969 ( .A(n1053), .ZN(n1101) );
NAND2_X1 U970 ( .A1(G214), .A2(n1287), .ZN(n1053) );
XOR2_X1 U971 ( .A(n1067), .B(KEYINPUT18), .Z(n1080) );
XOR2_X1 U972 ( .A(n1288), .B(n1200), .Z(n1067) );
NAND2_X1 U973 ( .A1(G210), .A2(n1287), .ZN(n1200) );
NAND2_X1 U974 ( .A1(n1289), .A2(n1201), .ZN(n1287) );
INV_X1 U975 ( .A(G237), .ZN(n1289) );
NAND2_X1 U976 ( .A1(n1290), .A2(n1201), .ZN(n1288) );
XNOR2_X1 U977 ( .A(n1291), .B(n1292), .ZN(n1290) );
INV_X1 U978 ( .A(n1135), .ZN(n1292) );
XNOR2_X1 U979 ( .A(n1293), .B(n1294), .ZN(n1135) );
XOR2_X1 U980 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U981 ( .A(n1267), .B(G101), .ZN(n1296) );
XNOR2_X1 U982 ( .A(KEYINPUT32), .B(n1297), .ZN(n1295) );
XNOR2_X1 U983 ( .A(n1298), .B(n1299), .ZN(n1293) );
XOR2_X1 U984 ( .A(n1300), .B(n1283), .Z(n1299) );
XNOR2_X1 U985 ( .A(G113), .B(n1301), .ZN(n1283) );
NOR2_X1 U986 ( .A1(KEYINPUT13), .A2(n1251), .ZN(n1300) );
INV_X1 U987 ( .A(G119), .ZN(n1251) );
XNOR2_X1 U988 ( .A(KEYINPUT59), .B(n1302), .ZN(n1291) );
NOR2_X1 U989 ( .A1(KEYINPUT22), .A2(n1303), .ZN(n1302) );
XOR2_X1 U990 ( .A(n1304), .B(KEYINPUT14), .Z(n1303) );
NAND2_X1 U991 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND3_X1 U992 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1306) );
XNOR2_X1 U993 ( .A(KEYINPUT52), .B(n1197), .ZN(n1309) );
NAND2_X1 U994 ( .A1(G125), .A2(n1281), .ZN(n1308) );
XNOR2_X1 U995 ( .A(n1310), .B(n1311), .ZN(n1307) );
NAND3_X1 U996 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(n1305) );
XOR2_X1 U997 ( .A(KEYINPUT52), .B(n1197), .Z(n1314) );
NOR2_X1 U998 ( .A1(n1128), .A2(G953), .ZN(n1197) );
INV_X1 U999 ( .A(G224), .ZN(n1128) );
NAND2_X1 U1000 ( .A1(n1311), .A2(n1310), .ZN(n1313) );
INV_X1 U1001 ( .A(KEYINPUT43), .ZN(n1310) );
NAND2_X1 U1002 ( .A1(n1198), .A2(KEYINPUT43), .ZN(n1312) );
NOR2_X1 U1003 ( .A1(n1311), .A2(n1315), .ZN(n1198) );
AND2_X1 U1004 ( .A1(G125), .A2(n1281), .ZN(n1315) );
NOR2_X1 U1005 ( .A1(n1281), .A2(G125), .ZN(n1311) );
NAND3_X1 U1006 ( .A1(n1316), .A2(n1317), .A3(n1318), .ZN(n1281) );
NAND2_X1 U1007 ( .A1(n1319), .A2(n1275), .ZN(n1318) );
NAND2_X1 U1008 ( .A1(KEYINPUT61), .A2(n1320), .ZN(n1317) );
NAND2_X1 U1009 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
INV_X1 U1010 ( .A(n1319), .ZN(n1322) );
XNOR2_X1 U1011 ( .A(KEYINPUT27), .B(n1275), .ZN(n1321) );
NAND2_X1 U1012 ( .A1(n1323), .A2(n1324), .ZN(n1316) );
INV_X1 U1013 ( .A(KEYINPUT61), .ZN(n1324) );
NAND2_X1 U1014 ( .A1(n1325), .A2(n1326), .ZN(n1323) );
NAND2_X1 U1015 ( .A1(KEYINPUT27), .A2(n1275), .ZN(n1326) );
OR3_X1 U1016 ( .A1(n1319), .A2(KEYINPUT27), .A3(n1275), .ZN(n1325) );
XOR2_X1 U1017 ( .A(G143), .B(n1327), .Z(n1319) );
INV_X1 U1018 ( .A(G146), .ZN(n1327) );
NAND2_X1 U1019 ( .A1(n1103), .A2(n1328), .ZN(n1219) );
NAND2_X1 U1020 ( .A1(n1246), .A2(n1129), .ZN(n1328) );
INV_X1 U1021 ( .A(G898), .ZN(n1129) );
AND3_X1 U1022 ( .A1(G953), .A2(n1329), .A3(n1330), .ZN(n1246) );
XNOR2_X1 U1023 ( .A(G902), .B(KEYINPUT7), .ZN(n1330) );
NAND3_X1 U1024 ( .A1(n1329), .A2(n1052), .A3(G952), .ZN(n1103) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1329) );
INV_X1 U1026 ( .A(n1090), .ZN(n1235) );
NAND2_X1 U1027 ( .A1(n1093), .A2(n1331), .ZN(n1090) );
NAND2_X1 U1028 ( .A1(n1092), .A2(n1054), .ZN(n1331) );
NAND3_X1 U1029 ( .A1(n1192), .A2(n1201), .A3(n1332), .ZN(n1054) );
INV_X1 U1030 ( .A(G469), .ZN(n1192) );
XNOR2_X1 U1031 ( .A(n1072), .B(KEYINPUT28), .ZN(n1092) );
AND2_X1 U1032 ( .A1(G469), .A2(n1333), .ZN(n1072) );
NAND2_X1 U1033 ( .A1(n1332), .A2(n1201), .ZN(n1333) );
XNOR2_X1 U1034 ( .A(n1334), .B(n1335), .ZN(n1332) );
XNOR2_X1 U1035 ( .A(KEYINPUT35), .B(n1176), .ZN(n1335) );
NAND2_X1 U1036 ( .A1(G227), .A2(n1052), .ZN(n1176) );
XOR2_X1 U1037 ( .A(n1190), .B(n1336), .Z(n1334) );
NOR2_X1 U1038 ( .A1(n1186), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1039 ( .A(n1185), .B(KEYINPUT30), .Z(n1337) );
NAND2_X1 U1040 ( .A1(n1189), .A2(n1267), .ZN(n1185) );
NOR2_X1 U1041 ( .A1(n1189), .A2(n1267), .ZN(n1186) );
INV_X1 U1042 ( .A(G110), .ZN(n1267) );
XOR2_X1 U1043 ( .A(G140), .B(KEYINPUT17), .Z(n1189) );
XNOR2_X1 U1044 ( .A(n1338), .B(n1339), .ZN(n1190) );
INV_X1 U1045 ( .A(n1117), .ZN(n1339) );
XOR2_X1 U1046 ( .A(G146), .B(n1340), .Z(n1117) );
XOR2_X1 U1047 ( .A(n1341), .B(n1282), .Z(n1338) );
XNOR2_X1 U1048 ( .A(n1123), .B(n1122), .ZN(n1282) );
XOR2_X1 U1049 ( .A(G131), .B(G134), .Z(n1122) );
INV_X1 U1050 ( .A(G137), .ZN(n1123) );
NAND2_X1 U1051 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NAND2_X1 U1052 ( .A1(G101), .A2(n1298), .ZN(n1343) );
XOR2_X1 U1053 ( .A(KEYINPUT20), .B(n1344), .Z(n1342) );
NOR2_X1 U1054 ( .A1(G101), .A2(n1298), .ZN(n1344) );
XOR2_X1 U1055 ( .A(G104), .B(G107), .Z(n1298) );
NAND2_X1 U1056 ( .A1(G221), .A2(n1262), .ZN(n1093) );
NAND2_X1 U1057 ( .A1(G234), .A2(n1201), .ZN(n1262) );
INV_X1 U1058 ( .A(G902), .ZN(n1201) );
NOR2_X1 U1059 ( .A1(n1058), .A2(n1250), .ZN(n1088) );
XNOR2_X1 U1060 ( .A(n1069), .B(n1071), .ZN(n1250) );
INV_X1 U1061 ( .A(G475), .ZN(n1071) );
NOR2_X1 U1062 ( .A1(n1150), .A2(G902), .ZN(n1069) );
XOR2_X1 U1063 ( .A(n1345), .B(n1346), .Z(n1150) );
XOR2_X1 U1064 ( .A(G104), .B(n1347), .Z(n1346) );
XOR2_X1 U1065 ( .A(G131), .B(G113), .Z(n1347) );
XOR2_X1 U1066 ( .A(n1348), .B(n1349), .Z(n1345) );
XOR2_X1 U1067 ( .A(n1350), .B(n1351), .Z(n1349) );
NAND3_X1 U1068 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1351) );
OR2_X1 U1069 ( .A1(n1118), .A2(KEYINPUT19), .ZN(n1354) );
NAND3_X1 U1070 ( .A1(KEYINPUT19), .A2(n1118), .A3(n1355), .ZN(n1353) );
NAND2_X1 U1071 ( .A1(n1356), .A2(n1357), .ZN(n1352) );
NAND2_X1 U1072 ( .A1(n1358), .A2(KEYINPUT19), .ZN(n1357) );
XNOR2_X1 U1073 ( .A(n1118), .B(KEYINPUT12), .ZN(n1358) );
XOR2_X1 U1074 ( .A(G140), .B(G125), .Z(n1118) );
INV_X1 U1075 ( .A(n1355), .ZN(n1356) );
XOR2_X1 U1076 ( .A(G146), .B(KEYINPUT24), .Z(n1355) );
NAND2_X1 U1077 ( .A1(n1359), .A2(KEYINPUT23), .ZN(n1350) );
XOR2_X1 U1078 ( .A(n1360), .B(G143), .Z(n1359) );
NAND2_X1 U1079 ( .A1(n1286), .A2(G214), .ZN(n1360) );
NOR2_X1 U1080 ( .A1(G953), .A2(G237), .ZN(n1286) );
NAND2_X1 U1081 ( .A1(KEYINPUT45), .A2(n1297), .ZN(n1348) );
XOR2_X1 U1082 ( .A(G478), .B(n1361), .Z(n1058) );
NOR2_X1 U1083 ( .A1(G902), .A2(n1145), .ZN(n1361) );
NAND2_X1 U1084 ( .A1(n1362), .A2(n1363), .ZN(n1145) );
NAND2_X1 U1085 ( .A1(n1364), .A2(n1365), .ZN(n1363) );
NAND2_X1 U1086 ( .A1(n1366), .A2(n1367), .ZN(n1365) );
NAND4_X1 U1087 ( .A1(KEYINPUT33), .A2(G217), .A3(G234), .A4(n1052), .ZN(n1367) );
XNOR2_X1 U1088 ( .A(KEYINPUT29), .B(n1368), .ZN(n1364) );
NAND2_X1 U1089 ( .A1(n1369), .A2(n1370), .ZN(n1362) );
NAND3_X1 U1090 ( .A1(G234), .A2(n1052), .A3(G217), .ZN(n1370) );
INV_X1 U1091 ( .A(G953), .ZN(n1052) );
NAND2_X1 U1092 ( .A1(n1366), .A2(KEYINPUT33), .ZN(n1369) );
XNOR2_X1 U1093 ( .A(n1371), .B(KEYINPUT37), .ZN(n1366) );
INV_X1 U1094 ( .A(n1368), .ZN(n1371) );
NAND2_X1 U1095 ( .A1(n1372), .A2(n1373), .ZN(n1368) );
NAND2_X1 U1096 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
XNOR2_X1 U1097 ( .A(n1376), .B(n1377), .ZN(n1375) );
XOR2_X1 U1098 ( .A(G134), .B(n1340), .Z(n1374) );
XOR2_X1 U1099 ( .A(n1378), .B(KEYINPUT26), .Z(n1372) );
NAND2_X1 U1100 ( .A1(n1379), .A2(n1380), .ZN(n1378) );
XOR2_X1 U1101 ( .A(n1376), .B(n1377), .Z(n1380) );
XNOR2_X1 U1102 ( .A(G107), .B(n1297), .ZN(n1377) );
INV_X1 U1103 ( .A(G122), .ZN(n1297) );
NAND2_X1 U1104 ( .A1(KEYINPUT25), .A2(n1301), .ZN(n1376) );
INV_X1 U1105 ( .A(G116), .ZN(n1301) );
XNOR2_X1 U1106 ( .A(G134), .B(n1340), .ZN(n1379) );
XNOR2_X1 U1107 ( .A(G143), .B(n1275), .ZN(n1340) );
INV_X1 U1108 ( .A(G128), .ZN(n1275) );
endmodule


