//Key = 0001110110001011110100000111010101101110100110000100101001001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348;

XOR2_X1 U738 ( .A(G107), .B(n1032), .Z(G9) );
NOR2_X1 U739 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR2_X1 U740 ( .A1(n1035), .A2(n1036), .ZN(G75) );
NOR4_X1 U741 ( .A1(n1037), .A2(n1038), .A3(G953), .A4(n1039), .ZN(n1036) );
NOR4_X1 U742 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1038) );
NAND3_X1 U743 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1040) );
OR2_X1 U744 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND3_X1 U745 ( .A1(n1034), .A2(n1049), .A3(n1047), .ZN(n1044) );
NAND2_X1 U746 ( .A1(n1050), .A2(n1051), .ZN(n1037) );
NAND3_X1 U747 ( .A1(n1046), .A2(n1052), .A3(n1048), .ZN(n1051) );
NAND2_X1 U748 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND3_X1 U749 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NAND2_X1 U750 ( .A1(n1058), .A2(n1059), .ZN(n1053) );
NAND2_X1 U751 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U752 ( .A1(n1055), .A2(n1062), .ZN(n1061) );
NAND2_X1 U753 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U754 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U755 ( .A1(n1056), .A2(n1067), .ZN(n1060) );
NAND2_X1 U756 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND3_X1 U757 ( .A1(G214), .A2(n1070), .A3(n1071), .ZN(n1069) );
INV_X1 U758 ( .A(n1072), .ZN(n1046) );
NOR3_X1 U759 ( .A1(n1039), .A2(G953), .A3(G952), .ZN(n1035) );
AND4_X1 U760 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1039) );
NOR3_X1 U761 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1076) );
NOR2_X1 U762 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
INV_X1 U763 ( .A(n1082), .ZN(n1078) );
XNOR2_X1 U764 ( .A(n1083), .B(n1084), .ZN(n1077) );
XOR2_X1 U765 ( .A(KEYINPUT52), .B(G472), .Z(n1084) );
XNOR2_X1 U766 ( .A(n1085), .B(n1086), .ZN(n1075) );
XNOR2_X1 U767 ( .A(KEYINPUT56), .B(KEYINPUT55), .ZN(n1085) );
XOR2_X1 U768 ( .A(KEYINPUT18), .B(n1087), .Z(n1074) );
NOR3_X1 U769 ( .A1(n1088), .A2(n1089), .A3(n1043), .ZN(n1087) );
XNOR2_X1 U770 ( .A(G469), .B(n1090), .ZN(n1088) );
NAND2_X1 U771 ( .A1(n1091), .A2(n1092), .ZN(G72) );
NAND2_X1 U772 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U773 ( .A1(KEYINPUT27), .A2(n1095), .ZN(n1093) );
NAND2_X1 U774 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U775 ( .A(n1098), .B(n1099), .Z(n1091) );
NOR3_X1 U776 ( .A1(n1097), .A2(n1100), .A3(n1096), .ZN(n1099) );
XOR2_X1 U777 ( .A(n1101), .B(n1102), .Z(n1096) );
XNOR2_X1 U778 ( .A(n1103), .B(KEYINPUT54), .ZN(n1102) );
NAND3_X1 U779 ( .A1(n1104), .A2(n1105), .A3(KEYINPUT14), .ZN(n1103) );
NAND2_X1 U780 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U781 ( .A(n1108), .B(n1109), .Z(n1106) );
OR3_X1 U782 ( .A1(n1109), .A2(n1108), .A3(n1107), .ZN(n1104) );
INV_X1 U783 ( .A(KEYINPUT6), .ZN(n1107) );
XOR2_X1 U784 ( .A(G131), .B(KEYINPUT43), .Z(n1109) );
XNOR2_X1 U785 ( .A(n1110), .B(n1111), .ZN(n1101) );
NAND2_X1 U786 ( .A1(n1112), .A2(KEYINPUT27), .ZN(n1098) );
INV_X1 U787 ( .A(n1094), .ZN(n1112) );
NAND2_X1 U788 ( .A1(G953), .A2(n1113), .ZN(n1094) );
NAND2_X1 U789 ( .A1(G900), .A2(G227), .ZN(n1113) );
XOR2_X1 U790 ( .A(n1114), .B(n1115), .Z(G69) );
XOR2_X1 U791 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U792 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U793 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
NAND2_X1 U794 ( .A1(n1122), .A2(n1123), .ZN(n1116) );
NAND2_X1 U795 ( .A1(G953), .A2(n1121), .ZN(n1123) );
XOR2_X1 U796 ( .A(n1124), .B(n1125), .Z(n1122) );
NAND2_X1 U797 ( .A1(n1119), .A2(n1126), .ZN(n1114) );
NOR2_X1 U798 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XOR2_X1 U799 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U800 ( .A1(n1081), .A2(n1131), .ZN(n1130) );
INV_X1 U801 ( .A(n1132), .ZN(n1131) );
NAND2_X1 U802 ( .A1(KEYINPUT38), .A2(n1133), .ZN(n1129) );
NOR3_X1 U803 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(G63) );
AND3_X1 U804 ( .A1(KEYINPUT2), .A2(G953), .A3(G952), .ZN(n1136) );
NOR2_X1 U805 ( .A1(KEYINPUT2), .A2(n1137), .ZN(n1135) );
INV_X1 U806 ( .A(n1127), .ZN(n1137) );
XOR2_X1 U807 ( .A(n1138), .B(n1139), .Z(n1134) );
NAND2_X1 U808 ( .A1(n1132), .A2(G478), .ZN(n1138) );
NOR2_X1 U809 ( .A1(n1127), .A2(n1140), .ZN(G60) );
XOR2_X1 U810 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U811 ( .A1(n1132), .A2(G475), .ZN(n1141) );
XOR2_X1 U812 ( .A(G104), .B(n1143), .Z(G6) );
NOR2_X1 U813 ( .A1(n1127), .A2(n1144), .ZN(G57) );
XOR2_X1 U814 ( .A(n1145), .B(n1146), .Z(n1144) );
XNOR2_X1 U815 ( .A(n1147), .B(n1148), .ZN(n1146) );
XNOR2_X1 U816 ( .A(n1149), .B(n1150), .ZN(n1148) );
NAND3_X1 U817 ( .A1(n1151), .A2(n1152), .A3(G472), .ZN(n1149) );
OR2_X1 U818 ( .A1(n1132), .A2(KEYINPUT10), .ZN(n1152) );
NAND2_X1 U819 ( .A1(KEYINPUT10), .A2(n1153), .ZN(n1151) );
NAND2_X1 U820 ( .A1(n1050), .A2(G902), .ZN(n1153) );
XOR2_X1 U821 ( .A(n1154), .B(n1155), .Z(n1145) );
XOR2_X1 U822 ( .A(KEYINPUT32), .B(KEYINPUT26), .Z(n1155) );
XOR2_X1 U823 ( .A(n1156), .B(n1157), .Z(n1154) );
NOR2_X1 U824 ( .A1(KEYINPUT45), .A2(n1158), .ZN(n1157) );
XNOR2_X1 U825 ( .A(n1159), .B(n1160), .ZN(n1158) );
NOR2_X1 U826 ( .A1(n1161), .A2(n1162), .ZN(n1159) );
AND2_X1 U827 ( .A1(KEYINPUT53), .A2(n1163), .ZN(n1162) );
NOR2_X1 U828 ( .A1(KEYINPUT11), .A2(n1163), .ZN(n1161) );
NOR2_X1 U829 ( .A1(n1127), .A2(n1164), .ZN(G54) );
XOR2_X1 U830 ( .A(n1165), .B(n1166), .Z(n1164) );
XNOR2_X1 U831 ( .A(n1167), .B(n1168), .ZN(n1166) );
XNOR2_X1 U832 ( .A(n1169), .B(n1170), .ZN(n1168) );
NAND2_X1 U833 ( .A1(KEYINPUT34), .A2(n1171), .ZN(n1169) );
XOR2_X1 U834 ( .A(n1172), .B(n1173), .Z(n1165) );
XOR2_X1 U835 ( .A(KEYINPUT17), .B(n1174), .Z(n1173) );
NOR3_X1 U836 ( .A1(n1175), .A2(KEYINPUT30), .A3(n1176), .ZN(n1174) );
NOR2_X1 U837 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XNOR2_X1 U838 ( .A(KEYINPUT51), .B(n1179), .ZN(n1178) );
NOR2_X1 U839 ( .A1(n1180), .A2(G110), .ZN(n1177) );
NOR2_X1 U840 ( .A1(G140), .A2(n1181), .ZN(n1180) );
NOR2_X1 U841 ( .A1(n1182), .A2(n1183), .ZN(n1175) );
NOR2_X1 U842 ( .A1(G110), .A2(n1181), .ZN(n1182) );
INV_X1 U843 ( .A(KEYINPUT36), .ZN(n1181) );
XNOR2_X1 U844 ( .A(n1184), .B(n1185), .ZN(n1172) );
NAND2_X1 U845 ( .A1(n1132), .A2(G469), .ZN(n1184) );
NOR2_X1 U846 ( .A1(n1127), .A2(n1186), .ZN(G51) );
XOR2_X1 U847 ( .A(n1187), .B(n1188), .Z(n1186) );
XNOR2_X1 U848 ( .A(n1189), .B(n1190), .ZN(n1188) );
NAND2_X1 U849 ( .A1(KEYINPUT29), .A2(n1160), .ZN(n1189) );
XNOR2_X1 U850 ( .A(n1191), .B(n1192), .ZN(n1187) );
NAND2_X1 U851 ( .A1(n1132), .A2(G210), .ZN(n1191) );
NOR2_X1 U852 ( .A1(n1193), .A2(n1050), .ZN(n1132) );
NOR2_X1 U853 ( .A1(n1126), .A2(n1097), .ZN(n1050) );
NAND2_X1 U854 ( .A1(n1194), .A2(n1195), .ZN(n1097) );
NOR4_X1 U855 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1195) );
NOR4_X1 U856 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1194) );
NOR2_X1 U857 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NOR3_X1 U858 ( .A1(n1206), .A2(n1034), .A3(n1043), .ZN(n1202) );
NAND4_X1 U859 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1126) );
NOR4_X1 U860 ( .A1(n1211), .A2(n1143), .A3(n1212), .A4(n1213), .ZN(n1210) );
NOR4_X1 U861 ( .A1(n1214), .A2(n1215), .A3(n1042), .A4(n1034), .ZN(n1213) );
INV_X1 U862 ( .A(n1056), .ZN(n1042) );
NOR2_X1 U863 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
INV_X1 U864 ( .A(KEYINPUT47), .ZN(n1217) );
NOR3_X1 U865 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1216) );
INV_X1 U866 ( .A(n1221), .ZN(n1219) );
NOR2_X1 U867 ( .A1(KEYINPUT47), .A2(n1222), .ZN(n1214) );
NOR2_X1 U868 ( .A1(n1063), .A2(n1223), .ZN(n1212) );
INV_X1 U869 ( .A(n1224), .ZN(n1063) );
NOR2_X1 U870 ( .A1(n1049), .A2(n1033), .ZN(n1143) );
NAND2_X1 U871 ( .A1(n1222), .A2(n1056), .ZN(n1033) );
NOR2_X1 U872 ( .A1(n1225), .A2(n1226), .ZN(n1209) );
NOR2_X1 U873 ( .A1(n1119), .A2(G952), .ZN(n1127) );
XNOR2_X1 U874 ( .A(n1227), .B(n1228), .ZN(G48) );
NOR2_X1 U875 ( .A1(n1229), .A2(n1205), .ZN(n1228) );
NAND3_X1 U876 ( .A1(n1230), .A2(n1231), .A3(n1057), .ZN(n1205) );
XNOR2_X1 U877 ( .A(n1204), .B(KEYINPUT40), .ZN(n1229) );
XOR2_X1 U878 ( .A(G143), .B(n1199), .Z(G45) );
NOR4_X1 U879 ( .A1(n1206), .A2(n1068), .A3(n1086), .A4(n1073), .ZN(n1199) );
XNOR2_X1 U880 ( .A(n1183), .B(n1201), .ZN(G42) );
AND3_X1 U881 ( .A1(n1231), .A2(n1065), .A3(n1232), .ZN(n1201) );
XOR2_X1 U882 ( .A(G137), .B(n1200), .Z(G39) );
AND3_X1 U883 ( .A1(n1233), .A2(n1048), .A3(n1232), .ZN(n1200) );
AND4_X1 U884 ( .A1(n1057), .A2(n1055), .A3(n1234), .A4(n1066), .ZN(n1232) );
XOR2_X1 U885 ( .A(n1235), .B(n1236), .Z(G36) );
XOR2_X1 U886 ( .A(KEYINPUT42), .B(G134), .Z(n1236) );
NOR3_X1 U887 ( .A1(n1206), .A2(n1237), .A3(n1034), .ZN(n1235) );
INV_X1 U888 ( .A(n1238), .ZN(n1034) );
XNOR2_X1 U889 ( .A(n1055), .B(KEYINPUT28), .ZN(n1237) );
INV_X1 U890 ( .A(n1043), .ZN(n1055) );
NAND2_X1 U891 ( .A1(n1239), .A2(n1240), .ZN(G33) );
NAND2_X1 U892 ( .A1(n1198), .A2(n1241), .ZN(n1240) );
XOR2_X1 U893 ( .A(KEYINPUT5), .B(n1242), .Z(n1239) );
NOR2_X1 U894 ( .A1(n1198), .A2(n1241), .ZN(n1242) );
NOR3_X1 U895 ( .A1(n1049), .A2(n1043), .A3(n1206), .ZN(n1198) );
NAND3_X1 U896 ( .A1(n1224), .A2(n1234), .A3(n1057), .ZN(n1206) );
XNOR2_X1 U897 ( .A(n1243), .B(KEYINPUT37), .ZN(n1057) );
NAND2_X1 U898 ( .A1(n1071), .A2(n1244), .ZN(n1043) );
INV_X1 U899 ( .A(n1245), .ZN(n1071) );
INV_X1 U900 ( .A(n1231), .ZN(n1049) );
XOR2_X1 U901 ( .A(G128), .B(n1197), .Z(G30) );
AND4_X1 U902 ( .A1(n1230), .A2(n1238), .A3(n1243), .A4(n1234), .ZN(n1197) );
NOR3_X1 U903 ( .A1(n1068), .A2(n1246), .A3(n1065), .ZN(n1230) );
XOR2_X1 U904 ( .A(G101), .B(n1211), .Z(G3) );
AND3_X1 U905 ( .A1(n1048), .A2(n1222), .A3(n1224), .ZN(n1211) );
XOR2_X1 U906 ( .A(n1196), .B(n1247), .Z(G27) );
NOR2_X1 U907 ( .A1(KEYINPUT58), .A2(n1192), .ZN(n1247) );
AND4_X1 U908 ( .A1(n1058), .A2(n1248), .A3(n1231), .A4(n1249), .ZN(n1196) );
NOR3_X1 U909 ( .A1(n1233), .A2(n1246), .A3(n1204), .ZN(n1249) );
INV_X1 U910 ( .A(n1234), .ZN(n1204) );
NAND2_X1 U911 ( .A1(n1072), .A2(n1250), .ZN(n1234) );
NAND3_X1 U912 ( .A1(G902), .A2(n1251), .A3(n1100), .ZN(n1250) );
NOR2_X1 U913 ( .A1(n1119), .A2(G900), .ZN(n1100) );
INV_X1 U914 ( .A(n1066), .ZN(n1246) );
XOR2_X1 U915 ( .A(G122), .B(n1226), .Z(G24) );
AND4_X1 U916 ( .A1(n1252), .A2(n1056), .A3(n1253), .A4(n1254), .ZN(n1226) );
NOR2_X1 U917 ( .A1(n1066), .A2(n1233), .ZN(n1056) );
XNOR2_X1 U918 ( .A(n1225), .B(n1255), .ZN(G21) );
NAND2_X1 U919 ( .A1(KEYINPUT16), .A2(n1256), .ZN(n1255) );
XOR2_X1 U920 ( .A(KEYINPUT22), .B(G119), .Z(n1256) );
AND4_X1 U921 ( .A1(n1233), .A2(n1252), .A3(n1048), .A4(n1066), .ZN(n1225) );
INV_X1 U922 ( .A(n1065), .ZN(n1233) );
XNOR2_X1 U923 ( .A(G116), .B(n1207), .ZN(G18) );
NAND3_X1 U924 ( .A1(n1252), .A2(n1238), .A3(n1224), .ZN(n1207) );
NOR2_X1 U925 ( .A1(n1254), .A2(n1086), .ZN(n1238) );
INV_X1 U926 ( .A(n1253), .ZN(n1086) );
AND3_X1 U927 ( .A1(n1248), .A2(n1218), .A3(n1058), .ZN(n1252) );
XNOR2_X1 U928 ( .A(G113), .B(n1257), .ZN(G15) );
NAND3_X1 U929 ( .A1(KEYINPUT15), .A2(n1258), .A3(n1259), .ZN(n1257) );
XNOR2_X1 U930 ( .A(n1224), .B(KEYINPUT4), .ZN(n1259) );
NOR2_X1 U931 ( .A1(n1065), .A2(n1066), .ZN(n1224) );
INV_X1 U932 ( .A(n1223), .ZN(n1258) );
NAND4_X1 U933 ( .A1(n1231), .A2(n1058), .A3(n1221), .A4(n1218), .ZN(n1223) );
NOR2_X1 U934 ( .A1(n1041), .A2(n1089), .ZN(n1058) );
INV_X1 U935 ( .A(n1047), .ZN(n1089) );
NOR2_X1 U936 ( .A1(n1253), .A2(n1073), .ZN(n1231) );
INV_X1 U937 ( .A(n1254), .ZN(n1073) );
XNOR2_X1 U938 ( .A(G110), .B(n1208), .ZN(G12) );
NAND4_X1 U939 ( .A1(n1048), .A2(n1222), .A3(n1065), .A4(n1066), .ZN(n1208) );
NAND3_X1 U940 ( .A1(n1260), .A2(n1261), .A3(n1082), .ZN(n1066) );
NAND2_X1 U941 ( .A1(n1080), .A2(n1081), .ZN(n1082) );
NAND2_X1 U942 ( .A1(n1081), .A2(n1262), .ZN(n1261) );
OR3_X1 U943 ( .A1(n1081), .A2(n1080), .A3(n1262), .ZN(n1260) );
INV_X1 U944 ( .A(KEYINPUT31), .ZN(n1262) );
AND2_X1 U945 ( .A1(n1133), .A2(n1193), .ZN(n1080) );
XNOR2_X1 U946 ( .A(n1263), .B(n1264), .ZN(n1133) );
XNOR2_X1 U947 ( .A(n1265), .B(n1266), .ZN(n1264) );
NOR2_X1 U948 ( .A1(KEYINPUT35), .A2(n1267), .ZN(n1266) );
XOR2_X1 U949 ( .A(n1268), .B(n1269), .Z(n1267) );
NAND2_X1 U950 ( .A1(G221), .A2(n1270), .ZN(n1268) );
NAND2_X1 U951 ( .A1(KEYINPUT25), .A2(n1271), .ZN(n1265) );
XNOR2_X1 U952 ( .A(KEYINPUT3), .B(n1227), .ZN(n1271) );
XOR2_X1 U953 ( .A(n1272), .B(n1111), .Z(n1263) );
NAND2_X1 U954 ( .A1(KEYINPUT44), .A2(n1273), .ZN(n1272) );
XOR2_X1 U955 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U956 ( .A(G119), .B(n1179), .ZN(n1275) );
INV_X1 U957 ( .A(G110), .ZN(n1179) );
NAND2_X1 U958 ( .A1(G217), .A2(n1276), .ZN(n1081) );
XOR2_X1 U959 ( .A(G472), .B(n1277), .Z(n1065) );
NOR2_X1 U960 ( .A1(n1083), .A2(KEYINPUT46), .ZN(n1277) );
AND2_X1 U961 ( .A1(n1278), .A2(n1193), .ZN(n1083) );
XOR2_X1 U962 ( .A(n1279), .B(n1280), .Z(n1278) );
XNOR2_X1 U963 ( .A(n1150), .B(n1147), .ZN(n1280) );
XOR2_X1 U964 ( .A(n1156), .B(n1281), .Z(n1279) );
NOR2_X1 U965 ( .A1(KEYINPUT59), .A2(n1282), .ZN(n1281) );
XNOR2_X1 U966 ( .A(n1160), .B(n1163), .ZN(n1282) );
NAND3_X1 U967 ( .A1(n1283), .A2(n1119), .A3(G210), .ZN(n1156) );
AND3_X1 U968 ( .A1(n1221), .A2(n1218), .A3(n1243), .ZN(n1222) );
INV_X1 U969 ( .A(n1220), .ZN(n1243) );
NAND2_X1 U970 ( .A1(n1047), .A2(n1041), .ZN(n1220) );
NAND3_X1 U971 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1041) );
NAND2_X1 U972 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
INV_X1 U973 ( .A(G469), .ZN(n1288) );
NAND2_X1 U974 ( .A1(n1289), .A2(KEYINPUT7), .ZN(n1287) );
XOR2_X1 U975 ( .A(n1090), .B(KEYINPUT24), .Z(n1289) );
NAND3_X1 U976 ( .A1(KEYINPUT7), .A2(G469), .A3(n1090), .ZN(n1285) );
OR2_X1 U977 ( .A1(n1090), .A2(KEYINPUT7), .ZN(n1284) );
NAND3_X1 U978 ( .A1(n1290), .A2(n1291), .A3(n1193), .ZN(n1090) );
NAND3_X1 U979 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n1291) );
INV_X1 U980 ( .A(KEYINPUT12), .ZN(n1294) );
NAND2_X1 U981 ( .A1(n1295), .A2(KEYINPUT12), .ZN(n1290) );
XOR2_X1 U982 ( .A(n1293), .B(n1292), .Z(n1295) );
XOR2_X1 U983 ( .A(n1296), .B(n1167), .Z(n1292) );
INV_X1 U984 ( .A(n1110), .ZN(n1167) );
XNOR2_X1 U985 ( .A(n1297), .B(n1298), .ZN(n1110) );
XNOR2_X1 U986 ( .A(G146), .B(n1299), .ZN(n1297) );
XNOR2_X1 U987 ( .A(n1300), .B(n1163), .ZN(n1296) );
INV_X1 U988 ( .A(n1170), .ZN(n1163) );
XOR2_X1 U989 ( .A(G131), .B(n1108), .Z(n1170) );
XOR2_X1 U990 ( .A(G134), .B(n1269), .Z(n1108) );
XOR2_X1 U991 ( .A(G137), .B(KEYINPUT62), .Z(n1269) );
NAND2_X1 U992 ( .A1(KEYINPUT49), .A2(n1171), .ZN(n1300) );
XNOR2_X1 U993 ( .A(n1301), .B(n1302), .ZN(n1171) );
XNOR2_X1 U994 ( .A(n1185), .B(n1303), .ZN(n1293) );
XNOR2_X1 U995 ( .A(n1183), .B(G110), .ZN(n1303) );
INV_X1 U996 ( .A(G140), .ZN(n1183) );
NAND2_X1 U997 ( .A1(G227), .A2(n1119), .ZN(n1185) );
NAND2_X1 U998 ( .A1(G221), .A2(n1276), .ZN(n1047) );
NAND2_X1 U999 ( .A1(G234), .A2(n1193), .ZN(n1276) );
NAND2_X1 U1000 ( .A1(n1072), .A2(n1304), .ZN(n1218) );
NAND4_X1 U1001 ( .A1(G953), .A2(G902), .A3(n1251), .A4(n1121), .ZN(n1304) );
INV_X1 U1002 ( .A(G898), .ZN(n1121) );
NAND3_X1 U1003 ( .A1(n1251), .A2(n1119), .A3(G952), .ZN(n1072) );
NAND2_X1 U1004 ( .A1(G237), .A2(G234), .ZN(n1251) );
XOR2_X1 U1005 ( .A(n1248), .B(KEYINPUT21), .Z(n1221) );
INV_X1 U1006 ( .A(n1068), .ZN(n1248) );
NAND2_X1 U1007 ( .A1(n1245), .A2(n1244), .ZN(n1068) );
NAND2_X1 U1008 ( .A1(G214), .A2(n1070), .ZN(n1244) );
NAND2_X1 U1009 ( .A1(n1193), .A2(n1283), .ZN(n1070) );
NAND3_X1 U1010 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1245) );
NAND2_X1 U1011 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
OR3_X1 U1012 ( .A1(n1309), .A2(n1308), .A3(G902), .ZN(n1306) );
AND2_X1 U1013 ( .A1(G210), .A2(G237), .ZN(n1308) );
XOR2_X1 U1014 ( .A(n1310), .B(n1311), .Z(n1309) );
INV_X1 U1015 ( .A(n1190), .ZN(n1311) );
XNOR2_X1 U1016 ( .A(n1312), .B(n1313), .ZN(n1190) );
NOR2_X1 U1017 ( .A1(G953), .A2(n1120), .ZN(n1313) );
INV_X1 U1018 ( .A(G224), .ZN(n1120) );
NAND2_X1 U1019 ( .A1(n1314), .A2(n1315), .ZN(n1312) );
NAND2_X1 U1020 ( .A1(n1125), .A2(n1124), .ZN(n1315) );
XOR2_X1 U1021 ( .A(n1316), .B(KEYINPUT50), .Z(n1314) );
OR2_X1 U1022 ( .A1(n1124), .A2(n1125), .ZN(n1316) );
XOR2_X1 U1023 ( .A(n1317), .B(n1318), .Z(n1125) );
INV_X1 U1024 ( .A(n1319), .ZN(n1318) );
XNOR2_X1 U1025 ( .A(G110), .B(KEYINPUT33), .ZN(n1317) );
XOR2_X1 U1026 ( .A(n1320), .B(n1321), .Z(n1124) );
INV_X1 U1027 ( .A(n1150), .ZN(n1321) );
XNOR2_X1 U1028 ( .A(n1322), .B(n1302), .ZN(n1150) );
XOR2_X1 U1029 ( .A(G101), .B(KEYINPUT60), .Z(n1302) );
XNOR2_X1 U1030 ( .A(G113), .B(G119), .ZN(n1322) );
XNOR2_X1 U1031 ( .A(n1323), .B(n1324), .ZN(n1320) );
NOR2_X1 U1032 ( .A1(KEYINPUT48), .A2(n1147), .ZN(n1324) );
XNOR2_X1 U1033 ( .A(G116), .B(KEYINPUT61), .ZN(n1147) );
NOR2_X1 U1034 ( .A1(KEYINPUT20), .A2(n1301), .ZN(n1323) );
XNOR2_X1 U1035 ( .A(G104), .B(G107), .ZN(n1301) );
XNOR2_X1 U1036 ( .A(n1160), .B(n1192), .ZN(n1310) );
INV_X1 U1037 ( .A(G125), .ZN(n1192) );
XNOR2_X1 U1038 ( .A(n1299), .B(n1325), .ZN(n1160) );
NOR2_X1 U1039 ( .A1(KEYINPUT13), .A2(n1326), .ZN(n1325) );
XNOR2_X1 U1040 ( .A(n1298), .B(n1327), .ZN(n1326) );
NOR2_X1 U1041 ( .A1(G146), .A2(KEYINPUT23), .ZN(n1327) );
XOR2_X1 U1042 ( .A(G143), .B(KEYINPUT57), .Z(n1298) );
XOR2_X1 U1043 ( .A(n1274), .B(KEYINPUT1), .Z(n1299) );
NAND2_X1 U1044 ( .A1(G210), .A2(G902), .ZN(n1305) );
NOR2_X1 U1045 ( .A1(n1253), .A2(n1254), .ZN(n1048) );
XNOR2_X1 U1046 ( .A(n1328), .B(G475), .ZN(n1254) );
NAND2_X1 U1047 ( .A1(n1142), .A2(n1193), .ZN(n1328) );
XNOR2_X1 U1048 ( .A(n1329), .B(n1330), .ZN(n1142) );
XNOR2_X1 U1049 ( .A(n1331), .B(n1332), .ZN(n1330) );
NOR2_X1 U1050 ( .A1(KEYINPUT39), .A2(n1333), .ZN(n1332) );
XOR2_X1 U1051 ( .A(n1334), .B(n1335), .Z(n1333) );
XNOR2_X1 U1052 ( .A(n1111), .B(n1336), .ZN(n1335) );
XOR2_X1 U1053 ( .A(n1337), .B(n1338), .Z(n1336) );
AND3_X1 U1054 ( .A1(G214), .A2(n1119), .A3(n1283), .ZN(n1338) );
INV_X1 U1055 ( .A(G237), .ZN(n1283) );
NAND2_X1 U1056 ( .A1(KEYINPUT8), .A2(n1227), .ZN(n1337) );
INV_X1 U1057 ( .A(G146), .ZN(n1227) );
XOR2_X1 U1058 ( .A(G125), .B(G140), .Z(n1111) );
XNOR2_X1 U1059 ( .A(n1241), .B(n1339), .ZN(n1334) );
XOR2_X1 U1060 ( .A(KEYINPUT19), .B(G143), .Z(n1339) );
INV_X1 U1061 ( .A(G131), .ZN(n1241) );
INV_X1 U1062 ( .A(G113), .ZN(n1331) );
XNOR2_X1 U1063 ( .A(n1319), .B(n1340), .ZN(n1329) );
NOR2_X1 U1064 ( .A1(G104), .A2(KEYINPUT9), .ZN(n1340) );
XNOR2_X1 U1065 ( .A(n1341), .B(G478), .ZN(n1253) );
NAND2_X1 U1066 ( .A1(n1139), .A2(n1193), .ZN(n1341) );
INV_X1 U1067 ( .A(G902), .ZN(n1193) );
XNOR2_X1 U1068 ( .A(n1342), .B(n1343), .ZN(n1139) );
XNOR2_X1 U1069 ( .A(n1319), .B(n1344), .ZN(n1343) );
XOR2_X1 U1070 ( .A(n1345), .B(n1274), .Z(n1344) );
XOR2_X1 U1071 ( .A(G128), .B(KEYINPUT41), .Z(n1274) );
NAND2_X1 U1072 ( .A1(KEYINPUT63), .A2(G143), .ZN(n1345) );
XOR2_X1 U1073 ( .A(G122), .B(KEYINPUT0), .Z(n1319) );
XOR2_X1 U1074 ( .A(n1346), .B(n1347), .Z(n1342) );
XOR2_X1 U1075 ( .A(G134), .B(G116), .Z(n1347) );
XOR2_X1 U1076 ( .A(n1348), .B(G107), .Z(n1346) );
NAND2_X1 U1077 ( .A1(G217), .A2(n1270), .ZN(n1348) );
AND2_X1 U1078 ( .A1(G234), .A2(n1119), .ZN(n1270) );
INV_X1 U1079 ( .A(G953), .ZN(n1119) );
endmodule


