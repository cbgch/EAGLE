//Key = 0101010110011101000100110001000110000001101110100001101100110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375;

XNOR2_X1 U748 ( .A(n1048), .B(n1049), .ZN(G9) );
NOR4_X1 U749 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1049) );
INV_X1 U750 ( .A(n1054), .ZN(n1053) );
OR2_X1 U751 ( .A1(n1055), .A2(n1056), .ZN(n1051) );
XNOR2_X1 U752 ( .A(n1057), .B(KEYINPUT50), .ZN(n1050) );
NOR2_X1 U753 ( .A1(n1058), .A2(n1059), .ZN(G75) );
NOR3_X1 U754 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NOR2_X1 U755 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR3_X1 U756 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1063) );
NOR2_X1 U757 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
INV_X1 U758 ( .A(n1070), .ZN(n1069) );
NOR2_X1 U759 ( .A1(n1071), .A2(n1072), .ZN(n1068) );
NOR2_X1 U760 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR3_X1 U761 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1066) );
NOR3_X1 U762 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1076) );
NOR2_X1 U763 ( .A1(n1081), .A2(n1052), .ZN(n1080) );
NOR2_X1 U764 ( .A1(n1054), .A2(n1082), .ZN(n1081) );
NOR2_X1 U765 ( .A1(KEYINPUT17), .A2(n1083), .ZN(n1078) );
NOR2_X1 U766 ( .A1(n1084), .A2(n1085), .ZN(n1065) );
INV_X1 U767 ( .A(KEYINPUT17), .ZN(n1085) );
NOR3_X1 U768 ( .A1(n1083), .A2(n1077), .A3(n1075), .ZN(n1084) );
NAND3_X1 U769 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1060) );
NAND3_X1 U770 ( .A1(n1089), .A2(n1090), .A3(n1070), .ZN(n1088) );
NOR3_X1 U771 ( .A1(n1075), .A2(n1052), .A3(n1091), .ZN(n1070) );
INV_X1 U772 ( .A(n1092), .ZN(n1052) );
NAND2_X1 U773 ( .A1(n1093), .A2(n1094), .ZN(n1090) );
NAND2_X1 U774 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR3_X1 U775 ( .A1(n1097), .A2(G953), .A3(G952), .ZN(n1058) );
INV_X1 U776 ( .A(n1086), .ZN(n1097) );
NAND4_X1 U777 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1086) );
NOR4_X1 U778 ( .A1(n1102), .A2(n1103), .A3(n1077), .A4(n1104), .ZN(n1101) );
XNOR2_X1 U779 ( .A(n1105), .B(KEYINPUT19), .ZN(n1102) );
NOR2_X1 U780 ( .A1(n1095), .A2(n1106), .ZN(n1100) );
XNOR2_X1 U781 ( .A(n1107), .B(n1108), .ZN(n1099) );
NAND2_X1 U782 ( .A1(KEYINPUT62), .A2(n1109), .ZN(n1108) );
XOR2_X1 U783 ( .A(G475), .B(n1110), .Z(n1098) );
NOR2_X1 U784 ( .A1(n1111), .A2(KEYINPUT61), .ZN(n1110) );
XOR2_X1 U785 ( .A(n1112), .B(n1113), .Z(G72) );
NOR2_X1 U786 ( .A1(n1114), .A2(n1087), .ZN(n1113) );
NOR2_X1 U787 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U788 ( .A1(n1117), .A2(n1118), .ZN(n1112) );
NAND2_X1 U789 ( .A1(n1119), .A2(n1087), .ZN(n1118) );
XNOR2_X1 U790 ( .A(n1120), .B(n1121), .ZN(n1119) );
NAND3_X1 U791 ( .A1(G900), .A2(n1121), .A3(G953), .ZN(n1117) );
XOR2_X1 U792 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U793 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U794 ( .A1(KEYINPUT34), .A2(n1126), .ZN(n1124) );
XOR2_X1 U795 ( .A(n1127), .B(n1128), .Z(n1122) );
NOR2_X1 U796 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XOR2_X1 U797 ( .A(KEYINPUT30), .B(n1131), .Z(n1130) );
NOR2_X1 U798 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NOR2_X1 U799 ( .A1(G125), .A2(n1134), .ZN(n1129) );
XNOR2_X1 U800 ( .A(KEYINPUT2), .B(n1132), .ZN(n1134) );
NAND2_X1 U801 ( .A1(KEYINPUT32), .A2(n1135), .ZN(n1127) );
XNOR2_X1 U802 ( .A(KEYINPUT11), .B(n1136), .ZN(n1135) );
NAND3_X1 U803 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(G69) );
XOR2_X1 U804 ( .A(KEYINPUT7), .B(n1140), .Z(n1139) );
NOR3_X1 U805 ( .A1(n1087), .A2(n1141), .A3(n1142), .ZN(n1140) );
NOR2_X1 U806 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U807 ( .A1(n1145), .A2(n1087), .ZN(n1138) );
XOR2_X1 U808 ( .A(n1146), .B(n1141), .Z(n1145) );
NAND2_X1 U809 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND3_X1 U810 ( .A1(n1141), .A2(G224), .A3(G953), .ZN(n1137) );
AND2_X1 U811 ( .A1(n1149), .A2(n1150), .ZN(n1141) );
NAND2_X1 U812 ( .A1(G953), .A2(n1144), .ZN(n1150) );
XOR2_X1 U813 ( .A(n1151), .B(n1152), .Z(n1149) );
NAND2_X1 U814 ( .A1(KEYINPUT31), .A2(n1153), .ZN(n1151) );
NOR2_X1 U815 ( .A1(n1154), .A2(n1155), .ZN(G66) );
XOR2_X1 U816 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U817 ( .A1(n1158), .A2(n1159), .ZN(n1156) );
NOR2_X1 U818 ( .A1(n1154), .A2(n1160), .ZN(G63) );
XOR2_X1 U819 ( .A(n1161), .B(n1162), .Z(n1160) );
NAND2_X1 U820 ( .A1(n1158), .A2(G478), .ZN(n1161) );
NOR2_X1 U821 ( .A1(n1154), .A2(n1163), .ZN(G60) );
NOR3_X1 U822 ( .A1(n1111), .A2(n1164), .A3(n1165), .ZN(n1163) );
AND3_X1 U823 ( .A1(n1166), .A2(G475), .A3(n1158), .ZN(n1165) );
NOR2_X1 U824 ( .A1(n1167), .A2(n1166), .ZN(n1164) );
AND2_X1 U825 ( .A1(n1062), .A2(G475), .ZN(n1167) );
XOR2_X1 U826 ( .A(G104), .B(n1168), .Z(G6) );
NOR2_X1 U827 ( .A1(n1154), .A2(n1169), .ZN(G57) );
XOR2_X1 U828 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U829 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U830 ( .A1(KEYINPUT14), .A2(n1174), .ZN(n1173) );
XOR2_X1 U831 ( .A(n1175), .B(KEYINPUT9), .Z(n1174) );
NAND2_X1 U832 ( .A1(n1176), .A2(n1177), .ZN(n1172) );
NAND2_X1 U833 ( .A1(n1158), .A2(G472), .ZN(n1170) );
NOR2_X1 U834 ( .A1(n1154), .A2(n1178), .ZN(G54) );
XOR2_X1 U835 ( .A(n1179), .B(n1180), .Z(n1178) );
XNOR2_X1 U836 ( .A(n1181), .B(n1182), .ZN(n1180) );
XNOR2_X1 U837 ( .A(n1183), .B(n1184), .ZN(n1181) );
XOR2_X1 U838 ( .A(n1185), .B(n1186), .Z(n1179) );
XNOR2_X1 U839 ( .A(n1187), .B(n1132), .ZN(n1186) );
XOR2_X1 U840 ( .A(n1188), .B(KEYINPUT58), .Z(n1185) );
NAND2_X1 U841 ( .A1(n1158), .A2(G469), .ZN(n1188) );
NOR2_X1 U842 ( .A1(n1154), .A2(n1189), .ZN(G51) );
XOR2_X1 U843 ( .A(n1190), .B(n1191), .Z(n1189) );
XNOR2_X1 U844 ( .A(n1192), .B(n1193), .ZN(n1191) );
NAND2_X1 U845 ( .A1(n1158), .A2(n1107), .ZN(n1192) );
INV_X1 U846 ( .A(n1194), .ZN(n1107) );
AND2_X1 U847 ( .A1(G902), .A2(n1062), .ZN(n1158) );
NAND3_X1 U848 ( .A1(n1120), .A2(n1147), .A3(n1195), .ZN(n1062) );
XOR2_X1 U849 ( .A(n1148), .B(KEYINPUT29), .Z(n1195) );
AND4_X1 U850 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1147) );
NOR4_X1 U851 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1168), .ZN(n1199) );
AND3_X1 U852 ( .A1(n1082), .A2(n1092), .A3(n1203), .ZN(n1168) );
NOR3_X1 U853 ( .A1(n1083), .A2(n1204), .A3(n1205), .ZN(n1202) );
NOR2_X1 U854 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NOR2_X1 U855 ( .A1(n1057), .A2(n1056), .ZN(n1206) );
NOR2_X1 U856 ( .A1(n1203), .A2(n1208), .ZN(n1204) );
NOR2_X1 U857 ( .A1(n1055), .A2(n1207), .ZN(n1208) );
INV_X1 U858 ( .A(KEYINPUT48), .ZN(n1207) );
INV_X1 U859 ( .A(n1209), .ZN(n1201) );
NAND2_X1 U860 ( .A1(n1203), .A2(n1210), .ZN(n1198) );
NAND2_X1 U861 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
OR2_X1 U862 ( .A1(n1213), .A2(KEYINPUT37), .ZN(n1212) );
NAND2_X1 U863 ( .A1(n1054), .A2(n1092), .ZN(n1211) );
INV_X1 U864 ( .A(n1214), .ZN(n1203) );
NAND3_X1 U865 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1197) );
XNOR2_X1 U866 ( .A(KEYINPUT4), .B(n1091), .ZN(n1216) );
NAND4_X1 U867 ( .A1(KEYINPUT37), .A2(n1056), .A3(n1079), .A4(n1218), .ZN(n1196) );
INV_X1 U868 ( .A(n1213), .ZN(n1079) );
AND4_X1 U869 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1120) );
NOR4_X1 U870 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1222) );
INV_X1 U871 ( .A(n1227), .ZN(n1223) );
OR2_X1 U872 ( .A1(n1228), .A2(n1064), .ZN(n1221) );
NAND2_X1 U873 ( .A1(n1229), .A2(n1230), .ZN(n1219) );
NAND2_X1 U874 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND2_X1 U875 ( .A1(n1233), .A2(n1089), .ZN(n1232) );
XNOR2_X1 U876 ( .A(n1057), .B(KEYINPUT44), .ZN(n1233) );
NAND2_X1 U877 ( .A1(n1234), .A2(n1072), .ZN(n1231) );
INV_X1 U878 ( .A(n1235), .ZN(n1229) );
NAND2_X1 U879 ( .A1(n1236), .A2(n1237), .ZN(n1190) );
OR2_X1 U880 ( .A1(KEYINPUT28), .A2(n1238), .ZN(n1237) );
NAND2_X1 U881 ( .A1(KEYINPUT20), .A2(n1238), .ZN(n1236) );
XOR2_X1 U882 ( .A(n1239), .B(n1240), .Z(n1238) );
NAND2_X1 U883 ( .A1(KEYINPUT22), .A2(n1241), .ZN(n1239) );
AND2_X1 U884 ( .A1(n1242), .A2(G953), .ZN(n1154) );
XNOR2_X1 U885 ( .A(G952), .B(KEYINPUT47), .ZN(n1242) );
NAND2_X1 U886 ( .A1(n1243), .A2(n1244), .ZN(G48) );
NAND2_X1 U887 ( .A1(G146), .A2(n1220), .ZN(n1244) );
XOR2_X1 U888 ( .A(KEYINPUT12), .B(n1245), .Z(n1243) );
NOR2_X1 U889 ( .A1(G146), .A2(n1220), .ZN(n1245) );
NAND3_X1 U890 ( .A1(n1082), .A2(n1215), .A3(n1246), .ZN(n1220) );
AND3_X1 U891 ( .A1(n1057), .A2(n1247), .A3(n1072), .ZN(n1246) );
XOR2_X1 U892 ( .A(G143), .B(n1226), .Z(G45) );
AND4_X1 U893 ( .A1(n1248), .A2(n1057), .A3(n1104), .A4(n1249), .ZN(n1226) );
XOR2_X1 U894 ( .A(G140), .B(n1250), .Z(G42) );
NOR3_X1 U895 ( .A1(n1235), .A2(n1251), .A3(n1064), .ZN(n1250) );
XNOR2_X1 U896 ( .A(n1072), .B(KEYINPUT10), .ZN(n1251) );
XOR2_X1 U897 ( .A(G137), .B(n1225), .Z(G39) );
AND4_X1 U898 ( .A1(n1072), .A2(n1247), .A3(n1215), .A4(n1252), .ZN(n1225) );
NOR2_X1 U899 ( .A1(n1064), .A2(n1091), .ZN(n1252) );
INV_X1 U900 ( .A(n1253), .ZN(n1091) );
XOR2_X1 U901 ( .A(G134), .B(n1224), .Z(G36) );
AND3_X1 U902 ( .A1(n1234), .A2(n1054), .A3(n1248), .ZN(n1224) );
XNOR2_X1 U903 ( .A(G131), .B(n1254), .ZN(G33) );
NAND3_X1 U904 ( .A1(KEYINPUT3), .A2(n1234), .A3(n1255), .ZN(n1254) );
XOR2_X1 U905 ( .A(n1228), .B(KEYINPUT15), .Z(n1255) );
NAND2_X1 U906 ( .A1(n1082), .A2(n1248), .ZN(n1228) );
AND3_X1 U907 ( .A1(n1072), .A2(n1247), .A3(n1256), .ZN(n1248) );
INV_X1 U908 ( .A(n1064), .ZN(n1234) );
NAND2_X1 U909 ( .A1(n1096), .A2(n1257), .ZN(n1064) );
XNOR2_X1 U910 ( .A(G128), .B(n1227), .ZN(G30) );
NAND4_X1 U911 ( .A1(n1218), .A2(n1215), .A3(n1054), .A4(n1247), .ZN(n1227) );
XNOR2_X1 U912 ( .A(n1258), .B(n1259), .ZN(G3) );
NOR3_X1 U913 ( .A1(n1214), .A2(KEYINPUT33), .A3(n1083), .ZN(n1259) );
NAND2_X1 U914 ( .A1(n1253), .A2(n1256), .ZN(n1083) );
XNOR2_X1 U915 ( .A(n1133), .B(n1260), .ZN(G27) );
NOR3_X1 U916 ( .A1(n1235), .A2(n1093), .A3(n1077), .ZN(n1260) );
NAND4_X1 U917 ( .A1(n1082), .A2(n1261), .A3(n1262), .A4(n1247), .ZN(n1235) );
NAND2_X1 U918 ( .A1(n1263), .A2(n1264), .ZN(n1247) );
NAND4_X1 U919 ( .A1(G953), .A2(G902), .A3(n1265), .A4(n1116), .ZN(n1264) );
INV_X1 U920 ( .A(G900), .ZN(n1116) );
XOR2_X1 U921 ( .A(n1075), .B(KEYINPUT26), .Z(n1263) );
XOR2_X1 U922 ( .A(n1266), .B(n1267), .Z(G24) );
NOR2_X1 U923 ( .A1(KEYINPUT63), .A2(n1209), .ZN(n1267) );
NAND4_X1 U924 ( .A1(n1217), .A2(n1092), .A3(n1104), .A4(n1249), .ZN(n1209) );
NOR2_X1 U925 ( .A1(n1268), .A2(n1262), .ZN(n1092) );
XNOR2_X1 U926 ( .A(G122), .B(KEYINPUT27), .ZN(n1266) );
XOR2_X1 U927 ( .A(n1269), .B(n1270), .Z(G21) );
NOR2_X1 U928 ( .A1(n1271), .A2(n1093), .ZN(n1270) );
XOR2_X1 U929 ( .A(n1272), .B(KEYINPUT56), .Z(n1271) );
NAND4_X1 U930 ( .A1(n1253), .A2(n1215), .A3(n1089), .A4(n1273), .ZN(n1272) );
INV_X1 U931 ( .A(n1077), .ZN(n1089) );
AND2_X1 U932 ( .A1(n1262), .A2(n1268), .ZN(n1215) );
XNOR2_X1 U933 ( .A(G119), .B(KEYINPUT52), .ZN(n1269) );
XOR2_X1 U934 ( .A(G116), .B(n1200), .Z(G18) );
AND3_X1 U935 ( .A1(n1256), .A2(n1054), .A3(n1217), .ZN(n1200) );
NOR2_X1 U936 ( .A1(n1249), .A2(n1274), .ZN(n1054) );
XOR2_X1 U937 ( .A(n1148), .B(n1275), .Z(G15) );
XNOR2_X1 U938 ( .A(KEYINPUT55), .B(n1276), .ZN(n1275) );
NAND3_X1 U939 ( .A1(n1082), .A2(n1256), .A3(n1217), .ZN(n1148) );
NOR3_X1 U940 ( .A1(n1093), .A2(n1056), .A3(n1077), .ZN(n1217) );
NAND2_X1 U941 ( .A1(n1277), .A2(n1074), .ZN(n1077) );
INV_X1 U942 ( .A(n1073), .ZN(n1277) );
INV_X1 U943 ( .A(n1273), .ZN(n1056) );
NOR2_X1 U944 ( .A1(n1262), .A2(n1278), .ZN(n1256) );
AND2_X1 U945 ( .A1(n1274), .A2(n1249), .ZN(n1082) );
INV_X1 U946 ( .A(n1104), .ZN(n1274) );
XOR2_X1 U947 ( .A(G110), .B(n1279), .Z(G12) );
NOR2_X1 U948 ( .A1(n1214), .A2(n1213), .ZN(n1279) );
NAND3_X1 U949 ( .A1(n1261), .A2(n1262), .A3(n1253), .ZN(n1213) );
NOR2_X1 U950 ( .A1(n1104), .A2(n1249), .ZN(n1253) );
XOR2_X1 U951 ( .A(n1111), .B(n1280), .Z(n1249) );
XOR2_X1 U952 ( .A(KEYINPUT18), .B(G475), .Z(n1280) );
NOR2_X1 U953 ( .A1(n1166), .A2(G902), .ZN(n1111) );
XOR2_X1 U954 ( .A(n1281), .B(n1282), .Z(n1166) );
XOR2_X1 U955 ( .A(n1283), .B(n1284), .Z(n1282) );
XNOR2_X1 U956 ( .A(n1276), .B(G104), .ZN(n1284) );
XOR2_X1 U957 ( .A(G131), .B(G122), .Z(n1283) );
XOR2_X1 U958 ( .A(n1285), .B(n1286), .Z(n1281) );
XNOR2_X1 U959 ( .A(n1287), .B(n1288), .ZN(n1285) );
AND3_X1 U960 ( .A1(G214), .A2(n1087), .A3(n1289), .ZN(n1288) );
XNOR2_X1 U961 ( .A(n1290), .B(G478), .ZN(n1104) );
NAND2_X1 U962 ( .A1(n1162), .A2(n1291), .ZN(n1290) );
XOR2_X1 U963 ( .A(n1292), .B(n1293), .Z(n1162) );
XOR2_X1 U964 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U965 ( .A(G122), .B(G116), .Z(n1295) );
XNOR2_X1 U966 ( .A(G134), .B(n1296), .ZN(n1294) );
XOR2_X1 U967 ( .A(n1297), .B(n1298), .Z(n1292) );
XNOR2_X1 U968 ( .A(n1299), .B(n1048), .ZN(n1297) );
NAND2_X1 U969 ( .A1(G217), .A2(n1300), .ZN(n1299) );
XOR2_X1 U970 ( .A(n1103), .B(KEYINPUT41), .Z(n1262) );
XNOR2_X1 U971 ( .A(n1301), .B(n1159), .ZN(n1103) );
AND2_X1 U972 ( .A1(G217), .A2(n1302), .ZN(n1159) );
NAND2_X1 U973 ( .A1(n1157), .A2(n1291), .ZN(n1301) );
XNOR2_X1 U974 ( .A(n1303), .B(n1304), .ZN(n1157) );
XOR2_X1 U975 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U976 ( .A(G146), .B(G110), .Z(n1306) );
XOR2_X1 U977 ( .A(KEYINPUT5), .B(KEYINPUT38), .Z(n1305) );
XOR2_X1 U978 ( .A(n1307), .B(n1308), .Z(n1303) );
XOR2_X1 U979 ( .A(n1309), .B(n1286), .Z(n1308) );
XNOR2_X1 U980 ( .A(G125), .B(n1132), .ZN(n1286) );
AND2_X1 U981 ( .A1(n1300), .A2(G221), .ZN(n1309) );
AND2_X1 U982 ( .A1(G234), .A2(n1087), .ZN(n1300) );
XOR2_X1 U983 ( .A(n1310), .B(n1311), .Z(n1307) );
NOR2_X1 U984 ( .A1(KEYINPUT24), .A2(G137), .ZN(n1311) );
NAND2_X1 U985 ( .A1(n1312), .A2(n1313), .ZN(n1310) );
NAND2_X1 U986 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
XOR2_X1 U987 ( .A(KEYINPUT40), .B(n1316), .Z(n1312) );
NOR2_X1 U988 ( .A1(n1315), .A2(n1314), .ZN(n1316) );
XNOR2_X1 U989 ( .A(KEYINPUT35), .B(n1296), .ZN(n1314) );
INV_X1 U990 ( .A(G119), .ZN(n1315) );
XNOR2_X1 U991 ( .A(n1268), .B(KEYINPUT53), .ZN(n1261) );
INV_X1 U992 ( .A(n1278), .ZN(n1268) );
NOR2_X1 U993 ( .A1(n1105), .A2(n1106), .ZN(n1278) );
NOR3_X1 U994 ( .A1(G472), .A2(G902), .A3(n1317), .ZN(n1106) );
XNOR2_X1 U995 ( .A(n1175), .B(n1318), .ZN(n1317) );
AND2_X1 U996 ( .A1(G472), .A2(n1319), .ZN(n1105) );
NAND2_X1 U997 ( .A1(n1320), .A2(n1291), .ZN(n1319) );
XOR2_X1 U998 ( .A(n1175), .B(n1318), .Z(n1320) );
AND2_X1 U999 ( .A1(n1321), .A2(n1176), .ZN(n1318) );
NAND2_X1 U1000 ( .A1(n1258), .A2(n1322), .ZN(n1176) );
NAND3_X1 U1001 ( .A1(n1289), .A2(n1087), .A3(G210), .ZN(n1322) );
XNOR2_X1 U1002 ( .A(KEYINPUT23), .B(n1177), .ZN(n1321) );
NAND4_X1 U1003 ( .A1(G101), .A2(G210), .A3(n1289), .A4(n1087), .ZN(n1177) );
XOR2_X1 U1004 ( .A(n1323), .B(n1324), .Z(n1175) );
XOR2_X1 U1005 ( .A(n1241), .B(n1325), .Z(n1324) );
NAND2_X1 U1006 ( .A1(KEYINPUT1), .A2(n1276), .ZN(n1325) );
XNOR2_X1 U1007 ( .A(n1326), .B(n1327), .ZN(n1323) );
INV_X1 U1008 ( .A(n1183), .ZN(n1327) );
NAND2_X1 U1009 ( .A1(n1218), .A2(n1273), .ZN(n1214) );
NAND2_X1 U1010 ( .A1(n1075), .A2(n1328), .ZN(n1273) );
NAND4_X1 U1011 ( .A1(G953), .A2(G902), .A3(n1265), .A4(n1144), .ZN(n1328) );
INV_X1 U1012 ( .A(G898), .ZN(n1144) );
NAND3_X1 U1013 ( .A1(n1265), .A2(n1087), .A3(G952), .ZN(n1075) );
INV_X1 U1014 ( .A(G953), .ZN(n1087) );
NAND2_X1 U1015 ( .A1(n1329), .A2(G237), .ZN(n1265) );
XNOR2_X1 U1016 ( .A(G234), .B(KEYINPUT51), .ZN(n1329) );
NOR2_X1 U1017 ( .A1(n1093), .A2(n1055), .ZN(n1218) );
XNOR2_X1 U1018 ( .A(n1072), .B(KEYINPUT45), .ZN(n1055) );
AND2_X1 U1019 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U1020 ( .A1(G221), .A2(n1302), .ZN(n1074) );
NAND2_X1 U1021 ( .A1(G234), .A2(n1291), .ZN(n1302) );
XNOR2_X1 U1022 ( .A(n1330), .B(G469), .ZN(n1073) );
NAND2_X1 U1023 ( .A1(n1331), .A2(n1291), .ZN(n1330) );
XNOR2_X1 U1024 ( .A(n1332), .B(n1333), .ZN(n1331) );
INV_X1 U1025 ( .A(n1187), .ZN(n1333) );
XOR2_X1 U1026 ( .A(G110), .B(n1334), .Z(n1187) );
NOR2_X1 U1027 ( .A1(G953), .A2(n1115), .ZN(n1334) );
INV_X1 U1028 ( .A(G227), .ZN(n1115) );
XNOR2_X1 U1029 ( .A(n1335), .B(n1336), .ZN(n1332) );
NOR2_X1 U1030 ( .A1(KEYINPUT6), .A2(n1132), .ZN(n1336) );
XNOR2_X1 U1031 ( .A(G140), .B(KEYINPUT54), .ZN(n1132) );
NOR2_X1 U1032 ( .A1(KEYINPUT0), .A2(n1337), .ZN(n1335) );
XNOR2_X1 U1033 ( .A(n1338), .B(n1183), .ZN(n1337) );
XOR2_X1 U1034 ( .A(n1125), .B(n1126), .Z(n1183) );
XOR2_X1 U1035 ( .A(G131), .B(KEYINPUT25), .Z(n1126) );
XOR2_X1 U1036 ( .A(G134), .B(G137), .Z(n1125) );
NAND2_X1 U1037 ( .A1(KEYINPUT59), .A2(n1339), .ZN(n1338) );
NAND3_X1 U1038 ( .A1(n1340), .A2(n1341), .A3(n1342), .ZN(n1339) );
NAND2_X1 U1039 ( .A1(n1182), .A2(n1343), .ZN(n1342) );
NAND2_X1 U1040 ( .A1(n1344), .A2(KEYINPUT13), .ZN(n1343) );
XNOR2_X1 U1041 ( .A(n1184), .B(KEYINPUT49), .ZN(n1344) );
INV_X1 U1042 ( .A(n1345), .ZN(n1182) );
NAND3_X1 U1043 ( .A1(KEYINPUT13), .A2(n1345), .A3(n1136), .ZN(n1341) );
XNOR2_X1 U1044 ( .A(n1346), .B(n1347), .ZN(n1345) );
XNOR2_X1 U1045 ( .A(G101), .B(G107), .ZN(n1346) );
OR2_X1 U1046 ( .A1(n1136), .A2(KEYINPUT13), .ZN(n1340) );
INV_X1 U1047 ( .A(n1184), .ZN(n1136) );
XOR2_X1 U1048 ( .A(n1348), .B(n1349), .Z(n1184) );
XNOR2_X1 U1049 ( .A(G128), .B(KEYINPUT57), .ZN(n1348) );
INV_X1 U1050 ( .A(n1057), .ZN(n1093) );
NOR2_X1 U1051 ( .A1(n1096), .A2(n1095), .ZN(n1057) );
INV_X1 U1052 ( .A(n1257), .ZN(n1095) );
NAND2_X1 U1053 ( .A1(G214), .A2(n1350), .ZN(n1257) );
XNOR2_X1 U1054 ( .A(n1351), .B(n1194), .ZN(n1096) );
NAND2_X1 U1055 ( .A1(G210), .A2(n1350), .ZN(n1194) );
NAND2_X1 U1056 ( .A1(n1289), .A2(n1291), .ZN(n1350) );
INV_X1 U1057 ( .A(G237), .ZN(n1289) );
XOR2_X1 U1058 ( .A(n1109), .B(KEYINPUT16), .Z(n1351) );
NAND2_X1 U1059 ( .A1(n1352), .A2(n1291), .ZN(n1109) );
INV_X1 U1060 ( .A(G902), .ZN(n1291) );
XOR2_X1 U1061 ( .A(n1240), .B(n1353), .Z(n1352) );
XNOR2_X1 U1062 ( .A(n1241), .B(n1193), .ZN(n1353) );
XOR2_X1 U1063 ( .A(n1153), .B(n1152), .Z(n1193) );
XNOR2_X1 U1064 ( .A(n1326), .B(n1354), .ZN(n1152) );
XOR2_X1 U1065 ( .A(n1355), .B(n1356), .Z(n1354) );
NAND2_X1 U1066 ( .A1(KEYINPUT39), .A2(n1276), .ZN(n1356) );
INV_X1 U1067 ( .A(G113), .ZN(n1276) );
NAND3_X1 U1068 ( .A1(n1357), .A2(n1358), .A3(n1359), .ZN(n1355) );
OR2_X1 U1069 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NAND4_X1 U1070 ( .A1(n1361), .A2(n1360), .A3(KEYINPUT46), .A4(n1258), .ZN(n1358) );
INV_X1 U1071 ( .A(G101), .ZN(n1258) );
INV_X1 U1072 ( .A(KEYINPUT60), .ZN(n1360) );
NAND2_X1 U1073 ( .A1(G101), .A2(n1362), .ZN(n1357) );
NAND2_X1 U1074 ( .A1(KEYINPUT46), .A2(n1361), .ZN(n1362) );
NAND3_X1 U1075 ( .A1(n1363), .A2(n1364), .A3(n1365), .ZN(n1361) );
OR2_X1 U1076 ( .A1(n1347), .A2(n1048), .ZN(n1365) );
NAND2_X1 U1077 ( .A1(n1366), .A2(n1367), .ZN(n1364) );
INV_X1 U1078 ( .A(KEYINPUT8), .ZN(n1367) );
NAND2_X1 U1079 ( .A1(n1368), .A2(n1048), .ZN(n1366) );
XNOR2_X1 U1080 ( .A(KEYINPUT43), .B(n1347), .ZN(n1368) );
NAND2_X1 U1081 ( .A1(KEYINPUT8), .A2(n1369), .ZN(n1363) );
NAND2_X1 U1082 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
OR2_X1 U1083 ( .A1(n1347), .A2(KEYINPUT43), .ZN(n1371) );
NAND3_X1 U1084 ( .A1(n1347), .A2(n1048), .A3(KEYINPUT43), .ZN(n1370) );
INV_X1 U1085 ( .A(G107), .ZN(n1048) );
XOR2_X1 U1086 ( .A(G104), .B(KEYINPUT36), .Z(n1347) );
XNOR2_X1 U1087 ( .A(G116), .B(G119), .ZN(n1326) );
XOR2_X1 U1088 ( .A(G110), .B(G122), .Z(n1153) );
NAND2_X1 U1089 ( .A1(n1372), .A2(n1373), .ZN(n1241) );
NAND2_X1 U1090 ( .A1(G128), .A2(n1349), .ZN(n1373) );
INV_X1 U1091 ( .A(n1287), .ZN(n1349) );
XOR2_X1 U1092 ( .A(n1374), .B(KEYINPUT21), .Z(n1372) );
NAND2_X1 U1093 ( .A1(n1287), .A2(n1296), .ZN(n1374) );
INV_X1 U1094 ( .A(G128), .ZN(n1296) );
XOR2_X1 U1095 ( .A(G146), .B(n1298), .Z(n1287) );
XOR2_X1 U1096 ( .A(G143), .B(KEYINPUT42), .Z(n1298) );
XNOR2_X1 U1097 ( .A(n1133), .B(n1375), .ZN(n1240) );
NOR2_X1 U1098 ( .A1(G953), .A2(n1143), .ZN(n1375) );
INV_X1 U1099 ( .A(G224), .ZN(n1143) );
INV_X1 U1100 ( .A(G125), .ZN(n1133) );
endmodule


