//Key = 0100010000011011000011101111011101010110101011010001111110110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366;

XNOR2_X1 U765 ( .A(G107), .B(n1042), .ZN(G9) );
NOR2_X1 U766 ( .A1(n1043), .A2(n1044), .ZN(G75) );
NOR4_X1 U767 ( .A1(G953), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1044) );
INV_X1 U768 ( .A(n1048), .ZN(n1047) );
NOR2_X1 U769 ( .A1(n1049), .A2(n1050), .ZN(n1046) );
NOR2_X1 U770 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR4_X1 U771 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
AND2_X1 U772 ( .A1(n1057), .A2(n1058), .ZN(n1054) );
NOR2_X1 U773 ( .A1(n1057), .A2(n1059), .ZN(n1053) );
NOR4_X1 U774 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1051) );
NOR2_X1 U775 ( .A1(n1055), .A2(n1064), .ZN(n1061) );
NOR2_X1 U776 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR3_X1 U777 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
NOR2_X1 U778 ( .A1(n1058), .A2(n1070), .ZN(n1069) );
NOR3_X1 U779 ( .A1(n1062), .A2(n1071), .A3(n1072), .ZN(n1058) );
NOR2_X1 U780 ( .A1(n1073), .A2(n1074), .ZN(n1068) );
NOR2_X1 U781 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NOR2_X1 U782 ( .A1(n1077), .A2(n1078), .ZN(n1065) );
NOR2_X1 U783 ( .A1(n1074), .A2(n1070), .ZN(n1077) );
INV_X1 U784 ( .A(n1079), .ZN(n1074) );
AND2_X1 U785 ( .A1(n1056), .A2(n1055), .ZN(n1060) );
NAND3_X1 U786 ( .A1(n1079), .A2(n1078), .A3(n1080), .ZN(n1056) );
NOR3_X1 U787 ( .A1(n1045), .A2(G953), .A3(G952), .ZN(n1043) );
AND4_X1 U788 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1045) );
NOR4_X1 U789 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1084) );
XOR2_X1 U790 ( .A(n1089), .B(n1090), .Z(n1088) );
XNOR2_X1 U791 ( .A(n1091), .B(G475), .ZN(n1090) );
XNOR2_X1 U792 ( .A(KEYINPUT57), .B(KEYINPUT50), .ZN(n1089) );
XOR2_X1 U793 ( .A(n1092), .B(n1093), .Z(n1086) );
XNOR2_X1 U794 ( .A(G469), .B(KEYINPUT32), .ZN(n1093) );
NAND4_X1 U795 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1085) );
NAND3_X1 U796 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1097) );
NAND2_X1 U797 ( .A1(n1101), .A2(n1102), .ZN(n1096) );
INV_X1 U798 ( .A(n1100), .ZN(n1102) );
NAND2_X1 U799 ( .A1(n1103), .A2(n1099), .ZN(n1101) );
XNOR2_X1 U800 ( .A(KEYINPUT52), .B(n1098), .ZN(n1103) );
NAND2_X1 U801 ( .A1(KEYINPUT8), .A2(n1104), .ZN(n1095) );
NAND2_X1 U802 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XNOR2_X1 U803 ( .A(n1107), .B(KEYINPUT15), .ZN(n1105) );
NAND2_X1 U804 ( .A1(n1108), .A2(n1109), .ZN(n1094) );
INV_X1 U805 ( .A(KEYINPUT8), .ZN(n1109) );
NAND2_X1 U806 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
OR2_X1 U807 ( .A1(n1107), .A2(KEYINPUT15), .ZN(n1111) );
NAND3_X1 U808 ( .A1(n1107), .A2(n1106), .A3(KEYINPUT15), .ZN(n1110) );
NOR3_X1 U809 ( .A1(n1112), .A2(n1067), .A3(n1113), .ZN(n1083) );
NOR2_X1 U810 ( .A1(n1107), .A2(n1106), .ZN(n1113) );
INV_X1 U811 ( .A(n1078), .ZN(n1067) );
XNOR2_X1 U812 ( .A(n1062), .B(KEYINPUT24), .ZN(n1112) );
INV_X1 U813 ( .A(n1059), .ZN(n1062) );
OR2_X1 U814 ( .A1(n1099), .A2(n1098), .ZN(n1082) );
XOR2_X1 U815 ( .A(n1114), .B(KEYINPUT48), .Z(n1098) );
INV_X1 U816 ( .A(KEYINPUT46), .ZN(n1099) );
XOR2_X1 U817 ( .A(n1115), .B(n1116), .Z(G72) );
NAND2_X1 U818 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U819 ( .A1(G900), .A2(G227), .ZN(n1118) );
NAND3_X1 U820 ( .A1(KEYINPUT40), .A2(n1119), .A3(n1120), .ZN(n1115) );
XOR2_X1 U821 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U822 ( .A1(KEYINPUT28), .A2(n1123), .ZN(n1122) );
XOR2_X1 U823 ( .A(n1124), .B(n1125), .Z(n1123) );
XNOR2_X1 U824 ( .A(n1126), .B(n1127), .ZN(n1125) );
NOR2_X1 U825 ( .A1(G131), .A2(KEYINPUT49), .ZN(n1127) );
NAND2_X1 U826 ( .A1(KEYINPUT21), .A2(n1128), .ZN(n1126) );
XOR2_X1 U827 ( .A(KEYINPUT6), .B(n1129), .Z(n1128) );
XOR2_X1 U828 ( .A(n1130), .B(n1131), .Z(n1124) );
XOR2_X1 U829 ( .A(G137), .B(n1132), .Z(n1131) );
NOR2_X1 U830 ( .A1(KEYINPUT2), .A2(n1133), .ZN(n1132) );
XNOR2_X1 U831 ( .A(n1134), .B(n1135), .ZN(n1133) );
XNOR2_X1 U832 ( .A(KEYINPUT61), .B(n1136), .ZN(n1135) );
NAND2_X1 U833 ( .A1(KEYINPUT35), .A2(n1137), .ZN(n1130) );
INV_X1 U834 ( .A(G134), .ZN(n1137) );
OR2_X1 U835 ( .A1(n1138), .A2(G900), .ZN(n1119) );
XOR2_X1 U836 ( .A(n1139), .B(n1140), .Z(G69) );
XOR2_X1 U837 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U838 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
OR2_X1 U839 ( .A1(n1138), .A2(G898), .ZN(n1144) );
XOR2_X1 U840 ( .A(n1145), .B(n1146), .Z(n1143) );
NAND2_X1 U841 ( .A1(KEYINPUT31), .A2(n1147), .ZN(n1145) );
NAND2_X1 U842 ( .A1(n1148), .A2(n1117), .ZN(n1141) );
XNOR2_X1 U843 ( .A(KEYINPUT19), .B(n1138), .ZN(n1117) );
XOR2_X1 U844 ( .A(KEYINPUT53), .B(n1149), .Z(n1148) );
AND2_X1 U845 ( .A1(G898), .A2(G224), .ZN(n1149) );
NOR2_X1 U846 ( .A1(n1150), .A2(G953), .ZN(n1139) );
NOR2_X1 U847 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U848 ( .A1(n1153), .A2(n1154), .ZN(G66) );
NOR3_X1 U849 ( .A1(n1100), .A2(n1155), .A3(n1156), .ZN(n1154) );
NOR2_X1 U850 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NOR2_X1 U851 ( .A1(n1048), .A2(n1114), .ZN(n1157) );
NOR3_X1 U852 ( .A1(n1159), .A2(n1114), .A3(n1160), .ZN(n1155) );
INV_X1 U853 ( .A(n1158), .ZN(n1159) );
NOR2_X1 U854 ( .A1(n1153), .A2(n1161), .ZN(G63) );
XOR2_X1 U855 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U856 ( .A1(n1164), .A2(G478), .ZN(n1162) );
NOR2_X1 U857 ( .A1(n1153), .A2(n1165), .ZN(G60) );
NOR3_X1 U858 ( .A1(n1091), .A2(n1166), .A3(n1167), .ZN(n1165) );
NOR3_X1 U859 ( .A1(n1168), .A2(n1169), .A3(n1160), .ZN(n1167) );
INV_X1 U860 ( .A(n1164), .ZN(n1160) );
NOR2_X1 U861 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
NOR2_X1 U862 ( .A1(n1048), .A2(n1169), .ZN(n1170) );
XNOR2_X1 U863 ( .A(G104), .B(n1172), .ZN(G6) );
NOR2_X1 U864 ( .A1(n1153), .A2(n1173), .ZN(G57) );
NOR3_X1 U865 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1173) );
NOR2_X1 U866 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR2_X1 U867 ( .A1(n1179), .A2(n1180), .ZN(n1177) );
XNOR2_X1 U868 ( .A(n1181), .B(KEYINPUT12), .ZN(n1179) );
NOR3_X1 U869 ( .A1(n1182), .A2(n1181), .A3(n1180), .ZN(n1175) );
INV_X1 U870 ( .A(KEYINPUT51), .ZN(n1180) );
NOR2_X1 U871 ( .A1(KEYINPUT51), .A2(n1183), .ZN(n1174) );
INV_X1 U872 ( .A(n1181), .ZN(n1183) );
XNOR2_X1 U873 ( .A(n1184), .B(n1185), .ZN(n1181) );
XOR2_X1 U874 ( .A(n1186), .B(n1187), .Z(n1184) );
NAND2_X1 U875 ( .A1(n1164), .A2(G472), .ZN(n1186) );
NOR2_X1 U876 ( .A1(n1153), .A2(n1188), .ZN(G54) );
XOR2_X1 U877 ( .A(n1189), .B(n1190), .Z(n1188) );
XNOR2_X1 U878 ( .A(n1191), .B(n1192), .ZN(n1190) );
XOR2_X1 U879 ( .A(n1193), .B(KEYINPUT44), .Z(n1189) );
NAND2_X1 U880 ( .A1(n1164), .A2(G469), .ZN(n1193) );
NOR2_X1 U881 ( .A1(n1153), .A2(n1194), .ZN(G51) );
XOR2_X1 U882 ( .A(n1195), .B(n1196), .Z(n1194) );
XNOR2_X1 U883 ( .A(n1197), .B(n1198), .ZN(n1196) );
NAND2_X1 U884 ( .A1(n1164), .A2(n1199), .ZN(n1197) );
NOR2_X1 U885 ( .A1(n1200), .A2(n1048), .ZN(n1164) );
NOR3_X1 U886 ( .A1(n1152), .A2(n1201), .A3(n1121), .ZN(n1048) );
NAND4_X1 U887 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1121) );
NOR4_X1 U888 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1205) );
INV_X1 U889 ( .A(n1210), .ZN(n1208) );
NOR3_X1 U890 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1207) );
XNOR2_X1 U891 ( .A(n1071), .B(KEYINPUT43), .ZN(n1212) );
AND2_X1 U892 ( .A1(n1214), .A2(n1215), .ZN(n1204) );
XOR2_X1 U893 ( .A(KEYINPUT9), .B(n1151), .Z(n1201) );
NAND4_X1 U894 ( .A1(n1172), .A2(n1216), .A3(n1217), .A4(n1042), .ZN(n1151) );
NAND3_X1 U895 ( .A1(n1079), .A2(n1075), .A3(n1218), .ZN(n1042) );
NAND3_X1 U896 ( .A1(n1218), .A2(n1079), .A3(n1076), .ZN(n1172) );
NAND4_X1 U897 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1152) );
NOR2_X1 U898 ( .A1(n1223), .A2(n1224), .ZN(n1195) );
NOR3_X1 U899 ( .A1(n1225), .A2(KEYINPUT36), .A3(n1226), .ZN(n1224) );
INV_X1 U900 ( .A(n1227), .ZN(n1225) );
NOR2_X1 U901 ( .A1(n1228), .A2(n1227), .ZN(n1223) );
NOR2_X1 U902 ( .A1(KEYINPUT36), .A2(n1226), .ZN(n1228) );
NOR2_X1 U903 ( .A1(n1138), .A2(G952), .ZN(n1153) );
XNOR2_X1 U904 ( .A(n1229), .B(n1230), .ZN(G48) );
NOR2_X1 U905 ( .A1(KEYINPUT60), .A2(n1215), .ZN(n1230) );
NAND2_X1 U906 ( .A1(n1076), .A2(n1231), .ZN(n1215) );
XOR2_X1 U907 ( .A(G143), .B(n1232), .Z(G45) );
NOR2_X1 U908 ( .A1(KEYINPUT39), .A2(n1214), .ZN(n1232) );
NAND4_X1 U909 ( .A1(n1055), .A2(n1087), .A3(n1233), .A4(n1234), .ZN(n1214) );
NOR2_X1 U910 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XNOR2_X1 U911 ( .A(G140), .B(n1202), .ZN(G42) );
NAND3_X1 U912 ( .A1(n1072), .A2(n1237), .A3(n1076), .ZN(n1202) );
XNOR2_X1 U913 ( .A(G137), .B(n1203), .ZN(G39) );
NAND2_X1 U914 ( .A1(n1238), .A2(n1237), .ZN(n1203) );
XNOR2_X1 U915 ( .A(G134), .B(n1239), .ZN(G36) );
NAND2_X1 U916 ( .A1(n1240), .A2(n1237), .ZN(n1239) );
XOR2_X1 U917 ( .A(G131), .B(n1209), .Z(G33) );
AND3_X1 U918 ( .A1(n1237), .A2(n1071), .A3(n1076), .ZN(n1209) );
INV_X1 U919 ( .A(n1211), .ZN(n1237) );
NAND3_X1 U920 ( .A1(n1055), .A2(n1057), .A3(n1241), .ZN(n1211) );
XNOR2_X1 U921 ( .A(n1242), .B(n1206), .ZN(G30) );
AND2_X1 U922 ( .A1(n1231), .A2(n1075), .ZN(n1206) );
INV_X1 U923 ( .A(n1213), .ZN(n1075) );
AND4_X1 U924 ( .A1(n1233), .A2(n1055), .A3(n1243), .A4(n1244), .ZN(n1231) );
XNOR2_X1 U925 ( .A(G101), .B(n1245), .ZN(G3) );
NOR2_X1 U926 ( .A1(n1246), .A2(KEYINPUT17), .ZN(n1245) );
INV_X1 U927 ( .A(n1216), .ZN(n1246) );
NAND3_X1 U928 ( .A1(n1071), .A2(n1218), .A3(n1080), .ZN(n1216) );
XNOR2_X1 U929 ( .A(G125), .B(n1210), .ZN(G27) );
NAND4_X1 U930 ( .A1(n1076), .A2(n1072), .A3(n1233), .A4(n1247), .ZN(n1210) );
AND2_X1 U931 ( .A1(n1241), .A2(n1063), .ZN(n1233) );
AND3_X1 U932 ( .A1(n1248), .A2(n1078), .A3(n1249), .ZN(n1241) );
NAND2_X1 U933 ( .A1(G900), .A2(n1050), .ZN(n1248) );
XNOR2_X1 U934 ( .A(G122), .B(n1219), .ZN(G24) );
NAND4_X1 U935 ( .A1(n1250), .A2(n1251), .A3(n1079), .A4(n1087), .ZN(n1219) );
NOR2_X1 U936 ( .A1(n1244), .A2(n1243), .ZN(n1079) );
INV_X1 U937 ( .A(n1236), .ZN(n1250) );
XNOR2_X1 U938 ( .A(G119), .B(n1220), .ZN(G21) );
NAND2_X1 U939 ( .A1(n1251), .A2(n1238), .ZN(n1220) );
AND3_X1 U940 ( .A1(n1243), .A2(n1244), .A3(n1080), .ZN(n1238) );
XNOR2_X1 U941 ( .A(G116), .B(n1221), .ZN(G18) );
NAND2_X1 U942 ( .A1(n1240), .A2(n1251), .ZN(n1221) );
NOR2_X1 U943 ( .A1(n1235), .A2(n1213), .ZN(n1240) );
NAND2_X1 U944 ( .A1(n1252), .A2(n1236), .ZN(n1213) );
XNOR2_X1 U945 ( .A(n1087), .B(KEYINPUT1), .ZN(n1252) );
INV_X1 U946 ( .A(n1071), .ZN(n1235) );
XNOR2_X1 U947 ( .A(G113), .B(n1222), .ZN(G15) );
NAND3_X1 U948 ( .A1(n1076), .A2(n1071), .A3(n1251), .ZN(n1222) );
AND3_X1 U949 ( .A1(n1078), .A2(n1247), .A3(n1253), .ZN(n1251) );
NOR2_X1 U950 ( .A1(n1243), .A2(n1081), .ZN(n1071) );
NOR2_X1 U951 ( .A1(n1236), .A2(n1087), .ZN(n1076) );
NAND2_X1 U952 ( .A1(n1254), .A2(n1255), .ZN(G12) );
NAND2_X1 U953 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND2_X1 U954 ( .A1(G110), .A2(n1258), .ZN(n1254) );
NAND2_X1 U955 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
OR2_X1 U956 ( .A1(n1217), .A2(KEYINPUT14), .ZN(n1260) );
NAND2_X1 U957 ( .A1(KEYINPUT14), .A2(n1261), .ZN(n1259) );
INV_X1 U958 ( .A(n1256), .ZN(n1261) );
NOR2_X1 U959 ( .A1(KEYINPUT18), .A2(n1217), .ZN(n1256) );
NAND3_X1 U960 ( .A1(n1072), .A2(n1218), .A3(n1080), .ZN(n1217) );
INV_X1 U961 ( .A(n1070), .ZN(n1080) );
NAND2_X1 U962 ( .A1(n1262), .A2(n1236), .ZN(n1070) );
XOR2_X1 U963 ( .A(n1263), .B(n1169), .Z(n1236) );
INV_X1 U964 ( .A(G475), .ZN(n1169) );
NAND2_X1 U965 ( .A1(KEYINPUT45), .A2(n1264), .ZN(n1263) );
INV_X1 U966 ( .A(n1091), .ZN(n1264) );
NOR2_X1 U967 ( .A1(n1171), .A2(G902), .ZN(n1091) );
INV_X1 U968 ( .A(n1168), .ZN(n1171) );
XNOR2_X1 U969 ( .A(n1265), .B(n1266), .ZN(n1168) );
XOR2_X1 U970 ( .A(KEYINPUT47), .B(G143), .Z(n1266) );
XOR2_X1 U971 ( .A(n1267), .B(n1268), .Z(n1265) );
XOR2_X1 U972 ( .A(n1269), .B(n1270), .Z(n1268) );
XNOR2_X1 U973 ( .A(n1271), .B(n1272), .ZN(n1270) );
NAND2_X1 U974 ( .A1(n1273), .A2(G214), .ZN(n1271) );
XNOR2_X1 U975 ( .A(G125), .B(G131), .ZN(n1269) );
XOR2_X1 U976 ( .A(n1274), .B(n1275), .Z(n1267) );
XNOR2_X1 U977 ( .A(n1276), .B(n1277), .ZN(n1275) );
INV_X1 U978 ( .A(n1278), .ZN(n1276) );
XOR2_X1 U979 ( .A(n1279), .B(n1280), .Z(n1274) );
NAND2_X1 U980 ( .A1(KEYINPUT30), .A2(n1136), .ZN(n1279) );
XOR2_X1 U981 ( .A(KEYINPUT56), .B(n1087), .Z(n1262) );
XNOR2_X1 U982 ( .A(n1281), .B(G478), .ZN(n1087) );
NAND2_X1 U983 ( .A1(n1163), .A2(n1200), .ZN(n1281) );
XOR2_X1 U984 ( .A(n1282), .B(n1283), .Z(n1163) );
XOR2_X1 U985 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U986 ( .A(G107), .B(G134), .ZN(n1285) );
NAND3_X1 U987 ( .A1(G217), .A2(n1286), .A3(KEYINPUT5), .ZN(n1284) );
XOR2_X1 U988 ( .A(n1287), .B(n1288), .Z(n1282) );
XOR2_X1 U989 ( .A(n1289), .B(n1277), .Z(n1288) );
NOR2_X1 U990 ( .A1(G116), .A2(KEYINPUT4), .ZN(n1289) );
AND3_X1 U991 ( .A1(n1253), .A2(n1078), .A3(n1055), .ZN(n1218) );
INV_X1 U992 ( .A(n1247), .ZN(n1055) );
NAND3_X1 U993 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1247) );
OR2_X1 U994 ( .A1(n1092), .A2(KEYINPUT38), .ZN(n1292) );
OR3_X1 U995 ( .A1(n1293), .A2(n1294), .A3(G469), .ZN(n1291) );
INV_X1 U996 ( .A(KEYINPUT38), .ZN(n1293) );
NAND2_X1 U997 ( .A1(G469), .A2(n1294), .ZN(n1290) );
NAND2_X1 U998 ( .A1(KEYINPUT42), .A2(n1092), .ZN(n1294) );
NAND2_X1 U999 ( .A1(n1295), .A2(n1200), .ZN(n1092) );
XNOR2_X1 U1000 ( .A(n1296), .B(n1192), .ZN(n1295) );
XNOR2_X1 U1001 ( .A(n1297), .B(n1298), .ZN(n1192) );
NAND2_X1 U1002 ( .A1(G227), .A2(n1138), .ZN(n1297) );
NAND2_X1 U1003 ( .A1(KEYINPUT11), .A2(n1191), .ZN(n1296) );
XNOR2_X1 U1004 ( .A(n1299), .B(n1300), .ZN(n1191) );
XOR2_X1 U1005 ( .A(n1301), .B(n1302), .Z(n1300) );
XNOR2_X1 U1006 ( .A(G101), .B(n1303), .ZN(n1302) );
NOR2_X1 U1007 ( .A1(KEYINPUT3), .A2(G107), .ZN(n1303) );
XNOR2_X1 U1008 ( .A(n1129), .B(n1278), .ZN(n1299) );
XOR2_X1 U1009 ( .A(n1304), .B(n1242), .Z(n1129) );
NAND3_X1 U1010 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1304) );
NAND2_X1 U1011 ( .A1(G143), .A2(n1308), .ZN(n1307) );
INV_X1 U1012 ( .A(KEYINPUT22), .ZN(n1308) );
NAND3_X1 U1013 ( .A1(KEYINPUT22), .A2(n1309), .A3(n1229), .ZN(n1306) );
OR2_X1 U1014 ( .A1(n1229), .A2(n1309), .ZN(n1305) );
NOR2_X1 U1015 ( .A1(G143), .A2(KEYINPUT0), .ZN(n1309) );
NAND2_X1 U1016 ( .A1(G221), .A2(n1310), .ZN(n1078) );
AND3_X1 U1017 ( .A1(n1063), .A2(n1311), .A3(n1249), .ZN(n1253) );
AND2_X1 U1018 ( .A1(n1059), .A2(n1312), .ZN(n1249) );
NAND2_X1 U1019 ( .A1(n1313), .A2(n1050), .ZN(n1312) );
NAND3_X1 U1020 ( .A1(G902), .A2(n1314), .A3(G953), .ZN(n1313) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1315), .ZN(n1059) );
NAND2_X1 U1022 ( .A1(G898), .A2(n1050), .ZN(n1311) );
NAND3_X1 U1023 ( .A1(n1314), .A2(n1138), .A3(G952), .ZN(n1050) );
NAND2_X1 U1024 ( .A1(G237), .A2(G234), .ZN(n1314) );
INV_X1 U1025 ( .A(n1057), .ZN(n1063) );
XOR2_X1 U1026 ( .A(n1107), .B(n1316), .Z(n1057) );
NOR2_X1 U1027 ( .A1(n1199), .A2(KEYINPUT41), .ZN(n1316) );
INV_X1 U1028 ( .A(n1106), .ZN(n1199) );
NAND2_X1 U1029 ( .A1(G210), .A2(n1315), .ZN(n1106) );
NAND2_X1 U1030 ( .A1(n1317), .A2(n1200), .ZN(n1315) );
INV_X1 U1031 ( .A(G237), .ZN(n1317) );
AND2_X1 U1032 ( .A1(n1318), .A2(n1200), .ZN(n1107) );
XNOR2_X1 U1033 ( .A(n1319), .B(n1320), .ZN(n1318) );
INV_X1 U1034 ( .A(n1198), .ZN(n1320) );
XOR2_X1 U1035 ( .A(n1321), .B(n1147), .Z(n1198) );
XOR2_X1 U1036 ( .A(n1257), .B(n1277), .Z(n1147) );
XOR2_X1 U1037 ( .A(G122), .B(KEYINPUT10), .Z(n1277) );
INV_X1 U1038 ( .A(G110), .ZN(n1257) );
XNOR2_X1 U1039 ( .A(n1146), .B(KEYINPUT26), .ZN(n1321) );
XNOR2_X1 U1040 ( .A(n1322), .B(n1323), .ZN(n1146) );
XNOR2_X1 U1041 ( .A(n1324), .B(n1278), .ZN(n1323) );
XOR2_X1 U1042 ( .A(G104), .B(KEYINPUT33), .Z(n1278) );
NAND2_X1 U1043 ( .A1(KEYINPUT59), .A2(n1272), .ZN(n1324) );
XOR2_X1 U1044 ( .A(n1325), .B(n1326), .Z(n1322) );
XOR2_X1 U1045 ( .A(G107), .B(G101), .Z(n1326) );
NAND3_X1 U1046 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1325) );
NAND2_X1 U1047 ( .A1(G116), .A2(n1330), .ZN(n1329) );
NAND2_X1 U1048 ( .A1(n1331), .A2(n1332), .ZN(n1328) );
INV_X1 U1049 ( .A(KEYINPUT27), .ZN(n1332) );
NAND2_X1 U1050 ( .A1(n1333), .A2(n1334), .ZN(n1331) );
XNOR2_X1 U1051 ( .A(KEYINPUT34), .B(n1330), .ZN(n1333) );
NAND2_X1 U1052 ( .A1(KEYINPUT27), .A2(n1335), .ZN(n1327) );
NAND2_X1 U1053 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
OR3_X1 U1054 ( .A1(n1330), .A2(G116), .A3(KEYINPUT34), .ZN(n1337) );
NAND2_X1 U1055 ( .A1(KEYINPUT34), .A2(n1330), .ZN(n1336) );
NAND2_X1 U1056 ( .A1(n1338), .A2(KEYINPUT55), .ZN(n1319) );
XNOR2_X1 U1057 ( .A(n1226), .B(n1227), .ZN(n1338) );
NAND2_X1 U1058 ( .A1(G224), .A2(n1138), .ZN(n1227) );
XNOR2_X1 U1059 ( .A(n1339), .B(G125), .ZN(n1226) );
AND2_X1 U1060 ( .A1(n1081), .A2(n1243), .ZN(n1072) );
XNOR2_X1 U1061 ( .A(n1100), .B(n1114), .ZN(n1243) );
NAND2_X1 U1062 ( .A1(G217), .A2(n1310), .ZN(n1114) );
NAND2_X1 U1063 ( .A1(G234), .A2(n1200), .ZN(n1310) );
NOR2_X1 U1064 ( .A1(n1158), .A2(G902), .ZN(n1100) );
XNOR2_X1 U1065 ( .A(n1340), .B(n1341), .ZN(n1158) );
XOR2_X1 U1066 ( .A(n1342), .B(n1343), .Z(n1341) );
XNOR2_X1 U1067 ( .A(n1298), .B(n1280), .ZN(n1343) );
XNOR2_X1 U1068 ( .A(n1229), .B(KEYINPUT54), .ZN(n1280) );
INV_X1 U1069 ( .A(G146), .ZN(n1229) );
XNOR2_X1 U1070 ( .A(G110), .B(n1136), .ZN(n1298) );
INV_X1 U1071 ( .A(G140), .ZN(n1136) );
NAND2_X1 U1072 ( .A1(n1344), .A2(n1345), .ZN(n1342) );
NAND2_X1 U1073 ( .A1(n1346), .A2(n1242), .ZN(n1345) );
INV_X1 U1074 ( .A(G128), .ZN(n1242) );
XNOR2_X1 U1075 ( .A(KEYINPUT20), .B(n1347), .ZN(n1346) );
NAND2_X1 U1076 ( .A1(n1348), .A2(G128), .ZN(n1344) );
XNOR2_X1 U1077 ( .A(KEYINPUT23), .B(n1347), .ZN(n1348) );
INV_X1 U1078 ( .A(n1330), .ZN(n1347) );
XOR2_X1 U1079 ( .A(n1349), .B(n1350), .Z(n1340) );
XOR2_X1 U1080 ( .A(n1351), .B(n1352), .Z(n1350) );
NOR2_X1 U1081 ( .A1(KEYINPUT13), .A2(n1134), .ZN(n1352) );
INV_X1 U1082 ( .A(G125), .ZN(n1134) );
NOR2_X1 U1083 ( .A1(G137), .A2(n1353), .ZN(n1351) );
XNOR2_X1 U1084 ( .A(KEYINPUT7), .B(KEYINPUT58), .ZN(n1353) );
NAND2_X1 U1085 ( .A1(n1286), .A2(G221), .ZN(n1349) );
AND2_X1 U1086 ( .A1(G234), .A2(n1138), .ZN(n1286) );
INV_X1 U1087 ( .A(G953), .ZN(n1138) );
INV_X1 U1088 ( .A(n1244), .ZN(n1081) );
XNOR2_X1 U1089 ( .A(n1354), .B(G472), .ZN(n1244) );
NAND2_X1 U1090 ( .A1(n1355), .A2(n1200), .ZN(n1354) );
INV_X1 U1091 ( .A(G902), .ZN(n1200) );
XNOR2_X1 U1092 ( .A(n1182), .B(n1356), .ZN(n1355) );
XOR2_X1 U1093 ( .A(n1357), .B(n1187), .Z(n1356) );
XNOR2_X1 U1094 ( .A(n1301), .B(n1339), .ZN(n1187) );
XNOR2_X1 U1095 ( .A(G146), .B(n1287), .ZN(n1339) );
XNOR2_X1 U1096 ( .A(G128), .B(G143), .ZN(n1287) );
NAND2_X1 U1097 ( .A1(n1358), .A2(n1359), .ZN(n1301) );
NAND2_X1 U1098 ( .A1(n1360), .A2(G131), .ZN(n1359) );
XOR2_X1 U1099 ( .A(KEYINPUT29), .B(n1361), .Z(n1358) );
NOR2_X1 U1100 ( .A1(G131), .A2(n1360), .ZN(n1361) );
XNOR2_X1 U1101 ( .A(G134), .B(n1362), .ZN(n1360) );
NOR2_X1 U1102 ( .A1(G137), .A2(KEYINPUT16), .ZN(n1362) );
NOR2_X1 U1103 ( .A1(KEYINPUT63), .A2(n1363), .ZN(n1357) );
XOR2_X1 U1104 ( .A(KEYINPUT25), .B(n1185), .Z(n1363) );
XNOR2_X1 U1105 ( .A(n1272), .B(n1364), .ZN(n1185) );
NOR2_X1 U1106 ( .A1(KEYINPUT62), .A2(n1365), .ZN(n1364) );
XNOR2_X1 U1107 ( .A(n1334), .B(n1330), .ZN(n1365) );
XOR2_X1 U1108 ( .A(G119), .B(KEYINPUT37), .Z(n1330) );
INV_X1 U1109 ( .A(G116), .ZN(n1334) );
INV_X1 U1110 ( .A(G113), .ZN(n1272) );
INV_X1 U1111 ( .A(n1178), .ZN(n1182) );
XNOR2_X1 U1112 ( .A(n1366), .B(G101), .ZN(n1178) );
NAND2_X1 U1113 ( .A1(n1273), .A2(G210), .ZN(n1366) );
NOR2_X1 U1114 ( .A1(G953), .A2(G237), .ZN(n1273) );
endmodule


