//Key = 1111001010100110001010010011100101111010000011010111010111011101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394;

XOR2_X1 U743 ( .A(n1056), .B(n1057), .Z(G9) );
NOR2_X1 U744 ( .A1(KEYINPUT17), .A2(n1058), .ZN(n1057) );
NOR3_X1 U745 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1056) );
NOR2_X1 U746 ( .A1(KEYINPUT34), .A2(n1062), .ZN(n1061) );
NOR3_X1 U747 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
AND2_X1 U748 ( .A1(n1066), .A2(KEYINPUT34), .ZN(n1060) );
NOR2_X1 U749 ( .A1(n1067), .A2(n1068), .ZN(G75) );
NOR4_X1 U750 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1068) );
XOR2_X1 U751 ( .A(n1073), .B(KEYINPUT47), .Z(n1072) );
NAND3_X1 U752 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
INV_X1 U753 ( .A(n1077), .ZN(n1076) );
NOR2_X1 U754 ( .A1(n1078), .A2(n1077), .ZN(n1071) );
NAND3_X1 U755 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1077) );
NOR3_X1 U756 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1078) );
AND3_X1 U757 ( .A1(KEYINPUT44), .A2(n1085), .A3(n1086), .ZN(n1084) );
AND2_X1 U758 ( .A1(n1087), .A2(n1075), .ZN(n1082) );
NAND4_X1 U759 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1069) );
NAND4_X1 U760 ( .A1(n1081), .A2(n1075), .A3(n1085), .A4(n1092), .ZN(n1089) );
NAND2_X1 U761 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U762 ( .A1(n1080), .A2(n1095), .ZN(n1094) );
NAND2_X1 U763 ( .A1(n1063), .A2(n1096), .ZN(n1095) );
NAND3_X1 U764 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
INV_X1 U765 ( .A(KEYINPUT48), .ZN(n1098) );
INV_X1 U766 ( .A(n1100), .ZN(n1063) );
NAND2_X1 U767 ( .A1(n1079), .A2(n1101), .ZN(n1093) );
NAND3_X1 U768 ( .A1(n1102), .A2(n1064), .A3(n1103), .ZN(n1101) );
NAND2_X1 U769 ( .A1(KEYINPUT48), .A2(n1080), .ZN(n1103) );
NAND2_X1 U770 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
XNOR2_X1 U771 ( .A(KEYINPUT59), .B(n1106), .ZN(n1105) );
XOR2_X1 U772 ( .A(n1107), .B(KEYINPUT27), .Z(n1104) );
NAND3_X1 U773 ( .A1(n1108), .A2(n1109), .A3(n1080), .ZN(n1088) );
INV_X1 U774 ( .A(KEYINPUT44), .ZN(n1109) );
NAND4_X1 U775 ( .A1(n1081), .A2(n1079), .A3(n1086), .A4(n1085), .ZN(n1108) );
INV_X1 U776 ( .A(n1110), .ZN(n1081) );
NOR3_X1 U777 ( .A1(n1111), .A2(G953), .A3(G952), .ZN(n1067) );
INV_X1 U778 ( .A(n1090), .ZN(n1111) );
NAND4_X1 U779 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1090) );
NOR4_X1 U780 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1115) );
XNOR2_X1 U781 ( .A(n1120), .B(KEYINPUT51), .ZN(n1117) );
XNOR2_X1 U782 ( .A(n1121), .B(KEYINPUT10), .ZN(n1116) );
AND3_X1 U783 ( .A1(n1107), .A2(n1122), .A3(n1123), .ZN(n1114) );
OR2_X1 U784 ( .A1(n1124), .A2(n1125), .ZN(n1113) );
XOR2_X1 U785 ( .A(n1126), .B(n1127), .Z(n1112) );
NAND2_X1 U786 ( .A1(KEYINPUT50), .A2(n1128), .ZN(n1127) );
XOR2_X1 U787 ( .A(n1129), .B(n1130), .Z(G72) );
NOR2_X1 U788 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U789 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U790 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U791 ( .A(n1137), .B(n1138), .Z(n1135) );
NAND3_X1 U792 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1137) );
NAND2_X1 U793 ( .A1(G140), .A2(n1142), .ZN(n1141) );
NAND2_X1 U794 ( .A1(KEYINPUT4), .A2(n1143), .ZN(n1140) );
NAND2_X1 U795 ( .A1(G125), .A2(n1144), .ZN(n1143) );
XNOR2_X1 U796 ( .A(KEYINPUT8), .B(n1145), .ZN(n1144) );
NAND2_X1 U797 ( .A1(n1146), .A2(n1147), .ZN(n1139) );
INV_X1 U798 ( .A(KEYINPUT4), .ZN(n1147) );
NAND2_X1 U799 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
NAND3_X1 U800 ( .A1(KEYINPUT8), .A2(G125), .A3(n1145), .ZN(n1149) );
OR2_X1 U801 ( .A1(n1145), .A2(KEYINPUT8), .ZN(n1148) );
XOR2_X1 U802 ( .A(n1150), .B(n1151), .Z(n1133) );
XOR2_X1 U803 ( .A(KEYINPUT11), .B(G143), .Z(n1151) );
XNOR2_X1 U804 ( .A(G134), .B(G137), .ZN(n1150) );
NAND2_X1 U805 ( .A1(n1152), .A2(n1153), .ZN(n1129) );
NAND2_X1 U806 ( .A1(n1154), .A2(n1091), .ZN(n1153) );
NAND2_X1 U807 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND2_X1 U808 ( .A1(KEYINPUT45), .A2(n1157), .ZN(n1152) );
NAND2_X1 U809 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U810 ( .A1(G953), .A2(n1160), .ZN(n1159) );
INV_X1 U811 ( .A(n1131), .ZN(n1158) );
NAND2_X1 U812 ( .A1(n1161), .A2(n1162), .ZN(G69) );
NAND4_X1 U813 ( .A1(KEYINPUT28), .A2(G953), .A3(n1163), .A4(n1164), .ZN(n1162) );
NAND2_X1 U814 ( .A1(n1165), .A2(n1166), .ZN(n1161) );
NAND2_X1 U815 ( .A1(G953), .A2(n1163), .ZN(n1166) );
NAND2_X1 U816 ( .A1(G898), .A2(G224), .ZN(n1163) );
XOR2_X1 U817 ( .A(n1167), .B(n1168), .Z(n1165) );
AND2_X1 U818 ( .A1(n1164), .A2(KEYINPUT28), .ZN(n1168) );
NAND4_X1 U819 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1164) );
NAND2_X1 U820 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XNOR2_X1 U821 ( .A(n1175), .B(n1176), .ZN(n1173) );
NAND3_X1 U822 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1171) );
NAND2_X1 U823 ( .A1(G953), .A2(n1179), .ZN(n1169) );
NAND2_X1 U824 ( .A1(n1180), .A2(n1091), .ZN(n1167) );
NAND2_X1 U825 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NOR2_X1 U826 ( .A1(n1183), .A2(n1184), .ZN(G66) );
XOR2_X1 U827 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U828 ( .A1(n1187), .A2(n1188), .ZN(n1185) );
NOR2_X1 U829 ( .A1(n1183), .A2(n1189), .ZN(G63) );
XOR2_X1 U830 ( .A(n1190), .B(n1191), .Z(n1189) );
NOR2_X1 U831 ( .A1(n1124), .A2(n1188), .ZN(n1190) );
NOR2_X1 U832 ( .A1(n1183), .A2(n1192), .ZN(G60) );
NOR2_X1 U833 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NOR2_X1 U834 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NOR2_X1 U835 ( .A1(n1197), .A2(n1198), .ZN(n1193) );
XOR2_X1 U836 ( .A(KEYINPUT38), .B(n1195), .Z(n1198) );
AND2_X1 U837 ( .A1(n1199), .A2(G475), .ZN(n1195) );
XNOR2_X1 U838 ( .A(n1196), .B(KEYINPUT16), .ZN(n1197) );
XNOR2_X1 U839 ( .A(G104), .B(n1200), .ZN(G6) );
NAND4_X1 U840 ( .A1(KEYINPUT18), .A2(n1201), .A3(n1086), .A4(n1202), .ZN(n1200) );
XOR2_X1 U841 ( .A(KEYINPUT24), .B(n1085), .Z(n1202) );
NOR2_X1 U842 ( .A1(n1183), .A2(n1203), .ZN(G57) );
XOR2_X1 U843 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U844 ( .A(n1206), .B(n1207), .Z(n1205) );
NAND2_X1 U845 ( .A1(n1208), .A2(n1209), .ZN(n1206) );
XOR2_X1 U846 ( .A(n1210), .B(n1211), .Z(n1209) );
NAND3_X1 U847 ( .A1(n1212), .A2(n1213), .A3(KEYINPUT1), .ZN(n1211) );
NAND2_X1 U848 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
INV_X1 U849 ( .A(KEYINPUT29), .ZN(n1215) );
XNOR2_X1 U850 ( .A(n1216), .B(n1217), .ZN(n1214) );
NAND2_X1 U851 ( .A1(n1218), .A2(KEYINPUT29), .ZN(n1212) );
XOR2_X1 U852 ( .A(n1219), .B(n1220), .Z(n1218) );
XNOR2_X1 U853 ( .A(KEYINPUT35), .B(KEYINPUT33), .ZN(n1208) );
XOR2_X1 U854 ( .A(n1221), .B(KEYINPUT40), .Z(n1204) );
NAND3_X1 U855 ( .A1(n1222), .A2(n1223), .A3(G472), .ZN(n1221) );
OR2_X1 U856 ( .A1(n1199), .A2(KEYINPUT19), .ZN(n1223) );
INV_X1 U857 ( .A(n1188), .ZN(n1199) );
NAND2_X1 U858 ( .A1(KEYINPUT19), .A2(n1224), .ZN(n1222) );
OR2_X1 U859 ( .A1(n1070), .A2(n1225), .ZN(n1224) );
NOR2_X1 U860 ( .A1(n1183), .A2(n1226), .ZN(G54) );
XOR2_X1 U861 ( .A(n1227), .B(n1228), .Z(n1226) );
XOR2_X1 U862 ( .A(KEYINPUT43), .B(n1229), .Z(n1228) );
NOR2_X1 U863 ( .A1(n1128), .A2(n1188), .ZN(n1229) );
NOR2_X1 U864 ( .A1(n1183), .A2(n1230), .ZN(G51) );
XOR2_X1 U865 ( .A(n1231), .B(n1232), .Z(n1230) );
XNOR2_X1 U866 ( .A(n1233), .B(n1234), .ZN(n1232) );
XOR2_X1 U867 ( .A(n1219), .B(KEYINPUT52), .Z(n1234) );
XOR2_X1 U868 ( .A(n1235), .B(n1236), .Z(n1231) );
XOR2_X1 U869 ( .A(n1237), .B(n1238), .Z(n1235) );
NOR2_X1 U870 ( .A1(n1239), .A2(n1188), .ZN(n1238) );
NAND2_X1 U871 ( .A1(G902), .A2(n1070), .ZN(n1188) );
NAND4_X1 U872 ( .A1(n1155), .A2(n1181), .A3(n1240), .A4(n1241), .ZN(n1070) );
XOR2_X1 U873 ( .A(KEYINPUT9), .B(n1156), .Z(n1241) );
NOR4_X1 U874 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1156) );
INV_X1 U875 ( .A(n1246), .ZN(n1243) );
XNOR2_X1 U876 ( .A(KEYINPUT3), .B(n1182), .ZN(n1240) );
NAND3_X1 U877 ( .A1(n1086), .A2(n1085), .A3(n1201), .ZN(n1182) );
AND4_X1 U878 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1181) );
NOR4_X1 U879 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1250) );
NOR2_X1 U880 ( .A1(n1064), .A2(n1255), .ZN(n1254) );
XNOR2_X1 U881 ( .A(KEYINPUT2), .B(n1256), .ZN(n1255) );
NOR2_X1 U882 ( .A1(n1257), .A2(n1066), .ZN(n1253) );
NOR2_X1 U883 ( .A1(n1258), .A2(n1083), .ZN(n1257) );
INV_X1 U884 ( .A(n1059), .ZN(n1083) );
NAND2_X1 U885 ( .A1(n1259), .A2(n1085), .ZN(n1059) );
NOR2_X1 U886 ( .A1(n1260), .A2(n1261), .ZN(n1258) );
XNOR2_X1 U887 ( .A(n1087), .B(KEYINPUT30), .ZN(n1260) );
AND3_X1 U888 ( .A1(KEYINPUT39), .A2(n1262), .A3(n1263), .ZN(n1252) );
INV_X1 U889 ( .A(n1086), .ZN(n1262) );
NOR2_X1 U890 ( .A1(KEYINPUT39), .A2(n1264), .ZN(n1251) );
AND3_X1 U891 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1155) );
NAND2_X1 U892 ( .A1(n1080), .A2(n1268), .ZN(n1267) );
NAND2_X1 U893 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
NAND2_X1 U894 ( .A1(n1075), .A2(n1271), .ZN(n1270) );
NAND2_X1 U895 ( .A1(n1272), .A2(n1100), .ZN(n1269) );
NOR2_X1 U896 ( .A1(n1091), .A2(G952), .ZN(n1183) );
XNOR2_X1 U897 ( .A(G146), .B(n1265), .ZN(G48) );
NAND3_X1 U898 ( .A1(n1271), .A2(n1273), .A3(n1086), .ZN(n1265) );
XNOR2_X1 U899 ( .A(G143), .B(n1266), .ZN(G45) );
NAND4_X1 U900 ( .A1(n1274), .A2(n1273), .A3(n1120), .A4(n1275), .ZN(n1266) );
XNOR2_X1 U901 ( .A(G140), .B(n1276), .ZN(G42) );
NAND4_X1 U902 ( .A1(KEYINPUT14), .A2(n1272), .A3(n1100), .A4(n1080), .ZN(n1276) );
XNOR2_X1 U903 ( .A(G137), .B(n1277), .ZN(G39) );
NAND2_X1 U904 ( .A1(n1278), .A2(n1080), .ZN(n1277) );
XOR2_X1 U905 ( .A(KEYINPUT21), .B(n1279), .Z(n1278) );
NOR2_X1 U906 ( .A1(n1280), .A2(n1261), .ZN(n1279) );
INV_X1 U907 ( .A(n1075), .ZN(n1261) );
XOR2_X1 U908 ( .A(n1281), .B(G134), .Z(G36) );
NAND2_X1 U909 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U910 ( .A1(n1242), .A2(n1284), .ZN(n1283) );
INV_X1 U911 ( .A(KEYINPUT42), .ZN(n1284) );
NOR2_X1 U912 ( .A1(n1285), .A2(n1286), .ZN(n1242) );
INV_X1 U913 ( .A(n1080), .ZN(n1286) );
NAND3_X1 U914 ( .A1(n1080), .A2(n1285), .A3(KEYINPUT42), .ZN(n1282) );
NAND2_X1 U915 ( .A1(n1274), .A2(n1259), .ZN(n1285) );
XNOR2_X1 U916 ( .A(G131), .B(n1246), .ZN(G33) );
NAND3_X1 U917 ( .A1(n1274), .A2(n1080), .A3(n1086), .ZN(n1246) );
NAND2_X1 U918 ( .A1(n1287), .A2(n1288), .ZN(n1080) );
OR2_X1 U919 ( .A1(n1064), .A2(KEYINPUT59), .ZN(n1288) );
NAND3_X1 U920 ( .A1(n1106), .A2(n1107), .A3(KEYINPUT59), .ZN(n1287) );
INV_X1 U921 ( .A(n1121), .ZN(n1106) );
AND3_X1 U922 ( .A1(n1100), .A2(n1289), .A3(n1087), .ZN(n1274) );
XOR2_X1 U923 ( .A(G128), .B(n1244), .Z(G30) );
AND3_X1 U924 ( .A1(n1273), .A2(n1259), .A3(n1271), .ZN(n1244) );
INV_X1 U925 ( .A(n1280), .ZN(n1271) );
NAND4_X1 U926 ( .A1(n1100), .A2(n1290), .A3(n1289), .A4(n1118), .ZN(n1280) );
XNOR2_X1 U927 ( .A(G101), .B(n1291), .ZN(G3) );
NAND3_X1 U928 ( .A1(n1075), .A2(n1087), .A3(n1201), .ZN(n1291) );
INV_X1 U929 ( .A(n1066), .ZN(n1201) );
NAND3_X1 U930 ( .A1(n1273), .A2(n1065), .A3(n1100), .ZN(n1066) );
NAND2_X1 U931 ( .A1(n1292), .A2(n1293), .ZN(G27) );
NAND2_X1 U932 ( .A1(n1245), .A2(n1142), .ZN(n1293) );
INV_X1 U933 ( .A(n1294), .ZN(n1245) );
XOR2_X1 U934 ( .A(n1295), .B(KEYINPUT15), .Z(n1292) );
NAND2_X1 U935 ( .A1(G125), .A2(n1294), .ZN(n1295) );
NAND3_X1 U936 ( .A1(n1272), .A2(n1273), .A3(n1079), .ZN(n1294) );
AND3_X1 U937 ( .A1(n1086), .A2(n1289), .A3(n1074), .ZN(n1272) );
NAND2_X1 U938 ( .A1(n1110), .A2(n1296), .ZN(n1289) );
NAND3_X1 U939 ( .A1(G902), .A2(n1297), .A3(n1131), .ZN(n1296) );
NOR2_X1 U940 ( .A1(G900), .A2(n1091), .ZN(n1131) );
XNOR2_X1 U941 ( .A(G122), .B(n1249), .ZN(G24) );
NAND4_X1 U942 ( .A1(n1298), .A2(n1085), .A3(n1120), .A4(n1275), .ZN(n1249) );
NOR2_X1 U943 ( .A1(n1118), .A2(n1290), .ZN(n1085) );
XNOR2_X1 U944 ( .A(G119), .B(n1247), .ZN(G21) );
NAND4_X1 U945 ( .A1(n1298), .A2(n1075), .A3(n1290), .A4(n1118), .ZN(n1247) );
XNOR2_X1 U946 ( .A(n1299), .B(n1248), .ZN(G18) );
NAND2_X1 U947 ( .A1(n1263), .A2(n1259), .ZN(n1248) );
AND2_X1 U948 ( .A1(n1300), .A2(n1275), .ZN(n1259) );
XNOR2_X1 U949 ( .A(G116), .B(KEYINPUT61), .ZN(n1299) );
XOR2_X1 U950 ( .A(n1264), .B(n1301), .Z(G15) );
NAND2_X1 U951 ( .A1(KEYINPUT53), .A2(G113), .ZN(n1301) );
NAND2_X1 U952 ( .A1(n1263), .A2(n1086), .ZN(n1264) );
NOR2_X1 U953 ( .A1(n1275), .A2(n1300), .ZN(n1086) );
INV_X1 U954 ( .A(n1120), .ZN(n1300) );
AND2_X1 U955 ( .A1(n1298), .A2(n1087), .ZN(n1263) );
NOR2_X1 U956 ( .A1(n1118), .A2(n1302), .ZN(n1087) );
AND3_X1 U957 ( .A1(n1273), .A2(n1065), .A3(n1079), .ZN(n1298) );
AND2_X1 U958 ( .A1(n1097), .A2(n1123), .ZN(n1079) );
INV_X1 U959 ( .A(n1064), .ZN(n1273) );
XNOR2_X1 U960 ( .A(n1303), .B(n1304), .ZN(G12) );
NOR2_X1 U961 ( .A1(n1064), .A2(n1256), .ZN(n1304) );
NAND4_X1 U962 ( .A1(n1074), .A2(n1075), .A3(n1100), .A4(n1065), .ZN(n1256) );
NAND2_X1 U963 ( .A1(n1110), .A2(n1305), .ZN(n1065) );
NAND4_X1 U964 ( .A1(G953), .A2(G902), .A3(n1297), .A4(n1179), .ZN(n1305) );
INV_X1 U965 ( .A(G898), .ZN(n1179) );
NAND3_X1 U966 ( .A1(n1297), .A2(n1091), .A3(G952), .ZN(n1110) );
NAND2_X1 U967 ( .A1(G237), .A2(G234), .ZN(n1297) );
NOR2_X1 U968 ( .A1(n1097), .A2(n1099), .ZN(n1100) );
INV_X1 U969 ( .A(n1123), .ZN(n1099) );
NAND2_X1 U970 ( .A1(G221), .A2(n1306), .ZN(n1123) );
NAND2_X1 U971 ( .A1(G234), .A2(n1225), .ZN(n1306) );
XOR2_X1 U972 ( .A(n1307), .B(n1128), .Z(n1097) );
INV_X1 U973 ( .A(G469), .ZN(n1128) );
NAND2_X1 U974 ( .A1(KEYINPUT31), .A2(n1308), .ZN(n1307) );
XNOR2_X1 U975 ( .A(KEYINPUT26), .B(n1126), .ZN(n1308) );
NAND2_X1 U976 ( .A1(n1309), .A2(n1225), .ZN(n1126) );
XOR2_X1 U977 ( .A(n1227), .B(n1310), .Z(n1309) );
XOR2_X1 U978 ( .A(KEYINPUT49), .B(KEYINPUT41), .Z(n1310) );
XOR2_X1 U979 ( .A(n1311), .B(n1312), .Z(n1227) );
XOR2_X1 U980 ( .A(n1313), .B(n1314), .Z(n1312) );
XNOR2_X1 U981 ( .A(n1303), .B(G101), .ZN(n1314) );
NOR2_X1 U982 ( .A1(G953), .A2(n1160), .ZN(n1313) );
INV_X1 U983 ( .A(G227), .ZN(n1160) );
XOR2_X1 U984 ( .A(n1315), .B(n1316), .Z(n1311) );
XOR2_X1 U985 ( .A(n1220), .B(n1317), .Z(n1315) );
XOR2_X1 U986 ( .A(n1216), .B(n1138), .Z(n1220) );
NOR2_X1 U987 ( .A1(n1275), .A2(n1120), .ZN(n1075) );
XNOR2_X1 U988 ( .A(n1318), .B(G475), .ZN(n1120) );
NAND2_X1 U989 ( .A1(n1319), .A2(n1225), .ZN(n1318) );
INV_X1 U990 ( .A(n1196), .ZN(n1319) );
XNOR2_X1 U991 ( .A(n1320), .B(n1321), .ZN(n1196) );
XOR2_X1 U992 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U993 ( .A(n1324), .B(G122), .Z(n1323) );
NAND2_X1 U994 ( .A1(G214), .A2(n1325), .ZN(n1324) );
XNOR2_X1 U995 ( .A(G131), .B(G125), .ZN(n1322) );
XOR2_X1 U996 ( .A(n1326), .B(n1327), .Z(n1320) );
XNOR2_X1 U997 ( .A(n1328), .B(n1329), .ZN(n1327) );
NOR2_X1 U998 ( .A1(KEYINPUT58), .A2(n1330), .ZN(n1329) );
INV_X1 U999 ( .A(G104), .ZN(n1330) );
NAND2_X1 U1000 ( .A1(KEYINPUT63), .A2(n1331), .ZN(n1328) );
XOR2_X1 U1001 ( .A(n1332), .B(n1316), .Z(n1326) );
XNOR2_X1 U1002 ( .A(G143), .B(n1145), .ZN(n1316) );
NAND2_X1 U1003 ( .A1(KEYINPUT57), .A2(G113), .ZN(n1332) );
NAND3_X1 U1004 ( .A1(n1333), .A2(n1334), .A3(n1122), .ZN(n1275) );
NAND2_X1 U1005 ( .A1(n1125), .A2(n1124), .ZN(n1122) );
OR3_X1 U1006 ( .A1(n1124), .A2(n1125), .A3(KEYINPUT5), .ZN(n1334) );
NOR2_X1 U1007 ( .A1(n1191), .A2(G902), .ZN(n1125) );
XNOR2_X1 U1008 ( .A(n1335), .B(n1336), .ZN(n1191) );
XOR2_X1 U1009 ( .A(G128), .B(n1337), .Z(n1336) );
XOR2_X1 U1010 ( .A(G143), .B(G134), .Z(n1337) );
XNOR2_X1 U1011 ( .A(n1338), .B(n1339), .ZN(n1335) );
NAND3_X1 U1012 ( .A1(G217), .A2(n1340), .A3(KEYINPUT55), .ZN(n1339) );
NAND2_X1 U1013 ( .A1(n1341), .A2(KEYINPUT20), .ZN(n1338) );
XNOR2_X1 U1014 ( .A(G107), .B(n1342), .ZN(n1341) );
XNOR2_X1 U1015 ( .A(G122), .B(n1343), .ZN(n1342) );
NAND2_X1 U1016 ( .A1(KEYINPUT5), .A2(n1124), .ZN(n1333) );
INV_X1 U1017 ( .A(G478), .ZN(n1124) );
AND2_X1 U1018 ( .A1(n1302), .A2(n1118), .ZN(n1074) );
NAND3_X1 U1019 ( .A1(n1344), .A2(n1345), .A3(n1346), .ZN(n1118) );
NAND2_X1 U1020 ( .A1(n1347), .A2(n1186), .ZN(n1346) );
OR3_X1 U1021 ( .A1(n1186), .A2(n1347), .A3(G902), .ZN(n1345) );
NOR2_X1 U1022 ( .A1(n1187), .A2(G234), .ZN(n1347) );
INV_X1 U1023 ( .A(G217), .ZN(n1187) );
XNOR2_X1 U1024 ( .A(n1348), .B(n1349), .ZN(n1186) );
XNOR2_X1 U1025 ( .A(n1350), .B(n1351), .ZN(n1349) );
XNOR2_X1 U1026 ( .A(n1145), .B(G137), .ZN(n1351) );
INV_X1 U1027 ( .A(G140), .ZN(n1145) );
XNOR2_X1 U1028 ( .A(n1236), .B(n1352), .ZN(n1348) );
XOR2_X1 U1029 ( .A(n1353), .B(n1354), .Z(n1352) );
NAND2_X1 U1030 ( .A1(G221), .A2(n1340), .ZN(n1354) );
AND2_X1 U1031 ( .A1(G234), .A2(n1091), .ZN(n1340) );
NAND2_X1 U1032 ( .A1(KEYINPUT36), .A2(n1355), .ZN(n1353) );
XNOR2_X1 U1033 ( .A(KEYINPUT60), .B(n1303), .ZN(n1355) );
XOR2_X1 U1034 ( .A(G125), .B(n1138), .Z(n1236) );
NAND2_X1 U1035 ( .A1(G902), .A2(G217), .ZN(n1344) );
INV_X1 U1036 ( .A(n1290), .ZN(n1302) );
XOR2_X1 U1037 ( .A(n1119), .B(KEYINPUT54), .Z(n1290) );
XNOR2_X1 U1038 ( .A(n1356), .B(G472), .ZN(n1119) );
NAND2_X1 U1039 ( .A1(n1357), .A2(n1225), .ZN(n1356) );
XOR2_X1 U1040 ( .A(n1358), .B(n1359), .Z(n1357) );
XNOR2_X1 U1041 ( .A(n1210), .B(n1360), .ZN(n1359) );
NOR2_X1 U1042 ( .A1(KEYINPUT12), .A2(n1217), .ZN(n1360) );
NAND2_X1 U1043 ( .A1(n1361), .A2(n1362), .ZN(n1210) );
NAND2_X1 U1044 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
XOR2_X1 U1045 ( .A(n1365), .B(KEYINPUT22), .Z(n1361) );
OR2_X1 U1046 ( .A1(n1364), .A2(n1363), .ZN(n1365) );
XNOR2_X1 U1047 ( .A(G116), .B(n1350), .ZN(n1363) );
XOR2_X1 U1048 ( .A(n1216), .B(n1207), .Z(n1358) );
XNOR2_X1 U1049 ( .A(n1366), .B(G101), .ZN(n1207) );
NAND2_X1 U1050 ( .A1(G210), .A2(n1325), .ZN(n1366) );
NOR2_X1 U1051 ( .A1(G953), .A2(G237), .ZN(n1325) );
XOR2_X1 U1052 ( .A(n1367), .B(n1136), .Z(n1216) );
XNOR2_X1 U1053 ( .A(n1368), .B(KEYINPUT13), .ZN(n1136) );
INV_X1 U1054 ( .A(G131), .ZN(n1368) );
NAND2_X1 U1055 ( .A1(n1369), .A2(n1370), .ZN(n1367) );
NAND2_X1 U1056 ( .A1(G134), .A2(n1371), .ZN(n1370) );
XOR2_X1 U1057 ( .A(KEYINPUT56), .B(n1372), .Z(n1369) );
NOR2_X1 U1058 ( .A1(G134), .A2(n1371), .ZN(n1372) );
INV_X1 U1059 ( .A(G137), .ZN(n1371) );
NAND2_X1 U1060 ( .A1(n1121), .A2(n1107), .ZN(n1064) );
NAND2_X1 U1061 ( .A1(G214), .A2(n1373), .ZN(n1107) );
XOR2_X1 U1062 ( .A(n1374), .B(n1239), .Z(n1121) );
NAND2_X1 U1063 ( .A1(G210), .A2(n1373), .ZN(n1239) );
NAND2_X1 U1064 ( .A1(n1375), .A2(n1225), .ZN(n1373) );
XNOR2_X1 U1065 ( .A(G237), .B(KEYINPUT7), .ZN(n1375) );
NAND2_X1 U1066 ( .A1(n1376), .A2(n1225), .ZN(n1374) );
INV_X1 U1067 ( .A(G902), .ZN(n1225) );
XOR2_X1 U1068 ( .A(n1377), .B(n1378), .Z(n1376) );
XOR2_X1 U1069 ( .A(n1237), .B(n1379), .Z(n1378) );
NAND2_X1 U1070 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
NAND2_X1 U1071 ( .A1(n1217), .A2(n1382), .ZN(n1381) );
NAND2_X1 U1072 ( .A1(KEYINPUT0), .A2(n1383), .ZN(n1382) );
NAND2_X1 U1073 ( .A1(KEYINPUT23), .A2(G125), .ZN(n1383) );
INV_X1 U1074 ( .A(n1384), .ZN(n1217) );
NAND2_X1 U1075 ( .A1(n1385), .A2(n1142), .ZN(n1380) );
INV_X1 U1076 ( .A(G125), .ZN(n1142) );
NAND2_X1 U1077 ( .A1(KEYINPUT23), .A2(n1386), .ZN(n1385) );
NAND2_X1 U1078 ( .A1(KEYINPUT0), .A2(n1384), .ZN(n1386) );
XNOR2_X1 U1079 ( .A(n1219), .B(n1138), .ZN(n1384) );
XNOR2_X1 U1080 ( .A(G128), .B(n1331), .ZN(n1138) );
INV_X1 U1081 ( .A(G146), .ZN(n1331) );
OR2_X1 U1082 ( .A1(KEYINPUT25), .A2(G143), .ZN(n1219) );
NAND2_X1 U1083 ( .A1(G224), .A2(n1091), .ZN(n1237) );
INV_X1 U1084 ( .A(G953), .ZN(n1091) );
NOR2_X1 U1085 ( .A1(n1233), .A2(KEYINPUT37), .ZN(n1377) );
AND3_X1 U1086 ( .A1(n1387), .A2(n1388), .A3(n1170), .ZN(n1233) );
OR3_X1 U1087 ( .A1(n1177), .A2(n1174), .A3(n1176), .ZN(n1170) );
NAND2_X1 U1088 ( .A1(n1389), .A2(n1177), .ZN(n1388) );
INV_X1 U1089 ( .A(n1175), .ZN(n1177) );
XOR2_X1 U1090 ( .A(n1176), .B(n1390), .Z(n1389) );
NOR2_X1 U1091 ( .A1(KEYINPUT46), .A2(n1178), .ZN(n1390) );
NAND3_X1 U1092 ( .A1(n1391), .A2(n1174), .A3(n1175), .ZN(n1387) );
XOR2_X1 U1093 ( .A(G110), .B(G122), .Z(n1175) );
INV_X1 U1094 ( .A(n1178), .ZN(n1174) );
XOR2_X1 U1095 ( .A(n1317), .B(n1392), .Z(n1178) );
NOR2_X1 U1096 ( .A1(G101), .A2(KEYINPUT32), .ZN(n1392) );
XNOR2_X1 U1097 ( .A(G104), .B(n1058), .ZN(n1317) );
INV_X1 U1098 ( .A(G107), .ZN(n1058) );
XOR2_X1 U1099 ( .A(n1176), .B(KEYINPUT46), .Z(n1391) );
XOR2_X1 U1100 ( .A(n1393), .B(n1364), .Z(n1176) );
XOR2_X1 U1101 ( .A(G113), .B(KEYINPUT62), .Z(n1364) );
XNOR2_X1 U1102 ( .A(n1394), .B(n1350), .ZN(n1393) );
INV_X1 U1103 ( .A(G119), .ZN(n1350) );
NAND2_X1 U1104 ( .A1(KEYINPUT6), .A2(n1343), .ZN(n1394) );
INV_X1 U1105 ( .A(G116), .ZN(n1343) );
INV_X1 U1106 ( .A(G110), .ZN(n1303) );
endmodule


