//Key = 0111100001010010100100110100000100000001010111101011011111111111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370;

XNOR2_X1 U751 ( .A(n1039), .B(n1040), .ZN(G9) );
NOR3_X1 U752 ( .A1(n1041), .A2(KEYINPUT35), .A3(n1042), .ZN(n1040) );
NOR2_X1 U753 ( .A1(n1043), .A2(n1044), .ZN(G75) );
XOR2_X1 U754 ( .A(n1045), .B(KEYINPUT50), .Z(n1044) );
NAND4_X1 U755 ( .A1(G952), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1045) );
NOR3_X1 U756 ( .A1(n1049), .A2(G953), .A3(n1050), .ZN(n1048) );
NOR3_X1 U757 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1049) );
NOR2_X1 U758 ( .A1(KEYINPUT3), .A2(n1054), .ZN(n1053) );
NAND4_X1 U759 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NOR2_X1 U760 ( .A1(n1059), .A2(n1060), .ZN(n1052) );
INV_X1 U761 ( .A(KEYINPUT3), .ZN(n1060) );
NOR4_X1 U762 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1059) );
NOR2_X1 U763 ( .A1(n1057), .A2(n1065), .ZN(n1061) );
INV_X1 U764 ( .A(n1066), .ZN(n1051) );
NAND3_X1 U765 ( .A1(n1067), .A2(n1068), .A3(n1055), .ZN(n1046) );
INV_X1 U766 ( .A(n1064), .ZN(n1055) );
NAND2_X1 U767 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U768 ( .A1(n1066), .A2(n1071), .ZN(n1070) );
NAND2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U770 ( .A1(n1056), .A2(n1074), .ZN(n1073) );
OR2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U772 ( .A1(n1058), .A2(n1077), .ZN(n1072) );
NAND2_X1 U773 ( .A1(n1058), .A2(n1078), .ZN(n1069) );
NAND2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND3_X1 U775 ( .A1(n1077), .A2(n1081), .A3(n1082), .ZN(n1080) );
INV_X1 U776 ( .A(KEYINPUT39), .ZN(n1081) );
NAND3_X1 U777 ( .A1(n1083), .A2(n1084), .A3(n1066), .ZN(n1077) );
NAND2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U779 ( .A1(KEYINPUT39), .A2(n1082), .ZN(n1083) );
NAND2_X1 U780 ( .A1(n1056), .A2(n1087), .ZN(n1079) );
NAND2_X1 U781 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U782 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR3_X1 U783 ( .A1(n1092), .A2(G953), .A3(n1093), .ZN(n1043) );
XNOR2_X1 U784 ( .A(G952), .B(KEYINPUT59), .ZN(n1093) );
XNOR2_X1 U785 ( .A(n1050), .B(KEYINPUT56), .ZN(n1092) );
AND4_X1 U786 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1050) );
NOR4_X1 U787 ( .A1(n1063), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1097) );
XNOR2_X1 U788 ( .A(KEYINPUT15), .B(n1091), .ZN(n1100) );
XNOR2_X1 U789 ( .A(KEYINPUT30), .B(n1101), .ZN(n1099) );
NOR3_X1 U790 ( .A1(n1102), .A2(n1103), .A3(n1090), .ZN(n1096) );
NAND2_X1 U791 ( .A1(n1104), .A2(n1105), .ZN(n1095) );
XNOR2_X1 U792 ( .A(n1106), .B(n1107), .ZN(n1104) );
XNOR2_X1 U793 ( .A(KEYINPUT38), .B(KEYINPUT1), .ZN(n1106) );
XOR2_X1 U794 ( .A(n1108), .B(n1109), .Z(G72) );
NOR2_X1 U795 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U796 ( .A(KEYINPUT20), .B(n1112), .Z(n1111) );
NOR2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1108) );
NAND2_X1 U799 ( .A1(n1117), .A2(n1110), .ZN(n1116) );
XNOR2_X1 U800 ( .A(n1118), .B(n1119), .ZN(n1117) );
NAND3_X1 U801 ( .A1(G900), .A2(n1118), .A3(G953), .ZN(n1115) );
XNOR2_X1 U802 ( .A(n1120), .B(n1121), .ZN(n1118) );
XNOR2_X1 U803 ( .A(n1122), .B(n1123), .ZN(n1121) );
NOR2_X1 U804 ( .A1(KEYINPUT5), .A2(G137), .ZN(n1123) );
NAND2_X1 U805 ( .A1(n1124), .A2(KEYINPUT45), .ZN(n1122) );
XNOR2_X1 U806 ( .A(G125), .B(G140), .ZN(n1124) );
XOR2_X1 U807 ( .A(n1125), .B(n1126), .Z(n1120) );
NAND2_X1 U808 ( .A1(n1127), .A2(n1128), .ZN(G69) );
NAND2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND3_X1 U810 ( .A1(n1131), .A2(n1132), .A3(G953), .ZN(n1130) );
NAND3_X1 U811 ( .A1(n1133), .A2(n1132), .A3(n1134), .ZN(n1127) );
INV_X1 U812 ( .A(n1129), .ZN(n1134) );
XNOR2_X1 U813 ( .A(n1135), .B(n1136), .ZN(n1129) );
NOR3_X1 U814 ( .A1(n1137), .A2(KEYINPUT28), .A3(G953), .ZN(n1136) );
AND2_X1 U815 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NAND2_X1 U816 ( .A1(n1140), .A2(n1141), .ZN(n1135) );
XOR2_X1 U817 ( .A(n1142), .B(n1143), .Z(n1140) );
NAND2_X1 U818 ( .A1(n1144), .A2(n1145), .ZN(n1142) );
NAND2_X1 U819 ( .A1(KEYINPUT48), .A2(n1146), .ZN(n1145) );
XNOR2_X1 U820 ( .A(n1147), .B(n1148), .ZN(n1146) );
NAND3_X1 U821 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1144) );
INV_X1 U822 ( .A(KEYINPUT48), .ZN(n1151) );
XNOR2_X1 U823 ( .A(n1147), .B(n1152), .ZN(n1149) );
INV_X1 U824 ( .A(KEYINPUT10), .ZN(n1132) );
NAND2_X1 U825 ( .A1(n1141), .A2(n1153), .ZN(n1133) );
NAND2_X1 U826 ( .A1(G953), .A2(n1131), .ZN(n1153) );
INV_X1 U827 ( .A(n1154), .ZN(n1141) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1156), .ZN(G66) );
XOR2_X1 U829 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U830 ( .A1(n1159), .A2(G217), .ZN(n1157) );
NOR2_X1 U831 ( .A1(n1155), .A2(n1160), .ZN(G63) );
XOR2_X1 U832 ( .A(n1161), .B(n1162), .Z(n1160) );
NAND2_X1 U833 ( .A1(n1159), .A2(G478), .ZN(n1161) );
NOR2_X1 U834 ( .A1(n1155), .A2(n1163), .ZN(G60) );
XNOR2_X1 U835 ( .A(n1164), .B(n1165), .ZN(n1163) );
NOR3_X1 U836 ( .A1(n1166), .A2(KEYINPUT32), .A3(n1107), .ZN(n1165) );
INV_X1 U837 ( .A(G475), .ZN(n1107) );
XNOR2_X1 U838 ( .A(G104), .B(n1167), .ZN(G6) );
NAND2_X1 U839 ( .A1(n1065), .A2(n1168), .ZN(n1167) );
INV_X1 U840 ( .A(n1042), .ZN(n1168) );
NAND2_X1 U841 ( .A1(n1058), .A2(n1169), .ZN(n1042) );
NOR2_X1 U842 ( .A1(n1155), .A2(n1170), .ZN(G57) );
XOR2_X1 U843 ( .A(n1171), .B(n1172), .Z(n1170) );
XNOR2_X1 U844 ( .A(n1173), .B(n1174), .ZN(n1172) );
NOR4_X1 U845 ( .A1(KEYINPUT49), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1173) );
NOR2_X1 U846 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XNOR2_X1 U847 ( .A(n1180), .B(n1181), .ZN(n1179) );
XOR2_X1 U848 ( .A(n1182), .B(n1183), .Z(n1171) );
AND2_X1 U849 ( .A1(G472), .A2(n1159), .ZN(n1183) );
NAND2_X1 U850 ( .A1(KEYINPUT44), .A2(G101), .ZN(n1182) );
NOR2_X1 U851 ( .A1(n1155), .A2(n1184), .ZN(G54) );
XOR2_X1 U852 ( .A(n1185), .B(n1186), .Z(n1184) );
XNOR2_X1 U853 ( .A(n1187), .B(n1178), .ZN(n1186) );
XOR2_X1 U854 ( .A(n1188), .B(n1189), .Z(n1185) );
XOR2_X1 U855 ( .A(n1190), .B(n1191), .Z(n1189) );
NAND2_X1 U856 ( .A1(KEYINPUT16), .A2(n1192), .ZN(n1191) );
NAND2_X1 U857 ( .A1(KEYINPUT11), .A2(n1193), .ZN(n1190) );
XNOR2_X1 U858 ( .A(KEYINPUT42), .B(n1194), .ZN(n1193) );
NAND2_X1 U859 ( .A1(n1159), .A2(G469), .ZN(n1188) );
NOR2_X1 U860 ( .A1(n1155), .A2(n1195), .ZN(G51) );
XOR2_X1 U861 ( .A(n1196), .B(n1197), .Z(n1195) );
NAND3_X1 U862 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1196) );
NAND2_X1 U863 ( .A1(KEYINPUT51), .A2(n1166), .ZN(n1199) );
INV_X1 U864 ( .A(n1159), .ZN(n1166) );
NOR2_X1 U865 ( .A1(n1201), .A2(n1047), .ZN(n1159) );
NAND2_X1 U866 ( .A1(n1202), .A2(n1203), .ZN(n1198) );
INV_X1 U867 ( .A(KEYINPUT51), .ZN(n1203) );
NAND2_X1 U868 ( .A1(n1047), .A2(G902), .ZN(n1202) );
AND3_X1 U869 ( .A1(n1119), .A2(n1204), .A3(n1139), .ZN(n1047) );
AND4_X1 U870 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1139) );
NAND3_X1 U871 ( .A1(n1209), .A2(n1210), .A3(KEYINPUT23), .ZN(n1208) );
AND2_X1 U872 ( .A1(n1211), .A2(n1212), .ZN(n1207) );
NAND2_X1 U873 ( .A1(n1169), .A2(n1213), .ZN(n1206) );
NAND3_X1 U874 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1213) );
NAND2_X1 U875 ( .A1(n1057), .A2(n1058), .ZN(n1216) );
NAND3_X1 U876 ( .A1(n1075), .A2(n1067), .A3(KEYINPUT60), .ZN(n1215) );
NAND2_X1 U877 ( .A1(n1065), .A2(n1217), .ZN(n1214) );
XNOR2_X1 U878 ( .A(KEYINPUT40), .B(n1062), .ZN(n1217) );
NAND2_X1 U879 ( .A1(n1218), .A2(n1219), .ZN(n1205) );
NAND2_X1 U880 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NAND2_X1 U881 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NAND2_X1 U882 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NAND4_X1 U883 ( .A1(n1075), .A2(n1067), .A3(n1082), .A4(n1226), .ZN(n1225) );
INV_X1 U884 ( .A(KEYINPUT60), .ZN(n1226) );
OR3_X1 U885 ( .A1(n1063), .A2(KEYINPUT23), .A3(n1227), .ZN(n1224) );
XOR2_X1 U886 ( .A(n1228), .B(KEYINPUT8), .Z(n1220) );
NAND4_X1 U887 ( .A1(n1229), .A2(n1230), .A3(n1067), .A4(n1231), .ZN(n1228) );
XNOR2_X1 U888 ( .A(n1056), .B(KEYINPUT46), .ZN(n1229) );
XNOR2_X1 U889 ( .A(KEYINPUT22), .B(n1138), .ZN(n1204) );
AND2_X1 U890 ( .A1(n1232), .A2(n1233), .ZN(n1119) );
AND4_X1 U891 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1233) );
NOR4_X1 U892 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1232) );
INV_X1 U893 ( .A(n1242), .ZN(n1241) );
NOR2_X1 U894 ( .A1(n1110), .A2(G952), .ZN(n1155) );
XOR2_X1 U895 ( .A(G146), .B(n1238), .Z(G48) );
AND3_X1 U896 ( .A1(n1065), .A2(n1218), .A3(n1243), .ZN(n1238) );
XNOR2_X1 U897 ( .A(G143), .B(n1242), .ZN(G45) );
NAND4_X1 U898 ( .A1(n1218), .A2(n1082), .A3(n1076), .A4(n1244), .ZN(n1242) );
AND3_X1 U899 ( .A1(n1098), .A2(n1245), .A3(n1246), .ZN(n1244) );
NAND2_X1 U900 ( .A1(n1247), .A2(n1248), .ZN(G42) );
NAND2_X1 U901 ( .A1(n1249), .A2(n1192), .ZN(n1248) );
XOR2_X1 U902 ( .A(n1237), .B(KEYINPUT4), .Z(n1249) );
NAND2_X1 U903 ( .A1(n1250), .A2(G140), .ZN(n1247) );
XNOR2_X1 U904 ( .A(KEYINPUT62), .B(n1237), .ZN(n1250) );
NAND3_X1 U905 ( .A1(n1065), .A2(n1075), .A3(n1251), .ZN(n1237) );
XNOR2_X1 U906 ( .A(G137), .B(n1236), .ZN(G39) );
NAND3_X1 U907 ( .A1(n1230), .A2(n1067), .A3(n1251), .ZN(n1236) );
XOR2_X1 U908 ( .A(G134), .B(n1240), .Z(G36) );
AND2_X1 U909 ( .A1(n1251), .A2(n1209), .ZN(n1240) );
XNOR2_X1 U910 ( .A(G131), .B(n1235), .ZN(G33) );
NAND3_X1 U911 ( .A1(n1065), .A2(n1076), .A3(n1251), .ZN(n1235) );
AND3_X1 U912 ( .A1(n1082), .A2(n1246), .A3(n1066), .ZN(n1251) );
NOR2_X1 U913 ( .A1(n1252), .A2(n1090), .ZN(n1066) );
XOR2_X1 U914 ( .A(n1253), .B(n1254), .Z(G30) );
NOR2_X1 U915 ( .A1(KEYINPUT21), .A2(n1255), .ZN(n1254) );
NAND2_X1 U916 ( .A1(n1256), .A2(n1257), .ZN(n1253) );
OR2_X1 U917 ( .A1(n1234), .A2(KEYINPUT18), .ZN(n1257) );
NAND3_X1 U918 ( .A1(n1057), .A2(n1218), .A3(n1243), .ZN(n1234) );
NAND3_X1 U919 ( .A1(n1218), .A2(n1258), .A3(KEYINPUT18), .ZN(n1256) );
NAND2_X1 U920 ( .A1(n1243), .A2(n1057), .ZN(n1258) );
AND3_X1 U921 ( .A1(n1082), .A2(n1246), .A3(n1230), .ZN(n1243) );
XNOR2_X1 U922 ( .A(G101), .B(n1212), .ZN(G3) );
NAND3_X1 U923 ( .A1(n1067), .A2(n1169), .A3(n1076), .ZN(n1212) );
XOR2_X1 U924 ( .A(G125), .B(n1239), .Z(G27) );
AND4_X1 U925 ( .A1(n1218), .A2(n1246), .A3(n1056), .A4(n1259), .ZN(n1239) );
AND2_X1 U926 ( .A1(n1075), .A2(n1065), .ZN(n1259) );
INV_X1 U927 ( .A(n1063), .ZN(n1056) );
NAND2_X1 U928 ( .A1(n1064), .A2(n1260), .ZN(n1246) );
NAND4_X1 U929 ( .A1(G953), .A2(n1261), .A3(n1262), .A4(n1114), .ZN(n1260) );
INV_X1 U930 ( .A(G900), .ZN(n1114) );
XNOR2_X1 U931 ( .A(KEYINPUT43), .B(n1263), .ZN(n1261) );
XNOR2_X1 U932 ( .A(G122), .B(n1211), .ZN(G24) );
NAND4_X1 U933 ( .A1(n1210), .A2(n1058), .A3(n1098), .A4(n1245), .ZN(n1211) );
INV_X1 U934 ( .A(n1062), .ZN(n1058) );
NAND2_X1 U935 ( .A1(n1264), .A2(n1094), .ZN(n1062) );
XNOR2_X1 U936 ( .A(n1265), .B(n1266), .ZN(G21) );
AND3_X1 U937 ( .A1(n1230), .A2(n1210), .A3(n1067), .ZN(n1266) );
NOR2_X1 U938 ( .A1(n1094), .A2(n1264), .ZN(n1230) );
INV_X1 U939 ( .A(n1267), .ZN(n1264) );
XOR2_X1 U940 ( .A(G116), .B(n1268), .Z(G18) );
AND2_X1 U941 ( .A1(n1210), .A2(n1209), .ZN(n1268) );
INV_X1 U942 ( .A(n1227), .ZN(n1209) );
NAND2_X1 U943 ( .A1(n1076), .A2(n1057), .ZN(n1227) );
INV_X1 U944 ( .A(n1041), .ZN(n1057) );
NAND2_X1 U945 ( .A1(n1269), .A2(n1098), .ZN(n1041) );
XNOR2_X1 U946 ( .A(G113), .B(n1138), .ZN(G15) );
NAND3_X1 U947 ( .A1(n1076), .A2(n1210), .A3(n1065), .ZN(n1138) );
NOR2_X1 U948 ( .A1(n1098), .A2(n1269), .ZN(n1065) );
NOR3_X1 U949 ( .A1(n1088), .A2(n1222), .A3(n1063), .ZN(n1210) );
NAND2_X1 U950 ( .A1(n1086), .A2(n1270), .ZN(n1063) );
INV_X1 U951 ( .A(n1231), .ZN(n1222) );
INV_X1 U952 ( .A(n1218), .ZN(n1088) );
NOR2_X1 U953 ( .A1(n1267), .A2(n1094), .ZN(n1076) );
XNOR2_X1 U954 ( .A(G110), .B(n1271), .ZN(G12) );
NAND3_X1 U955 ( .A1(n1067), .A2(n1169), .A3(n1075), .ZN(n1271) );
AND2_X1 U956 ( .A1(n1094), .A2(n1267), .ZN(n1075) );
NAND3_X1 U957 ( .A1(n1272), .A2(n1273), .A3(n1101), .ZN(n1267) );
NAND3_X1 U958 ( .A1(n1274), .A2(n1201), .A3(n1158), .ZN(n1101) );
NAND2_X1 U959 ( .A1(KEYINPUT24), .A2(n1274), .ZN(n1273) );
NAND2_X1 U960 ( .A1(n1102), .A2(n1275), .ZN(n1272) );
INV_X1 U961 ( .A(KEYINPUT24), .ZN(n1275) );
NOR2_X1 U962 ( .A1(n1274), .A2(n1276), .ZN(n1102) );
AND2_X1 U963 ( .A1(n1158), .A2(n1201), .ZN(n1276) );
XNOR2_X1 U964 ( .A(n1277), .B(n1278), .ZN(n1158) );
XNOR2_X1 U965 ( .A(n1279), .B(n1280), .ZN(n1278) );
XOR2_X1 U966 ( .A(n1281), .B(n1282), .Z(n1280) );
NAND2_X1 U967 ( .A1(KEYINPUT9), .A2(n1283), .ZN(n1281) );
XNOR2_X1 U968 ( .A(G137), .B(n1284), .ZN(n1283) );
NAND2_X1 U969 ( .A1(G221), .A2(n1285), .ZN(n1284) );
XOR2_X1 U970 ( .A(n1286), .B(n1287), .Z(n1277) );
NOR2_X1 U971 ( .A1(G125), .A2(KEYINPUT34), .ZN(n1287) );
XOR2_X1 U972 ( .A(n1288), .B(KEYINPUT19), .Z(n1286) );
NAND2_X1 U973 ( .A1(n1289), .A2(KEYINPUT58), .ZN(n1288) );
XNOR2_X1 U974 ( .A(G128), .B(n1290), .ZN(n1289) );
NOR2_X1 U975 ( .A1(G119), .A2(KEYINPUT7), .ZN(n1290) );
NAND2_X1 U976 ( .A1(G217), .A2(n1291), .ZN(n1274) );
XOR2_X1 U977 ( .A(KEYINPUT57), .B(n1292), .Z(n1291) );
NOR2_X1 U978 ( .A1(G902), .A2(n1293), .ZN(n1292) );
XOR2_X1 U979 ( .A(n1294), .B(G472), .Z(n1094) );
NAND3_X1 U980 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1294) );
XNOR2_X1 U981 ( .A(G902), .B(KEYINPUT0), .ZN(n1297) );
NAND2_X1 U982 ( .A1(KEYINPUT54), .A2(n1298), .ZN(n1296) );
XOR2_X1 U983 ( .A(n1299), .B(n1300), .Z(n1298) );
OR3_X1 U984 ( .A1(n1299), .A2(n1300), .A3(KEYINPUT54), .ZN(n1295) );
XNOR2_X1 U985 ( .A(n1174), .B(G101), .ZN(n1300) );
NAND2_X1 U986 ( .A1(G210), .A2(n1301), .ZN(n1174) );
NAND4_X1 U987 ( .A1(n1302), .A2(n1303), .A3(n1304), .A4(n1305), .ZN(n1299) );
NAND3_X1 U988 ( .A1(n1306), .A2(n1180), .A3(n1307), .ZN(n1305) );
XNOR2_X1 U989 ( .A(n1178), .B(KEYINPUT6), .ZN(n1306) );
INV_X1 U990 ( .A(n1308), .ZN(n1178) );
NAND3_X1 U991 ( .A1(n1308), .A2(n1309), .A3(n1181), .ZN(n1304) );
NAND2_X1 U992 ( .A1(n1180), .A2(n1310), .ZN(n1309) );
INV_X1 U993 ( .A(n1176), .ZN(n1303) );
NOR3_X1 U994 ( .A1(n1181), .A2(n1180), .A3(n1308), .ZN(n1176) );
INV_X1 U995 ( .A(n1311), .ZN(n1180) );
NAND2_X1 U996 ( .A1(n1175), .A2(n1310), .ZN(n1302) );
INV_X1 U997 ( .A(KEYINPUT6), .ZN(n1310) );
NOR3_X1 U998 ( .A1(n1308), .A2(n1307), .A3(n1311), .ZN(n1175) );
INV_X1 U999 ( .A(n1181), .ZN(n1307) );
XOR2_X1 U1000 ( .A(G119), .B(n1312), .Z(n1181) );
AND3_X1 U1001 ( .A1(n1082), .A2(n1231), .A3(n1218), .ZN(n1169) );
NOR2_X1 U1002 ( .A1(n1091), .A2(n1090), .ZN(n1218) );
AND2_X1 U1003 ( .A1(G214), .A2(n1313), .ZN(n1090) );
INV_X1 U1004 ( .A(n1252), .ZN(n1091) );
XNOR2_X1 U1005 ( .A(n1314), .B(n1200), .ZN(n1252) );
AND2_X1 U1006 ( .A1(G210), .A2(n1313), .ZN(n1200) );
NAND2_X1 U1007 ( .A1(n1315), .A2(n1201), .ZN(n1313) );
INV_X1 U1008 ( .A(G237), .ZN(n1315) );
NAND2_X1 U1009 ( .A1(n1316), .A2(n1201), .ZN(n1314) );
XNOR2_X1 U1010 ( .A(n1197), .B(n1317), .ZN(n1316) );
XOR2_X1 U1011 ( .A(KEYINPUT2), .B(KEYINPUT12), .Z(n1317) );
XNOR2_X1 U1012 ( .A(n1318), .B(n1319), .ZN(n1197) );
XNOR2_X1 U1013 ( .A(n1311), .B(n1320), .ZN(n1319) );
XOR2_X1 U1014 ( .A(n1321), .B(n1322), .Z(n1320) );
NOR2_X1 U1015 ( .A1(G953), .A2(n1131), .ZN(n1322) );
INV_X1 U1016 ( .A(G224), .ZN(n1131) );
NAND2_X1 U1017 ( .A1(KEYINPUT55), .A2(n1143), .ZN(n1321) );
XOR2_X1 U1018 ( .A(n1323), .B(n1282), .Z(n1143) );
XNOR2_X1 U1019 ( .A(G122), .B(KEYINPUT17), .ZN(n1323) );
XNOR2_X1 U1020 ( .A(n1324), .B(n1325), .ZN(n1311) );
XNOR2_X1 U1021 ( .A(G143), .B(KEYINPUT63), .ZN(n1324) );
XNOR2_X1 U1022 ( .A(n1148), .B(n1326), .ZN(n1318) );
XOR2_X1 U1023 ( .A(n1150), .B(n1152), .Z(n1148) );
XNOR2_X1 U1024 ( .A(n1039), .B(G101), .ZN(n1152) );
AND2_X1 U1025 ( .A1(n1327), .A2(n1328), .ZN(n1150) );
NAND2_X1 U1026 ( .A1(n1329), .A2(n1265), .ZN(n1328) );
INV_X1 U1027 ( .A(G119), .ZN(n1265) );
XOR2_X1 U1028 ( .A(KEYINPUT61), .B(n1312), .Z(n1329) );
NAND2_X1 U1029 ( .A1(n1312), .A2(G119), .ZN(n1327) );
XOR2_X1 U1030 ( .A(G113), .B(G116), .Z(n1312) );
NAND2_X1 U1031 ( .A1(n1064), .A2(n1330), .ZN(n1231) );
NAND3_X1 U1032 ( .A1(n1263), .A2(n1262), .A3(n1154), .ZN(n1330) );
NOR2_X1 U1033 ( .A1(G898), .A2(n1110), .ZN(n1154) );
XOR2_X1 U1034 ( .A(n1201), .B(KEYINPUT14), .Z(n1263) );
NAND3_X1 U1035 ( .A1(n1262), .A2(n1110), .A3(G952), .ZN(n1064) );
INV_X1 U1036 ( .A(G953), .ZN(n1110) );
NAND2_X1 U1037 ( .A1(G237), .A2(G234), .ZN(n1262) );
NOR2_X1 U1038 ( .A1(n1086), .A2(n1085), .ZN(n1082) );
INV_X1 U1039 ( .A(n1270), .ZN(n1085) );
NAND2_X1 U1040 ( .A1(G221), .A2(n1331), .ZN(n1270) );
NAND2_X1 U1041 ( .A1(G234), .A2(n1201), .ZN(n1331) );
XOR2_X1 U1042 ( .A(n1332), .B(G469), .Z(n1086) );
NAND2_X1 U1043 ( .A1(n1333), .A2(n1201), .ZN(n1332) );
XOR2_X1 U1044 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1045 ( .A(n1187), .B(n1336), .Z(n1335) );
XOR2_X1 U1046 ( .A(n1194), .B(n1337), .Z(n1336) );
NAND2_X1 U1047 ( .A1(KEYINPUT31), .A2(n1308), .ZN(n1337) );
NAND2_X1 U1048 ( .A1(n1338), .A2(n1339), .ZN(n1308) );
NAND2_X1 U1049 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
INV_X1 U1050 ( .A(G137), .ZN(n1341) );
XOR2_X1 U1051 ( .A(KEYINPUT36), .B(n1126), .Z(n1340) );
NAND2_X1 U1052 ( .A1(G137), .A2(n1342), .ZN(n1338) );
XNOR2_X1 U1053 ( .A(n1126), .B(KEYINPUT26), .ZN(n1342) );
XOR2_X1 U1054 ( .A(G131), .B(G134), .Z(n1126) );
NAND3_X1 U1055 ( .A1(n1343), .A2(n1344), .A3(n1345), .ZN(n1194) );
OR2_X1 U1056 ( .A1(n1346), .A2(KEYINPUT53), .ZN(n1345) );
OR3_X1 U1057 ( .A1(n1347), .A2(n1348), .A3(G101), .ZN(n1344) );
INV_X1 U1058 ( .A(KEYINPUT53), .ZN(n1347) );
NAND2_X1 U1059 ( .A1(G101), .A2(n1348), .ZN(n1343) );
NAND2_X1 U1060 ( .A1(KEYINPUT41), .A2(n1346), .ZN(n1348) );
XOR2_X1 U1061 ( .A(G107), .B(n1349), .Z(n1346) );
NOR2_X1 U1062 ( .A1(KEYINPUT33), .A2(n1147), .ZN(n1349) );
XOR2_X1 U1063 ( .A(n1350), .B(n1282), .Z(n1187) );
XOR2_X1 U1064 ( .A(G110), .B(KEYINPUT37), .Z(n1282) );
XOR2_X1 U1065 ( .A(n1125), .B(n1351), .Z(n1350) );
NOR2_X1 U1066 ( .A1(G953), .A2(n1113), .ZN(n1351) );
INV_X1 U1067 ( .A(G227), .ZN(n1113) );
XOR2_X1 U1068 ( .A(n1352), .B(n1325), .Z(n1125) );
XOR2_X1 U1069 ( .A(G146), .B(G128), .Z(n1325) );
NAND2_X1 U1070 ( .A1(KEYINPUT25), .A2(n1353), .ZN(n1352) );
XNOR2_X1 U1071 ( .A(n1354), .B(n1192), .ZN(n1334) );
XNOR2_X1 U1072 ( .A(KEYINPUT52), .B(KEYINPUT13), .ZN(n1354) );
NOR2_X1 U1073 ( .A1(n1098), .A2(n1245), .ZN(n1067) );
INV_X1 U1074 ( .A(n1269), .ZN(n1245) );
NOR2_X1 U1075 ( .A1(n1355), .A2(n1103), .ZN(n1269) );
NOR2_X1 U1076 ( .A1(n1105), .A2(G475), .ZN(n1103) );
AND2_X1 U1077 ( .A1(G475), .A2(n1105), .ZN(n1355) );
NAND2_X1 U1078 ( .A1(n1164), .A2(n1201), .ZN(n1105) );
XNOR2_X1 U1079 ( .A(n1356), .B(n1357), .ZN(n1164) );
XOR2_X1 U1080 ( .A(n1358), .B(n1359), .Z(n1357) );
XOR2_X1 U1081 ( .A(G131), .B(G113), .Z(n1359) );
XOR2_X1 U1082 ( .A(KEYINPUT47), .B(KEYINPUT27), .Z(n1358) );
XOR2_X1 U1083 ( .A(n1360), .B(n1361), .Z(n1356) );
XOR2_X1 U1084 ( .A(n1279), .B(n1362), .Z(n1361) );
XNOR2_X1 U1085 ( .A(G146), .B(n1192), .ZN(n1279) );
INV_X1 U1086 ( .A(G140), .ZN(n1192) );
XOR2_X1 U1087 ( .A(n1363), .B(n1326), .Z(n1360) );
XNOR2_X1 U1088 ( .A(n1147), .B(G125), .ZN(n1326) );
INV_X1 U1089 ( .A(G104), .ZN(n1147) );
NAND2_X1 U1090 ( .A1(G214), .A2(n1301), .ZN(n1363) );
NOR2_X1 U1091 ( .A1(G953), .A2(G237), .ZN(n1301) );
XNOR2_X1 U1092 ( .A(n1364), .B(G478), .ZN(n1098) );
NAND2_X1 U1093 ( .A1(n1162), .A2(n1201), .ZN(n1364) );
INV_X1 U1094 ( .A(G902), .ZN(n1201) );
XNOR2_X1 U1095 ( .A(n1365), .B(n1366), .ZN(n1162) );
XOR2_X1 U1096 ( .A(n1362), .B(n1367), .Z(n1366) );
XNOR2_X1 U1097 ( .A(n1039), .B(n1368), .ZN(n1367) );
AND3_X1 U1098 ( .A1(G217), .A2(n1369), .A3(n1285), .ZN(n1368) );
NOR2_X1 U1099 ( .A1(n1293), .A2(G953), .ZN(n1285) );
INV_X1 U1100 ( .A(G234), .ZN(n1293) );
INV_X1 U1101 ( .A(KEYINPUT29), .ZN(n1369) );
INV_X1 U1102 ( .A(G107), .ZN(n1039) );
XNOR2_X1 U1103 ( .A(G122), .B(n1353), .ZN(n1362) );
INV_X1 U1104 ( .A(G143), .ZN(n1353) );
XNOR2_X1 U1105 ( .A(G116), .B(n1370), .ZN(n1365) );
XNOR2_X1 U1106 ( .A(G134), .B(n1255), .ZN(n1370) );
INV_X1 U1107 ( .A(G128), .ZN(n1255) );
endmodule


