//Key = 0011101010000010010010110100011000010011110000011111111000001010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408;

XOR2_X1 U774 ( .A(n1073), .B(n1074), .Z(G9) );
NOR3_X1 U775 ( .A1(n1075), .A2(KEYINPUT7), .A3(n1076), .ZN(n1074) );
XNOR2_X1 U776 ( .A(G107), .B(KEYINPUT23), .ZN(n1073) );
NOR2_X1 U777 ( .A1(n1077), .A2(n1078), .ZN(G75) );
NOR2_X1 U778 ( .A1(G952), .A2(n1079), .ZN(n1078) );
NOR4_X1 U779 ( .A1(n1080), .A2(n1081), .A3(KEYINPUT19), .A4(n1082), .ZN(n1077) );
NOR2_X1 U780 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
INV_X1 U781 ( .A(n1085), .ZN(n1084) );
NOR2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(n1083) );
NOR2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR2_X1 U784 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
XNOR2_X1 U785 ( .A(n1092), .B(KEYINPUT51), .ZN(n1091) );
NOR2_X1 U786 ( .A1(KEYINPUT63), .A2(n1093), .ZN(n1090) );
NOR2_X1 U787 ( .A1(n1094), .A2(n1095), .ZN(n1086) );
NOR2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NOR2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
NOR4_X1 U790 ( .A1(n1100), .A2(n1101), .A3(n1095), .A4(n1089), .ZN(n1081) );
INV_X1 U791 ( .A(n1102), .ZN(n1095) );
NOR2_X1 U792 ( .A1(n1103), .A2(n1104), .ZN(n1100) );
NOR2_X1 U793 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NOR2_X1 U794 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
NOR2_X1 U795 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
NOR2_X1 U796 ( .A1(n1111), .A2(n1112), .ZN(n1103) );
NOR2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NAND3_X1 U799 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1080) );
NAND2_X1 U800 ( .A1(KEYINPUT63), .A2(n1120), .ZN(n1118) );
NAND3_X1 U801 ( .A1(n1121), .A2(n1122), .A3(n1085), .ZN(n1120) );
NOR3_X1 U802 ( .A1(n1112), .A2(n1106), .A3(n1101), .ZN(n1085) );
INV_X1 U803 ( .A(n1123), .ZN(n1106) );
INV_X1 U804 ( .A(n1079), .ZN(n1117) );
NAND2_X1 U805 ( .A1(n1124), .A2(n1125), .ZN(n1079) );
NAND4_X1 U806 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n1125) );
NOR4_X1 U807 ( .A1(n1130), .A2(n1131), .A3(n1112), .A4(n1132), .ZN(n1129) );
XNOR2_X1 U808 ( .A(n1133), .B(n1134), .ZN(n1132) );
XNOR2_X1 U809 ( .A(n1135), .B(n1136), .ZN(n1131) );
NAND2_X1 U810 ( .A1(KEYINPUT3), .A2(n1137), .ZN(n1135) );
XNOR2_X1 U811 ( .A(n1138), .B(n1139), .ZN(n1128) );
XOR2_X1 U812 ( .A(n1140), .B(n1141), .Z(n1127) );
XNOR2_X1 U813 ( .A(n1098), .B(KEYINPUT36), .ZN(n1126) );
XOR2_X1 U814 ( .A(n1142), .B(n1143), .Z(G72) );
NOR2_X1 U815 ( .A1(n1144), .A2(n1124), .ZN(n1143) );
NOR2_X1 U816 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U817 ( .A(KEYINPUT47), .B(G227), .Z(n1146) );
NAND2_X1 U818 ( .A1(n1147), .A2(n1148), .ZN(n1142) );
NAND2_X1 U819 ( .A1(n1149), .A2(n1124), .ZN(n1148) );
XOR2_X1 U820 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U821 ( .A(n1152), .B(KEYINPUT34), .Z(n1150) );
NAND3_X1 U822 ( .A1(n1151), .A2(G900), .A3(G953), .ZN(n1147) );
NOR2_X1 U823 ( .A1(KEYINPUT26), .A2(n1153), .ZN(n1151) );
XOR2_X1 U824 ( .A(n1154), .B(n1155), .Z(n1153) );
XNOR2_X1 U825 ( .A(n1156), .B(n1157), .ZN(n1155) );
XOR2_X1 U826 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U827 ( .A1(G137), .A2(KEYINPUT59), .ZN(n1159) );
NOR2_X1 U828 ( .A1(G125), .A2(KEYINPUT18), .ZN(n1158) );
XNOR2_X1 U829 ( .A(n1160), .B(n1161), .ZN(n1154) );
XOR2_X1 U830 ( .A(G140), .B(G134), .Z(n1161) );
XOR2_X1 U831 ( .A(n1162), .B(n1163), .Z(G69) );
XOR2_X1 U832 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U833 ( .A1(n1166), .A2(KEYINPUT61), .ZN(n1165) );
AND2_X1 U834 ( .A1(n1124), .A2(n1167), .ZN(n1166) );
NOR2_X1 U835 ( .A1(n1168), .A2(n1169), .ZN(n1164) );
XOR2_X1 U836 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U837 ( .A1(KEYINPUT22), .A2(n1172), .ZN(n1170) );
NOR2_X1 U838 ( .A1(G898), .A2(n1124), .ZN(n1168) );
NAND2_X1 U839 ( .A1(G953), .A2(n1173), .ZN(n1162) );
NAND2_X1 U840 ( .A1(G898), .A2(G224), .ZN(n1173) );
NOR2_X1 U841 ( .A1(n1174), .A2(n1175), .ZN(G66) );
NOR3_X1 U842 ( .A1(n1140), .A2(n1176), .A3(n1177), .ZN(n1175) );
NOR3_X1 U843 ( .A1(n1178), .A2(n1141), .A3(n1179), .ZN(n1177) );
NOR2_X1 U844 ( .A1(n1180), .A2(n1181), .ZN(n1176) );
NOR2_X1 U845 ( .A1(n1119), .A2(n1141), .ZN(n1180) );
NOR2_X1 U846 ( .A1(n1174), .A2(n1182), .ZN(G63) );
XOR2_X1 U847 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U848 ( .A1(n1139), .A2(n1179), .ZN(n1184) );
NAND2_X1 U849 ( .A1(KEYINPUT4), .A2(n1185), .ZN(n1183) );
NOR2_X1 U850 ( .A1(n1174), .A2(n1186), .ZN(G60) );
NOR3_X1 U851 ( .A1(n1134), .A2(n1187), .A3(n1188), .ZN(n1186) );
NOR2_X1 U852 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NOR3_X1 U853 ( .A1(n1133), .A2(KEYINPUT45), .A3(n1119), .ZN(n1189) );
NOR4_X1 U854 ( .A1(n1191), .A2(n1179), .A3(KEYINPUT45), .A4(n1133), .ZN(n1187) );
INV_X1 U855 ( .A(n1192), .ZN(n1179) );
INV_X1 U856 ( .A(n1190), .ZN(n1191) );
XNOR2_X1 U857 ( .A(n1193), .B(n1194), .ZN(G6) );
NOR3_X1 U858 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(G57) );
NOR2_X1 U859 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NOR2_X1 U860 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
AND2_X1 U861 ( .A1(KEYINPUT10), .A2(n1202), .ZN(n1201) );
NOR3_X1 U862 ( .A1(KEYINPUT10), .A2(n1202), .A3(n1203), .ZN(n1200) );
NOR2_X1 U863 ( .A1(n1204), .A2(n1205), .ZN(n1196) );
INV_X1 U864 ( .A(n1198), .ZN(n1205) );
XNOR2_X1 U865 ( .A(n1206), .B(n1207), .ZN(n1198) );
XOR2_X1 U866 ( .A(n1208), .B(n1209), .Z(n1206) );
NOR2_X1 U867 ( .A1(KEYINPUT43), .A2(n1210), .ZN(n1209) );
XNOR2_X1 U868 ( .A(n1211), .B(n1212), .ZN(n1210) );
NOR2_X1 U869 ( .A1(KEYINPUT46), .A2(n1213), .ZN(n1212) );
NAND2_X1 U870 ( .A1(n1192), .A2(G472), .ZN(n1208) );
NOR2_X1 U871 ( .A1(n1202), .A2(n1203), .ZN(n1204) );
INV_X1 U872 ( .A(KEYINPUT20), .ZN(n1203) );
XOR2_X1 U873 ( .A(n1214), .B(n1215), .Z(n1202) );
XOR2_X1 U874 ( .A(KEYINPUT44), .B(n1174), .Z(n1195) );
NOR2_X1 U875 ( .A1(n1174), .A2(n1216), .ZN(G54) );
XOR2_X1 U876 ( .A(n1217), .B(n1218), .Z(n1216) );
XNOR2_X1 U877 ( .A(n1211), .B(n1219), .ZN(n1218) );
NAND2_X1 U878 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NAND2_X1 U879 ( .A1(G110), .A2(n1222), .ZN(n1221) );
NAND2_X1 U880 ( .A1(n1223), .A2(n1224), .ZN(n1220) );
XNOR2_X1 U881 ( .A(KEYINPUT21), .B(n1222), .ZN(n1223) );
XOR2_X1 U882 ( .A(n1225), .B(n1226), .Z(n1217) );
NAND2_X1 U883 ( .A1(n1192), .A2(G469), .ZN(n1226) );
NAND2_X1 U884 ( .A1(KEYINPUT25), .A2(n1227), .ZN(n1225) );
XOR2_X1 U885 ( .A(n1228), .B(n1229), .Z(n1227) );
NOR2_X1 U886 ( .A1(KEYINPUT12), .A2(n1156), .ZN(n1228) );
NOR2_X1 U887 ( .A1(n1174), .A2(n1230), .ZN(G51) );
NOR2_X1 U888 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XOR2_X1 U889 ( .A(n1233), .B(KEYINPUT17), .Z(n1232) );
NAND2_X1 U890 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NOR2_X1 U891 ( .A1(n1234), .A2(n1235), .ZN(n1231) );
XOR2_X1 U892 ( .A(n1236), .B(n1237), .Z(n1235) );
XNOR2_X1 U893 ( .A(n1238), .B(n1239), .ZN(n1237) );
NOR3_X1 U894 ( .A1(n1240), .A2(KEYINPUT33), .A3(G953), .ZN(n1239) );
NAND2_X1 U895 ( .A1(KEYINPUT41), .A2(n1241), .ZN(n1238) );
XNOR2_X1 U896 ( .A(n1242), .B(n1213), .ZN(n1236) );
AND2_X1 U897 ( .A1(n1192), .A2(n1243), .ZN(n1234) );
NOR2_X1 U898 ( .A1(n1244), .A2(n1119), .ZN(n1192) );
NOR2_X1 U899 ( .A1(n1167), .A2(n1152), .ZN(n1119) );
NAND2_X1 U900 ( .A1(n1245), .A2(n1246), .ZN(n1152) );
NOR4_X1 U901 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1246) );
AND4_X1 U902 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1245) );
NAND4_X1 U903 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1167) );
AND4_X1 U904 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1258) );
INV_X1 U905 ( .A(n1263), .ZN(n1260) );
NAND2_X1 U906 ( .A1(n1092), .A2(n1264), .ZN(n1257) );
NAND2_X1 U907 ( .A1(n1265), .A2(n1076), .ZN(n1264) );
INV_X1 U908 ( .A(n1194), .ZN(n1255) );
NOR2_X1 U909 ( .A1(n1093), .A2(n1076), .ZN(n1194) );
NAND2_X1 U910 ( .A1(n1266), .A2(n1123), .ZN(n1076) );
NOR2_X1 U911 ( .A1(n1124), .A2(G952), .ZN(n1174) );
XNOR2_X1 U912 ( .A(G146), .B(n1254), .ZN(G48) );
NAND3_X1 U913 ( .A1(n1122), .A2(n1108), .A3(n1267), .ZN(n1254) );
XNOR2_X1 U914 ( .A(G143), .B(n1253), .ZN(G45) );
NAND4_X1 U915 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1253) );
AND3_X1 U916 ( .A1(n1114), .A2(n1108), .A3(n1097), .ZN(n1271) );
NAND2_X1 U917 ( .A1(n1272), .A2(n1273), .ZN(G42) );
OR2_X1 U918 ( .A1(n1252), .A2(G140), .ZN(n1273) );
XOR2_X1 U919 ( .A(n1274), .B(KEYINPUT58), .Z(n1272) );
NAND2_X1 U920 ( .A1(G140), .A2(n1252), .ZN(n1274) );
NAND3_X1 U921 ( .A1(n1275), .A2(n1097), .A3(n1276), .ZN(n1252) );
XNOR2_X1 U922 ( .A(G137), .B(n1251), .ZN(G39) );
NAND3_X1 U923 ( .A1(n1102), .A2(n1275), .A3(n1267), .ZN(n1251) );
XOR2_X1 U924 ( .A(n1249), .B(n1277), .Z(G36) );
XOR2_X1 U925 ( .A(KEYINPUT11), .B(G134), .Z(n1277) );
AND2_X1 U926 ( .A1(n1278), .A2(n1092), .ZN(n1249) );
XOR2_X1 U927 ( .A(n1248), .B(n1279), .Z(G33) );
NOR2_X1 U928 ( .A1(KEYINPUT27), .A2(n1160), .ZN(n1279) );
AND2_X1 U929 ( .A1(n1278), .A2(n1122), .ZN(n1248) );
AND4_X1 U930 ( .A1(n1114), .A2(n1275), .A3(n1097), .A4(n1268), .ZN(n1278) );
INV_X1 U931 ( .A(n1112), .ZN(n1275) );
NAND2_X1 U932 ( .A1(n1280), .A2(n1110), .ZN(n1112) );
INV_X1 U933 ( .A(n1109), .ZN(n1280) );
NAND3_X1 U934 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(G30) );
OR2_X1 U935 ( .A1(G128), .A2(KEYINPUT14), .ZN(n1283) );
NAND3_X1 U936 ( .A1(KEYINPUT14), .A2(G128), .A3(n1284), .ZN(n1282) );
NAND2_X1 U937 ( .A1(n1250), .A2(n1285), .ZN(n1281) );
NAND2_X1 U938 ( .A1(n1286), .A2(KEYINPUT14), .ZN(n1285) );
XNOR2_X1 U939 ( .A(G128), .B(KEYINPUT60), .ZN(n1286) );
INV_X1 U940 ( .A(n1284), .ZN(n1250) );
NAND3_X1 U941 ( .A1(n1092), .A2(n1108), .A3(n1267), .ZN(n1284) );
AND4_X1 U942 ( .A1(n1287), .A2(n1097), .A3(n1115), .A4(n1268), .ZN(n1267) );
INV_X1 U943 ( .A(n1075), .ZN(n1092) );
XNOR2_X1 U944 ( .A(G101), .B(n1256), .ZN(G3) );
NAND3_X1 U945 ( .A1(n1102), .A2(n1266), .A3(n1114), .ZN(n1256) );
XOR2_X1 U946 ( .A(n1288), .B(n1289), .Z(G27) );
XNOR2_X1 U947 ( .A(G125), .B(KEYINPUT42), .ZN(n1289) );
NAND2_X1 U948 ( .A1(KEYINPUT8), .A2(n1247), .ZN(n1288) );
AND3_X1 U949 ( .A1(n1121), .A2(n1108), .A3(n1276), .ZN(n1247) );
AND4_X1 U950 ( .A1(n1287), .A2(n1122), .A3(n1290), .A4(n1268), .ZN(n1276) );
NAND2_X1 U951 ( .A1(n1101), .A2(n1291), .ZN(n1268) );
NAND4_X1 U952 ( .A1(G953), .A2(G902), .A3(n1292), .A4(n1145), .ZN(n1291) );
INV_X1 U953 ( .A(G900), .ZN(n1145) );
XNOR2_X1 U954 ( .A(G122), .B(n1262), .ZN(G24) );
NAND4_X1 U955 ( .A1(n1293), .A2(n1123), .A3(n1270), .A4(n1269), .ZN(n1262) );
NOR2_X1 U956 ( .A1(n1115), .A2(n1287), .ZN(n1123) );
XNOR2_X1 U957 ( .A(G119), .B(n1261), .ZN(G21) );
NAND4_X1 U958 ( .A1(n1293), .A2(n1287), .A3(n1102), .A4(n1115), .ZN(n1261) );
NAND2_X1 U959 ( .A1(n1294), .A2(n1295), .ZN(G18) );
OR2_X1 U960 ( .A1(n1296), .A2(G116), .ZN(n1295) );
NAND2_X1 U961 ( .A1(G116), .A2(n1297), .ZN(n1294) );
NAND2_X1 U962 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NAND2_X1 U963 ( .A1(KEYINPUT32), .A2(n1300), .ZN(n1299) );
NAND2_X1 U964 ( .A1(n1296), .A2(n1301), .ZN(n1298) );
INV_X1 U965 ( .A(KEYINPUT32), .ZN(n1301) );
NAND2_X1 U966 ( .A1(KEYINPUT53), .A2(n1300), .ZN(n1296) );
AND4_X1 U967 ( .A1(n1302), .A2(n1114), .A3(n1303), .A4(n1121), .ZN(n1300) );
NOR2_X1 U968 ( .A1(n1304), .A2(n1075), .ZN(n1303) );
NAND2_X1 U969 ( .A1(n1305), .A2(n1269), .ZN(n1075) );
XNOR2_X1 U970 ( .A(n1108), .B(KEYINPUT6), .ZN(n1302) );
INV_X1 U971 ( .A(n1306), .ZN(n1108) );
XNOR2_X1 U972 ( .A(n1307), .B(n1263), .ZN(G15) );
NOR2_X1 U973 ( .A1(n1265), .A2(n1093), .ZN(n1263) );
INV_X1 U974 ( .A(n1122), .ZN(n1093) );
NOR2_X1 U975 ( .A1(n1269), .A2(n1305), .ZN(n1122) );
INV_X1 U976 ( .A(n1270), .ZN(n1305) );
NAND2_X1 U977 ( .A1(n1293), .A2(n1114), .ZN(n1265) );
NOR2_X1 U978 ( .A1(n1290), .A2(n1287), .ZN(n1114) );
NOR3_X1 U979 ( .A1(n1306), .A2(n1304), .A3(n1089), .ZN(n1293) );
INV_X1 U980 ( .A(n1121), .ZN(n1089) );
NOR2_X1 U981 ( .A1(n1098), .A2(n1130), .ZN(n1121) );
XOR2_X1 U982 ( .A(n1259), .B(n1308), .Z(G12) );
XNOR2_X1 U983 ( .A(G110), .B(KEYINPUT13), .ZN(n1308) );
NAND4_X1 U984 ( .A1(n1287), .A2(n1102), .A3(n1290), .A4(n1266), .ZN(n1259) );
NOR3_X1 U985 ( .A1(n1306), .A2(n1304), .A3(n1309), .ZN(n1266) );
INV_X1 U986 ( .A(n1097), .ZN(n1309) );
NOR2_X1 U987 ( .A1(n1310), .A2(n1130), .ZN(n1097) );
INV_X1 U988 ( .A(n1099), .ZN(n1130) );
NAND2_X1 U989 ( .A1(G221), .A2(n1311), .ZN(n1099) );
INV_X1 U990 ( .A(n1098), .ZN(n1310) );
XNOR2_X1 U991 ( .A(n1312), .B(G469), .ZN(n1098) );
NAND4_X1 U992 ( .A1(n1313), .A2(n1244), .A3(n1314), .A4(n1315), .ZN(n1312) );
NAND3_X1 U993 ( .A1(KEYINPUT48), .A2(n1316), .A3(n1317), .ZN(n1315) );
OR2_X1 U994 ( .A1(n1317), .A2(n1316), .ZN(n1314) );
AND2_X1 U995 ( .A1(KEYINPUT62), .A2(n1318), .ZN(n1316) );
XOR2_X1 U996 ( .A(n1319), .B(n1320), .Z(n1317) );
XNOR2_X1 U997 ( .A(KEYINPUT50), .B(n1321), .ZN(n1319) );
NOR2_X1 U998 ( .A1(KEYINPUT57), .A2(n1322), .ZN(n1321) );
XNOR2_X1 U999 ( .A(n1156), .B(n1229), .ZN(n1322) );
XNOR2_X1 U1000 ( .A(n1323), .B(n1324), .ZN(n1229) );
NAND2_X1 U1001 ( .A1(KEYINPUT2), .A2(n1215), .ZN(n1323) );
OR2_X1 U1002 ( .A1(n1318), .A2(KEYINPUT48), .ZN(n1313) );
XNOR2_X1 U1003 ( .A(G110), .B(n1222), .ZN(n1318) );
XNOR2_X1 U1004 ( .A(G140), .B(n1325), .ZN(n1222) );
AND2_X1 U1005 ( .A1(n1124), .A2(G227), .ZN(n1325) );
AND2_X1 U1006 ( .A1(n1326), .A2(n1101), .ZN(n1304) );
NAND3_X1 U1007 ( .A1(n1292), .A2(n1124), .A3(G952), .ZN(n1101) );
NAND4_X1 U1008 ( .A1(G953), .A2(G902), .A3(n1292), .A4(n1327), .ZN(n1326) );
INV_X1 U1009 ( .A(G898), .ZN(n1327) );
NAND2_X1 U1010 ( .A1(G237), .A2(G234), .ZN(n1292) );
NAND2_X1 U1011 ( .A1(n1109), .A2(n1110), .ZN(n1306) );
NAND2_X1 U1012 ( .A1(G214), .A2(n1328), .ZN(n1110) );
XNOR2_X1 U1013 ( .A(n1329), .B(n1243), .ZN(n1109) );
AND2_X1 U1014 ( .A1(G210), .A2(n1328), .ZN(n1243) );
NAND2_X1 U1015 ( .A1(n1330), .A2(n1244), .ZN(n1328) );
INV_X1 U1016 ( .A(G237), .ZN(n1330) );
NAND2_X1 U1017 ( .A1(n1331), .A2(n1244), .ZN(n1329) );
XNOR2_X1 U1018 ( .A(n1332), .B(n1333), .ZN(n1331) );
INV_X1 U1019 ( .A(n1242), .ZN(n1333) );
XOR2_X1 U1020 ( .A(n1172), .B(n1171), .Z(n1242) );
XNOR2_X1 U1021 ( .A(n1334), .B(n1335), .ZN(n1171) );
XNOR2_X1 U1022 ( .A(G122), .B(n1224), .ZN(n1335) );
XNOR2_X1 U1023 ( .A(G101), .B(n1324), .ZN(n1334) );
XNOR2_X1 U1024 ( .A(n1193), .B(G107), .ZN(n1324) );
AND2_X1 U1025 ( .A1(n1336), .A2(n1337), .ZN(n1172) );
NAND2_X1 U1026 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
INV_X1 U1027 ( .A(G119), .ZN(n1339) );
NAND2_X1 U1028 ( .A1(n1340), .A2(G119), .ZN(n1336) );
XOR2_X1 U1029 ( .A(KEYINPUT39), .B(n1338), .Z(n1340) );
NOR2_X1 U1030 ( .A1(KEYINPUT56), .A2(n1341), .ZN(n1332) );
XNOR2_X1 U1031 ( .A(n1156), .B(n1342), .ZN(n1341) );
XNOR2_X1 U1032 ( .A(n1240), .B(G125), .ZN(n1342) );
INV_X1 U1033 ( .A(G224), .ZN(n1240) );
INV_X1 U1034 ( .A(n1213), .ZN(n1156) );
INV_X1 U1035 ( .A(n1115), .ZN(n1290) );
XOR2_X1 U1036 ( .A(n1136), .B(n1137), .Z(n1115) );
INV_X1 U1037 ( .A(G472), .ZN(n1137) );
NAND2_X1 U1038 ( .A1(n1343), .A2(n1244), .ZN(n1136) );
XOR2_X1 U1039 ( .A(n1344), .B(n1345), .Z(n1343) );
XNOR2_X1 U1040 ( .A(n1207), .B(n1320), .ZN(n1345) );
INV_X1 U1041 ( .A(n1211), .ZN(n1320) );
XNOR2_X1 U1042 ( .A(n1346), .B(n1347), .ZN(n1211) );
XOR2_X1 U1043 ( .A(G137), .B(G134), .Z(n1347) );
NAND2_X1 U1044 ( .A1(KEYINPUT38), .A2(n1160), .ZN(n1346) );
XNOR2_X1 U1045 ( .A(n1348), .B(n1338), .ZN(n1207) );
XNOR2_X1 U1046 ( .A(n1307), .B(G116), .ZN(n1338) );
XNOR2_X1 U1047 ( .A(G119), .B(KEYINPUT16), .ZN(n1348) );
XNOR2_X1 U1048 ( .A(n1349), .B(n1213), .ZN(n1344) );
XOR2_X1 U1049 ( .A(G146), .B(n1350), .Z(n1213) );
NAND3_X1 U1050 ( .A1(n1351), .A2(n1352), .A3(n1353), .ZN(n1349) );
NAND2_X1 U1051 ( .A1(n1214), .A2(n1354), .ZN(n1353) );
INV_X1 U1052 ( .A(KEYINPUT49), .ZN(n1354) );
NAND3_X1 U1053 ( .A1(KEYINPUT49), .A2(n1355), .A3(n1215), .ZN(n1352) );
OR2_X1 U1054 ( .A1(n1215), .A2(n1355), .ZN(n1351) );
NOR2_X1 U1055 ( .A1(n1356), .A2(n1214), .ZN(n1355) );
NAND2_X1 U1056 ( .A1(G210), .A2(n1357), .ZN(n1214) );
INV_X1 U1057 ( .A(KEYINPUT54), .ZN(n1356) );
INV_X1 U1058 ( .A(G101), .ZN(n1215) );
NOR2_X1 U1059 ( .A1(n1269), .A2(n1270), .ZN(n1102) );
XNOR2_X1 U1060 ( .A(n1358), .B(n1359), .ZN(n1270) );
NOR2_X1 U1061 ( .A1(KEYINPUT24), .A2(n1133), .ZN(n1359) );
INV_X1 U1062 ( .A(G475), .ZN(n1133) );
XNOR2_X1 U1063 ( .A(n1134), .B(KEYINPUT28), .ZN(n1358) );
NOR2_X1 U1064 ( .A1(n1190), .A2(G902), .ZN(n1134) );
XNOR2_X1 U1065 ( .A(n1360), .B(n1361), .ZN(n1190) );
XOR2_X1 U1066 ( .A(n1362), .B(n1363), .Z(n1361) );
XOR2_X1 U1067 ( .A(n1364), .B(n1365), .Z(n1363) );
NOR2_X1 U1068 ( .A1(n1366), .A2(n1367), .ZN(n1365) );
AND2_X1 U1069 ( .A1(KEYINPUT0), .A2(n1307), .ZN(n1367) );
NOR2_X1 U1070 ( .A1(KEYINPUT1), .A2(n1307), .ZN(n1366) );
INV_X1 U1071 ( .A(G113), .ZN(n1307) );
NAND2_X1 U1072 ( .A1(KEYINPUT40), .A2(n1193), .ZN(n1364) );
INV_X1 U1073 ( .A(G104), .ZN(n1193) );
XOR2_X1 U1074 ( .A(n1368), .B(n1369), .Z(n1362) );
NOR4_X1 U1075 ( .A1(n1370), .A2(n1371), .A3(KEYINPUT31), .A4(n1372), .ZN(n1369) );
NOR2_X1 U1076 ( .A1(G125), .A2(n1373), .ZN(n1372) );
NOR2_X1 U1077 ( .A1(KEYINPUT9), .A2(n1374), .ZN(n1373) );
XOR2_X1 U1078 ( .A(KEYINPUT52), .B(n1375), .Z(n1374) );
NOR2_X1 U1079 ( .A1(n1375), .A2(n1376), .ZN(n1371) );
AND3_X1 U1080 ( .A1(n1376), .A2(n1375), .A3(G125), .ZN(n1370) );
INV_X1 U1081 ( .A(KEYINPUT9), .ZN(n1376) );
NAND2_X1 U1082 ( .A1(G214), .A2(n1357), .ZN(n1368) );
NOR2_X1 U1083 ( .A1(G953), .A2(G237), .ZN(n1357) );
XOR2_X1 U1084 ( .A(n1377), .B(n1378), .Z(n1360) );
XNOR2_X1 U1085 ( .A(n1160), .B(G122), .ZN(n1378) );
INV_X1 U1086 ( .A(G131), .ZN(n1160) );
XNOR2_X1 U1087 ( .A(G143), .B(G146), .ZN(n1377) );
NAND3_X1 U1088 ( .A1(n1379), .A2(n1380), .A3(n1381), .ZN(n1269) );
OR2_X1 U1089 ( .A1(n1382), .A2(n1138), .ZN(n1381) );
NAND3_X1 U1090 ( .A1(n1138), .A2(n1382), .A3(G478), .ZN(n1380) );
NAND2_X1 U1091 ( .A1(n1383), .A2(n1139), .ZN(n1379) );
INV_X1 U1092 ( .A(G478), .ZN(n1139) );
NAND2_X1 U1093 ( .A1(n1384), .A2(n1382), .ZN(n1383) );
INV_X1 U1094 ( .A(KEYINPUT5), .ZN(n1382) );
XNOR2_X1 U1095 ( .A(KEYINPUT35), .B(n1138), .ZN(n1384) );
NAND2_X1 U1096 ( .A1(n1185), .A2(n1244), .ZN(n1138) );
XNOR2_X1 U1097 ( .A(n1385), .B(n1386), .ZN(n1185) );
XOR2_X1 U1098 ( .A(n1350), .B(n1387), .Z(n1386) );
XOR2_X1 U1099 ( .A(G107), .B(n1388), .Z(n1387) );
AND3_X1 U1100 ( .A1(G234), .A2(n1124), .A3(G217), .ZN(n1388) );
XNOR2_X1 U1101 ( .A(n1389), .B(G128), .ZN(n1350) );
INV_X1 U1102 ( .A(G143), .ZN(n1389) );
XNOR2_X1 U1103 ( .A(G116), .B(n1390), .ZN(n1385) );
XOR2_X1 U1104 ( .A(G134), .B(G122), .Z(n1390) );
INV_X1 U1105 ( .A(n1116), .ZN(n1287) );
NAND2_X1 U1106 ( .A1(n1391), .A2(n1392), .ZN(n1116) );
NAND2_X1 U1107 ( .A1(n1393), .A2(n1394), .ZN(n1392) );
NAND2_X1 U1108 ( .A1(n1395), .A2(n1396), .ZN(n1394) );
OR2_X1 U1109 ( .A1(n1140), .A2(KEYINPUT55), .ZN(n1396) );
INV_X1 U1110 ( .A(KEYINPUT15), .ZN(n1395) );
NAND2_X1 U1111 ( .A1(n1140), .A2(n1397), .ZN(n1391) );
NAND2_X1 U1112 ( .A1(n1398), .A2(n1399), .ZN(n1397) );
OR2_X1 U1113 ( .A1(n1393), .A2(KEYINPUT15), .ZN(n1399) );
XOR2_X1 U1114 ( .A(n1141), .B(KEYINPUT37), .Z(n1393) );
NAND2_X1 U1115 ( .A1(G217), .A2(n1311), .ZN(n1141) );
NAND2_X1 U1116 ( .A1(G234), .A2(n1244), .ZN(n1311) );
INV_X1 U1117 ( .A(G902), .ZN(n1244) );
INV_X1 U1118 ( .A(KEYINPUT55), .ZN(n1398) );
NOR2_X1 U1119 ( .A1(n1181), .A2(G902), .ZN(n1140) );
INV_X1 U1120 ( .A(n1178), .ZN(n1181) );
XOR2_X1 U1121 ( .A(n1400), .B(n1401), .Z(n1178) );
XOR2_X1 U1122 ( .A(n1402), .B(n1403), .Z(n1401) );
XNOR2_X1 U1123 ( .A(n1404), .B(n1224), .ZN(n1403) );
INV_X1 U1124 ( .A(G110), .ZN(n1224) );
NAND3_X1 U1125 ( .A1(G234), .A2(n1124), .A3(G221), .ZN(n1404) );
INV_X1 U1126 ( .A(G953), .ZN(n1124) );
NAND2_X1 U1127 ( .A1(KEYINPUT29), .A2(n1405), .ZN(n1402) );
XNOR2_X1 U1128 ( .A(n1241), .B(n1375), .ZN(n1405) );
XOR2_X1 U1129 ( .A(G140), .B(KEYINPUT30), .Z(n1375) );
INV_X1 U1130 ( .A(G125), .ZN(n1241) );
XOR2_X1 U1131 ( .A(n1406), .B(n1407), .Z(n1400) );
XNOR2_X1 U1132 ( .A(n1408), .B(G137), .ZN(n1407) );
INV_X1 U1133 ( .A(G146), .ZN(n1408) );
XNOR2_X1 U1134 ( .A(G119), .B(G128), .ZN(n1406) );
endmodule


