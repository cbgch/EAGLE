//Key = 1111011011000000100101100111100011010100000001100011010110011101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337;

XNOR2_X1 U734 ( .A(n1012), .B(n1013), .ZN(G9) );
NOR2_X1 U735 ( .A1(KEYINPUT47), .A2(n1014), .ZN(n1013) );
INV_X1 U736 ( .A(n1015), .ZN(n1014) );
NOR2_X1 U737 ( .A1(n1016), .A2(n1017), .ZN(G75) );
XOR2_X1 U738 ( .A(KEYINPUT40), .B(n1018), .Z(n1017) );
NOR4_X1 U739 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
NOR2_X1 U740 ( .A1(n1023), .A2(n1024), .ZN(n1019) );
NOR2_X1 U741 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U742 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NOR2_X1 U743 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U744 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U745 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U746 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1033) );
XNOR2_X1 U750 ( .A(KEYINPUT56), .B(n1043), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1044), .A2(n1043), .ZN(n1029) );
NOR2_X1 U752 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U753 ( .A1(n1036), .A2(n1047), .ZN(n1045) );
NOR4_X1 U754 ( .A1(n1048), .A2(n1032), .A3(n1043), .A4(n1036), .ZN(n1025) );
NOR2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U756 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U757 ( .A1(G952), .A2(n1020), .ZN(n1016) );
NAND2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1020) );
NAND4_X1 U759 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NOR2_X1 U760 ( .A1(n1028), .A2(n1036), .ZN(n1058) );
INV_X1 U761 ( .A(n1043), .ZN(n1057) );
XOR2_X1 U762 ( .A(n1059), .B(n1060), .Z(n1056) );
NAND2_X1 U763 ( .A1(KEYINPUT50), .A2(n1061), .ZN(n1060) );
XOR2_X1 U764 ( .A(n1062), .B(n1063), .Z(G72) );
XOR2_X1 U765 ( .A(n1064), .B(n1065), .Z(n1063) );
NOR3_X1 U766 ( .A1(n1066), .A2(KEYINPUT52), .A3(G953), .ZN(n1065) );
NOR2_X1 U767 ( .A1(n1067), .A2(n1068), .ZN(n1064) );
XNOR2_X1 U768 ( .A(n1069), .B(n1070), .ZN(n1068) );
XNOR2_X1 U769 ( .A(n1071), .B(n1072), .ZN(n1069) );
NAND3_X1 U770 ( .A1(n1073), .A2(n1074), .A3(KEYINPUT6), .ZN(n1071) );
OR3_X1 U771 ( .A1(n1075), .A2(n1076), .A3(KEYINPUT3), .ZN(n1074) );
NAND2_X1 U772 ( .A1(n1077), .A2(KEYINPUT3), .ZN(n1073) );
XOR2_X1 U773 ( .A(n1076), .B(n1075), .Z(n1077) );
XOR2_X1 U774 ( .A(G134), .B(n1078), .Z(n1075) );
NOR2_X1 U775 ( .A1(KEYINPUT44), .A2(n1079), .ZN(n1078) );
NOR2_X1 U776 ( .A1(G900), .A2(n1053), .ZN(n1067) );
NOR2_X1 U777 ( .A1(n1080), .A2(n1053), .ZN(n1062) );
AND2_X1 U778 ( .A1(G227), .A2(G900), .ZN(n1080) );
NAND2_X1 U779 ( .A1(n1081), .A2(n1082), .ZN(G69) );
NAND2_X1 U780 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U781 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NAND3_X1 U782 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NAND2_X1 U783 ( .A1(G953), .A2(n1090), .ZN(n1088) );
NAND3_X1 U784 ( .A1(n1091), .A2(n1085), .A3(n1092), .ZN(n1081) );
NAND2_X1 U785 ( .A1(n1089), .A2(n1087), .ZN(n1092) );
NAND3_X1 U786 ( .A1(n1021), .A2(n1053), .A3(n1093), .ZN(n1085) );
XOR2_X1 U787 ( .A(KEYINPUT55), .B(n1089), .Z(n1093) );
AND3_X1 U788 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1089) );
INV_X1 U789 ( .A(n1097), .ZN(n1096) );
NAND2_X1 U790 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
NAND2_X1 U791 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND3_X1 U792 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1094) );
XNOR2_X1 U793 ( .A(KEYINPUT26), .B(n1103), .ZN(n1100) );
NAND2_X1 U794 ( .A1(n1104), .A2(n1084), .ZN(n1091) );
INV_X1 U795 ( .A(KEYINPUT24), .ZN(n1084) );
NAND2_X1 U796 ( .A1(G953), .A2(n1105), .ZN(n1104) );
NAND2_X1 U797 ( .A1(G898), .A2(G224), .ZN(n1105) );
NOR2_X1 U798 ( .A1(n1106), .A2(n1107), .ZN(G66) );
XOR2_X1 U799 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U800 ( .A1(KEYINPUT49), .A2(n1110), .ZN(n1109) );
OR2_X1 U801 ( .A1(n1111), .A2(n1061), .ZN(n1108) );
NOR2_X1 U802 ( .A1(n1106), .A2(n1112), .ZN(G63) );
XOR2_X1 U803 ( .A(n1113), .B(n1114), .Z(n1112) );
AND2_X1 U804 ( .A1(G478), .A2(n1115), .ZN(n1113) );
NOR2_X1 U805 ( .A1(n1106), .A2(n1116), .ZN(G60) );
XOR2_X1 U806 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR3_X1 U807 ( .A1(n1111), .A2(KEYINPUT4), .A3(n1119), .ZN(n1117) );
NAND2_X1 U808 ( .A1(n1120), .A2(n1121), .ZN(G6) );
NAND2_X1 U809 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XOR2_X1 U810 ( .A(KEYINPUT1), .B(n1124), .Z(n1120) );
NOR2_X1 U811 ( .A1(n1122), .A2(n1123), .ZN(n1124) );
NAND4_X1 U812 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1123) );
XNOR2_X1 U813 ( .A(n1050), .B(KEYINPUT19), .ZN(n1125) );
XNOR2_X1 U814 ( .A(KEYINPUT45), .B(G104), .ZN(n1122) );
NOR2_X1 U815 ( .A1(n1106), .A2(n1129), .ZN(G57) );
XOR2_X1 U816 ( .A(n1130), .B(n1131), .Z(n1129) );
XNOR2_X1 U817 ( .A(n1132), .B(n1133), .ZN(n1131) );
NAND3_X1 U818 ( .A1(n1115), .A2(G472), .A3(KEYINPUT33), .ZN(n1132) );
NOR2_X1 U819 ( .A1(n1106), .A2(n1134), .ZN(G54) );
XOR2_X1 U820 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U821 ( .A(n1137), .B(n1138), .Z(n1136) );
XNOR2_X1 U822 ( .A(n1139), .B(n1140), .ZN(n1138) );
NOR2_X1 U823 ( .A1(KEYINPUT14), .A2(n1141), .ZN(n1140) );
XOR2_X1 U824 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U825 ( .A(n1144), .B(G110), .Z(n1143) );
XNOR2_X1 U826 ( .A(G140), .B(KEYINPUT7), .ZN(n1142) );
NAND2_X1 U827 ( .A1(KEYINPUT63), .A2(n1145), .ZN(n1139) );
NOR2_X1 U828 ( .A1(KEYINPUT18), .A2(n1146), .ZN(n1137) );
XOR2_X1 U829 ( .A(n1147), .B(n1148), .Z(n1135) );
NAND2_X1 U830 ( .A1(n1115), .A2(G469), .ZN(n1147) );
NOR2_X1 U831 ( .A1(n1106), .A2(n1149), .ZN(G51) );
XOR2_X1 U832 ( .A(n1150), .B(n1151), .Z(n1149) );
XNOR2_X1 U833 ( .A(n1072), .B(n1152), .ZN(n1151) );
XOR2_X1 U834 ( .A(n1153), .B(n1154), .Z(n1150) );
NOR2_X1 U835 ( .A1(KEYINPUT11), .A2(n1155), .ZN(n1154) );
XOR2_X1 U836 ( .A(n1156), .B(n1157), .Z(n1153) );
NAND2_X1 U837 ( .A1(n1115), .A2(n1158), .ZN(n1156) );
INV_X1 U838 ( .A(n1111), .ZN(n1115) );
NAND2_X1 U839 ( .A1(G902), .A2(n1159), .ZN(n1111) );
NAND2_X1 U840 ( .A1(n1066), .A2(n1087), .ZN(n1159) );
INV_X1 U841 ( .A(n1021), .ZN(n1087) );
NAND4_X1 U842 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1021) );
NOR4_X1 U843 ( .A1(n1164), .A2(n1015), .A3(n1165), .A4(n1166), .ZN(n1163) );
INV_X1 U844 ( .A(n1167), .ZN(n1166) );
NOR3_X1 U845 ( .A1(n1032), .A2(n1168), .A3(n1041), .ZN(n1015) );
NAND2_X1 U846 ( .A1(n1169), .A2(n1046), .ZN(n1162) );
NAND2_X1 U847 ( .A1(n1170), .A2(n1171), .ZN(n1046) );
NAND2_X1 U848 ( .A1(n1126), .A2(n1128), .ZN(n1171) );
NAND2_X1 U849 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
INV_X1 U850 ( .A(n1168), .ZN(n1169) );
INV_X1 U851 ( .A(n1022), .ZN(n1066) );
NAND4_X1 U852 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1022) );
NOR4_X1 U853 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1177) );
NOR2_X1 U854 ( .A1(n1182), .A2(n1183), .ZN(n1176) );
NOR2_X1 U855 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR3_X1 U856 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1182) );
XNOR2_X1 U857 ( .A(KEYINPUT32), .B(n1036), .ZN(n1186) );
NOR2_X1 U858 ( .A1(n1053), .A2(G952), .ZN(n1106) );
NAND2_X1 U859 ( .A1(n1189), .A2(n1190), .ZN(G48) );
NAND2_X1 U860 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U861 ( .A(KEYINPUT9), .B(n1193), .Z(n1189) );
NOR2_X1 U862 ( .A1(n1191), .A2(n1192), .ZN(n1193) );
INV_X1 U863 ( .A(n1175), .ZN(n1191) );
NAND3_X1 U864 ( .A1(n1194), .A2(n1128), .A3(n1195), .ZN(n1175) );
XNOR2_X1 U865 ( .A(G143), .B(n1174), .ZN(G45) );
NAND4_X1 U866 ( .A1(n1196), .A2(n1195), .A3(n1197), .A4(n1198), .ZN(n1174) );
XNOR2_X1 U867 ( .A(G140), .B(n1199), .ZN(G42) );
NAND2_X1 U868 ( .A1(KEYINPUT35), .A2(n1181), .ZN(n1199) );
AND3_X1 U869 ( .A1(n1200), .A2(n1128), .A3(n1172), .ZN(n1181) );
XNOR2_X1 U870 ( .A(G137), .B(n1201), .ZN(G39) );
NAND2_X1 U871 ( .A1(n1202), .A2(n1200), .ZN(n1201) );
XNOR2_X1 U872 ( .A(n1203), .B(n1180), .ZN(G36) );
NOR3_X1 U873 ( .A1(n1047), .A2(n1041), .A3(n1188), .ZN(n1180) );
INV_X1 U874 ( .A(n1200), .ZN(n1188) );
INV_X1 U875 ( .A(n1204), .ZN(n1041) );
XOR2_X1 U876 ( .A(n1179), .B(n1205), .Z(G33) );
NOR2_X1 U877 ( .A1(KEYINPUT38), .A2(n1206), .ZN(n1205) );
INV_X1 U878 ( .A(G131), .ZN(n1206) );
AND3_X1 U879 ( .A1(n1196), .A2(n1128), .A3(n1200), .ZN(n1179) );
NOR3_X1 U880 ( .A1(n1207), .A2(n1184), .A3(n1043), .ZN(n1200) );
NAND2_X1 U881 ( .A1(n1208), .A2(n1040), .ZN(n1043) );
INV_X1 U882 ( .A(n1039), .ZN(n1208) );
XNOR2_X1 U883 ( .A(n1178), .B(n1209), .ZN(G30) );
XNOR2_X1 U884 ( .A(G128), .B(KEYINPUT10), .ZN(n1209) );
AND3_X1 U885 ( .A1(n1194), .A2(n1204), .A3(n1195), .ZN(n1178) );
AND3_X1 U886 ( .A1(n1038), .A2(n1210), .A3(n1050), .ZN(n1195) );
INV_X1 U887 ( .A(n1187), .ZN(n1194) );
XNOR2_X1 U888 ( .A(n1211), .B(n1164), .ZN(G3) );
NOR3_X1 U889 ( .A1(n1036), .A2(n1168), .A3(n1047), .ZN(n1164) );
XNOR2_X1 U890 ( .A(n1155), .B(n1212), .ZN(G27) );
NOR2_X1 U891 ( .A1(n1213), .A2(n1185), .ZN(n1212) );
NAND4_X1 U892 ( .A1(n1172), .A2(n1214), .A3(n1038), .A4(n1128), .ZN(n1185) );
INV_X1 U893 ( .A(n1215), .ZN(n1172) );
XNOR2_X1 U894 ( .A(n1184), .B(KEYINPUT51), .ZN(n1213) );
INV_X1 U895 ( .A(n1210), .ZN(n1184) );
NAND2_X1 U896 ( .A1(n1024), .A2(n1216), .ZN(n1210) );
NAND4_X1 U897 ( .A1(G902), .A2(G953), .A3(n1217), .A4(n1218), .ZN(n1216) );
INV_X1 U898 ( .A(G900), .ZN(n1218) );
XNOR2_X1 U899 ( .A(G122), .B(n1160), .ZN(G24) );
NAND4_X1 U900 ( .A1(n1219), .A2(n1126), .A3(n1197), .A4(n1198), .ZN(n1160) );
INV_X1 U901 ( .A(n1032), .ZN(n1126) );
NAND2_X1 U902 ( .A1(n1055), .A2(n1220), .ZN(n1032) );
XNOR2_X1 U903 ( .A(G119), .B(n1161), .ZN(G21) );
NAND2_X1 U904 ( .A1(n1202), .A2(n1219), .ZN(n1161) );
NOR2_X1 U905 ( .A1(n1187), .A2(n1036), .ZN(n1202) );
NAND2_X1 U906 ( .A1(n1221), .A2(n1222), .ZN(n1187) );
XOR2_X1 U907 ( .A(G116), .B(n1223), .Z(G18) );
NOR2_X1 U908 ( .A1(KEYINPUT36), .A2(n1167), .ZN(n1223) );
NAND3_X1 U909 ( .A1(n1196), .A2(n1204), .A3(n1219), .ZN(n1167) );
NOR2_X1 U910 ( .A1(n1198), .A2(n1224), .ZN(n1204) );
XOR2_X1 U911 ( .A(G113), .B(n1165), .Z(G15) );
AND3_X1 U912 ( .A1(n1196), .A2(n1128), .A3(n1219), .ZN(n1165) );
AND2_X1 U913 ( .A1(n1214), .A2(n1127), .ZN(n1219) );
INV_X1 U914 ( .A(n1028), .ZN(n1214) );
NAND2_X1 U915 ( .A1(n1225), .A2(n1052), .ZN(n1028) );
INV_X1 U916 ( .A(n1051), .ZN(n1225) );
NAND2_X1 U917 ( .A1(n1226), .A2(n1227), .ZN(n1128) );
NAND3_X1 U918 ( .A1(n1198), .A2(n1224), .A3(n1228), .ZN(n1227) );
INV_X1 U919 ( .A(KEYINPUT13), .ZN(n1228) );
INV_X1 U920 ( .A(n1197), .ZN(n1224) );
NAND2_X1 U921 ( .A1(KEYINPUT13), .A2(n1173), .ZN(n1226) );
INV_X1 U922 ( .A(n1047), .ZN(n1196) );
NAND2_X1 U923 ( .A1(n1229), .A2(n1220), .ZN(n1047) );
INV_X1 U924 ( .A(n1222), .ZN(n1220) );
XNOR2_X1 U925 ( .A(n1221), .B(KEYINPUT46), .ZN(n1229) );
XNOR2_X1 U926 ( .A(n1055), .B(KEYINPUT17), .ZN(n1221) );
XOR2_X1 U927 ( .A(G110), .B(n1230), .Z(G12) );
NOR4_X1 U928 ( .A1(KEYINPUT54), .A2(n1168), .A3(n1036), .A4(n1215), .ZN(n1230) );
NAND2_X1 U929 ( .A1(n1055), .A2(n1222), .ZN(n1215) );
XOR2_X1 U930 ( .A(n1059), .B(n1061), .Z(n1222) );
NAND2_X1 U931 ( .A1(G217), .A2(n1231), .ZN(n1061) );
OR2_X1 U932 ( .A1(n1110), .A2(G902), .ZN(n1059) );
XOR2_X1 U933 ( .A(n1232), .B(n1233), .Z(n1110) );
XOR2_X1 U934 ( .A(n1234), .B(n1235), .Z(n1233) );
NAND2_X1 U935 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U936 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
XOR2_X1 U937 ( .A(KEYINPUT21), .B(n1079), .Z(n1238) );
NAND2_X1 U938 ( .A1(n1079), .A2(n1240), .ZN(n1236) );
INV_X1 U939 ( .A(n1239), .ZN(n1240) );
NAND3_X1 U940 ( .A1(G221), .A2(G234), .A3(n1241), .ZN(n1239) );
XNOR2_X1 U941 ( .A(G953), .B(KEYINPUT43), .ZN(n1241) );
NAND3_X1 U942 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1234) );
NAND2_X1 U943 ( .A1(KEYINPUT62), .A2(G146), .ZN(n1244) );
OR3_X1 U944 ( .A1(n1245), .A2(KEYINPUT62), .A3(n1246), .ZN(n1243) );
NAND2_X1 U945 ( .A1(n1246), .A2(n1245), .ZN(n1242) );
NAND2_X1 U946 ( .A1(KEYINPUT16), .A2(n1192), .ZN(n1245) );
INV_X1 U947 ( .A(G146), .ZN(n1192) );
XOR2_X1 U948 ( .A(n1247), .B(KEYINPUT59), .Z(n1246) );
XOR2_X1 U949 ( .A(n1248), .B(n1249), .Z(n1232) );
NOR2_X1 U950 ( .A1(G110), .A2(KEYINPUT15), .ZN(n1249) );
XNOR2_X1 U951 ( .A(G119), .B(G128), .ZN(n1248) );
XOR2_X1 U952 ( .A(n1250), .B(G472), .Z(n1055) );
NAND3_X1 U953 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1250) );
NAND2_X1 U954 ( .A1(n1254), .A2(n1255), .ZN(n1252) );
XNOR2_X1 U955 ( .A(n1256), .B(n1257), .ZN(n1254) );
INV_X1 U956 ( .A(n1133), .ZN(n1256) );
OR3_X1 U957 ( .A1(n1257), .A2(n1133), .A3(n1255), .ZN(n1251) );
INV_X1 U958 ( .A(KEYINPUT20), .ZN(n1255) );
XOR2_X1 U959 ( .A(n1258), .B(n1211), .Z(n1133) );
INV_X1 U960 ( .A(G101), .ZN(n1211) );
NAND3_X1 U961 ( .A1(G210), .A2(n1053), .A3(n1259), .ZN(n1258) );
XOR2_X1 U962 ( .A(n1260), .B(KEYINPUT34), .Z(n1259) );
XOR2_X1 U963 ( .A(n1130), .B(KEYINPUT48), .Z(n1257) );
XOR2_X1 U964 ( .A(n1261), .B(n1262), .Z(n1130) );
INV_X1 U965 ( .A(n1263), .ZN(n1262) );
XNOR2_X1 U966 ( .A(G113), .B(n1264), .ZN(n1261) );
INV_X1 U967 ( .A(n1173), .ZN(n1036) );
NOR2_X1 U968 ( .A1(n1197), .A2(n1198), .ZN(n1173) );
XOR2_X1 U969 ( .A(n1265), .B(n1119), .Z(n1198) );
INV_X1 U970 ( .A(G475), .ZN(n1119) );
OR2_X1 U971 ( .A1(n1118), .A2(G902), .ZN(n1265) );
XNOR2_X1 U972 ( .A(n1266), .B(n1267), .ZN(n1118) );
XOR2_X1 U973 ( .A(G113), .B(G104), .Z(n1267) );
XOR2_X1 U974 ( .A(n1268), .B(n1269), .Z(n1266) );
NOR2_X1 U975 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NOR2_X1 U976 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NOR2_X1 U977 ( .A1(KEYINPUT57), .A2(n1070), .ZN(n1273) );
NOR2_X1 U978 ( .A1(G146), .A2(n1274), .ZN(n1272) );
NOR2_X1 U979 ( .A1(KEYINPUT8), .A2(n1247), .ZN(n1274) );
NOR4_X1 U980 ( .A1(KEYINPUT57), .A2(G146), .A3(n1070), .A4(n1275), .ZN(n1270) );
INV_X1 U981 ( .A(KEYINPUT8), .ZN(n1275) );
INV_X1 U982 ( .A(n1247), .ZN(n1070) );
XNOR2_X1 U983 ( .A(G140), .B(n1155), .ZN(n1247) );
XOR2_X1 U984 ( .A(n1276), .B(n1277), .Z(n1268) );
XNOR2_X1 U985 ( .A(G143), .B(n1278), .ZN(n1277) );
XNOR2_X1 U986 ( .A(KEYINPUT28), .B(KEYINPUT12), .ZN(n1278) );
XOR2_X1 U987 ( .A(n1279), .B(n1076), .Z(n1276) );
XNOR2_X1 U988 ( .A(n1280), .B(n1281), .ZN(n1279) );
NAND3_X1 U989 ( .A1(n1260), .A2(n1053), .A3(G214), .ZN(n1280) );
XNOR2_X1 U990 ( .A(G237), .B(KEYINPUT41), .ZN(n1260) );
XNOR2_X1 U991 ( .A(n1282), .B(G478), .ZN(n1197) );
OR2_X1 U992 ( .A1(n1114), .A2(G902), .ZN(n1282) );
XNOR2_X1 U993 ( .A(n1283), .B(n1284), .ZN(n1114) );
XOR2_X1 U994 ( .A(n1285), .B(n1286), .Z(n1284) );
NAND3_X1 U995 ( .A1(G217), .A2(n1053), .A3(G234), .ZN(n1286) );
NAND2_X1 U996 ( .A1(n1287), .A2(KEYINPUT27), .ZN(n1285) );
XNOR2_X1 U997 ( .A(G134), .B(n1288), .ZN(n1287) );
XNOR2_X1 U998 ( .A(G107), .B(n1289), .ZN(n1283) );
XNOR2_X1 U999 ( .A(n1281), .B(G116), .ZN(n1289) );
INV_X1 U1000 ( .A(G122), .ZN(n1281) );
NAND2_X1 U1001 ( .A1(n1050), .A2(n1127), .ZN(n1168) );
AND2_X1 U1002 ( .A1(n1038), .A2(n1290), .ZN(n1127) );
NAND2_X1 U1003 ( .A1(n1024), .A2(n1291), .ZN(n1290) );
NAND3_X1 U1004 ( .A1(n1097), .A2(n1217), .A3(G902), .ZN(n1291) );
NOR2_X1 U1005 ( .A1(n1053), .A2(G898), .ZN(n1097) );
NAND3_X1 U1006 ( .A1(n1217), .A2(n1053), .A3(G952), .ZN(n1024) );
NAND2_X1 U1007 ( .A1(G234), .A2(G237), .ZN(n1217) );
AND2_X1 U1008 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U1009 ( .A1(G214), .A2(n1292), .ZN(n1040) );
XNOR2_X1 U1010 ( .A(n1293), .B(n1158), .ZN(n1039) );
AND2_X1 U1011 ( .A1(G210), .A2(n1292), .ZN(n1158) );
NAND2_X1 U1012 ( .A1(n1253), .A2(n1294), .ZN(n1292) );
INV_X1 U1013 ( .A(G237), .ZN(n1294) );
NAND2_X1 U1014 ( .A1(n1295), .A2(n1253), .ZN(n1293) );
XOR2_X1 U1015 ( .A(n1296), .B(n1152), .Z(n1295) );
XNOR2_X1 U1016 ( .A(n1297), .B(n1098), .ZN(n1152) );
INV_X1 U1017 ( .A(n1102), .ZN(n1098) );
XNOR2_X1 U1018 ( .A(G122), .B(G110), .ZN(n1102) );
NAND2_X1 U1019 ( .A1(n1101), .A2(n1103), .ZN(n1297) );
NAND2_X1 U1020 ( .A1(n1298), .A2(n1299), .ZN(n1103) );
XNOR2_X1 U1021 ( .A(n1264), .B(n1300), .ZN(n1299) );
INV_X1 U1022 ( .A(n1301), .ZN(n1264) );
XNOR2_X1 U1023 ( .A(n1302), .B(n1303), .ZN(n1298) );
NAND2_X1 U1024 ( .A1(n1304), .A2(n1305), .ZN(n1101) );
XNOR2_X1 U1025 ( .A(n1300), .B(n1301), .ZN(n1305) );
XNOR2_X1 U1026 ( .A(G116), .B(G119), .ZN(n1301) );
NOR2_X1 U1027 ( .A1(KEYINPUT31), .A2(n1306), .ZN(n1300) );
XOR2_X1 U1028 ( .A(KEYINPUT30), .B(G113), .Z(n1306) );
XNOR2_X1 U1029 ( .A(n1302), .B(n1307), .ZN(n1304) );
NAND2_X1 U1030 ( .A1(KEYINPUT2), .A2(n1308), .ZN(n1302) );
NAND2_X1 U1031 ( .A1(n1309), .A2(n1310), .ZN(n1296) );
NAND2_X1 U1032 ( .A1(n1072), .A2(n1311), .ZN(n1310) );
NAND2_X1 U1033 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NAND2_X1 U1034 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
XNOR2_X1 U1035 ( .A(KEYINPUT23), .B(n1155), .ZN(n1314) );
NAND2_X1 U1036 ( .A1(n1316), .A2(n1317), .ZN(n1312) );
XNOR2_X1 U1037 ( .A(KEYINPUT23), .B(G125), .ZN(n1316) );
INV_X1 U1038 ( .A(n1145), .ZN(n1072) );
NAND2_X1 U1039 ( .A1(n1318), .A2(n1145), .ZN(n1309) );
NAND2_X1 U1040 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
NAND2_X1 U1041 ( .A1(n1315), .A2(n1155), .ZN(n1320) );
INV_X1 U1042 ( .A(G125), .ZN(n1155) );
XOR2_X1 U1043 ( .A(KEYINPUT37), .B(n1157), .Z(n1315) );
NAND2_X1 U1044 ( .A1(n1317), .A2(G125), .ZN(n1319) );
XNOR2_X1 U1045 ( .A(KEYINPUT0), .B(n1157), .ZN(n1317) );
NOR2_X1 U1046 ( .A1(n1090), .A2(G953), .ZN(n1157) );
INV_X1 U1047 ( .A(G224), .ZN(n1090) );
INV_X1 U1048 ( .A(n1207), .ZN(n1050) );
NAND2_X1 U1049 ( .A1(n1051), .A2(n1052), .ZN(n1207) );
NAND2_X1 U1050 ( .A1(G221), .A2(n1231), .ZN(n1052) );
NAND2_X1 U1051 ( .A1(G234), .A2(n1253), .ZN(n1231) );
XNOR2_X1 U1052 ( .A(n1321), .B(G469), .ZN(n1051) );
NAND2_X1 U1053 ( .A1(n1322), .A2(n1253), .ZN(n1321) );
INV_X1 U1054 ( .A(G902), .ZN(n1253) );
XNOR2_X1 U1055 ( .A(n1323), .B(n1144), .ZN(n1322) );
NAND2_X1 U1056 ( .A1(n1324), .A2(n1053), .ZN(n1144) );
INV_X1 U1057 ( .A(G953), .ZN(n1053) );
XNOR2_X1 U1058 ( .A(G227), .B(KEYINPUT5), .ZN(n1324) );
XOR2_X1 U1059 ( .A(n1325), .B(n1326), .Z(n1323) );
NOR3_X1 U1060 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1326) );
NOR2_X1 U1061 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
AND3_X1 U1062 ( .A1(n1331), .A2(n1330), .A3(KEYINPUT25), .ZN(n1328) );
NOR2_X1 U1063 ( .A1(G110), .A2(KEYINPUT29), .ZN(n1330) );
INV_X1 U1064 ( .A(G140), .ZN(n1331) );
NOR2_X1 U1065 ( .A1(KEYINPUT25), .A2(n1332), .ZN(n1327) );
INV_X1 U1066 ( .A(G110), .ZN(n1332) );
NAND2_X1 U1067 ( .A1(n1333), .A2(KEYINPUT60), .ZN(n1325) );
XNOR2_X1 U1068 ( .A(n1263), .B(n1334), .ZN(n1333) );
XOR2_X1 U1069 ( .A(KEYINPUT39), .B(n1148), .Z(n1334) );
XNOR2_X1 U1070 ( .A(n1308), .B(n1335), .ZN(n1148) );
XNOR2_X1 U1071 ( .A(KEYINPUT53), .B(n1303), .ZN(n1335) );
INV_X1 U1072 ( .A(n1307), .ZN(n1303) );
XNOR2_X1 U1073 ( .A(G101), .B(n1012), .ZN(n1307) );
INV_X1 U1074 ( .A(G107), .ZN(n1012) );
XNOR2_X1 U1075 ( .A(G104), .B(KEYINPUT42), .ZN(n1308) );
XOR2_X1 U1076 ( .A(n1145), .B(n1146), .Z(n1263) );
XNOR2_X1 U1077 ( .A(n1336), .B(n1076), .ZN(n1146) );
XOR2_X1 U1078 ( .A(G131), .B(KEYINPUT22), .Z(n1076) );
NAND2_X1 U1079 ( .A1(KEYINPUT61), .A2(n1337), .ZN(n1336) );
XNOR2_X1 U1080 ( .A(n1203), .B(n1079), .ZN(n1337) );
XOR2_X1 U1081 ( .A(G137), .B(KEYINPUT58), .Z(n1079) );
INV_X1 U1082 ( .A(G134), .ZN(n1203) );
XOR2_X1 U1083 ( .A(G146), .B(n1288), .Z(n1145) );
XOR2_X1 U1084 ( .A(G128), .B(G143), .Z(n1288) );
endmodule


