//Key = 1000011100001001110010000010110101011011001100010001110111100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347;

XOR2_X1 U740 ( .A(n1024), .B(G107), .Z(G9) );
NAND2_X1 U741 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
OR2_X1 U742 ( .A1(n1027), .A2(KEYINPUT44), .ZN(n1026) );
NAND3_X1 U743 ( .A1(n1028), .A2(n1029), .A3(KEYINPUT44), .ZN(n1025) );
NOR2_X1 U744 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U745 ( .A1(G953), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1031) );
NOR2_X1 U746 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR3_X1 U750 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1028), .A2(n1046), .ZN(n1044) );
NOR3_X1 U752 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
XNOR2_X1 U753 ( .A(KEYINPUT11), .B(n1050), .ZN(n1047) );
NOR2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1041) );
NOR2_X1 U755 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U756 ( .A1(n1055), .A2(n1043), .ZN(n1054) );
NOR2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U758 ( .A1(n1058), .A2(n1045), .ZN(n1053) );
NOR2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR4_X1 U760 ( .A1(n1061), .A2(n1045), .A3(n1052), .A4(n1043), .ZN(n1037) );
INV_X1 U761 ( .A(n1062), .ZN(n1043) );
INV_X1 U762 ( .A(n1063), .ZN(n1045) );
NOR2_X1 U763 ( .A1(n1064), .A2(n1065), .ZN(n1061) );
NOR2_X1 U764 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
INV_X1 U765 ( .A(n1068), .ZN(n1035) );
NOR3_X1 U766 ( .A1(n1032), .A2(G953), .A3(G952), .ZN(n1030) );
AND4_X1 U767 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1032) );
NOR3_X1 U768 ( .A1(n1052), .A2(n1073), .A3(n1074), .ZN(n1072) );
XOR2_X1 U769 ( .A(n1075), .B(n1076), .Z(n1073) );
XNOR2_X1 U770 ( .A(KEYINPUT36), .B(n1077), .ZN(n1076) );
XOR2_X1 U771 ( .A(n1078), .B(KEYINPUT58), .Z(n1071) );
NAND2_X1 U772 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XNOR2_X1 U773 ( .A(KEYINPUT31), .B(n1081), .ZN(n1079) );
XNOR2_X1 U774 ( .A(n1082), .B(KEYINPUT21), .ZN(n1069) );
XOR2_X1 U775 ( .A(n1083), .B(n1084), .Z(G72) );
NOR2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
AND3_X1 U777 ( .A1(G953), .A2(G227), .A3(G900), .ZN(n1086) );
NOR2_X1 U778 ( .A1(G953), .A2(n1087), .ZN(n1085) );
NOR2_X1 U779 ( .A1(n1088), .A2(KEYINPUT34), .ZN(n1087) );
NOR2_X1 U780 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1083) );
XOR2_X1 U782 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U783 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND2_X1 U784 ( .A1(KEYINPUT47), .A2(n1097), .ZN(n1096) );
INV_X1 U785 ( .A(G131), .ZN(n1097) );
XNOR2_X1 U786 ( .A(n1098), .B(n1099), .ZN(n1093) );
NOR2_X1 U787 ( .A1(G900), .A2(n1100), .ZN(n1091) );
NAND2_X1 U788 ( .A1(n1101), .A2(n1102), .ZN(G69) );
NAND2_X1 U789 ( .A1(n1103), .A2(G953), .ZN(n1102) );
XOR2_X1 U790 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U791 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U792 ( .A1(n1108), .A2(n1100), .ZN(n1101) );
NAND2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U794 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
OR2_X1 U795 ( .A1(n1104), .A2(n1111), .ZN(n1109) );
NAND3_X1 U796 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1111) );
XOR2_X1 U797 ( .A(n1116), .B(KEYINPUT17), .Z(n1115) );
INV_X1 U798 ( .A(n1117), .ZN(n1113) );
XOR2_X1 U799 ( .A(n1112), .B(KEYINPUT3), .Z(n1104) );
NAND2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(n1112) );
NAND2_X1 U801 ( .A1(G953), .A2(n1107), .ZN(n1119) );
XNOR2_X1 U802 ( .A(n1120), .B(n1121), .ZN(n1118) );
NAND2_X1 U803 ( .A1(KEYINPUT6), .A2(n1122), .ZN(n1120) );
XOR2_X1 U804 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U805 ( .A(KEYINPUT43), .B(KEYINPUT41), .Z(n1124) );
NOR3_X1 U806 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(G66) );
AND2_X1 U807 ( .A1(KEYINPUT51), .A2(n1128), .ZN(n1127) );
NOR3_X1 U808 ( .A1(KEYINPUT51), .A2(n1100), .A3(n1129), .ZN(n1126) );
INV_X1 U809 ( .A(G952), .ZN(n1129) );
XNOR2_X1 U810 ( .A(n1130), .B(n1131), .ZN(n1125) );
XOR2_X1 U811 ( .A(KEYINPUT25), .B(n1132), .Z(n1131) );
NOR2_X1 U812 ( .A1(n1077), .A2(n1133), .ZN(n1132) );
NOR2_X1 U813 ( .A1(n1128), .A2(n1134), .ZN(G63) );
XOR2_X1 U814 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U815 ( .A1(n1137), .A2(KEYINPUT37), .ZN(n1136) );
NOR2_X1 U816 ( .A1(n1138), .A2(n1133), .ZN(n1137) );
NOR2_X1 U817 ( .A1(n1128), .A2(n1139), .ZN(G60) );
XOR2_X1 U818 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U819 ( .A1(n1142), .A2(n1133), .ZN(n1140) );
NAND2_X1 U820 ( .A1(n1143), .A2(n1144), .ZN(G6) );
OR2_X1 U821 ( .A1(n1145), .A2(G104), .ZN(n1144) );
NAND2_X1 U822 ( .A1(G104), .A2(n1146), .ZN(n1143) );
NAND2_X1 U823 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
OR2_X1 U824 ( .A1(n1149), .A2(KEYINPUT5), .ZN(n1148) );
NAND2_X1 U825 ( .A1(KEYINPUT5), .A2(n1145), .ZN(n1147) );
OR2_X1 U826 ( .A1(KEYINPUT23), .A2(n1149), .ZN(n1145) );
NOR2_X1 U827 ( .A1(n1128), .A2(n1150), .ZN(G57) );
XOR2_X1 U828 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U829 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U830 ( .A(n1155), .B(n1156), .Z(n1151) );
NOR2_X1 U831 ( .A1(n1157), .A2(n1133), .ZN(n1156) );
NAND2_X1 U832 ( .A1(n1158), .A2(KEYINPUT56), .ZN(n1155) );
XNOR2_X1 U833 ( .A(n1159), .B(KEYINPUT22), .ZN(n1158) );
NOR2_X1 U834 ( .A1(n1128), .A2(n1160), .ZN(G54) );
XOR2_X1 U835 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U836 ( .A1(n1163), .A2(n1133), .ZN(n1162) );
NAND2_X1 U837 ( .A1(n1164), .A2(KEYINPUT61), .ZN(n1161) );
XOR2_X1 U838 ( .A(n1165), .B(n1166), .Z(n1164) );
XNOR2_X1 U839 ( .A(n1167), .B(n1168), .ZN(n1165) );
NOR2_X1 U840 ( .A1(n1128), .A2(n1169), .ZN(G51) );
XOR2_X1 U841 ( .A(n1170), .B(n1171), .Z(n1169) );
XNOR2_X1 U842 ( .A(n1159), .B(n1172), .ZN(n1171) );
XOR2_X1 U843 ( .A(n1173), .B(n1174), .Z(n1170) );
NOR3_X1 U844 ( .A1(n1133), .A2(n1048), .A3(n1175), .ZN(n1173) );
NAND2_X1 U845 ( .A1(G902), .A2(n1034), .ZN(n1133) );
NAND3_X1 U846 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1034) );
NOR3_X1 U847 ( .A1(n1090), .A2(n1117), .A3(n1116), .ZN(n1178) );
NAND4_X1 U848 ( .A1(n1149), .A2(n1179), .A3(n1180), .A4(n1027), .ZN(n1116) );
OR2_X1 U849 ( .A1(n1029), .A2(n1181), .ZN(n1027) );
NAND4_X1 U850 ( .A1(n1182), .A2(n1063), .A3(n1059), .A4(n1183), .ZN(n1029) );
NAND3_X1 U851 ( .A1(n1060), .A2(n1063), .A3(n1184), .ZN(n1149) );
NAND3_X1 U852 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1117) );
NAND4_X1 U853 ( .A1(n1188), .A2(n1063), .A3(n1082), .A4(n1189), .ZN(n1187) );
NAND4_X1 U854 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1090) );
AND4_X1 U855 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
NAND2_X1 U856 ( .A1(n1028), .A2(n1198), .ZN(n1190) );
XNOR2_X1 U857 ( .A(KEYINPUT54), .B(n1199), .ZN(n1198) );
XNOR2_X1 U858 ( .A(n1089), .B(KEYINPUT48), .ZN(n1177) );
INV_X1 U859 ( .A(n1200), .ZN(n1089) );
XOR2_X1 U860 ( .A(n1114), .B(KEYINPUT30), .Z(n1176) );
NOR2_X1 U861 ( .A1(n1100), .A2(G952), .ZN(n1128) );
XNOR2_X1 U862 ( .A(G146), .B(n1191), .ZN(G48) );
NAND3_X1 U863 ( .A1(n1201), .A2(n1060), .A3(n1202), .ZN(n1191) );
XNOR2_X1 U864 ( .A(G143), .B(n1200), .ZN(G45) );
NAND4_X1 U865 ( .A1(n1202), .A2(n1057), .A3(n1082), .A4(n1189), .ZN(n1200) );
AND3_X1 U866 ( .A1(n1203), .A2(n1028), .A3(n1065), .ZN(n1202) );
NAND3_X1 U867 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(G42) );
NAND2_X1 U868 ( .A1(G140), .A2(n1197), .ZN(n1206) );
NAND2_X1 U869 ( .A1(n1207), .A2(n1208), .ZN(n1205) );
INV_X1 U870 ( .A(KEYINPUT16), .ZN(n1208) );
NAND2_X1 U871 ( .A1(n1209), .A2(n1210), .ZN(n1207) );
XNOR2_X1 U872 ( .A(KEYINPUT35), .B(n1211), .ZN(n1210) );
NAND2_X1 U873 ( .A1(KEYINPUT16), .A2(n1212), .ZN(n1204) );
NAND2_X1 U874 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND3_X1 U875 ( .A1(KEYINPUT35), .A2(n1209), .A3(n1211), .ZN(n1214) );
INV_X1 U876 ( .A(n1197), .ZN(n1209) );
NAND3_X1 U877 ( .A1(n1060), .A2(n1056), .A3(n1215), .ZN(n1197) );
OR2_X1 U878 ( .A1(n1211), .A2(KEYINPUT35), .ZN(n1213) );
XNOR2_X1 U879 ( .A(G137), .B(n1196), .ZN(G39) );
NAND3_X1 U880 ( .A1(n1201), .A2(n1215), .A3(n1062), .ZN(n1196) );
XNOR2_X1 U881 ( .A(n1216), .B(n1217), .ZN(G36) );
NOR2_X1 U882 ( .A1(KEYINPUT2), .A2(n1192), .ZN(n1217) );
NAND3_X1 U883 ( .A1(n1057), .A2(n1059), .A3(n1215), .ZN(n1192) );
XNOR2_X1 U884 ( .A(G131), .B(n1195), .ZN(G33) );
NAND3_X1 U885 ( .A1(n1057), .A2(n1060), .A3(n1215), .ZN(n1195) );
AND3_X1 U886 ( .A1(n1203), .A2(n1218), .A3(n1065), .ZN(n1215) );
XNOR2_X1 U887 ( .A(n1182), .B(KEYINPUT57), .ZN(n1065) );
INV_X1 U888 ( .A(n1052), .ZN(n1218) );
NAND2_X1 U889 ( .A1(n1050), .A2(n1219), .ZN(n1052) );
XOR2_X1 U890 ( .A(G128), .B(n1220), .Z(G30) );
NOR2_X1 U891 ( .A1(n1181), .A2(n1199), .ZN(n1220) );
NAND4_X1 U892 ( .A1(n1201), .A2(n1203), .A3(n1182), .A4(n1059), .ZN(n1199) );
XNOR2_X1 U893 ( .A(G101), .B(n1179), .ZN(G3) );
NAND3_X1 U894 ( .A1(n1062), .A2(n1057), .A3(n1184), .ZN(n1179) );
XNOR2_X1 U895 ( .A(G125), .B(n1194), .ZN(G27) );
NAND4_X1 U896 ( .A1(n1060), .A2(n1203), .A3(n1221), .A4(n1056), .ZN(n1194) );
NOR2_X1 U897 ( .A1(n1181), .A2(n1040), .ZN(n1221) );
INV_X1 U898 ( .A(n1070), .ZN(n1040) );
AND3_X1 U899 ( .A1(n1222), .A2(n1068), .A3(n1223), .ZN(n1203) );
NAND2_X1 U900 ( .A1(n1224), .A2(n1225), .ZN(n1222) );
OR2_X1 U901 ( .A1(n1226), .A2(G900), .ZN(n1225) );
NAND2_X1 U902 ( .A1(G952), .A2(n1227), .ZN(n1224) );
NAND2_X1 U903 ( .A1(G953), .A2(n1228), .ZN(n1227) );
XNOR2_X1 U904 ( .A(G122), .B(n1229), .ZN(G24) );
NAND4_X1 U905 ( .A1(n1230), .A2(n1188), .A3(n1082), .A4(n1189), .ZN(n1229) );
XNOR2_X1 U906 ( .A(n1063), .B(KEYINPUT12), .ZN(n1230) );
NOR2_X1 U907 ( .A1(n1074), .A2(n1231), .ZN(n1063) );
XNOR2_X1 U908 ( .A(G119), .B(n1185), .ZN(G21) );
NAND3_X1 U909 ( .A1(n1062), .A2(n1201), .A3(n1188), .ZN(n1185) );
AND2_X1 U910 ( .A1(n1232), .A2(n1233), .ZN(n1201) );
XNOR2_X1 U911 ( .A(n1074), .B(KEYINPUT52), .ZN(n1232) );
NAND2_X1 U912 ( .A1(n1234), .A2(n1235), .ZN(G18) );
OR2_X1 U913 ( .A1(n1236), .A2(G116), .ZN(n1235) );
NAND2_X1 U914 ( .A1(G116), .A2(n1237), .ZN(n1234) );
NAND2_X1 U915 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
OR2_X1 U916 ( .A1(n1186), .A2(KEYINPUT53), .ZN(n1239) );
NAND2_X1 U917 ( .A1(KEYINPUT53), .A2(n1236), .ZN(n1238) );
OR2_X1 U918 ( .A1(KEYINPUT59), .A2(n1186), .ZN(n1236) );
NAND3_X1 U919 ( .A1(n1057), .A2(n1059), .A3(n1188), .ZN(n1186) );
AND2_X1 U920 ( .A1(n1240), .A2(n1189), .ZN(n1059) );
XNOR2_X1 U921 ( .A(n1082), .B(KEYINPUT60), .ZN(n1240) );
XNOR2_X1 U922 ( .A(G113), .B(n1114), .ZN(G15) );
NAND3_X1 U923 ( .A1(n1057), .A2(n1060), .A3(n1188), .ZN(n1114) );
AND3_X1 U924 ( .A1(n1028), .A2(n1183), .A3(n1070), .ZN(n1188) );
NOR2_X1 U925 ( .A1(n1066), .A2(n1241), .ZN(n1070) );
INV_X1 U926 ( .A(n1067), .ZN(n1241) );
NOR2_X1 U927 ( .A1(n1189), .A2(n1242), .ZN(n1060) );
INV_X1 U928 ( .A(n1082), .ZN(n1242) );
AND2_X1 U929 ( .A1(n1243), .A2(n1074), .ZN(n1057) );
XNOR2_X1 U930 ( .A(KEYINPUT45), .B(n1231), .ZN(n1243) );
INV_X1 U931 ( .A(n1244), .ZN(n1231) );
NAND2_X1 U932 ( .A1(n1245), .A2(n1246), .ZN(G12) );
NAND2_X1 U933 ( .A1(G110), .A2(n1180), .ZN(n1246) );
XOR2_X1 U934 ( .A(n1247), .B(KEYINPUT10), .Z(n1245) );
OR2_X1 U935 ( .A1(n1180), .A2(G110), .ZN(n1247) );
NAND3_X1 U936 ( .A1(n1062), .A2(n1056), .A3(n1184), .ZN(n1180) );
AND3_X1 U937 ( .A1(n1182), .A2(n1183), .A3(n1028), .ZN(n1184) );
INV_X1 U938 ( .A(n1181), .ZN(n1028) );
NAND2_X1 U939 ( .A1(n1248), .A2(n1219), .ZN(n1181) );
NAND2_X1 U940 ( .A1(G214), .A2(n1249), .ZN(n1219) );
XNOR2_X1 U941 ( .A(KEYINPUT4), .B(n1050), .ZN(n1248) );
XOR2_X1 U942 ( .A(n1250), .B(n1251), .Z(n1050) );
NOR2_X1 U943 ( .A1(n1048), .A2(n1175), .ZN(n1251) );
INV_X1 U944 ( .A(G210), .ZN(n1175) );
INV_X1 U945 ( .A(n1249), .ZN(n1048) );
NAND2_X1 U946 ( .A1(n1252), .A2(n1253), .ZN(n1249) );
NAND2_X1 U947 ( .A1(n1254), .A2(n1226), .ZN(n1250) );
XOR2_X1 U948 ( .A(n1172), .B(n1255), .Z(n1254) );
XOR2_X1 U949 ( .A(n1256), .B(n1257), .Z(n1255) );
NOR2_X1 U950 ( .A1(KEYINPUT32), .A2(n1174), .ZN(n1257) );
NOR2_X1 U951 ( .A1(n1106), .A2(G953), .ZN(n1174) );
INV_X1 U952 ( .A(G224), .ZN(n1106) );
NAND2_X1 U953 ( .A1(KEYINPUT15), .A2(n1159), .ZN(n1256) );
XOR2_X1 U954 ( .A(n1258), .B(n1123), .Z(n1172) );
XNOR2_X1 U955 ( .A(n1259), .B(n1260), .ZN(n1123) );
XOR2_X1 U956 ( .A(n1261), .B(KEYINPUT18), .Z(n1259) );
NAND3_X1 U957 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1261) );
INV_X1 U958 ( .A(n1265), .ZN(n1264) );
NAND3_X1 U959 ( .A1(KEYINPUT39), .A2(n1266), .A3(n1267), .ZN(n1263) );
OR2_X1 U960 ( .A1(n1267), .A2(KEYINPUT39), .ZN(n1262) );
XNOR2_X1 U961 ( .A(G125), .B(n1121), .ZN(n1258) );
XNOR2_X1 U962 ( .A(G110), .B(n1268), .ZN(n1121) );
NAND2_X1 U963 ( .A1(n1269), .A2(n1270), .ZN(n1183) );
NAND3_X1 U964 ( .A1(n1271), .A2(n1223), .A3(n1068), .ZN(n1270) );
NAND2_X1 U965 ( .A1(n1272), .A2(n1100), .ZN(n1223) );
NAND2_X1 U966 ( .A1(G952), .A2(n1228), .ZN(n1272) );
INV_X1 U967 ( .A(KEYINPUT62), .ZN(n1228) );
NAND3_X1 U968 ( .A1(n1273), .A2(n1274), .A3(G953), .ZN(n1271) );
NAND3_X1 U969 ( .A1(G902), .A2(n1107), .A3(KEYINPUT7), .ZN(n1274) );
NAND2_X1 U970 ( .A1(KEYINPUT62), .A2(G952), .ZN(n1273) );
NAND2_X1 U971 ( .A1(n1275), .A2(n1276), .ZN(n1269) );
INV_X1 U972 ( .A(KEYINPUT7), .ZN(n1276) );
NAND4_X1 U973 ( .A1(G953), .A2(G902), .A3(n1068), .A4(n1107), .ZN(n1275) );
INV_X1 U974 ( .A(G898), .ZN(n1107) );
NAND2_X1 U975 ( .A1(G237), .A2(G234), .ZN(n1068) );
AND2_X1 U976 ( .A1(n1066), .A2(n1067), .ZN(n1182) );
NAND2_X1 U977 ( .A1(G221), .A2(n1277), .ZN(n1067) );
XOR2_X1 U978 ( .A(n1278), .B(n1163), .Z(n1066) );
INV_X1 U979 ( .A(G469), .ZN(n1163) );
NAND2_X1 U980 ( .A1(n1279), .A2(n1226), .ZN(n1278) );
XNOR2_X1 U981 ( .A(n1280), .B(n1281), .ZN(n1279) );
INV_X1 U982 ( .A(n1167), .ZN(n1281) );
XNOR2_X1 U983 ( .A(n1282), .B(n1283), .ZN(n1167) );
XNOR2_X1 U984 ( .A(n1211), .B(G110), .ZN(n1283) );
INV_X1 U985 ( .A(G140), .ZN(n1211) );
NAND2_X1 U986 ( .A1(G227), .A2(n1100), .ZN(n1282) );
NAND3_X1 U987 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1280) );
NAND2_X1 U988 ( .A1(n1168), .A2(n1287), .ZN(n1286) );
OR3_X1 U989 ( .A1(n1287), .A2(n1168), .A3(KEYINPUT14), .ZN(n1285) );
NAND2_X1 U990 ( .A1(KEYINPUT55), .A2(n1288), .ZN(n1287) );
NAND2_X1 U991 ( .A1(n1166), .A2(KEYINPUT14), .ZN(n1284) );
INV_X1 U992 ( .A(n1288), .ZN(n1166) );
XOR2_X1 U993 ( .A(n1095), .B(n1289), .Z(n1288) );
NOR2_X1 U994 ( .A1(n1265), .A2(n1290), .ZN(n1289) );
XOR2_X1 U995 ( .A(KEYINPUT27), .B(n1291), .Z(n1290) );
AND2_X1 U996 ( .A1(n1266), .A2(n1267), .ZN(n1291) );
NOR2_X1 U997 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XNOR2_X1 U998 ( .A(G107), .B(G104), .ZN(n1267) );
NAND2_X1 U999 ( .A1(n1292), .A2(n1293), .ZN(n1095) );
NAND2_X1 U1000 ( .A1(G128), .A2(n1294), .ZN(n1293) );
XOR2_X1 U1001 ( .A(KEYINPUT28), .B(n1295), .Z(n1292) );
NOR2_X1 U1002 ( .A1(G128), .A2(n1294), .ZN(n1295) );
AND2_X1 U1003 ( .A1(n1233), .A2(n1296), .ZN(n1056) );
INV_X1 U1004 ( .A(n1074), .ZN(n1296) );
XOR2_X1 U1005 ( .A(n1297), .B(n1157), .Z(n1074) );
INV_X1 U1006 ( .A(G472), .ZN(n1157) );
NAND2_X1 U1007 ( .A1(n1298), .A2(n1226), .ZN(n1297) );
XNOR2_X1 U1008 ( .A(n1299), .B(n1300), .ZN(n1298) );
XOR2_X1 U1009 ( .A(n1301), .B(n1153), .Z(n1300) );
XOR2_X1 U1010 ( .A(n1302), .B(n1168), .Z(n1153) );
XNOR2_X1 U1011 ( .A(n1303), .B(n1098), .ZN(n1168) );
XOR2_X1 U1012 ( .A(G137), .B(G134), .Z(n1098) );
XNOR2_X1 U1013 ( .A(G131), .B(KEYINPUT26), .ZN(n1303) );
XNOR2_X1 U1014 ( .A(n1304), .B(n1266), .ZN(n1302) );
INV_X1 U1015 ( .A(G101), .ZN(n1266) );
NAND3_X1 U1016 ( .A1(n1305), .A2(n1253), .A3(G210), .ZN(n1304) );
INV_X1 U1017 ( .A(G237), .ZN(n1253) );
XNOR2_X1 U1018 ( .A(KEYINPUT0), .B(n1100), .ZN(n1305) );
NAND2_X1 U1019 ( .A1(KEYINPUT29), .A2(n1154), .ZN(n1301) );
XOR2_X1 U1020 ( .A(n1260), .B(KEYINPUT50), .Z(n1154) );
XOR2_X1 U1021 ( .A(n1306), .B(n1307), .Z(n1260) );
XNOR2_X1 U1022 ( .A(G119), .B(G113), .ZN(n1306) );
INV_X1 U1023 ( .A(n1159), .ZN(n1299) );
XNOR2_X1 U1024 ( .A(n1308), .B(n1309), .ZN(n1159) );
NOR2_X1 U1025 ( .A1(KEYINPUT46), .A2(n1294), .ZN(n1309) );
XNOR2_X1 U1026 ( .A(G128), .B(KEYINPUT13), .ZN(n1308) );
XNOR2_X1 U1027 ( .A(n1244), .B(KEYINPUT19), .ZN(n1233) );
XOR2_X1 U1028 ( .A(n1310), .B(n1077), .Z(n1244) );
NAND2_X1 U1029 ( .A1(G217), .A2(n1277), .ZN(n1077) );
NAND2_X1 U1030 ( .A1(G234), .A2(n1252), .ZN(n1277) );
XNOR2_X1 U1031 ( .A(G902), .B(KEYINPUT49), .ZN(n1252) );
NAND2_X1 U1032 ( .A1(KEYINPUT20), .A2(n1075), .ZN(n1310) );
NAND2_X1 U1033 ( .A1(n1130), .A2(n1226), .ZN(n1075) );
XNOR2_X1 U1034 ( .A(n1311), .B(n1312), .ZN(n1130) );
XNOR2_X1 U1035 ( .A(n1313), .B(n1314), .ZN(n1312) );
XNOR2_X1 U1036 ( .A(n1315), .B(G128), .ZN(n1314) );
INV_X1 U1037 ( .A(G137), .ZN(n1315) );
INV_X1 U1038 ( .A(G119), .ZN(n1313) );
XOR2_X1 U1039 ( .A(n1316), .B(n1317), .Z(n1311) );
AND3_X1 U1040 ( .A1(G221), .A2(n1100), .A3(G234), .ZN(n1317) );
XOR2_X1 U1041 ( .A(n1318), .B(G110), .Z(n1316) );
NAND2_X1 U1042 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
NAND2_X1 U1043 ( .A1(G146), .A2(n1099), .ZN(n1320) );
XOR2_X1 U1044 ( .A(KEYINPUT33), .B(n1321), .Z(n1319) );
NOR2_X1 U1045 ( .A1(G146), .A2(n1099), .ZN(n1321) );
NOR2_X1 U1046 ( .A1(n1189), .A2(n1082), .ZN(n1062) );
XOR2_X1 U1047 ( .A(n1322), .B(n1142), .Z(n1082) );
INV_X1 U1048 ( .A(G475), .ZN(n1142) );
OR2_X1 U1049 ( .A1(n1141), .A2(G902), .ZN(n1322) );
XNOR2_X1 U1050 ( .A(n1323), .B(n1324), .ZN(n1141) );
XOR2_X1 U1051 ( .A(G104), .B(n1325), .Z(n1324) );
NOR2_X1 U1052 ( .A1(KEYINPUT24), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1053 ( .A(n1327), .B(n1328), .Z(n1326) );
XOR2_X1 U1054 ( .A(n1294), .B(n1099), .Z(n1328) );
XNOR2_X1 U1055 ( .A(n1329), .B(G140), .ZN(n1099) );
INV_X1 U1056 ( .A(G125), .ZN(n1329) );
XOR2_X1 U1057 ( .A(G143), .B(G146), .Z(n1294) );
XOR2_X1 U1058 ( .A(n1330), .B(n1331), .Z(n1327) );
NOR3_X1 U1059 ( .A1(n1049), .A2(G953), .A3(G237), .ZN(n1331) );
INV_X1 U1060 ( .A(G214), .ZN(n1049) );
XNOR2_X1 U1061 ( .A(G131), .B(KEYINPUT8), .ZN(n1330) );
NAND2_X1 U1062 ( .A1(n1332), .A2(n1333), .ZN(n1323) );
NAND2_X1 U1063 ( .A1(G113), .A2(n1268), .ZN(n1333) );
XOR2_X1 U1064 ( .A(n1334), .B(KEYINPUT1), .Z(n1332) );
OR2_X1 U1065 ( .A1(n1268), .A2(G113), .ZN(n1334) );
INV_X1 U1066 ( .A(G122), .ZN(n1268) );
NAND2_X1 U1067 ( .A1(n1081), .A2(n1080), .ZN(n1189) );
NAND3_X1 U1068 ( .A1(n1138), .A2(n1226), .A3(n1135), .ZN(n1080) );
INV_X1 U1069 ( .A(G478), .ZN(n1138) );
NAND2_X1 U1070 ( .A1(G478), .A2(n1335), .ZN(n1081) );
NAND2_X1 U1071 ( .A1(n1135), .A2(n1226), .ZN(n1335) );
INV_X1 U1072 ( .A(G902), .ZN(n1226) );
XOR2_X1 U1073 ( .A(n1336), .B(n1337), .Z(n1135) );
XNOR2_X1 U1074 ( .A(n1338), .B(n1339), .ZN(n1337) );
NOR2_X1 U1075 ( .A1(G107), .A2(KEYINPUT9), .ZN(n1339) );
NAND2_X1 U1076 ( .A1(KEYINPUT38), .A2(n1307), .ZN(n1338) );
XNOR2_X1 U1077 ( .A(G116), .B(KEYINPUT63), .ZN(n1307) );
XOR2_X1 U1078 ( .A(n1340), .B(n1341), .Z(n1336) );
AND3_X1 U1079 ( .A1(G217), .A2(n1100), .A3(G234), .ZN(n1341) );
INV_X1 U1080 ( .A(G953), .ZN(n1100) );
XNOR2_X1 U1081 ( .A(G122), .B(n1342), .ZN(n1340) );
NOR2_X1 U1082 ( .A1(KEYINPUT40), .A2(n1343), .ZN(n1342) );
NOR2_X1 U1083 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
XOR2_X1 U1084 ( .A(n1346), .B(KEYINPUT42), .Z(n1345) );
NAND2_X1 U1085 ( .A1(n1347), .A2(n1216), .ZN(n1346) );
NOR2_X1 U1086 ( .A1(n1347), .A2(n1216), .ZN(n1344) );
INV_X1 U1087 ( .A(G134), .ZN(n1216) );
XNOR2_X1 U1088 ( .A(G143), .B(G128), .ZN(n1347) );
endmodule


