//Key = 1111001100000101010001001111010010010010000110101010100000110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279;

XOR2_X1 U712 ( .A(G107), .B(n980), .Z(G9) );
NOR2_X1 U713 ( .A1(n981), .A2(n982), .ZN(G75) );
NOR4_X1 U714 ( .A1(n983), .A2(n984), .A3(G953), .A4(n985), .ZN(n982) );
NOR2_X1 U715 ( .A1(n986), .A2(n987), .ZN(n984) );
NOR2_X1 U716 ( .A1(n988), .A2(n989), .ZN(n986) );
NOR3_X1 U717 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n989) );
NOR2_X1 U718 ( .A1(n993), .A2(n994), .ZN(n991) );
NOR2_X1 U719 ( .A1(n995), .A2(n996), .ZN(n994) );
NOR3_X1 U720 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n993) );
NOR4_X1 U721 ( .A1(n1000), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(n999) );
AND2_X1 U722 ( .A1(n1004), .A2(KEYINPUT55), .ZN(n1001) );
NOR2_X1 U723 ( .A1(n1005), .A2(n1006), .ZN(n998) );
NOR2_X1 U724 ( .A1(KEYINPUT55), .A2(n996), .ZN(n1005) );
NOR4_X1 U725 ( .A1(n1000), .A2(n1007), .A3(n997), .A4(n996), .ZN(n988) );
INV_X1 U726 ( .A(n1004), .ZN(n996) );
INV_X1 U727 ( .A(n1008), .ZN(n997) );
NOR2_X1 U728 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U729 ( .A1(n1011), .A2(n992), .ZN(n1010) );
NOR3_X1 U730 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1011) );
AND3_X1 U731 ( .A1(KEYINPUT52), .A2(n1015), .A3(n1016), .ZN(n1014) );
NOR2_X1 U732 ( .A1(KEYINPUT52), .A2(n990), .ZN(n1013) );
NOR2_X1 U733 ( .A1(n1017), .A2(n990), .ZN(n1009) );
INV_X1 U734 ( .A(n1018), .ZN(n990) );
NOR2_X1 U735 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NAND2_X1 U736 ( .A1(n1021), .A2(G952), .ZN(n983) );
NOR3_X1 U737 ( .A1(n1022), .A2(G953), .A3(n985), .ZN(n981) );
AND4_X1 U738 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n985) );
NOR4_X1 U739 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
XOR2_X1 U740 ( .A(n1031), .B(n1032), .Z(n1030) );
XNOR2_X1 U741 ( .A(n1033), .B(KEYINPUT5), .ZN(n1032) );
XNOR2_X1 U742 ( .A(G472), .B(n1034), .ZN(n1029) );
XNOR2_X1 U743 ( .A(KEYINPUT57), .B(n1035), .ZN(n1028) );
INV_X1 U744 ( .A(n1036), .ZN(n1035) );
XOR2_X1 U745 ( .A(n1037), .B(KEYINPUT2), .Z(n1027) );
NOR3_X1 U746 ( .A1(n1038), .A2(n1016), .A3(n1000), .ZN(n1025) );
NAND2_X1 U747 ( .A1(n1039), .A2(n1040), .ZN(n1024) );
XOR2_X1 U748 ( .A(KEYINPUT36), .B(G475), .Z(n1039) );
XNOR2_X1 U749 ( .A(KEYINPUT6), .B(n1015), .ZN(n1023) );
XOR2_X1 U750 ( .A(KEYINPUT23), .B(G952), .Z(n1022) );
XOR2_X1 U751 ( .A(n1041), .B(n1042), .Z(G72) );
NOR2_X1 U752 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
AND2_X1 U753 ( .A1(G227), .A2(G900), .ZN(n1043) );
NAND2_X1 U754 ( .A1(n1045), .A2(n1046), .ZN(n1041) );
NAND3_X1 U755 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND2_X1 U756 ( .A1(G953), .A2(n1050), .ZN(n1048) );
OR2_X1 U757 ( .A1(n1047), .A2(n1049), .ZN(n1045) );
NAND2_X1 U758 ( .A1(n1044), .A2(n1051), .ZN(n1049) );
NAND2_X1 U759 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XOR2_X1 U760 ( .A(KEYINPUT56), .B(n1054), .Z(n1053) );
XOR2_X1 U761 ( .A(n1055), .B(n1056), .Z(n1047) );
XOR2_X1 U762 ( .A(KEYINPUT28), .B(n1057), .Z(n1056) );
NOR2_X1 U763 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
XOR2_X1 U764 ( .A(KEYINPUT11), .B(n1060), .Z(n1059) );
NOR2_X1 U765 ( .A1(G140), .A2(n1061), .ZN(n1060) );
XOR2_X1 U766 ( .A(n1062), .B(n1063), .Z(G69) );
NOR2_X1 U767 ( .A1(n1064), .A2(n1044), .ZN(n1063) );
NOR2_X1 U768 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1062) );
NAND2_X1 U770 ( .A1(n1069), .A2(n1044), .ZN(n1068) );
XNOR2_X1 U771 ( .A(n1070), .B(n1071), .ZN(n1069) );
NAND3_X1 U772 ( .A1(G898), .A2(n1071), .A3(G953), .ZN(n1067) );
NOR2_X1 U773 ( .A1(n1072), .A2(n1073), .ZN(G66) );
XOR2_X1 U774 ( .A(n1074), .B(n1075), .Z(n1073) );
NAND2_X1 U775 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U776 ( .A1(n1072), .A2(n1078), .ZN(G63) );
XOR2_X1 U777 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND2_X1 U778 ( .A1(n1076), .A2(G478), .ZN(n1079) );
NOR2_X1 U779 ( .A1(n1072), .A2(n1081), .ZN(G60) );
XOR2_X1 U780 ( .A(n1082), .B(n1083), .Z(n1081) );
NAND2_X1 U781 ( .A1(n1076), .A2(G475), .ZN(n1082) );
XNOR2_X1 U782 ( .A(G104), .B(n1084), .ZN(G6) );
NOR2_X1 U783 ( .A1(n1085), .A2(n1086), .ZN(G57) );
XOR2_X1 U784 ( .A(n1087), .B(n1088), .Z(n1086) );
XOR2_X1 U785 ( .A(n1089), .B(n1090), .Z(n1088) );
NAND2_X1 U786 ( .A1(n1076), .A2(G472), .ZN(n1090) );
NAND3_X1 U787 ( .A1(n1091), .A2(n1092), .A3(KEYINPUT58), .ZN(n1089) );
NAND3_X1 U788 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
INV_X1 U789 ( .A(KEYINPUT32), .ZN(n1095) );
NAND2_X1 U790 ( .A1(n1096), .A2(KEYINPUT32), .ZN(n1091) );
XOR2_X1 U791 ( .A(n1094), .B(n1093), .Z(n1096) );
XNOR2_X1 U792 ( .A(n1097), .B(n1098), .ZN(n1093) );
NOR2_X1 U793 ( .A1(KEYINPUT39), .A2(n1099), .ZN(n1098) );
XNOR2_X1 U794 ( .A(n1072), .B(KEYINPUT3), .ZN(n1085) );
NOR2_X1 U795 ( .A1(n1072), .A2(n1100), .ZN(G54) );
XOR2_X1 U796 ( .A(n1101), .B(n1102), .Z(n1100) );
XNOR2_X1 U797 ( .A(n1103), .B(KEYINPUT47), .ZN(n1102) );
NAND2_X1 U798 ( .A1(n1104), .A2(KEYINPUT44), .ZN(n1103) );
XNOR2_X1 U799 ( .A(n1105), .B(n1106), .ZN(n1104) );
NAND2_X1 U800 ( .A1(n1076), .A2(G469), .ZN(n1101) );
NOR2_X1 U801 ( .A1(n1072), .A2(n1107), .ZN(G51) );
XNOR2_X1 U802 ( .A(n1108), .B(n1071), .ZN(n1107) );
XOR2_X1 U803 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U804 ( .A1(KEYINPUT63), .A2(n1111), .ZN(n1110) );
XNOR2_X1 U805 ( .A(n1112), .B(G125), .ZN(n1111) );
NAND2_X1 U806 ( .A1(n1076), .A2(n1033), .ZN(n1109) );
NOR2_X1 U807 ( .A1(n1113), .A2(n1021), .ZN(n1076) );
AND3_X1 U808 ( .A1(n1054), .A2(n1052), .A3(n1070), .ZN(n1021) );
AND4_X1 U809 ( .A1(n1114), .A2(n1084), .A3(n1115), .A4(n1116), .ZN(n1070) );
NOR4_X1 U810 ( .A1(n980), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1116) );
INV_X1 U811 ( .A(n1120), .ZN(n1119) );
AND3_X1 U812 ( .A1(n1019), .A2(n1004), .A3(n1121), .ZN(n980) );
NOR2_X1 U813 ( .A1(n1122), .A2(n1123), .ZN(n1115) );
INV_X1 U814 ( .A(n1124), .ZN(n1122) );
NAND3_X1 U815 ( .A1(n1121), .A2(n1004), .A3(n1020), .ZN(n1084) );
NAND2_X1 U816 ( .A1(n1125), .A2(n1126), .ZN(n1114) );
XOR2_X1 U817 ( .A(n1127), .B(KEYINPUT50), .Z(n1125) );
AND4_X1 U818 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1052) );
AND4_X1 U819 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1054) );
NAND2_X1 U820 ( .A1(n1136), .A2(n1126), .ZN(n1132) );
XOR2_X1 U821 ( .A(n1137), .B(KEYINPUT46), .Z(n1136) );
NAND4_X1 U822 ( .A1(n1138), .A2(n1020), .A3(n1012), .A4(n1139), .ZN(n1137) );
NOR2_X1 U823 ( .A1(n1044), .A2(G952), .ZN(n1072) );
XNOR2_X1 U824 ( .A(G146), .B(n1140), .ZN(G48) );
NAND3_X1 U825 ( .A1(n1020), .A2(n1141), .A3(n1142), .ZN(n1140) );
XOR2_X1 U826 ( .A(KEYINPUT4), .B(n1138), .Z(n1141) );
XNOR2_X1 U827 ( .A(G143), .B(n1133), .ZN(G45) );
NAND4_X1 U828 ( .A1(n1142), .A2(n1003), .A3(n1036), .A4(n1143), .ZN(n1133) );
XNOR2_X1 U829 ( .A(G140), .B(n1134), .ZN(G42) );
NAND3_X1 U830 ( .A1(n1020), .A2(n1002), .A3(n1144), .ZN(n1134) );
XNOR2_X1 U831 ( .A(G137), .B(n1135), .ZN(G39) );
NAND3_X1 U832 ( .A1(n1138), .A2(n1145), .A3(n1144), .ZN(n1135) );
XNOR2_X1 U833 ( .A(G134), .B(n1128), .ZN(G36) );
NAND3_X1 U834 ( .A1(n1003), .A2(n1019), .A3(n1144), .ZN(n1128) );
XNOR2_X1 U835 ( .A(G131), .B(n1129), .ZN(G33) );
NAND3_X1 U836 ( .A1(n1003), .A2(n1020), .A3(n1144), .ZN(n1129) );
AND4_X1 U837 ( .A1(n1012), .A2(n1008), .A3(n1139), .A4(n1006), .ZN(n1144) );
XNOR2_X1 U838 ( .A(G128), .B(n1130), .ZN(G30) );
NAND3_X1 U839 ( .A1(n1138), .A2(n1019), .A3(n1142), .ZN(n1130) );
AND3_X1 U840 ( .A1(n1126), .A2(n1139), .A3(n1012), .ZN(n1142) );
XNOR2_X1 U841 ( .A(n1146), .B(n1123), .ZN(G3) );
AND3_X1 U842 ( .A1(n1145), .A2(n1121), .A3(n1003), .ZN(n1123) );
XNOR2_X1 U843 ( .A(G125), .B(n1131), .ZN(G27) );
NAND4_X1 U844 ( .A1(n1020), .A2(n1018), .A3(n1147), .A4(n1002), .ZN(n1131) );
AND2_X1 U845 ( .A1(n1139), .A2(n1126), .ZN(n1147) );
NAND2_X1 U846 ( .A1(n987), .A2(n1148), .ZN(n1139) );
NAND4_X1 U847 ( .A1(G953), .A2(G902), .A3(n1149), .A4(n1050), .ZN(n1148) );
INV_X1 U848 ( .A(G900), .ZN(n1050) );
XNOR2_X1 U849 ( .A(G122), .B(n1124), .ZN(G24) );
NAND4_X1 U850 ( .A1(n1150), .A2(n1004), .A3(n1036), .A4(n1143), .ZN(n1124) );
NOR2_X1 U851 ( .A1(n1151), .A2(n1152), .ZN(n1004) );
XNOR2_X1 U852 ( .A(G119), .B(n1120), .ZN(G21) );
NAND3_X1 U853 ( .A1(n1150), .A2(n1145), .A3(n1138), .ZN(n1120) );
AND2_X1 U854 ( .A1(n1153), .A2(n1152), .ZN(n1138) );
XOR2_X1 U855 ( .A(KEYINPUT12), .B(n1154), .Z(n1153) );
XOR2_X1 U856 ( .A(G116), .B(n1155), .Z(G18) );
NOR2_X1 U857 ( .A1(n995), .A2(n1127), .ZN(n1155) );
NAND4_X1 U858 ( .A1(n1003), .A2(n1018), .A3(n1019), .A4(n1156), .ZN(n1127) );
AND2_X1 U859 ( .A1(n1157), .A2(n1036), .ZN(n1019) );
INV_X1 U860 ( .A(n1126), .ZN(n995) );
XNOR2_X1 U861 ( .A(n1158), .B(n1118), .ZN(G15) );
AND3_X1 U862 ( .A1(n1020), .A2(n1150), .A3(n1003), .ZN(n1118) );
NOR2_X1 U863 ( .A1(n1159), .A2(n1152), .ZN(n1003) );
INV_X1 U864 ( .A(n1037), .ZN(n1152) );
XOR2_X1 U865 ( .A(n1154), .B(KEYINPUT26), .Z(n1159) );
XNOR2_X1 U866 ( .A(n1151), .B(KEYINPUT24), .ZN(n1154) );
AND3_X1 U867 ( .A1(n1126), .A2(n1156), .A3(n1018), .ZN(n1150) );
NOR2_X1 U868 ( .A1(n1160), .A2(n1016), .ZN(n1018) );
AND2_X1 U869 ( .A1(n1161), .A2(n1143), .ZN(n1020) );
XOR2_X1 U870 ( .A(G110), .B(n1117), .Z(G12) );
AND3_X1 U871 ( .A1(n1145), .A2(n1121), .A3(n1002), .ZN(n1117) );
NOR2_X1 U872 ( .A1(n1151), .A2(n1037), .ZN(n1002) );
XOR2_X1 U873 ( .A(n1162), .B(n1077), .Z(n1037) );
AND2_X1 U874 ( .A1(G217), .A2(n1163), .ZN(n1077) );
NAND2_X1 U875 ( .A1(n1164), .A2(n1113), .ZN(n1162) );
XNOR2_X1 U876 ( .A(n1075), .B(KEYINPUT17), .ZN(n1164) );
XNOR2_X1 U877 ( .A(n1165), .B(n1166), .ZN(n1075) );
XOR2_X1 U878 ( .A(G137), .B(n1167), .Z(n1166) );
NOR2_X1 U879 ( .A1(KEYINPUT40), .A2(n1168), .ZN(n1167) );
XOR2_X1 U880 ( .A(n1169), .B(n1170), .Z(n1168) );
XNOR2_X1 U881 ( .A(n1171), .B(n1172), .ZN(n1170) );
XNOR2_X1 U882 ( .A(KEYINPUT62), .B(n1173), .ZN(n1172) );
INV_X1 U883 ( .A(G128), .ZN(n1171) );
XOR2_X1 U884 ( .A(n1174), .B(n1175), .Z(n1169) );
XNOR2_X1 U885 ( .A(n1176), .B(G110), .ZN(n1175) );
INV_X1 U886 ( .A(G119), .ZN(n1176) );
NAND3_X1 U887 ( .A1(G234), .A2(n1044), .A3(G221), .ZN(n1165) );
NAND3_X1 U888 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1151) );
OR2_X1 U889 ( .A1(G472), .A2(KEYINPUT43), .ZN(n1179) );
NAND3_X1 U890 ( .A1(KEYINPUT43), .A2(G472), .A3(n1034), .ZN(n1178) );
NAND2_X1 U891 ( .A1(n1180), .A2(n1181), .ZN(n1177) );
NAND2_X1 U892 ( .A1(KEYINPUT43), .A2(n1182), .ZN(n1181) );
XOR2_X1 U893 ( .A(KEYINPUT10), .B(G472), .Z(n1182) );
INV_X1 U894 ( .A(n1034), .ZN(n1180) );
NAND2_X1 U895 ( .A1(n1183), .A2(n1113), .ZN(n1034) );
XNOR2_X1 U896 ( .A(n1184), .B(n1087), .ZN(n1183) );
XOR2_X1 U897 ( .A(n1185), .B(n1146), .Z(n1087) );
NAND2_X1 U898 ( .A1(n1186), .A2(G210), .ZN(n1185) );
NAND2_X1 U899 ( .A1(n1187), .A2(KEYINPUT35), .ZN(n1184) );
XOR2_X1 U900 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U901 ( .A(n1099), .B(n1097), .Z(n1189) );
XNOR2_X1 U902 ( .A(KEYINPUT27), .B(n1190), .ZN(n1099) );
XNOR2_X1 U903 ( .A(n1094), .B(KEYINPUT48), .ZN(n1188) );
XNOR2_X1 U904 ( .A(n1191), .B(n1192), .ZN(n1094) );
XOR2_X1 U905 ( .A(KEYINPUT45), .B(n1193), .Z(n1192) );
NOR2_X1 U906 ( .A1(KEYINPUT37), .A2(n1158), .ZN(n1193) );
AND3_X1 U907 ( .A1(n1126), .A2(n1156), .A3(n1012), .ZN(n1121) );
NOR2_X1 U908 ( .A1(n1015), .A2(n1016), .ZN(n1012) );
AND2_X1 U909 ( .A1(G221), .A2(n1163), .ZN(n1016) );
NAND2_X1 U910 ( .A1(G234), .A2(n1113), .ZN(n1163) );
INV_X1 U911 ( .A(n1160), .ZN(n1015) );
XNOR2_X1 U912 ( .A(n1194), .B(G469), .ZN(n1160) );
NAND2_X1 U913 ( .A1(n1195), .A2(n1113), .ZN(n1194) );
XOR2_X1 U914 ( .A(n1105), .B(n1196), .Z(n1195) );
XOR2_X1 U915 ( .A(n1197), .B(KEYINPUT8), .Z(n1196) );
NAND2_X1 U916 ( .A1(KEYINPUT38), .A2(n1106), .ZN(n1197) );
XOR2_X1 U917 ( .A(n1198), .B(n1199), .Z(n1105) );
XNOR2_X1 U918 ( .A(n1146), .B(n1200), .ZN(n1199) );
XOR2_X1 U919 ( .A(KEYINPUT27), .B(G110), .Z(n1200) );
XOR2_X1 U920 ( .A(n1055), .B(n1201), .Z(n1198) );
XOR2_X1 U921 ( .A(n1202), .B(n1203), .Z(n1201) );
NAND2_X1 U922 ( .A1(KEYINPUT59), .A2(n1204), .ZN(n1203) );
NAND2_X1 U923 ( .A1(n1205), .A2(n1044), .ZN(n1202) );
XOR2_X1 U924 ( .A(KEYINPUT51), .B(G227), .Z(n1205) );
XOR2_X1 U925 ( .A(n1206), .B(n1207), .Z(n1055) );
XNOR2_X1 U926 ( .A(n1173), .B(n1208), .ZN(n1207) );
NOR2_X1 U927 ( .A1(KEYINPUT22), .A2(n1209), .ZN(n1208) );
XNOR2_X1 U928 ( .A(n1210), .B(n1190), .ZN(n1206) );
XNOR2_X1 U929 ( .A(n1211), .B(n1212), .ZN(n1190) );
XOR2_X1 U930 ( .A(KEYINPUT61), .B(G137), .Z(n1212) );
XNOR2_X1 U931 ( .A(G131), .B(G134), .ZN(n1211) );
NAND2_X1 U932 ( .A1(n1213), .A2(n987), .ZN(n1156) );
NAND3_X1 U933 ( .A1(n1149), .A2(n1044), .A3(G952), .ZN(n987) );
XOR2_X1 U934 ( .A(n1214), .B(KEYINPUT14), .Z(n1213) );
NAND4_X1 U935 ( .A1(G953), .A2(G902), .A3(n1149), .A4(n1066), .ZN(n1214) );
INV_X1 U936 ( .A(G898), .ZN(n1066) );
NAND2_X1 U937 ( .A1(G237), .A2(G234), .ZN(n1149) );
NOR2_X1 U938 ( .A1(n1008), .A2(n1000), .ZN(n1126) );
INV_X1 U939 ( .A(n1006), .ZN(n1000) );
NAND2_X1 U940 ( .A1(G214), .A2(n1215), .ZN(n1006) );
XNOR2_X1 U941 ( .A(n1031), .B(n1216), .ZN(n1008) );
NOR2_X1 U942 ( .A1(n1033), .A2(KEYINPUT30), .ZN(n1216) );
AND2_X1 U943 ( .A1(G210), .A2(n1215), .ZN(n1033) );
NAND2_X1 U944 ( .A1(n1217), .A2(n1113), .ZN(n1215) );
INV_X1 U945 ( .A(G237), .ZN(n1217) );
NAND2_X1 U946 ( .A1(n1218), .A2(n1113), .ZN(n1031) );
XNOR2_X1 U947 ( .A(n1219), .B(n1071), .ZN(n1218) );
XOR2_X1 U948 ( .A(n1220), .B(n1221), .Z(n1071) );
XOR2_X1 U949 ( .A(n1222), .B(n1191), .Z(n1221) );
XNOR2_X1 U950 ( .A(G119), .B(n1223), .ZN(n1191) );
NAND2_X1 U951 ( .A1(n1224), .A2(n1225), .ZN(n1222) );
OR2_X1 U952 ( .A1(n1146), .A2(n1204), .ZN(n1225) );
XOR2_X1 U953 ( .A(n1226), .B(KEYINPUT41), .Z(n1224) );
NAND2_X1 U954 ( .A1(n1204), .A2(n1146), .ZN(n1226) );
INV_X1 U955 ( .A(G101), .ZN(n1146) );
XNOR2_X1 U956 ( .A(G104), .B(G107), .ZN(n1204) );
XNOR2_X1 U957 ( .A(n1227), .B(n1158), .ZN(n1220) );
INV_X1 U958 ( .A(G113), .ZN(n1158) );
NAND3_X1 U959 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1227) );
NAND2_X1 U960 ( .A1(G110), .A2(n1231), .ZN(n1230) );
INV_X1 U961 ( .A(KEYINPUT0), .ZN(n1231) );
NAND3_X1 U962 ( .A1(KEYINPUT0), .A2(n1232), .A3(n1233), .ZN(n1229) );
OR2_X1 U963 ( .A1(n1233), .A2(n1232), .ZN(n1228) );
NOR2_X1 U964 ( .A1(G110), .A2(KEYINPUT54), .ZN(n1232) );
NAND2_X1 U965 ( .A1(n1234), .A2(n1235), .ZN(n1219) );
NAND2_X1 U966 ( .A1(n1112), .A2(n1061), .ZN(n1235) );
INV_X1 U967 ( .A(G125), .ZN(n1061) );
NAND2_X1 U968 ( .A1(n1236), .A2(G125), .ZN(n1234) );
XNOR2_X1 U969 ( .A(n1112), .B(KEYINPUT18), .ZN(n1236) );
XNOR2_X1 U970 ( .A(n1097), .B(n1237), .ZN(n1112) );
NOR2_X1 U971 ( .A1(G953), .A2(n1065), .ZN(n1237) );
INV_X1 U972 ( .A(G224), .ZN(n1065) );
XOR2_X1 U973 ( .A(n1238), .B(n1239), .Z(n1097) );
XNOR2_X1 U974 ( .A(KEYINPUT33), .B(n1173), .ZN(n1239) );
XNOR2_X1 U975 ( .A(G143), .B(n1210), .ZN(n1238) );
XOR2_X1 U976 ( .A(G128), .B(KEYINPUT53), .Z(n1210) );
INV_X1 U977 ( .A(n992), .ZN(n1145) );
NAND2_X1 U978 ( .A1(n1161), .A2(n1157), .ZN(n992) );
XNOR2_X1 U979 ( .A(KEYINPUT19), .B(n1143), .ZN(n1157) );
NAND2_X1 U980 ( .A1(n1240), .A2(n1241), .ZN(n1143) );
NAND2_X1 U981 ( .A1(G475), .A2(n1040), .ZN(n1241) );
INV_X1 U982 ( .A(n1038), .ZN(n1240) );
NOR2_X1 U983 ( .A1(n1040), .A2(G475), .ZN(n1038) );
NAND2_X1 U984 ( .A1(n1083), .A2(n1113), .ZN(n1040) );
XNOR2_X1 U985 ( .A(n1242), .B(n1243), .ZN(n1083) );
XOR2_X1 U986 ( .A(n1244), .B(n1245), .Z(n1243) );
XOR2_X1 U987 ( .A(n1246), .B(n1247), .Z(n1245) );
NAND2_X1 U988 ( .A1(KEYINPUT29), .A2(n1248), .ZN(n1247) );
INV_X1 U989 ( .A(G131), .ZN(n1248) );
NAND3_X1 U990 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1246) );
XNOR2_X1 U991 ( .A(KEYINPUT15), .B(KEYINPUT13), .ZN(n1251) );
NAND2_X1 U992 ( .A1(n1252), .A2(n1253), .ZN(n1250) );
NAND2_X1 U993 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U994 ( .A1(G122), .A2(n1256), .ZN(n1255) );
INV_X1 U995 ( .A(KEYINPUT34), .ZN(n1254) );
NAND2_X1 U996 ( .A1(n1257), .A2(n1233), .ZN(n1249) );
NAND2_X1 U997 ( .A1(n1256), .A2(n1258), .ZN(n1257) );
OR2_X1 U998 ( .A1(n1252), .A2(KEYINPUT34), .ZN(n1258) );
XNOR2_X1 U999 ( .A(G113), .B(KEYINPUT1), .ZN(n1252) );
INV_X1 U1000 ( .A(KEYINPUT31), .ZN(n1256) );
AND2_X1 U1001 ( .A1(G214), .A2(n1186), .ZN(n1244) );
NOR2_X1 U1002 ( .A1(G953), .A2(G237), .ZN(n1186) );
XOR2_X1 U1003 ( .A(n1259), .B(n1260), .Z(n1242) );
XNOR2_X1 U1004 ( .A(n1209), .B(G104), .ZN(n1260) );
INV_X1 U1005 ( .A(G143), .ZN(n1209) );
NAND3_X1 U1006 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1259) );
NAND2_X1 U1007 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
INV_X1 U1008 ( .A(KEYINPUT25), .ZN(n1265) );
NAND3_X1 U1009 ( .A1(KEYINPUT25), .A2(n1266), .A3(n1173), .ZN(n1262) );
OR2_X1 U1010 ( .A1(n1173), .A2(n1266), .ZN(n1261) );
NOR2_X1 U1011 ( .A1(KEYINPUT60), .A2(n1264), .ZN(n1266) );
XNOR2_X1 U1012 ( .A(n1174), .B(KEYINPUT20), .ZN(n1264) );
NAND2_X1 U1013 ( .A1(n1267), .A2(n1268), .ZN(n1174) );
NAND2_X1 U1014 ( .A1(G125), .A2(n1106), .ZN(n1268) );
INV_X1 U1015 ( .A(n1058), .ZN(n1267) );
NOR2_X1 U1016 ( .A1(n1106), .A2(G125), .ZN(n1058) );
INV_X1 U1017 ( .A(G140), .ZN(n1106) );
INV_X1 U1018 ( .A(G146), .ZN(n1173) );
XNOR2_X1 U1019 ( .A(n1036), .B(KEYINPUT16), .ZN(n1161) );
XNOR2_X1 U1020 ( .A(n1269), .B(G478), .ZN(n1036) );
NAND2_X1 U1021 ( .A1(n1270), .A2(n1113), .ZN(n1269) );
INV_X1 U1022 ( .A(G902), .ZN(n1113) );
XOR2_X1 U1023 ( .A(n1080), .B(KEYINPUT42), .Z(n1270) );
XOR2_X1 U1024 ( .A(n1271), .B(n1272), .Z(n1080) );
XOR2_X1 U1025 ( .A(n1273), .B(n1274), .Z(n1272) );
XOR2_X1 U1026 ( .A(G134), .B(G107), .Z(n1274) );
NOR2_X1 U1027 ( .A1(KEYINPUT9), .A2(n1275), .ZN(n1273) );
XNOR2_X1 U1028 ( .A(G128), .B(G143), .ZN(n1275) );
XNOR2_X1 U1029 ( .A(n1276), .B(n1277), .ZN(n1271) );
NAND2_X1 U1030 ( .A1(KEYINPUT21), .A2(n1278), .ZN(n1277) );
NAND3_X1 U1031 ( .A1(G234), .A2(n1044), .A3(G217), .ZN(n1278) );
INV_X1 U1032 ( .A(G953), .ZN(n1044) );
NAND2_X1 U1033 ( .A1(KEYINPUT7), .A2(n1279), .ZN(n1276) );
XNOR2_X1 U1034 ( .A(n1233), .B(n1223), .ZN(n1279) );
XOR2_X1 U1035 ( .A(G116), .B(KEYINPUT49), .Z(n1223) );
INV_X1 U1036 ( .A(G122), .ZN(n1233) );
endmodule


