//Key = 1101010010001010101000011100101110001011111001001100001110001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332;

NAND2_X1 U734 ( .A1(n1015), .A2(n1016), .ZN(G9) );
OR2_X1 U735 ( .A1(n1017), .A2(G107), .ZN(n1016) );
XOR2_X1 U736 ( .A(n1018), .B(KEYINPUT27), .Z(n1015) );
NAND2_X1 U737 ( .A1(n1019), .A2(n1017), .ZN(n1018) );
NAND2_X1 U738 ( .A1(n1020), .A2(n1021), .ZN(n1017) );
XOR2_X1 U739 ( .A(KEYINPUT2), .B(n1022), .Z(n1021) );
NOR2_X1 U740 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
XOR2_X1 U741 ( .A(KEYINPUT22), .B(G107), .Z(n1019) );
NOR2_X1 U742 ( .A1(n1025), .A2(n1026), .ZN(G75) );
NOR4_X1 U743 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
NOR2_X1 U744 ( .A1(n1031), .A2(n1032), .ZN(n1028) );
NOR2_X1 U745 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR3_X1 U746 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NOR3_X1 U747 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1036) );
NOR3_X1 U748 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NOR3_X1 U749 ( .A1(n1044), .A2(n1045), .A3(n1042), .ZN(n1039) );
NOR2_X1 U750 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR4_X1 U751 ( .A1(n1044), .A2(n1048), .A3(n1042), .A4(n1043), .ZN(n1033) );
INV_X1 U752 ( .A(n1049), .ZN(n1043) );
NOR2_X1 U753 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR2_X1 U754 ( .A1(n1052), .A2(n1035), .ZN(n1051) );
NOR2_X1 U755 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR2_X1 U756 ( .A1(n1055), .A2(n1037), .ZN(n1050) );
INV_X1 U757 ( .A(n1056), .ZN(n1037) );
NOR2_X1 U758 ( .A1(n1057), .A2(n1020), .ZN(n1055) );
NOR2_X1 U759 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR3_X1 U760 ( .A1(n1030), .A2(G952), .A3(n1027), .ZN(n1025) );
AND4_X1 U761 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1027) );
NOR3_X1 U762 ( .A1(n1064), .A2(n1065), .A3(n1044), .ZN(n1063) );
NAND3_X1 U763 ( .A1(n1058), .A2(n1066), .A3(n1067), .ZN(n1064) );
NOR3_X1 U764 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1062) );
XNOR2_X1 U765 ( .A(n1071), .B(n1072), .ZN(n1069) );
NOR2_X1 U766 ( .A1(n1073), .A2(KEYINPUT50), .ZN(n1072) );
XNOR2_X1 U767 ( .A(n1074), .B(n1075), .ZN(n1068) );
XNOR2_X1 U768 ( .A(G469), .B(KEYINPUT15), .ZN(n1075) );
XNOR2_X1 U769 ( .A(n1076), .B(KEYINPUT46), .ZN(n1061) );
XNOR2_X1 U770 ( .A(n1077), .B(G475), .ZN(n1060) );
XOR2_X1 U771 ( .A(n1078), .B(n1079), .Z(G72) );
XOR2_X1 U772 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U773 ( .A1(G953), .A2(n1082), .ZN(n1081) );
XOR2_X1 U774 ( .A(KEYINPUT33), .B(n1083), .Z(n1082) );
NOR2_X1 U775 ( .A1(n1084), .A2(n1085), .ZN(n1080) );
NOR2_X1 U776 ( .A1(n1086), .A2(KEYINPUT31), .ZN(n1085) );
NOR2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR3_X1 U778 ( .A1(n1088), .A2(KEYINPUT17), .A3(n1087), .ZN(n1084) );
AND2_X1 U779 ( .A1(G900), .A2(G227), .ZN(n1087) );
NAND2_X1 U780 ( .A1(n1089), .A2(n1090), .ZN(n1078) );
NAND2_X1 U781 ( .A1(n1091), .A2(G953), .ZN(n1090) );
XOR2_X1 U782 ( .A(n1092), .B(n1093), .Z(n1089) );
XOR2_X1 U783 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U784 ( .A1(KEYINPUT16), .A2(n1096), .ZN(n1095) );
NAND3_X1 U785 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1094) );
OR2_X1 U786 ( .A1(n1100), .A2(KEYINPUT28), .ZN(n1099) );
NAND3_X1 U787 ( .A1(KEYINPUT28), .A2(n1100), .A3(G140), .ZN(n1098) );
NAND2_X1 U788 ( .A1(n1101), .A2(n1102), .ZN(n1097) );
NAND2_X1 U789 ( .A1(n1103), .A2(KEYINPUT28), .ZN(n1101) );
XNOR2_X1 U790 ( .A(G125), .B(KEYINPUT29), .ZN(n1103) );
XNOR2_X1 U791 ( .A(n1104), .B(n1105), .ZN(n1092) );
XOR2_X1 U792 ( .A(n1106), .B(n1107), .Z(G69) );
XOR2_X1 U793 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U794 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
INV_X1 U795 ( .A(n1112), .ZN(n1111) );
XOR2_X1 U796 ( .A(n1113), .B(n1114), .Z(n1110) );
XOR2_X1 U797 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U798 ( .A1(n1088), .A2(n1117), .ZN(n1108) );
NAND2_X1 U799 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XNOR2_X1 U800 ( .A(n1120), .B(KEYINPUT1), .ZN(n1118) );
NOR2_X1 U801 ( .A1(n1121), .A2(n1088), .ZN(n1106) );
AND2_X1 U802 ( .A1(G224), .A2(G898), .ZN(n1121) );
NOR2_X1 U803 ( .A1(n1122), .A2(n1123), .ZN(G66) );
NOR3_X1 U804 ( .A1(n1071), .A2(n1124), .A3(n1125), .ZN(n1123) );
AND3_X1 U805 ( .A1(n1126), .A2(n1073), .A3(n1127), .ZN(n1125) );
INV_X1 U806 ( .A(n1128), .ZN(n1073) );
NOR2_X1 U807 ( .A1(n1129), .A2(n1126), .ZN(n1124) );
NOR2_X1 U808 ( .A1(n1130), .A2(n1128), .ZN(n1129) );
NOR2_X1 U809 ( .A1(n1122), .A2(n1131), .ZN(G63) );
XNOR2_X1 U810 ( .A(n1132), .B(n1133), .ZN(n1131) );
NAND2_X1 U811 ( .A1(n1127), .A2(G478), .ZN(n1132) );
NOR2_X1 U812 ( .A1(n1122), .A2(n1134), .ZN(G60) );
NOR3_X1 U813 ( .A1(n1077), .A2(n1135), .A3(n1136), .ZN(n1134) );
AND3_X1 U814 ( .A1(n1137), .A2(G475), .A3(n1127), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
AND2_X1 U816 ( .A1(n1029), .A2(G475), .ZN(n1138) );
XNOR2_X1 U817 ( .A(n1139), .B(n1140), .ZN(G6) );
NOR3_X1 U818 ( .A1(n1141), .A2(n1023), .A3(n1142), .ZN(n1140) );
XNOR2_X1 U819 ( .A(KEYINPUT42), .B(n1143), .ZN(n1141) );
NOR2_X1 U820 ( .A1(n1122), .A2(n1144), .ZN(G57) );
XOR2_X1 U821 ( .A(n1145), .B(n1146), .Z(n1144) );
XNOR2_X1 U822 ( .A(n1147), .B(n1148), .ZN(n1146) );
XOR2_X1 U823 ( .A(n1149), .B(n1150), .Z(n1145) );
NAND2_X1 U824 ( .A1(n1127), .A2(G472), .ZN(n1149) );
NOR2_X1 U825 ( .A1(n1122), .A2(n1151), .ZN(G54) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U827 ( .A1(n1127), .A2(G469), .ZN(n1153) );
NAND2_X1 U828 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NAND2_X1 U829 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
OR2_X1 U830 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U831 ( .A(KEYINPUT12), .B(n1160), .Z(n1154) );
NOR3_X1 U832 ( .A1(n1158), .A2(n1159), .A3(n1156), .ZN(n1160) );
XOR2_X1 U833 ( .A(n1161), .B(n1162), .Z(n1156) );
XNOR2_X1 U834 ( .A(KEYINPUT18), .B(n1163), .ZN(n1162) );
NAND2_X1 U835 ( .A1(KEYINPUT14), .A2(n1164), .ZN(n1161) );
AND2_X1 U836 ( .A1(n1165), .A2(n1166), .ZN(n1159) );
XNOR2_X1 U837 ( .A(n1167), .B(KEYINPUT7), .ZN(n1158) );
OR2_X1 U838 ( .A1(n1165), .A2(n1166), .ZN(n1167) );
XNOR2_X1 U839 ( .A(n1168), .B(n1116), .ZN(n1165) );
XOR2_X1 U840 ( .A(n1169), .B(KEYINPUT13), .Z(n1168) );
NAND2_X1 U841 ( .A1(KEYINPUT0), .A2(n1104), .ZN(n1169) );
NOR2_X1 U842 ( .A1(n1122), .A2(n1170), .ZN(G51) );
XOR2_X1 U843 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR3_X1 U844 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1172) );
AND3_X1 U845 ( .A1(KEYINPUT40), .A2(n1176), .A3(n1177), .ZN(n1175) );
NOR2_X1 U846 ( .A1(KEYINPUT40), .A2(n1177), .ZN(n1174) );
XOR2_X1 U847 ( .A(n1178), .B(KEYINPUT30), .Z(n1171) );
NAND2_X1 U848 ( .A1(n1127), .A2(n1179), .ZN(n1178) );
XNOR2_X1 U849 ( .A(KEYINPUT4), .B(n1180), .ZN(n1179) );
NOR2_X1 U850 ( .A1(n1181), .A2(n1130), .ZN(n1127) );
INV_X1 U851 ( .A(n1029), .ZN(n1130) );
NAND3_X1 U852 ( .A1(n1083), .A2(n1119), .A3(n1120), .ZN(n1029) );
AND4_X1 U853 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1120) );
NAND2_X1 U854 ( .A1(n1020), .A2(n1186), .ZN(n1119) );
NAND3_X1 U855 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1186) );
NAND2_X1 U856 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND2_X1 U857 ( .A1(n1142), .A2(n1024), .ZN(n1191) );
INV_X1 U858 ( .A(n1046), .ZN(n1024) );
INV_X1 U859 ( .A(n1023), .ZN(n1190) );
NAND4_X1 U860 ( .A1(n1042), .A2(n1056), .A3(n1192), .A4(n1041), .ZN(n1023) );
NAND3_X1 U861 ( .A1(n1054), .A2(n1192), .A3(n1038), .ZN(n1187) );
AND4_X1 U862 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1083) );
AND4_X1 U863 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1196) );
AND2_X1 U864 ( .A1(n1201), .A2(n1202), .ZN(n1195) );
NOR2_X1 U865 ( .A1(n1088), .A2(G952), .ZN(n1122) );
NAND3_X1 U866 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(G48) );
OR2_X1 U867 ( .A1(n1206), .A2(n1202), .ZN(n1205) );
NAND3_X1 U868 ( .A1(n1202), .A2(n1206), .A3(G146), .ZN(n1204) );
NAND2_X1 U869 ( .A1(n1207), .A2(n1208), .ZN(n1203) );
NAND2_X1 U870 ( .A1(n1209), .A2(n1206), .ZN(n1207) );
INV_X1 U871 ( .A(KEYINPUT53), .ZN(n1206) );
XNOR2_X1 U872 ( .A(KEYINPUT3), .B(n1202), .ZN(n1209) );
NAND3_X1 U873 ( .A1(n1047), .A2(n1020), .A3(n1210), .ZN(n1202) );
NAND2_X1 U874 ( .A1(n1211), .A2(n1212), .ZN(G45) );
NAND2_X1 U875 ( .A1(G143), .A2(n1201), .ZN(n1212) );
XOR2_X1 U876 ( .A(n1213), .B(KEYINPUT52), .Z(n1211) );
OR2_X1 U877 ( .A1(n1201), .A2(G143), .ZN(n1213) );
NAND4_X1 U878 ( .A1(n1214), .A2(n1215), .A3(n1020), .A4(n1216), .ZN(n1201) );
AND2_X1 U879 ( .A1(n1053), .A2(n1217), .ZN(n1216) );
XNOR2_X1 U880 ( .A(G140), .B(n1193), .ZN(G42) );
NAND2_X1 U881 ( .A1(n1218), .A2(n1054), .ZN(n1193) );
XNOR2_X1 U882 ( .A(G137), .B(n1219), .ZN(G39) );
NAND2_X1 U883 ( .A1(KEYINPUT23), .A2(n1220), .ZN(n1219) );
INV_X1 U884 ( .A(n1194), .ZN(n1220) );
NAND3_X1 U885 ( .A1(n1210), .A2(n1049), .A3(n1221), .ZN(n1194) );
XNOR2_X1 U886 ( .A(n1222), .B(n1200), .ZN(G36) );
NAND4_X1 U887 ( .A1(n1221), .A2(n1217), .A3(n1053), .A4(n1046), .ZN(n1200) );
NAND2_X1 U888 ( .A1(KEYINPUT54), .A2(n1096), .ZN(n1222) );
XNOR2_X1 U889 ( .A(G131), .B(n1199), .ZN(G33) );
NAND2_X1 U890 ( .A1(n1218), .A2(n1053), .ZN(n1199) );
NOR3_X1 U891 ( .A1(n1223), .A2(n1142), .A3(n1035), .ZN(n1218) );
INV_X1 U892 ( .A(n1221), .ZN(n1035) );
NOR2_X1 U893 ( .A1(n1059), .A2(n1224), .ZN(n1221) );
XOR2_X1 U894 ( .A(KEYINPUT41), .B(n1058), .Z(n1224) );
XNOR2_X1 U895 ( .A(G128), .B(n1198), .ZN(G30) );
NAND3_X1 U896 ( .A1(n1020), .A2(n1046), .A3(n1210), .ZN(n1198) );
AND3_X1 U897 ( .A1(n1070), .A2(n1225), .A3(n1217), .ZN(n1210) );
INV_X1 U898 ( .A(n1223), .ZN(n1217) );
NAND2_X1 U899 ( .A1(n1226), .A2(n1042), .ZN(n1223) );
INV_X1 U900 ( .A(n1143), .ZN(n1020) );
XOR2_X1 U901 ( .A(G101), .B(n1227), .Z(G3) );
NOR2_X1 U902 ( .A1(n1143), .A2(n1228), .ZN(n1227) );
XNOR2_X1 U903 ( .A(KEYINPUT49), .B(n1188), .ZN(n1228) );
NAND3_X1 U904 ( .A1(n1053), .A2(n1192), .A3(n1038), .ZN(n1188) );
XNOR2_X1 U905 ( .A(G125), .B(n1197), .ZN(G27) );
NAND3_X1 U906 ( .A1(n1054), .A2(n1226), .A3(n1229), .ZN(n1197) );
NOR3_X1 U907 ( .A1(n1142), .A2(n1042), .A3(n1143), .ZN(n1229) );
AND2_X1 U908 ( .A1(n1041), .A2(n1230), .ZN(n1226) );
NAND2_X1 U909 ( .A1(n1231), .A2(n1032), .ZN(n1230) );
NAND4_X1 U910 ( .A1(n1091), .A2(G902), .A3(G953), .A4(n1232), .ZN(n1231) );
XNOR2_X1 U911 ( .A(G900), .B(KEYINPUT51), .ZN(n1091) );
XNOR2_X1 U912 ( .A(G122), .B(n1182), .ZN(G24) );
NAND4_X1 U913 ( .A1(n1233), .A2(n1056), .A3(n1214), .A4(n1215), .ZN(n1182) );
NOR2_X1 U914 ( .A1(n1225), .A2(n1070), .ZN(n1056) );
NAND2_X1 U915 ( .A1(n1234), .A2(n1235), .ZN(G21) );
OR2_X1 U916 ( .A1(n1183), .A2(G119), .ZN(n1235) );
XOR2_X1 U917 ( .A(n1236), .B(KEYINPUT57), .Z(n1234) );
NAND2_X1 U918 ( .A1(G119), .A2(n1183), .ZN(n1236) );
NAND4_X1 U919 ( .A1(n1233), .A2(n1049), .A3(n1070), .A4(n1225), .ZN(n1183) );
XNOR2_X1 U920 ( .A(G116), .B(n1184), .ZN(G18) );
NAND3_X1 U921 ( .A1(n1053), .A2(n1046), .A3(n1233), .ZN(n1184) );
NAND2_X1 U922 ( .A1(n1237), .A2(n1238), .ZN(G15) );
NAND2_X1 U923 ( .A1(G113), .A2(n1185), .ZN(n1238) );
XOR2_X1 U924 ( .A(KEYINPUT5), .B(n1239), .Z(n1237) );
NOR2_X1 U925 ( .A1(G113), .A2(n1185), .ZN(n1239) );
NAND3_X1 U926 ( .A1(n1047), .A2(n1053), .A3(n1233), .ZN(n1185) );
NOR4_X1 U927 ( .A1(n1143), .A2(n1042), .A3(n1240), .A4(n1044), .ZN(n1233) );
INV_X1 U928 ( .A(n1041), .ZN(n1044) );
NOR2_X1 U929 ( .A1(n1225), .A2(n1241), .ZN(n1053) );
INV_X1 U930 ( .A(n1142), .ZN(n1047) );
XNOR2_X1 U931 ( .A(G110), .B(n1242), .ZN(G12) );
NAND3_X1 U932 ( .A1(n1243), .A2(n1038), .A3(n1244), .ZN(n1242) );
NOR3_X1 U933 ( .A1(n1143), .A2(KEYINPUT9), .A3(n1240), .ZN(n1244) );
INV_X1 U934 ( .A(n1192), .ZN(n1240) );
NAND2_X1 U935 ( .A1(n1032), .A2(n1245), .ZN(n1192) );
NAND3_X1 U936 ( .A1(n1112), .A2(n1232), .A3(G902), .ZN(n1245) );
NOR2_X1 U937 ( .A1(n1088), .A2(G898), .ZN(n1112) );
NAND3_X1 U938 ( .A1(n1246), .A2(n1232), .A3(G952), .ZN(n1032) );
NAND2_X1 U939 ( .A1(G237), .A2(G234), .ZN(n1232) );
INV_X1 U940 ( .A(n1030), .ZN(n1246) );
XOR2_X1 U941 ( .A(G953), .B(KEYINPUT59), .Z(n1030) );
NAND2_X1 U942 ( .A1(n1058), .A2(n1059), .ZN(n1143) );
NAND2_X1 U943 ( .A1(n1247), .A2(n1066), .ZN(n1059) );
NAND3_X1 U944 ( .A1(n1180), .A2(n1181), .A3(n1248), .ZN(n1066) );
XNOR2_X1 U945 ( .A(KEYINPUT39), .B(n1067), .ZN(n1247) );
NAND2_X1 U946 ( .A1(n1249), .A2(n1250), .ZN(n1067) );
NAND2_X1 U947 ( .A1(n1248), .A2(n1181), .ZN(n1250) );
NAND2_X1 U948 ( .A1(n1251), .A2(n1252), .ZN(n1248) );
NAND2_X1 U949 ( .A1(n1177), .A2(n1176), .ZN(n1252) );
INV_X1 U950 ( .A(n1173), .ZN(n1251) );
NOR2_X1 U951 ( .A1(n1176), .A2(n1177), .ZN(n1173) );
XNOR2_X1 U952 ( .A(n1253), .B(n1254), .ZN(n1177) );
XOR2_X1 U953 ( .A(n1255), .B(n1113), .Z(n1254) );
XNOR2_X1 U954 ( .A(n1256), .B(G113), .ZN(n1113) );
XNOR2_X1 U955 ( .A(n1257), .B(n1100), .ZN(n1253) );
NAND2_X1 U956 ( .A1(KEYINPUT8), .A2(n1115), .ZN(n1257) );
XNOR2_X1 U957 ( .A(G110), .B(n1258), .ZN(n1115) );
NAND2_X1 U958 ( .A1(G224), .A2(n1088), .ZN(n1176) );
INV_X1 U959 ( .A(n1180), .ZN(n1249) );
NAND2_X1 U960 ( .A1(G210), .A2(n1259), .ZN(n1180) );
NAND2_X1 U961 ( .A1(G214), .A2(n1259), .ZN(n1058) );
NAND2_X1 U962 ( .A1(n1260), .A2(n1181), .ZN(n1259) );
INV_X1 U963 ( .A(G237), .ZN(n1260) );
AND3_X1 U964 ( .A1(n1049), .A2(n1041), .A3(n1042), .ZN(n1038) );
XNOR2_X1 U965 ( .A(G469), .B(n1261), .ZN(n1042) );
NOR2_X1 U966 ( .A1(n1074), .A2(KEYINPUT43), .ZN(n1261) );
AND2_X1 U967 ( .A1(n1262), .A2(n1181), .ZN(n1074) );
XOR2_X1 U968 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U969 ( .A(n1255), .B(n1164), .ZN(n1264) );
XNOR2_X1 U970 ( .A(G110), .B(n1102), .ZN(n1164) );
INV_X1 U971 ( .A(G140), .ZN(n1102) );
XNOR2_X1 U972 ( .A(n1116), .B(n1104), .ZN(n1255) );
XOR2_X1 U973 ( .A(G101), .B(n1265), .Z(n1116) );
XNOR2_X1 U974 ( .A(G107), .B(n1139), .ZN(n1265) );
XOR2_X1 U975 ( .A(n1266), .B(n1267), .Z(n1263) );
XNOR2_X1 U976 ( .A(KEYINPUT13), .B(n1163), .ZN(n1267) );
NAND2_X1 U977 ( .A1(G227), .A2(n1268), .ZN(n1163) );
XNOR2_X1 U978 ( .A(KEYINPUT24), .B(n1088), .ZN(n1268) );
NAND2_X1 U979 ( .A1(KEYINPUT61), .A2(n1269), .ZN(n1266) );
NAND2_X1 U980 ( .A1(G221), .A2(n1270), .ZN(n1041) );
NAND2_X1 U981 ( .A1(n1271), .A2(n1272), .ZN(n1049) );
OR2_X1 U982 ( .A1(n1142), .A2(KEYINPUT62), .ZN(n1272) );
NAND2_X1 U983 ( .A1(n1273), .A2(n1214), .ZN(n1142) );
XNOR2_X1 U984 ( .A(KEYINPUT10), .B(n1215), .ZN(n1273) );
NAND2_X1 U985 ( .A1(KEYINPUT62), .A2(n1274), .ZN(n1271) );
NAND2_X1 U986 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
OR3_X1 U987 ( .A1(n1215), .A2(n1214), .A3(KEYINPUT10), .ZN(n1276) );
INV_X1 U988 ( .A(n1277), .ZN(n1215) );
NAND2_X1 U989 ( .A1(KEYINPUT10), .A2(n1046), .ZN(n1275) );
NOR2_X1 U990 ( .A1(n1214), .A2(n1277), .ZN(n1046) );
NOR2_X1 U991 ( .A1(n1076), .A2(n1065), .ZN(n1277) );
NOR3_X1 U992 ( .A1(G478), .A2(G902), .A3(n1133), .ZN(n1065) );
AND2_X1 U993 ( .A1(G478), .A2(n1278), .ZN(n1076) );
OR2_X1 U994 ( .A1(n1133), .A2(G902), .ZN(n1278) );
XOR2_X1 U995 ( .A(n1279), .B(n1280), .Z(n1133) );
XOR2_X1 U996 ( .A(G107), .B(n1281), .Z(n1280) );
XNOR2_X1 U997 ( .A(n1096), .B(G116), .ZN(n1281) );
XOR2_X1 U998 ( .A(n1282), .B(n1258), .Z(n1279) );
XOR2_X1 U999 ( .A(n1283), .B(n1284), .Z(n1282) );
NAND3_X1 U1000 ( .A1(G217), .A2(n1088), .A3(G234), .ZN(n1283) );
XNOR2_X1 U1001 ( .A(n1285), .B(n1286), .ZN(n1214) );
XOR2_X1 U1002 ( .A(KEYINPUT25), .B(n1077), .Z(n1286) );
NOR2_X1 U1003 ( .A1(n1137), .A2(G902), .ZN(n1077) );
AND2_X1 U1004 ( .A1(n1287), .A2(n1288), .ZN(n1137) );
NAND2_X1 U1005 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XOR2_X1 U1006 ( .A(n1291), .B(KEYINPUT35), .Z(n1287) );
OR2_X1 U1007 ( .A1(n1290), .A2(n1289), .ZN(n1291) );
XOR2_X1 U1008 ( .A(n1292), .B(n1293), .Z(n1289) );
XNOR2_X1 U1009 ( .A(n1208), .B(n1294), .ZN(n1293) );
NOR2_X1 U1010 ( .A1(KEYINPUT47), .A2(n1295), .ZN(n1294) );
NAND2_X1 U1011 ( .A1(KEYINPUT55), .A2(n1296), .ZN(n1292) );
XOR2_X1 U1012 ( .A(n1297), .B(n1298), .Z(n1296) );
XNOR2_X1 U1013 ( .A(n1299), .B(n1300), .ZN(n1298) );
AND2_X1 U1014 ( .A1(G214), .A2(n1301), .ZN(n1300) );
INV_X1 U1015 ( .A(G131), .ZN(n1299) );
XOR2_X1 U1016 ( .A(KEYINPUT21), .B(G143), .Z(n1297) );
NAND3_X1 U1017 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1290) );
NAND2_X1 U1018 ( .A1(KEYINPUT20), .A2(n1305), .ZN(n1304) );
NAND3_X1 U1019 ( .A1(n1306), .A2(n1307), .A3(n1139), .ZN(n1303) );
INV_X1 U1020 ( .A(KEYINPUT20), .ZN(n1307) );
OR2_X1 U1021 ( .A1(n1139), .A2(n1306), .ZN(n1302) );
NOR2_X1 U1022 ( .A1(KEYINPUT6), .A2(n1305), .ZN(n1306) );
XNOR2_X1 U1023 ( .A(n1308), .B(n1258), .ZN(n1305) );
XOR2_X1 U1024 ( .A(G122), .B(KEYINPUT26), .Z(n1258) );
NAND2_X1 U1025 ( .A1(KEYINPUT56), .A2(n1309), .ZN(n1308) );
INV_X1 U1026 ( .A(G113), .ZN(n1309) );
INV_X1 U1027 ( .A(G104), .ZN(n1139) );
NAND2_X1 U1028 ( .A1(n1310), .A2(KEYINPUT36), .ZN(n1285) );
XNOR2_X1 U1029 ( .A(G475), .B(KEYINPUT58), .ZN(n1310) );
XNOR2_X1 U1030 ( .A(n1054), .B(KEYINPUT38), .ZN(n1243) );
AND2_X1 U1031 ( .A1(n1241), .A2(n1225), .ZN(n1054) );
XNOR2_X1 U1032 ( .A(n1071), .B(n1128), .ZN(n1225) );
NAND2_X1 U1033 ( .A1(G217), .A2(n1270), .ZN(n1128) );
NAND2_X1 U1034 ( .A1(G234), .A2(n1181), .ZN(n1270) );
NOR2_X1 U1035 ( .A1(n1126), .A2(G902), .ZN(n1071) );
XOR2_X1 U1036 ( .A(n1311), .B(n1312), .Z(n1126) );
XOR2_X1 U1037 ( .A(G119), .B(n1313), .Z(n1312) );
XOR2_X1 U1038 ( .A(G137), .B(G128), .Z(n1313) );
XOR2_X1 U1039 ( .A(n1314), .B(n1315), .Z(n1311) );
XNOR2_X1 U1040 ( .A(G110), .B(n1316), .ZN(n1315) );
NAND3_X1 U1041 ( .A1(G234), .A2(n1088), .A3(G221), .ZN(n1316) );
NAND3_X1 U1042 ( .A1(KEYINPUT32), .A2(n1317), .A3(n1318), .ZN(n1314) );
XOR2_X1 U1043 ( .A(n1319), .B(KEYINPUT19), .Z(n1318) );
NAND2_X1 U1044 ( .A1(G146), .A2(n1320), .ZN(n1319) );
NAND2_X1 U1045 ( .A1(n1295), .A2(n1208), .ZN(n1317) );
INV_X1 U1046 ( .A(G146), .ZN(n1208) );
INV_X1 U1047 ( .A(n1320), .ZN(n1295) );
XNOR2_X1 U1048 ( .A(G140), .B(n1100), .ZN(n1320) );
INV_X1 U1049 ( .A(G125), .ZN(n1100) );
INV_X1 U1050 ( .A(n1070), .ZN(n1241) );
XNOR2_X1 U1051 ( .A(n1321), .B(G472), .ZN(n1070) );
NAND2_X1 U1052 ( .A1(n1322), .A2(n1181), .ZN(n1321) );
INV_X1 U1053 ( .A(G902), .ZN(n1181) );
XOR2_X1 U1054 ( .A(n1150), .B(n1323), .Z(n1322) );
XNOR2_X1 U1055 ( .A(n1324), .B(n1325), .ZN(n1323) );
NOR2_X1 U1056 ( .A1(KEYINPUT44), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1057 ( .A(KEYINPUT11), .B(n1148), .Z(n1326) );
XNOR2_X1 U1058 ( .A(n1327), .B(G101), .ZN(n1148) );
NAND2_X1 U1059 ( .A1(n1301), .A2(G210), .ZN(n1327) );
AND2_X1 U1060 ( .A1(n1328), .A2(n1088), .ZN(n1301) );
INV_X1 U1061 ( .A(G953), .ZN(n1088) );
XNOR2_X1 U1062 ( .A(G237), .B(KEYINPUT63), .ZN(n1328) );
NAND2_X1 U1063 ( .A1(KEYINPUT48), .A2(n1147), .ZN(n1324) );
XNOR2_X1 U1064 ( .A(n1104), .B(KEYINPUT34), .ZN(n1147) );
XOR2_X1 U1065 ( .A(G146), .B(n1284), .Z(n1104) );
XOR2_X1 U1066 ( .A(G128), .B(G143), .Z(n1284) );
XNOR2_X1 U1067 ( .A(n1166), .B(n1329), .ZN(n1150) );
XNOR2_X1 U1068 ( .A(G113), .B(n1330), .ZN(n1329) );
NAND2_X1 U1069 ( .A1(KEYINPUT60), .A2(n1256), .ZN(n1330) );
XOR2_X1 U1070 ( .A(G116), .B(n1331), .Z(n1256) );
XOR2_X1 U1071 ( .A(KEYINPUT45), .B(G119), .Z(n1331) );
INV_X1 U1072 ( .A(n1269), .ZN(n1166) );
XOR2_X1 U1073 ( .A(n1105), .B(n1096), .Z(n1269) );
INV_X1 U1074 ( .A(G134), .ZN(n1096) );
XOR2_X1 U1075 ( .A(G131), .B(n1332), .Z(n1105) );
XOR2_X1 U1076 ( .A(KEYINPUT37), .B(G137), .Z(n1332) );
endmodule


