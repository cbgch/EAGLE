//Key = 0111100110001010110001110000110100001001111111001100000011111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311;

XNOR2_X1 U729 ( .A(G107), .B(n1000), .ZN(G9) );
NAND4_X1 U730 ( .A1(KEYINPUT56), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(n1000) );
NAND3_X1 U731 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(G75) );
NAND2_X1 U732 ( .A1(G952), .A2(n1007), .ZN(n1006) );
NAND4_X1 U733 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1007) );
NAND2_X1 U734 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND2_X1 U735 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND3_X1 U736 ( .A1(n1001), .A2(n1016), .A3(n1017), .ZN(n1015) );
NAND2_X1 U737 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NAND2_X1 U738 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U739 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND3_X1 U740 ( .A1(n1024), .A2(n1025), .A3(KEYINPUT8), .ZN(n1023) );
NAND3_X1 U741 ( .A1(n1026), .A2(n1027), .A3(n1024), .ZN(n1014) );
NAND2_X1 U742 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NAND3_X1 U743 ( .A1(n1001), .A2(n1025), .A3(n1017), .ZN(n1029) );
NAND3_X1 U744 ( .A1(n1030), .A2(n1027), .A3(n1031), .ZN(n1025) );
NAND2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
OR2_X1 U746 ( .A1(n1034), .A2(KEYINPUT8), .ZN(n1030) );
NAND2_X1 U747 ( .A1(n1020), .A2(n1035), .ZN(n1028) );
NAND2_X1 U748 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U749 ( .A1(n1001), .A2(n1038), .ZN(n1037) );
NAND2_X1 U750 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U751 ( .A1(n1017), .A2(n1041), .ZN(n1036) );
OR2_X1 U752 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
INV_X1 U753 ( .A(n1044), .ZN(n1012) );
XNOR2_X1 U754 ( .A(G953), .B(KEYINPUT55), .ZN(n1008) );
INV_X1 U755 ( .A(n1045), .ZN(n1005) );
NAND4_X1 U756 ( .A1(n1024), .A2(n1046), .A3(n1020), .A4(n1047), .ZN(n1004) );
NOR4_X1 U757 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
XNOR2_X1 U758 ( .A(n1052), .B(n1053), .ZN(n1050) );
NOR2_X1 U759 ( .A1(n1054), .A2(KEYINPUT53), .ZN(n1053) );
XNOR2_X1 U760 ( .A(G472), .B(n1055), .ZN(n1049) );
NOR2_X1 U761 ( .A1(n1056), .A2(KEYINPUT32), .ZN(n1055) );
INV_X1 U762 ( .A(n1057), .ZN(n1056) );
NAND2_X1 U763 ( .A1(n1058), .A2(n1059), .ZN(G72) );
NAND3_X1 U764 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
XNOR2_X1 U765 ( .A(KEYINPUT36), .B(n1063), .ZN(n1062) );
NAND2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1058) );
NAND2_X1 U767 ( .A1(n1060), .A2(n1061), .ZN(n1065) );
XOR2_X1 U768 ( .A(n1066), .B(n1067), .Z(n1064) );
XOR2_X1 U769 ( .A(n1063), .B(KEYINPUT12), .Z(n1067) );
NAND2_X1 U770 ( .A1(n1068), .A2(n1069), .ZN(n1063) );
XOR2_X1 U771 ( .A(n1070), .B(n1071), .Z(n1068) );
XNOR2_X1 U772 ( .A(G125), .B(G140), .ZN(n1071) );
NAND2_X1 U773 ( .A1(KEYINPUT62), .A2(n1072), .ZN(n1070) );
XOR2_X1 U774 ( .A(n1073), .B(n1074), .Z(n1072) );
XNOR2_X1 U775 ( .A(n1075), .B(n1076), .ZN(n1074) );
NAND2_X1 U776 ( .A1(KEYINPUT4), .A2(n1077), .ZN(n1075) );
XNOR2_X1 U777 ( .A(n1078), .B(G131), .ZN(n1073) );
NAND2_X1 U778 ( .A1(n1069), .A2(n1079), .ZN(n1066) );
NAND2_X1 U779 ( .A1(G953), .A2(n1080), .ZN(n1079) );
INV_X1 U780 ( .A(n1081), .ZN(n1069) );
NAND2_X1 U781 ( .A1(n1082), .A2(n1083), .ZN(G69) );
NAND2_X1 U782 ( .A1(n1084), .A2(n1061), .ZN(n1083) );
XNOR2_X1 U783 ( .A(n1085), .B(n1086), .ZN(n1084) );
NOR2_X1 U784 ( .A1(n1009), .A2(KEYINPUT26), .ZN(n1086) );
NAND2_X1 U785 ( .A1(n1087), .A2(G953), .ZN(n1082) );
XOR2_X1 U786 ( .A(n1085), .B(n1088), .Z(n1087) );
AND2_X1 U787 ( .A1(G224), .A2(G898), .ZN(n1088) );
NAND2_X1 U788 ( .A1(n1089), .A2(n1090), .ZN(n1085) );
NAND2_X1 U789 ( .A1(G953), .A2(n1091), .ZN(n1090) );
XOR2_X1 U790 ( .A(n1092), .B(KEYINPUT11), .Z(n1089) );
NOR2_X1 U791 ( .A1(n1045), .A2(n1093), .ZN(G66) );
XOR2_X1 U792 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U793 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NOR2_X1 U794 ( .A1(n1045), .A2(n1098), .ZN(G63) );
NOR2_X1 U795 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U796 ( .A(n1101), .B(n1102), .Z(n1100) );
AND2_X1 U797 ( .A1(G478), .A2(n1096), .ZN(n1102) );
AND2_X1 U798 ( .A1(n1103), .A2(KEYINPUT22), .ZN(n1101) );
NOR2_X1 U799 ( .A1(KEYINPUT22), .A2(n1103), .ZN(n1099) );
NOR2_X1 U800 ( .A1(n1045), .A2(n1104), .ZN(G60) );
NOR3_X1 U801 ( .A1(n1054), .A2(n1105), .A3(n1106), .ZN(n1104) );
NOR4_X1 U802 ( .A1(n1107), .A2(n1108), .A3(KEYINPUT18), .A4(n1109), .ZN(n1106) );
INV_X1 U803 ( .A(n1110), .ZN(n1107) );
NOR2_X1 U804 ( .A1(n1111), .A2(n1110), .ZN(n1105) );
NOR3_X1 U805 ( .A1(n1109), .A2(KEYINPUT18), .A3(n1112), .ZN(n1111) );
NOR2_X1 U806 ( .A1(n1060), .A2(n1113), .ZN(n1112) );
INV_X1 U807 ( .A(G475), .ZN(n1109) );
XOR2_X1 U808 ( .A(G104), .B(n1114), .Z(G6) );
NOR2_X1 U809 ( .A1(n1045), .A2(n1115), .ZN(G57) );
XOR2_X1 U810 ( .A(n1116), .B(n1117), .Z(n1115) );
XNOR2_X1 U811 ( .A(n1118), .B(n1119), .ZN(n1117) );
XOR2_X1 U812 ( .A(n1120), .B(n1121), .Z(n1116) );
XNOR2_X1 U813 ( .A(G101), .B(n1122), .ZN(n1121) );
AND2_X1 U814 ( .A1(G472), .A2(n1096), .ZN(n1120) );
NOR2_X1 U815 ( .A1(n1045), .A2(n1123), .ZN(G54) );
XOR2_X1 U816 ( .A(n1124), .B(n1125), .Z(n1123) );
XNOR2_X1 U817 ( .A(n1126), .B(n1127), .ZN(n1125) );
NOR3_X1 U818 ( .A1(n1108), .A2(KEYINPUT51), .A3(n1128), .ZN(n1127) );
INV_X1 U819 ( .A(G469), .ZN(n1128) );
NAND2_X1 U820 ( .A1(KEYINPUT14), .A2(n1129), .ZN(n1126) );
XNOR2_X1 U821 ( .A(n1130), .B(n1131), .ZN(n1124) );
NOR2_X1 U822 ( .A1(n1045), .A2(n1132), .ZN(G51) );
XOR2_X1 U823 ( .A(n1133), .B(n1134), .Z(n1132) );
XNOR2_X1 U824 ( .A(n1135), .B(n1136), .ZN(n1134) );
XOR2_X1 U825 ( .A(n1137), .B(n1138), .Z(n1135) );
NOR2_X1 U826 ( .A1(KEYINPUT35), .A2(n1092), .ZN(n1138) );
NAND2_X1 U827 ( .A1(n1096), .A2(n1139), .ZN(n1137) );
INV_X1 U828 ( .A(n1108), .ZN(n1096) );
NAND2_X1 U829 ( .A1(G902), .A2(n1140), .ZN(n1108) );
NAND2_X1 U830 ( .A1(n1009), .A2(n1010), .ZN(n1140) );
INV_X1 U831 ( .A(n1060), .ZN(n1010) );
NAND2_X1 U832 ( .A1(n1141), .A2(n1142), .ZN(n1060) );
AND4_X1 U833 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1142) );
NOR4_X1 U834 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1141) );
NOR2_X1 U835 ( .A1(n1039), .A2(n1151), .ZN(n1150) );
NOR2_X1 U836 ( .A1(n1034), .A2(n1152), .ZN(n1149) );
NOR2_X1 U837 ( .A1(n1153), .A2(n1154), .ZN(n1148) );
XNOR2_X1 U838 ( .A(KEYINPUT1), .B(n1155), .ZN(n1154) );
INV_X1 U839 ( .A(n1156), .ZN(n1153) );
INV_X1 U840 ( .A(n1113), .ZN(n1009) );
NAND4_X1 U841 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1113) );
NOR4_X1 U842 ( .A1(n1161), .A2(n1162), .A3(n1114), .A4(n1163), .ZN(n1160) );
AND3_X1 U843 ( .A1(n1001), .A2(n1002), .A3(n1164), .ZN(n1114) );
NAND2_X1 U844 ( .A1(n1165), .A2(n1166), .ZN(n1159) );
NAND2_X1 U845 ( .A1(n1167), .A2(n1168), .ZN(n1158) );
NAND2_X1 U846 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND3_X1 U847 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1170) );
XNOR2_X1 U848 ( .A(n1001), .B(KEYINPUT43), .ZN(n1173) );
NAND2_X1 U849 ( .A1(n1164), .A2(n1043), .ZN(n1169) );
NAND3_X1 U850 ( .A1(n1002), .A2(n1003), .A3(n1001), .ZN(n1157) );
XOR2_X1 U851 ( .A(n1174), .B(n1175), .Z(n1133) );
XNOR2_X1 U852 ( .A(n1176), .B(n1177), .ZN(n1175) );
NAND2_X1 U853 ( .A1(KEYINPUT29), .A2(n1178), .ZN(n1177) );
INV_X1 U854 ( .A(G125), .ZN(n1178) );
XNOR2_X1 U855 ( .A(KEYINPUT7), .B(KEYINPUT45), .ZN(n1174) );
NOR2_X1 U856 ( .A1(n1061), .A2(G952), .ZN(n1045) );
XOR2_X1 U857 ( .A(n1179), .B(n1180), .Z(G48) );
NOR2_X1 U858 ( .A1(KEYINPUT37), .A2(n1181), .ZN(n1180) );
INV_X1 U859 ( .A(G146), .ZN(n1181) );
NOR2_X1 U860 ( .A1(n1182), .A2(n1151), .ZN(n1179) );
XNOR2_X1 U861 ( .A(n1164), .B(KEYINPUT52), .ZN(n1182) );
XNOR2_X1 U862 ( .A(n1147), .B(n1183), .ZN(G45) );
NOR2_X1 U863 ( .A1(G143), .A2(KEYINPUT50), .ZN(n1183) );
AND4_X1 U864 ( .A1(n1166), .A2(n1172), .A3(n1043), .A4(n1184), .ZN(n1147) );
NOR2_X1 U865 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U866 ( .A(n1187), .B(n1188), .Z(G42) );
XNOR2_X1 U867 ( .A(G140), .B(KEYINPUT27), .ZN(n1188) );
NAND2_X1 U868 ( .A1(n1156), .A2(n1042), .ZN(n1187) );
XOR2_X1 U869 ( .A(n1143), .B(n1189), .Z(G39) );
NAND2_X1 U870 ( .A1(KEYINPUT58), .A2(G137), .ZN(n1189) );
NAND4_X1 U871 ( .A1(n1020), .A2(n1051), .A3(n1190), .A4(n1191), .ZN(n1143) );
NOR2_X1 U872 ( .A1(n1192), .A2(n1185), .ZN(n1191) );
NAND2_X1 U873 ( .A1(n1193), .A2(n1194), .ZN(G36) );
NAND2_X1 U874 ( .A1(G134), .A2(n1195), .ZN(n1194) );
XOR2_X1 U875 ( .A(n1196), .B(KEYINPUT47), .Z(n1193) );
OR2_X1 U876 ( .A1(n1195), .A2(G134), .ZN(n1196) );
NAND2_X1 U877 ( .A1(n1197), .A2(n1020), .ZN(n1195) );
INV_X1 U878 ( .A(n1034), .ZN(n1020) );
XOR2_X1 U879 ( .A(n1152), .B(KEYINPUT42), .Z(n1197) );
NAND3_X1 U880 ( .A1(n1043), .A2(n1003), .A3(n1198), .ZN(n1152) );
XNOR2_X1 U881 ( .A(G131), .B(n1146), .ZN(G33) );
NAND2_X1 U882 ( .A1(n1156), .A2(n1043), .ZN(n1146) );
NOR3_X1 U883 ( .A1(n1039), .A2(n1034), .A3(n1185), .ZN(n1156) );
NAND2_X1 U884 ( .A1(n1033), .A2(n1199), .ZN(n1034) );
INV_X1 U885 ( .A(n1164), .ZN(n1039) );
XNOR2_X1 U886 ( .A(n1145), .B(n1200), .ZN(G30) );
NOR2_X1 U887 ( .A1(KEYINPUT20), .A2(n1201), .ZN(n1200) );
INV_X1 U888 ( .A(G128), .ZN(n1201) );
OR2_X1 U889 ( .A1(n1151), .A2(n1040), .ZN(n1145) );
INV_X1 U890 ( .A(n1003), .ZN(n1040) );
NAND4_X1 U891 ( .A1(n1190), .A2(n1198), .A3(n1166), .A4(n1051), .ZN(n1151) );
INV_X1 U892 ( .A(n1185), .ZN(n1198) );
NAND2_X1 U893 ( .A1(n1202), .A2(n1203), .ZN(n1185) );
XNOR2_X1 U894 ( .A(n1204), .B(n1162), .ZN(G3) );
AND3_X1 U895 ( .A1(n1043), .A2(n1002), .A3(n1017), .ZN(n1162) );
AND3_X1 U896 ( .A1(n1202), .A2(n1205), .A3(n1166), .ZN(n1002) );
XNOR2_X1 U897 ( .A(G125), .B(n1144), .ZN(G27) );
NAND4_X1 U898 ( .A1(n1042), .A2(n1164), .A3(n1206), .A4(n1203), .ZN(n1144) );
NAND2_X1 U899 ( .A1(n1044), .A2(n1207), .ZN(n1203) );
NAND3_X1 U900 ( .A1(G902), .A2(n1208), .A3(n1081), .ZN(n1207) );
NOR2_X1 U901 ( .A1(G900), .A2(n1061), .ZN(n1081) );
INV_X1 U902 ( .A(n1155), .ZN(n1042) );
XOR2_X1 U903 ( .A(n1209), .B(n1210), .Z(G24) );
XNOR2_X1 U904 ( .A(G122), .B(KEYINPUT33), .ZN(n1210) );
NAND4_X1 U905 ( .A1(n1171), .A2(KEYINPUT23), .A3(n1211), .A4(n1167), .ZN(n1209) );
AND2_X1 U906 ( .A1(n1172), .A2(n1001), .ZN(n1211) );
NOR2_X1 U907 ( .A1(n1051), .A2(n1190), .ZN(n1001) );
NAND2_X1 U908 ( .A1(n1212), .A2(n1213), .ZN(G21) );
NAND2_X1 U909 ( .A1(n1163), .A2(n1214), .ZN(n1213) );
INV_X1 U910 ( .A(n1215), .ZN(n1163) );
XOR2_X1 U911 ( .A(n1216), .B(KEYINPUT54), .Z(n1212) );
NAND2_X1 U912 ( .A1(G119), .A2(n1215), .ZN(n1216) );
NAND4_X1 U913 ( .A1(n1017), .A2(n1167), .A3(n1190), .A4(n1051), .ZN(n1215) );
INV_X1 U914 ( .A(n1217), .ZN(n1190) );
XOR2_X1 U915 ( .A(G116), .B(n1161), .Z(G18) );
AND3_X1 U916 ( .A1(n1167), .A2(n1003), .A3(n1043), .ZN(n1161) );
NOR2_X1 U917 ( .A1(n1046), .A2(n1171), .ZN(n1003) );
INV_X1 U918 ( .A(n1172), .ZN(n1046) );
NOR2_X1 U919 ( .A1(n1018), .A2(n1218), .ZN(n1167) );
XNOR2_X1 U920 ( .A(G113), .B(n1219), .ZN(G15) );
NAND4_X1 U921 ( .A1(n1164), .A2(n1043), .A3(n1206), .A4(n1220), .ZN(n1219) );
XNOR2_X1 U922 ( .A(KEYINPUT17), .B(n1205), .ZN(n1220) );
INV_X1 U923 ( .A(n1018), .ZN(n1206) );
NAND3_X1 U924 ( .A1(n1166), .A2(n1027), .A3(n1024), .ZN(n1018) );
NOR2_X1 U925 ( .A1(n1217), .A2(n1051), .ZN(n1043) );
NOR2_X1 U926 ( .A1(n1186), .A2(n1172), .ZN(n1164) );
XNOR2_X1 U927 ( .A(G110), .B(n1221), .ZN(G12) );
NAND3_X1 U928 ( .A1(n1166), .A2(n1222), .A3(KEYINPUT61), .ZN(n1221) );
XOR2_X1 U929 ( .A(KEYINPUT9), .B(n1165), .Z(n1222) );
NOR4_X1 U930 ( .A1(n1155), .A2(n1192), .A3(n1022), .A4(n1218), .ZN(n1165) );
INV_X1 U931 ( .A(n1205), .ZN(n1218) );
NAND2_X1 U932 ( .A1(n1044), .A2(n1223), .ZN(n1205) );
NAND4_X1 U933 ( .A1(G953), .A2(G902), .A3(n1208), .A4(n1091), .ZN(n1223) );
INV_X1 U934 ( .A(G898), .ZN(n1091) );
NAND3_X1 U935 ( .A1(n1208), .A2(n1061), .A3(G952), .ZN(n1044) );
NAND2_X1 U936 ( .A1(G237), .A2(G234), .ZN(n1208) );
INV_X1 U937 ( .A(n1202), .ZN(n1022) );
NOR2_X1 U938 ( .A1(n1024), .A2(n1048), .ZN(n1202) );
INV_X1 U939 ( .A(n1027), .ZN(n1048) );
NAND2_X1 U940 ( .A1(G221), .A2(n1224), .ZN(n1027) );
XOR2_X1 U941 ( .A(n1225), .B(G469), .Z(n1024) );
NAND2_X1 U942 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
XOR2_X1 U943 ( .A(n1228), .B(n1129), .Z(n1226) );
AND2_X1 U944 ( .A1(n1229), .A2(n1230), .ZN(n1129) );
NAND2_X1 U945 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND2_X1 U946 ( .A1(G227), .A2(n1061), .ZN(n1232) );
OR3_X1 U947 ( .A1(n1080), .A2(G953), .A3(n1231), .ZN(n1229) );
INV_X1 U948 ( .A(G227), .ZN(n1080) );
XNOR2_X1 U949 ( .A(n1233), .B(n1131), .ZN(n1228) );
INV_X1 U950 ( .A(n1118), .ZN(n1131) );
NAND2_X1 U951 ( .A1(KEYINPUT41), .A2(n1130), .ZN(n1233) );
XNOR2_X1 U952 ( .A(n1234), .B(n1136), .ZN(n1130) );
NAND2_X1 U953 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NAND2_X1 U954 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XNOR2_X1 U955 ( .A(KEYINPUT25), .B(n1204), .ZN(n1238) );
XNOR2_X1 U956 ( .A(n1239), .B(KEYINPUT3), .ZN(n1237) );
XOR2_X1 U957 ( .A(KEYINPUT48), .B(n1240), .Z(n1235) );
NOR2_X1 U958 ( .A1(G101), .A2(n1239), .ZN(n1240) );
INV_X1 U959 ( .A(n1017), .ZN(n1192) );
NOR2_X1 U960 ( .A1(n1172), .A2(n1171), .ZN(n1017) );
INV_X1 U961 ( .A(n1186), .ZN(n1171) );
XOR2_X1 U962 ( .A(n1241), .B(n1242), .Z(n1186) );
INV_X1 U963 ( .A(n1052), .ZN(n1242) );
XOR2_X1 U964 ( .A(G475), .B(KEYINPUT19), .Z(n1052) );
XNOR2_X1 U965 ( .A(n1054), .B(KEYINPUT39), .ZN(n1241) );
NOR2_X1 U966 ( .A1(n1110), .A2(G902), .ZN(n1054) );
XNOR2_X1 U967 ( .A(n1243), .B(n1244), .ZN(n1110) );
XOR2_X1 U968 ( .A(n1245), .B(n1246), .Z(n1244) );
XNOR2_X1 U969 ( .A(G140), .B(n1247), .ZN(n1246) );
NOR2_X1 U970 ( .A1(KEYINPUT6), .A2(n1248), .ZN(n1247) );
XOR2_X1 U971 ( .A(n1249), .B(n1250), .Z(n1248) );
NOR2_X1 U972 ( .A1(KEYINPUT15), .A2(n1251), .ZN(n1250) );
XNOR2_X1 U973 ( .A(G104), .B(G113), .ZN(n1249) );
NAND3_X1 U974 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1245) );
NAND2_X1 U975 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
OR3_X1 U976 ( .A1(n1256), .A2(n1255), .A3(n1257), .ZN(n1253) );
INV_X1 U977 ( .A(KEYINPUT59), .ZN(n1256) );
NAND2_X1 U978 ( .A1(n1258), .A2(n1257), .ZN(n1252) );
INV_X1 U979 ( .A(G143), .ZN(n1257) );
NAND2_X1 U980 ( .A1(KEYINPUT59), .A2(n1259), .ZN(n1258) );
XNOR2_X1 U981 ( .A(KEYINPUT46), .B(n1255), .ZN(n1259) );
NAND3_X1 U982 ( .A1(n1260), .A2(n1061), .A3(G214), .ZN(n1255) );
XNOR2_X1 U983 ( .A(n1261), .B(n1262), .ZN(n1243) );
NOR2_X1 U984 ( .A1(KEYINPUT63), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U985 ( .A(n1264), .B(G478), .ZN(n1172) );
NAND2_X1 U986 ( .A1(n1103), .A2(n1227), .ZN(n1264) );
XNOR2_X1 U987 ( .A(n1265), .B(n1266), .ZN(n1103) );
NOR2_X1 U988 ( .A1(KEYINPUT0), .A2(n1267), .ZN(n1266) );
XOR2_X1 U989 ( .A(n1268), .B(n1269), .Z(n1267) );
XNOR2_X1 U990 ( .A(n1270), .B(n1251), .ZN(n1269) );
NAND2_X1 U991 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND2_X1 U992 ( .A1(n1273), .A2(n1078), .ZN(n1272) );
XOR2_X1 U993 ( .A(n1274), .B(KEYINPUT13), .Z(n1271) );
OR2_X1 U994 ( .A1(n1273), .A2(n1078), .ZN(n1274) );
INV_X1 U995 ( .A(G134), .ZN(n1078) );
XOR2_X1 U996 ( .A(n1275), .B(KEYINPUT21), .Z(n1273) );
XNOR2_X1 U997 ( .A(G107), .B(G116), .ZN(n1268) );
NAND3_X1 U998 ( .A1(G234), .A2(n1061), .A3(G217), .ZN(n1265) );
NAND2_X1 U999 ( .A1(n1051), .A2(n1217), .ZN(n1155) );
XNOR2_X1 U1000 ( .A(n1276), .B(n1277), .ZN(n1217) );
NOR2_X1 U1001 ( .A1(KEYINPUT34), .A2(n1057), .ZN(n1277) );
NAND2_X1 U1002 ( .A1(n1278), .A2(n1227), .ZN(n1057) );
XOR2_X1 U1003 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U1004 ( .A(n1119), .B(n1281), .Z(n1280) );
NOR2_X1 U1005 ( .A1(KEYINPUT10), .A2(n1122), .ZN(n1281) );
NAND3_X1 U1006 ( .A1(n1260), .A2(n1061), .A3(G210), .ZN(n1122) );
XNOR2_X1 U1007 ( .A(n1282), .B(n1283), .ZN(n1119) );
INV_X1 U1008 ( .A(n1284), .ZN(n1283) );
XNOR2_X1 U1009 ( .A(n1076), .B(KEYINPUT5), .ZN(n1282) );
XNOR2_X1 U1010 ( .A(G101), .B(n1285), .ZN(n1279) );
NOR2_X1 U1011 ( .A1(KEYINPUT30), .A2(n1118), .ZN(n1285) );
XOR2_X1 U1012 ( .A(n1286), .B(n1263), .Z(n1118) );
INV_X1 U1013 ( .A(G131), .ZN(n1263) );
NAND2_X1 U1014 ( .A1(n1287), .A2(KEYINPUT31), .ZN(n1286) );
XNOR2_X1 U1015 ( .A(G137), .B(G134), .ZN(n1287) );
XNOR2_X1 U1016 ( .A(G472), .B(KEYINPUT49), .ZN(n1276) );
XNOR2_X1 U1017 ( .A(n1288), .B(n1097), .ZN(n1051) );
AND2_X1 U1018 ( .A1(G217), .A2(n1224), .ZN(n1097) );
NAND2_X1 U1019 ( .A1(G234), .A2(n1227), .ZN(n1224) );
NAND2_X1 U1020 ( .A1(n1095), .A2(n1227), .ZN(n1288) );
XNOR2_X1 U1021 ( .A(n1289), .B(n1290), .ZN(n1095) );
XOR2_X1 U1022 ( .A(n1261), .B(n1231), .Z(n1290) );
XOR2_X1 U1023 ( .A(G110), .B(G140), .Z(n1231) );
XOR2_X1 U1024 ( .A(G146), .B(G125), .Z(n1261) );
XOR2_X1 U1025 ( .A(n1291), .B(n1292), .Z(n1289) );
XNOR2_X1 U1026 ( .A(n1077), .B(n1293), .ZN(n1292) );
AND3_X1 U1027 ( .A1(G221), .A2(n1061), .A3(G234), .ZN(n1293) );
INV_X1 U1028 ( .A(G137), .ZN(n1077) );
NAND3_X1 U1029 ( .A1(n1294), .A2(n1295), .A3(KEYINPUT57), .ZN(n1291) );
NAND2_X1 U1030 ( .A1(KEYINPUT44), .A2(n1296), .ZN(n1295) );
XNOR2_X1 U1031 ( .A(G119), .B(n1297), .ZN(n1296) );
OR3_X1 U1032 ( .A1(n1214), .A2(n1297), .A3(KEYINPUT44), .ZN(n1294) );
XOR2_X1 U1033 ( .A(G128), .B(KEYINPUT38), .Z(n1297) );
NOR2_X1 U1034 ( .A1(n1033), .A2(n1032), .ZN(n1166) );
INV_X1 U1035 ( .A(n1199), .ZN(n1032) );
NAND2_X1 U1036 ( .A1(G214), .A2(n1298), .ZN(n1199) );
XOR2_X1 U1037 ( .A(n1299), .B(n1139), .Z(n1033) );
AND2_X1 U1038 ( .A1(G210), .A2(n1298), .ZN(n1139) );
NAND2_X1 U1039 ( .A1(n1227), .A2(n1260), .ZN(n1298) );
INV_X1 U1040 ( .A(G237), .ZN(n1260) );
NAND2_X1 U1041 ( .A1(n1300), .A2(n1227), .ZN(n1299) );
INV_X1 U1042 ( .A(G902), .ZN(n1227) );
XOR2_X1 U1043 ( .A(n1301), .B(n1302), .Z(n1300) );
XNOR2_X1 U1044 ( .A(G125), .B(n1303), .ZN(n1302) );
XNOR2_X1 U1045 ( .A(KEYINPUT60), .B(KEYINPUT2), .ZN(n1303) );
XOR2_X1 U1046 ( .A(n1092), .B(n1304), .Z(n1301) );
XNOR2_X1 U1047 ( .A(n1305), .B(n1136), .ZN(n1304) );
INV_X1 U1048 ( .A(n1076), .ZN(n1136) );
XOR2_X1 U1049 ( .A(G146), .B(n1275), .Z(n1076) );
XOR2_X1 U1050 ( .A(G128), .B(G143), .Z(n1275) );
NOR2_X1 U1051 ( .A1(n1176), .A2(KEYINPUT24), .ZN(n1305) );
AND2_X1 U1052 ( .A1(n1306), .A2(n1061), .ZN(n1176) );
INV_X1 U1053 ( .A(G953), .ZN(n1061) );
XNOR2_X1 U1054 ( .A(G224), .B(KEYINPUT28), .ZN(n1306) );
XOR2_X1 U1055 ( .A(n1307), .B(n1308), .Z(n1092) );
XOR2_X1 U1056 ( .A(n1251), .B(n1309), .Z(n1308) );
XOR2_X1 U1057 ( .A(n1310), .B(G110), .Z(n1309) );
NAND2_X1 U1058 ( .A1(KEYINPUT40), .A2(n1204), .ZN(n1310) );
INV_X1 U1059 ( .A(G101), .ZN(n1204) );
XNOR2_X1 U1060 ( .A(G122), .B(KEYINPUT16), .ZN(n1251) );
XNOR2_X1 U1061 ( .A(n1284), .B(n1239), .ZN(n1307) );
XOR2_X1 U1062 ( .A(G104), .B(G107), .Z(n1239) );
XOR2_X1 U1063 ( .A(G113), .B(n1311), .Z(n1284) );
XNOR2_X1 U1064 ( .A(n1214), .B(G116), .ZN(n1311) );
INV_X1 U1065 ( .A(G119), .ZN(n1214) );
endmodule


