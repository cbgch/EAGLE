//Key = 1111010011111101111100001010101001001000111000111001110111001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360;

XNOR2_X1 U742 ( .A(G107), .B(n1035), .ZN(G9) );
NAND4_X1 U743 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
NOR2_X1 U744 ( .A1(KEYINPUT20), .A2(n1040), .ZN(n1038) );
NOR2_X1 U745 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR4_X1 U746 ( .A1(G953), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1042) );
INV_X1 U747 ( .A(n1046), .ZN(n1045) );
NOR2_X1 U748 ( .A1(n1047), .A2(n1048), .ZN(n1044) );
NOR2_X1 U749 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U751 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
AND2_X1 U752 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U753 ( .A1(n1057), .A2(n1058), .ZN(n1053) );
NOR2_X1 U754 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
AND2_X1 U755 ( .A1(n1056), .A2(n1061), .ZN(n1060) );
NOR2_X1 U756 ( .A1(n1062), .A2(n1040), .ZN(n1059) );
NOR2_X1 U757 ( .A1(n1063), .A2(n1037), .ZN(n1062) );
NOR2_X1 U758 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR4_X1 U759 ( .A1(n1066), .A2(n1040), .A3(n1067), .A4(n1058), .ZN(n1049) );
NOR2_X1 U760 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U761 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR3_X1 U762 ( .A1(n1043), .A2(G953), .A3(G952), .ZN(n1041) );
AND4_X1 U763 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1043) );
NOR3_X1 U764 ( .A1(n1076), .A2(n1067), .A3(n1052), .ZN(n1075) );
XNOR2_X1 U765 ( .A(G478), .B(n1077), .ZN(n1076) );
XNOR2_X1 U766 ( .A(KEYINPUT12), .B(n1078), .ZN(n1074) );
XNOR2_X1 U767 ( .A(n1079), .B(n1080), .ZN(n1073) );
XOR2_X1 U768 ( .A(KEYINPUT49), .B(KEYINPUT42), .Z(n1080) );
XOR2_X1 U769 ( .A(n1081), .B(n1082), .Z(n1072) );
XNOR2_X1 U770 ( .A(KEYINPUT36), .B(n1083), .ZN(n1082) );
XOR2_X1 U771 ( .A(n1084), .B(n1085), .Z(G72) );
XOR2_X1 U772 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND2_X1 U773 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NAND2_X1 U774 ( .A1(G900), .A2(G227), .ZN(n1088) );
NAND2_X1 U775 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
XOR2_X1 U776 ( .A(KEYINPUT57), .B(n1091), .Z(n1090) );
NOR2_X1 U777 ( .A1(G900), .A2(n1092), .ZN(n1091) );
XOR2_X1 U778 ( .A(n1093), .B(n1094), .Z(n1089) );
XOR2_X1 U779 ( .A(n1095), .B(n1096), .Z(n1093) );
AND2_X1 U780 ( .A1(n1097), .A2(n1092), .ZN(n1084) );
XOR2_X1 U781 ( .A(n1098), .B(n1099), .Z(G69) );
NOR2_X1 U782 ( .A1(KEYINPUT27), .A2(n1100), .ZN(n1099) );
XOR2_X1 U783 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U784 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U785 ( .A(n1105), .B(n1106), .ZN(n1104) );
NAND2_X1 U786 ( .A1(n1092), .A2(n1107), .ZN(n1101) );
NAND2_X1 U787 ( .A1(n1108), .A2(n1109), .ZN(n1098) );
NAND2_X1 U788 ( .A1(G953), .A2(n1110), .ZN(n1109) );
XOR2_X1 U789 ( .A(KEYINPUT15), .B(G224), .Z(n1110) );
INV_X1 U790 ( .A(n1103), .ZN(n1108) );
NOR2_X1 U791 ( .A1(n1111), .A2(n1112), .ZN(G66) );
XOR2_X1 U792 ( .A(n1113), .B(n1114), .Z(n1112) );
AND2_X1 U793 ( .A1(G217), .A2(n1115), .ZN(n1114) );
NOR2_X1 U794 ( .A1(KEYINPUT7), .A2(n1116), .ZN(n1113) );
NOR2_X1 U795 ( .A1(n1111), .A2(n1117), .ZN(G63) );
NOR3_X1 U796 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1117) );
NOR4_X1 U797 ( .A1(n1121), .A2(n1122), .A3(KEYINPUT23), .A4(n1123), .ZN(n1120) );
NOR2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1119) );
NOR3_X1 U799 ( .A1(n1123), .A2(KEYINPUT23), .A3(n1046), .ZN(n1124) );
NOR2_X1 U800 ( .A1(n1111), .A2(n1126), .ZN(G60) );
NOR3_X1 U801 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1126) );
AND2_X1 U802 ( .A1(n1130), .A2(KEYINPUT4), .ZN(n1129) );
NOR2_X1 U803 ( .A1(KEYINPUT4), .A2(n1131), .ZN(n1128) );
NOR2_X1 U804 ( .A1(n1132), .A2(n1081), .ZN(n1131) );
NOR2_X1 U805 ( .A1(n1133), .A2(n1130), .ZN(n1132) );
NOR2_X1 U806 ( .A1(n1046), .A2(n1083), .ZN(n1133) );
NOR3_X1 U807 ( .A1(n1122), .A2(n1134), .A3(n1083), .ZN(n1127) );
NOR2_X1 U808 ( .A1(KEYINPUT4), .A2(n1130), .ZN(n1134) );
INV_X1 U809 ( .A(n1115), .ZN(n1122) );
XNOR2_X1 U810 ( .A(G104), .B(n1135), .ZN(G6) );
NAND2_X1 U811 ( .A1(n1136), .A2(n1069), .ZN(n1135) );
XOR2_X1 U812 ( .A(n1137), .B(KEYINPUT18), .Z(n1136) );
NAND4_X1 U813 ( .A1(n1138), .A2(n1037), .A3(n1139), .A4(n1140), .ZN(n1137) );
XNOR2_X1 U814 ( .A(KEYINPUT58), .B(n1040), .ZN(n1139) );
INV_X1 U815 ( .A(n1141), .ZN(n1040) );
NOR4_X1 U816 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(G57) );
NOR2_X1 U817 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U818 ( .A(n1148), .B(KEYINPUT45), .Z(n1147) );
NOR2_X1 U819 ( .A1(n1149), .A2(n1150), .ZN(n1144) );
XOR2_X1 U820 ( .A(n1148), .B(KEYINPUT19), .Z(n1150) );
XOR2_X1 U821 ( .A(n1151), .B(n1152), .Z(n1148) );
XOR2_X1 U822 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U823 ( .A1(n1115), .A2(G472), .ZN(n1154) );
NAND2_X1 U824 ( .A1(KEYINPUT11), .A2(n1155), .ZN(n1151) );
INV_X1 U825 ( .A(G101), .ZN(n1155) );
INV_X1 U826 ( .A(n1146), .ZN(n1149) );
XNOR2_X1 U827 ( .A(n1156), .B(n1157), .ZN(n1146) );
XNOR2_X1 U828 ( .A(KEYINPUT56), .B(n1158), .ZN(n1157) );
XOR2_X1 U829 ( .A(n1159), .B(n1160), .Z(n1156) );
NOR2_X1 U830 ( .A1(KEYINPUT54), .A2(n1161), .ZN(n1160) );
AND3_X1 U831 ( .A1(KEYINPUT22), .A2(G953), .A3(G952), .ZN(n1143) );
NOR2_X1 U832 ( .A1(KEYINPUT22), .A2(n1162), .ZN(n1142) );
INV_X1 U833 ( .A(n1111), .ZN(n1162) );
NOR2_X1 U834 ( .A1(n1111), .A2(n1163), .ZN(G54) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U836 ( .A(n1166), .B(n1167), .Z(n1165) );
NAND2_X1 U837 ( .A1(n1168), .A2(KEYINPUT1), .ZN(n1166) );
XOR2_X1 U838 ( .A(n1169), .B(n1096), .Z(n1168) );
NAND2_X1 U839 ( .A1(KEYINPUT13), .A2(n1170), .ZN(n1169) );
XOR2_X1 U840 ( .A(n1171), .B(n1172), .Z(n1164) );
XNOR2_X1 U841 ( .A(G110), .B(G140), .ZN(n1172) );
NAND2_X1 U842 ( .A1(n1115), .A2(G469), .ZN(n1171) );
NOR2_X1 U843 ( .A1(n1111), .A2(n1173), .ZN(G51) );
XOR2_X1 U844 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U845 ( .A(n1176), .B(n1177), .ZN(n1174) );
NAND2_X1 U846 ( .A1(n1115), .A2(n1178), .ZN(n1176) );
NOR2_X1 U847 ( .A1(n1179), .A2(n1046), .ZN(n1115) );
NOR2_X1 U848 ( .A1(n1107), .A2(n1097), .ZN(n1046) );
NAND2_X1 U849 ( .A1(n1180), .A2(n1181), .ZN(n1097) );
AND4_X1 U850 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181) );
NOR4_X1 U851 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1180) );
AND3_X1 U852 ( .A1(n1190), .A2(n1191), .A3(n1039), .ZN(n1188) );
XNOR2_X1 U853 ( .A(n1192), .B(KEYINPUT47), .ZN(n1191) );
INV_X1 U854 ( .A(n1193), .ZN(n1186) );
NAND3_X1 U855 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1107) );
NOR3_X1 U856 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1196) );
NAND4_X1 U857 ( .A1(n1200), .A2(n1141), .A3(n1201), .A4(n1202), .ZN(n1195) );
NAND2_X1 U858 ( .A1(n1037), .A2(n1203), .ZN(n1194) );
NAND2_X1 U859 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NAND4_X1 U860 ( .A1(n1061), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1205) );
OR2_X1 U861 ( .A1(n1209), .A2(n1036), .ZN(n1208) );
NAND2_X1 U862 ( .A1(n1210), .A2(n1209), .ZN(n1207) );
INV_X1 U863 ( .A(KEYINPUT53), .ZN(n1209) );
NAND2_X1 U864 ( .A1(n1140), .A2(n1211), .ZN(n1210) );
NAND2_X1 U865 ( .A1(n1036), .A2(n1055), .ZN(n1204) );
NAND2_X1 U866 ( .A1(n1212), .A2(n1213), .ZN(n1055) );
NAND2_X1 U867 ( .A1(n1141), .A2(n1214), .ZN(n1213) );
OR2_X1 U868 ( .A1(n1138), .A2(n1039), .ZN(n1214) );
NAND2_X1 U869 ( .A1(n1206), .A2(n1215), .ZN(n1212) );
NOR2_X1 U870 ( .A1(n1092), .A2(G952), .ZN(n1111) );
NAND2_X1 U871 ( .A1(n1216), .A2(n1217), .ZN(G48) );
NAND2_X1 U872 ( .A1(G146), .A2(n1218), .ZN(n1217) );
NAND2_X1 U873 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NAND2_X1 U874 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
INV_X1 U875 ( .A(KEYINPUT33), .ZN(n1222) );
XOR2_X1 U876 ( .A(KEYINPUT31), .B(n1187), .Z(n1219) );
NAND3_X1 U877 ( .A1(KEYINPUT33), .A2(n1221), .A3(n1223), .ZN(n1216) );
XOR2_X1 U878 ( .A(n1187), .B(KEYINPUT29), .Z(n1221) );
AND3_X1 U879 ( .A1(n1138), .A2(n1192), .A3(n1190), .ZN(n1187) );
XNOR2_X1 U880 ( .A(G143), .B(n1224), .ZN(G45) );
NAND2_X1 U881 ( .A1(KEYINPUT63), .A2(n1189), .ZN(n1224) );
AND4_X1 U882 ( .A1(n1201), .A2(n1037), .A3(n1215), .A4(n1225), .ZN(n1189) );
NOR3_X1 U883 ( .A1(n1211), .A2(n1226), .A3(n1227), .ZN(n1225) );
XNOR2_X1 U884 ( .A(G140), .B(n1193), .ZN(G42) );
NAND3_X1 U885 ( .A1(n1061), .A2(n1138), .A3(n1228), .ZN(n1193) );
XNOR2_X1 U886 ( .A(G137), .B(n1185), .ZN(G39) );
NAND2_X1 U887 ( .A1(n1228), .A2(n1229), .ZN(n1185) );
XNOR2_X1 U888 ( .A(G134), .B(n1184), .ZN(G36) );
NAND3_X1 U889 ( .A1(n1215), .A2(n1039), .A3(n1228), .ZN(n1184) );
XNOR2_X1 U890 ( .A(G131), .B(n1183), .ZN(G33) );
NAND3_X1 U891 ( .A1(n1215), .A2(n1138), .A3(n1228), .ZN(n1183) );
NOR3_X1 U892 ( .A1(n1230), .A2(n1226), .A3(n1052), .ZN(n1228) );
NAND2_X1 U893 ( .A1(n1231), .A2(n1071), .ZN(n1052) );
XNOR2_X1 U894 ( .A(G128), .B(n1232), .ZN(G30) );
NAND4_X1 U895 ( .A1(KEYINPUT51), .A2(n1190), .A3(n1039), .A4(n1192), .ZN(n1232) );
NOR4_X1 U896 ( .A1(n1230), .A2(n1211), .A3(n1079), .A4(n1078), .ZN(n1190) );
XNOR2_X1 U897 ( .A(G101), .B(n1233), .ZN(G3) );
NAND4_X1 U898 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1215), .ZN(n1233) );
NOR2_X1 U899 ( .A1(n1237), .A2(n1230), .ZN(n1236) );
XNOR2_X1 U900 ( .A(n1069), .B(KEYINPUT9), .ZN(n1235) );
INV_X1 U901 ( .A(n1211), .ZN(n1069) );
XNOR2_X1 U902 ( .A(n1206), .B(KEYINPUT52), .ZN(n1234) );
XNOR2_X1 U903 ( .A(G125), .B(n1182), .ZN(G27) );
NAND3_X1 U904 ( .A1(n1061), .A2(n1138), .A3(n1238), .ZN(n1182) );
NOR3_X1 U905 ( .A1(n1067), .A2(n1226), .A3(n1211), .ZN(n1238) );
INV_X1 U906 ( .A(n1192), .ZN(n1226) );
NAND2_X1 U907 ( .A1(n1048), .A2(n1239), .ZN(n1192) );
NAND4_X1 U908 ( .A1(G902), .A2(G953), .A3(n1240), .A4(n1241), .ZN(n1239) );
INV_X1 U909 ( .A(G900), .ZN(n1241) );
NAND2_X1 U910 ( .A1(n1242), .A2(n1243), .ZN(G24) );
NAND2_X1 U911 ( .A1(G122), .A2(n1244), .ZN(n1243) );
XOR2_X1 U912 ( .A(n1245), .B(KEYINPUT6), .Z(n1242) );
OR2_X1 U913 ( .A1(n1244), .A2(G122), .ZN(n1245) );
NAND4_X1 U914 ( .A1(n1246), .A2(n1036), .A3(n1247), .A4(n1141), .ZN(n1244) );
NOR2_X1 U915 ( .A1(n1248), .A2(n1249), .ZN(n1141) );
NOR2_X1 U916 ( .A1(n1227), .A2(n1250), .ZN(n1247) );
XNOR2_X1 U917 ( .A(n1056), .B(KEYINPUT61), .ZN(n1246) );
XNOR2_X1 U918 ( .A(n1251), .B(n1197), .ZN(G21) );
AND2_X1 U919 ( .A1(n1229), .A2(n1200), .ZN(n1197) );
NOR3_X1 U920 ( .A1(n1079), .A2(n1078), .A3(n1058), .ZN(n1229) );
INV_X1 U921 ( .A(n1206), .ZN(n1058) );
XOR2_X1 U922 ( .A(G116), .B(n1199), .Z(G18) );
AND3_X1 U923 ( .A1(n1200), .A2(n1039), .A3(n1215), .ZN(n1199) );
NOR2_X1 U924 ( .A1(n1250), .A2(n1252), .ZN(n1039) );
NAND2_X1 U925 ( .A1(n1253), .A2(n1254), .ZN(G15) );
NAND2_X1 U926 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
NAND2_X1 U927 ( .A1(n1257), .A2(n1258), .ZN(n1255) );
OR2_X1 U928 ( .A1(n1198), .A2(KEYINPUT48), .ZN(n1258) );
INV_X1 U929 ( .A(n1259), .ZN(n1198) );
NAND2_X1 U930 ( .A1(KEYINPUT48), .A2(n1260), .ZN(n1257) );
OR2_X1 U931 ( .A1(n1260), .A2(n1256), .ZN(n1253) );
NAND2_X1 U932 ( .A1(KEYINPUT60), .A2(n1259), .ZN(n1260) );
NAND3_X1 U933 ( .A1(n1138), .A2(n1200), .A3(n1215), .ZN(n1259) );
NOR2_X1 U934 ( .A1(n1248), .A2(n1079), .ZN(n1215) );
INV_X1 U935 ( .A(n1249), .ZN(n1079) );
AND2_X1 U936 ( .A1(n1056), .A2(n1036), .ZN(n1200) );
INV_X1 U937 ( .A(n1067), .ZN(n1056) );
NAND2_X1 U938 ( .A1(n1261), .A2(n1065), .ZN(n1067) );
INV_X1 U939 ( .A(n1064), .ZN(n1261) );
NOR2_X1 U940 ( .A1(n1227), .A2(n1201), .ZN(n1138) );
INV_X1 U941 ( .A(n1202), .ZN(n1227) );
XOR2_X1 U942 ( .A(n1262), .B(KEYINPUT8), .Z(n1202) );
XNOR2_X1 U943 ( .A(G110), .B(n1263), .ZN(G12) );
NAND4_X1 U944 ( .A1(n1061), .A2(n1206), .A3(n1036), .A4(n1037), .ZN(n1263) );
INV_X1 U945 ( .A(n1230), .ZN(n1037) );
NAND2_X1 U946 ( .A1(n1064), .A2(n1065), .ZN(n1230) );
NAND2_X1 U947 ( .A1(G221), .A2(n1264), .ZN(n1065) );
XNOR2_X1 U948 ( .A(n1265), .B(G469), .ZN(n1064) );
NAND2_X1 U949 ( .A1(n1266), .A2(n1179), .ZN(n1265) );
XOR2_X1 U950 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U951 ( .A(n1167), .B(n1269), .Z(n1268) );
XNOR2_X1 U952 ( .A(n1161), .B(n1270), .ZN(n1167) );
AND2_X1 U953 ( .A1(n1271), .A2(G227), .ZN(n1270) );
XOR2_X1 U954 ( .A(n1272), .B(n1096), .Z(n1267) );
NAND2_X1 U955 ( .A1(KEYINPUT17), .A2(n1273), .ZN(n1272) );
NOR2_X1 U956 ( .A1(n1211), .A2(n1237), .ZN(n1036) );
INV_X1 U957 ( .A(n1140), .ZN(n1237) );
NAND2_X1 U958 ( .A1(n1048), .A2(n1274), .ZN(n1140) );
NAND3_X1 U959 ( .A1(n1103), .A2(n1240), .A3(G902), .ZN(n1274) );
NOR2_X1 U960 ( .A1(G898), .A2(n1092), .ZN(n1103) );
NAND3_X1 U961 ( .A1(n1240), .A2(n1092), .A3(G952), .ZN(n1048) );
INV_X1 U962 ( .A(G953), .ZN(n1092) );
NAND2_X1 U963 ( .A1(G237), .A2(G234), .ZN(n1240) );
NAND2_X1 U964 ( .A1(n1070), .A2(n1071), .ZN(n1211) );
NAND2_X1 U965 ( .A1(G214), .A2(n1275), .ZN(n1071) );
INV_X1 U966 ( .A(n1231), .ZN(n1070) );
XOR2_X1 U967 ( .A(n1276), .B(n1178), .Z(n1231) );
AND2_X1 U968 ( .A1(G210), .A2(n1275), .ZN(n1178) );
NAND2_X1 U969 ( .A1(n1277), .A2(n1179), .ZN(n1275) );
NAND3_X1 U970 ( .A1(n1278), .A2(n1279), .A3(n1179), .ZN(n1276) );
NAND2_X1 U971 ( .A1(n1280), .A2(n1177), .ZN(n1279) );
NAND2_X1 U972 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND2_X1 U973 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
INV_X1 U974 ( .A(KEYINPUT62), .ZN(n1284) );
NAND2_X1 U975 ( .A1(KEYINPUT62), .A2(n1175), .ZN(n1281) );
OR2_X1 U976 ( .A1(n1177), .A2(n1283), .ZN(n1278) );
NAND2_X1 U977 ( .A1(KEYINPUT2), .A2(n1175), .ZN(n1283) );
XNOR2_X1 U978 ( .A(n1159), .B(n1285), .ZN(n1175) );
XOR2_X1 U979 ( .A(G125), .B(n1286), .Z(n1285) );
AND2_X1 U980 ( .A1(n1271), .A2(G224), .ZN(n1286) );
XOR2_X1 U981 ( .A(n1105), .B(n1287), .Z(n1177) );
NOR2_X1 U982 ( .A1(KEYINPUT39), .A2(n1106), .ZN(n1287) );
NAND2_X1 U983 ( .A1(n1288), .A2(n1289), .ZN(n1106) );
NAND2_X1 U984 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NAND2_X1 U985 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND2_X1 U986 ( .A1(KEYINPUT3), .A2(n1256), .ZN(n1293) );
NAND2_X1 U987 ( .A1(G113), .A2(n1294), .ZN(n1288) );
NAND2_X1 U988 ( .A1(KEYINPUT3), .A2(n1295), .ZN(n1294) );
NAND2_X1 U989 ( .A1(n1296), .A2(n1292), .ZN(n1295) );
INV_X1 U990 ( .A(KEYINPUT25), .ZN(n1292) );
XNOR2_X1 U991 ( .A(n1269), .B(G122), .ZN(n1105) );
XNOR2_X1 U992 ( .A(n1170), .B(G110), .ZN(n1269) );
XNOR2_X1 U993 ( .A(G101), .B(n1297), .ZN(n1170) );
XOR2_X1 U994 ( .A(G107), .B(G104), .Z(n1297) );
NOR2_X1 U995 ( .A1(n1201), .A2(n1252), .ZN(n1206) );
INV_X1 U996 ( .A(n1262), .ZN(n1252) );
XNOR2_X1 U997 ( .A(n1298), .B(n1081), .ZN(n1262) );
NOR2_X1 U998 ( .A1(n1130), .A2(G902), .ZN(n1081) );
XOR2_X1 U999 ( .A(n1299), .B(n1300), .Z(n1130) );
XOR2_X1 U1000 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1001 ( .A(n1303), .B(n1304), .Z(n1302) );
NOR2_X1 U1002 ( .A1(KEYINPUT59), .A2(n1305), .ZN(n1304) );
XOR2_X1 U1003 ( .A(n1306), .B(n1307), .Z(n1305) );
XNOR2_X1 U1004 ( .A(n1223), .B(G140), .ZN(n1307) );
NAND2_X1 U1005 ( .A1(KEYINPUT16), .A2(G125), .ZN(n1306) );
NAND3_X1 U1006 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1303) );
NAND2_X1 U1007 ( .A1(G113), .A2(n1311), .ZN(n1310) );
OR3_X1 U1008 ( .A1(n1311), .A2(n1312), .A3(G122), .ZN(n1309) );
INV_X1 U1009 ( .A(KEYINPUT5), .ZN(n1311) );
NAND2_X1 U1010 ( .A1(G122), .A2(n1312), .ZN(n1308) );
NAND2_X1 U1011 ( .A1(KEYINPUT26), .A2(n1256), .ZN(n1312) );
NAND3_X1 U1012 ( .A1(G214), .A2(n1277), .A3(n1271), .ZN(n1301) );
XOR2_X1 U1013 ( .A(n1313), .B(n1314), .Z(n1299) );
XOR2_X1 U1014 ( .A(KEYINPUT32), .B(G143), .Z(n1314) );
XNOR2_X1 U1015 ( .A(G104), .B(G131), .ZN(n1313) );
NAND2_X1 U1016 ( .A1(KEYINPUT28), .A2(n1083), .ZN(n1298) );
INV_X1 U1017 ( .A(G475), .ZN(n1083) );
INV_X1 U1018 ( .A(n1250), .ZN(n1201) );
XOR2_X1 U1019 ( .A(n1315), .B(n1077), .Z(n1250) );
INV_X1 U1020 ( .A(n1118), .ZN(n1077) );
NOR2_X1 U1021 ( .A1(n1125), .A2(G902), .ZN(n1118) );
INV_X1 U1022 ( .A(n1121), .ZN(n1125) );
XNOR2_X1 U1023 ( .A(n1316), .B(n1317), .ZN(n1121) );
XOR2_X1 U1024 ( .A(G116), .B(n1318), .Z(n1317) );
XOR2_X1 U1025 ( .A(n1319), .B(n1320), .Z(n1318) );
XOR2_X1 U1026 ( .A(n1321), .B(n1322), .Z(n1320) );
AND3_X1 U1027 ( .A1(G217), .A2(G234), .A3(n1271), .ZN(n1322) );
XNOR2_X1 U1028 ( .A(G107), .B(G134), .ZN(n1321) );
XOR2_X1 U1029 ( .A(n1323), .B(G143), .Z(n1319) );
XNOR2_X1 U1030 ( .A(KEYINPUT41), .B(KEYINPUT0), .ZN(n1323) );
XNOR2_X1 U1031 ( .A(G128), .B(G122), .ZN(n1316) );
NAND2_X1 U1032 ( .A1(KEYINPUT10), .A2(n1123), .ZN(n1315) );
INV_X1 U1033 ( .A(G478), .ZN(n1123) );
NOR2_X1 U1034 ( .A1(n1249), .A2(n1078), .ZN(n1061) );
INV_X1 U1035 ( .A(n1248), .ZN(n1078) );
XNOR2_X1 U1036 ( .A(n1324), .B(n1325), .ZN(n1248) );
NOR2_X1 U1037 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
XOR2_X1 U1038 ( .A(KEYINPUT55), .B(G217), .Z(n1327) );
INV_X1 U1039 ( .A(n1264), .ZN(n1326) );
NAND2_X1 U1040 ( .A1(G234), .A2(n1179), .ZN(n1264) );
NAND2_X1 U1041 ( .A1(n1116), .A2(n1179), .ZN(n1324) );
XNOR2_X1 U1042 ( .A(n1328), .B(n1329), .ZN(n1116) );
XOR2_X1 U1043 ( .A(n1330), .B(n1331), .Z(n1329) );
XNOR2_X1 U1044 ( .A(G110), .B(n1332), .ZN(n1331) );
NOR3_X1 U1045 ( .A1(n1333), .A2(KEYINPUT38), .A3(n1334), .ZN(n1332) );
NOR2_X1 U1046 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
XOR2_X1 U1047 ( .A(KEYINPUT35), .B(n1337), .Z(n1333) );
AND2_X1 U1048 ( .A1(n1336), .A2(n1335), .ZN(n1337) );
NAND3_X1 U1049 ( .A1(n1271), .A2(G234), .A3(G221), .ZN(n1336) );
NAND2_X1 U1050 ( .A1(n1338), .A2(KEYINPUT40), .ZN(n1330) );
XNOR2_X1 U1051 ( .A(n1094), .B(n1339), .ZN(n1338) );
NOR2_X1 U1052 ( .A1(G146), .A2(KEYINPUT50), .ZN(n1339) );
XNOR2_X1 U1053 ( .A(G125), .B(n1273), .ZN(n1094) );
INV_X1 U1054 ( .A(G140), .ZN(n1273) );
XNOR2_X1 U1055 ( .A(G119), .B(n1340), .ZN(n1328) );
XNOR2_X1 U1056 ( .A(KEYINPUT21), .B(n1341), .ZN(n1340) );
XNOR2_X1 U1057 ( .A(n1342), .B(G472), .ZN(n1249) );
NAND2_X1 U1058 ( .A1(n1343), .A2(n1179), .ZN(n1342) );
INV_X1 U1059 ( .A(G902), .ZN(n1179) );
XOR2_X1 U1060 ( .A(n1344), .B(n1345), .Z(n1343) );
XNOR2_X1 U1061 ( .A(n1346), .B(n1159), .ZN(n1345) );
NAND2_X1 U1062 ( .A1(n1347), .A2(n1348), .ZN(n1159) );
NAND2_X1 U1063 ( .A1(n1096), .A2(KEYINPUT46), .ZN(n1348) );
XNOR2_X1 U1064 ( .A(n1349), .B(n1350), .ZN(n1096) );
XNOR2_X1 U1065 ( .A(G128), .B(G146), .ZN(n1349) );
NAND2_X1 U1066 ( .A1(n1351), .A2(n1352), .ZN(n1347) );
INV_X1 U1067 ( .A(KEYINPUT46), .ZN(n1352) );
XNOR2_X1 U1068 ( .A(n1353), .B(n1341), .ZN(n1351) );
INV_X1 U1069 ( .A(G128), .ZN(n1341) );
NAND2_X1 U1070 ( .A1(n1350), .A2(n1223), .ZN(n1353) );
INV_X1 U1071 ( .A(G146), .ZN(n1223) );
XOR2_X1 U1072 ( .A(G143), .B(KEYINPUT34), .Z(n1350) );
XOR2_X1 U1073 ( .A(n1354), .B(n1161), .Z(n1346) );
XNOR2_X1 U1074 ( .A(n1095), .B(KEYINPUT24), .ZN(n1161) );
XNOR2_X1 U1075 ( .A(G131), .B(n1355), .ZN(n1095) );
XNOR2_X1 U1076 ( .A(n1335), .B(G134), .ZN(n1355) );
INV_X1 U1077 ( .A(G137), .ZN(n1335) );
NAND2_X1 U1078 ( .A1(KEYINPUT30), .A2(n1158), .ZN(n1354) );
NAND2_X1 U1079 ( .A1(n1356), .A2(n1357), .ZN(n1158) );
NAND2_X1 U1080 ( .A1(n1296), .A2(n1256), .ZN(n1357) );
INV_X1 U1081 ( .A(G113), .ZN(n1256) );
XOR2_X1 U1082 ( .A(n1358), .B(KEYINPUT14), .Z(n1356) );
NAND2_X1 U1083 ( .A1(G113), .A2(n1290), .ZN(n1358) );
INV_X1 U1084 ( .A(n1296), .ZN(n1290) );
XOR2_X1 U1085 ( .A(G116), .B(n1251), .Z(n1296) );
INV_X1 U1086 ( .A(G119), .ZN(n1251) );
XOR2_X1 U1087 ( .A(n1359), .B(n1360), .Z(n1344) );
NOR2_X1 U1088 ( .A1(G101), .A2(KEYINPUT44), .ZN(n1360) );
XOR2_X1 U1089 ( .A(n1153), .B(KEYINPUT37), .Z(n1359) );
NAND3_X1 U1090 ( .A1(n1271), .A2(n1277), .A3(G210), .ZN(n1153) );
INV_X1 U1091 ( .A(G237), .ZN(n1277) );
XNOR2_X1 U1092 ( .A(G953), .B(KEYINPUT43), .ZN(n1271) );
endmodule


