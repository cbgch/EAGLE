//Key = 1101110111100001101010111111111111111100000001011101000110111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373;

XOR2_X1 U743 ( .A(G107), .B(n1039), .Z(G9) );
NOR2_X1 U744 ( .A1(n1040), .A2(n1041), .ZN(G75) );
NOR4_X1 U745 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1041) );
NOR2_X1 U746 ( .A1(n1046), .A2(n1047), .ZN(n1043) );
NOR2_X1 U747 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U748 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U749 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U750 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR3_X1 U751 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1054) );
NOR3_X1 U752 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
NOR2_X1 U753 ( .A1(n1062), .A2(n1063), .ZN(n1056) );
XNOR2_X1 U754 ( .A(n1064), .B(n1065), .ZN(n1063) );
AND2_X1 U755 ( .A1(KEYINPUT45), .A2(n1066), .ZN(n1065) );
NOR3_X1 U756 ( .A1(n1062), .A2(n1067), .A3(n1060), .ZN(n1052) );
NOR2_X1 U757 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR4_X1 U758 ( .A1(n1070), .A2(n1055), .A3(n1060), .A4(n1062), .ZN(n1048) );
INV_X1 U759 ( .A(n1071), .ZN(n1062) );
NOR2_X1 U760 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR3_X1 U761 ( .A1(n1044), .A2(G952), .A3(n1042), .ZN(n1040) );
AND4_X1 U762 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1042) );
NOR4_X1 U763 ( .A1(n1078), .A2(n1066), .A3(n1055), .A4(n1079), .ZN(n1077) );
XOR2_X1 U764 ( .A(n1080), .B(n1081), .Z(n1079) );
XOR2_X1 U765 ( .A(n1082), .B(KEYINPUT61), .Z(n1081) );
NAND2_X1 U766 ( .A1(KEYINPUT30), .A2(n1083), .ZN(n1080) );
XNOR2_X1 U767 ( .A(KEYINPUT29), .B(n1084), .ZN(n1083) );
INV_X1 U768 ( .A(n1085), .ZN(n1066) );
NOR3_X1 U769 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1076) );
NOR2_X1 U770 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XOR2_X1 U771 ( .A(KEYINPUT57), .B(n1091), .Z(n1090) );
NOR2_X1 U772 ( .A1(G475), .A2(n1092), .ZN(n1087) );
XOR2_X1 U773 ( .A(KEYINPUT23), .B(n1091), .Z(n1092) );
XNOR2_X1 U774 ( .A(G469), .B(n1093), .ZN(n1086) );
NAND2_X1 U775 ( .A1(n1094), .A2(n1095), .ZN(n1075) );
NAND2_X1 U776 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NAND2_X1 U777 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
INV_X1 U778 ( .A(KEYINPUT32), .ZN(n1099) );
NAND2_X1 U779 ( .A1(KEYINPUT32), .A2(n1100), .ZN(n1096) );
NAND2_X1 U780 ( .A1(n1098), .A2(n1101), .ZN(n1100) );
NAND3_X1 U781 ( .A1(n1098), .A2(n1101), .A3(n1102), .ZN(n1074) );
INV_X1 U782 ( .A(KEYINPUT44), .ZN(n1101) );
INV_X1 U783 ( .A(n1103), .ZN(n1044) );
XOR2_X1 U784 ( .A(n1104), .B(n1105), .Z(G72) );
NOR2_X1 U785 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U786 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U787 ( .A(n1110), .B(n1111), .Z(n1109) );
XNOR2_X1 U788 ( .A(G125), .B(G140), .ZN(n1108) );
AND2_X1 U789 ( .A1(n1112), .A2(n1113), .ZN(n1106) );
NAND2_X1 U790 ( .A1(n1114), .A2(n1115), .ZN(n1104) );
NAND2_X1 U791 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U792 ( .A1(G953), .A2(n1118), .ZN(n1114) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1118) );
XOR2_X1 U794 ( .A(n1119), .B(n1120), .Z(G69) );
XOR2_X1 U795 ( .A(n1121), .B(n1122), .Z(n1120) );
NAND2_X1 U796 ( .A1(G953), .A2(n1123), .ZN(n1122) );
NAND2_X1 U797 ( .A1(G898), .A2(G224), .ZN(n1123) );
NAND2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1121) );
NAND2_X1 U799 ( .A1(n1113), .A2(n1126), .ZN(n1125) );
XNOR2_X1 U800 ( .A(n1127), .B(n1128), .ZN(n1124) );
XNOR2_X1 U801 ( .A(n1129), .B(n1130), .ZN(n1127) );
AND2_X1 U802 ( .A1(n1131), .A2(n1117), .ZN(n1119) );
NOR2_X1 U803 ( .A1(n1132), .A2(n1133), .ZN(G66) );
XNOR2_X1 U804 ( .A(n1134), .B(n1135), .ZN(n1133) );
NAND4_X1 U805 ( .A1(KEYINPUT37), .A2(G902), .A3(G217), .A4(n1136), .ZN(n1134) );
XNOR2_X1 U806 ( .A(KEYINPUT51), .B(n1045), .ZN(n1136) );
NOR2_X1 U807 ( .A1(n1132), .A2(n1137), .ZN(G63) );
XOR2_X1 U808 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U809 ( .A1(n1084), .A2(n1140), .ZN(n1139) );
NAND2_X1 U810 ( .A1(n1141), .A2(KEYINPUT49), .ZN(n1138) );
XNOR2_X1 U811 ( .A(n1142), .B(KEYINPUT0), .ZN(n1141) );
NOR2_X1 U812 ( .A1(n1132), .A2(n1143), .ZN(G60) );
NOR3_X1 U813 ( .A1(n1091), .A2(n1144), .A3(n1145), .ZN(n1143) );
NOR3_X1 U814 ( .A1(n1146), .A2(n1089), .A3(n1140), .ZN(n1145) );
NOR2_X1 U815 ( .A1(n1147), .A2(n1148), .ZN(n1144) );
NOR2_X1 U816 ( .A1(n1149), .A2(n1089), .ZN(n1148) );
NAND2_X1 U817 ( .A1(n1150), .A2(n1151), .ZN(G6) );
NAND2_X1 U818 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U819 ( .A(KEYINPUT36), .B(n1154), .Z(n1150) );
NOR2_X1 U820 ( .A1(n1152), .A2(n1153), .ZN(n1154) );
NOR2_X1 U821 ( .A1(n1132), .A2(n1155), .ZN(G57) );
XOR2_X1 U822 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U823 ( .A1(n1158), .A2(KEYINPUT22), .ZN(n1156) );
XOR2_X1 U824 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U825 ( .A1(n1161), .A2(n1140), .ZN(n1160) );
NOR2_X1 U826 ( .A1(n1132), .A2(n1162), .ZN(G54) );
XOR2_X1 U827 ( .A(n1163), .B(n1164), .Z(n1162) );
XNOR2_X1 U828 ( .A(n1165), .B(n1166), .ZN(n1164) );
XOR2_X1 U829 ( .A(n1167), .B(n1168), .Z(n1163) );
NOR2_X1 U830 ( .A1(KEYINPUT19), .A2(n1169), .ZN(n1168) );
XOR2_X1 U831 ( .A(n1170), .B(n1171), .Z(n1167) );
NOR2_X1 U832 ( .A1(n1172), .A2(n1140), .ZN(n1171) );
INV_X1 U833 ( .A(G469), .ZN(n1172) );
NOR2_X1 U834 ( .A1(n1132), .A2(n1173), .ZN(G51) );
XOR2_X1 U835 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U836 ( .A1(n1098), .A2(n1140), .ZN(n1175) );
NAND2_X1 U837 ( .A1(G902), .A2(n1045), .ZN(n1140) );
INV_X1 U838 ( .A(n1149), .ZN(n1045) );
NOR2_X1 U839 ( .A1(n1131), .A2(n1116), .ZN(n1149) );
NAND4_X1 U840 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1116) );
AND4_X1 U841 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1179) );
NAND2_X1 U842 ( .A1(n1184), .A2(n1185), .ZN(n1178) );
NAND2_X1 U843 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NAND2_X1 U844 ( .A1(n1072), .A2(n1188), .ZN(n1187) );
XNOR2_X1 U845 ( .A(KEYINPUT14), .B(n1189), .ZN(n1188) );
NAND2_X1 U846 ( .A1(n1073), .A2(n1190), .ZN(n1186) );
XNOR2_X1 U847 ( .A(KEYINPUT21), .B(n1189), .ZN(n1190) );
INV_X1 U848 ( .A(n1191), .ZN(n1184) );
NAND4_X1 U849 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1177) );
NAND2_X1 U850 ( .A1(n1196), .A2(n1071), .ZN(n1176) );
XOR2_X1 U851 ( .A(n1197), .B(KEYINPUT15), .Z(n1196) );
NAND3_X1 U852 ( .A1(n1072), .A2(n1198), .A3(n1199), .ZN(n1197) );
XNOR2_X1 U853 ( .A(KEYINPUT41), .B(n1200), .ZN(n1198) );
NAND4_X1 U854 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1131) );
NOR4_X1 U855 ( .A1(n1205), .A2(n1039), .A3(n1152), .A4(n1206), .ZN(n1204) );
INV_X1 U856 ( .A(n1207), .ZN(n1206) );
NOR3_X1 U857 ( .A1(n1055), .A2(n1208), .A3(n1209), .ZN(n1152) );
NOR3_X1 U858 ( .A1(n1210), .A2(n1208), .A3(n1055), .ZN(n1039) );
INV_X1 U859 ( .A(n1211), .ZN(n1205) );
NOR2_X1 U860 ( .A1(n1212), .A2(n1213), .ZN(n1203) );
NAND4_X1 U861 ( .A1(n1072), .A2(n1068), .A3(n1214), .A4(n1215), .ZN(n1202) );
OR2_X1 U862 ( .A1(n1216), .A2(KEYINPUT2), .ZN(n1215) );
NAND2_X1 U863 ( .A1(KEYINPUT2), .A2(n1217), .ZN(n1214) );
NAND3_X1 U864 ( .A1(n1218), .A2(n1189), .A3(n1219), .ZN(n1217) );
INV_X1 U865 ( .A(n1060), .ZN(n1219) );
NAND3_X1 U866 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1201) );
XNOR2_X1 U867 ( .A(n1069), .B(KEYINPUT9), .ZN(n1222) );
NAND2_X1 U868 ( .A1(KEYINPUT47), .A2(n1223), .ZN(n1174) );
XOR2_X1 U869 ( .A(n1224), .B(n1225), .Z(n1223) );
XOR2_X1 U870 ( .A(n1226), .B(n1227), .Z(n1225) );
NAND2_X1 U871 ( .A1(KEYINPUT18), .A2(n1228), .ZN(n1226) );
XOR2_X1 U872 ( .A(n1229), .B(n1230), .Z(n1224) );
XNOR2_X1 U873 ( .A(KEYINPUT56), .B(n1231), .ZN(n1230) );
NOR2_X1 U874 ( .A1(n1117), .A2(G952), .ZN(n1132) );
INV_X1 U875 ( .A(G953), .ZN(n1117) );
XOR2_X1 U876 ( .A(n1232), .B(n1233), .Z(G48) );
XOR2_X1 U877 ( .A(KEYINPUT17), .B(G146), .Z(n1233) );
NOR3_X1 U878 ( .A1(n1191), .A2(n1189), .A3(n1209), .ZN(n1232) );
XNOR2_X1 U879 ( .A(G143), .B(n1234), .ZN(G45) );
NAND4_X1 U880 ( .A1(n1235), .A2(KEYINPUT28), .A3(n1236), .A4(n1192), .ZN(n1234) );
NOR2_X1 U881 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XNOR2_X1 U882 ( .A(n1193), .B(KEYINPUT33), .ZN(n1235) );
XNOR2_X1 U883 ( .A(G140), .B(n1239), .ZN(G42) );
NAND3_X1 U884 ( .A1(n1071), .A2(n1199), .A3(n1240), .ZN(n1239) );
NOR3_X1 U885 ( .A1(n1200), .A2(KEYINPUT40), .A3(n1209), .ZN(n1240) );
INV_X1 U886 ( .A(n1072), .ZN(n1209) );
NAND2_X1 U887 ( .A1(n1241), .A2(n1242), .ZN(G39) );
OR2_X1 U888 ( .A1(n1183), .A2(G137), .ZN(n1242) );
XOR2_X1 U889 ( .A(n1243), .B(KEYINPUT6), .Z(n1241) );
NAND2_X1 U890 ( .A1(G137), .A2(n1183), .ZN(n1243) );
NAND3_X1 U891 ( .A1(n1199), .A2(n1244), .A3(n1071), .ZN(n1183) );
XNOR2_X1 U892 ( .A(n1182), .B(n1245), .ZN(G36) );
NOR2_X1 U893 ( .A1(KEYINPUT43), .A2(n1246), .ZN(n1245) );
NAND3_X1 U894 ( .A1(n1192), .A2(n1073), .A3(n1071), .ZN(n1182) );
XOR2_X1 U895 ( .A(n1181), .B(n1247), .Z(G33) );
XNOR2_X1 U896 ( .A(G131), .B(KEYINPUT12), .ZN(n1247) );
NAND3_X1 U897 ( .A1(n1192), .A2(n1072), .A3(n1071), .ZN(n1181) );
NOR2_X1 U898 ( .A1(n1061), .A2(n1078), .ZN(n1071) );
INV_X1 U899 ( .A(n1059), .ZN(n1078) );
AND2_X1 U900 ( .A1(n1199), .A2(n1068), .ZN(n1192) );
XNOR2_X1 U901 ( .A(n1248), .B(n1249), .ZN(G30) );
NOR3_X1 U902 ( .A1(n1191), .A2(n1189), .A3(n1210), .ZN(n1249) );
NAND3_X1 U903 ( .A1(n1250), .A2(n1251), .A3(n1199), .ZN(n1191) );
AND3_X1 U904 ( .A1(n1085), .A2(n1064), .A3(n1252), .ZN(n1199) );
NAND2_X1 U905 ( .A1(n1253), .A2(n1254), .ZN(G3) );
NAND2_X1 U906 ( .A1(G101), .A2(n1211), .ZN(n1254) );
XOR2_X1 U907 ( .A(KEYINPUT1), .B(n1255), .Z(n1253) );
NOR2_X1 U908 ( .A1(G101), .A2(n1211), .ZN(n1255) );
NAND3_X1 U909 ( .A1(n1220), .A2(n1221), .A3(n1068), .ZN(n1211) );
INV_X1 U910 ( .A(n1208), .ZN(n1220) );
XNOR2_X1 U911 ( .A(G125), .B(n1180), .ZN(G27) );
NAND4_X1 U912 ( .A1(n1069), .A2(n1057), .A3(n1072), .A4(n1252), .ZN(n1180) );
NAND2_X1 U913 ( .A1(n1047), .A2(n1256), .ZN(n1252) );
NAND2_X1 U914 ( .A1(n1257), .A2(n1112), .ZN(n1256) );
INV_X1 U915 ( .A(G900), .ZN(n1112) );
INV_X1 U916 ( .A(n1200), .ZN(n1069) );
XNOR2_X1 U917 ( .A(n1258), .B(n1213), .ZN(G24) );
NOR4_X1 U918 ( .A1(n1259), .A2(n1055), .A3(n1238), .A4(n1237), .ZN(n1213) );
OR2_X1 U919 ( .A1(n1251), .A2(n1250), .ZN(n1055) );
XOR2_X1 U920 ( .A(G119), .B(n1212), .Z(G21) );
AND2_X1 U921 ( .A1(n1244), .A2(n1216), .ZN(n1212) );
AND3_X1 U922 ( .A1(n1250), .A2(n1251), .A3(n1221), .ZN(n1244) );
XNOR2_X1 U923 ( .A(G116), .B(n1207), .ZN(G18) );
NAND2_X1 U924 ( .A1(n1260), .A2(n1073), .ZN(n1207) );
XNOR2_X1 U925 ( .A(G113), .B(n1261), .ZN(G15) );
NAND2_X1 U926 ( .A1(n1260), .A2(n1072), .ZN(n1261) );
NOR2_X1 U927 ( .A1(n1195), .A2(n1238), .ZN(n1072) );
AND2_X1 U928 ( .A1(n1216), .A2(n1068), .ZN(n1260) );
NOR2_X1 U929 ( .A1(n1251), .A2(n1262), .ZN(n1068) );
INV_X1 U930 ( .A(n1259), .ZN(n1216) );
NAND2_X1 U931 ( .A1(n1057), .A2(n1218), .ZN(n1259) );
NOR2_X1 U932 ( .A1(n1060), .A2(n1189), .ZN(n1057) );
NAND2_X1 U933 ( .A1(n1263), .A2(n1085), .ZN(n1060) );
XOR2_X1 U934 ( .A(KEYINPUT45), .B(n1064), .Z(n1263) );
XOR2_X1 U935 ( .A(G110), .B(n1264), .Z(G12) );
NOR3_X1 U936 ( .A1(n1200), .A2(n1051), .A3(n1208), .ZN(n1264) );
NAND4_X1 U937 ( .A1(n1193), .A2(n1218), .A3(n1085), .A4(n1064), .ZN(n1208) );
NAND2_X1 U938 ( .A1(n1265), .A2(n1266), .ZN(n1064) );
NAND2_X1 U939 ( .A1(G469), .A2(n1093), .ZN(n1266) );
XOR2_X1 U940 ( .A(n1267), .B(KEYINPUT54), .Z(n1265) );
OR2_X1 U941 ( .A1(n1093), .A2(G469), .ZN(n1267) );
NAND2_X1 U942 ( .A1(n1268), .A2(n1269), .ZN(n1093) );
XOR2_X1 U943 ( .A(n1270), .B(n1271), .Z(n1268) );
XOR2_X1 U944 ( .A(n1170), .B(n1272), .Z(n1271) );
NAND2_X1 U945 ( .A1(KEYINPUT58), .A2(n1165), .ZN(n1272) );
XOR2_X1 U946 ( .A(n1273), .B(n1274), .Z(n1165) );
XNOR2_X1 U947 ( .A(G101), .B(KEYINPUT39), .ZN(n1273) );
NAND2_X1 U948 ( .A1(G227), .A2(n1275), .ZN(n1170) );
XNOR2_X1 U949 ( .A(n1166), .B(n1276), .ZN(n1270) );
INV_X1 U950 ( .A(n1169), .ZN(n1276) );
XNOR2_X1 U951 ( .A(n1110), .B(n1277), .ZN(n1166) );
XOR2_X1 U952 ( .A(KEYINPUT52), .B(n1111), .Z(n1277) );
XOR2_X1 U953 ( .A(n1278), .B(KEYINPUT46), .Z(n1110) );
NAND3_X1 U954 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1278) );
OR2_X1 U955 ( .A1(n1248), .A2(n1282), .ZN(n1281) );
NAND2_X1 U956 ( .A1(n1283), .A2(n1284), .ZN(n1280) );
INV_X1 U957 ( .A(KEYINPUT24), .ZN(n1284) );
NAND2_X1 U958 ( .A1(n1285), .A2(n1248), .ZN(n1283) );
XNOR2_X1 U959 ( .A(KEYINPUT8), .B(n1282), .ZN(n1285) );
NAND2_X1 U960 ( .A1(KEYINPUT24), .A2(n1286), .ZN(n1279) );
NAND2_X1 U961 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
NAND3_X1 U962 ( .A1(KEYINPUT8), .A2(n1248), .A3(n1282), .ZN(n1288) );
OR2_X1 U963 ( .A1(n1282), .A2(KEYINPUT8), .ZN(n1287) );
NAND2_X1 U964 ( .A1(G221), .A2(n1289), .ZN(n1085) );
NAND2_X1 U965 ( .A1(G234), .A2(n1269), .ZN(n1289) );
NAND2_X1 U966 ( .A1(n1047), .A2(n1290), .ZN(n1218) );
NAND2_X1 U967 ( .A1(n1257), .A2(n1126), .ZN(n1290) );
INV_X1 U968 ( .A(G898), .ZN(n1126) );
AND3_X1 U969 ( .A1(G902), .A2(n1291), .A3(n1113), .ZN(n1257) );
XNOR2_X1 U970 ( .A(G953), .B(KEYINPUT5), .ZN(n1113) );
NAND3_X1 U971 ( .A1(n1103), .A2(n1291), .A3(G952), .ZN(n1047) );
NAND2_X1 U972 ( .A1(G237), .A2(G234), .ZN(n1291) );
XOR2_X1 U973 ( .A(G953), .B(KEYINPUT3), .Z(n1103) );
INV_X1 U974 ( .A(n1189), .ZN(n1193) );
NAND2_X1 U975 ( .A1(n1061), .A2(n1059), .ZN(n1189) );
NAND2_X1 U976 ( .A1(n1292), .A2(n1293), .ZN(n1059) );
XNOR2_X1 U977 ( .A(KEYINPUT53), .B(n1294), .ZN(n1292) );
XNOR2_X1 U978 ( .A(n1102), .B(n1098), .ZN(n1061) );
NAND2_X1 U979 ( .A1(G210), .A2(n1293), .ZN(n1098) );
NAND2_X1 U980 ( .A1(n1295), .A2(n1269), .ZN(n1293) );
INV_X1 U981 ( .A(n1095), .ZN(n1102) );
NAND2_X1 U982 ( .A1(n1296), .A2(n1269), .ZN(n1095) );
XOR2_X1 U983 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U984 ( .A(n1229), .B(n1299), .Z(n1298) );
NAND2_X1 U985 ( .A1(KEYINPUT20), .A2(n1227), .ZN(n1299) );
NAND2_X1 U986 ( .A1(n1300), .A2(n1301), .ZN(n1229) );
NAND2_X1 U987 ( .A1(n1130), .A2(n1302), .ZN(n1301) );
XOR2_X1 U988 ( .A(KEYINPUT27), .B(n1303), .Z(n1300) );
NOR2_X1 U989 ( .A1(n1130), .A2(n1302), .ZN(n1303) );
XNOR2_X1 U990 ( .A(n1128), .B(n1304), .ZN(n1302) );
NOR2_X1 U991 ( .A1(KEYINPUT38), .A2(n1129), .ZN(n1304) );
XOR2_X1 U992 ( .A(n1305), .B(n1306), .Z(n1129) );
XOR2_X1 U993 ( .A(n1307), .B(KEYINPUT34), .Z(n1305) );
NAND2_X1 U994 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND2_X1 U995 ( .A1(G119), .A2(n1310), .ZN(n1309) );
XOR2_X1 U996 ( .A(KEYINPUT55), .B(n1311), .Z(n1308) );
NOR2_X1 U997 ( .A1(G119), .A2(n1310), .ZN(n1311) );
NAND2_X1 U998 ( .A1(n1312), .A2(n1313), .ZN(n1128) );
NAND2_X1 U999 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
INV_X1 U1000 ( .A(G101), .ZN(n1315) );
XNOR2_X1 U1001 ( .A(n1274), .B(KEYINPUT48), .ZN(n1314) );
NAND2_X1 U1002 ( .A1(n1316), .A2(G101), .ZN(n1312) );
XNOR2_X1 U1003 ( .A(n1274), .B(KEYINPUT50), .ZN(n1316) );
XNOR2_X1 U1004 ( .A(G107), .B(n1153), .ZN(n1274) );
INV_X1 U1005 ( .A(G104), .ZN(n1153) );
XNOR2_X1 U1006 ( .A(G110), .B(G122), .ZN(n1130) );
XNOR2_X1 U1007 ( .A(G125), .B(n1228), .ZN(n1297) );
NAND2_X1 U1008 ( .A1(G224), .A2(n1275), .ZN(n1228) );
INV_X1 U1009 ( .A(n1221), .ZN(n1051) );
NAND2_X1 U1010 ( .A1(n1317), .A2(n1318), .ZN(n1221) );
OR2_X1 U1011 ( .A1(n1210), .A2(KEYINPUT16), .ZN(n1318) );
INV_X1 U1012 ( .A(n1073), .ZN(n1210) );
NOR2_X1 U1013 ( .A1(n1194), .A2(n1237), .ZN(n1073) );
INV_X1 U1014 ( .A(n1238), .ZN(n1194) );
NAND3_X1 U1015 ( .A1(n1238), .A2(n1237), .A3(KEYINPUT16), .ZN(n1317) );
INV_X1 U1016 ( .A(n1195), .ZN(n1237) );
XOR2_X1 U1017 ( .A(n1082), .B(n1084), .Z(n1195) );
INV_X1 U1018 ( .A(G478), .ZN(n1084) );
NAND2_X1 U1019 ( .A1(n1142), .A2(n1269), .ZN(n1082) );
XNOR2_X1 U1020 ( .A(n1319), .B(n1320), .ZN(n1142) );
XOR2_X1 U1021 ( .A(n1321), .B(n1322), .Z(n1320) );
NOR2_X1 U1022 ( .A1(G116), .A2(KEYINPUT13), .ZN(n1322) );
AND3_X1 U1023 ( .A1(G234), .A2(n1275), .A3(G217), .ZN(n1321) );
XOR2_X1 U1024 ( .A(n1323), .B(n1324), .Z(n1319) );
NOR2_X1 U1025 ( .A1(KEYINPUT62), .A2(n1325), .ZN(n1324) );
XNOR2_X1 U1026 ( .A(n1248), .B(n1326), .ZN(n1325) );
XNOR2_X1 U1027 ( .A(G143), .B(n1246), .ZN(n1326) );
XNOR2_X1 U1028 ( .A(G107), .B(G122), .ZN(n1323) );
XOR2_X1 U1029 ( .A(n1091), .B(n1089), .Z(n1238) );
INV_X1 U1030 ( .A(G475), .ZN(n1089) );
NOR2_X1 U1031 ( .A1(n1147), .A2(G902), .ZN(n1091) );
INV_X1 U1032 ( .A(n1146), .ZN(n1147) );
NAND2_X1 U1033 ( .A1(n1327), .A2(n1328), .ZN(n1146) );
OR2_X1 U1034 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XOR2_X1 U1035 ( .A(n1331), .B(KEYINPUT11), .Z(n1327) );
NAND2_X1 U1036 ( .A1(n1330), .A2(n1329), .ZN(n1331) );
NAND2_X1 U1037 ( .A1(n1332), .A2(n1333), .ZN(n1329) );
NAND4_X1 U1038 ( .A1(KEYINPUT59), .A2(n1334), .A3(n1335), .A4(n1336), .ZN(n1333) );
NAND2_X1 U1039 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
NAND2_X1 U1040 ( .A1(n1339), .A2(n1340), .ZN(n1335) );
NAND3_X1 U1041 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1332) );
NAND2_X1 U1042 ( .A1(KEYINPUT59), .A2(n1334), .ZN(n1343) );
NAND2_X1 U1043 ( .A1(n1339), .A2(n1338), .ZN(n1342) );
XNOR2_X1 U1044 ( .A(KEYINPUT60), .B(n1344), .ZN(n1339) );
NAND2_X1 U1045 ( .A1(n1340), .A2(n1337), .ZN(n1341) );
XNOR2_X1 U1046 ( .A(n1344), .B(n1345), .ZN(n1337) );
XOR2_X1 U1047 ( .A(KEYINPUT63), .B(KEYINPUT10), .Z(n1345) );
XOR2_X1 U1048 ( .A(n1346), .B(n1347), .Z(n1344) );
NOR2_X1 U1049 ( .A1(n1348), .A2(n1294), .ZN(n1347) );
INV_X1 U1050 ( .A(G214), .ZN(n1294) );
XNOR2_X1 U1051 ( .A(G131), .B(G143), .ZN(n1346) );
XNOR2_X1 U1052 ( .A(n1349), .B(n1350), .ZN(n1330) );
XNOR2_X1 U1053 ( .A(KEYINPUT4), .B(n1258), .ZN(n1350) );
INV_X1 U1054 ( .A(G122), .ZN(n1258) );
XNOR2_X1 U1055 ( .A(G104), .B(n1306), .ZN(n1349) );
NAND2_X1 U1056 ( .A1(n1262), .A2(n1251), .ZN(n1200) );
NAND3_X1 U1057 ( .A1(n1351), .A2(n1352), .A3(n1353), .ZN(n1251) );
NAND2_X1 U1058 ( .A1(n1354), .A2(n1135), .ZN(n1353) );
OR3_X1 U1059 ( .A1(n1135), .A2(n1354), .A3(G902), .ZN(n1352) );
NOR2_X1 U1060 ( .A1(n1355), .A2(G234), .ZN(n1354) );
INV_X1 U1061 ( .A(G217), .ZN(n1355) );
XNOR2_X1 U1062 ( .A(n1356), .B(n1357), .ZN(n1135) );
XNOR2_X1 U1063 ( .A(n1340), .B(n1358), .ZN(n1357) );
XNOR2_X1 U1064 ( .A(n1359), .B(n1169), .ZN(n1358) );
XOR2_X1 U1065 ( .A(G110), .B(n1334), .Z(n1169) );
INV_X1 U1066 ( .A(G140), .ZN(n1334) );
NAND2_X1 U1067 ( .A1(KEYINPUT26), .A2(G128), .ZN(n1359) );
INV_X1 U1068 ( .A(n1338), .ZN(n1340) );
XOR2_X1 U1069 ( .A(G146), .B(n1231), .Z(n1338) );
INV_X1 U1070 ( .A(G125), .ZN(n1231) );
XOR2_X1 U1071 ( .A(n1360), .B(n1361), .Z(n1356) );
XOR2_X1 U1072 ( .A(KEYINPUT7), .B(G137), .Z(n1361) );
XOR2_X1 U1073 ( .A(n1362), .B(G119), .Z(n1360) );
NAND3_X1 U1074 ( .A1(G221), .A2(n1275), .A3(G234), .ZN(n1362) );
NAND2_X1 U1075 ( .A1(G902), .A2(G217), .ZN(n1351) );
INV_X1 U1076 ( .A(n1250), .ZN(n1262) );
XOR2_X1 U1077 ( .A(n1363), .B(n1161), .Z(n1250) );
INV_X1 U1078 ( .A(G472), .ZN(n1161) );
NAND2_X1 U1079 ( .A1(n1364), .A2(n1269), .ZN(n1363) );
INV_X1 U1080 ( .A(G902), .ZN(n1269) );
XOR2_X1 U1081 ( .A(n1159), .B(n1157), .Z(n1364) );
XNOR2_X1 U1082 ( .A(G101), .B(n1365), .ZN(n1157) );
NOR2_X1 U1083 ( .A1(n1348), .A2(n1366), .ZN(n1365) );
INV_X1 U1084 ( .A(G210), .ZN(n1366) );
NAND2_X1 U1085 ( .A1(n1275), .A2(n1295), .ZN(n1348) );
INV_X1 U1086 ( .A(G237), .ZN(n1295) );
XOR2_X1 U1087 ( .A(G953), .B(KEYINPUT31), .Z(n1275) );
XOR2_X1 U1088 ( .A(n1367), .B(n1368), .Z(n1159) );
XNOR2_X1 U1089 ( .A(n1310), .B(n1369), .ZN(n1368) );
XOR2_X1 U1090 ( .A(KEYINPUT42), .B(G119), .Z(n1369) );
INV_X1 U1091 ( .A(G116), .ZN(n1310) );
XOR2_X1 U1092 ( .A(n1370), .B(n1306), .Z(n1367) );
XOR2_X1 U1093 ( .A(G113), .B(KEYINPUT35), .Z(n1306) );
XNOR2_X1 U1094 ( .A(n1227), .B(n1111), .ZN(n1370) );
XNOR2_X1 U1095 ( .A(n1371), .B(n1372), .ZN(n1111) );
XNOR2_X1 U1096 ( .A(G137), .B(n1246), .ZN(n1372) );
INV_X1 U1097 ( .A(G134), .ZN(n1246) );
INV_X1 U1098 ( .A(G131), .ZN(n1371) );
XOR2_X1 U1099 ( .A(n1373), .B(n1248), .Z(n1227) );
INV_X1 U1100 ( .A(G128), .ZN(n1248) );
NAND2_X1 U1101 ( .A1(KEYINPUT25), .A2(n1282), .ZN(n1373) );
XNOR2_X1 U1102 ( .A(G146), .B(G143), .ZN(n1282) );
endmodule


