//Key = 0100010100011011011101100000011000110011010011000111000110011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394;

XNOR2_X1 U763 ( .A(G107), .B(n1050), .ZN(G9) );
NOR2_X1 U764 ( .A1(n1051), .A2(n1052), .ZN(G75) );
NOR4_X1 U765 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
XOR2_X1 U766 ( .A(n1057), .B(KEYINPUT9), .Z(n1055) );
NAND3_X1 U767 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
XOR2_X1 U768 ( .A(n1061), .B(KEYINPUT40), .Z(n1060) );
NAND3_X1 U769 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
NAND3_X1 U770 ( .A1(n1065), .A2(n1066), .A3(n1064), .ZN(n1059) );
NAND4_X1 U771 ( .A1(n1063), .A2(n1065), .A3(n1067), .A4(n1068), .ZN(n1058) );
NAND2_X1 U772 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NAND2_X1 U773 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XOR2_X1 U774 ( .A(KEYINPUT16), .B(n1073), .Z(n1072) );
NAND2_X1 U775 ( .A1(n1074), .A2(n1075), .ZN(n1069) );
NAND4_X1 U776 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1053) );
NAND3_X1 U777 ( .A1(n1063), .A2(n1080), .A3(n1064), .ZN(n1077) );
AND3_X1 U778 ( .A1(n1071), .A2(n1068), .A3(n1074), .ZN(n1064) );
NAND3_X1 U779 ( .A1(n1081), .A2(n1068), .A3(n1065), .ZN(n1076) );
NAND2_X1 U780 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND4_X1 U781 ( .A1(n1074), .A2(n1084), .A3(n1071), .A4(n1085), .ZN(n1083) );
INV_X1 U782 ( .A(n1086), .ZN(n1085) );
NAND2_X1 U783 ( .A1(n1063), .A2(n1087), .ZN(n1082) );
NAND2_X1 U784 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U785 ( .A1(n1090), .A2(n1071), .A3(n1091), .ZN(n1089) );
NAND2_X1 U786 ( .A1(n1074), .A2(n1092), .ZN(n1088) );
AND3_X1 U787 ( .A1(n1078), .A2(n1079), .A3(n1093), .ZN(n1051) );
NAND4_X1 U788 ( .A1(n1094), .A2(n1086), .A3(n1095), .A4(n1096), .ZN(n1078) );
NOR4_X1 U789 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
XNOR2_X1 U790 ( .A(n1101), .B(n1102), .ZN(n1098) );
XNOR2_X1 U791 ( .A(n1103), .B(KEYINPUT18), .ZN(n1101) );
XNOR2_X1 U792 ( .A(n1104), .B(n1105), .ZN(n1097) );
NAND2_X1 U793 ( .A1(KEYINPUT22), .A2(n1106), .ZN(n1104) );
NOR2_X1 U794 ( .A1(n1107), .A2(n1091), .ZN(n1095) );
NAND2_X1 U795 ( .A1(G469), .A2(n1108), .ZN(n1094) );
NAND3_X1 U796 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(G72) );
OR2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND3_X1 U798 ( .A1(n1113), .A2(n1112), .A3(G953), .ZN(n1110) );
NAND2_X1 U799 ( .A1(G900), .A2(G227), .ZN(n1113) );
NAND2_X1 U800 ( .A1(n1114), .A2(n1079), .ZN(n1109) );
NAND2_X1 U801 ( .A1(n1112), .A2(n1115), .ZN(n1114) );
NAND2_X1 U802 ( .A1(n1116), .A2(n1056), .ZN(n1115) );
OR2_X1 U803 ( .A1(n1116), .A2(n1117), .ZN(n1112) );
XNOR2_X1 U804 ( .A(KEYINPUT60), .B(n1118), .ZN(n1117) );
NOR2_X1 U805 ( .A1(n1119), .A2(G953), .ZN(n1118) );
NAND3_X1 U806 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1116) );
XOR2_X1 U807 ( .A(n1123), .B(KEYINPUT43), .Z(n1122) );
OR2_X1 U808 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND2_X1 U809 ( .A1(n1124), .A2(n1125), .ZN(n1121) );
XOR2_X1 U810 ( .A(n1126), .B(n1127), .Z(n1124) );
XNOR2_X1 U811 ( .A(n1128), .B(n1129), .ZN(n1127) );
NAND2_X1 U812 ( .A1(G953), .A2(n1130), .ZN(n1120) );
XOR2_X1 U813 ( .A(n1131), .B(n1132), .Z(G69) );
XOR2_X1 U814 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U815 ( .A1(n1135), .A2(G953), .ZN(n1134) );
NOR2_X1 U816 ( .A1(n1136), .A2(n1137), .ZN(n1133) );
XOR2_X1 U817 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U818 ( .A(n1140), .B(KEYINPUT10), .Z(n1139) );
NAND2_X1 U819 ( .A1(n1141), .A2(n1142), .ZN(n1138) );
NAND2_X1 U820 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U821 ( .A(KEYINPUT39), .B(n1145), .Z(n1141) );
NOR2_X1 U822 ( .A1(n1143), .A2(n1144), .ZN(n1145) );
NOR2_X1 U823 ( .A1(n1079), .A2(n1146), .ZN(n1136) );
XOR2_X1 U824 ( .A(KEYINPUT27), .B(G898), .Z(n1146) );
NOR2_X1 U825 ( .A1(n1147), .A2(n1079), .ZN(n1131) );
AND2_X1 U826 ( .A1(G224), .A2(G898), .ZN(n1147) );
NOR2_X1 U827 ( .A1(n1148), .A2(n1149), .ZN(G66) );
NOR3_X1 U828 ( .A1(n1103), .A2(n1150), .A3(n1151), .ZN(n1149) );
NOR3_X1 U829 ( .A1(n1152), .A2(n1102), .A3(n1153), .ZN(n1151) );
INV_X1 U830 ( .A(n1154), .ZN(n1152) );
NOR2_X1 U831 ( .A1(n1155), .A2(n1154), .ZN(n1150) );
NOR2_X1 U832 ( .A1(n1156), .A2(n1102), .ZN(n1155) );
NOR2_X1 U833 ( .A1(n1056), .A2(n1054), .ZN(n1156) );
NOR2_X1 U834 ( .A1(n1148), .A2(n1157), .ZN(G63) );
XNOR2_X1 U835 ( .A(n1158), .B(n1159), .ZN(n1157) );
NOR2_X1 U836 ( .A1(n1160), .A2(n1153), .ZN(n1159) );
NOR2_X1 U837 ( .A1(n1148), .A2(n1161), .ZN(G60) );
XOR2_X1 U838 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U839 ( .A1(n1164), .A2(n1153), .ZN(n1162) );
NAND2_X1 U840 ( .A1(n1165), .A2(n1166), .ZN(G6) );
NAND3_X1 U841 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1166) );
NAND2_X1 U842 ( .A1(G104), .A2(n1170), .ZN(n1165) );
NAND2_X1 U843 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND2_X1 U844 ( .A1(n1167), .A2(n1173), .ZN(n1172) );
INV_X1 U845 ( .A(KEYINPUT12), .ZN(n1173) );
NAND2_X1 U846 ( .A1(KEYINPUT12), .A2(n1174), .ZN(n1171) );
NAND2_X1 U847 ( .A1(n1167), .A2(n1168), .ZN(n1174) );
INV_X1 U848 ( .A(KEYINPUT63), .ZN(n1168) );
AND3_X1 U849 ( .A1(n1175), .A2(n1176), .A3(n1062), .ZN(n1167) );
XOR2_X1 U850 ( .A(KEYINPUT53), .B(n1071), .Z(n1176) );
NOR2_X1 U851 ( .A1(n1148), .A2(n1177), .ZN(G57) );
XOR2_X1 U852 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U853 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U854 ( .A1(KEYINPUT32), .A2(n1182), .ZN(n1181) );
NAND2_X1 U855 ( .A1(n1183), .A2(n1184), .ZN(n1180) );
XOR2_X1 U856 ( .A(n1185), .B(KEYINPUT26), .Z(n1183) );
XOR2_X1 U857 ( .A(n1186), .B(n1187), .Z(n1178) );
NOR2_X1 U858 ( .A1(KEYINPUT33), .A2(n1188), .ZN(n1187) );
NOR2_X1 U859 ( .A1(n1189), .A2(n1153), .ZN(n1188) );
NOR2_X1 U860 ( .A1(n1148), .A2(n1190), .ZN(G54) );
XOR2_X1 U861 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U862 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U863 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XOR2_X1 U864 ( .A(n1197), .B(KEYINPUT62), .Z(n1196) );
NAND2_X1 U865 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NOR2_X1 U866 ( .A1(n1199), .A2(n1198), .ZN(n1195) );
XNOR2_X1 U867 ( .A(G140), .B(n1200), .ZN(n1198) );
NOR2_X1 U868 ( .A1(KEYINPUT57), .A2(n1201), .ZN(n1200) );
NOR2_X1 U869 ( .A1(n1202), .A2(n1153), .ZN(n1193) );
INV_X1 U870 ( .A(G469), .ZN(n1202) );
NOR3_X1 U871 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(G51) );
AND2_X1 U872 ( .A1(KEYINPUT55), .A2(n1148), .ZN(n1205) );
NOR2_X1 U873 ( .A1(n1079), .A2(G952), .ZN(n1148) );
NOR3_X1 U874 ( .A1(KEYINPUT55), .A2(n1079), .A3(n1093), .ZN(n1204) );
INV_X1 U875 ( .A(G952), .ZN(n1093) );
XNOR2_X1 U876 ( .A(n1206), .B(n1207), .ZN(n1203) );
XOR2_X1 U877 ( .A(n1208), .B(n1209), .Z(n1207) );
NOR2_X1 U878 ( .A1(KEYINPUT6), .A2(n1210), .ZN(n1209) );
NOR2_X1 U879 ( .A1(n1105), .A2(n1153), .ZN(n1208) );
NAND2_X1 U880 ( .A1(G902), .A2(n1211), .ZN(n1153) );
NAND2_X1 U881 ( .A1(n1135), .A2(n1119), .ZN(n1211) );
INV_X1 U882 ( .A(n1056), .ZN(n1119) );
NAND4_X1 U883 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1056) );
NOR4_X1 U884 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1215) );
NOR2_X1 U885 ( .A1(n1220), .A2(n1221), .ZN(n1214) );
NOR2_X1 U886 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NOR2_X1 U887 ( .A1(n1224), .A2(n1225), .ZN(n1220) );
NOR2_X1 U888 ( .A1(n1226), .A2(n1227), .ZN(n1224) );
NOR3_X1 U889 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1226) );
NAND3_X1 U890 ( .A1(n1231), .A2(n1223), .A3(n1065), .ZN(n1228) );
INV_X1 U891 ( .A(KEYINPUT30), .ZN(n1223) );
INV_X1 U892 ( .A(n1054), .ZN(n1135) );
NAND4_X1 U893 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1054) );
AND4_X1 U894 ( .A1(n1236), .A2(n1237), .A3(n1050), .A4(n1238), .ZN(n1235) );
OR3_X1 U895 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(n1238) );
NOR2_X1 U896 ( .A1(KEYINPUT41), .A2(n1242), .ZN(n1241) );
NOR2_X1 U897 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
AND2_X1 U898 ( .A1(n1245), .A2(KEYINPUT41), .ZN(n1240) );
NAND3_X1 U899 ( .A1(n1175), .A2(n1080), .A3(n1071), .ZN(n1050) );
NOR2_X1 U900 ( .A1(n1246), .A2(n1247), .ZN(n1234) );
INV_X1 U901 ( .A(n1248), .ZN(n1247) );
NOR3_X1 U902 ( .A1(n1229), .A2(n1099), .A3(n1245), .ZN(n1246) );
NAND3_X1 U903 ( .A1(n1071), .A2(n1175), .A3(n1062), .ZN(n1232) );
XNOR2_X1 U904 ( .A(G146), .B(n1212), .ZN(G48) );
NAND3_X1 U905 ( .A1(n1249), .A2(n1062), .A3(n1250), .ZN(n1212) );
XNOR2_X1 U906 ( .A(G143), .B(n1213), .ZN(G45) );
NAND4_X1 U907 ( .A1(n1250), .A2(n1075), .A3(n1251), .A4(n1252), .ZN(n1213) );
XNOR2_X1 U908 ( .A(n1253), .B(n1218), .ZN(G42) );
AND2_X1 U909 ( .A1(n1254), .A2(n1092), .ZN(n1218) );
XNOR2_X1 U910 ( .A(G137), .B(n1222), .ZN(G39) );
NAND4_X1 U911 ( .A1(n1074), .A2(n1255), .A3(n1249), .A4(n1065), .ZN(n1222) );
XOR2_X1 U912 ( .A(n1256), .B(n1257), .Z(G36) );
NOR2_X1 U913 ( .A1(n1258), .A2(n1225), .ZN(n1257) );
XNOR2_X1 U914 ( .A(n1227), .B(KEYINPUT8), .ZN(n1258) );
AND2_X1 U915 ( .A1(n1255), .A2(n1259), .ZN(n1227) );
NAND2_X1 U916 ( .A1(KEYINPUT21), .A2(n1260), .ZN(n1256) );
XNOR2_X1 U917 ( .A(n1261), .B(n1217), .ZN(G33) );
AND2_X1 U918 ( .A1(n1254), .A2(n1075), .ZN(n1217) );
AND3_X1 U919 ( .A1(n1255), .A2(n1062), .A3(n1074), .ZN(n1254) );
INV_X1 U920 ( .A(n1225), .ZN(n1074) );
NAND2_X1 U921 ( .A1(n1090), .A2(n1262), .ZN(n1225) );
XOR2_X1 U922 ( .A(G128), .B(n1219), .Z(G30) );
AND3_X1 U923 ( .A1(n1249), .A2(n1080), .A3(n1250), .ZN(n1219) );
AND2_X1 U924 ( .A1(n1255), .A2(n1073), .ZN(n1250) );
NOR2_X1 U925 ( .A1(n1230), .A2(n1231), .ZN(n1255) );
INV_X1 U926 ( .A(n1066), .ZN(n1231) );
INV_X1 U927 ( .A(n1229), .ZN(n1249) );
XNOR2_X1 U928 ( .A(G101), .B(n1237), .ZN(G3) );
NAND3_X1 U929 ( .A1(n1175), .A2(n1065), .A3(n1075), .ZN(n1237) );
XNOR2_X1 U930 ( .A(n1263), .B(n1216), .ZN(G27) );
AND4_X1 U931 ( .A1(n1264), .A2(n1092), .A3(n1062), .A4(n1265), .ZN(n1216) );
INV_X1 U932 ( .A(n1230), .ZN(n1264) );
NAND3_X1 U933 ( .A1(n1266), .A2(n1068), .A3(n1267), .ZN(n1230) );
NAND2_X1 U934 ( .A1(n1268), .A2(n1079), .ZN(n1267) );
NAND2_X1 U935 ( .A1(G952), .A2(KEYINPUT5), .ZN(n1268) );
NAND2_X1 U936 ( .A1(n1269), .A2(n1270), .ZN(n1266) );
NAND2_X1 U937 ( .A1(G902), .A2(n1130), .ZN(n1270) );
INV_X1 U938 ( .A(G900), .ZN(n1130) );
NAND2_X1 U939 ( .A1(G952), .A2(n1271), .ZN(n1269) );
NAND2_X1 U940 ( .A1(G953), .A2(KEYINPUT5), .ZN(n1271) );
XNOR2_X1 U941 ( .A(G122), .B(n1233), .ZN(G24) );
NAND4_X1 U942 ( .A1(n1272), .A2(n1071), .A3(n1251), .A4(n1252), .ZN(n1233) );
NOR2_X1 U943 ( .A1(n1273), .A2(n1274), .ZN(n1071) );
XNOR2_X1 U944 ( .A(G119), .B(n1275), .ZN(G21) );
NAND3_X1 U945 ( .A1(n1065), .A2(n1276), .A3(n1272), .ZN(n1275) );
XNOR2_X1 U946 ( .A(KEYINPUT13), .B(n1229), .ZN(n1276) );
NAND2_X1 U947 ( .A1(n1274), .A2(n1273), .ZN(n1229) );
XOR2_X1 U948 ( .A(n1277), .B(G116), .Z(G18) );
NAND2_X1 U949 ( .A1(KEYINPUT19), .A2(n1278), .ZN(n1277) );
NAND2_X1 U950 ( .A1(n1259), .A2(n1272), .ZN(n1278) );
INV_X1 U951 ( .A(n1239), .ZN(n1259) );
NAND2_X1 U952 ( .A1(n1075), .A2(n1080), .ZN(n1239) );
NAND2_X1 U953 ( .A1(n1279), .A2(n1280), .ZN(n1080) );
OR2_X1 U954 ( .A1(n1099), .A2(KEYINPUT59), .ZN(n1280) );
INV_X1 U955 ( .A(n1065), .ZN(n1099) );
NAND3_X1 U956 ( .A1(n1252), .A2(n1281), .A3(KEYINPUT59), .ZN(n1279) );
XNOR2_X1 U957 ( .A(G113), .B(n1236), .ZN(G15) );
NAND3_X1 U958 ( .A1(n1272), .A2(n1075), .A3(n1062), .ZN(n1236) );
NOR2_X1 U959 ( .A1(n1252), .A2(n1281), .ZN(n1062) );
INV_X1 U960 ( .A(n1251), .ZN(n1281) );
AND2_X1 U961 ( .A1(n1282), .A2(n1274), .ZN(n1075) );
INV_X1 U962 ( .A(n1245), .ZN(n1272) );
NAND2_X1 U963 ( .A1(n1265), .A2(n1244), .ZN(n1245) );
INV_X1 U964 ( .A(n1243), .ZN(n1265) );
NAND2_X1 U965 ( .A1(n1063), .A2(n1073), .ZN(n1243) );
AND2_X1 U966 ( .A1(n1084), .A2(n1283), .ZN(n1063) );
XNOR2_X1 U967 ( .A(G110), .B(n1248), .ZN(G12) );
NAND3_X1 U968 ( .A1(n1175), .A2(n1065), .A3(n1092), .ZN(n1248) );
NOR2_X1 U969 ( .A1(n1274), .A2(n1282), .ZN(n1092) );
INV_X1 U970 ( .A(n1273), .ZN(n1282) );
NAND3_X1 U971 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1273) );
OR2_X1 U972 ( .A1(n1102), .A2(KEYINPUT7), .ZN(n1286) );
NAND3_X1 U973 ( .A1(KEYINPUT7), .A2(n1102), .A3(n1287), .ZN(n1285) );
NAND2_X1 U974 ( .A1(n1288), .A2(n1289), .ZN(n1284) );
NAND2_X1 U975 ( .A1(n1290), .A2(KEYINPUT7), .ZN(n1289) );
XOR2_X1 U976 ( .A(n1102), .B(KEYINPUT25), .Z(n1290) );
NAND2_X1 U977 ( .A1(G217), .A2(n1291), .ZN(n1102) );
INV_X1 U978 ( .A(n1287), .ZN(n1288) );
XOR2_X1 U979 ( .A(n1103), .B(KEYINPUT4), .Z(n1287) );
NOR2_X1 U980 ( .A1(n1154), .A2(G902), .ZN(n1103) );
XNOR2_X1 U981 ( .A(n1292), .B(n1293), .ZN(n1154) );
XNOR2_X1 U982 ( .A(n1294), .B(n1295), .ZN(n1293) );
XOR2_X1 U983 ( .A(n1296), .B(n1297), .Z(n1295) );
NOR2_X1 U984 ( .A1(KEYINPUT42), .A2(n1298), .ZN(n1297) );
XNOR2_X1 U985 ( .A(G146), .B(n1125), .ZN(n1298) );
XNOR2_X1 U986 ( .A(G125), .B(n1253), .ZN(n1125) );
NAND3_X1 U987 ( .A1(n1299), .A2(n1079), .A3(G221), .ZN(n1296) );
XOR2_X1 U988 ( .A(KEYINPUT47), .B(G234), .Z(n1299) );
XNOR2_X1 U989 ( .A(G110), .B(n1300), .ZN(n1292) );
XNOR2_X1 U990 ( .A(n1301), .B(G128), .ZN(n1300) );
XOR2_X1 U991 ( .A(n1100), .B(KEYINPUT20), .Z(n1274) );
XOR2_X1 U992 ( .A(n1302), .B(n1189), .Z(n1100) );
INV_X1 U993 ( .A(G472), .ZN(n1189) );
NAND4_X1 U994 ( .A1(n1303), .A2(n1304), .A3(n1305), .A4(n1306), .ZN(n1302) );
NAND3_X1 U995 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1306) );
INV_X1 U996 ( .A(KEYINPUT58), .ZN(n1308) );
OR2_X1 U997 ( .A1(n1309), .A2(n1307), .ZN(n1305) );
NOR2_X1 U998 ( .A1(KEYINPUT23), .A2(n1310), .ZN(n1307) );
NAND2_X1 U999 ( .A1(n1311), .A2(n1312), .ZN(n1309) );
NAND2_X1 U1000 ( .A1(KEYINPUT0), .A2(n1313), .ZN(n1312) );
NAND2_X1 U1001 ( .A1(n1184), .A2(n1185), .ZN(n1313) );
NAND2_X1 U1002 ( .A1(n1314), .A2(n1315), .ZN(n1185) );
OR2_X1 U1003 ( .A1(n1315), .A2(n1314), .ZN(n1184) );
NAND2_X1 U1004 ( .A1(n1316), .A2(n1317), .ZN(n1311) );
INV_X1 U1005 ( .A(KEYINPUT0), .ZN(n1317) );
XOR2_X1 U1006 ( .A(n1315), .B(n1314), .Z(n1316) );
XOR2_X1 U1007 ( .A(n1318), .B(n1319), .Z(n1314) );
XNOR2_X1 U1008 ( .A(G113), .B(KEYINPUT49), .ZN(n1318) );
XNOR2_X1 U1009 ( .A(n1320), .B(n1321), .ZN(n1315) );
NAND2_X1 U1010 ( .A1(KEYINPUT58), .A2(n1310), .ZN(n1303) );
XNOR2_X1 U1011 ( .A(n1186), .B(n1182), .ZN(n1310) );
NAND2_X1 U1012 ( .A1(G210), .A2(n1322), .ZN(n1186) );
NOR2_X1 U1013 ( .A1(n1252), .A2(n1251), .ZN(n1065) );
XOR2_X1 U1014 ( .A(n1323), .B(n1164), .Z(n1251) );
INV_X1 U1015 ( .A(G475), .ZN(n1164) );
OR2_X1 U1016 ( .A1(n1163), .A2(G902), .ZN(n1323) );
XNOR2_X1 U1017 ( .A(n1324), .B(n1325), .ZN(n1163) );
XOR2_X1 U1018 ( .A(n1321), .B(n1326), .Z(n1325) );
XNOR2_X1 U1019 ( .A(n1327), .B(n1328), .ZN(n1326) );
NOR2_X1 U1020 ( .A1(G125), .A2(KEYINPUT2), .ZN(n1328) );
NAND2_X1 U1021 ( .A1(KEYINPUT56), .A2(n1261), .ZN(n1327) );
XOR2_X1 U1022 ( .A(n1329), .B(n1330), .Z(n1324) );
XNOR2_X1 U1023 ( .A(G140), .B(n1331), .ZN(n1330) );
NAND2_X1 U1024 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
XNOR2_X1 U1025 ( .A(G104), .B(n1334), .ZN(n1333) );
XNOR2_X1 U1026 ( .A(n1335), .B(G113), .ZN(n1334) );
XNOR2_X1 U1027 ( .A(KEYINPUT50), .B(KEYINPUT14), .ZN(n1332) );
NAND2_X1 U1028 ( .A1(G214), .A2(n1322), .ZN(n1329) );
NOR2_X1 U1029 ( .A1(G953), .A2(G237), .ZN(n1322) );
XOR2_X1 U1030 ( .A(n1336), .B(n1160), .Z(n1252) );
INV_X1 U1031 ( .A(G478), .ZN(n1160) );
NAND2_X1 U1032 ( .A1(n1158), .A2(n1304), .ZN(n1336) );
XNOR2_X1 U1033 ( .A(n1337), .B(n1338), .ZN(n1158) );
XOR2_X1 U1034 ( .A(G128), .B(n1339), .Z(n1338) );
XNOR2_X1 U1035 ( .A(n1340), .B(G134), .ZN(n1339) );
XOR2_X1 U1036 ( .A(n1341), .B(n1342), .Z(n1337) );
AND3_X1 U1037 ( .A1(G217), .A2(n1079), .A3(G234), .ZN(n1342) );
XNOR2_X1 U1038 ( .A(n1343), .B(n1344), .ZN(n1341) );
NAND3_X1 U1039 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1343) );
NAND2_X1 U1040 ( .A1(G116), .A2(n1348), .ZN(n1347) );
INV_X1 U1041 ( .A(KEYINPUT38), .ZN(n1348) );
NAND3_X1 U1042 ( .A1(KEYINPUT38), .A2(n1349), .A3(n1335), .ZN(n1346) );
OR2_X1 U1043 ( .A1(n1335), .A2(n1349), .ZN(n1345) );
NOR2_X1 U1044 ( .A1(G116), .A2(KEYINPUT28), .ZN(n1349) );
INV_X1 U1045 ( .A(G122), .ZN(n1335) );
AND3_X1 U1046 ( .A1(n1066), .A2(n1244), .A3(n1073), .ZN(n1175) );
NOR2_X1 U1047 ( .A1(n1090), .A2(n1091), .ZN(n1073) );
INV_X1 U1048 ( .A(n1262), .ZN(n1091) );
NAND2_X1 U1049 ( .A1(G214), .A2(n1350), .ZN(n1262) );
XOR2_X1 U1050 ( .A(n1351), .B(n1352), .Z(n1090) );
XNOR2_X1 U1051 ( .A(KEYINPUT1), .B(n1106), .ZN(n1352) );
NAND2_X1 U1052 ( .A1(n1353), .A2(n1304), .ZN(n1106) );
XNOR2_X1 U1053 ( .A(n1210), .B(n1206), .ZN(n1353) );
XNOR2_X1 U1054 ( .A(n1354), .B(n1355), .ZN(n1206) );
XNOR2_X1 U1055 ( .A(n1144), .B(n1143), .ZN(n1355) );
XNOR2_X1 U1056 ( .A(G113), .B(n1356), .ZN(n1143) );
NOR2_X1 U1057 ( .A1(KEYINPUT24), .A2(n1319), .ZN(n1356) );
XOR2_X1 U1058 ( .A(G116), .B(n1294), .Z(n1319) );
XOR2_X1 U1059 ( .A(G119), .B(KEYINPUT44), .Z(n1294) );
XNOR2_X1 U1060 ( .A(n1357), .B(G101), .ZN(n1144) );
NAND3_X1 U1061 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1357) );
NAND2_X1 U1062 ( .A1(n1344), .A2(n1361), .ZN(n1360) );
OR3_X1 U1063 ( .A1(n1361), .A2(n1344), .A3(n1362), .ZN(n1359) );
INV_X1 U1064 ( .A(KEYINPUT11), .ZN(n1361) );
NAND2_X1 U1065 ( .A1(n1362), .A2(n1363), .ZN(n1358) );
NAND2_X1 U1066 ( .A1(KEYINPUT11), .A2(n1364), .ZN(n1363) );
XNOR2_X1 U1067 ( .A(KEYINPUT36), .B(n1344), .ZN(n1364) );
XOR2_X1 U1068 ( .A(G104), .B(KEYINPUT46), .Z(n1362) );
XOR2_X1 U1069 ( .A(n1365), .B(KEYINPUT61), .Z(n1354) );
NAND2_X1 U1070 ( .A1(KEYINPUT34), .A2(n1140), .ZN(n1365) );
NAND3_X1 U1071 ( .A1(n1366), .A2(n1367), .A3(n1368), .ZN(n1140) );
NAND2_X1 U1072 ( .A1(KEYINPUT54), .A2(G110), .ZN(n1368) );
OR3_X1 U1073 ( .A1(n1369), .A2(KEYINPUT54), .A3(G122), .ZN(n1367) );
NAND2_X1 U1074 ( .A1(G122), .A2(n1369), .ZN(n1366) );
NAND2_X1 U1075 ( .A1(KEYINPUT35), .A2(n1201), .ZN(n1369) );
XOR2_X1 U1076 ( .A(n1370), .B(n1371), .Z(n1210) );
XNOR2_X1 U1077 ( .A(G128), .B(n1263), .ZN(n1371) );
INV_X1 U1078 ( .A(G125), .ZN(n1263) );
XOR2_X1 U1079 ( .A(n1372), .B(n1321), .Z(n1370) );
XNOR2_X1 U1080 ( .A(n1340), .B(G146), .ZN(n1321) );
INV_X1 U1081 ( .A(G143), .ZN(n1340) );
NAND2_X1 U1082 ( .A1(G224), .A2(n1079), .ZN(n1372) );
NAND2_X1 U1083 ( .A1(KEYINPUT51), .A2(n1105), .ZN(n1351) );
NAND2_X1 U1084 ( .A1(G210), .A2(n1350), .ZN(n1105) );
NAND2_X1 U1085 ( .A1(n1373), .A2(n1374), .ZN(n1350) );
INV_X1 U1086 ( .A(G237), .ZN(n1374) );
XNOR2_X1 U1087 ( .A(KEYINPUT29), .B(n1304), .ZN(n1373) );
NAND2_X1 U1088 ( .A1(n1375), .A2(n1376), .ZN(n1244) );
NAND3_X1 U1089 ( .A1(n1377), .A2(n1068), .A3(G952), .ZN(n1376) );
XNOR2_X1 U1090 ( .A(KEYINPUT5), .B(n1079), .ZN(n1377) );
XOR2_X1 U1091 ( .A(n1378), .B(KEYINPUT31), .Z(n1375) );
NAND4_X1 U1092 ( .A1(n1379), .A2(G953), .A3(G902), .A4(n1068), .ZN(n1378) );
NAND2_X1 U1093 ( .A1(G237), .A2(n1380), .ZN(n1068) );
XOR2_X1 U1094 ( .A(KEYINPUT3), .B(G234), .Z(n1380) );
XNOR2_X1 U1095 ( .A(G898), .B(KEYINPUT27), .ZN(n1379) );
NOR2_X1 U1096 ( .A1(n1381), .A2(n1084), .ZN(n1066) );
NOR2_X1 U1097 ( .A1(n1382), .A2(n1107), .ZN(n1084) );
NOR2_X1 U1098 ( .A1(n1108), .A2(G469), .ZN(n1107) );
AND2_X1 U1099 ( .A1(n1383), .A2(G469), .ZN(n1382) );
XOR2_X1 U1100 ( .A(n1108), .B(KEYINPUT52), .Z(n1383) );
NAND2_X1 U1101 ( .A1(n1384), .A2(n1304), .ZN(n1108) );
XOR2_X1 U1102 ( .A(n1385), .B(n1386), .Z(n1384) );
XNOR2_X1 U1103 ( .A(n1201), .B(n1387), .ZN(n1386) );
XNOR2_X1 U1104 ( .A(KEYINPUT17), .B(n1253), .ZN(n1387) );
INV_X1 U1105 ( .A(G140), .ZN(n1253) );
INV_X1 U1106 ( .A(G110), .ZN(n1201) );
XNOR2_X1 U1107 ( .A(n1191), .B(n1199), .ZN(n1385) );
AND2_X1 U1108 ( .A1(G227), .A2(n1079), .ZN(n1199) );
INV_X1 U1109 ( .A(G953), .ZN(n1079) );
XNOR2_X1 U1110 ( .A(n1388), .B(n1389), .ZN(n1191) );
XNOR2_X1 U1111 ( .A(n1169), .B(n1390), .ZN(n1389) );
XNOR2_X1 U1112 ( .A(KEYINPUT48), .B(n1344), .ZN(n1390) );
INV_X1 U1113 ( .A(G107), .ZN(n1344) );
INV_X1 U1114 ( .A(G104), .ZN(n1169) );
XNOR2_X1 U1115 ( .A(n1391), .B(n1392), .ZN(n1388) );
INV_X1 U1116 ( .A(n1126), .ZN(n1392) );
XOR2_X1 U1117 ( .A(G143), .B(n1393), .Z(n1126) );
NOR2_X1 U1118 ( .A1(G146), .A2(KEYINPUT37), .ZN(n1393) );
XNOR2_X1 U1119 ( .A(n1320), .B(n1182), .ZN(n1391) );
INV_X1 U1120 ( .A(G101), .ZN(n1182) );
XOR2_X1 U1121 ( .A(n1394), .B(n1128), .Z(n1320) );
XNOR2_X1 U1122 ( .A(n1261), .B(G128), .ZN(n1128) );
INV_X1 U1123 ( .A(G131), .ZN(n1261) );
NAND2_X1 U1124 ( .A1(KEYINPUT15), .A2(n1129), .ZN(n1394) );
XNOR2_X1 U1125 ( .A(n1260), .B(n1301), .ZN(n1129) );
INV_X1 U1126 ( .A(G137), .ZN(n1301) );
INV_X1 U1127 ( .A(G134), .ZN(n1260) );
INV_X1 U1128 ( .A(n1283), .ZN(n1381) );
XNOR2_X1 U1129 ( .A(n1086), .B(KEYINPUT45), .ZN(n1283) );
NAND2_X1 U1130 ( .A1(G221), .A2(n1291), .ZN(n1086) );
NAND2_X1 U1131 ( .A1(G234), .A2(n1304), .ZN(n1291) );
INV_X1 U1132 ( .A(G902), .ZN(n1304) );
endmodule


