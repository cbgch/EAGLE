//Key = 0001111001100111001110110101010111110001010000010110100001100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369;

XOR2_X1 U741 ( .A(n1037), .B(n1038), .Z(G9) );
NAND2_X1 U742 ( .A1(KEYINPUT47), .A2(G107), .ZN(n1038) );
NOR2_X1 U743 ( .A1(n1039), .A2(n1040), .ZN(G75) );
NOR3_X1 U744 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NAND3_X1 U745 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1041) );
NAND2_X1 U746 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U747 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND4_X1 U748 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1050) );
NOR3_X1 U749 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NAND2_X1 U750 ( .A1(n1058), .A2(n1059), .ZN(n1053) );
NAND3_X1 U751 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1052) );
NAND2_X1 U752 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U753 ( .A1(n1058), .A2(n1065), .ZN(n1064) );
INV_X1 U754 ( .A(n1066), .ZN(n1058) );
OR2_X1 U755 ( .A1(n1067), .A2(n1063), .ZN(n1051) );
NAND3_X1 U756 ( .A1(n1063), .A2(n1068), .A3(n1067), .ZN(n1049) );
NAND2_X1 U757 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U758 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NAND2_X1 U759 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
OR2_X1 U760 ( .A1(n1056), .A2(n1075), .ZN(n1074) );
INV_X1 U761 ( .A(n1076), .ZN(n1056) );
NAND2_X1 U762 ( .A1(n1077), .A2(n1078), .ZN(n1073) );
OR2_X1 U763 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
INV_X1 U764 ( .A(n1081), .ZN(n1047) );
NOR3_X1 U765 ( .A1(n1082), .A2(G953), .A3(G952), .ZN(n1039) );
INV_X1 U766 ( .A(n1044), .ZN(n1082) );
NAND4_X1 U767 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1044) );
NOR3_X1 U768 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NOR2_X1 U769 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U770 ( .A1(n1092), .A2(n1093), .ZN(n1088) );
NOR2_X1 U771 ( .A1(n1094), .A2(G469), .ZN(n1093) );
NOR2_X1 U772 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U773 ( .A1(n1097), .A2(KEYINPUT0), .ZN(n1095) );
NOR2_X1 U774 ( .A1(n1098), .A2(n1099), .ZN(n1092) );
NOR2_X1 U775 ( .A1(n1100), .A2(KEYINPUT0), .ZN(n1098) );
NOR2_X1 U776 ( .A1(n1101), .A2(n1096), .ZN(n1100) );
INV_X1 U777 ( .A(KEYINPUT23), .ZN(n1096) );
NAND3_X1 U778 ( .A1(n1065), .A2(n1075), .A3(n1102), .ZN(n1087) );
NOR3_X1 U779 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1085) );
XOR2_X1 U780 ( .A(n1106), .B(KEYINPUT3), .Z(n1105) );
XNOR2_X1 U781 ( .A(n1107), .B(KEYINPUT20), .ZN(n1104) );
XOR2_X1 U782 ( .A(n1108), .B(KEYINPUT38), .Z(n1083) );
NAND2_X1 U783 ( .A1(n1109), .A2(n1091), .ZN(n1108) );
XOR2_X1 U784 ( .A(KEYINPUT2), .B(n1090), .Z(n1109) );
XOR2_X1 U785 ( .A(n1110), .B(n1111), .Z(G72) );
XOR2_X1 U786 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND2_X1 U787 ( .A1(G953), .A2(n1114), .ZN(n1113) );
NAND2_X1 U788 ( .A1(G900), .A2(G227), .ZN(n1114) );
NAND2_X1 U789 ( .A1(n1115), .A2(n1116), .ZN(n1112) );
NAND2_X1 U790 ( .A1(G953), .A2(n1117), .ZN(n1116) );
XOR2_X1 U791 ( .A(n1118), .B(n1119), .Z(n1115) );
XOR2_X1 U792 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U793 ( .A1(KEYINPUT25), .A2(n1122), .ZN(n1121) );
NAND2_X1 U794 ( .A1(n1123), .A2(n1124), .ZN(n1120) );
NAND2_X1 U795 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XOR2_X1 U796 ( .A(n1127), .B(KEYINPUT11), .Z(n1123) );
OR2_X1 U797 ( .A1(n1125), .A2(n1126), .ZN(n1127) );
XNOR2_X1 U798 ( .A(n1128), .B(n1129), .ZN(n1125) );
XOR2_X1 U799 ( .A(G137), .B(G134), .Z(n1129) );
NAND2_X1 U800 ( .A1(KEYINPUT50), .A2(n1130), .ZN(n1128) );
XNOR2_X1 U801 ( .A(G125), .B(KEYINPUT31), .ZN(n1118) );
AND2_X1 U802 ( .A1(n1042), .A2(n1045), .ZN(n1110) );
XOR2_X1 U803 ( .A(n1131), .B(n1132), .Z(G69) );
XOR2_X1 U804 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U805 ( .A1(n1135), .A2(n1045), .ZN(n1134) );
NOR2_X1 U806 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XNOR2_X1 U807 ( .A(G224), .B(KEYINPUT7), .ZN(n1136) );
NAND2_X1 U808 ( .A1(n1138), .A2(n1139), .ZN(n1133) );
NAND2_X1 U809 ( .A1(G953), .A2(n1137), .ZN(n1139) );
XOR2_X1 U810 ( .A(n1140), .B(KEYINPUT32), .Z(n1138) );
NAND2_X1 U811 ( .A1(n1045), .A2(n1043), .ZN(n1131) );
NOR2_X1 U812 ( .A1(n1141), .A2(n1142), .ZN(G66) );
XOR2_X1 U813 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U814 ( .A1(n1145), .A2(n1090), .ZN(n1143) );
NOR2_X1 U815 ( .A1(n1141), .A2(n1146), .ZN(G63) );
XOR2_X1 U816 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U817 ( .A1(n1149), .A2(KEYINPUT59), .ZN(n1148) );
INV_X1 U818 ( .A(n1150), .ZN(n1149) );
AND2_X1 U819 ( .A1(G478), .A2(n1145), .ZN(n1147) );
NOR2_X1 U820 ( .A1(n1141), .A2(n1151), .ZN(G60) );
XOR2_X1 U821 ( .A(n1152), .B(n1153), .Z(n1151) );
AND2_X1 U822 ( .A1(G475), .A2(n1145), .ZN(n1153) );
NAND2_X1 U823 ( .A1(KEYINPUT18), .A2(n1154), .ZN(n1152) );
NAND2_X1 U824 ( .A1(n1155), .A2(n1156), .ZN(G6) );
NAND2_X1 U825 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND2_X1 U826 ( .A1(G104), .A2(n1159), .ZN(n1158) );
NAND2_X1 U827 ( .A1(KEYINPUT54), .A2(KEYINPUT15), .ZN(n1159) );
NAND3_X1 U828 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1155) );
INV_X1 U829 ( .A(KEYINPUT54), .ZN(n1162) );
OR2_X1 U830 ( .A1(n1163), .A2(KEYINPUT15), .ZN(n1161) );
NAND2_X1 U831 ( .A1(KEYINPUT15), .A2(n1164), .ZN(n1160) );
NAND2_X1 U832 ( .A1(G104), .A2(n1165), .ZN(n1164) );
NOR2_X1 U833 ( .A1(n1141), .A2(n1166), .ZN(G57) );
XOR2_X1 U834 ( .A(n1167), .B(n1168), .Z(n1166) );
XNOR2_X1 U835 ( .A(n1169), .B(n1170), .ZN(n1168) );
XOR2_X1 U836 ( .A(n1171), .B(n1172), .Z(n1167) );
NOR2_X1 U837 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U838 ( .A(n1175), .B(KEYINPUT9), .Z(n1174) );
NAND2_X1 U839 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NOR2_X1 U840 ( .A1(n1177), .A2(n1176), .ZN(n1173) );
XNOR2_X1 U841 ( .A(KEYINPUT5), .B(n1178), .ZN(n1176) );
NAND2_X1 U842 ( .A1(n1145), .A2(G472), .ZN(n1171) );
NOR2_X1 U843 ( .A1(n1141), .A2(n1179), .ZN(G54) );
XOR2_X1 U844 ( .A(n1180), .B(n1181), .Z(n1179) );
XNOR2_X1 U845 ( .A(n1182), .B(KEYINPUT63), .ZN(n1181) );
NAND2_X1 U846 ( .A1(KEYINPUT22), .A2(n1183), .ZN(n1182) );
XOR2_X1 U847 ( .A(n1184), .B(n1185), .Z(n1180) );
NAND2_X1 U848 ( .A1(n1145), .A2(G469), .ZN(n1184) );
NOR2_X1 U849 ( .A1(n1141), .A2(n1186), .ZN(G51) );
NOR2_X1 U850 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U851 ( .A(n1189), .B(KEYINPUT58), .Z(n1188) );
NAND2_X1 U852 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U853 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
XOR2_X1 U854 ( .A(n1192), .B(n1193), .Z(n1191) );
NAND2_X1 U855 ( .A1(n1194), .A2(n1195), .ZN(n1192) );
INV_X1 U856 ( .A(n1196), .ZN(n1195) );
NAND2_X1 U857 ( .A1(G125), .A2(n1197), .ZN(n1194) );
XNOR2_X1 U858 ( .A(n1198), .B(KEYINPUT56), .ZN(n1197) );
AND3_X1 U859 ( .A1(G210), .A2(n1199), .A3(n1145), .ZN(n1190) );
AND2_X1 U860 ( .A1(G902), .A2(n1200), .ZN(n1145) );
OR2_X1 U861 ( .A1(n1043), .A2(n1042), .ZN(n1200) );
NAND4_X1 U862 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1042) );
NOR4_X1 U863 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
NOR2_X1 U864 ( .A1(n1209), .A2(n1210), .ZN(n1203) );
NAND4_X1 U865 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1043) );
AND4_X1 U866 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
NOR3_X1 U867 ( .A1(n1157), .A2(n1219), .A3(n1220), .ZN(n1213) );
NOR2_X1 U868 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
OR4_X1 U869 ( .A1(n1223), .A2(n1070), .A3(n1060), .A4(n1224), .ZN(n1222) );
INV_X1 U870 ( .A(n1225), .ZN(n1060) );
NAND2_X1 U871 ( .A1(n1076), .A2(n1226), .ZN(n1070) );
INV_X1 U872 ( .A(KEYINPUT44), .ZN(n1221) );
NOR2_X1 U873 ( .A1(KEYINPUT44), .A2(n1037), .ZN(n1219) );
NAND3_X1 U874 ( .A1(n1225), .A2(n1076), .A3(n1227), .ZN(n1037) );
INV_X1 U875 ( .A(n1165), .ZN(n1157) );
NAND3_X1 U876 ( .A1(n1227), .A2(n1076), .A3(n1228), .ZN(n1165) );
NOR2_X1 U877 ( .A1(n1045), .A2(G952), .ZN(n1141) );
NAND3_X1 U878 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(G48) );
OR2_X1 U879 ( .A1(n1232), .A2(G146), .ZN(n1231) );
NAND3_X1 U880 ( .A1(G146), .A2(n1232), .A3(n1201), .ZN(n1230) );
NAND2_X1 U881 ( .A1(n1233), .A2(n1234), .ZN(n1229) );
NAND2_X1 U882 ( .A1(n1235), .A2(n1232), .ZN(n1234) );
INV_X1 U883 ( .A(KEYINPUT17), .ZN(n1232) );
XOR2_X1 U884 ( .A(KEYINPUT28), .B(G146), .Z(n1235) );
INV_X1 U885 ( .A(n1201), .ZN(n1233) );
NAND3_X1 U886 ( .A1(n1236), .A2(n1066), .A3(n1237), .ZN(n1201) );
XNOR2_X1 U887 ( .A(G143), .B(n1238), .ZN(G45) );
NOR2_X1 U888 ( .A1(n1210), .A2(KEYINPUT43), .ZN(n1238) );
AND4_X1 U889 ( .A1(n1103), .A2(n1239), .A3(n1107), .A4(n1240), .ZN(n1210) );
AND3_X1 U890 ( .A1(n1080), .A2(n1066), .A3(n1226), .ZN(n1240) );
XNOR2_X1 U891 ( .A(n1122), .B(n1209), .ZN(G42) );
AND3_X1 U892 ( .A1(n1228), .A2(n1079), .A3(n1241), .ZN(n1209) );
XOR2_X1 U893 ( .A(G137), .B(n1208), .Z(G39) );
AND3_X1 U894 ( .A1(n1063), .A2(n1236), .A3(n1241), .ZN(n1208) );
XOR2_X1 U895 ( .A(G134), .B(n1207), .Z(G36) );
AND3_X1 U896 ( .A1(n1080), .A2(n1225), .A3(n1241), .ZN(n1207) );
XNOR2_X1 U897 ( .A(n1130), .B(n1206), .ZN(G33) );
AND3_X1 U898 ( .A1(n1080), .A2(n1228), .A3(n1241), .ZN(n1206) );
AND4_X1 U899 ( .A1(n1077), .A2(n1071), .A3(n1066), .A4(n1239), .ZN(n1241) );
XOR2_X1 U900 ( .A(n1242), .B(KEYINPUT30), .Z(n1066) );
INV_X1 U901 ( .A(n1057), .ZN(n1077) );
INV_X1 U902 ( .A(G131), .ZN(n1130) );
NAND2_X1 U903 ( .A1(n1243), .A2(n1244), .ZN(G30) );
NAND2_X1 U904 ( .A1(n1205), .A2(n1245), .ZN(n1244) );
XOR2_X1 U905 ( .A(KEYINPUT10), .B(n1246), .Z(n1243) );
NOR2_X1 U906 ( .A1(n1205), .A2(n1245), .ZN(n1246) );
AND3_X1 U907 ( .A1(n1225), .A2(n1242), .A3(n1247), .ZN(n1205) );
AND3_X1 U908 ( .A1(n1226), .A2(n1239), .A3(n1236), .ZN(n1247) );
XNOR2_X1 U909 ( .A(n1248), .B(n1211), .ZN(G3) );
NAND3_X1 U910 ( .A1(n1063), .A2(n1227), .A3(n1080), .ZN(n1211) );
NOR2_X1 U911 ( .A1(KEYINPUT53), .A2(n1249), .ZN(n1248) );
XNOR2_X1 U912 ( .A(G101), .B(KEYINPUT55), .ZN(n1249) );
XNOR2_X1 U913 ( .A(G125), .B(n1202), .ZN(G27) );
NAND3_X1 U914 ( .A1(n1067), .A2(n1079), .A3(n1237), .ZN(n1202) );
AND3_X1 U915 ( .A1(n1226), .A2(n1239), .A3(n1228), .ZN(n1237) );
NAND2_X1 U916 ( .A1(n1250), .A2(n1081), .ZN(n1239) );
NAND4_X1 U917 ( .A1(G953), .A2(G902), .A3(n1251), .A4(n1117), .ZN(n1250) );
INV_X1 U918 ( .A(G900), .ZN(n1117) );
XNOR2_X1 U919 ( .A(G122), .B(n1212), .ZN(G24) );
NAND4_X1 U920 ( .A1(n1252), .A2(n1076), .A3(n1107), .A4(n1103), .ZN(n1212) );
XNOR2_X1 U921 ( .A(G119), .B(n1218), .ZN(G21) );
NAND3_X1 U922 ( .A1(n1063), .A2(n1236), .A3(n1252), .ZN(n1218) );
NAND2_X1 U923 ( .A1(n1253), .A2(n1254), .ZN(n1236) );
NAND2_X1 U924 ( .A1(n1080), .A2(n1255), .ZN(n1254) );
NAND3_X1 U925 ( .A1(n1256), .A2(n1257), .A3(KEYINPUT33), .ZN(n1253) );
XNOR2_X1 U926 ( .A(G116), .B(n1217), .ZN(G18) );
NAND3_X1 U927 ( .A1(n1252), .A2(n1225), .A3(n1080), .ZN(n1217) );
NOR2_X1 U928 ( .A1(n1103), .A2(n1258), .ZN(n1225) );
XNOR2_X1 U929 ( .A(G113), .B(n1216), .ZN(G15) );
NAND3_X1 U930 ( .A1(n1228), .A2(n1252), .A3(n1080), .ZN(n1216) );
NOR2_X1 U931 ( .A1(n1256), .A2(n1084), .ZN(n1080) );
AND3_X1 U932 ( .A1(n1226), .A2(n1223), .A3(n1067), .ZN(n1252) );
NOR2_X1 U933 ( .A1(n1059), .A2(n1259), .ZN(n1067) );
INV_X1 U934 ( .A(n1065), .ZN(n1259) );
INV_X1 U935 ( .A(n1061), .ZN(n1228) );
NAND2_X1 U936 ( .A1(n1258), .A2(n1103), .ZN(n1061) );
INV_X1 U937 ( .A(n1107), .ZN(n1258) );
XNOR2_X1 U938 ( .A(G110), .B(n1215), .ZN(G12) );
NAND3_X1 U939 ( .A1(n1227), .A2(n1079), .A3(n1063), .ZN(n1215) );
NOR2_X1 U940 ( .A1(n1107), .A2(n1103), .ZN(n1063) );
XNOR2_X1 U941 ( .A(n1260), .B(G475), .ZN(n1103) );
NAND2_X1 U942 ( .A1(n1154), .A2(n1261), .ZN(n1260) );
XNOR2_X1 U943 ( .A(n1262), .B(n1263), .ZN(n1154) );
XOR2_X1 U944 ( .A(n1264), .B(n1265), .Z(n1263) );
NAND2_X1 U945 ( .A1(KEYINPUT13), .A2(G104), .ZN(n1265) );
NAND2_X1 U946 ( .A1(n1266), .A2(n1267), .ZN(n1264) );
NAND2_X1 U947 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XOR2_X1 U948 ( .A(KEYINPUT6), .B(n1270), .Z(n1266) );
NOR2_X1 U949 ( .A1(n1269), .A2(n1268), .ZN(n1270) );
XOR2_X1 U950 ( .A(n1271), .B(n1272), .Z(n1268) );
XOR2_X1 U951 ( .A(n1273), .B(G125), .Z(n1271) );
NAND2_X1 U952 ( .A1(KEYINPUT35), .A2(n1122), .ZN(n1273) );
XOR2_X1 U953 ( .A(n1274), .B(n1275), .Z(n1269) );
XNOR2_X1 U954 ( .A(n1276), .B(G131), .ZN(n1275) );
NAND2_X1 U955 ( .A1(n1277), .A2(G214), .ZN(n1274) );
XNOR2_X1 U956 ( .A(G113), .B(G122), .ZN(n1262) );
XOR2_X1 U957 ( .A(G478), .B(n1278), .Z(n1107) );
NOR2_X1 U958 ( .A1(G902), .A2(n1150), .ZN(n1278) );
NAND3_X1 U959 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1150) );
NAND2_X1 U960 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
INV_X1 U961 ( .A(KEYINPUT49), .ZN(n1283) );
NAND3_X1 U962 ( .A1(KEYINPUT49), .A2(n1284), .A3(n1285), .ZN(n1280) );
OR2_X1 U963 ( .A1(n1285), .A2(n1284), .ZN(n1279) );
NOR2_X1 U964 ( .A1(n1286), .A2(n1282), .ZN(n1284) );
NAND3_X1 U965 ( .A1(G234), .A2(n1045), .A3(G217), .ZN(n1282) );
INV_X1 U966 ( .A(KEYINPUT19), .ZN(n1286) );
XNOR2_X1 U967 ( .A(n1287), .B(n1288), .ZN(n1285) );
XOR2_X1 U968 ( .A(G116), .B(n1289), .Z(n1288) );
XNOR2_X1 U969 ( .A(G134), .B(n1290), .ZN(n1289) );
INV_X1 U970 ( .A(G122), .ZN(n1290) );
XNOR2_X1 U971 ( .A(G107), .B(n1291), .ZN(n1287) );
NAND2_X1 U972 ( .A1(n1292), .A2(n1293), .ZN(n1079) );
NAND2_X1 U973 ( .A1(n1076), .A2(n1255), .ZN(n1293) );
INV_X1 U974 ( .A(KEYINPUT33), .ZN(n1255) );
NOR2_X1 U975 ( .A1(n1257), .A2(n1256), .ZN(n1076) );
NAND3_X1 U976 ( .A1(n1256), .A2(n1084), .A3(KEYINPUT33), .ZN(n1292) );
INV_X1 U977 ( .A(n1257), .ZN(n1084) );
XNOR2_X1 U978 ( .A(n1294), .B(G472), .ZN(n1257) );
NAND2_X1 U979 ( .A1(n1295), .A2(n1261), .ZN(n1294) );
XNOR2_X1 U980 ( .A(n1296), .B(n1297), .ZN(n1295) );
XOR2_X1 U981 ( .A(n1178), .B(n1298), .Z(n1297) );
NAND2_X1 U982 ( .A1(n1277), .A2(G210), .ZN(n1178) );
NOR2_X1 U983 ( .A1(G953), .A2(G237), .ZN(n1277) );
INV_X1 U984 ( .A(n1169), .ZN(n1296) );
XNOR2_X1 U985 ( .A(n1299), .B(n1300), .ZN(n1169) );
XNOR2_X1 U986 ( .A(n1091), .B(n1090), .ZN(n1256) );
AND2_X1 U987 ( .A1(G217), .A2(n1301), .ZN(n1090) );
NAND2_X1 U988 ( .A1(n1144), .A2(n1302), .ZN(n1091) );
XNOR2_X1 U989 ( .A(KEYINPUT29), .B(n1261), .ZN(n1302) );
XOR2_X1 U990 ( .A(n1303), .B(n1304), .Z(n1144) );
XOR2_X1 U991 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U992 ( .A(KEYINPUT46), .B(G137), .Z(n1306) );
NOR2_X1 U993 ( .A1(n1307), .A2(n1308), .ZN(n1305) );
XOR2_X1 U994 ( .A(n1309), .B(KEYINPUT14), .Z(n1308) );
NAND2_X1 U995 ( .A1(G128), .A2(n1310), .ZN(n1309) );
XNOR2_X1 U996 ( .A(KEYINPUT34), .B(n1311), .ZN(n1310) );
NOR2_X1 U997 ( .A1(G128), .A2(n1311), .ZN(n1307) );
XOR2_X1 U998 ( .A(n1312), .B(n1313), .Z(n1303) );
XOR2_X1 U999 ( .A(n1314), .B(n1315), .Z(n1313) );
NAND2_X1 U1000 ( .A1(KEYINPUT62), .A2(n1183), .ZN(n1315) );
NAND2_X1 U1001 ( .A1(n1316), .A2(n1317), .ZN(n1314) );
NAND2_X1 U1002 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
XNOR2_X1 U1003 ( .A(G140), .B(n1320), .ZN(n1319) );
XNOR2_X1 U1004 ( .A(KEYINPUT40), .B(n1272), .ZN(n1318) );
XOR2_X1 U1005 ( .A(n1321), .B(KEYINPUT51), .Z(n1316) );
NAND2_X1 U1006 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XNOR2_X1 U1007 ( .A(n1122), .B(n1320), .ZN(n1323) );
NOR2_X1 U1008 ( .A1(G125), .A2(KEYINPUT12), .ZN(n1320) );
XOR2_X1 U1009 ( .A(KEYINPUT40), .B(n1272), .Z(n1322) );
NAND3_X1 U1010 ( .A1(G234), .A2(n1045), .A3(G221), .ZN(n1312) );
AND3_X1 U1011 ( .A1(n1226), .A2(n1223), .A3(n1242), .ZN(n1227) );
INV_X1 U1012 ( .A(n1224), .ZN(n1242) );
NAND2_X1 U1013 ( .A1(n1059), .A2(n1065), .ZN(n1224) );
NAND2_X1 U1014 ( .A1(G221), .A2(n1301), .ZN(n1065) );
NAND2_X1 U1015 ( .A1(G234), .A2(n1324), .ZN(n1301) );
XNOR2_X1 U1016 ( .A(n1097), .B(n1101), .ZN(n1059) );
INV_X1 U1017 ( .A(G469), .ZN(n1101) );
INV_X1 U1018 ( .A(n1099), .ZN(n1097) );
NAND2_X1 U1019 ( .A1(n1325), .A2(n1261), .ZN(n1099) );
XOR2_X1 U1020 ( .A(n1185), .B(n1326), .Z(n1325) );
XOR2_X1 U1021 ( .A(KEYINPUT4), .B(n1183), .Z(n1326) );
XNOR2_X1 U1022 ( .A(n1327), .B(n1328), .ZN(n1185) );
XNOR2_X1 U1023 ( .A(n1299), .B(n1126), .ZN(n1328) );
XOR2_X1 U1024 ( .A(n1291), .B(n1329), .Z(n1126) );
XOR2_X1 U1025 ( .A(KEYINPUT60), .B(n1272), .Z(n1329) );
XNOR2_X1 U1026 ( .A(G143), .B(n1245), .ZN(n1291) );
INV_X1 U1027 ( .A(G128), .ZN(n1245) );
XOR2_X1 U1028 ( .A(n1330), .B(n1331), .Z(n1299) );
NOR2_X1 U1029 ( .A1(KEYINPUT36), .A2(G134), .ZN(n1331) );
XNOR2_X1 U1030 ( .A(G131), .B(G137), .ZN(n1330) );
XOR2_X1 U1031 ( .A(n1332), .B(n1333), .Z(n1327) );
AND2_X1 U1032 ( .A1(n1045), .A2(G227), .ZN(n1333) );
XNOR2_X1 U1033 ( .A(n1334), .B(n1122), .ZN(n1332) );
INV_X1 U1034 ( .A(G140), .ZN(n1122) );
NAND3_X1 U1035 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1334) );
OR2_X1 U1036 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
NAND3_X1 U1037 ( .A1(n1340), .A2(n1338), .A3(n1177), .ZN(n1336) );
INV_X1 U1038 ( .A(KEYINPUT24), .ZN(n1338) );
OR2_X1 U1039 ( .A1(n1177), .A2(n1340), .ZN(n1335) );
AND2_X1 U1040 ( .A1(KEYINPUT61), .A2(n1339), .ZN(n1340) );
XNOR2_X1 U1041 ( .A(n1341), .B(n1342), .ZN(n1339) );
NOR2_X1 U1042 ( .A1(KEYINPUT8), .A2(n1163), .ZN(n1342) );
XNOR2_X1 U1043 ( .A(G107), .B(KEYINPUT48), .ZN(n1341) );
NAND2_X1 U1044 ( .A1(n1081), .A2(n1343), .ZN(n1223) );
NAND4_X1 U1045 ( .A1(G953), .A2(G902), .A3(n1251), .A4(n1137), .ZN(n1343) );
INV_X1 U1046 ( .A(G898), .ZN(n1137) );
NAND3_X1 U1047 ( .A1(n1251), .A2(n1045), .A3(G952), .ZN(n1081) );
NAND2_X1 U1048 ( .A1(G237), .A2(G234), .ZN(n1251) );
NOR2_X1 U1049 ( .A1(n1057), .A2(n1071), .ZN(n1226) );
INV_X1 U1050 ( .A(n1055), .ZN(n1071) );
NAND2_X1 U1051 ( .A1(n1102), .A2(n1106), .ZN(n1055) );
NAND3_X1 U1052 ( .A1(n1344), .A2(n1261), .A3(n1345), .ZN(n1106) );
NAND2_X1 U1053 ( .A1(G210), .A2(n1199), .ZN(n1345) );
NAND3_X1 U1054 ( .A1(n1346), .A2(n1199), .A3(G210), .ZN(n1102) );
NAND2_X1 U1055 ( .A1(n1344), .A2(n1261), .ZN(n1346) );
INV_X1 U1056 ( .A(G902), .ZN(n1261) );
NAND3_X1 U1057 ( .A1(n1347), .A2(n1348), .A3(n1349), .ZN(n1344) );
NAND2_X1 U1058 ( .A1(n1196), .A2(n1193), .ZN(n1349) );
NOR2_X1 U1059 ( .A1(n1350), .A2(G125), .ZN(n1196) );
OR3_X1 U1060 ( .A1(n1198), .A2(n1193), .A3(G125), .ZN(n1348) );
NAND2_X1 U1061 ( .A1(n1351), .A2(G125), .ZN(n1347) );
XNOR2_X1 U1062 ( .A(n1193), .B(n1350), .ZN(n1351) );
INV_X1 U1063 ( .A(n1198), .ZN(n1350) );
XNOR2_X1 U1064 ( .A(n1352), .B(n1300), .ZN(n1198) );
XNOR2_X1 U1065 ( .A(n1353), .B(G128), .ZN(n1300) );
NAND2_X1 U1066 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NAND3_X1 U1067 ( .A1(G143), .A2(n1272), .A3(n1356), .ZN(n1355) );
INV_X1 U1068 ( .A(KEYINPUT52), .ZN(n1356) );
NAND2_X1 U1069 ( .A1(n1357), .A2(KEYINPUT52), .ZN(n1354) );
XNOR2_X1 U1070 ( .A(n1276), .B(n1272), .ZN(n1357) );
XOR2_X1 U1071 ( .A(G146), .B(KEYINPUT27), .Z(n1272) );
INV_X1 U1072 ( .A(G143), .ZN(n1276) );
NAND2_X1 U1073 ( .A1(G224), .A2(n1045), .ZN(n1352) );
INV_X1 U1074 ( .A(G953), .ZN(n1045) );
XNOR2_X1 U1075 ( .A(n1140), .B(KEYINPUT26), .ZN(n1193) );
XOR2_X1 U1076 ( .A(n1358), .B(n1359), .Z(n1140) );
XNOR2_X1 U1077 ( .A(G122), .B(n1360), .ZN(n1359) );
XNOR2_X1 U1078 ( .A(KEYINPUT41), .B(KEYINPUT21), .ZN(n1360) );
XOR2_X1 U1079 ( .A(n1298), .B(n1361), .Z(n1358) );
XNOR2_X1 U1080 ( .A(n1362), .B(n1183), .ZN(n1361) );
XOR2_X1 U1081 ( .A(G110), .B(KEYINPUT37), .Z(n1183) );
NAND2_X1 U1082 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
NAND2_X1 U1083 ( .A1(G107), .A2(n1163), .ZN(n1364) );
XOR2_X1 U1084 ( .A(KEYINPUT57), .B(n1365), .Z(n1363) );
NOR2_X1 U1085 ( .A1(G107), .A2(n1163), .ZN(n1365) );
INV_X1 U1086 ( .A(G104), .ZN(n1163) );
XNOR2_X1 U1087 ( .A(n1177), .B(n1170), .ZN(n1298) );
XNOR2_X1 U1088 ( .A(n1366), .B(n1367), .ZN(n1170) );
XNOR2_X1 U1089 ( .A(KEYINPUT16), .B(n1311), .ZN(n1367) );
INV_X1 U1090 ( .A(G119), .ZN(n1311) );
XNOR2_X1 U1091 ( .A(G113), .B(G116), .ZN(n1366) );
XOR2_X1 U1092 ( .A(G101), .B(KEYINPUT39), .Z(n1177) );
XNOR2_X1 U1093 ( .A(n1075), .B(KEYINPUT45), .ZN(n1057) );
NAND2_X1 U1094 ( .A1(G214), .A2(n1199), .ZN(n1075) );
NAND2_X1 U1095 ( .A1(n1368), .A2(n1369), .ZN(n1199) );
INV_X1 U1096 ( .A(G237), .ZN(n1369) );
XOR2_X1 U1097 ( .A(n1324), .B(KEYINPUT1), .Z(n1368) );
XNOR2_X1 U1098 ( .A(G902), .B(KEYINPUT42), .ZN(n1324) );
endmodule


