//Key = 1010101110011101111011011111111100010011011101101110110110110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377;

XNOR2_X1 U746 ( .A(G107), .B(n1043), .ZN(G9) );
NOR2_X1 U747 ( .A1(n1044), .A2(n1045), .ZN(G75) );
NOR4_X1 U748 ( .A1(G953), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1045) );
NOR2_X1 U749 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR3_X1 U751 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NOR2_X1 U752 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U753 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U754 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U755 ( .A1(n1062), .A2(n1063), .ZN(n1056) );
NOR2_X1 U756 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U757 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR3_X1 U758 ( .A1(n1063), .A2(n1068), .A3(n1059), .ZN(n1051) );
NOR3_X1 U759 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1068) );
NOR2_X1 U760 ( .A1(n1072), .A2(n1053), .ZN(n1071) );
NOR2_X1 U761 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U762 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NOR3_X1 U763 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1070) );
XOR2_X1 U764 ( .A(KEYINPUT28), .B(n1080), .Z(n1077) );
NOR2_X1 U765 ( .A1(n1081), .A2(n1055), .ZN(n1069) );
NOR3_X1 U766 ( .A1(n1046), .A2(G953), .A3(G952), .ZN(n1044) );
AND4_X1 U767 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1046) );
NOR4_X1 U768 ( .A1(n1086), .A2(n1075), .A3(n1087), .A4(n1088), .ZN(n1085) );
XOR2_X1 U769 ( .A(n1089), .B(KEYINPUT17), .Z(n1088) );
XNOR2_X1 U770 ( .A(n1090), .B(n1091), .ZN(n1087) );
NOR2_X1 U771 ( .A1(G475), .A2(KEYINPUT62), .ZN(n1091) );
INV_X1 U772 ( .A(n1092), .ZN(n1086) );
XOR2_X1 U773 ( .A(n1093), .B(n1094), .Z(n1083) );
XOR2_X1 U774 ( .A(n1095), .B(KEYINPUT11), .Z(n1094) );
NAND2_X1 U775 ( .A1(n1096), .A2(n1097), .ZN(G72) );
NAND2_X1 U776 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
INV_X1 U777 ( .A(n1100), .ZN(n1098) );
NAND2_X1 U778 ( .A1(n1100), .A2(n1101), .ZN(n1096) );
NAND2_X1 U779 ( .A1(n1102), .A2(n1099), .ZN(n1101) );
NAND2_X1 U780 ( .A1(G953), .A2(n1103), .ZN(n1099) );
INV_X1 U781 ( .A(G227), .ZN(n1103) );
XOR2_X1 U782 ( .A(n1104), .B(n1105), .Z(n1100) );
NOR2_X1 U783 ( .A1(n1106), .A2(G953), .ZN(n1105) );
NOR2_X1 U784 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U785 ( .A(KEYINPUT45), .B(n1109), .ZN(n1108) );
NAND2_X1 U786 ( .A1(n1110), .A2(n1102), .ZN(n1104) );
INV_X1 U787 ( .A(n1111), .ZN(n1102) );
XOR2_X1 U788 ( .A(n1112), .B(n1113), .Z(n1110) );
XOR2_X1 U789 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U790 ( .A1(KEYINPUT9), .A2(n1116), .ZN(n1115) );
NOR2_X1 U791 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
XOR2_X1 U792 ( .A(KEYINPUT44), .B(n1119), .Z(n1118) );
AND2_X1 U793 ( .A1(n1120), .A2(G125), .ZN(n1119) );
NOR2_X1 U794 ( .A1(G125), .A2(n1120), .ZN(n1117) );
XOR2_X1 U795 ( .A(n1121), .B(n1122), .Z(G69) );
XOR2_X1 U796 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U797 ( .A1(G953), .A2(n1125), .ZN(n1124) );
NOR2_X1 U798 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U799 ( .A1(n1128), .A2(n1129), .ZN(n1123) );
NAND2_X1 U800 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U801 ( .A(KEYINPUT36), .B(G953), .Z(n1130) );
XOR2_X1 U802 ( .A(n1132), .B(n1133), .Z(n1128) );
XOR2_X1 U803 ( .A(KEYINPUT51), .B(n1134), .Z(n1133) );
NOR2_X1 U804 ( .A1(KEYINPUT40), .A2(n1135), .ZN(n1134) );
XOR2_X1 U805 ( .A(n1136), .B(n1137), .Z(n1132) );
NAND2_X1 U806 ( .A1(KEYINPUT59), .A2(n1138), .ZN(n1136) );
NAND2_X1 U807 ( .A1(G953), .A2(n1139), .ZN(n1121) );
NAND2_X1 U808 ( .A1(G898), .A2(G224), .ZN(n1139) );
NOR2_X1 U809 ( .A1(n1140), .A2(n1141), .ZN(G66) );
NOR3_X1 U810 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1141) );
NOR3_X1 U811 ( .A1(n1145), .A2(n1093), .A3(n1146), .ZN(n1144) );
NOR2_X1 U812 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
NOR2_X1 U813 ( .A1(n1149), .A2(n1093), .ZN(n1147) );
NOR2_X1 U814 ( .A1(n1140), .A2(n1150), .ZN(G63) );
NOR2_X1 U815 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U816 ( .A(n1153), .B(n1154), .Z(n1152) );
AND2_X1 U817 ( .A1(n1155), .A2(KEYINPUT0), .ZN(n1154) );
NOR2_X1 U818 ( .A1(n1156), .A2(n1146), .ZN(n1153) );
NOR2_X1 U819 ( .A1(KEYINPUT0), .A2(n1155), .ZN(n1151) );
NOR2_X1 U820 ( .A1(n1140), .A2(n1157), .ZN(G60) );
NOR3_X1 U821 ( .A1(n1090), .A2(n1158), .A3(n1159), .ZN(n1157) );
AND3_X1 U822 ( .A1(n1160), .A2(G475), .A3(n1161), .ZN(n1159) );
NOR2_X1 U823 ( .A1(n1162), .A2(n1160), .ZN(n1158) );
AND2_X1 U824 ( .A1(n1048), .A2(G475), .ZN(n1162) );
NAND2_X1 U825 ( .A1(n1163), .A2(n1164), .ZN(G6) );
NAND2_X1 U826 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XOR2_X1 U827 ( .A(KEYINPUT48), .B(n1167), .Z(n1163) );
NOR2_X1 U828 ( .A1(n1165), .A2(n1166), .ZN(n1167) );
INV_X1 U829 ( .A(n1168), .ZN(n1165) );
NOR2_X1 U830 ( .A1(n1140), .A2(n1169), .ZN(G57) );
NOR2_X1 U831 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U832 ( .A(n1172), .B(KEYINPUT30), .Z(n1171) );
NAND2_X1 U833 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
OR2_X1 U834 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NOR3_X1 U835 ( .A1(n1175), .A2(n1176), .A3(n1173), .ZN(n1170) );
AND2_X1 U836 ( .A1(n1177), .A2(n1178), .ZN(n1173) );
NAND2_X1 U837 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XNOR2_X1 U838 ( .A(n1181), .B(n1182), .ZN(n1179) );
NAND2_X1 U839 ( .A1(n1183), .A2(n1184), .ZN(n1177) );
XOR2_X1 U840 ( .A(KEYINPUT13), .B(n1180), .Z(n1184) );
AND2_X1 U841 ( .A1(n1161), .A2(G472), .ZN(n1180) );
XOR2_X1 U842 ( .A(n1182), .B(n1181), .Z(n1183) );
NAND2_X1 U843 ( .A1(KEYINPUT12), .A2(n1185), .ZN(n1182) );
AND2_X1 U844 ( .A1(n1186), .A2(n1187), .ZN(n1176) );
NOR2_X1 U845 ( .A1(n1186), .A2(n1187), .ZN(n1175) );
NOR2_X1 U846 ( .A1(n1140), .A2(n1188), .ZN(G54) );
XOR2_X1 U847 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U848 ( .A(n1191), .B(n1192), .Z(n1190) );
AND2_X1 U849 ( .A1(G469), .A2(n1161), .ZN(n1191) );
INV_X1 U850 ( .A(n1146), .ZN(n1161) );
XOR2_X1 U851 ( .A(n1193), .B(KEYINPUT50), .Z(n1189) );
NAND2_X1 U852 ( .A1(KEYINPUT53), .A2(n1194), .ZN(n1193) );
NAND2_X1 U853 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NAND3_X1 U854 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1196) );
XOR2_X1 U855 ( .A(KEYINPUT58), .B(n1200), .Z(n1195) );
NOR2_X1 U856 ( .A1(n1201), .A2(n1199), .ZN(n1200) );
AND2_X1 U857 ( .A1(n1198), .A2(n1197), .ZN(n1201) );
NAND2_X1 U858 ( .A1(n1202), .A2(n1203), .ZN(n1197) );
XOR2_X1 U859 ( .A(KEYINPUT27), .B(n1204), .Z(n1203) );
NOR2_X1 U860 ( .A1(n1205), .A2(n1206), .ZN(G51) );
XOR2_X1 U861 ( .A(n1207), .B(n1208), .Z(n1206) );
XOR2_X1 U862 ( .A(n1209), .B(n1210), .Z(n1208) );
XOR2_X1 U863 ( .A(G125), .B(n1211), .Z(n1207) );
NOR2_X1 U864 ( .A1(n1212), .A2(n1146), .ZN(n1211) );
NAND2_X1 U865 ( .A1(G902), .A2(n1048), .ZN(n1146) );
INV_X1 U866 ( .A(n1149), .ZN(n1048) );
NOR4_X1 U867 ( .A1(n1213), .A2(n1109), .A3(n1107), .A4(n1127), .ZN(n1149) );
NAND4_X1 U868 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1127) );
NAND2_X1 U869 ( .A1(n1218), .A2(n1065), .ZN(n1214) );
NAND4_X1 U870 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1107) );
NAND3_X1 U871 ( .A1(n1223), .A2(n1224), .A3(n1075), .ZN(n1221) );
XOR2_X1 U872 ( .A(KEYINPUT47), .B(n1225), .Z(n1224) );
NAND3_X1 U873 ( .A1(n1065), .A2(n1225), .A3(n1226), .ZN(n1220) );
INV_X1 U874 ( .A(n1227), .ZN(n1226) );
NAND2_X1 U875 ( .A1(n1082), .A2(n1228), .ZN(n1219) );
XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n1229), .ZN(n1228) );
NAND4_X1 U877 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1109) );
XNOR2_X1 U878 ( .A(n1126), .B(KEYINPUT18), .ZN(n1213) );
NAND4_X1 U879 ( .A1(n1168), .A2(n1234), .A3(n1235), .A4(n1043), .ZN(n1126) );
NAND3_X1 U880 ( .A1(n1060), .A2(n1080), .A3(n1236), .ZN(n1043) );
NAND3_X1 U881 ( .A1(n1236), .A2(n1080), .A3(n1061), .ZN(n1168) );
XNOR2_X1 U882 ( .A(n1140), .B(KEYINPUT35), .ZN(n1205) );
NOR2_X1 U883 ( .A1(n1237), .A2(G952), .ZN(n1140) );
XNOR2_X1 U884 ( .A(G146), .B(n1238), .ZN(G48) );
NAND4_X1 U885 ( .A1(n1075), .A2(KEYINPUT7), .A3(n1223), .A4(n1225), .ZN(n1238) );
XOR2_X1 U886 ( .A(G143), .B(n1239), .Z(G45) );
NOR3_X1 U887 ( .A1(n1240), .A2(n1227), .A3(n1241), .ZN(n1239) );
XOR2_X1 U888 ( .A(KEYINPUT26), .B(n1225), .Z(n1241) );
NAND4_X1 U889 ( .A1(n1074), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1227) );
XOR2_X1 U890 ( .A(KEYINPUT23), .B(n1065), .Z(n1240) );
XOR2_X1 U891 ( .A(n1120), .B(n1222), .Z(G42) );
NAND4_X1 U892 ( .A1(n1245), .A2(n1061), .A3(n1246), .A4(n1247), .ZN(n1222) );
INV_X1 U893 ( .A(G140), .ZN(n1120) );
XOR2_X1 U894 ( .A(G137), .B(n1248), .Z(G39) );
NOR2_X1 U895 ( .A1(n1059), .A2(n1229), .ZN(n1248) );
NAND4_X1 U896 ( .A1(n1075), .A2(n1249), .A3(n1225), .A4(n1243), .ZN(n1229) );
XNOR2_X1 U897 ( .A(G134), .B(n1230), .ZN(G36) );
NAND3_X1 U898 ( .A1(n1245), .A2(n1060), .A3(n1074), .ZN(n1230) );
XNOR2_X1 U899 ( .A(n1231), .B(n1250), .ZN(G33) );
NOR2_X1 U900 ( .A1(KEYINPUT60), .A2(n1251), .ZN(n1250) );
NAND3_X1 U901 ( .A1(n1245), .A2(n1061), .A3(n1074), .ZN(n1231) );
AND3_X1 U902 ( .A1(n1225), .A2(n1243), .A3(n1082), .ZN(n1245) );
INV_X1 U903 ( .A(n1059), .ZN(n1082) );
NAND2_X1 U904 ( .A1(n1252), .A2(n1067), .ZN(n1059) );
XOR2_X1 U905 ( .A(n1232), .B(n1253), .Z(G30) );
NAND2_X1 U906 ( .A1(n1254), .A2(KEYINPUT25), .ZN(n1253) );
XNOR2_X1 U907 ( .A(G128), .B(KEYINPUT6), .ZN(n1254) );
NAND4_X1 U908 ( .A1(n1075), .A2(n1255), .A3(n1060), .A4(n1256), .ZN(n1232) );
INV_X1 U909 ( .A(n1257), .ZN(n1255) );
NAND3_X1 U910 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(G3) );
OR2_X1 U911 ( .A1(n1234), .A2(G101), .ZN(n1260) );
NAND2_X1 U912 ( .A1(n1261), .A2(n1262), .ZN(n1259) );
INV_X1 U913 ( .A(KEYINPUT4), .ZN(n1262) );
NAND2_X1 U914 ( .A1(G101), .A2(n1263), .ZN(n1261) );
XNOR2_X1 U915 ( .A(KEYINPUT2), .B(n1234), .ZN(n1263) );
NAND2_X1 U916 ( .A1(KEYINPUT4), .A2(n1264), .ZN(n1258) );
NAND2_X1 U917 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
OR2_X1 U918 ( .A1(n1234), .A2(KEYINPUT2), .ZN(n1266) );
NAND3_X1 U919 ( .A1(G101), .A2(n1234), .A3(KEYINPUT2), .ZN(n1265) );
NAND3_X1 U920 ( .A1(n1074), .A2(n1236), .A3(n1267), .ZN(n1234) );
XOR2_X1 U921 ( .A(n1268), .B(G125), .Z(G27) );
NAND2_X1 U922 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
NAND4_X1 U923 ( .A1(n1247), .A2(n1271), .A3(n1272), .A4(n1273), .ZN(n1270) );
NOR2_X1 U924 ( .A1(n1053), .A2(n1257), .ZN(n1272) );
OR2_X1 U925 ( .A1(n1233), .A2(n1273), .ZN(n1269) );
INV_X1 U926 ( .A(KEYINPUT15), .ZN(n1273) );
NAND3_X1 U927 ( .A1(n1084), .A2(n1247), .A3(n1223), .ZN(n1233) );
NOR2_X1 U928 ( .A1(n1271), .A2(n1257), .ZN(n1223) );
NAND3_X1 U929 ( .A1(n1065), .A2(n1243), .A3(n1246), .ZN(n1257) );
NAND2_X1 U930 ( .A1(n1050), .A2(n1274), .ZN(n1243) );
NAND3_X1 U931 ( .A1(G902), .A2(n1275), .A3(n1111), .ZN(n1274) );
NOR2_X1 U932 ( .A1(G900), .A2(n1237), .ZN(n1111) );
XNOR2_X1 U933 ( .A(G122), .B(n1215), .ZN(G24) );
NAND4_X1 U934 ( .A1(n1276), .A2(n1080), .A3(n1242), .A4(n1244), .ZN(n1215) );
INV_X1 U935 ( .A(n1055), .ZN(n1080) );
NAND2_X1 U936 ( .A1(n1247), .A2(n1076), .ZN(n1055) );
XNOR2_X1 U937 ( .A(G119), .B(n1216), .ZN(G21) );
NAND3_X1 U938 ( .A1(n1075), .A2(n1249), .A3(n1276), .ZN(n1216) );
XOR2_X1 U939 ( .A(n1277), .B(n1278), .Z(G18) );
XOR2_X1 U940 ( .A(KEYINPUT8), .B(G116), .Z(n1278) );
NAND2_X1 U941 ( .A1(n1279), .A2(n1065), .ZN(n1277) );
XNOR2_X1 U942 ( .A(n1218), .B(KEYINPUT46), .ZN(n1279) );
AND4_X1 U943 ( .A1(n1074), .A2(n1084), .A3(n1060), .A4(n1280), .ZN(n1218) );
NOR2_X1 U944 ( .A1(n1242), .A2(n1281), .ZN(n1060) );
XNOR2_X1 U945 ( .A(G113), .B(n1217), .ZN(G15) );
NAND3_X1 U946 ( .A1(n1074), .A2(n1061), .A3(n1276), .ZN(n1217) );
AND3_X1 U947 ( .A1(n1065), .A2(n1280), .A3(n1084), .ZN(n1276) );
INV_X1 U948 ( .A(n1053), .ZN(n1084) );
NAND2_X1 U949 ( .A1(n1282), .A2(n1078), .ZN(n1053) );
INV_X1 U950 ( .A(n1271), .ZN(n1061) );
NAND2_X1 U951 ( .A1(n1281), .A2(n1242), .ZN(n1271) );
INV_X1 U952 ( .A(n1244), .ZN(n1281) );
NOR2_X1 U953 ( .A1(n1247), .A2(n1246), .ZN(n1074) );
XNOR2_X1 U954 ( .A(G110), .B(n1235), .ZN(G12) );
NAND3_X1 U955 ( .A1(n1236), .A2(n1247), .A3(n1249), .ZN(n1235) );
NOR2_X1 U956 ( .A1(n1063), .A2(n1076), .ZN(n1249) );
INV_X1 U957 ( .A(n1246), .ZN(n1076) );
XOR2_X1 U958 ( .A(n1283), .B(n1142), .Z(n1246) );
INV_X1 U959 ( .A(n1095), .ZN(n1142) );
NAND2_X1 U960 ( .A1(n1145), .A2(n1284), .ZN(n1095) );
INV_X1 U961 ( .A(n1148), .ZN(n1145) );
XOR2_X1 U962 ( .A(n1285), .B(n1286), .Z(n1148) );
XOR2_X1 U963 ( .A(n1287), .B(n1288), .Z(n1286) );
NAND2_X1 U964 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
NAND2_X1 U965 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XOR2_X1 U966 ( .A(n1293), .B(KEYINPUT33), .Z(n1289) );
OR2_X1 U967 ( .A1(n1292), .A2(n1291), .ZN(n1293) );
XNOR2_X1 U968 ( .A(G110), .B(KEYINPUT10), .ZN(n1291) );
XNOR2_X1 U969 ( .A(n1294), .B(n1295), .ZN(n1292) );
XNOR2_X1 U970 ( .A(G119), .B(KEYINPUT3), .ZN(n1294) );
NAND2_X1 U971 ( .A1(n1296), .A2(KEYINPUT42), .ZN(n1287) );
XNOR2_X1 U972 ( .A(G146), .B(n1297), .ZN(n1296) );
XOR2_X1 U973 ( .A(n1298), .B(n1299), .Z(n1285) );
NAND3_X1 U974 ( .A1(G234), .A2(n1237), .A3(G221), .ZN(n1298) );
NAND2_X1 U975 ( .A1(KEYINPUT38), .A2(n1093), .ZN(n1283) );
NAND2_X1 U976 ( .A1(G217), .A2(n1300), .ZN(n1093) );
INV_X1 U977 ( .A(n1267), .ZN(n1063) );
NOR2_X1 U978 ( .A1(n1244), .A2(n1242), .ZN(n1267) );
XOR2_X1 U979 ( .A(n1090), .B(G475), .Z(n1242) );
NOR2_X1 U980 ( .A1(n1160), .A2(G902), .ZN(n1090) );
XOR2_X1 U981 ( .A(n1301), .B(n1302), .Z(n1160) );
XOR2_X1 U982 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U983 ( .A(G122), .B(G113), .Z(n1304) );
XOR2_X1 U984 ( .A(G143), .B(G131), .Z(n1303) );
XOR2_X1 U985 ( .A(n1305), .B(n1306), .Z(n1301) );
XOR2_X1 U986 ( .A(n1166), .B(n1307), .Z(n1306) );
NAND2_X1 U987 ( .A1(KEYINPUT52), .A2(G146), .ZN(n1307) );
XOR2_X1 U988 ( .A(n1308), .B(n1297), .Z(n1305) );
XOR2_X1 U989 ( .A(G140), .B(G125), .Z(n1297) );
NAND2_X1 U990 ( .A1(n1309), .A2(G214), .ZN(n1308) );
NAND2_X1 U991 ( .A1(n1092), .A2(n1089), .ZN(n1244) );
NAND3_X1 U992 ( .A1(n1156), .A2(n1284), .A3(n1155), .ZN(n1089) );
INV_X1 U993 ( .A(G478), .ZN(n1156) );
NAND2_X1 U994 ( .A1(G478), .A2(n1310), .ZN(n1092) );
NAND2_X1 U995 ( .A1(n1155), .A2(n1284), .ZN(n1310) );
XOR2_X1 U996 ( .A(n1311), .B(n1312), .Z(n1155) );
XOR2_X1 U997 ( .A(G116), .B(n1313), .Z(n1312) );
XOR2_X1 U998 ( .A(G134), .B(G122), .Z(n1313) );
XOR2_X1 U999 ( .A(n1314), .B(n1315), .Z(n1311) );
XOR2_X1 U1000 ( .A(n1316), .B(G107), .Z(n1314) );
NAND3_X1 U1001 ( .A1(G234), .A2(n1317), .A3(G217), .ZN(n1316) );
XOR2_X1 U1002 ( .A(KEYINPUT49), .B(G953), .Z(n1317) );
INV_X1 U1003 ( .A(n1075), .ZN(n1247) );
XOR2_X1 U1004 ( .A(n1318), .B(n1319), .Z(n1075) );
XOR2_X1 U1005 ( .A(KEYINPUT20), .B(G472), .Z(n1319) );
NAND2_X1 U1006 ( .A1(n1320), .A2(n1284), .ZN(n1318) );
XOR2_X1 U1007 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1008 ( .A(n1323), .B(n1186), .Z(n1322) );
NAND2_X1 U1009 ( .A1(n1309), .A2(G210), .ZN(n1186) );
NOR2_X1 U1010 ( .A1(G953), .A2(G237), .ZN(n1309) );
NAND2_X1 U1011 ( .A1(n1324), .A2(n1187), .ZN(n1323) );
XOR2_X1 U1012 ( .A(KEYINPUT41), .B(KEYINPUT19), .Z(n1324) );
XOR2_X1 U1013 ( .A(n1325), .B(n1185), .Z(n1321) );
XOR2_X1 U1014 ( .A(n1209), .B(n1199), .Z(n1185) );
NAND2_X1 U1015 ( .A1(KEYINPUT31), .A2(n1181), .ZN(n1325) );
XOR2_X1 U1016 ( .A(n1326), .B(KEYINPUT39), .Z(n1181) );
NAND3_X1 U1017 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1326) );
NAND2_X1 U1018 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
NAND2_X1 U1019 ( .A1(n1332), .A2(n1333), .ZN(n1328) );
INV_X1 U1020 ( .A(KEYINPUT16), .ZN(n1333) );
NAND2_X1 U1021 ( .A1(n1334), .A2(n1335), .ZN(n1332) );
INV_X1 U1022 ( .A(n1330), .ZN(n1335) );
XOR2_X1 U1023 ( .A(KEYINPUT43), .B(n1331), .Z(n1334) );
NAND2_X1 U1024 ( .A1(KEYINPUT16), .A2(n1336), .ZN(n1327) );
NAND2_X1 U1025 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
NAND2_X1 U1026 ( .A1(n1331), .A2(n1339), .ZN(n1338) );
OR3_X1 U1027 ( .A1(n1330), .A2(n1331), .A3(n1339), .ZN(n1337) );
INV_X1 U1028 ( .A(KEYINPUT43), .ZN(n1339) );
XNOR2_X1 U1029 ( .A(G113), .B(KEYINPUT21), .ZN(n1330) );
AND3_X1 U1030 ( .A1(n1256), .A2(n1280), .A3(n1065), .ZN(n1236) );
AND2_X1 U1031 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U1032 ( .A1(G214), .A2(n1340), .ZN(n1067) );
INV_X1 U1033 ( .A(n1252), .ZN(n1066) );
XNOR2_X1 U1034 ( .A(n1341), .B(n1212), .ZN(n1252) );
NAND2_X1 U1035 ( .A1(G210), .A2(n1340), .ZN(n1212) );
NAND2_X1 U1036 ( .A1(n1342), .A2(n1284), .ZN(n1340) );
INV_X1 U1037 ( .A(G237), .ZN(n1342) );
NAND2_X1 U1038 ( .A1(n1343), .A2(n1284), .ZN(n1341) );
XOR2_X1 U1039 ( .A(n1210), .B(n1344), .Z(n1343) );
XOR2_X1 U1040 ( .A(n1345), .B(KEYINPUT1), .Z(n1344) );
NAND3_X1 U1041 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1345) );
NAND2_X1 U1042 ( .A1(KEYINPUT32), .A2(n1209), .ZN(n1348) );
OR3_X1 U1043 ( .A1(n1349), .A2(KEYINPUT32), .A3(G125), .ZN(n1347) );
NAND2_X1 U1044 ( .A1(G125), .A2(n1349), .ZN(n1346) );
NAND2_X1 U1045 ( .A1(KEYINPUT61), .A2(n1350), .ZN(n1349) );
INV_X1 U1046 ( .A(n1209), .ZN(n1350) );
XOR2_X1 U1047 ( .A(n1351), .B(n1295), .Z(n1209) );
NAND2_X1 U1048 ( .A1(KEYINPUT55), .A2(n1352), .ZN(n1351) );
XOR2_X1 U1049 ( .A(G146), .B(G143), .Z(n1352) );
XOR2_X1 U1050 ( .A(n1353), .B(n1354), .Z(n1210) );
XNOR2_X1 U1051 ( .A(n1135), .B(n1355), .ZN(n1354) );
XOR2_X1 U1052 ( .A(KEYINPUT37), .B(n1356), .Z(n1355) );
AND2_X1 U1053 ( .A1(n1237), .A2(G224), .ZN(n1356) );
XNOR2_X1 U1054 ( .A(G110), .B(G122), .ZN(n1135) );
XNOR2_X1 U1055 ( .A(n1138), .B(n1137), .ZN(n1353) );
XNOR2_X1 U1056 ( .A(n1357), .B(n1331), .ZN(n1137) );
XOR2_X1 U1057 ( .A(G116), .B(G119), .Z(n1331) );
XNOR2_X1 U1058 ( .A(G113), .B(KEYINPUT5), .ZN(n1357) );
AND2_X1 U1059 ( .A1(n1358), .A2(n1359), .ZN(n1138) );
NAND2_X1 U1060 ( .A1(n1360), .A2(n1187), .ZN(n1359) );
XOR2_X1 U1061 ( .A(G104), .B(n1361), .Z(n1360) );
NAND2_X1 U1062 ( .A1(n1362), .A2(G101), .ZN(n1358) );
XOR2_X1 U1063 ( .A(n1166), .B(n1361), .Z(n1362) );
NOR2_X1 U1064 ( .A1(G107), .A2(KEYINPUT22), .ZN(n1361) );
INV_X1 U1065 ( .A(G104), .ZN(n1166) );
NAND2_X1 U1066 ( .A1(n1050), .A2(n1363), .ZN(n1280) );
NAND4_X1 U1067 ( .A1(G953), .A2(G902), .A3(n1275), .A4(n1131), .ZN(n1363) );
INV_X1 U1068 ( .A(G898), .ZN(n1131) );
NAND3_X1 U1069 ( .A1(n1275), .A2(n1237), .A3(n1364), .ZN(n1050) );
XOR2_X1 U1070 ( .A(KEYINPUT14), .B(G952), .Z(n1364) );
NAND2_X1 U1071 ( .A1(G237), .A2(G234), .ZN(n1275) );
XOR2_X1 U1072 ( .A(n1225), .B(KEYINPUT57), .Z(n1256) );
INV_X1 U1073 ( .A(n1081), .ZN(n1225) );
NAND2_X1 U1074 ( .A1(n1079), .A2(n1078), .ZN(n1081) );
NAND2_X1 U1075 ( .A1(G221), .A2(n1300), .ZN(n1078) );
NAND2_X1 U1076 ( .A1(G234), .A2(n1284), .ZN(n1300) );
INV_X1 U1077 ( .A(n1282), .ZN(n1079) );
XOR2_X1 U1078 ( .A(n1365), .B(G469), .Z(n1282) );
NAND4_X1 U1079 ( .A1(n1366), .A2(n1284), .A3(n1367), .A4(n1368), .ZN(n1365) );
NAND3_X1 U1080 ( .A1(n1202), .A2(n1369), .A3(n1204), .ZN(n1368) );
NAND2_X1 U1081 ( .A1(n1370), .A2(n1116), .ZN(n1367) );
XOR2_X1 U1082 ( .A(n1369), .B(n1202), .Z(n1370) );
INV_X1 U1083 ( .A(G902), .ZN(n1284) );
OR2_X1 U1084 ( .A1(n1198), .A2(n1369), .ZN(n1366) );
XNOR2_X1 U1085 ( .A(n1192), .B(n1371), .ZN(n1369) );
XNOR2_X1 U1086 ( .A(KEYINPUT54), .B(n1199), .ZN(n1371) );
XOR2_X1 U1087 ( .A(n1112), .B(KEYINPUT63), .Z(n1199) );
XOR2_X1 U1088 ( .A(n1372), .B(n1299), .Z(n1112) );
XOR2_X1 U1089 ( .A(G137), .B(KEYINPUT29), .Z(n1299) );
XOR2_X1 U1090 ( .A(n1251), .B(G134), .Z(n1372) );
INV_X1 U1091 ( .A(G131), .ZN(n1251) );
XNOR2_X1 U1092 ( .A(n1373), .B(n1374), .ZN(n1192) );
XOR2_X1 U1093 ( .A(G140), .B(G110), .Z(n1374) );
NAND2_X1 U1094 ( .A1(G227), .A2(n1237), .ZN(n1373) );
INV_X1 U1095 ( .A(G953), .ZN(n1237) );
NAND2_X1 U1096 ( .A1(n1204), .A2(n1375), .ZN(n1198) );
INV_X1 U1097 ( .A(n1202), .ZN(n1375) );
XOR2_X1 U1098 ( .A(n1187), .B(n1376), .Z(n1202) );
XOR2_X1 U1099 ( .A(G107), .B(G104), .Z(n1376) );
INV_X1 U1100 ( .A(G101), .ZN(n1187) );
INV_X1 U1101 ( .A(n1116), .ZN(n1204) );
XOR2_X1 U1102 ( .A(n1377), .B(n1315), .Z(n1116) );
XOR2_X1 U1103 ( .A(G143), .B(n1295), .Z(n1315) );
XOR2_X1 U1104 ( .A(G128), .B(KEYINPUT56), .Z(n1295) );
XNOR2_X1 U1105 ( .A(G146), .B(KEYINPUT24), .ZN(n1377) );
endmodule


