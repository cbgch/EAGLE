//Key = 1110011100010110011111010100000010000111110101010000001001110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342;

XOR2_X1 U732 ( .A(n1017), .B(n1018), .Z(G9) );
NOR2_X1 U733 ( .A1(n1019), .A2(n1020), .ZN(G75) );
NOR4_X1 U734 ( .A1(G953), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1020) );
NOR2_X1 U735 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U736 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR3_X1 U737 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
NOR2_X1 U738 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U739 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR3_X1 U740 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1031) );
NOR2_X1 U741 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
XNOR2_X1 U742 ( .A(n1040), .B(KEYINPUT61), .ZN(n1039) );
NOR4_X1 U743 ( .A1(n1041), .A2(n1042), .A3(n1034), .A4(n1035), .ZN(n1026) );
NOR3_X1 U744 ( .A1(n1037), .A2(n1043), .A3(n1044), .ZN(n1042) );
NOR2_X1 U745 ( .A1(n1045), .A2(n1030), .ZN(n1044) );
NOR2_X1 U746 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U747 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U748 ( .A1(n1050), .A2(n1028), .ZN(n1043) );
NOR2_X1 U749 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U750 ( .A1(n1053), .A2(n1054), .ZN(n1041) );
NOR2_X1 U751 ( .A1(n1030), .A2(n1028), .ZN(n1053) );
NOR3_X1 U752 ( .A1(n1021), .A2(G953), .A3(G952), .ZN(n1019) );
AND4_X1 U753 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1021) );
NOR4_X1 U754 ( .A1(n1028), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1058) );
XNOR2_X1 U755 ( .A(G472), .B(n1062), .ZN(n1061) );
XOR2_X1 U756 ( .A(KEYINPUT48), .B(n1063), .Z(n1060) );
XOR2_X1 U757 ( .A(KEYINPUT35), .B(n1064), .Z(n1059) );
AND2_X1 U758 ( .A1(n1065), .A2(G469), .ZN(n1064) );
NOR3_X1 U759 ( .A1(n1066), .A2(n1037), .A3(n1067), .ZN(n1057) );
NOR2_X1 U760 ( .A1(G469), .A2(n1065), .ZN(n1066) );
XOR2_X1 U761 ( .A(KEYINPUT18), .B(n1068), .Z(n1055) );
XOR2_X1 U762 ( .A(n1069), .B(n1070), .Z(G72) );
XOR2_X1 U763 ( .A(n1071), .B(n1072), .Z(n1070) );
NOR2_X1 U764 ( .A1(n1073), .A2(G953), .ZN(n1072) );
NOR2_X1 U765 ( .A1(n1074), .A2(n1075), .ZN(n1071) );
XOR2_X1 U766 ( .A(n1076), .B(n1077), .Z(n1075) );
XOR2_X1 U767 ( .A(G134), .B(n1078), .Z(n1077) );
XOR2_X1 U768 ( .A(G140), .B(G137), .Z(n1078) );
XOR2_X1 U769 ( .A(n1079), .B(n1080), .Z(n1076) );
XOR2_X1 U770 ( .A(n1081), .B(n1082), .Z(n1079) );
NOR2_X1 U771 ( .A1(G125), .A2(KEYINPUT51), .ZN(n1082) );
NOR2_X1 U772 ( .A1(G900), .A2(n1083), .ZN(n1074) );
NOR2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1069) );
AND2_X1 U774 ( .A1(G227), .A2(G900), .ZN(n1084) );
XOR2_X1 U775 ( .A(n1086), .B(n1087), .Z(G69) );
XOR2_X1 U776 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U778 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND2_X1 U779 ( .A1(KEYINPUT43), .A2(n1094), .ZN(n1092) );
NOR2_X1 U780 ( .A1(G898), .A2(n1083), .ZN(n1090) );
INV_X1 U781 ( .A(n1095), .ZN(n1083) );
NAND2_X1 U782 ( .A1(n1085), .A2(n1096), .ZN(n1088) );
NAND3_X1 U783 ( .A1(n1097), .A2(n1018), .A3(n1098), .ZN(n1096) );
XOR2_X1 U784 ( .A(n1099), .B(KEYINPUT34), .Z(n1098) );
NAND2_X1 U785 ( .A1(G953), .A2(n1100), .ZN(n1086) );
NAND2_X1 U786 ( .A1(G224), .A2(G898), .ZN(n1100) );
NOR2_X1 U787 ( .A1(n1101), .A2(n1102), .ZN(G66) );
XOR2_X1 U788 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR2_X1 U789 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NOR2_X1 U790 ( .A1(n1101), .A2(n1107), .ZN(G63) );
XNOR2_X1 U791 ( .A(n1108), .B(n1109), .ZN(n1107) );
AND2_X1 U792 ( .A1(G478), .A2(n1110), .ZN(n1109) );
NOR2_X1 U793 ( .A1(n1101), .A2(n1111), .ZN(G60) );
XOR2_X1 U794 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U795 ( .A1(KEYINPUT46), .A2(n1114), .ZN(n1113) );
XOR2_X1 U796 ( .A(n1115), .B(KEYINPUT8), .Z(n1114) );
NAND2_X1 U797 ( .A1(n1110), .A2(G475), .ZN(n1112) );
XOR2_X1 U798 ( .A(n1116), .B(n1117), .Z(G6) );
NOR2_X1 U799 ( .A1(n1101), .A2(n1118), .ZN(G57) );
XOR2_X1 U800 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U801 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U802 ( .A(n1123), .B(n1124), .Z(n1119) );
AND2_X1 U803 ( .A1(G472), .A2(n1110), .ZN(n1124) );
NOR2_X1 U804 ( .A1(n1101), .A2(n1125), .ZN(G54) );
XOR2_X1 U805 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U806 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND2_X1 U807 ( .A1(KEYINPUT58), .A2(n1130), .ZN(n1128) );
XOR2_X1 U808 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U809 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U810 ( .A1(KEYINPUT31), .A2(n1135), .ZN(n1134) );
NAND2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(n1126) );
NAND2_X1 U812 ( .A1(KEYINPUT38), .A2(n1138), .ZN(n1137) );
NAND2_X1 U813 ( .A1(KEYINPUT22), .A2(n1139), .ZN(n1136) );
INV_X1 U814 ( .A(n1138), .ZN(n1139) );
NAND2_X1 U815 ( .A1(n1110), .A2(G469), .ZN(n1138) );
INV_X1 U816 ( .A(n1106), .ZN(n1110) );
NOR2_X1 U817 ( .A1(n1085), .A2(G952), .ZN(n1101) );
NOR2_X1 U818 ( .A1(n1140), .A2(n1141), .ZN(G51) );
XOR2_X1 U819 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U820 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U821 ( .A(n1146), .B(KEYINPUT45), .Z(n1145) );
NAND2_X1 U822 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NOR2_X1 U823 ( .A1(n1147), .A2(n1148), .ZN(n1144) );
NAND3_X1 U824 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1148) );
NAND2_X1 U825 ( .A1(n1152), .A2(G125), .ZN(n1150) );
XOR2_X1 U826 ( .A(n1153), .B(n1080), .Z(n1152) );
NAND3_X1 U827 ( .A1(n1154), .A2(n1135), .A3(n1155), .ZN(n1149) );
NOR2_X1 U828 ( .A1(n1156), .A2(n1106), .ZN(n1142) );
NAND2_X1 U829 ( .A1(G902), .A2(n1023), .ZN(n1106) );
NAND4_X1 U830 ( .A1(n1073), .A2(n1097), .A3(n1157), .A4(n1099), .ZN(n1023) );
XNOR2_X1 U831 ( .A(KEYINPUT11), .B(n1018), .ZN(n1157) );
NAND3_X1 U832 ( .A1(n1158), .A2(n1052), .A3(n1159), .ZN(n1018) );
AND4_X1 U833 ( .A1(n1160), .A2(n1117), .A3(n1161), .A4(n1162), .ZN(n1097) );
NOR4_X1 U834 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1162) );
AND3_X1 U835 ( .A1(n1040), .A2(n1167), .A3(n1158), .ZN(n1166) );
NOR4_X1 U836 ( .A1(n1168), .A2(n1169), .A3(n1047), .A4(n1034), .ZN(n1164) );
NAND2_X1 U837 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
INV_X1 U838 ( .A(KEYINPUT15), .ZN(n1168) );
NOR2_X1 U839 ( .A1(KEYINPUT15), .A2(n1172), .ZN(n1163) );
NAND3_X1 U840 ( .A1(n1159), .A2(n1158), .A3(n1051), .ZN(n1117) );
AND2_X1 U841 ( .A1(n1173), .A2(n1174), .ZN(n1073) );
AND4_X1 U842 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1174) );
NOR4_X1 U843 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1173) );
NOR2_X1 U844 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XNOR2_X1 U845 ( .A(n1185), .B(KEYINPUT16), .ZN(n1183) );
INV_X1 U846 ( .A(n1186), .ZN(n1181) );
INV_X1 U847 ( .A(n1187), .ZN(n1180) );
NOR3_X1 U848 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1179) );
NOR2_X1 U849 ( .A1(KEYINPUT14), .A2(n1191), .ZN(n1190) );
NOR3_X1 U850 ( .A1(n1028), .A2(n1192), .A3(n1193), .ZN(n1191) );
AND2_X1 U851 ( .A1(n1194), .A2(KEYINPUT14), .ZN(n1189) );
NOR2_X1 U852 ( .A1(n1085), .A2(n1195), .ZN(n1140) );
XOR2_X1 U853 ( .A(KEYINPUT27), .B(G952), .Z(n1195) );
XNOR2_X1 U854 ( .A(G146), .B(n1178), .ZN(G48) );
NAND3_X1 U855 ( .A1(n1185), .A2(n1196), .A3(n1051), .ZN(n1178) );
XOR2_X1 U856 ( .A(n1197), .B(n1198), .Z(G45) );
NOR2_X1 U857 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NOR3_X1 U858 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
AND4_X1 U859 ( .A1(n1204), .A2(n1192), .A3(n1038), .A4(n1171), .ZN(n1202) );
INV_X1 U860 ( .A(KEYINPUT53), .ZN(n1201) );
NOR2_X1 U861 ( .A1(KEYINPUT53), .A2(n1177), .ZN(n1199) );
NAND3_X1 U862 ( .A1(n1038), .A2(n1196), .A3(n1171), .ZN(n1177) );
XOR2_X1 U863 ( .A(n1205), .B(n1186), .Z(G42) );
NAND3_X1 U864 ( .A1(n1051), .A2(n1206), .A3(n1040), .ZN(n1186) );
XOR2_X1 U865 ( .A(n1207), .B(n1208), .Z(G39) );
XOR2_X1 U866 ( .A(KEYINPUT39), .B(G137), .Z(n1208) );
NAND3_X1 U867 ( .A1(n1209), .A2(n1185), .A3(KEYINPUT62), .ZN(n1207) );
INV_X1 U868 ( .A(n1184), .ZN(n1209) );
NAND2_X1 U869 ( .A1(n1206), .A2(n1167), .ZN(n1184) );
XOR2_X1 U870 ( .A(G134), .B(n1210), .Z(G36) );
NOR2_X1 U871 ( .A1(n1194), .A2(n1188), .ZN(n1210) );
INV_X1 U872 ( .A(n1206), .ZN(n1194) );
XNOR2_X1 U873 ( .A(G131), .B(n1176), .ZN(G33) );
NAND3_X1 U874 ( .A1(n1038), .A2(n1206), .A3(n1051), .ZN(n1176) );
NOR3_X1 U875 ( .A1(n1033), .A2(n1193), .A3(n1028), .ZN(n1206) );
NAND2_X1 U876 ( .A1(n1211), .A2(n1049), .ZN(n1028) );
XNOR2_X1 U877 ( .A(n1175), .B(n1212), .ZN(G30) );
NOR2_X1 U878 ( .A1(KEYINPUT33), .A2(n1213), .ZN(n1212) );
NAND3_X1 U879 ( .A1(n1196), .A2(n1052), .A3(n1185), .ZN(n1175) );
NOR3_X1 U880 ( .A1(n1203), .A2(n1193), .A3(n1033), .ZN(n1196) );
XOR2_X1 U881 ( .A(G101), .B(n1165), .Z(G3) );
AND3_X1 U882 ( .A1(n1158), .A2(n1167), .A3(n1038), .ZN(n1165) );
XOR2_X1 U883 ( .A(n1155), .B(n1187), .Z(G27) );
NAND4_X1 U884 ( .A1(n1214), .A2(n1051), .A3(n1040), .A4(n1215), .ZN(n1187) );
NOR3_X1 U885 ( .A1(n1203), .A2(n1037), .A3(n1193), .ZN(n1215) );
INV_X1 U886 ( .A(n1204), .ZN(n1193) );
NAND2_X1 U887 ( .A1(n1025), .A2(n1216), .ZN(n1204) );
NAND4_X1 U888 ( .A1(n1095), .A2(G902), .A3(n1217), .A4(n1218), .ZN(n1216) );
INV_X1 U889 ( .A(G900), .ZN(n1218) );
INV_X1 U890 ( .A(n1054), .ZN(n1037) );
XNOR2_X1 U891 ( .A(n1172), .B(n1219), .ZN(G24) );
NOR2_X1 U892 ( .A1(KEYINPUT26), .A2(n1220), .ZN(n1219) );
INV_X1 U893 ( .A(G122), .ZN(n1220) );
NAND4_X1 U894 ( .A1(n1170), .A2(n1171), .A3(n1159), .A4(n1047), .ZN(n1172) );
INV_X1 U895 ( .A(n1034), .ZN(n1159) );
NAND2_X1 U896 ( .A1(n1221), .A2(n1222), .ZN(n1034) );
NOR2_X1 U897 ( .A1(n1056), .A2(n1223), .ZN(n1171) );
XNOR2_X1 U898 ( .A(G119), .B(n1099), .ZN(G21) );
NAND4_X1 U899 ( .A1(n1170), .A2(n1185), .A3(n1167), .A4(n1047), .ZN(n1099) );
NOR2_X1 U900 ( .A1(n1222), .A2(n1221), .ZN(n1185) );
XNOR2_X1 U901 ( .A(G116), .B(n1161), .ZN(G18) );
NAND3_X1 U902 ( .A1(n1224), .A2(n1047), .A3(n1170), .ZN(n1161) );
INV_X1 U903 ( .A(n1188), .ZN(n1224) );
NAND2_X1 U904 ( .A1(n1038), .A2(n1052), .ZN(n1188) );
NAND2_X1 U905 ( .A1(n1225), .A2(n1226), .ZN(n1052) );
OR2_X1 U906 ( .A1(n1030), .A2(KEYINPUT1), .ZN(n1226) );
NAND3_X1 U907 ( .A1(n1223), .A2(n1227), .A3(KEYINPUT1), .ZN(n1225) );
XNOR2_X1 U908 ( .A(G113), .B(n1160), .ZN(G15) );
NAND4_X1 U909 ( .A1(n1170), .A2(n1051), .A3(n1038), .A4(n1228), .ZN(n1160) );
NOR2_X1 U910 ( .A1(n1063), .A2(n1221), .ZN(n1038) );
INV_X1 U911 ( .A(n1229), .ZN(n1221) );
INV_X1 U912 ( .A(n1222), .ZN(n1063) );
NOR2_X1 U913 ( .A1(n1227), .A2(n1223), .ZN(n1051) );
AND3_X1 U914 ( .A1(n1230), .A2(n1054), .A3(n1214), .ZN(n1170) );
XNOR2_X1 U915 ( .A(G110), .B(n1231), .ZN(G12) );
NAND3_X1 U916 ( .A1(n1158), .A2(n1232), .A3(n1040), .ZN(n1231) );
NOR2_X1 U917 ( .A1(n1229), .A2(n1222), .ZN(n1040) );
XNOR2_X1 U918 ( .A(n1233), .B(n1105), .ZN(n1222) );
NAND2_X1 U919 ( .A1(G217), .A2(n1234), .ZN(n1105) );
OR2_X1 U920 ( .A1(n1104), .A2(n1235), .ZN(n1233) );
XNOR2_X1 U921 ( .A(n1236), .B(n1237), .ZN(n1104) );
XOR2_X1 U922 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U923 ( .A(n1240), .B(KEYINPUT23), .Z(n1239) );
NAND3_X1 U924 ( .A1(n1241), .A2(n1085), .A3(G221), .ZN(n1240) );
XOR2_X1 U925 ( .A(KEYINPUT40), .B(n1242), .Z(n1241) );
NAND2_X1 U926 ( .A1(n1243), .A2(KEYINPUT32), .ZN(n1238) );
XOR2_X1 U927 ( .A(G119), .B(n1213), .Z(n1243) );
XOR2_X1 U928 ( .A(n1244), .B(n1245), .Z(n1236) );
XOR2_X1 U929 ( .A(n1246), .B(n1247), .Z(n1244) );
NAND2_X1 U930 ( .A1(KEYINPUT41), .A2(n1248), .ZN(n1246) );
NAND2_X1 U931 ( .A1(n1249), .A2(n1250), .ZN(n1229) );
NAND2_X1 U932 ( .A1(G472), .A2(n1062), .ZN(n1250) );
XOR2_X1 U933 ( .A(KEYINPUT59), .B(n1251), .Z(n1249) );
NOR2_X1 U934 ( .A1(G472), .A2(n1062), .ZN(n1251) );
NAND2_X1 U935 ( .A1(n1252), .A2(n1253), .ZN(n1062) );
XOR2_X1 U936 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U937 ( .A(n1256), .B(n1080), .Z(n1255) );
XOR2_X1 U938 ( .A(n1257), .B(n1258), .Z(n1254) );
NOR2_X1 U939 ( .A1(KEYINPUT24), .A2(n1131), .ZN(n1258) );
XNOR2_X1 U940 ( .A(KEYINPUT21), .B(n1259), .ZN(n1257) );
NOR2_X1 U941 ( .A1(KEYINPUT9), .A2(n1260), .ZN(n1259) );
XOR2_X1 U942 ( .A(n1123), .B(n1261), .Z(n1260) );
XOR2_X1 U943 ( .A(KEYINPUT47), .B(G101), .Z(n1261) );
NAND3_X1 U944 ( .A1(n1262), .A2(n1085), .A3(G210), .ZN(n1123) );
XOR2_X1 U945 ( .A(KEYINPUT42), .B(n1167), .Z(n1232) );
INV_X1 U946 ( .A(n1030), .ZN(n1167) );
NAND2_X1 U947 ( .A1(n1223), .A2(n1056), .ZN(n1030) );
INV_X1 U948 ( .A(n1227), .ZN(n1056) );
XOR2_X1 U949 ( .A(n1263), .B(n1264), .Z(n1227) );
XOR2_X1 U950 ( .A(KEYINPUT0), .B(G478), .Z(n1264) );
NAND2_X1 U951 ( .A1(n1252), .A2(n1108), .ZN(n1263) );
XNOR2_X1 U952 ( .A(n1265), .B(n1266), .ZN(n1108) );
NOR3_X1 U953 ( .A1(n1242), .A2(G953), .A3(n1267), .ZN(n1266) );
INV_X1 U954 ( .A(G217), .ZN(n1267) );
XOR2_X1 U955 ( .A(G234), .B(KEYINPUT13), .Z(n1242) );
NAND3_X1 U956 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1265) );
NAND2_X1 U957 ( .A1(KEYINPUT52), .A2(n1271), .ZN(n1270) );
NAND3_X1 U958 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n1269) );
INV_X1 U959 ( .A(KEYINPUT52), .ZN(n1273) );
OR2_X1 U960 ( .A1(n1274), .A2(n1272), .ZN(n1268) );
NOR2_X1 U961 ( .A1(KEYINPUT49), .A2(n1271), .ZN(n1272) );
XOR2_X1 U962 ( .A(n1275), .B(G134), .Z(n1271) );
NAND2_X1 U963 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND2_X1 U964 ( .A1(G128), .A2(n1197), .ZN(n1277) );
XOR2_X1 U965 ( .A(n1278), .B(KEYINPUT10), .Z(n1276) );
NAND2_X1 U966 ( .A1(G143), .A2(n1213), .ZN(n1278) );
XNOR2_X1 U967 ( .A(G107), .B(n1279), .ZN(n1274) );
XOR2_X1 U968 ( .A(G122), .B(G116), .Z(n1279) );
NOR2_X1 U969 ( .A1(n1068), .A2(n1067), .ZN(n1223) );
AND2_X1 U970 ( .A1(n1280), .A2(G475), .ZN(n1067) );
NOR2_X1 U971 ( .A1(n1280), .A2(G475), .ZN(n1068) );
OR2_X1 U972 ( .A1(n1115), .A2(n1235), .ZN(n1280) );
NAND3_X1 U973 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1115) );
NAND2_X1 U974 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
INV_X1 U975 ( .A(KEYINPUT57), .ZN(n1285) );
NAND3_X1 U976 ( .A1(KEYINPUT57), .A2(n1286), .A3(n1287), .ZN(n1282) );
OR2_X1 U977 ( .A1(n1287), .A2(n1286), .ZN(n1281) );
NOR2_X1 U978 ( .A1(n1288), .A2(n1284), .ZN(n1286) );
XNOR2_X1 U979 ( .A(n1116), .B(n1289), .ZN(n1284) );
XOR2_X1 U980 ( .A(G122), .B(G113), .Z(n1289) );
INV_X1 U981 ( .A(KEYINPUT19), .ZN(n1288) );
XNOR2_X1 U982 ( .A(n1290), .B(n1291), .ZN(n1287) );
XOR2_X1 U983 ( .A(n1292), .B(n1293), .Z(n1291) );
NAND2_X1 U984 ( .A1(KEYINPUT6), .A2(n1205), .ZN(n1293) );
INV_X1 U985 ( .A(G140), .ZN(n1205) );
NAND2_X1 U986 ( .A1(n1294), .A2(n1295), .ZN(n1292) );
NAND2_X1 U987 ( .A1(n1296), .A2(n1197), .ZN(n1295) );
XOR2_X1 U988 ( .A(n1297), .B(KEYINPUT50), .Z(n1294) );
NAND2_X1 U989 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
INV_X1 U990 ( .A(n1296), .ZN(n1299) );
NAND3_X1 U991 ( .A1(n1262), .A2(n1085), .A3(G214), .ZN(n1296) );
XOR2_X1 U992 ( .A(n1197), .B(KEYINPUT25), .Z(n1298) );
INV_X1 U993 ( .A(G143), .ZN(n1197) );
XOR2_X1 U994 ( .A(n1247), .B(n1081), .Z(n1290) );
XOR2_X1 U995 ( .A(G146), .B(G125), .Z(n1247) );
AND3_X1 U996 ( .A1(n1228), .A2(n1230), .A3(n1192), .ZN(n1158) );
INV_X1 U997 ( .A(n1033), .ZN(n1192) );
NAND2_X1 U998 ( .A1(n1035), .A2(n1054), .ZN(n1033) );
NAND2_X1 U999 ( .A1(G221), .A2(n1234), .ZN(n1054) );
NAND2_X1 U1000 ( .A1(G234), .A2(n1300), .ZN(n1234) );
INV_X1 U1001 ( .A(n1214), .ZN(n1035) );
XNOR2_X1 U1002 ( .A(G469), .B(n1301), .ZN(n1214) );
NOR2_X1 U1003 ( .A1(KEYINPUT56), .A2(n1065), .ZN(n1301) );
NAND2_X1 U1004 ( .A1(n1252), .A2(n1302), .ZN(n1065) );
XOR2_X1 U1005 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U1006 ( .A(n1305), .B(n1122), .Z(n1304) );
XOR2_X1 U1007 ( .A(n1080), .B(n1306), .Z(n1122) );
INV_X1 U1008 ( .A(n1131), .ZN(n1306) );
XOR2_X1 U1009 ( .A(n1307), .B(n1308), .Z(n1131) );
INV_X1 U1010 ( .A(n1081), .ZN(n1308) );
XNOR2_X1 U1011 ( .A(G131), .B(KEYINPUT4), .ZN(n1081) );
NAND4_X1 U1012 ( .A1(KEYINPUT63), .A2(n1309), .A3(n1310), .A4(n1311), .ZN(n1307) );
NAND3_X1 U1013 ( .A1(n1312), .A2(n1313), .A3(n1248), .ZN(n1311) );
INV_X1 U1014 ( .A(KEYINPUT28), .ZN(n1313) );
OR2_X1 U1015 ( .A1(n1248), .A2(n1312), .ZN(n1310) );
NOR2_X1 U1016 ( .A1(n1314), .A2(G134), .ZN(n1312) );
INV_X1 U1017 ( .A(KEYINPUT2), .ZN(n1314) );
INV_X1 U1018 ( .A(G137), .ZN(n1248) );
NAND2_X1 U1019 ( .A1(KEYINPUT28), .A2(G134), .ZN(n1309) );
INV_X1 U1020 ( .A(n1133), .ZN(n1305) );
XOR2_X1 U1021 ( .A(n1315), .B(n1316), .Z(n1133) );
XOR2_X1 U1022 ( .A(KEYINPUT30), .B(G101), .Z(n1316) );
NAND3_X1 U1023 ( .A1(n1317), .A2(n1318), .A3(n1319), .ZN(n1315) );
OR2_X1 U1024 ( .A1(n1116), .A2(KEYINPUT7), .ZN(n1319) );
NAND3_X1 U1025 ( .A1(KEYINPUT7), .A2(n1320), .A3(n1017), .ZN(n1318) );
OR2_X1 U1026 ( .A1(n1017), .A2(n1320), .ZN(n1317) );
NOR2_X1 U1027 ( .A1(G104), .A2(KEYINPUT29), .ZN(n1320) );
XOR2_X1 U1028 ( .A(KEYINPUT3), .B(n1321), .Z(n1303) );
INV_X1 U1029 ( .A(n1129), .ZN(n1321) );
XOR2_X1 U1030 ( .A(n1322), .B(n1245), .Z(n1129) );
XOR2_X1 U1031 ( .A(G110), .B(G140), .Z(n1245) );
NAND2_X1 U1032 ( .A1(G227), .A2(n1085), .ZN(n1322) );
NAND2_X1 U1033 ( .A1(n1323), .A2(n1025), .ZN(n1230) );
NAND3_X1 U1034 ( .A1(n1217), .A2(n1085), .A3(G952), .ZN(n1025) );
NAND4_X1 U1035 ( .A1(n1095), .A2(G902), .A3(n1324), .A4(n1217), .ZN(n1323) );
NAND2_X1 U1036 ( .A1(G237), .A2(G234), .ZN(n1217) );
XOR2_X1 U1037 ( .A(KEYINPUT54), .B(G898), .Z(n1324) );
XOR2_X1 U1038 ( .A(n1085), .B(KEYINPUT20), .Z(n1095) );
XOR2_X1 U1039 ( .A(n1047), .B(KEYINPUT44), .Z(n1228) );
INV_X1 U1040 ( .A(n1203), .ZN(n1047) );
NAND2_X1 U1041 ( .A1(n1325), .A2(n1049), .ZN(n1203) );
NAND2_X1 U1042 ( .A1(G214), .A2(n1326), .ZN(n1049) );
XOR2_X1 U1043 ( .A(KEYINPUT60), .B(n1048), .Z(n1325) );
INV_X1 U1044 ( .A(n1211), .ZN(n1048) );
XOR2_X1 U1045 ( .A(n1156), .B(n1327), .Z(n1211) );
NOR2_X1 U1046 ( .A1(n1328), .A2(n1235), .ZN(n1327) );
INV_X1 U1047 ( .A(n1252), .ZN(n1235) );
XOR2_X1 U1048 ( .A(n1300), .B(KEYINPUT12), .Z(n1252) );
XNOR2_X1 U1049 ( .A(n1147), .B(n1329), .ZN(n1328) );
NOR4_X1 U1050 ( .A1(n1330), .A2(n1331), .A3(KEYINPUT55), .A4(n1332), .ZN(n1329) );
INV_X1 U1051 ( .A(n1151), .ZN(n1332) );
NAND3_X1 U1052 ( .A1(n1153), .A2(n1155), .A3(n1080), .ZN(n1151) );
INV_X1 U1053 ( .A(G125), .ZN(n1155) );
NOR3_X1 U1054 ( .A1(n1153), .A2(n1333), .A3(n1334), .ZN(n1331) );
NOR2_X1 U1055 ( .A1(G125), .A2(n1135), .ZN(n1334) );
INV_X1 U1056 ( .A(n1335), .ZN(n1333) );
NOR2_X1 U1057 ( .A1(n1154), .A2(n1335), .ZN(n1330) );
NAND2_X1 U1058 ( .A1(G125), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1059 ( .A(KEYINPUT5), .B(n1080), .Z(n1336) );
INV_X1 U1060 ( .A(n1135), .ZN(n1080) );
XOR2_X1 U1061 ( .A(n1213), .B(n1337), .Z(n1135) );
XOR2_X1 U1062 ( .A(G146), .B(G143), .Z(n1337) );
INV_X1 U1063 ( .A(G128), .ZN(n1213) );
INV_X1 U1064 ( .A(n1153), .ZN(n1154) );
NAND2_X1 U1065 ( .A1(n1338), .A2(n1085), .ZN(n1153) );
INV_X1 U1066 ( .A(G953), .ZN(n1085) );
XNOR2_X1 U1067 ( .A(G224), .B(KEYINPUT37), .ZN(n1338) );
XOR2_X1 U1068 ( .A(n1094), .B(n1093), .Z(n1147) );
XOR2_X1 U1069 ( .A(G110), .B(n1339), .Z(n1093) );
XOR2_X1 U1070 ( .A(KEYINPUT36), .B(G122), .Z(n1339) );
XOR2_X1 U1071 ( .A(n1121), .B(n1340), .Z(n1094) );
XOR2_X1 U1072 ( .A(n1017), .B(n1341), .Z(n1340) );
NAND2_X1 U1073 ( .A1(KEYINPUT17), .A2(n1116), .ZN(n1341) );
INV_X1 U1074 ( .A(G104), .ZN(n1116) );
INV_X1 U1075 ( .A(G107), .ZN(n1017) );
XNOR2_X1 U1076 ( .A(n1256), .B(G101), .ZN(n1121) );
XNOR2_X1 U1077 ( .A(G113), .B(n1342), .ZN(n1256) );
XOR2_X1 U1078 ( .A(G119), .B(G116), .Z(n1342) );
NAND2_X1 U1079 ( .A1(G210), .A2(n1326), .ZN(n1156) );
NAND2_X1 U1080 ( .A1(n1262), .A2(n1300), .ZN(n1326) );
INV_X1 U1081 ( .A(G902), .ZN(n1300) );
INV_X1 U1082 ( .A(G237), .ZN(n1262) );
endmodule


