//Key = 1101011000000001000100010011000110001011011000010010000011100011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338;

XNOR2_X1 U737 ( .A(G107), .B(n1019), .ZN(G9) );
NOR2_X1 U738 ( .A1(n1020), .A2(n1021), .ZN(G75) );
NOR4_X1 U739 ( .A1(n1022), .A2(n1023), .A3(G953), .A4(n1024), .ZN(n1021) );
INV_X1 U740 ( .A(G952), .ZN(n1023) );
NAND2_X1 U741 ( .A1(n1025), .A2(n1026), .ZN(n1022) );
XOR2_X1 U742 ( .A(n1027), .B(KEYINPUT1), .Z(n1025) );
NAND2_X1 U743 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND3_X1 U744 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NAND2_X1 U745 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NAND2_X1 U746 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(n1028) );
NAND3_X1 U748 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
XOR2_X1 U749 ( .A(n1042), .B(KEYINPUT48), .Z(n1041) );
NAND3_X1 U750 ( .A1(n1032), .A2(n1043), .A3(n1044), .ZN(n1042) );
NAND2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1040) );
NAND2_X1 U752 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U753 ( .A1(n1049), .A2(n1050), .A3(n1030), .ZN(n1048) );
OR2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U755 ( .A1(n1053), .A2(n1054), .ZN(n1047) );
NAND3_X1 U756 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NAND2_X1 U757 ( .A1(n1030), .A2(n1058), .ZN(n1057) );
NAND3_X1 U758 ( .A1(n1059), .A2(n1060), .A3(n1049), .ZN(n1056) );
INV_X1 U759 ( .A(KEYINPUT37), .ZN(n1060) );
NAND2_X1 U760 ( .A1(n1061), .A2(n1062), .ZN(n1055) );
XOR2_X1 U761 ( .A(KEYINPUT49), .B(n1030), .Z(n1062) );
NAND2_X1 U762 ( .A1(KEYINPUT37), .A2(n1063), .ZN(n1039) );
NAND2_X1 U763 ( .A1(n1032), .A2(n1059), .ZN(n1063) );
AND3_X1 U764 ( .A1(n1053), .A2(n1049), .A3(n1045), .ZN(n1032) );
INV_X1 U765 ( .A(n1064), .ZN(n1045) );
NOR3_X1 U766 ( .A1(n1024), .A2(n1065), .A3(n1066), .ZN(n1020) );
NOR2_X1 U767 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
INV_X1 U768 ( .A(KEYINPUT0), .ZN(n1068) );
NOR2_X1 U769 ( .A1(G953), .A2(G952), .ZN(n1067) );
NOR2_X1 U770 ( .A1(KEYINPUT0), .A2(n1069), .ZN(n1065) );
AND4_X1 U771 ( .A1(n1070), .A2(n1037), .A3(n1071), .A4(n1072), .ZN(n1024) );
NOR4_X1 U772 ( .A1(n1044), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1072) );
XNOR2_X1 U773 ( .A(n1076), .B(n1077), .ZN(n1074) );
XNOR2_X1 U774 ( .A(n1078), .B(KEYINPUT15), .ZN(n1076) );
XNOR2_X1 U775 ( .A(n1079), .B(KEYINPUT41), .ZN(n1073) );
XNOR2_X1 U776 ( .A(n1080), .B(n1081), .ZN(n1071) );
XOR2_X1 U777 ( .A(n1082), .B(n1083), .Z(G72) );
XOR2_X1 U778 ( .A(n1084), .B(n1085), .Z(n1083) );
NOR2_X1 U779 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U780 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U781 ( .A1(KEYINPUT24), .A2(n1090), .ZN(n1089) );
XOR2_X1 U782 ( .A(n1091), .B(n1092), .Z(n1090) );
XNOR2_X1 U783 ( .A(n1093), .B(n1094), .ZN(n1092) );
XNOR2_X1 U784 ( .A(KEYINPUT57), .B(n1095), .ZN(n1091) );
NOR2_X1 U785 ( .A1(G134), .A2(KEYINPUT60), .ZN(n1095) );
NOR2_X1 U786 ( .A1(G900), .A2(n1096), .ZN(n1086) );
NAND2_X1 U787 ( .A1(n1097), .A2(n1096), .ZN(n1084) );
NAND2_X1 U788 ( .A1(n1098), .A2(n1099), .ZN(n1082) );
NAND2_X1 U789 ( .A1(G900), .A2(G227), .ZN(n1099) );
INV_X1 U790 ( .A(n1100), .ZN(n1098) );
XOR2_X1 U791 ( .A(n1101), .B(n1102), .Z(G69) );
NOR2_X1 U792 ( .A1(n1103), .A2(n1100), .ZN(n1102) );
XOR2_X1 U793 ( .A(G953), .B(KEYINPUT39), .Z(n1100) );
AND2_X1 U794 ( .A1(G224), .A2(G898), .ZN(n1103) );
NAND2_X1 U795 ( .A1(n1104), .A2(n1105), .ZN(n1101) );
NAND3_X1 U796 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
XOR2_X1 U797 ( .A(n1109), .B(KEYINPUT10), .Z(n1104) );
NAND2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1108), .A2(n1106), .ZN(n1111) );
INV_X1 U800 ( .A(n1112), .ZN(n1106) );
XOR2_X1 U801 ( .A(n1113), .B(n1114), .Z(n1108) );
XNOR2_X1 U802 ( .A(KEYINPUT53), .B(n1107), .ZN(n1110) );
NAND2_X1 U803 ( .A1(n1115), .A2(n1116), .ZN(n1107) );
XNOR2_X1 U804 ( .A(G953), .B(KEYINPUT2), .ZN(n1115) );
NOR2_X1 U805 ( .A1(n1069), .A2(n1117), .ZN(G66) );
NOR3_X1 U806 ( .A1(n1078), .A2(n1118), .A3(n1119), .ZN(n1117) );
AND4_X1 U807 ( .A1(n1120), .A2(KEYINPUT56), .A3(n1121), .A4(n1122), .ZN(n1119) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1120), .ZN(n1118) );
NOR3_X1 U809 ( .A1(n1124), .A2(n1026), .A3(n1077), .ZN(n1123) );
INV_X1 U810 ( .A(KEYINPUT56), .ZN(n1124) );
NOR2_X1 U811 ( .A1(n1069), .A2(n1125), .ZN(G63) );
XOR2_X1 U812 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U813 ( .A1(n1122), .A2(G478), .ZN(n1126) );
NOR2_X1 U814 ( .A1(n1069), .A2(n1128), .ZN(G60) );
XOR2_X1 U815 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U816 ( .A1(n1122), .A2(G475), .ZN(n1129) );
XNOR2_X1 U817 ( .A(G104), .B(n1131), .ZN(G6) );
NOR2_X1 U818 ( .A1(n1069), .A2(n1132), .ZN(G57) );
XOR2_X1 U819 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U820 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U821 ( .A(n1137), .B(n1138), .Z(n1133) );
XOR2_X1 U822 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U823 ( .A1(n1122), .A2(G472), .ZN(n1140) );
NAND2_X1 U824 ( .A1(KEYINPUT19), .A2(n1141), .ZN(n1137) );
NOR3_X1 U825 ( .A1(n1069), .A2(n1142), .A3(n1143), .ZN(G54) );
NOR2_X1 U826 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U827 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U828 ( .A1(KEYINPUT47), .A2(n1148), .ZN(n1146) );
NOR2_X1 U829 ( .A1(n1093), .A2(n1149), .ZN(n1142) );
XOR2_X1 U830 ( .A(n1150), .B(n1147), .Z(n1149) );
NAND2_X1 U831 ( .A1(n1151), .A2(n1152), .ZN(n1147) );
NAND2_X1 U832 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XNOR2_X1 U833 ( .A(n1155), .B(KEYINPUT18), .ZN(n1153) );
NAND2_X1 U834 ( .A1(n1156), .A2(n1157), .ZN(n1151) );
XNOR2_X1 U835 ( .A(KEYINPUT8), .B(n1158), .ZN(n1156) );
INV_X1 U836 ( .A(n1155), .ZN(n1158) );
XNOR2_X1 U837 ( .A(n1159), .B(n1160), .ZN(n1155) );
NAND2_X1 U838 ( .A1(n1122), .A2(G469), .ZN(n1159) );
NAND2_X1 U839 ( .A1(n1161), .A2(KEYINPUT47), .ZN(n1150) );
INV_X1 U840 ( .A(n1148), .ZN(n1161) );
XOR2_X1 U841 ( .A(n1162), .B(n1163), .Z(n1148) );
NOR2_X1 U842 ( .A1(KEYINPUT4), .A2(n1164), .ZN(n1163) );
NOR2_X1 U843 ( .A1(n1069), .A2(n1165), .ZN(G51) );
XOR2_X1 U844 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U845 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U846 ( .A(n1170), .B(KEYINPUT29), .Z(n1169) );
NAND2_X1 U847 ( .A1(KEYINPUT62), .A2(n1171), .ZN(n1170) );
XOR2_X1 U848 ( .A(KEYINPUT40), .B(n1172), .Z(n1171) );
NAND2_X1 U849 ( .A1(n1122), .A2(n1173), .ZN(n1168) );
NOR2_X1 U850 ( .A1(n1174), .A2(n1026), .ZN(n1122) );
NOR2_X1 U851 ( .A1(n1116), .A2(n1097), .ZN(n1026) );
NAND4_X1 U852 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1097) );
NOR4_X1 U853 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1178) );
NOR3_X1 U854 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1177) );
NOR3_X1 U855 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1185) );
AND2_X1 U856 ( .A1(n1186), .A2(n1189), .ZN(n1184) );
INV_X1 U857 ( .A(KEYINPUT52), .ZN(n1186) );
NOR2_X1 U858 ( .A1(n1190), .A2(n1191), .ZN(n1183) );
NAND3_X1 U859 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1175) );
INV_X1 U860 ( .A(n1195), .ZN(n1194) );
XNOR2_X1 U861 ( .A(n1196), .B(KEYINPUT12), .ZN(n1192) );
NAND2_X1 U862 ( .A1(n1197), .A2(n1198), .ZN(n1116) );
AND4_X1 U863 ( .A1(n1019), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1198) );
NAND3_X1 U864 ( .A1(n1052), .A2(n1202), .A3(n1049), .ZN(n1019) );
AND4_X1 U865 ( .A1(n1203), .A2(n1204), .A3(n1131), .A4(n1205), .ZN(n1197) );
NAND3_X1 U866 ( .A1(n1053), .A2(n1202), .A3(n1061), .ZN(n1205) );
NAND3_X1 U867 ( .A1(n1049), .A2(n1202), .A3(n1051), .ZN(n1131) );
XOR2_X1 U868 ( .A(n1206), .B(n1207), .Z(n1166) );
NOR3_X1 U869 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1207) );
NOR3_X1 U870 ( .A1(n1211), .A2(n1144), .A3(n1212), .ZN(n1210) );
INV_X1 U871 ( .A(KEYINPUT27), .ZN(n1211) );
NOR2_X1 U872 ( .A1(KEYINPUT27), .A2(n1093), .ZN(n1209) );
NOR2_X1 U873 ( .A1(n1096), .A2(G952), .ZN(n1069) );
XNOR2_X1 U874 ( .A(G146), .B(n1176), .ZN(G48) );
NAND4_X1 U875 ( .A1(n1051), .A2(n1213), .A3(n1187), .A4(n1193), .ZN(n1176) );
XOR2_X1 U876 ( .A(G143), .B(n1214), .Z(G45) );
NOR3_X1 U877 ( .A1(n1215), .A2(n1196), .A3(n1195), .ZN(n1214) );
NAND3_X1 U878 ( .A1(n1216), .A2(n1079), .A3(n1213), .ZN(n1195) );
XNOR2_X1 U879 ( .A(KEYINPUT17), .B(n1193), .ZN(n1215) );
NAND2_X1 U880 ( .A1(n1217), .A2(n1218), .ZN(G42) );
NAND2_X1 U881 ( .A1(G140), .A2(n1219), .ZN(n1218) );
XOR2_X1 U882 ( .A(KEYINPUT6), .B(n1220), .Z(n1217) );
NOR2_X1 U883 ( .A1(G140), .A2(n1219), .ZN(n1220) );
NAND2_X1 U884 ( .A1(n1221), .A2(n1222), .ZN(n1219) );
XNOR2_X1 U885 ( .A(KEYINPUT34), .B(n1190), .ZN(n1222) );
INV_X1 U886 ( .A(n1191), .ZN(n1221) );
XOR2_X1 U887 ( .A(G137), .B(n1182), .Z(G39) );
AND3_X1 U888 ( .A1(n1053), .A2(n1187), .A3(n1223), .ZN(n1182) );
XOR2_X1 U889 ( .A(G134), .B(n1181), .Z(G36) );
AND3_X1 U890 ( .A1(n1052), .A2(n1058), .A3(n1223), .ZN(n1181) );
XOR2_X1 U891 ( .A(G131), .B(n1180), .Z(G33) );
NOR2_X1 U892 ( .A1(n1191), .A2(n1196), .ZN(n1180) );
INV_X1 U893 ( .A(n1058), .ZN(n1196) );
NAND2_X1 U894 ( .A1(n1223), .A2(n1051), .ZN(n1191) );
AND3_X1 U895 ( .A1(n1059), .A2(n1193), .A3(n1037), .ZN(n1223) );
NOR2_X1 U896 ( .A1(n1224), .A2(n1035), .ZN(n1037) );
XOR2_X1 U897 ( .A(G128), .B(n1189), .Z(G30) );
NOR2_X1 U898 ( .A1(n1188), .A2(n1225), .ZN(n1189) );
INV_X1 U899 ( .A(n1187), .ZN(n1225) );
NAND3_X1 U900 ( .A1(n1213), .A2(n1193), .A3(n1052), .ZN(n1188) );
XNOR2_X1 U901 ( .A(G101), .B(n1204), .ZN(G3) );
NAND3_X1 U902 ( .A1(n1202), .A2(n1058), .A3(n1053), .ZN(n1204) );
AND2_X1 U903 ( .A1(n1213), .A2(n1226), .ZN(n1202) );
AND2_X1 U904 ( .A1(n1059), .A2(n1227), .ZN(n1213) );
XOR2_X1 U905 ( .A(n1228), .B(G125), .Z(G27) );
NAND2_X1 U906 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NAND2_X1 U907 ( .A1(n1179), .A2(n1231), .ZN(n1230) );
INV_X1 U908 ( .A(KEYINPUT14), .ZN(n1231) );
AND2_X1 U909 ( .A1(n1232), .A2(n1061), .ZN(n1179) );
NAND3_X1 U910 ( .A1(n1232), .A2(n1190), .A3(KEYINPUT14), .ZN(n1229) );
INV_X1 U911 ( .A(n1061), .ZN(n1190) );
AND4_X1 U912 ( .A1(n1051), .A2(n1030), .A3(n1227), .A4(n1193), .ZN(n1232) );
NAND2_X1 U913 ( .A1(n1064), .A2(n1233), .ZN(n1193) );
NAND4_X1 U914 ( .A1(G902), .A2(G953), .A3(n1234), .A4(n1235), .ZN(n1233) );
INV_X1 U915 ( .A(G900), .ZN(n1235) );
XNOR2_X1 U916 ( .A(G122), .B(n1203), .ZN(G24) );
NAND4_X1 U917 ( .A1(n1236), .A2(n1049), .A3(n1216), .A4(n1079), .ZN(n1203) );
XNOR2_X1 U918 ( .A(G119), .B(n1201), .ZN(G21) );
NAND3_X1 U919 ( .A1(n1236), .A2(n1187), .A3(n1053), .ZN(n1201) );
NAND2_X1 U920 ( .A1(n1237), .A2(n1238), .ZN(n1187) );
NAND2_X1 U921 ( .A1(n1061), .A2(n1239), .ZN(n1238) );
NAND3_X1 U922 ( .A1(n1075), .A2(n1240), .A3(KEYINPUT32), .ZN(n1237) );
XOR2_X1 U923 ( .A(G116), .B(n1241), .Z(G18) );
NOR2_X1 U924 ( .A1(KEYINPUT44), .A2(n1200), .ZN(n1241) );
NAND3_X1 U925 ( .A1(n1052), .A2(n1058), .A3(n1236), .ZN(n1200) );
NOR2_X1 U926 ( .A1(n1079), .A2(n1070), .ZN(n1052) );
XNOR2_X1 U927 ( .A(G113), .B(n1199), .ZN(G15) );
NAND3_X1 U928 ( .A1(n1236), .A2(n1058), .A3(n1051), .ZN(n1199) );
AND2_X1 U929 ( .A1(n1070), .A2(n1079), .ZN(n1051) );
INV_X1 U930 ( .A(n1216), .ZN(n1070) );
NAND2_X1 U931 ( .A1(n1242), .A2(n1243), .ZN(n1058) );
NAND2_X1 U932 ( .A1(n1049), .A2(n1239), .ZN(n1243) );
INV_X1 U933 ( .A(KEYINPUT32), .ZN(n1239) );
NOR2_X1 U934 ( .A1(n1075), .A2(n1240), .ZN(n1049) );
INV_X1 U935 ( .A(n1244), .ZN(n1240) );
NAND3_X1 U936 ( .A1(n1244), .A2(n1075), .A3(KEYINPUT32), .ZN(n1242) );
AND3_X1 U937 ( .A1(n1227), .A2(n1226), .A3(n1030), .ZN(n1236) );
AND2_X1 U938 ( .A1(n1043), .A2(n1245), .ZN(n1030) );
XNOR2_X1 U939 ( .A(G110), .B(n1246), .ZN(G12) );
NAND4_X1 U940 ( .A1(n1053), .A2(n1061), .A3(n1247), .A4(n1248), .ZN(n1246) );
NOR3_X1 U941 ( .A1(n1033), .A2(KEYINPUT13), .A3(n1249), .ZN(n1248) );
INV_X1 U942 ( .A(n1226), .ZN(n1249) );
NAND2_X1 U943 ( .A1(n1250), .A2(n1064), .ZN(n1226) );
NAND3_X1 U944 ( .A1(n1234), .A2(n1096), .A3(G952), .ZN(n1064) );
NAND3_X1 U945 ( .A1(n1112), .A2(n1234), .A3(G902), .ZN(n1250) );
NAND2_X1 U946 ( .A1(G237), .A2(G234), .ZN(n1234) );
NOR2_X1 U947 ( .A1(n1096), .A2(G898), .ZN(n1112) );
INV_X1 U948 ( .A(n1227), .ZN(n1033) );
NOR2_X1 U949 ( .A1(n1036), .A2(n1035), .ZN(n1227) );
AND2_X1 U950 ( .A1(G214), .A2(n1251), .ZN(n1035) );
INV_X1 U951 ( .A(n1224), .ZN(n1036) );
XNOR2_X1 U952 ( .A(n1252), .B(n1173), .ZN(n1224) );
AND2_X1 U953 ( .A1(G210), .A2(n1251), .ZN(n1173) );
NAND2_X1 U954 ( .A1(n1174), .A2(n1253), .ZN(n1251) );
INV_X1 U955 ( .A(G237), .ZN(n1253) );
NAND2_X1 U956 ( .A1(n1254), .A2(n1174), .ZN(n1252) );
XOR2_X1 U957 ( .A(n1255), .B(n1256), .Z(n1254) );
XNOR2_X1 U958 ( .A(n1172), .B(n1257), .ZN(n1256) );
XNOR2_X1 U959 ( .A(KEYINPUT55), .B(KEYINPUT50), .ZN(n1257) );
AND2_X1 U960 ( .A1(G224), .A2(n1096), .ZN(n1172) );
XOR2_X1 U961 ( .A(n1206), .B(n1258), .Z(n1255) );
NOR3_X1 U962 ( .A1(n1208), .A2(n1259), .A3(n1260), .ZN(n1258) );
NOR2_X1 U963 ( .A1(KEYINPUT54), .A2(n1261), .ZN(n1260) );
NOR2_X1 U964 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
AND2_X1 U965 ( .A1(n1144), .A2(KEYINPUT30), .ZN(n1263) );
NOR3_X1 U966 ( .A1(KEYINPUT30), .A2(n1144), .A3(n1212), .ZN(n1262) );
NOR2_X1 U967 ( .A1(n1264), .A2(n1265), .ZN(n1259) );
INV_X1 U968 ( .A(KEYINPUT54), .ZN(n1265) );
NOR2_X1 U969 ( .A1(n1212), .A2(n1266), .ZN(n1264) );
XNOR2_X1 U970 ( .A(KEYINPUT30), .B(n1093), .ZN(n1266) );
AND2_X1 U971 ( .A1(n1212), .A2(n1144), .ZN(n1208) );
XNOR2_X1 U972 ( .A(G125), .B(KEYINPUT42), .ZN(n1212) );
XOR2_X1 U973 ( .A(n1114), .B(n1267), .Z(n1206) );
NOR2_X1 U974 ( .A1(KEYINPUT46), .A2(n1113), .ZN(n1267) );
NAND2_X1 U975 ( .A1(n1268), .A2(n1269), .ZN(n1113) );
NAND2_X1 U976 ( .A1(G122), .A2(n1270), .ZN(n1269) );
XOR2_X1 U977 ( .A(n1271), .B(KEYINPUT9), .Z(n1268) );
OR2_X1 U978 ( .A1(n1270), .A2(G122), .ZN(n1271) );
XOR2_X1 U979 ( .A(n1272), .B(n1273), .Z(n1114) );
XOR2_X1 U980 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U981 ( .A(KEYINPUT21), .B(n1276), .ZN(n1275) );
XOR2_X1 U982 ( .A(n1277), .B(n1278), .Z(n1272) );
NAND2_X1 U983 ( .A1(n1279), .A2(n1280), .ZN(n1277) );
NAND2_X1 U984 ( .A1(KEYINPUT38), .A2(n1281), .ZN(n1280) );
OR3_X1 U985 ( .A1(n1282), .A2(G107), .A3(KEYINPUT38), .ZN(n1279) );
XNOR2_X1 U986 ( .A(n1059), .B(KEYINPUT26), .ZN(n1247) );
NOR2_X1 U987 ( .A1(n1043), .A2(n1044), .ZN(n1059) );
INV_X1 U988 ( .A(n1245), .ZN(n1044) );
NAND2_X1 U989 ( .A1(G221), .A2(n1283), .ZN(n1245) );
XOR2_X1 U990 ( .A(n1284), .B(n1080), .Z(n1043) );
NAND2_X1 U991 ( .A1(n1285), .A2(n1174), .ZN(n1080) );
XOR2_X1 U992 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U993 ( .A(n1154), .B(n1164), .ZN(n1287) );
XOR2_X1 U994 ( .A(n1281), .B(n1278), .Z(n1164) );
XNOR2_X1 U995 ( .A(n1135), .B(KEYINPUT28), .ZN(n1278) );
XNOR2_X1 U996 ( .A(G104), .B(G107), .ZN(n1281) );
INV_X1 U997 ( .A(n1157), .ZN(n1154) );
XOR2_X1 U998 ( .A(G110), .B(n1288), .Z(n1157) );
XNOR2_X1 U999 ( .A(n1289), .B(n1290), .ZN(n1286) );
XOR2_X1 U1000 ( .A(n1291), .B(n1160), .Z(n1289) );
AND2_X1 U1001 ( .A1(G227), .A2(n1096), .ZN(n1160) );
NAND2_X1 U1002 ( .A1(n1292), .A2(KEYINPUT36), .ZN(n1291) );
XNOR2_X1 U1003 ( .A(n1093), .B(KEYINPUT51), .ZN(n1292) );
NAND2_X1 U1004 ( .A1(KEYINPUT63), .A2(n1081), .ZN(n1284) );
XNOR2_X1 U1005 ( .A(G469), .B(KEYINPUT61), .ZN(n1081) );
NOR2_X1 U1006 ( .A1(n1244), .A2(n1075), .ZN(n1061) );
XNOR2_X1 U1007 ( .A(n1293), .B(G472), .ZN(n1075) );
NAND2_X1 U1008 ( .A1(n1174), .A2(n1294), .ZN(n1293) );
NAND2_X1 U1009 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
NAND2_X1 U1010 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XOR2_X1 U1011 ( .A(n1299), .B(KEYINPUT20), .Z(n1295) );
OR2_X1 U1012 ( .A1(n1298), .A2(n1297), .ZN(n1299) );
XNOR2_X1 U1013 ( .A(n1136), .B(n1300), .ZN(n1297) );
XOR2_X1 U1014 ( .A(KEYINPUT23), .B(n1141), .Z(n1300) );
XNOR2_X1 U1015 ( .A(n1290), .B(n1301), .ZN(n1141) );
XNOR2_X1 U1016 ( .A(KEYINPUT31), .B(n1144), .ZN(n1301) );
INV_X1 U1017 ( .A(n1093), .ZN(n1144) );
XOR2_X1 U1018 ( .A(G146), .B(n1302), .Z(n1093) );
INV_X1 U1019 ( .A(n1162), .ZN(n1290) );
XNOR2_X1 U1020 ( .A(G134), .B(n1094), .ZN(n1162) );
XNOR2_X1 U1021 ( .A(G131), .B(G137), .ZN(n1094) );
XOR2_X1 U1022 ( .A(G113), .B(n1303), .Z(n1136) );
NOR3_X1 U1023 ( .A1(KEYINPUT43), .A2(n1304), .A3(n1305), .ZN(n1303) );
NOR3_X1 U1024 ( .A1(n1306), .A2(G116), .A3(n1307), .ZN(n1305) );
INV_X1 U1025 ( .A(KEYINPUT7), .ZN(n1306) );
NOR2_X1 U1026 ( .A1(KEYINPUT7), .A2(n1274), .ZN(n1304) );
XOR2_X1 U1027 ( .A(G116), .B(G119), .Z(n1274) );
XNOR2_X1 U1028 ( .A(n1135), .B(n1308), .ZN(n1298) );
NOR2_X1 U1029 ( .A1(KEYINPUT45), .A2(n1139), .ZN(n1308) );
NAND2_X1 U1030 ( .A1(G210), .A2(n1309), .ZN(n1139) );
XNOR2_X1 U1031 ( .A(G101), .B(KEYINPUT35), .ZN(n1135) );
XOR2_X1 U1032 ( .A(n1078), .B(n1310), .Z(n1244) );
NOR2_X1 U1033 ( .A1(n1121), .A2(KEYINPUT33), .ZN(n1310) );
INV_X1 U1034 ( .A(n1077), .ZN(n1121) );
NAND2_X1 U1035 ( .A1(G217), .A2(n1283), .ZN(n1077) );
NAND2_X1 U1036 ( .A1(G234), .A2(n1174), .ZN(n1283) );
NOR2_X1 U1037 ( .A1(n1120), .A2(G902), .ZN(n1078) );
XOR2_X1 U1038 ( .A(n1311), .B(n1312), .Z(n1120) );
XOR2_X1 U1039 ( .A(n1313), .B(n1314), .Z(n1312) );
XNOR2_X1 U1040 ( .A(G128), .B(n1307), .ZN(n1314) );
INV_X1 U1041 ( .A(G119), .ZN(n1307) );
XNOR2_X1 U1042 ( .A(n1315), .B(G137), .ZN(n1313) );
XOR2_X1 U1043 ( .A(n1088), .B(n1316), .Z(n1311) );
XOR2_X1 U1044 ( .A(n1317), .B(n1318), .Z(n1316) );
NAND2_X1 U1045 ( .A1(KEYINPUT58), .A2(n1270), .ZN(n1318) );
INV_X1 U1046 ( .A(G110), .ZN(n1270) );
NAND3_X1 U1047 ( .A1(G221), .A2(n1096), .A3(G234), .ZN(n1317) );
NOR2_X1 U1048 ( .A1(n1216), .A2(n1079), .ZN(n1053) );
XNOR2_X1 U1049 ( .A(n1319), .B(G475), .ZN(n1079) );
NAND2_X1 U1050 ( .A1(n1130), .A2(n1174), .ZN(n1319) );
XOR2_X1 U1051 ( .A(n1320), .B(n1321), .Z(n1130) );
XOR2_X1 U1052 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1053 ( .A(n1324), .B(n1325), .ZN(n1323) );
NOR2_X1 U1054 ( .A1(KEYINPUT16), .A2(n1276), .ZN(n1325) );
INV_X1 U1055 ( .A(G113), .ZN(n1276) );
NOR2_X1 U1056 ( .A1(KEYINPUT11), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1057 ( .A(n1327), .B(n1088), .Z(n1326) );
XNOR2_X1 U1058 ( .A(G125), .B(n1288), .ZN(n1088) );
XOR2_X1 U1059 ( .A(G140), .B(KEYINPUT3), .Z(n1288) );
NAND2_X1 U1060 ( .A1(KEYINPUT5), .A2(n1315), .ZN(n1327) );
INV_X1 U1061 ( .A(G146), .ZN(n1315) );
NAND2_X1 U1062 ( .A1(G214), .A2(n1309), .ZN(n1322) );
NOR2_X1 U1063 ( .A1(G953), .A2(G237), .ZN(n1309) );
XOR2_X1 U1064 ( .A(n1328), .B(n1329), .Z(n1320) );
XNOR2_X1 U1065 ( .A(G122), .B(n1282), .ZN(n1329) );
INV_X1 U1066 ( .A(G104), .ZN(n1282) );
XNOR2_X1 U1067 ( .A(G131), .B(G143), .ZN(n1328) );
XNOR2_X1 U1068 ( .A(n1330), .B(G478), .ZN(n1216) );
NAND2_X1 U1069 ( .A1(n1127), .A2(n1174), .ZN(n1330) );
INV_X1 U1070 ( .A(G902), .ZN(n1174) );
XOR2_X1 U1071 ( .A(n1331), .B(n1332), .Z(n1127) );
XOR2_X1 U1072 ( .A(n1333), .B(n1334), .Z(n1332) );
NOR2_X1 U1073 ( .A1(KEYINPUT22), .A2(n1335), .ZN(n1334) );
XNOR2_X1 U1074 ( .A(G107), .B(n1336), .ZN(n1335) );
XOR2_X1 U1075 ( .A(G122), .B(G116), .Z(n1336) );
NOR2_X1 U1076 ( .A1(G134), .A2(n1337), .ZN(n1333) );
XOR2_X1 U1077 ( .A(KEYINPUT59), .B(KEYINPUT25), .Z(n1337) );
XOR2_X1 U1078 ( .A(n1338), .B(n1302), .Z(n1331) );
XOR2_X1 U1079 ( .A(G128), .B(G143), .Z(n1302) );
NAND3_X1 U1080 ( .A1(G234), .A2(n1096), .A3(G217), .ZN(n1338) );
INV_X1 U1081 ( .A(G953), .ZN(n1096) );
endmodule


