//Key = 0101000001000111001110111101011110110100111011100101001100100101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368;

XOR2_X1 U766 ( .A(G107), .B(n1053), .Z(G9) );
NOR2_X1 U767 ( .A1(n1054), .A2(n1055), .ZN(G75) );
XOR2_X1 U768 ( .A(n1056), .B(KEYINPUT51), .Z(n1055) );
NAND4_X1 U769 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
NOR2_X1 U770 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
XNOR2_X1 U771 ( .A(KEYINPUT3), .B(n1063), .ZN(n1059) );
NAND2_X1 U772 ( .A1(n1064), .A2(n1065), .ZN(n1057) );
NAND2_X1 U773 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND4_X1 U774 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1067) );
OR2_X1 U775 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U776 ( .A1(n1074), .A2(n1075), .ZN(n1066) );
NAND2_X1 U777 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND3_X1 U778 ( .A1(n1069), .A2(n1078), .A3(n1068), .ZN(n1077) );
NAND2_X1 U779 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U780 ( .A1(n1070), .A2(n1081), .ZN(n1076) );
NAND3_X1 U781 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NAND2_X1 U782 ( .A1(n1085), .A2(n1068), .ZN(n1084) );
XNOR2_X1 U783 ( .A(n1086), .B(n1087), .ZN(n1085) );
NOR2_X1 U784 ( .A1(KEYINPUT11), .A2(n1088), .ZN(n1087) );
NAND3_X1 U785 ( .A1(n1069), .A2(n1089), .A3(n1090), .ZN(n1082) );
INV_X1 U786 ( .A(n1091), .ZN(n1064) );
AND3_X1 U787 ( .A1(n1058), .A2(n1063), .A3(n1061), .ZN(n1054) );
INV_X1 U788 ( .A(G952), .ZN(n1061) );
NAND4_X1 U789 ( .A1(n1092), .A2(n1069), .A3(n1093), .A4(n1094), .ZN(n1058) );
NOR4_X1 U790 ( .A1(n1095), .A2(n1090), .A3(n1096), .A4(n1097), .ZN(n1094) );
INV_X1 U791 ( .A(n1098), .ZN(n1095) );
NOR4_X1 U792 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1093) );
NOR3_X1 U793 ( .A1(G472), .A2(G902), .A3(n1103), .ZN(n1102) );
NOR2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(n1101) );
NOR2_X1 U795 ( .A1(G902), .A2(n1103), .ZN(n1104) );
NOR3_X1 U796 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1100) );
INV_X1 U797 ( .A(KEYINPUT63), .ZN(n1106) );
NOR2_X1 U798 ( .A1(KEYINPUT63), .A2(G475), .ZN(n1099) );
XNOR2_X1 U799 ( .A(n1109), .B(KEYINPUT12), .ZN(n1092) );
XOR2_X1 U800 ( .A(n1110), .B(n1111), .Z(G72) );
NOR2_X1 U801 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XOR2_X1 U802 ( .A(n1114), .B(KEYINPUT15), .Z(n1113) );
NAND4_X1 U803 ( .A1(n1115), .A2(n1116), .A3(n1117), .A4(n1118), .ZN(n1114) );
NAND2_X1 U804 ( .A1(G953), .A2(n1119), .ZN(n1117) );
NOR3_X1 U805 ( .A1(n1115), .A2(G953), .A3(n1120), .ZN(n1112) );
NOR2_X1 U806 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XNOR2_X1 U807 ( .A(n1123), .B(n1124), .ZN(n1115) );
XOR2_X1 U808 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND2_X1 U809 ( .A1(KEYINPUT44), .A2(n1127), .ZN(n1125) );
XNOR2_X1 U810 ( .A(n1128), .B(n1129), .ZN(n1123) );
NAND2_X1 U811 ( .A1(G953), .A2(n1130), .ZN(n1110) );
NAND2_X1 U812 ( .A1(G900), .A2(G227), .ZN(n1130) );
XOR2_X1 U813 ( .A(n1131), .B(n1132), .Z(G69) );
NAND2_X1 U814 ( .A1(G953), .A2(n1133), .ZN(n1132) );
NAND2_X1 U815 ( .A1(G898), .A2(G224), .ZN(n1133) );
NAND2_X1 U816 ( .A1(n1134), .A2(n1135), .ZN(n1131) );
NAND2_X1 U817 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U818 ( .A1(KEYINPUT18), .A2(n1138), .ZN(n1137) );
NAND2_X1 U819 ( .A1(KEYINPUT27), .A2(n1139), .ZN(n1138) );
INV_X1 U820 ( .A(n1140), .ZN(n1139) );
INV_X1 U821 ( .A(n1141), .ZN(n1136) );
NAND2_X1 U822 ( .A1(n1142), .A2(n1140), .ZN(n1134) );
NAND2_X1 U823 ( .A1(n1143), .A2(n1144), .ZN(n1140) );
NAND2_X1 U824 ( .A1(G953), .A2(n1145), .ZN(n1144) );
XOR2_X1 U825 ( .A(n1146), .B(n1147), .Z(n1143) );
XOR2_X1 U826 ( .A(KEYINPUT28), .B(n1148), .Z(n1147) );
NOR2_X1 U827 ( .A1(KEYINPUT16), .A2(n1149), .ZN(n1148) );
NAND2_X1 U828 ( .A1(KEYINPUT27), .A2(n1150), .ZN(n1142) );
NAND2_X1 U829 ( .A1(KEYINPUT18), .A2(n1141), .ZN(n1150) );
NAND2_X1 U830 ( .A1(n1063), .A2(n1151), .ZN(n1141) );
NAND2_X1 U831 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NOR2_X1 U832 ( .A1(n1154), .A2(n1155), .ZN(G66) );
XOR2_X1 U833 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U834 ( .A(KEYINPUT45), .B(n1158), .Z(n1157) );
NOR2_X1 U835 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U836 ( .A1(n1154), .A2(n1161), .ZN(G63) );
XOR2_X1 U837 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U838 ( .A1(n1164), .A2(n1160), .ZN(n1162) );
NOR2_X1 U839 ( .A1(n1154), .A2(n1165), .ZN(G60) );
XOR2_X1 U840 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U841 ( .A1(n1108), .A2(n1160), .ZN(n1166) );
NAND2_X1 U842 ( .A1(n1168), .A2(n1169), .ZN(G6) );
OR2_X1 U843 ( .A1(n1170), .A2(G104), .ZN(n1169) );
XOR2_X1 U844 ( .A(n1171), .B(KEYINPUT48), .Z(n1168) );
NAND2_X1 U845 ( .A1(G104), .A2(n1170), .ZN(n1171) );
NOR2_X1 U846 ( .A1(n1154), .A2(n1172), .ZN(G57) );
XOR2_X1 U847 ( .A(n1173), .B(n1103), .Z(n1172) );
NOR2_X1 U848 ( .A1(n1105), .A2(n1160), .ZN(n1173) );
INV_X1 U849 ( .A(G472), .ZN(n1105) );
NOR2_X1 U850 ( .A1(n1154), .A2(n1174), .ZN(G54) );
XOR2_X1 U851 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U852 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U853 ( .A(n1179), .B(n1180), .Z(n1175) );
XNOR2_X1 U854 ( .A(G110), .B(n1181), .ZN(n1179) );
NOR3_X1 U855 ( .A1(n1160), .A2(KEYINPUT36), .A3(n1182), .ZN(n1181) );
NOR2_X1 U856 ( .A1(n1154), .A2(n1183), .ZN(G51) );
XOR2_X1 U857 ( .A(n1184), .B(n1185), .Z(n1183) );
XOR2_X1 U858 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U859 ( .A1(n1188), .A2(n1160), .ZN(n1187) );
NAND2_X1 U860 ( .A1(G902), .A2(n1062), .ZN(n1160) );
NAND4_X1 U861 ( .A1(n1189), .A2(n1190), .A3(n1152), .A4(n1116), .ZN(n1062) );
INV_X1 U862 ( .A(n1122), .ZN(n1116) );
NAND4_X1 U863 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1122) );
NOR4_X1 U864 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1194) );
NOR3_X1 U865 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1198) );
XNOR2_X1 U866 ( .A(KEYINPUT23), .B(n1202), .ZN(n1199) );
NOR3_X1 U867 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1196) );
INV_X1 U868 ( .A(KEYINPUT8), .ZN(n1205) );
NOR2_X1 U869 ( .A1(n1206), .A2(n1079), .ZN(n1195) );
NOR2_X1 U870 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NOR2_X1 U871 ( .A1(KEYINPUT8), .A2(n1204), .ZN(n1208) );
AND3_X1 U872 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1207) );
AND4_X1 U873 ( .A1(n1170), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1152) );
NOR4_X1 U874 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1053), .ZN(n1214) );
AND3_X1 U875 ( .A1(n1070), .A2(n1072), .A3(n1218), .ZN(n1053) );
NAND2_X1 U876 ( .A1(n1219), .A2(n1210), .ZN(n1213) );
XOR2_X1 U877 ( .A(n1220), .B(KEYINPUT31), .Z(n1219) );
NAND3_X1 U878 ( .A1(n1218), .A2(n1070), .A3(n1073), .ZN(n1170) );
XOR2_X1 U879 ( .A(n1153), .B(KEYINPUT47), .Z(n1190) );
XNOR2_X1 U880 ( .A(n1121), .B(KEYINPUT39), .ZN(n1189) );
NOR2_X1 U881 ( .A1(KEYINPUT2), .A2(n1221), .ZN(n1186) );
XOR2_X1 U882 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR2_X1 U883 ( .A1(KEYINPUT57), .A2(n1224), .ZN(n1223) );
NOR2_X1 U884 ( .A1(n1063), .A2(G952), .ZN(n1154) );
XNOR2_X1 U885 ( .A(n1121), .B(n1225), .ZN(G48) );
XNOR2_X1 U886 ( .A(G146), .B(KEYINPUT60), .ZN(n1225) );
INV_X1 U887 ( .A(n1118), .ZN(n1121) );
NAND3_X1 U888 ( .A1(n1073), .A2(n1210), .A3(n1226), .ZN(n1118) );
XNOR2_X1 U889 ( .A(G143), .B(n1227), .ZN(G45) );
NAND4_X1 U890 ( .A1(n1228), .A2(n1209), .A3(n1203), .A4(n1211), .ZN(n1227) );
XNOR2_X1 U891 ( .A(n1210), .B(KEYINPUT34), .ZN(n1228) );
XOR2_X1 U892 ( .A(G140), .B(n1197), .Z(G42) );
NOR2_X1 U893 ( .A1(n1204), .A2(n1080), .ZN(n1197) );
XOR2_X1 U894 ( .A(G137), .B(n1229), .Z(G39) );
NOR4_X1 U895 ( .A1(KEYINPUT21), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1229) );
NAND2_X1 U896 ( .A1(n1230), .A2(n1231), .ZN(G36) );
NAND2_X1 U897 ( .A1(G134), .A2(n1193), .ZN(n1231) );
XOR2_X1 U898 ( .A(KEYINPUT24), .B(n1232), .Z(n1230) );
NOR2_X1 U899 ( .A1(G134), .A2(n1193), .ZN(n1232) );
NAND4_X1 U900 ( .A1(n1068), .A2(n1209), .A3(n1203), .A4(n1072), .ZN(n1193) );
XOR2_X1 U901 ( .A(n1233), .B(n1234), .Z(G33) );
NOR2_X1 U902 ( .A1(n1079), .A2(n1204), .ZN(n1234) );
NAND3_X1 U903 ( .A1(n1209), .A2(n1073), .A3(n1068), .ZN(n1204) );
INV_X1 U904 ( .A(n1202), .ZN(n1068) );
NAND2_X1 U905 ( .A1(n1089), .A2(n1235), .ZN(n1202) );
INV_X1 U906 ( .A(n1203), .ZN(n1079) );
NOR2_X1 U907 ( .A1(KEYINPUT0), .A2(n1127), .ZN(n1233) );
INV_X1 U908 ( .A(G131), .ZN(n1127) );
XNOR2_X1 U909 ( .A(n1236), .B(n1191), .ZN(G30) );
NAND3_X1 U910 ( .A1(n1210), .A2(n1072), .A3(n1226), .ZN(n1191) );
INV_X1 U911 ( .A(n1201), .ZN(n1226) );
NAND3_X1 U912 ( .A1(n1237), .A2(n1109), .A3(n1209), .ZN(n1201) );
AND3_X1 U913 ( .A1(n1238), .A2(n1239), .A3(n1088), .ZN(n1209) );
NAND2_X1 U914 ( .A1(KEYINPUT35), .A2(n1240), .ZN(n1236) );
XOR2_X1 U915 ( .A(n1212), .B(n1241), .Z(G3) );
NAND2_X1 U916 ( .A1(KEYINPUT25), .A2(G101), .ZN(n1241) );
NAND3_X1 U917 ( .A1(n1203), .A2(n1218), .A3(n1074), .ZN(n1212) );
NOR4_X1 U918 ( .A1(n1242), .A2(n1243), .A3(n1086), .A4(n1244), .ZN(n1218) );
XNOR2_X1 U919 ( .A(n1192), .B(n1245), .ZN(G27) );
NOR2_X1 U920 ( .A1(KEYINPUT59), .A2(n1246), .ZN(n1245) );
NAND4_X1 U921 ( .A1(n1247), .A2(n1073), .A3(n1248), .A4(n1238), .ZN(n1192) );
NAND2_X1 U922 ( .A1(n1091), .A2(n1249), .ZN(n1238) );
NAND4_X1 U923 ( .A1(G953), .A2(G902), .A3(n1250), .A4(n1119), .ZN(n1249) );
INV_X1 U924 ( .A(G900), .ZN(n1119) );
INV_X1 U925 ( .A(n1083), .ZN(n1248) );
XOR2_X1 U926 ( .A(G122), .B(n1217), .Z(G24) );
AND3_X1 U927 ( .A1(n1070), .A2(n1211), .A3(n1251), .ZN(n1217) );
NOR2_X1 U928 ( .A1(n1109), .A2(n1237), .ZN(n1070) );
XOR2_X1 U929 ( .A(G119), .B(n1216), .Z(G21) );
AND4_X1 U930 ( .A1(n1074), .A2(n1251), .A3(n1237), .A4(n1109), .ZN(n1216) );
XNOR2_X1 U931 ( .A(G116), .B(n1153), .ZN(G18) );
NAND3_X1 U932 ( .A1(n1251), .A2(n1072), .A3(n1203), .ZN(n1153) );
NAND2_X1 U933 ( .A1(n1252), .A2(n1253), .ZN(n1072) );
OR3_X1 U934 ( .A1(n1254), .A2(n1255), .A3(KEYINPUT6), .ZN(n1253) );
NAND2_X1 U935 ( .A1(KEYINPUT6), .A2(n1211), .ZN(n1252) );
NOR2_X1 U936 ( .A1(n1255), .A2(n1256), .ZN(n1211) );
XOR2_X1 U937 ( .A(G113), .B(n1215), .Z(G15) );
AND3_X1 U938 ( .A1(n1203), .A2(n1251), .A3(n1073), .ZN(n1215) );
NOR2_X1 U939 ( .A1(n1096), .A2(n1256), .ZN(n1073) );
INV_X1 U940 ( .A(n1254), .ZN(n1256) );
NOR2_X1 U941 ( .A1(n1083), .A2(n1244), .ZN(n1251) );
NAND2_X1 U942 ( .A1(n1069), .A2(n1210), .ZN(n1083) );
NOR2_X1 U943 ( .A1(n1088), .A2(n1086), .ZN(n1069) );
NOR2_X1 U944 ( .A1(n1109), .A2(n1257), .ZN(n1203) );
XNOR2_X1 U945 ( .A(n1258), .B(n1259), .ZN(G12) );
NOR2_X1 U946 ( .A1(n1242), .A2(n1220), .ZN(n1259) );
NAND3_X1 U947 ( .A1(n1247), .A2(n1074), .A3(n1260), .ZN(n1220) );
NOR3_X1 U948 ( .A1(n1243), .A2(n1244), .A3(n1086), .ZN(n1260) );
INV_X1 U949 ( .A(n1239), .ZN(n1086) );
NAND2_X1 U950 ( .A1(G221), .A2(n1261), .ZN(n1239) );
AND2_X1 U951 ( .A1(n1091), .A2(n1262), .ZN(n1244) );
NAND4_X1 U952 ( .A1(G953), .A2(G902), .A3(n1250), .A4(n1145), .ZN(n1262) );
INV_X1 U953 ( .A(G898), .ZN(n1145) );
NAND3_X1 U954 ( .A1(n1250), .A2(n1063), .A3(G952), .ZN(n1091) );
NAND2_X1 U955 ( .A1(G237), .A2(n1263), .ZN(n1250) );
INV_X1 U956 ( .A(n1088), .ZN(n1243) );
XOR2_X1 U957 ( .A(n1264), .B(n1182), .Z(n1088) );
INV_X1 U958 ( .A(G469), .ZN(n1182) );
NAND2_X1 U959 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
XOR2_X1 U960 ( .A(n1267), .B(n1268), .Z(n1265) );
NOR2_X1 U961 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
AND3_X1 U962 ( .A1(KEYINPUT7), .A2(n1128), .A3(n1271), .ZN(n1270) );
NOR2_X1 U963 ( .A1(KEYINPUT7), .A2(n1178), .ZN(n1269) );
XNOR2_X1 U964 ( .A(n1128), .B(n1271), .ZN(n1178) );
XNOR2_X1 U965 ( .A(n1272), .B(n1273), .ZN(n1271) );
NOR2_X1 U966 ( .A1(KEYINPUT38), .A2(n1274), .ZN(n1273) );
XNOR2_X1 U967 ( .A(G101), .B(G107), .ZN(n1272) );
NAND2_X1 U968 ( .A1(n1275), .A2(n1276), .ZN(n1128) );
NAND2_X1 U969 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
XOR2_X1 U970 ( .A(KEYINPUT55), .B(n1279), .Z(n1277) );
NAND2_X1 U971 ( .A1(n1279), .A2(G146), .ZN(n1275) );
XOR2_X1 U972 ( .A(n1280), .B(n1177), .Z(n1267) );
XNOR2_X1 U973 ( .A(n1281), .B(KEYINPUT13), .ZN(n1177) );
NAND2_X1 U974 ( .A1(n1282), .A2(n1283), .ZN(n1280) );
OR2_X1 U975 ( .A1(n1258), .A2(n1180), .ZN(n1283) );
NAND2_X1 U976 ( .A1(n1284), .A2(n1258), .ZN(n1282) );
XNOR2_X1 U977 ( .A(n1180), .B(KEYINPUT1), .ZN(n1284) );
XOR2_X1 U978 ( .A(G140), .B(n1285), .Z(n1180) );
AND2_X1 U979 ( .A1(n1063), .A2(G227), .ZN(n1285) );
INV_X1 U980 ( .A(n1200), .ZN(n1074) );
NAND2_X1 U981 ( .A1(n1255), .A2(n1286), .ZN(n1200) );
XNOR2_X1 U982 ( .A(KEYINPUT6), .B(n1254), .ZN(n1286) );
NAND3_X1 U983 ( .A1(n1287), .A2(n1288), .A3(n1098), .ZN(n1254) );
NAND2_X1 U984 ( .A1(n1107), .A2(n1108), .ZN(n1098) );
NAND2_X1 U985 ( .A1(KEYINPUT4), .A2(n1108), .ZN(n1288) );
OR3_X1 U986 ( .A1(n1107), .A2(KEYINPUT4), .A3(n1108), .ZN(n1287) );
INV_X1 U987 ( .A(G475), .ZN(n1108) );
NOR2_X1 U988 ( .A1(n1167), .A2(G902), .ZN(n1107) );
XNOR2_X1 U989 ( .A(n1289), .B(n1290), .ZN(n1167) );
XOR2_X1 U990 ( .A(n1291), .B(n1292), .Z(n1290) );
XNOR2_X1 U991 ( .A(G104), .B(G122), .ZN(n1292) );
NAND2_X1 U992 ( .A1(n1293), .A2(n1294), .ZN(n1291) );
XNOR2_X1 U993 ( .A(KEYINPUT49), .B(KEYINPUT32), .ZN(n1293) );
XOR2_X1 U994 ( .A(n1295), .B(n1296), .Z(n1289) );
NOR2_X1 U995 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XOR2_X1 U996 ( .A(n1299), .B(KEYINPUT37), .Z(n1298) );
NAND2_X1 U997 ( .A1(n1300), .A2(G140), .ZN(n1299) );
NOR2_X1 U998 ( .A1(G140), .A2(n1300), .ZN(n1297) );
XNOR2_X1 U999 ( .A(KEYINPUT5), .B(G125), .ZN(n1300) );
XOR2_X1 U1000 ( .A(n1301), .B(n1302), .Z(n1295) );
NOR2_X1 U1001 ( .A1(KEYINPUT17), .A2(n1278), .ZN(n1302) );
NAND2_X1 U1002 ( .A1(n1303), .A2(n1304), .ZN(n1301) );
NAND2_X1 U1003 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XOR2_X1 U1004 ( .A(n1307), .B(KEYINPUT33), .Z(n1303) );
OR2_X1 U1005 ( .A1(n1306), .A2(n1305), .ZN(n1307) );
XOR2_X1 U1006 ( .A(G131), .B(KEYINPUT9), .Z(n1305) );
XNOR2_X1 U1007 ( .A(n1308), .B(G143), .ZN(n1306) );
NAND3_X1 U1008 ( .A1(n1309), .A2(n1063), .A3(G214), .ZN(n1308) );
INV_X1 U1009 ( .A(n1096), .ZN(n1255) );
XOR2_X1 U1010 ( .A(n1310), .B(n1164), .Z(n1096) );
INV_X1 U1011 ( .A(G478), .ZN(n1164) );
OR2_X1 U1012 ( .A1(n1163), .A2(G902), .ZN(n1310) );
XNOR2_X1 U1013 ( .A(n1311), .B(n1312), .ZN(n1163) );
XNOR2_X1 U1014 ( .A(n1313), .B(n1314), .ZN(n1312) );
NOR2_X1 U1015 ( .A1(KEYINPUT26), .A2(n1315), .ZN(n1314) );
XOR2_X1 U1016 ( .A(G107), .B(n1316), .Z(n1315) );
NOR2_X1 U1017 ( .A1(KEYINPUT10), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1018 ( .A(G122), .B(n1318), .ZN(n1317) );
NOR2_X1 U1019 ( .A1(KEYINPUT53), .A2(n1319), .ZN(n1318) );
INV_X1 U1020 ( .A(G116), .ZN(n1319) );
XOR2_X1 U1021 ( .A(n1320), .B(n1279), .Z(n1311) );
XNOR2_X1 U1022 ( .A(n1240), .B(G143), .ZN(n1279) );
NAND2_X1 U1023 ( .A1(n1321), .A2(G217), .ZN(n1320) );
INV_X1 U1024 ( .A(n1080), .ZN(n1247) );
NAND2_X1 U1025 ( .A1(n1257), .A2(n1109), .ZN(n1080) );
XOR2_X1 U1026 ( .A(n1322), .B(n1159), .Z(n1109) );
NAND2_X1 U1027 ( .A1(G217), .A2(n1261), .ZN(n1159) );
NAND2_X1 U1028 ( .A1(n1263), .A2(n1266), .ZN(n1261) );
XNOR2_X1 U1029 ( .A(G234), .B(KEYINPUT46), .ZN(n1263) );
NAND2_X1 U1030 ( .A1(n1156), .A2(n1266), .ZN(n1322) );
XNOR2_X1 U1031 ( .A(n1323), .B(n1324), .ZN(n1156) );
XNOR2_X1 U1032 ( .A(G137), .B(n1325), .ZN(n1324) );
NAND2_X1 U1033 ( .A1(KEYINPUT42), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1034 ( .A(n1327), .B(n1328), .Z(n1326) );
XOR2_X1 U1035 ( .A(n1329), .B(n1330), .Z(n1328) );
NAND2_X1 U1036 ( .A1(KEYINPUT14), .A2(n1331), .ZN(n1330) );
NAND3_X1 U1037 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1329) );
NAND2_X1 U1038 ( .A1(KEYINPUT43), .A2(n1129), .ZN(n1334) );
NAND3_X1 U1039 ( .A1(n1335), .A2(n1336), .A3(G146), .ZN(n1333) );
INV_X1 U1040 ( .A(n1129), .ZN(n1335) );
NAND2_X1 U1041 ( .A1(n1337), .A2(n1278), .ZN(n1332) );
NAND2_X1 U1042 ( .A1(n1338), .A2(n1336), .ZN(n1337) );
INV_X1 U1043 ( .A(KEYINPUT43), .ZN(n1336) );
XNOR2_X1 U1044 ( .A(KEYINPUT50), .B(n1129), .ZN(n1338) );
XOR2_X1 U1045 ( .A(G140), .B(n1246), .Z(n1129) );
INV_X1 U1046 ( .A(G125), .ZN(n1246) );
XNOR2_X1 U1047 ( .A(n1240), .B(G110), .ZN(n1327) );
NAND2_X1 U1048 ( .A1(n1321), .A2(G221), .ZN(n1323) );
AND2_X1 U1049 ( .A1(G234), .A2(n1063), .ZN(n1321) );
INV_X1 U1050 ( .A(n1237), .ZN(n1257) );
XOR2_X1 U1051 ( .A(G472), .B(n1339), .Z(n1237) );
NOR3_X1 U1052 ( .A1(n1103), .A2(KEYINPUT56), .A3(G902), .ZN(n1339) );
XNOR2_X1 U1053 ( .A(n1340), .B(n1341), .ZN(n1103) );
XOR2_X1 U1054 ( .A(n1281), .B(n1224), .Z(n1341) );
XOR2_X1 U1055 ( .A(n1342), .B(G131), .Z(n1281) );
NAND3_X1 U1056 ( .A1(n1343), .A2(n1344), .A3(KEYINPUT58), .ZN(n1342) );
NAND2_X1 U1057 ( .A1(KEYINPUT41), .A2(n1126), .ZN(n1344) );
XNOR2_X1 U1058 ( .A(G134), .B(G137), .ZN(n1126) );
OR3_X1 U1059 ( .A1(n1313), .A2(G137), .A3(KEYINPUT41), .ZN(n1343) );
INV_X1 U1060 ( .A(G134), .ZN(n1313) );
XOR2_X1 U1061 ( .A(n1345), .B(n1346), .Z(n1340) );
XNOR2_X1 U1062 ( .A(G101), .B(n1347), .ZN(n1346) );
NAND3_X1 U1063 ( .A1(n1348), .A2(n1063), .A3(G210), .ZN(n1347) );
XNOR2_X1 U1064 ( .A(KEYINPUT20), .B(n1309), .ZN(n1348) );
NAND3_X1 U1065 ( .A1(n1349), .A2(n1350), .A3(n1351), .ZN(n1345) );
OR2_X1 U1066 ( .A1(n1352), .A2(n1294), .ZN(n1351) );
NAND3_X1 U1067 ( .A1(n1294), .A2(n1352), .A3(n1353), .ZN(n1350) );
NAND2_X1 U1068 ( .A1(n1354), .A2(n1355), .ZN(n1349) );
NAND2_X1 U1069 ( .A1(n1356), .A2(n1352), .ZN(n1355) );
INV_X1 U1070 ( .A(KEYINPUT62), .ZN(n1352) );
XNOR2_X1 U1071 ( .A(n1294), .B(KEYINPUT40), .ZN(n1356) );
INV_X1 U1072 ( .A(n1210), .ZN(n1242) );
NOR2_X1 U1073 ( .A1(n1089), .A2(n1090), .ZN(n1210) );
INV_X1 U1074 ( .A(n1235), .ZN(n1090) );
NAND2_X1 U1075 ( .A1(G214), .A2(n1357), .ZN(n1235) );
XOR2_X1 U1076 ( .A(n1097), .B(KEYINPUT19), .Z(n1089) );
XOR2_X1 U1077 ( .A(n1358), .B(n1188), .Z(n1097) );
NAND2_X1 U1078 ( .A1(G210), .A2(n1357), .ZN(n1188) );
NAND2_X1 U1079 ( .A1(n1309), .A2(n1266), .ZN(n1357) );
INV_X1 U1080 ( .A(G237), .ZN(n1309) );
NAND2_X1 U1081 ( .A1(n1359), .A2(n1266), .ZN(n1358) );
INV_X1 U1082 ( .A(G902), .ZN(n1266) );
XOR2_X1 U1083 ( .A(n1222), .B(n1360), .Z(n1359) );
XNOR2_X1 U1084 ( .A(n1184), .B(n1224), .ZN(n1360) );
XOR2_X1 U1085 ( .A(n1361), .B(n1362), .Z(n1224) );
XNOR2_X1 U1086 ( .A(n1278), .B(G143), .ZN(n1362) );
INV_X1 U1087 ( .A(G146), .ZN(n1278) );
NAND2_X1 U1088 ( .A1(KEYINPUT61), .A2(n1240), .ZN(n1361) );
INV_X1 U1089 ( .A(G128), .ZN(n1240) );
XOR2_X1 U1090 ( .A(n1146), .B(n1149), .Z(n1184) );
XOR2_X1 U1091 ( .A(G122), .B(G110), .Z(n1149) );
XOR2_X1 U1092 ( .A(n1363), .B(n1364), .Z(n1146) );
XOR2_X1 U1093 ( .A(n1365), .B(n1366), .Z(n1364) );
XNOR2_X1 U1094 ( .A(G101), .B(KEYINPUT22), .ZN(n1366) );
NAND2_X1 U1095 ( .A1(KEYINPUT54), .A2(n1367), .ZN(n1365) );
XOR2_X1 U1096 ( .A(G107), .B(n1274), .Z(n1367) );
XOR2_X1 U1097 ( .A(G104), .B(KEYINPUT52), .Z(n1274) );
XNOR2_X1 U1098 ( .A(n1353), .B(n1294), .ZN(n1363) );
XOR2_X1 U1099 ( .A(G113), .B(KEYINPUT29), .Z(n1294) );
INV_X1 U1100 ( .A(n1354), .ZN(n1353) );
XOR2_X1 U1101 ( .A(G116), .B(n1331), .Z(n1354) );
XNOR2_X1 U1102 ( .A(G119), .B(KEYINPUT30), .ZN(n1331) );
XNOR2_X1 U1103 ( .A(G125), .B(n1368), .ZN(n1222) );
AND2_X1 U1104 ( .A1(G224), .A2(n1063), .ZN(n1368) );
INV_X1 U1105 ( .A(G953), .ZN(n1063) );
INV_X1 U1106 ( .A(G110), .ZN(n1258) );
endmodule


