//Key = 1100110100001111110011111011110010101001010000101101000100001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313;

NAND2_X1 U733 ( .A1(n1010), .A2(n1011), .ZN(G9) );
NAND2_X1 U734 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND2_X1 U735 ( .A1(G107), .A2(n1014), .ZN(n1010) );
NAND2_X1 U736 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U737 ( .A1(KEYINPUT45), .A2(n1017), .ZN(n1016) );
OR2_X1 U738 ( .A1(n1012), .A2(KEYINPUT45), .ZN(n1015) );
AND2_X1 U739 ( .A1(KEYINPUT51), .A2(n1017), .ZN(n1012) );
NAND3_X1 U740 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(G75) );
NAND2_X1 U741 ( .A1(G952), .A2(n1021), .ZN(n1020) );
NAND3_X1 U742 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1021) );
NAND2_X1 U743 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NAND2_X1 U744 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND3_X1 U745 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NAND3_X1 U746 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1030) );
INV_X1 U747 ( .A(n1035), .ZN(n1034) );
NAND2_X1 U748 ( .A1(n1036), .A2(n1037), .ZN(n1033) );
NAND2_X1 U749 ( .A1(n1038), .A2(n1039), .ZN(n1032) );
NAND3_X1 U750 ( .A1(n1037), .A2(n1040), .A3(n1039), .ZN(n1027) );
NAND3_X1 U751 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NAND2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
XNOR2_X1 U753 ( .A(KEYINPUT44), .B(n1046), .ZN(n1045) );
NAND3_X1 U754 ( .A1(n1031), .A2(n1047), .A3(n1048), .ZN(n1042) );
NAND2_X1 U755 ( .A1(n1029), .A2(n1049), .ZN(n1041) );
NAND2_X1 U756 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND3_X1 U757 ( .A1(n1052), .A2(n1053), .A3(KEYINPUT41), .ZN(n1051) );
NAND2_X1 U758 ( .A1(n1054), .A2(n1055), .ZN(n1022) );
INV_X1 U759 ( .A(KEYINPUT41), .ZN(n1055) );
NAND4_X1 U760 ( .A1(n1039), .A2(n1029), .A3(n1053), .A4(n1056), .ZN(n1054) );
AND3_X1 U761 ( .A1(n1052), .A2(n1025), .A3(n1037), .ZN(n1056) );
XNOR2_X1 U762 ( .A(n1057), .B(KEYINPUT55), .ZN(n1025) );
NAND4_X1 U763 ( .A1(n1029), .A2(n1058), .A3(n1039), .A4(n1059), .ZN(n1018) );
NOR3_X1 U764 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NOR2_X1 U765 ( .A1(KEYINPUT14), .A2(n1063), .ZN(n1062) );
NOR3_X1 U766 ( .A1(n1064), .A2(n1053), .A3(n1065), .ZN(n1063) );
AND2_X1 U767 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
AND2_X1 U768 ( .A1(n1046), .A2(KEYINPUT14), .ZN(n1061) );
XNOR2_X1 U769 ( .A(n1068), .B(n1069), .ZN(n1060) );
XNOR2_X1 U770 ( .A(KEYINPUT36), .B(n1070), .ZN(n1058) );
NAND2_X1 U771 ( .A1(n1071), .A2(n1072), .ZN(G72) );
NAND2_X1 U772 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XOR2_X1 U773 ( .A(n1075), .B(KEYINPUT11), .Z(n1071) );
OR2_X1 U774 ( .A1(n1074), .A2(n1073), .ZN(n1075) );
XNOR2_X1 U775 ( .A(n1076), .B(n1077), .ZN(n1073) );
NOR2_X1 U776 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XNOR2_X1 U777 ( .A(G953), .B(KEYINPUT16), .ZN(n1079) );
NOR2_X1 U778 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
XOR2_X1 U779 ( .A(n1082), .B(KEYINPUT19), .Z(n1080) );
NAND2_X1 U780 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U781 ( .A(KEYINPUT28), .B(n1085), .Z(n1084) );
INV_X1 U782 ( .A(n1086), .ZN(n1083) );
NAND2_X1 U783 ( .A1(n1087), .A2(n1088), .ZN(n1076) );
NAND2_X1 U784 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
INV_X1 U785 ( .A(G900), .ZN(n1090) );
XOR2_X1 U786 ( .A(n1091), .B(n1092), .Z(n1087) );
XOR2_X1 U787 ( .A(n1093), .B(n1094), .Z(n1091) );
NAND2_X1 U788 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
XOR2_X1 U789 ( .A(KEYINPUT39), .B(n1097), .Z(n1095) );
NOR2_X1 U790 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XNOR2_X1 U791 ( .A(n1100), .B(KEYINPUT18), .ZN(n1099) );
NAND2_X1 U792 ( .A1(G953), .A2(n1101), .ZN(n1074) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1101) );
XOR2_X1 U794 ( .A(n1102), .B(n1103), .Z(G69) );
NOR2_X1 U795 ( .A1(n1104), .A2(n1019), .ZN(n1103) );
AND2_X1 U796 ( .A1(G224), .A2(G898), .ZN(n1104) );
NAND2_X1 U797 ( .A1(n1105), .A2(n1106), .ZN(n1102) );
NAND3_X1 U798 ( .A1(n1107), .A2(n1019), .A3(n1108), .ZN(n1106) );
XOR2_X1 U799 ( .A(KEYINPUT0), .B(n1109), .Z(n1105) );
NOR2_X1 U800 ( .A1(n1108), .A2(n1107), .ZN(n1109) );
NAND2_X1 U801 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
XNOR2_X1 U802 ( .A(n1112), .B(n1113), .ZN(n1110) );
XOR2_X1 U803 ( .A(KEYINPUT63), .B(n1114), .Z(n1113) );
NOR2_X1 U804 ( .A1(KEYINPUT57), .A2(n1115), .ZN(n1114) );
NOR2_X1 U805 ( .A1(n1116), .A2(n1117), .ZN(G66) );
XOR2_X1 U806 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U807 ( .A(KEYINPUT13), .B(n1120), .Z(n1119) );
NOR2_X1 U808 ( .A1(n1069), .A2(n1121), .ZN(n1120) );
NOR2_X1 U809 ( .A1(n1116), .A2(n1122), .ZN(G63) );
XNOR2_X1 U810 ( .A(n1123), .B(n1124), .ZN(n1122) );
AND2_X1 U811 ( .A1(G478), .A2(n1125), .ZN(n1124) );
NOR2_X1 U812 ( .A1(n1116), .A2(n1126), .ZN(G60) );
XOR2_X1 U813 ( .A(n1127), .B(n1128), .Z(n1126) );
AND2_X1 U814 ( .A1(G475), .A2(n1125), .ZN(n1128) );
XNOR2_X1 U815 ( .A(G104), .B(n1129), .ZN(G6) );
NAND4_X1 U816 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1037), .ZN(n1129) );
NOR2_X1 U817 ( .A1(n1133), .A2(n1050), .ZN(n1132) );
INV_X1 U818 ( .A(n1134), .ZN(n1050) );
XNOR2_X1 U819 ( .A(n1135), .B(KEYINPUT5), .ZN(n1130) );
NOR2_X1 U820 ( .A1(n1116), .A2(n1136), .ZN(G57) );
XOR2_X1 U821 ( .A(n1137), .B(n1138), .Z(n1136) );
XNOR2_X1 U822 ( .A(n1139), .B(n1140), .ZN(n1138) );
NOR3_X1 U823 ( .A1(n1121), .A2(KEYINPUT58), .A3(n1141), .ZN(n1140) );
INV_X1 U824 ( .A(n1125), .ZN(n1121) );
XOR2_X1 U825 ( .A(n1142), .B(n1143), .Z(n1137) );
NOR2_X1 U826 ( .A1(n1116), .A2(n1144), .ZN(G54) );
XOR2_X1 U827 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U828 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U829 ( .A(n1149), .B(n1150), .ZN(n1148) );
NAND2_X1 U830 ( .A1(KEYINPUT26), .A2(n1151), .ZN(n1149) );
XOR2_X1 U831 ( .A(n1152), .B(n1153), .Z(n1145) );
XOR2_X1 U832 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U833 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U834 ( .A(KEYINPUT9), .B(KEYINPUT61), .Z(n1157) );
NAND3_X1 U835 ( .A1(n1158), .A2(n1159), .A3(G469), .ZN(n1154) );
OR2_X1 U836 ( .A1(n1125), .A2(KEYINPUT54), .ZN(n1159) );
NAND2_X1 U837 ( .A1(KEYINPUT54), .A2(n1160), .ZN(n1158) );
OR2_X1 U838 ( .A1(G902), .A2(n1024), .ZN(n1160) );
NAND2_X1 U839 ( .A1(KEYINPUT4), .A2(n1094), .ZN(n1152) );
NOR2_X1 U840 ( .A1(n1116), .A2(n1161), .ZN(G51) );
XOR2_X1 U841 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U842 ( .A1(KEYINPUT3), .A2(n1164), .ZN(n1163) );
XOR2_X1 U843 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U844 ( .A(n1167), .B(n1168), .Z(n1165) );
NOR2_X1 U845 ( .A1(G125), .A2(KEYINPUT35), .ZN(n1168) );
NAND2_X1 U846 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
XNOR2_X1 U847 ( .A(KEYINPUT50), .B(KEYINPUT42), .ZN(n1169) );
NAND2_X1 U848 ( .A1(n1125), .A2(G210), .ZN(n1162) );
NOR2_X1 U849 ( .A1(n1066), .A2(n1024), .ZN(n1125) );
NOR4_X1 U850 ( .A1(n1108), .A2(n1086), .A3(n1081), .A4(n1085), .ZN(n1024) );
NOR2_X1 U851 ( .A1(n1171), .A2(n1133), .ZN(n1085) );
NAND4_X1 U852 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1081) );
NAND3_X1 U853 ( .A1(n1038), .A2(n1131), .A3(n1176), .ZN(n1172) );
NAND3_X1 U854 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1086) );
NAND3_X1 U855 ( .A1(n1180), .A2(n1036), .A3(n1181), .ZN(n1179) );
NAND4_X1 U856 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1108) );
NOR4_X1 U857 ( .A1(n1186), .A2(n1187), .A3(n1017), .A4(n1188), .ZN(n1185) );
AND3_X1 U858 ( .A1(n1037), .A2(n1189), .A3(n1036), .ZN(n1017) );
OR2_X1 U859 ( .A1(n1190), .A2(n1133), .ZN(n1184) );
NAND4_X1 U860 ( .A1(n1180), .A2(n1031), .A3(n1039), .A4(n1191), .ZN(n1183) );
NAND2_X1 U861 ( .A1(n1189), .A2(n1035), .ZN(n1182) );
NAND2_X1 U862 ( .A1(n1192), .A2(n1193), .ZN(n1035) );
NAND2_X1 U863 ( .A1(n1131), .A2(n1037), .ZN(n1193) );
NAND2_X1 U864 ( .A1(n1194), .A2(n1039), .ZN(n1192) );
NOR2_X1 U865 ( .A1(n1019), .A2(G952), .ZN(n1116) );
XOR2_X1 U866 ( .A(n1173), .B(n1195), .Z(G48) );
NAND2_X1 U867 ( .A1(KEYINPUT21), .A2(G146), .ZN(n1195) );
NAND3_X1 U868 ( .A1(n1180), .A2(n1131), .A3(n1181), .ZN(n1173) );
XNOR2_X1 U869 ( .A(G143), .B(n1174), .ZN(G45) );
NAND4_X1 U870 ( .A1(n1181), .A2(n1194), .A3(n1196), .A4(n1197), .ZN(n1174) );
XNOR2_X1 U871 ( .A(G140), .B(n1198), .ZN(G42) );
NAND3_X1 U872 ( .A1(n1134), .A2(n1199), .A3(n1200), .ZN(n1198) );
XOR2_X1 U873 ( .A(KEYINPUT52), .B(n1029), .Z(n1199) );
XNOR2_X1 U874 ( .A(n1175), .B(n1201), .ZN(G39) );
XOR2_X1 U875 ( .A(KEYINPUT62), .B(G137), .Z(n1201) );
NAND3_X1 U876 ( .A1(n1180), .A2(n1039), .A3(n1176), .ZN(n1175) );
XOR2_X1 U877 ( .A(n1177), .B(n1202), .Z(G36) );
NAND2_X1 U878 ( .A1(KEYINPUT23), .A2(G134), .ZN(n1202) );
NAND3_X1 U879 ( .A1(n1194), .A2(n1036), .A3(n1176), .ZN(n1177) );
XNOR2_X1 U880 ( .A(G131), .B(n1178), .ZN(G33) );
NAND3_X1 U881 ( .A1(n1194), .A2(n1131), .A3(n1176), .ZN(n1178) );
AND3_X1 U882 ( .A1(n1029), .A2(n1134), .A3(n1203), .ZN(n1176) );
NOR2_X1 U883 ( .A1(n1204), .A2(n1048), .ZN(n1029) );
XNOR2_X1 U884 ( .A(G128), .B(n1205), .ZN(G30) );
NAND4_X1 U885 ( .A1(KEYINPUT1), .A2(n1181), .A3(n1180), .A4(n1036), .ZN(n1205) );
AND3_X1 U886 ( .A1(n1134), .A2(n1044), .A3(n1203), .ZN(n1181) );
NAND2_X1 U887 ( .A1(n1206), .A2(n1207), .ZN(G3) );
NAND2_X1 U888 ( .A1(G101), .A2(n1208), .ZN(n1207) );
XOR2_X1 U889 ( .A(KEYINPUT46), .B(n1209), .Z(n1206) );
NOR2_X1 U890 ( .A1(G101), .A2(n1208), .ZN(n1209) );
NAND3_X1 U891 ( .A1(n1039), .A2(n1189), .A3(n1194), .ZN(n1208) );
NAND2_X1 U892 ( .A1(n1210), .A2(n1211), .ZN(G27) );
NAND2_X1 U893 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XOR2_X1 U894 ( .A(KEYINPUT34), .B(n1214), .Z(n1210) );
NOR2_X1 U895 ( .A1(n1212), .A2(n1213), .ZN(n1214) );
AND2_X1 U896 ( .A1(n1215), .A2(n1044), .ZN(n1212) );
XOR2_X1 U897 ( .A(n1171), .B(KEYINPUT49), .Z(n1215) );
NAND2_X1 U898 ( .A1(n1031), .A2(n1200), .ZN(n1171) );
AND3_X1 U899 ( .A1(n1131), .A2(n1203), .A3(n1038), .ZN(n1200) );
AND4_X1 U900 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1203) );
OR3_X1 U901 ( .A1(G952), .A2(G953), .A3(KEYINPUT2), .ZN(n1219) );
NAND2_X1 U902 ( .A1(KEYINPUT2), .A2(G953), .ZN(n1218) );
NAND2_X1 U903 ( .A1(G900), .A2(n1220), .ZN(n1217) );
XOR2_X1 U904 ( .A(G122), .B(n1188), .Z(G24) );
AND4_X1 U905 ( .A1(n1031), .A2(n1037), .A3(n1221), .A4(n1191), .ZN(n1188) );
NOR2_X1 U906 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NOR2_X1 U907 ( .A1(n1224), .A2(n1225), .ZN(n1037) );
XNOR2_X1 U908 ( .A(G119), .B(n1226), .ZN(G21) );
NAND4_X1 U909 ( .A1(n1227), .A2(n1180), .A3(n1039), .A4(n1191), .ZN(n1226) );
NOR2_X1 U910 ( .A1(n1228), .A2(n1070), .ZN(n1180) );
XNOR2_X1 U911 ( .A(n1031), .B(KEYINPUT60), .ZN(n1227) );
XNOR2_X1 U912 ( .A(n1229), .B(n1230), .ZN(G18) );
NAND2_X1 U913 ( .A1(KEYINPUT17), .A2(n1231), .ZN(n1229) );
NAND2_X1 U914 ( .A1(n1232), .A2(n1044), .ZN(n1231) );
XOR2_X1 U915 ( .A(n1190), .B(KEYINPUT20), .Z(n1232) );
NAND4_X1 U916 ( .A1(n1194), .A2(n1031), .A3(n1036), .A4(n1135), .ZN(n1190) );
INV_X1 U917 ( .A(n1233), .ZN(n1135) );
NOR2_X1 U918 ( .A1(n1197), .A2(n1223), .ZN(n1036) );
INV_X1 U919 ( .A(n1196), .ZN(n1223) );
XOR2_X1 U920 ( .A(G113), .B(n1187), .Z(G15) );
AND4_X1 U921 ( .A1(n1194), .A2(n1031), .A3(n1131), .A4(n1191), .ZN(n1187) );
NOR2_X1 U922 ( .A1(n1196), .A2(n1222), .ZN(n1131) );
INV_X1 U923 ( .A(n1197), .ZN(n1222) );
INV_X1 U924 ( .A(n1046), .ZN(n1031) );
NAND2_X1 U925 ( .A1(n1052), .A2(n1234), .ZN(n1046) );
NOR2_X1 U926 ( .A1(n1225), .A2(n1070), .ZN(n1194) );
INV_X1 U927 ( .A(n1224), .ZN(n1070) );
INV_X1 U928 ( .A(n1228), .ZN(n1225) );
XOR2_X1 U929 ( .A(G110), .B(n1186), .Z(G12) );
AND3_X1 U930 ( .A1(n1039), .A2(n1189), .A3(n1038), .ZN(n1186) );
NOR2_X1 U931 ( .A1(n1228), .A2(n1224), .ZN(n1038) );
XOR2_X1 U932 ( .A(n1235), .B(n1141), .Z(n1224) );
INV_X1 U933 ( .A(G472), .ZN(n1141) );
NAND2_X1 U934 ( .A1(n1236), .A2(n1066), .ZN(n1235) );
XOR2_X1 U935 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U936 ( .A(KEYINPUT59), .B(n1239), .Z(n1238) );
NOR2_X1 U937 ( .A1(KEYINPUT56), .A2(n1139), .ZN(n1239) );
NAND2_X1 U938 ( .A1(G210), .A2(n1240), .ZN(n1139) );
XOR2_X1 U939 ( .A(n1142), .B(n1241), .Z(n1237) );
NOR2_X1 U940 ( .A1(KEYINPUT47), .A2(n1143), .ZN(n1241) );
XNOR2_X1 U941 ( .A(n1242), .B(n1243), .ZN(n1143) );
XOR2_X1 U942 ( .A(KEYINPUT43), .B(G113), .Z(n1243) );
NAND2_X1 U943 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
NAND2_X1 U944 ( .A1(G119), .A2(n1230), .ZN(n1245) );
XOR2_X1 U945 ( .A(KEYINPUT32), .B(n1246), .Z(n1244) );
NOR2_X1 U946 ( .A1(G119), .A2(n1230), .ZN(n1246) );
XOR2_X1 U947 ( .A(n1247), .B(n1248), .Z(n1142) );
XNOR2_X1 U948 ( .A(G101), .B(n1156), .ZN(n1248) );
XNOR2_X1 U949 ( .A(n1069), .B(n1249), .ZN(n1228) );
NOR2_X1 U950 ( .A1(n1068), .A2(KEYINPUT31), .ZN(n1249) );
AND2_X1 U951 ( .A1(n1250), .A2(n1118), .ZN(n1068) );
XNOR2_X1 U952 ( .A(n1251), .B(n1252), .ZN(n1118) );
XOR2_X1 U953 ( .A(n1253), .B(n1092), .Z(n1252) );
XOR2_X1 U954 ( .A(n1254), .B(n1255), .Z(n1251) );
NOR2_X1 U955 ( .A1(KEYINPUT6), .A2(n1256), .ZN(n1255) );
XOR2_X1 U956 ( .A(n1257), .B(G137), .Z(n1256) );
NAND2_X1 U957 ( .A1(G221), .A2(n1258), .ZN(n1257) );
XNOR2_X1 U958 ( .A(G110), .B(G119), .ZN(n1254) );
XNOR2_X1 U959 ( .A(G902), .B(KEYINPUT33), .ZN(n1250) );
NAND2_X1 U960 ( .A1(G217), .A2(n1259), .ZN(n1069) );
AND2_X1 U961 ( .A1(n1191), .A2(n1134), .ZN(n1189) );
NOR2_X1 U962 ( .A1(n1052), .A2(n1053), .ZN(n1134) );
INV_X1 U963 ( .A(n1234), .ZN(n1053) );
NAND2_X1 U964 ( .A1(n1260), .A2(n1259), .ZN(n1234) );
NAND2_X1 U965 ( .A1(G234), .A2(n1066), .ZN(n1259) );
XNOR2_X1 U966 ( .A(G221), .B(KEYINPUT22), .ZN(n1260) );
XNOR2_X1 U967 ( .A(n1261), .B(n1064), .ZN(n1052) );
INV_X1 U968 ( .A(G469), .ZN(n1064) );
NAND2_X1 U969 ( .A1(n1067), .A2(n1066), .ZN(n1261) );
XNOR2_X1 U970 ( .A(n1262), .B(n1263), .ZN(n1067) );
XOR2_X1 U971 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U972 ( .A(n1151), .B(n1266), .Z(n1265) );
NOR2_X1 U973 ( .A1(KEYINPUT38), .A2(n1150), .ZN(n1266) );
XNOR2_X1 U974 ( .A(G140), .B(G110), .ZN(n1150) );
NAND2_X1 U975 ( .A1(G227), .A2(n1019), .ZN(n1151) );
NAND2_X1 U976 ( .A1(KEYINPUT15), .A2(n1094), .ZN(n1264) );
XNOR2_X1 U977 ( .A(n1267), .B(KEYINPUT10), .ZN(n1094) );
XNOR2_X1 U978 ( .A(n1147), .B(n1156), .ZN(n1262) );
NAND3_X1 U979 ( .A1(n1268), .A2(n1269), .A3(n1096), .ZN(n1156) );
NAND2_X1 U980 ( .A1(n1270), .A2(n1098), .ZN(n1096) );
INV_X1 U981 ( .A(n1271), .ZN(n1098) );
INV_X1 U982 ( .A(n1100), .ZN(n1270) );
OR2_X1 U983 ( .A1(n1100), .A2(KEYINPUT7), .ZN(n1269) );
NAND3_X1 U984 ( .A1(n1271), .A2(n1100), .A3(KEYINPUT7), .ZN(n1268) );
XOR2_X1 U985 ( .A(G131), .B(KEYINPUT8), .Z(n1100) );
XOR2_X1 U986 ( .A(G134), .B(G137), .Z(n1271) );
XOR2_X1 U987 ( .A(n1272), .B(KEYINPUT53), .Z(n1147) );
NOR2_X1 U988 ( .A1(n1133), .A2(n1233), .ZN(n1191) );
NAND2_X1 U989 ( .A1(n1216), .A2(n1273), .ZN(n1233) );
NAND2_X1 U990 ( .A1(n1220), .A2(n1111), .ZN(n1273) );
NAND2_X1 U991 ( .A1(n1089), .A2(n1274), .ZN(n1111) );
XOR2_X1 U992 ( .A(KEYINPUT12), .B(G898), .Z(n1274) );
XNOR2_X1 U993 ( .A(KEYINPUT2), .B(n1019), .ZN(n1089) );
AND2_X1 U994 ( .A1(n1057), .A2(n1275), .ZN(n1216) );
NAND2_X1 U995 ( .A1(n1220), .A2(n1066), .ZN(n1275) );
NAND2_X1 U996 ( .A1(G952), .A2(n1019), .ZN(n1220) );
NAND2_X1 U997 ( .A1(G237), .A2(G234), .ZN(n1057) );
INV_X1 U998 ( .A(n1044), .ZN(n1133) );
NOR2_X1 U999 ( .A1(n1047), .A2(n1048), .ZN(n1044) );
AND2_X1 U1000 ( .A1(G214), .A2(n1276), .ZN(n1048) );
OR2_X1 U1001 ( .A1(G902), .A2(G237), .ZN(n1276) );
INV_X1 U1002 ( .A(n1204), .ZN(n1047) );
NAND3_X1 U1003 ( .A1(n1277), .A2(n1278), .A3(n1279), .ZN(n1204) );
OR2_X1 U1004 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND3_X1 U1005 ( .A1(n1281), .A2(n1280), .A3(n1066), .ZN(n1278) );
NAND2_X1 U1006 ( .A1(G237), .A2(G210), .ZN(n1280) );
XNOR2_X1 U1007 ( .A(n1282), .B(n1166), .ZN(n1281) );
XNOR2_X1 U1008 ( .A(n1247), .B(n1283), .ZN(n1166) );
AND2_X1 U1009 ( .A1(n1019), .A2(G224), .ZN(n1283) );
XOR2_X1 U1010 ( .A(n1267), .B(KEYINPUT29), .Z(n1247) );
XNOR2_X1 U1011 ( .A(G143), .B(n1253), .ZN(n1267) );
XOR2_X1 U1012 ( .A(G128), .B(G146), .Z(n1253) );
XNOR2_X1 U1013 ( .A(n1170), .B(n1213), .ZN(n1282) );
NAND2_X1 U1014 ( .A1(n1284), .A2(n1285), .ZN(n1170) );
NAND2_X1 U1015 ( .A1(n1115), .A2(n1112), .ZN(n1285) );
XOR2_X1 U1016 ( .A(n1286), .B(KEYINPUT37), .Z(n1284) );
OR2_X1 U1017 ( .A1(n1112), .A2(n1115), .ZN(n1286) );
XOR2_X1 U1018 ( .A(G110), .B(n1287), .Z(n1115) );
XOR2_X1 U1019 ( .A(KEYINPUT40), .B(G122), .Z(n1287) );
XNOR2_X1 U1020 ( .A(n1288), .B(n1289), .ZN(n1112) );
XNOR2_X1 U1021 ( .A(n1230), .B(G113), .ZN(n1289) );
INV_X1 U1022 ( .A(G116), .ZN(n1230) );
XOR2_X1 U1023 ( .A(n1272), .B(n1290), .Z(n1288) );
NOR2_X1 U1024 ( .A1(G119), .A2(KEYINPUT30), .ZN(n1290) );
XNOR2_X1 U1025 ( .A(G101), .B(n1291), .ZN(n1272) );
XNOR2_X1 U1026 ( .A(n1013), .B(G104), .ZN(n1291) );
INV_X1 U1027 ( .A(G107), .ZN(n1013) );
NAND2_X1 U1028 ( .A1(G902), .A2(G210), .ZN(n1277) );
NOR2_X1 U1029 ( .A1(n1196), .A2(n1197), .ZN(n1039) );
XOR2_X1 U1030 ( .A(G475), .B(n1292), .Z(n1197) );
NOR2_X1 U1031 ( .A1(n1127), .A2(G902), .ZN(n1292) );
AND2_X1 U1032 ( .A1(n1293), .A2(n1294), .ZN(n1127) );
NAND2_X1 U1033 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
XOR2_X1 U1034 ( .A(KEYINPUT24), .B(n1297), .Z(n1293) );
NOR2_X1 U1035 ( .A1(n1295), .A2(n1296), .ZN(n1297) );
XOR2_X1 U1036 ( .A(G104), .B(n1298), .Z(n1296) );
XOR2_X1 U1037 ( .A(G122), .B(G113), .Z(n1298) );
XNOR2_X1 U1038 ( .A(n1299), .B(n1300), .ZN(n1295) );
XNOR2_X1 U1039 ( .A(n1301), .B(n1302), .ZN(n1300) );
XOR2_X1 U1040 ( .A(KEYINPUT27), .B(G146), .Z(n1302) );
XOR2_X1 U1041 ( .A(n1303), .B(n1092), .Z(n1299) );
XNOR2_X1 U1042 ( .A(G140), .B(n1213), .ZN(n1092) );
INV_X1 U1043 ( .A(G125), .ZN(n1213) );
XOR2_X1 U1044 ( .A(n1304), .B(G131), .Z(n1303) );
NAND2_X1 U1045 ( .A1(G214), .A2(n1240), .ZN(n1304) );
NOR2_X1 U1046 ( .A1(G953), .A2(G237), .ZN(n1240) );
XNOR2_X1 U1047 ( .A(n1305), .B(G478), .ZN(n1196) );
NAND2_X1 U1048 ( .A1(n1123), .A2(n1066), .ZN(n1305) );
INV_X1 U1049 ( .A(G902), .ZN(n1066) );
XNOR2_X1 U1050 ( .A(n1306), .B(n1307), .ZN(n1123) );
AND2_X1 U1051 ( .A1(n1258), .A2(G217), .ZN(n1307) );
AND2_X1 U1052 ( .A1(G234), .A2(n1019), .ZN(n1258) );
INV_X1 U1053 ( .A(G953), .ZN(n1019) );
NAND2_X1 U1054 ( .A1(n1308), .A2(KEYINPUT48), .ZN(n1306) );
XOR2_X1 U1055 ( .A(n1309), .B(n1310), .Z(n1308) );
XOR2_X1 U1056 ( .A(G128), .B(n1311), .Z(n1310) );
XNOR2_X1 U1057 ( .A(n1301), .B(G134), .ZN(n1311) );
INV_X1 U1058 ( .A(G143), .ZN(n1301) );
XOR2_X1 U1059 ( .A(n1312), .B(n1313), .Z(n1309) );
NOR2_X1 U1060 ( .A1(KEYINPUT25), .A2(G107), .ZN(n1313) );
XNOR2_X1 U1061 ( .A(G116), .B(G122), .ZN(n1312) );
endmodule


