//Key = 1011111000011011001101101111011001100110101101001101001000001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353;

XOR2_X1 U734 ( .A(G107), .B(n1021), .Z(G9) );
NAND3_X1 U735 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(G75) );
NAND2_X1 U736 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NAND2_X1 U737 ( .A1(G952), .A2(n1027), .ZN(n1022) );
NAND4_X1 U738 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1027) );
NAND2_X1 U739 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NAND2_X1 U740 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND3_X1 U741 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NAND2_X1 U742 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NAND2_X1 U743 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
OR2_X1 U744 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U745 ( .A1(n1045), .A2(n1046), .ZN(n1039) );
NAND3_X1 U746 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
OR3_X1 U747 ( .A1(n1050), .A2(n1051), .A3(KEYINPUT57), .ZN(n1048) );
NAND2_X1 U748 ( .A1(KEYINPUT57), .A2(n1041), .ZN(n1047) );
NAND3_X1 U749 ( .A1(n1052), .A2(n1053), .A3(n1041), .ZN(n1034) );
NAND2_X1 U750 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U751 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
INV_X1 U752 ( .A(KEYINPUT30), .ZN(n1057) );
NAND4_X1 U753 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1045), .ZN(n1052) );
NAND2_X1 U754 ( .A1(KEYINPUT30), .A2(n1056), .ZN(n1060) );
NAND3_X1 U755 ( .A1(n1061), .A2(n1036), .A3(n1062), .ZN(n1059) );
NAND2_X1 U756 ( .A1(n1038), .A2(n1063), .ZN(n1058) );
NAND2_X1 U757 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
INV_X1 U758 ( .A(n1066), .ZN(n1032) );
XOR2_X1 U759 ( .A(KEYINPUT38), .B(n1025), .Z(n1029) );
AND4_X1 U760 ( .A1(n1061), .A2(n1045), .A3(n1067), .A4(n1068), .ZN(n1025) );
NOR4_X1 U761 ( .A1(n1069), .A2(n1062), .A3(n1070), .A4(n1071), .ZN(n1068) );
XOR2_X1 U762 ( .A(n1072), .B(KEYINPUT59), .Z(n1070) );
NAND2_X1 U763 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XNOR2_X1 U764 ( .A(KEYINPUT25), .B(n1075), .ZN(n1073) );
XOR2_X1 U765 ( .A(n1076), .B(KEYINPUT28), .Z(n1067) );
NAND2_X1 U766 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U767 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U768 ( .A(n1081), .B(n1082), .Z(G72) );
NOR2_X1 U769 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U770 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U771 ( .A1(n1087), .A2(n1088), .ZN(n1083) );
XOR2_X1 U772 ( .A(n1089), .B(KEYINPUT1), .Z(n1088) );
NAND2_X1 U773 ( .A1(n1031), .A2(n1085), .ZN(n1089) );
INV_X1 U774 ( .A(n1086), .ZN(n1087) );
NAND2_X1 U775 ( .A1(n1090), .A2(n1091), .ZN(n1086) );
NAND2_X1 U776 ( .A1(G953), .A2(n1092), .ZN(n1091) );
XOR2_X1 U777 ( .A(n1093), .B(n1094), .Z(n1090) );
XOR2_X1 U778 ( .A(n1095), .B(n1096), .Z(n1093) );
NAND2_X1 U779 ( .A1(G953), .A2(n1097), .ZN(n1081) );
NAND2_X1 U780 ( .A1(G900), .A2(G227), .ZN(n1097) );
NAND2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(G69) );
NAND3_X1 U782 ( .A1(G953), .A2(n1100), .A3(n1101), .ZN(n1099) );
XOR2_X1 U783 ( .A(KEYINPUT14), .B(n1102), .Z(n1098) );
NOR2_X1 U784 ( .A1(n1101), .A2(n1103), .ZN(n1102) );
AND2_X1 U785 ( .A1(n1100), .A2(G953), .ZN(n1103) );
NAND2_X1 U786 ( .A1(G898), .A2(G224), .ZN(n1100) );
AND2_X1 U787 ( .A1(n1104), .A2(n1105), .ZN(n1101) );
NAND3_X1 U788 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
NAND2_X1 U789 ( .A1(n1109), .A2(n1110), .ZN(n1104) );
NAND2_X1 U790 ( .A1(n1108), .A2(n1107), .ZN(n1110) );
XOR2_X1 U791 ( .A(KEYINPUT63), .B(n1031), .Z(n1108) );
XOR2_X1 U792 ( .A(n1106), .B(KEYINPUT0), .Z(n1109) );
NAND2_X1 U793 ( .A1(n1111), .A2(n1112), .ZN(n1106) );
NAND2_X1 U794 ( .A1(G953), .A2(n1113), .ZN(n1112) );
XOR2_X1 U795 ( .A(n1114), .B(n1115), .Z(n1111) );
NOR2_X1 U796 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NOR2_X1 U797 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XNOR2_X1 U798 ( .A(n1120), .B(n1121), .ZN(n1119) );
NAND2_X1 U799 ( .A1(n1122), .A2(G217), .ZN(n1120) );
NOR2_X1 U800 ( .A1(n1118), .A2(n1123), .ZN(G63) );
XOR2_X1 U801 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U802 ( .A1(n1080), .A2(n1126), .ZN(n1125) );
NAND2_X1 U803 ( .A1(KEYINPUT48), .A2(n1127), .ZN(n1124) );
NOR2_X1 U804 ( .A1(n1118), .A2(n1128), .ZN(G60) );
XOR2_X1 U805 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U806 ( .A1(n1122), .A2(G475), .ZN(n1129) );
XOR2_X1 U807 ( .A(G104), .B(n1131), .Z(G6) );
NOR2_X1 U808 ( .A1(n1118), .A2(n1132), .ZN(G57) );
XOR2_X1 U809 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U810 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U811 ( .A(n1137), .B(KEYINPUT40), .Z(n1136) );
NAND3_X1 U812 ( .A1(G472), .A2(n1138), .A3(n1122), .ZN(n1137) );
NOR2_X1 U813 ( .A1(n1139), .A2(n1138), .ZN(n1135) );
XNOR2_X1 U814 ( .A(n1140), .B(n1096), .ZN(n1138) );
AND2_X1 U815 ( .A1(G472), .A2(n1122), .ZN(n1139) );
NOR2_X1 U816 ( .A1(n1118), .A2(n1141), .ZN(G54) );
XOR2_X1 U817 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U818 ( .A(n1144), .B(n1145), .Z(n1143) );
NAND2_X1 U819 ( .A1(KEYINPUT4), .A2(n1146), .ZN(n1144) );
XOR2_X1 U820 ( .A(KEYINPUT3), .B(n1147), .Z(n1146) );
XOR2_X1 U821 ( .A(n1148), .B(n1149), .Z(n1142) );
NOR3_X1 U822 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1149) );
NOR2_X1 U823 ( .A1(KEYINPUT51), .A2(n1153), .ZN(n1152) );
NOR2_X1 U824 ( .A1(n1028), .A2(G902), .ZN(n1153) );
AND2_X1 U825 ( .A1(n1126), .A2(KEYINPUT51), .ZN(n1151) );
INV_X1 U826 ( .A(n1122), .ZN(n1126) );
NOR2_X1 U827 ( .A1(KEYINPUT7), .A2(n1154), .ZN(n1148) );
XNOR2_X1 U828 ( .A(n1155), .B(KEYINPUT23), .ZN(n1154) );
NOR2_X1 U829 ( .A1(n1118), .A2(n1156), .ZN(G51) );
XOR2_X1 U830 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U831 ( .A(n1159), .B(n1160), .ZN(n1158) );
XOR2_X1 U832 ( .A(n1161), .B(n1155), .Z(n1160) );
NAND2_X1 U833 ( .A1(KEYINPUT29), .A2(n1162), .ZN(n1161) );
XOR2_X1 U834 ( .A(n1163), .B(n1164), .Z(n1157) );
XOR2_X1 U835 ( .A(KEYINPUT61), .B(G125), .Z(n1164) );
XOR2_X1 U836 ( .A(n1165), .B(n1166), .Z(n1163) );
NAND2_X1 U837 ( .A1(n1122), .A2(n1167), .ZN(n1165) );
NOR2_X1 U838 ( .A1(n1168), .A2(n1028), .ZN(n1122) );
NOR2_X1 U839 ( .A1(n1085), .A2(n1107), .ZN(n1028) );
NAND4_X1 U840 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1107) );
NOR4_X1 U841 ( .A1(n1021), .A2(n1173), .A3(n1174), .A4(n1131), .ZN(n1172) );
AND2_X1 U842 ( .A1(n1175), .A2(n1176), .ZN(n1131) );
AND2_X1 U843 ( .A1(n1177), .A2(n1176), .ZN(n1021) );
AND3_X1 U844 ( .A1(n1045), .A2(n1178), .A3(n1179), .ZN(n1176) );
NAND2_X1 U845 ( .A1(KEYINPUT12), .A2(n1180), .ZN(n1171) );
NAND4_X1 U846 ( .A1(n1056), .A2(n1043), .A3(n1181), .A4(n1182), .ZN(n1170) );
OR2_X1 U847 ( .A1(n1183), .A2(n1179), .ZN(n1182) );
NAND2_X1 U848 ( .A1(n1184), .A2(n1183), .ZN(n1181) );
INV_X1 U849 ( .A(KEYINPUT21), .ZN(n1183) );
NAND2_X1 U850 ( .A1(n1185), .A2(n1049), .ZN(n1184) );
NAND2_X1 U851 ( .A1(n1186), .A2(n1187), .ZN(n1169) );
NAND3_X1 U852 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
XOR2_X1 U853 ( .A(n1191), .B(KEYINPUT8), .Z(n1190) );
NAND4_X1 U854 ( .A1(n1038), .A2(n1036), .A3(n1192), .A4(n1193), .ZN(n1189) );
NOR3_X1 U855 ( .A1(n1194), .A2(KEYINPUT12), .A3(n1195), .ZN(n1193) );
XNOR2_X1 U856 ( .A(KEYINPUT42), .B(n1196), .ZN(n1188) );
NAND4_X1 U857 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1085) );
NOR3_X1 U858 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
INV_X1 U859 ( .A(n1204), .ZN(n1202) );
NOR2_X1 U860 ( .A1(n1205), .A2(n1049), .ZN(n1201) );
NOR3_X1 U861 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1205) );
NOR3_X1 U862 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1208) );
NOR2_X1 U863 ( .A1(n1065), .A2(n1212), .ZN(n1206) );
INV_X1 U864 ( .A(n1024), .ZN(n1118) );
NAND2_X1 U865 ( .A1(G953), .A2(n1026), .ZN(n1024) );
INV_X1 U866 ( .A(G952), .ZN(n1026) );
NAND3_X1 U867 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(G48) );
NAND2_X1 U868 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U869 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
XOR2_X1 U870 ( .A(n1220), .B(KEYINPUT31), .Z(n1218) );
NAND3_X1 U871 ( .A1(G146), .A2(n1220), .A3(n1219), .ZN(n1214) );
INV_X1 U872 ( .A(KEYINPUT50), .ZN(n1219) );
NAND2_X1 U873 ( .A1(n1203), .A2(KEYINPUT50), .ZN(n1213) );
INV_X1 U874 ( .A(n1220), .ZN(n1203) );
NAND3_X1 U875 ( .A1(n1175), .A2(n1186), .A3(n1221), .ZN(n1220) );
XNOR2_X1 U876 ( .A(G143), .B(n1222), .ZN(G45) );
NAND4_X1 U877 ( .A1(n1223), .A2(n1224), .A3(n1071), .A4(n1225), .ZN(n1222) );
XOR2_X1 U878 ( .A(KEYINPUT20), .B(n1186), .Z(n1224) );
XOR2_X1 U879 ( .A(n1226), .B(n1204), .Z(G42) );
NAND3_X1 U880 ( .A1(n1041), .A2(n1178), .A3(n1227), .ZN(n1204) );
XOR2_X1 U881 ( .A(n1228), .B(n1199), .Z(G39) );
NAND3_X1 U882 ( .A1(n1221), .A2(n1041), .A3(n1036), .ZN(n1199) );
XNOR2_X1 U883 ( .A(G134), .B(n1197), .ZN(G36) );
NAND3_X1 U884 ( .A1(n1041), .A2(n1177), .A3(n1223), .ZN(n1197) );
XNOR2_X1 U885 ( .A(G131), .B(n1198), .ZN(G33) );
NAND3_X1 U886 ( .A1(n1223), .A2(n1041), .A3(n1175), .ZN(n1198) );
NOR2_X1 U887 ( .A1(n1051), .A2(n1069), .ZN(n1041) );
INV_X1 U888 ( .A(n1050), .ZN(n1069) );
INV_X1 U889 ( .A(n1209), .ZN(n1223) );
NAND3_X1 U890 ( .A1(n1178), .A2(n1229), .A3(n1044), .ZN(n1209) );
NAND2_X1 U891 ( .A1(n1230), .A2(n1231), .ZN(G30) );
NAND2_X1 U892 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
XOR2_X1 U893 ( .A(n1234), .B(KEYINPUT17), .Z(n1230) );
OR2_X1 U894 ( .A1(n1233), .A2(n1232), .ZN(n1234) );
XNOR2_X1 U895 ( .A(G128), .B(KEYINPUT18), .ZN(n1232) );
NAND3_X1 U896 ( .A1(n1221), .A2(n1177), .A3(n1235), .ZN(n1233) );
XOR2_X1 U897 ( .A(n1049), .B(KEYINPUT6), .Z(n1235) );
INV_X1 U898 ( .A(n1212), .ZN(n1221) );
NAND4_X1 U899 ( .A1(n1178), .A2(n1236), .A3(n1229), .A4(n1237), .ZN(n1212) );
XOR2_X1 U900 ( .A(G101), .B(n1238), .Z(G3) );
NOR2_X1 U901 ( .A1(n1049), .A2(n1196), .ZN(n1238) );
NAND3_X1 U902 ( .A1(n1044), .A2(n1185), .A3(n1056), .ZN(n1196) );
XOR2_X1 U903 ( .A(n1239), .B(n1240), .Z(G27) );
NAND2_X1 U904 ( .A1(n1241), .A2(n1186), .ZN(n1240) );
INV_X1 U905 ( .A(n1049), .ZN(n1186) );
XNOR2_X1 U906 ( .A(n1207), .B(KEYINPUT22), .ZN(n1241) );
AND2_X1 U907 ( .A1(n1038), .A2(n1227), .ZN(n1207) );
AND3_X1 U908 ( .A1(n1175), .A2(n1229), .A3(n1043), .ZN(n1227) );
NAND2_X1 U909 ( .A1(n1066), .A2(n1242), .ZN(n1229) );
NAND4_X1 U910 ( .A1(G902), .A2(G953), .A3(n1243), .A4(n1092), .ZN(n1242) );
INV_X1 U911 ( .A(G900), .ZN(n1092) );
NAND3_X1 U912 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(G24) );
NAND2_X1 U913 ( .A1(G122), .A2(n1247), .ZN(n1246) );
NAND2_X1 U914 ( .A1(n1248), .A2(n1249), .ZN(n1245) );
INV_X1 U915 ( .A(KEYINPUT45), .ZN(n1249) );
NAND2_X1 U916 ( .A1(n1250), .A2(n1174), .ZN(n1248) );
INV_X1 U917 ( .A(n1247), .ZN(n1174) );
XNOR2_X1 U918 ( .A(KEYINPUT32), .B(G122), .ZN(n1250) );
NAND2_X1 U919 ( .A1(KEYINPUT45), .A2(n1251), .ZN(n1244) );
NAND2_X1 U920 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
OR3_X1 U921 ( .A1(n1247), .A2(G122), .A3(KEYINPUT32), .ZN(n1253) );
NAND4_X1 U922 ( .A1(n1254), .A2(n1045), .A3(n1071), .A4(n1225), .ZN(n1247) );
INV_X1 U923 ( .A(n1055), .ZN(n1045) );
NAND2_X1 U924 ( .A1(n1195), .A2(n1194), .ZN(n1055) );
NAND2_X1 U925 ( .A1(KEYINPUT32), .A2(G122), .ZN(n1252) );
NAND2_X1 U926 ( .A1(n1255), .A2(n1256), .ZN(G21) );
NAND2_X1 U927 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XNOR2_X1 U928 ( .A(n1180), .B(KEYINPUT54), .ZN(n1257) );
NAND2_X1 U929 ( .A1(G119), .A2(n1259), .ZN(n1255) );
XNOR2_X1 U930 ( .A(n1180), .B(KEYINPUT53), .ZN(n1259) );
AND4_X1 U931 ( .A1(n1254), .A2(n1036), .A3(n1236), .A4(n1237), .ZN(n1180) );
XOR2_X1 U932 ( .A(G116), .B(n1173), .Z(G18) );
AND3_X1 U933 ( .A1(n1044), .A2(n1177), .A3(n1254), .ZN(n1173) );
AND2_X1 U934 ( .A1(n1038), .A2(n1179), .ZN(n1254) );
INV_X1 U935 ( .A(n1065), .ZN(n1177) );
NAND2_X1 U936 ( .A1(n1211), .A2(n1225), .ZN(n1065) );
XOR2_X1 U937 ( .A(G113), .B(n1260), .Z(G15) );
NOR2_X1 U938 ( .A1(n1049), .A2(n1191), .ZN(n1260) );
NAND4_X1 U939 ( .A1(n1038), .A2(n1175), .A3(n1044), .A4(n1185), .ZN(n1191) );
NOR2_X1 U940 ( .A1(n1237), .A2(n1194), .ZN(n1044) );
INV_X1 U941 ( .A(n1064), .ZN(n1175) );
NAND2_X1 U942 ( .A1(n1210), .A2(n1071), .ZN(n1064) );
INV_X1 U943 ( .A(n1225), .ZN(n1210) );
AND2_X1 U944 ( .A1(n1261), .A2(n1262), .ZN(n1038) );
XNOR2_X1 U945 ( .A(KEYINPUT2), .B(n1061), .ZN(n1261) );
XOR2_X1 U946 ( .A(n1263), .B(n1264), .Z(G12) );
NAND3_X1 U947 ( .A1(n1043), .A2(n1179), .A3(n1056), .ZN(n1264) );
AND2_X1 U948 ( .A1(n1036), .A2(n1178), .ZN(n1056) );
NOR2_X1 U949 ( .A1(n1061), .A2(n1062), .ZN(n1178) );
INV_X1 U950 ( .A(n1262), .ZN(n1062) );
NAND2_X1 U951 ( .A1(G221), .A2(n1265), .ZN(n1262) );
NAND2_X1 U952 ( .A1(G234), .A2(n1168), .ZN(n1265) );
XNOR2_X1 U953 ( .A(n1266), .B(n1150), .ZN(n1061) );
INV_X1 U954 ( .A(G469), .ZN(n1150) );
NAND2_X1 U955 ( .A1(n1267), .A2(n1168), .ZN(n1266) );
XOR2_X1 U956 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U957 ( .A(KEYINPUT24), .B(n1270), .Z(n1269) );
XNOR2_X1 U958 ( .A(n1147), .B(n1155), .ZN(n1268) );
XNOR2_X1 U959 ( .A(n1271), .B(n1096), .ZN(n1155) );
XNOR2_X1 U960 ( .A(n1272), .B(n1273), .ZN(n1147) );
XOR2_X1 U961 ( .A(G140), .B(G110), .Z(n1273) );
NAND2_X1 U962 ( .A1(G227), .A2(n1031), .ZN(n1272) );
NOR2_X1 U963 ( .A1(n1225), .A2(n1071), .ZN(n1036) );
INV_X1 U964 ( .A(n1211), .ZN(n1071) );
XOR2_X1 U965 ( .A(n1274), .B(G475), .Z(n1211) );
NAND2_X1 U966 ( .A1(n1130), .A2(n1168), .ZN(n1274) );
XOR2_X1 U967 ( .A(n1275), .B(n1276), .Z(n1130) );
XOR2_X1 U968 ( .A(G104), .B(n1277), .Z(n1276) );
NOR2_X1 U969 ( .A1(KEYINPUT39), .A2(n1278), .ZN(n1277) );
XOR2_X1 U970 ( .A(n1279), .B(n1280), .Z(n1278) );
XNOR2_X1 U971 ( .A(n1281), .B(n1094), .ZN(n1280) );
XOR2_X1 U972 ( .A(n1239), .B(n1226), .Z(n1094) );
INV_X1 U973 ( .A(G140), .ZN(n1226) );
NAND2_X1 U974 ( .A1(G214), .A2(n1282), .ZN(n1281) );
XOR2_X1 U975 ( .A(n1283), .B(n1284), .Z(n1279) );
XOR2_X1 U976 ( .A(G146), .B(G131), .Z(n1284) );
NAND2_X1 U977 ( .A1(KEYINPUT11), .A2(n1285), .ZN(n1283) );
NAND2_X1 U978 ( .A1(KEYINPUT34), .A2(n1286), .ZN(n1275) );
XOR2_X1 U979 ( .A(G122), .B(G113), .Z(n1286) );
NAND3_X1 U980 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n1225) );
XOR2_X1 U981 ( .A(n1290), .B(KEYINPUT19), .Z(n1289) );
NAND2_X1 U982 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
OR2_X1 U983 ( .A1(n1077), .A2(KEYINPUT27), .ZN(n1292) );
NAND3_X1 U984 ( .A1(n1293), .A2(n1080), .A3(KEYINPUT27), .ZN(n1291) );
OR3_X1 U985 ( .A1(n1080), .A2(n1293), .A3(KEYINPUT13), .ZN(n1288) );
INV_X1 U986 ( .A(G478), .ZN(n1080) );
NAND2_X1 U987 ( .A1(KEYINPUT13), .A2(n1294), .ZN(n1287) );
INV_X1 U988 ( .A(n1077), .ZN(n1294) );
NAND2_X1 U989 ( .A1(G478), .A2(n1293), .ZN(n1077) );
INV_X1 U990 ( .A(n1079), .ZN(n1293) );
NAND2_X1 U991 ( .A1(n1127), .A2(n1168), .ZN(n1079) );
XOR2_X1 U992 ( .A(n1295), .B(n1296), .Z(n1127) );
XOR2_X1 U993 ( .A(G107), .B(n1297), .Z(n1296) );
XOR2_X1 U994 ( .A(G122), .B(G116), .Z(n1297) );
XNOR2_X1 U995 ( .A(n1298), .B(n1299), .ZN(n1295) );
NOR2_X1 U996 ( .A1(KEYINPUT9), .A2(n1300), .ZN(n1299) );
XOR2_X1 U997 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U998 ( .A(G134), .B(G128), .Z(n1302) );
INV_X1 U999 ( .A(n1285), .ZN(n1301) );
NOR4_X1 U1000 ( .A1(KEYINPUT52), .A2(n1303), .A3(n1304), .A4(n1305), .ZN(n1298) );
XOR2_X1 U1001 ( .A(KEYINPUT55), .B(G953), .Z(n1305) );
INV_X1 U1002 ( .A(G234), .ZN(n1304) );
NOR2_X1 U1003 ( .A1(n1049), .A2(n1192), .ZN(n1179) );
INV_X1 U1004 ( .A(n1185), .ZN(n1192) );
NAND2_X1 U1005 ( .A1(n1066), .A2(n1306), .ZN(n1185) );
NAND4_X1 U1006 ( .A1(G902), .A2(G953), .A3(n1243), .A4(n1113), .ZN(n1306) );
INV_X1 U1007 ( .A(G898), .ZN(n1113) );
NAND3_X1 U1008 ( .A1(n1243), .A2(n1031), .A3(G952), .ZN(n1066) );
NAND2_X1 U1009 ( .A1(G237), .A2(G234), .ZN(n1243) );
NAND2_X1 U1010 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U1011 ( .A1(n1075), .A2(n1074), .ZN(n1051) );
NAND2_X1 U1012 ( .A1(n1167), .A2(n1307), .ZN(n1074) );
NAND2_X1 U1013 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
INV_X1 U1014 ( .A(n1310), .ZN(n1167) );
NAND3_X1 U1015 ( .A1(n1309), .A2(n1310), .A3(n1308), .ZN(n1075) );
XOR2_X1 U1016 ( .A(KEYINPUT60), .B(G902), .Z(n1308) );
NAND2_X1 U1017 ( .A1(G210), .A2(n1311), .ZN(n1310) );
XNOR2_X1 U1018 ( .A(n1312), .B(n1313), .ZN(n1309) );
XOR2_X1 U1019 ( .A(n1115), .B(n1314), .Z(n1313) );
XNOR2_X1 U1020 ( .A(n1162), .B(n1096), .ZN(n1314) );
NAND2_X1 U1021 ( .A1(G224), .A2(n1031), .ZN(n1162) );
XNOR2_X1 U1022 ( .A(n1271), .B(n1159), .ZN(n1115) );
XOR2_X1 U1023 ( .A(G122), .B(n1315), .Z(n1159) );
NOR2_X1 U1024 ( .A1(KEYINPUT58), .A2(n1263), .ZN(n1315) );
XOR2_X1 U1025 ( .A(n1316), .B(n1317), .Z(n1271) );
XOR2_X1 U1026 ( .A(G107), .B(G104), .Z(n1317) );
INV_X1 U1027 ( .A(G101), .ZN(n1316) );
XOR2_X1 U1028 ( .A(n1318), .B(n1319), .Z(n1312) );
XOR2_X1 U1029 ( .A(KEYINPUT44), .B(n1166), .Z(n1319) );
NOR3_X1 U1030 ( .A1(KEYINPUT16), .A2(n1117), .A3(n1116), .ZN(n1166) );
AND2_X1 U1031 ( .A1(n1320), .A2(n1321), .ZN(n1116) );
XOR2_X1 U1032 ( .A(n1322), .B(KEYINPUT49), .Z(n1321) );
XNOR2_X1 U1033 ( .A(KEYINPUT47), .B(G113), .ZN(n1320) );
AND2_X1 U1034 ( .A1(n1323), .A2(n1324), .ZN(n1117) );
XOR2_X1 U1035 ( .A(KEYINPUT47), .B(G113), .Z(n1324) );
XOR2_X1 U1036 ( .A(n1322), .B(KEYINPUT36), .Z(n1323) );
XOR2_X1 U1037 ( .A(G116), .B(n1258), .Z(n1322) );
NAND2_X1 U1038 ( .A1(KEYINPUT33), .A2(n1239), .ZN(n1318) );
INV_X1 U1039 ( .A(G125), .ZN(n1239) );
NAND2_X1 U1040 ( .A1(G214), .A2(n1311), .ZN(n1050) );
NAND2_X1 U1041 ( .A1(n1325), .A2(n1168), .ZN(n1311) );
INV_X1 U1042 ( .A(G237), .ZN(n1325) );
NOR2_X1 U1043 ( .A1(n1236), .A2(n1195), .ZN(n1043) );
INV_X1 U1044 ( .A(n1237), .ZN(n1195) );
NAND3_X1 U1045 ( .A1(n1326), .A2(n1327), .A3(n1328), .ZN(n1237) );
NAND2_X1 U1046 ( .A1(n1329), .A2(n1121), .ZN(n1328) );
OR3_X1 U1047 ( .A1(n1121), .A2(n1329), .A3(G902), .ZN(n1327) );
NOR2_X1 U1048 ( .A1(n1303), .A2(G234), .ZN(n1329) );
INV_X1 U1049 ( .A(G217), .ZN(n1303) );
XNOR2_X1 U1050 ( .A(n1330), .B(n1331), .ZN(n1121) );
XOR2_X1 U1051 ( .A(n1332), .B(n1333), .Z(n1331) );
XOR2_X1 U1052 ( .A(G119), .B(G110), .Z(n1333) );
XOR2_X1 U1053 ( .A(KEYINPUT62), .B(G125), .Z(n1332) );
XOR2_X1 U1054 ( .A(n1334), .B(n1335), .Z(n1330) );
XOR2_X1 U1055 ( .A(n1336), .B(n1337), .Z(n1335) );
NAND2_X1 U1056 ( .A1(KEYINPUT43), .A2(G140), .ZN(n1336) );
XOR2_X1 U1057 ( .A(n1338), .B(n1339), .Z(n1334) );
AND3_X1 U1058 ( .A1(G221), .A2(n1031), .A3(G234), .ZN(n1339) );
INV_X1 U1059 ( .A(G953), .ZN(n1031) );
NAND2_X1 U1060 ( .A1(KEYINPUT5), .A2(n1228), .ZN(n1338) );
INV_X1 U1061 ( .A(G137), .ZN(n1228) );
NAND2_X1 U1062 ( .A1(G902), .A2(G217), .ZN(n1326) );
INV_X1 U1063 ( .A(n1194), .ZN(n1236) );
XOR2_X1 U1064 ( .A(n1340), .B(G472), .Z(n1194) );
NAND2_X1 U1065 ( .A1(n1341), .A2(n1168), .ZN(n1340) );
INV_X1 U1066 ( .A(G902), .ZN(n1168) );
XOR2_X1 U1067 ( .A(n1342), .B(n1343), .Z(n1341) );
XOR2_X1 U1068 ( .A(n1344), .B(n1345), .Z(n1343) );
INV_X1 U1069 ( .A(n1133), .ZN(n1345) );
XOR2_X1 U1070 ( .A(n1346), .B(G101), .Z(n1133) );
NAND2_X1 U1071 ( .A1(G210), .A2(n1282), .ZN(n1346) );
NOR2_X1 U1072 ( .A1(G953), .A2(G237), .ZN(n1282) );
NAND2_X1 U1073 ( .A1(n1347), .A2(KEYINPUT37), .ZN(n1344) );
XOR2_X1 U1074 ( .A(n1140), .B(n1348), .Z(n1347) );
NOR2_X1 U1075 ( .A1(KEYINPUT46), .A2(n1096), .ZN(n1348) );
XOR2_X1 U1076 ( .A(n1337), .B(n1285), .Z(n1096) );
XNOR2_X1 U1077 ( .A(G143), .B(KEYINPUT10), .ZN(n1285) );
XOR2_X1 U1078 ( .A(G128), .B(n1217), .Z(n1337) );
INV_X1 U1079 ( .A(G146), .ZN(n1217) );
XOR2_X1 U1080 ( .A(n1349), .B(n1350), .Z(n1140) );
XOR2_X1 U1081 ( .A(G116), .B(G113), .Z(n1350) );
XOR2_X1 U1082 ( .A(n1351), .B(n1270), .Z(n1349) );
INV_X1 U1083 ( .A(n1145), .ZN(n1270) );
XOR2_X1 U1084 ( .A(n1095), .B(KEYINPUT41), .Z(n1145) );
XNOR2_X1 U1085 ( .A(G131), .B(n1352), .ZN(n1095) );
XOR2_X1 U1086 ( .A(G137), .B(G134), .Z(n1352) );
NAND2_X1 U1087 ( .A1(n1353), .A2(KEYINPUT26), .ZN(n1351) );
XOR2_X1 U1088 ( .A(n1258), .B(KEYINPUT15), .Z(n1353) );
INV_X1 U1089 ( .A(G119), .ZN(n1258) );
XNOR2_X1 U1090 ( .A(KEYINPUT56), .B(KEYINPUT35), .ZN(n1342) );
INV_X1 U1091 ( .A(G110), .ZN(n1263) );
endmodule


