//Key = 1110000110001010101100110100101001111010111100110001011101000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347;

XNOR2_X1 U751 ( .A(G107), .B(n1026), .ZN(G9) );
NOR2_X1 U752 ( .A1(n1027), .A2(n1028), .ZN(G75) );
NOR4_X1 U753 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1028) );
NOR2_X1 U754 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U755 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR3_X1 U756 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NOR3_X1 U757 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
NOR2_X1 U758 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR3_X1 U759 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1043) );
NOR3_X1 U760 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
INV_X1 U761 ( .A(KEYINPUT0), .ZN(n1048) );
NOR2_X1 U762 ( .A1(KEYINPUT0), .A2(n1051), .ZN(n1046) );
AND2_X1 U763 ( .A1(n1052), .A2(KEYINPUT51), .ZN(n1045) );
NOR2_X1 U764 ( .A1(n1053), .A2(n1051), .ZN(n1041) );
NOR2_X1 U765 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U766 ( .A1(n1056), .A2(n1057), .ZN(n1038) );
NOR3_X1 U767 ( .A1(n1044), .A2(KEYINPUT51), .A3(n1058), .ZN(n1057) );
INV_X1 U768 ( .A(n1040), .ZN(n1056) );
NOR4_X1 U769 ( .A1(n1059), .A2(n1044), .A3(n1051), .A4(n1040), .ZN(n1035) );
INV_X1 U770 ( .A(n1060), .ZN(n1044) );
NOR2_X1 U771 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NAND3_X1 U772 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1029) );
NAND4_X1 U773 ( .A1(n1060), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1065) );
NOR2_X1 U774 ( .A1(n1037), .A2(n1040), .ZN(n1068) );
XNOR2_X1 U775 ( .A(n1069), .B(n1070), .ZN(n1066) );
NOR2_X1 U776 ( .A1(KEYINPUT59), .A2(n1071), .ZN(n1069) );
AND3_X1 U777 ( .A1(n1063), .A2(n1064), .A3(n1072), .ZN(n1027) );
NAND4_X1 U778 ( .A1(n1073), .A2(n1070), .A3(n1074), .A4(n1075), .ZN(n1063) );
NOR3_X1 U779 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NOR2_X1 U780 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XNOR2_X1 U781 ( .A(KEYINPUT35), .B(n1081), .ZN(n1080) );
NOR2_X1 U782 ( .A1(n1082), .A2(n1083), .ZN(n1077) );
XNOR2_X1 U783 ( .A(KEYINPUT22), .B(n1084), .ZN(n1083) );
NAND3_X1 U784 ( .A1(n1085), .A2(n1086), .A3(n1071), .ZN(n1076) );
NOR3_X1 U785 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1074) );
XOR2_X1 U786 ( .A(n1050), .B(KEYINPUT61), .Z(n1088) );
XOR2_X1 U787 ( .A(n1090), .B(n1091), .Z(G72) );
NOR2_X1 U788 ( .A1(n1092), .A2(n1064), .ZN(n1091) );
NOR2_X1 U789 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XNOR2_X1 U790 ( .A(G227), .B(KEYINPUT58), .ZN(n1093) );
NAND2_X1 U791 ( .A1(n1095), .A2(n1096), .ZN(n1090) );
NAND2_X1 U792 ( .A1(n1097), .A2(n1064), .ZN(n1096) );
XOR2_X1 U793 ( .A(n1030), .B(n1098), .Z(n1097) );
NAND3_X1 U794 ( .A1(G900), .A2(n1098), .A3(G953), .ZN(n1095) );
XNOR2_X1 U795 ( .A(n1099), .B(n1100), .ZN(n1098) );
XNOR2_X1 U796 ( .A(n1101), .B(n1102), .ZN(n1099) );
NOR2_X1 U797 ( .A1(KEYINPUT11), .A2(n1103), .ZN(n1102) );
XNOR2_X1 U798 ( .A(n1104), .B(n1105), .ZN(n1103) );
XOR2_X1 U799 ( .A(n1106), .B(n1107), .Z(G69) );
XOR2_X1 U800 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR3_X1 U801 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
NOR2_X1 U802 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U803 ( .A(KEYINPUT40), .B(n1115), .Z(n1114) );
NOR2_X1 U804 ( .A1(n1115), .A2(n1116), .ZN(n1111) );
AND2_X1 U805 ( .A1(n1117), .A2(n1118), .ZN(n1115) );
XOR2_X1 U806 ( .A(n1119), .B(KEYINPUT48), .Z(n1117) );
NAND2_X1 U807 ( .A1(n1120), .A2(n1032), .ZN(n1108) );
XNOR2_X1 U808 ( .A(G953), .B(KEYINPUT44), .ZN(n1120) );
NAND2_X1 U809 ( .A1(G953), .A2(n1121), .ZN(n1106) );
NAND2_X1 U810 ( .A1(G898), .A2(G224), .ZN(n1121) );
NOR2_X1 U811 ( .A1(n1122), .A2(n1123), .ZN(G66) );
XOR2_X1 U812 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U813 ( .A(KEYINPUT15), .B(n1126), .Z(n1125) );
NOR2_X1 U814 ( .A1(n1081), .A2(n1127), .ZN(n1126) );
NOR2_X1 U815 ( .A1(n1122), .A2(n1128), .ZN(G63) );
XNOR2_X1 U816 ( .A(n1129), .B(n1130), .ZN(n1128) );
NOR2_X1 U817 ( .A1(n1131), .A2(n1127), .ZN(n1130) );
NOR2_X1 U818 ( .A1(n1122), .A2(n1132), .ZN(G60) );
XOR2_X1 U819 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR3_X1 U820 ( .A1(n1127), .A2(KEYINPUT24), .A3(n1135), .ZN(n1133) );
XNOR2_X1 U821 ( .A(G104), .B(n1136), .ZN(G6) );
NOR2_X1 U822 ( .A1(n1122), .A2(n1137), .ZN(G57) );
XOR2_X1 U823 ( .A(n1138), .B(n1139), .Z(n1137) );
XNOR2_X1 U824 ( .A(n1140), .B(n1141), .ZN(n1139) );
NAND2_X1 U825 ( .A1(KEYINPUT57), .A2(n1142), .ZN(n1140) );
XOR2_X1 U826 ( .A(n1143), .B(n1144), .Z(n1138) );
NOR2_X1 U827 ( .A1(G101), .A2(KEYINPUT13), .ZN(n1144) );
XNOR2_X1 U828 ( .A(n1145), .B(n1146), .ZN(n1143) );
NOR3_X1 U829 ( .A1(n1127), .A2(KEYINPUT9), .A3(n1084), .ZN(n1146) );
NOR2_X1 U830 ( .A1(n1122), .A2(n1147), .ZN(G54) );
XOR2_X1 U831 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U832 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U833 ( .A(n1152), .B(n1153), .Z(n1148) );
NOR2_X1 U834 ( .A1(n1154), .A2(n1127), .ZN(n1153) );
NAND2_X1 U835 ( .A1(KEYINPUT12), .A2(n1155), .ZN(n1152) );
NOR2_X1 U836 ( .A1(n1122), .A2(n1156), .ZN(G51) );
XOR2_X1 U837 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U838 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U839 ( .A1(n1161), .A2(n1127), .ZN(n1160) );
NAND2_X1 U840 ( .A1(G902), .A2(n1162), .ZN(n1127) );
NAND2_X1 U841 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
INV_X1 U842 ( .A(n1032), .ZN(n1164) );
NAND4_X1 U843 ( .A1(n1165), .A2(n1136), .A3(n1166), .A4(n1167), .ZN(n1032) );
AND4_X1 U844 ( .A1(n1026), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1167) );
NAND3_X1 U845 ( .A1(n1060), .A2(n1061), .A3(n1171), .ZN(n1026) );
AND2_X1 U846 ( .A1(n1172), .A2(n1173), .ZN(n1166) );
NAND3_X1 U847 ( .A1(n1171), .A2(n1060), .A3(n1062), .ZN(n1136) );
NAND2_X1 U848 ( .A1(n1174), .A2(n1052), .ZN(n1165) );
XOR2_X1 U849 ( .A(n1175), .B(KEYINPUT30), .Z(n1174) );
NAND4_X1 U850 ( .A1(n1176), .A2(n1177), .A3(n1060), .A4(n1178), .ZN(n1175) );
XNOR2_X1 U851 ( .A(KEYINPUT38), .B(n1179), .ZN(n1176) );
XOR2_X1 U852 ( .A(n1030), .B(KEYINPUT34), .Z(n1163) );
NAND4_X1 U853 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1030) );
AND3_X1 U854 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1183) );
NAND2_X1 U855 ( .A1(n1187), .A2(n1188), .ZN(n1182) );
NAND2_X1 U856 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND3_X1 U857 ( .A1(n1191), .A2(n1192), .A3(n1062), .ZN(n1190) );
NAND2_X1 U858 ( .A1(n1193), .A2(n1194), .ZN(n1189) );
NAND2_X1 U859 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NAND2_X1 U860 ( .A1(n1052), .A2(n1197), .ZN(n1196) );
NAND2_X1 U861 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NAND2_X1 U862 ( .A1(n1062), .A2(n1191), .ZN(n1199) );
NAND2_X1 U863 ( .A1(n1192), .A2(n1200), .ZN(n1191) );
NAND2_X1 U864 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
INV_X1 U865 ( .A(KEYINPUT8), .ZN(n1192) );
NAND2_X1 U866 ( .A1(n1203), .A2(n1067), .ZN(n1195) );
NOR2_X1 U867 ( .A1(n1204), .A2(n1205), .ZN(n1159) );
NOR3_X1 U868 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1205) );
NOR2_X1 U869 ( .A1(n1100), .A2(n1209), .ZN(n1208) );
NOR2_X1 U870 ( .A1(n1210), .A2(n1211), .ZN(n1207) );
NOR2_X1 U871 ( .A1(KEYINPUT21), .A2(G125), .ZN(n1206) );
NOR4_X1 U872 ( .A1(n1212), .A2(n1213), .A3(KEYINPUT21), .A4(G125), .ZN(n1204) );
NOR2_X1 U873 ( .A1(n1209), .A2(n1211), .ZN(n1213) );
XOR2_X1 U874 ( .A(n1214), .B(n1210), .Z(n1209) );
XNOR2_X1 U875 ( .A(KEYINPUT63), .B(KEYINPUT52), .ZN(n1214) );
NOR2_X1 U876 ( .A1(n1100), .A2(n1210), .ZN(n1212) );
XNOR2_X1 U877 ( .A(n1215), .B(KEYINPUT62), .ZN(n1210) );
NOR2_X1 U878 ( .A1(KEYINPUT49), .A2(n1216), .ZN(n1157) );
AND2_X1 U879 ( .A1(n1217), .A2(n1072), .ZN(n1122) );
INV_X1 U880 ( .A(G952), .ZN(n1072) );
XNOR2_X1 U881 ( .A(KEYINPUT26), .B(n1064), .ZN(n1217) );
XOR2_X1 U882 ( .A(G146), .B(n1218), .Z(G48) );
NOR4_X1 U883 ( .A1(n1058), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1218) );
XNOR2_X1 U884 ( .A(KEYINPUT42), .B(n1222), .ZN(n1221) );
XNOR2_X1 U885 ( .A(G143), .B(n1180), .ZN(G45) );
NAND4_X1 U886 ( .A1(n1055), .A2(n1193), .A3(n1052), .A4(n1179), .ZN(n1180) );
XNOR2_X1 U887 ( .A(G140), .B(n1181), .ZN(G42) );
NAND3_X1 U888 ( .A1(n1062), .A2(n1054), .A3(n1223), .ZN(n1181) );
NAND2_X1 U889 ( .A1(n1224), .A2(n1225), .ZN(G39) );
NAND2_X1 U890 ( .A1(n1226), .A2(G137), .ZN(n1225) );
XOR2_X1 U891 ( .A(KEYINPUT7), .B(n1227), .Z(n1224) );
NOR2_X1 U892 ( .A1(G137), .A2(n1226), .ZN(n1227) );
AND2_X1 U893 ( .A1(n1228), .A2(n1229), .ZN(n1226) );
NAND4_X1 U894 ( .A1(n1203), .A2(n1223), .A3(n1187), .A4(n1230), .ZN(n1229) );
INV_X1 U895 ( .A(KEYINPUT3), .ZN(n1230) );
NAND3_X1 U896 ( .A1(n1067), .A2(n1231), .A3(KEYINPUT3), .ZN(n1228) );
NAND3_X1 U897 ( .A1(n1203), .A2(n1193), .A3(n1187), .ZN(n1231) );
INV_X1 U898 ( .A(n1220), .ZN(n1193) );
INV_X1 U899 ( .A(n1051), .ZN(n1067) );
XNOR2_X1 U900 ( .A(G134), .B(n1184), .ZN(G36) );
NAND3_X1 U901 ( .A1(n1223), .A2(n1061), .A3(n1055), .ZN(n1184) );
XNOR2_X1 U902 ( .A(G131), .B(n1186), .ZN(G33) );
NAND3_X1 U903 ( .A1(n1223), .A2(n1062), .A3(n1055), .ZN(n1186) );
NOR2_X1 U904 ( .A1(n1220), .A2(n1051), .ZN(n1223) );
NAND2_X1 U905 ( .A1(n1073), .A2(n1050), .ZN(n1051) );
INV_X1 U906 ( .A(n1049), .ZN(n1073) );
XOR2_X1 U907 ( .A(G128), .B(n1232), .Z(G30) );
NOR4_X1 U908 ( .A1(n1233), .A2(n1198), .A3(n1220), .A4(n1222), .ZN(n1232) );
NAND3_X1 U909 ( .A1(n1234), .A2(n1071), .A3(n1235), .ZN(n1220) );
INV_X1 U910 ( .A(n1061), .ZN(n1198) );
XNOR2_X1 U911 ( .A(n1052), .B(KEYINPUT6), .ZN(n1233) );
XOR2_X1 U912 ( .A(n1173), .B(n1236), .Z(G3) );
NAND2_X1 U913 ( .A1(KEYINPUT23), .A2(G101), .ZN(n1236) );
NAND3_X1 U914 ( .A1(n1055), .A2(n1171), .A3(n1203), .ZN(n1173) );
XNOR2_X1 U915 ( .A(G125), .B(n1185), .ZN(G27) );
NAND4_X1 U916 ( .A1(n1062), .A2(n1054), .A3(n1237), .A4(n1177), .ZN(n1185) );
NOR2_X1 U917 ( .A1(n1201), .A2(n1058), .ZN(n1237) );
INV_X1 U918 ( .A(n1234), .ZN(n1201) );
NAND2_X1 U919 ( .A1(n1040), .A2(n1238), .ZN(n1234) );
NAND4_X1 U920 ( .A1(G902), .A2(G953), .A3(n1239), .A4(n1094), .ZN(n1238) );
INV_X1 U921 ( .A(G900), .ZN(n1094) );
XOR2_X1 U922 ( .A(n1240), .B(n1241), .Z(G24) );
AND3_X1 U923 ( .A1(n1242), .A2(n1179), .A3(n1060), .ZN(n1241) );
NOR2_X1 U924 ( .A1(n1243), .A2(n1244), .ZN(n1060) );
NAND2_X1 U925 ( .A1(n1245), .A2(n1246), .ZN(n1179) );
OR3_X1 U926 ( .A1(n1247), .A2(n1248), .A3(KEYINPUT10), .ZN(n1246) );
NAND2_X1 U927 ( .A1(KEYINPUT10), .A2(n1061), .ZN(n1245) );
NOR2_X1 U928 ( .A1(KEYINPUT20), .A2(n1249), .ZN(n1240) );
XNOR2_X1 U929 ( .A(G119), .B(n1172), .ZN(G21) );
NAND3_X1 U930 ( .A1(n1187), .A2(n1203), .A3(n1242), .ZN(n1172) );
INV_X1 U931 ( .A(n1222), .ZN(n1187) );
NAND2_X1 U932 ( .A1(n1244), .A2(n1243), .ZN(n1222) );
XNOR2_X1 U933 ( .A(G116), .B(n1170), .ZN(G18) );
NAND3_X1 U934 ( .A1(n1055), .A2(n1061), .A3(n1242), .ZN(n1170) );
NOR2_X1 U935 ( .A1(n1247), .A2(n1250), .ZN(n1061) );
XNOR2_X1 U936 ( .A(G113), .B(n1169), .ZN(G15) );
NAND3_X1 U937 ( .A1(n1055), .A2(n1062), .A3(n1242), .ZN(n1169) );
AND3_X1 U938 ( .A1(n1052), .A2(n1178), .A3(n1177), .ZN(n1242) );
INV_X1 U939 ( .A(n1034), .ZN(n1177) );
NAND2_X1 U940 ( .A1(n1251), .A2(n1071), .ZN(n1034) );
XNOR2_X1 U941 ( .A(KEYINPUT41), .B(n1070), .ZN(n1251) );
INV_X1 U942 ( .A(n1235), .ZN(n1070) );
INV_X1 U943 ( .A(n1219), .ZN(n1062) );
NAND2_X1 U944 ( .A1(n1252), .A2(n1247), .ZN(n1219) );
XNOR2_X1 U945 ( .A(n1248), .B(KEYINPUT10), .ZN(n1252) );
NOR2_X1 U946 ( .A1(n1244), .A2(n1253), .ZN(n1055) );
XNOR2_X1 U947 ( .A(G110), .B(n1168), .ZN(G12) );
NAND3_X1 U948 ( .A1(n1054), .A2(n1171), .A3(n1203), .ZN(n1168) );
INV_X1 U949 ( .A(n1037), .ZN(n1203) );
NAND2_X1 U950 ( .A1(n1247), .A2(n1254), .ZN(n1037) );
XNOR2_X1 U951 ( .A(KEYINPUT60), .B(n1250), .ZN(n1254) );
INV_X1 U952 ( .A(n1248), .ZN(n1250) );
XOR2_X1 U953 ( .A(n1089), .B(KEYINPUT2), .Z(n1248) );
XOR2_X1 U954 ( .A(n1255), .B(n1135), .Z(n1089) );
INV_X1 U955 ( .A(G475), .ZN(n1135) );
OR2_X1 U956 ( .A1(n1134), .A2(G902), .ZN(n1255) );
XNOR2_X1 U957 ( .A(n1256), .B(n1257), .ZN(n1134) );
XNOR2_X1 U958 ( .A(n1105), .B(n1258), .ZN(n1257) );
XOR2_X1 U959 ( .A(n1259), .B(n1260), .Z(n1258) );
NAND2_X1 U960 ( .A1(n1261), .A2(G214), .ZN(n1259) );
XOR2_X1 U961 ( .A(n1262), .B(n1263), .Z(n1256) );
XNOR2_X1 U962 ( .A(n1264), .B(G104), .ZN(n1263) );
INV_X1 U963 ( .A(G113), .ZN(n1264) );
NAND2_X1 U964 ( .A1(KEYINPUT14), .A2(n1265), .ZN(n1262) );
INV_X1 U965 ( .A(n1087), .ZN(n1247) );
XNOR2_X1 U966 ( .A(n1266), .B(n1267), .ZN(n1087) );
XNOR2_X1 U967 ( .A(KEYINPUT39), .B(n1131), .ZN(n1267) );
INV_X1 U968 ( .A(G478), .ZN(n1131) );
NAND2_X1 U969 ( .A1(n1129), .A2(n1268), .ZN(n1266) );
XNOR2_X1 U970 ( .A(n1269), .B(n1270), .ZN(n1129) );
XOR2_X1 U971 ( .A(n1271), .B(n1272), .Z(n1270) );
XNOR2_X1 U972 ( .A(G116), .B(G107), .ZN(n1272) );
NAND2_X1 U973 ( .A1(KEYINPUT25), .A2(n1273), .ZN(n1271) );
XOR2_X1 U974 ( .A(n1274), .B(n1275), .Z(n1269) );
XOR2_X1 U975 ( .A(n1276), .B(n1260), .Z(n1274) );
XNOR2_X1 U976 ( .A(n1249), .B(G143), .ZN(n1260) );
INV_X1 U977 ( .A(G122), .ZN(n1249) );
NAND3_X1 U978 ( .A1(G234), .A2(n1064), .A3(G217), .ZN(n1276) );
AND2_X1 U979 ( .A1(n1202), .A2(n1178), .ZN(n1171) );
NAND2_X1 U980 ( .A1(n1040), .A2(n1277), .ZN(n1178) );
NAND3_X1 U981 ( .A1(n1110), .A2(n1239), .A3(G902), .ZN(n1277) );
NOR2_X1 U982 ( .A1(n1064), .A2(G898), .ZN(n1110) );
NAND3_X1 U983 ( .A1(n1239), .A2(n1064), .A3(G952), .ZN(n1040) );
NAND2_X1 U984 ( .A1(G237), .A2(G234), .ZN(n1239) );
AND3_X1 U985 ( .A1(n1235), .A2(n1071), .A3(n1052), .ZN(n1202) );
INV_X1 U986 ( .A(n1058), .ZN(n1052) );
NAND2_X1 U987 ( .A1(n1278), .A2(n1049), .ZN(n1058) );
XOR2_X1 U988 ( .A(n1279), .B(n1161), .Z(n1049) );
NAND2_X1 U989 ( .A1(G210), .A2(n1280), .ZN(n1161) );
NAND2_X1 U990 ( .A1(n1281), .A2(n1268), .ZN(n1279) );
XOR2_X1 U991 ( .A(n1282), .B(n1283), .Z(n1281) );
XOR2_X1 U992 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U993 ( .A(G125), .B(KEYINPUT19), .ZN(n1285) );
NAND2_X1 U994 ( .A1(KEYINPUT1), .A2(n1215), .ZN(n1284) );
AND2_X1 U995 ( .A1(G224), .A2(n1064), .ZN(n1215) );
XNOR2_X1 U996 ( .A(n1216), .B(n1211), .ZN(n1282) );
XNOR2_X1 U997 ( .A(n1286), .B(n1116), .ZN(n1216) );
INV_X1 U998 ( .A(n1113), .ZN(n1116) );
XNOR2_X1 U999 ( .A(G122), .B(n1287), .ZN(n1113) );
NAND2_X1 U1000 ( .A1(n1118), .A2(n1119), .ZN(n1286) );
NAND2_X1 U1001 ( .A1(n1288), .A2(n1289), .ZN(n1119) );
XNOR2_X1 U1002 ( .A(KEYINPUT56), .B(n1290), .ZN(n1289) );
XNOR2_X1 U1003 ( .A(G101), .B(n1291), .ZN(n1288) );
NAND2_X1 U1004 ( .A1(n1292), .A2(n1293), .ZN(n1118) );
XNOR2_X1 U1005 ( .A(n1141), .B(KEYINPUT56), .ZN(n1293) );
XNOR2_X1 U1006 ( .A(n1291), .B(n1294), .ZN(n1292) );
NAND2_X1 U1007 ( .A1(KEYINPUT28), .A2(n1295), .ZN(n1291) );
XNOR2_X1 U1008 ( .A(n1296), .B(G104), .ZN(n1295) );
XNOR2_X1 U1009 ( .A(KEYINPUT18), .B(n1050), .ZN(n1278) );
NAND2_X1 U1010 ( .A1(G214), .A2(n1280), .ZN(n1050) );
NAND2_X1 U1011 ( .A1(n1297), .A2(n1268), .ZN(n1280) );
INV_X1 U1012 ( .A(G237), .ZN(n1297) );
NAND2_X1 U1013 ( .A1(G221), .A2(n1298), .ZN(n1071) );
XOR2_X1 U1014 ( .A(n1299), .B(n1154), .Z(n1235) );
INV_X1 U1015 ( .A(G469), .ZN(n1154) );
NAND2_X1 U1016 ( .A1(n1300), .A2(n1268), .ZN(n1299) );
XOR2_X1 U1017 ( .A(n1301), .B(n1151), .Z(n1300) );
XNOR2_X1 U1018 ( .A(G140), .B(n1287), .ZN(n1151) );
INV_X1 U1019 ( .A(G110), .ZN(n1287) );
XNOR2_X1 U1020 ( .A(n1155), .B(n1302), .ZN(n1301) );
NOR2_X1 U1021 ( .A1(KEYINPUT5), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1022 ( .A(n1150), .B(n1304), .Z(n1303) );
XOR2_X1 U1023 ( .A(KEYINPUT4), .B(KEYINPUT29), .Z(n1304) );
XOR2_X1 U1024 ( .A(n1305), .B(n1306), .Z(n1150) );
XNOR2_X1 U1025 ( .A(n1296), .B(G101), .ZN(n1306) );
INV_X1 U1026 ( .A(G107), .ZN(n1296) );
XNOR2_X1 U1027 ( .A(n1307), .B(n1142), .ZN(n1305) );
NAND2_X1 U1028 ( .A1(KEYINPUT16), .A2(n1308), .ZN(n1307) );
INV_X1 U1029 ( .A(G104), .ZN(n1308) );
AND2_X1 U1030 ( .A1(G227), .A2(n1064), .ZN(n1155) );
AND2_X1 U1031 ( .A1(n1253), .A2(n1244), .ZN(n1054) );
NAND2_X1 U1032 ( .A1(n1309), .A2(n1085), .ZN(n1244) );
NAND2_X1 U1033 ( .A1(n1079), .A2(n1081), .ZN(n1085) );
OR2_X1 U1034 ( .A1(n1081), .A2(n1079), .ZN(n1309) );
NOR2_X1 U1035 ( .A1(n1124), .A2(G902), .ZN(n1079) );
XNOR2_X1 U1036 ( .A(n1310), .B(n1311), .ZN(n1124) );
XOR2_X1 U1037 ( .A(n1312), .B(n1265), .Z(n1311) );
XNOR2_X1 U1038 ( .A(G146), .B(n1101), .ZN(n1265) );
XOR2_X1 U1039 ( .A(G140), .B(G125), .Z(n1101) );
NAND2_X1 U1040 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
NAND4_X1 U1041 ( .A1(G221), .A2(G234), .A3(n1315), .A4(n1064), .ZN(n1314) );
NAND2_X1 U1042 ( .A1(n1316), .A2(n1317), .ZN(n1313) );
NAND3_X1 U1043 ( .A1(G234), .A2(n1064), .A3(G221), .ZN(n1317) );
INV_X1 U1044 ( .A(G953), .ZN(n1064) );
XOR2_X1 U1045 ( .A(KEYINPUT36), .B(n1315), .Z(n1316) );
XOR2_X1 U1046 ( .A(G137), .B(KEYINPUT31), .Z(n1315) );
XNOR2_X1 U1047 ( .A(KEYINPUT47), .B(n1318), .ZN(n1310) );
NOR2_X1 U1048 ( .A1(KEYINPUT17), .A2(n1319), .ZN(n1318) );
XNOR2_X1 U1049 ( .A(n1320), .B(n1321), .ZN(n1319) );
XNOR2_X1 U1050 ( .A(G110), .B(n1322), .ZN(n1321) );
NOR2_X1 U1051 ( .A1(G119), .A2(KEYINPUT32), .ZN(n1322) );
NAND2_X1 U1052 ( .A1(G217), .A2(n1298), .ZN(n1081) );
NAND2_X1 U1053 ( .A1(G234), .A2(n1268), .ZN(n1298) );
INV_X1 U1054 ( .A(n1243), .ZN(n1253) );
NAND2_X1 U1055 ( .A1(n1323), .A2(n1086), .ZN(n1243) );
NAND2_X1 U1056 ( .A1(n1082), .A2(n1084), .ZN(n1086) );
INV_X1 U1057 ( .A(G472), .ZN(n1084) );
INV_X1 U1058 ( .A(n1324), .ZN(n1082) );
NAND2_X1 U1059 ( .A1(n1325), .A2(n1324), .ZN(n1323) );
NAND2_X1 U1060 ( .A1(n1326), .A2(n1268), .ZN(n1324) );
INV_X1 U1061 ( .A(G902), .ZN(n1268) );
XOR2_X1 U1062 ( .A(n1327), .B(n1328), .Z(n1326) );
NOR2_X1 U1063 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XOR2_X1 U1064 ( .A(n1331), .B(KEYINPUT55), .Z(n1330) );
NAND2_X1 U1065 ( .A1(n1332), .A2(n1290), .ZN(n1331) );
NOR2_X1 U1066 ( .A1(n1290), .A2(n1332), .ZN(n1329) );
XNOR2_X1 U1067 ( .A(KEYINPUT46), .B(n1142), .ZN(n1332) );
XOR2_X1 U1068 ( .A(n1333), .B(n1334), .Z(n1142) );
XNOR2_X1 U1069 ( .A(n1105), .B(n1211), .ZN(n1334) );
INV_X1 U1070 ( .A(n1100), .ZN(n1211) );
XNOR2_X1 U1071 ( .A(n1335), .B(n1336), .ZN(n1100) );
XNOR2_X1 U1072 ( .A(G143), .B(n1273), .ZN(n1336) );
INV_X1 U1073 ( .A(n1320), .ZN(n1273) );
XOR2_X1 U1074 ( .A(G128), .B(KEYINPUT50), .Z(n1320) );
XNOR2_X1 U1075 ( .A(G146), .B(KEYINPUT27), .ZN(n1335) );
XOR2_X1 U1076 ( .A(G131), .B(KEYINPUT45), .Z(n1105) );
NAND2_X1 U1077 ( .A1(n1337), .A2(n1338), .ZN(n1333) );
OR3_X1 U1078 ( .A1(n1275), .A2(G137), .A3(KEYINPUT53), .ZN(n1338) );
NAND2_X1 U1079 ( .A1(n1104), .A2(KEYINPUT53), .ZN(n1337) );
XOR2_X1 U1080 ( .A(G137), .B(n1275), .Z(n1104) );
XOR2_X1 U1081 ( .A(G134), .B(KEYINPUT43), .Z(n1275) );
INV_X1 U1082 ( .A(n1141), .ZN(n1290) );
XOR2_X1 U1083 ( .A(G113), .B(n1339), .Z(n1141) );
XOR2_X1 U1084 ( .A(G119), .B(G116), .Z(n1339) );
NAND2_X1 U1085 ( .A1(n1340), .A2(n1341), .ZN(n1327) );
NAND2_X1 U1086 ( .A1(G101), .A2(n1342), .ZN(n1341) );
NAND2_X1 U1087 ( .A1(KEYINPUT54), .A2(n1343), .ZN(n1342) );
NAND2_X1 U1088 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
NAND2_X1 U1089 ( .A1(n1145), .A2(n1346), .ZN(n1340) );
NAND2_X1 U1090 ( .A1(n1347), .A2(n1345), .ZN(n1346) );
INV_X1 U1091 ( .A(KEYINPUT37), .ZN(n1345) );
NAND2_X1 U1092 ( .A1(KEYINPUT54), .A2(n1294), .ZN(n1347) );
INV_X1 U1093 ( .A(G101), .ZN(n1294) );
INV_X1 U1094 ( .A(n1344), .ZN(n1145) );
NAND2_X1 U1095 ( .A1(n1261), .A2(G210), .ZN(n1344) );
NOR2_X1 U1096 ( .A1(G953), .A2(G237), .ZN(n1261) );
XNOR2_X1 U1097 ( .A(G472), .B(KEYINPUT33), .ZN(n1325) );
endmodule


