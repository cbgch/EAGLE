//Key = 0110001110011010101010110100010101011011010111111000010100110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285;

XOR2_X1 U714 ( .A(G107), .B(n985), .Z(G9) );
NOR2_X1 U715 ( .A1(n986), .A2(n987), .ZN(G75) );
NOR4_X1 U716 ( .A1(n988), .A2(n989), .A3(n990), .A4(n991), .ZN(n987) );
XOR2_X1 U717 ( .A(KEYINPUT30), .B(n992), .Z(n989) );
NOR2_X1 U718 ( .A1(n993), .A2(n994), .ZN(n992) );
XOR2_X1 U719 ( .A(n995), .B(KEYINPUT52), .Z(n993) );
NAND4_X1 U720 ( .A1(n996), .A2(n997), .A3(n998), .A4(n999), .ZN(n995) );
XOR2_X1 U721 ( .A(KEYINPUT54), .B(n1000), .Z(n998) );
NAND3_X1 U722 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n988) );
NAND2_X1 U723 ( .A1(n996), .A2(n1004), .ZN(n1003) );
NAND2_X1 U724 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND3_X1 U725 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1006) );
NAND2_X1 U726 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NAND2_X1 U727 ( .A1(n1000), .A2(n1012), .ZN(n1011) );
OR2_X1 U728 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U729 ( .A1(n999), .A2(n1015), .ZN(n1010) );
NAND2_X1 U730 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U731 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND3_X1 U732 ( .A1(n999), .A2(n1020), .A3(n1000), .ZN(n1005) );
NAND2_X1 U733 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND3_X1 U734 ( .A1(n1023), .A2(n1024), .A3(n1009), .ZN(n1022) );
NAND2_X1 U735 ( .A1(n1007), .A2(n1025), .ZN(n1021) );
NAND2_X1 U736 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U737 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
INV_X1 U738 ( .A(n1030), .ZN(n1026) );
INV_X1 U739 ( .A(n1031), .ZN(n996) );
AND3_X1 U740 ( .A1(n1001), .A2(n1002), .A3(n1032), .ZN(n986) );
NAND4_X1 U741 ( .A1(n1033), .A2(n1007), .A3(n1034), .A4(n1035), .ZN(n1001) );
NOR4_X1 U742 ( .A1(n1028), .A2(n1018), .A3(n1036), .A4(n1037), .ZN(n1035) );
XNOR2_X1 U743 ( .A(n1038), .B(n1039), .ZN(n1036) );
XOR2_X1 U744 ( .A(n1040), .B(n1041), .Z(n1034) );
NOR2_X1 U745 ( .A1(KEYINPUT34), .A2(n1042), .ZN(n1041) );
NAND2_X1 U746 ( .A1(n1043), .A2(n1044), .ZN(G72) );
NAND3_X1 U747 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NAND2_X1 U748 ( .A1(n1048), .A2(n1049), .ZN(n1045) );
NAND3_X1 U749 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1043) );
XNOR2_X1 U750 ( .A(n1053), .B(n1048), .ZN(n1052) );
XNOR2_X1 U751 ( .A(n1054), .B(n1055), .ZN(n1048) );
XOR2_X1 U752 ( .A(n1056), .B(n1057), .Z(n1055) );
XNOR2_X1 U753 ( .A(G140), .B(KEYINPUT44), .ZN(n1057) );
NAND2_X1 U754 ( .A1(KEYINPUT53), .A2(n1058), .ZN(n1056) );
XOR2_X1 U755 ( .A(n1059), .B(n1060), .Z(n1054) );
NAND2_X1 U756 ( .A1(n1002), .A2(n1061), .ZN(n1053) );
NAND3_X1 U757 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
XNOR2_X1 U758 ( .A(n1065), .B(KEYINPUT8), .ZN(n1062) );
NAND2_X1 U759 ( .A1(G953), .A2(n1066), .ZN(n1051) );
NAND2_X1 U760 ( .A1(n1049), .A2(n1067), .ZN(n1066) );
NAND2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U762 ( .A1(n1069), .A2(n1070), .ZN(n1050) );
INV_X1 U763 ( .A(KEYINPUT45), .ZN(n1070) );
NAND2_X1 U764 ( .A1(n1047), .A2(n1071), .ZN(n1069) );
NAND2_X1 U765 ( .A1(KEYINPUT45), .A2(n1046), .ZN(n1071) );
INV_X1 U766 ( .A(KEYINPUT51), .ZN(n1046) );
AND2_X1 U767 ( .A1(G953), .A2(n1068), .ZN(n1047) );
NAND2_X1 U768 ( .A1(G900), .A2(G227), .ZN(n1068) );
NAND2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(G69) );
NAND2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U771 ( .A1(G953), .A2(n1076), .ZN(n1075) );
NAND2_X1 U772 ( .A1(G898), .A2(G224), .ZN(n1076) );
NAND2_X1 U773 ( .A1(n1077), .A2(n1078), .ZN(n1072) );
NAND2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U775 ( .A1(G953), .A2(n1081), .ZN(n1080) );
INV_X1 U776 ( .A(n1082), .ZN(n1079) );
INV_X1 U777 ( .A(n1074), .ZN(n1077) );
XNOR2_X1 U778 ( .A(n1083), .B(n1084), .ZN(n1074) );
NOR2_X1 U779 ( .A1(n1082), .A2(n1085), .ZN(n1084) );
XNOR2_X1 U780 ( .A(n1086), .B(n1087), .ZN(n1085) );
NAND3_X1 U781 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1083) );
XNOR2_X1 U782 ( .A(KEYINPUT58), .B(n1002), .ZN(n1090) );
NAND2_X1 U783 ( .A1(n985), .A2(n1091), .ZN(n1089) );
OR2_X1 U784 ( .A1(n1091), .A2(n990), .ZN(n1088) );
INV_X1 U785 ( .A(KEYINPUT38), .ZN(n1091) );
NOR2_X1 U786 ( .A1(n1092), .A2(n1093), .ZN(G66) );
XNOR2_X1 U787 ( .A(n1094), .B(n1095), .ZN(n1093) );
NOR2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NOR2_X1 U789 ( .A1(n1092), .A2(n1098), .ZN(G63) );
XOR2_X1 U790 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U791 ( .A1(n1101), .A2(n1097), .ZN(n1100) );
NOR2_X1 U792 ( .A1(KEYINPUT62), .A2(n1102), .ZN(n1099) );
NOR2_X1 U793 ( .A1(n1092), .A2(n1103), .ZN(G60) );
XOR2_X1 U794 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND4_X1 U795 ( .A1(KEYINPUT33), .A2(G475), .A3(G902), .A4(n1106), .ZN(n1104) );
XOR2_X1 U796 ( .A(KEYINPUT25), .B(n1107), .Z(n1106) );
XNOR2_X1 U797 ( .A(G104), .B(n1108), .ZN(G6) );
NOR2_X1 U798 ( .A1(n1092), .A2(n1109), .ZN(G57) );
XOR2_X1 U799 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U800 ( .A1(n1112), .A2(n1097), .ZN(n1111) );
XOR2_X1 U801 ( .A(n1113), .B(n1114), .Z(n1110) );
NOR2_X1 U802 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U803 ( .A(n1117), .B(KEYINPUT46), .Z(n1116) );
NAND2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U805 ( .A1(n1119), .A2(n1118), .ZN(n1115) );
XOR2_X1 U806 ( .A(n1120), .B(n1060), .Z(n1118) );
NOR2_X1 U807 ( .A1(KEYINPUT50), .A2(n1121), .ZN(n1120) );
NAND2_X1 U808 ( .A1(n1122), .A2(KEYINPUT2), .ZN(n1113) );
XOR2_X1 U809 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U810 ( .A1(KEYINPUT1), .A2(n1125), .ZN(n1123) );
NOR2_X1 U811 ( .A1(n1092), .A2(n1126), .ZN(G54) );
XOR2_X1 U812 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U813 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U814 ( .A(n1131), .B(n1060), .Z(n1130) );
NOR2_X1 U815 ( .A1(n1132), .A2(n1097), .ZN(n1131) );
XOR2_X1 U816 ( .A(n1133), .B(n1134), .Z(n1127) );
XOR2_X1 U817 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U818 ( .A1(KEYINPUT42), .A2(n1137), .ZN(n1135) );
XNOR2_X1 U819 ( .A(G140), .B(KEYINPUT59), .ZN(n1137) );
XNOR2_X1 U820 ( .A(KEYINPUT6), .B(n1138), .ZN(n1133) );
NOR3_X1 U821 ( .A1(n1092), .A2(n1139), .A3(n1140), .ZN(G51) );
NOR2_X1 U822 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XOR2_X1 U823 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U824 ( .A1(KEYINPUT29), .A2(n1145), .ZN(n1143) );
INV_X1 U825 ( .A(n1146), .ZN(n1145) );
INV_X1 U826 ( .A(KEYINPUT12), .ZN(n1141) );
NOR2_X1 U827 ( .A1(KEYINPUT12), .A2(n1147), .ZN(n1139) );
XOR2_X1 U828 ( .A(n1148), .B(n1144), .Z(n1147) );
XNOR2_X1 U829 ( .A(n1149), .B(n1150), .ZN(n1144) );
NOR2_X1 U830 ( .A1(n1040), .A2(n1097), .ZN(n1150) );
OR2_X1 U831 ( .A1(n1151), .A2(n1107), .ZN(n1097) );
NOR2_X1 U832 ( .A1(n991), .A2(n1152), .ZN(n1107) );
XOR2_X1 U833 ( .A(KEYINPUT3), .B(n990), .Z(n1152) );
NAND2_X1 U834 ( .A1(n1153), .A2(n1154), .ZN(n990) );
NOR4_X1 U835 ( .A1(n985), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1154) );
INV_X1 U836 ( .A(n1158), .ZN(n1155) );
AND3_X1 U837 ( .A1(n1014), .A2(n1007), .A3(n1159), .ZN(n985) );
AND4_X1 U838 ( .A1(n1160), .A2(n1161), .A3(n1108), .A4(n1162), .ZN(n1153) );
NAND2_X1 U839 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NAND3_X1 U840 ( .A1(n1159), .A2(n1007), .A3(n1013), .ZN(n1108) );
NAND3_X1 U841 ( .A1(n1165), .A2(n1065), .A3(n1064), .ZN(n991) );
NOR3_X1 U842 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1064) );
AND4_X1 U843 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1065) );
XOR2_X1 U844 ( .A(n1063), .B(KEYINPUT60), .Z(n1165) );
NAND2_X1 U845 ( .A1(KEYINPUT29), .A2(n1146), .ZN(n1148) );
AND2_X1 U846 ( .A1(n1173), .A2(n1032), .ZN(n1092) );
INV_X1 U847 ( .A(G952), .ZN(n1032) );
XNOR2_X1 U848 ( .A(KEYINPUT10), .B(n1002), .ZN(n1173) );
XNOR2_X1 U849 ( .A(G146), .B(n1170), .ZN(G48) );
NAND3_X1 U850 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1170) );
XOR2_X1 U851 ( .A(n1177), .B(G143), .Z(G45) );
NAND2_X1 U852 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
OR2_X1 U853 ( .A1(n1169), .A2(KEYINPUT21), .ZN(n1179) );
NAND2_X1 U854 ( .A1(n1180), .A2(n1174), .ZN(n1169) );
NAND3_X1 U855 ( .A1(n1180), .A2(n1016), .A3(KEYINPUT21), .ZN(n1178) );
INV_X1 U856 ( .A(n1174), .ZN(n1016) );
AND4_X1 U857 ( .A1(n997), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1180) );
XNOR2_X1 U858 ( .A(G140), .B(n1171), .ZN(G42) );
NAND4_X1 U859 ( .A1(n1013), .A2(n1184), .A3(n1023), .A4(n1024), .ZN(n1171) );
XNOR2_X1 U860 ( .A(G137), .B(n1185), .ZN(G39) );
NAND2_X1 U861 ( .A1(KEYINPUT41), .A2(n1186), .ZN(n1185) );
INV_X1 U862 ( .A(n1172), .ZN(n1186) );
NAND2_X1 U863 ( .A1(n1163), .A2(n1184), .ZN(n1172) );
XOR2_X1 U864 ( .A(G134), .B(n1166), .Z(G36) );
AND3_X1 U865 ( .A1(n1184), .A2(n1014), .A3(n997), .ZN(n1166) );
XNOR2_X1 U866 ( .A(n1168), .B(n1187), .ZN(G33) );
XOR2_X1 U867 ( .A(KEYINPUT55), .B(G131), .Z(n1187) );
AND3_X1 U868 ( .A1(n1013), .A2(n1184), .A3(n997), .ZN(n1168) );
AND3_X1 U869 ( .A1(n1174), .A2(n1188), .A3(n1009), .ZN(n1184) );
INV_X1 U870 ( .A(n994), .ZN(n1009) );
NAND2_X1 U871 ( .A1(n1029), .A2(n1189), .ZN(n994) );
XNOR2_X1 U872 ( .A(n1167), .B(n1190), .ZN(G30) );
XNOR2_X1 U873 ( .A(G128), .B(KEYINPUT32), .ZN(n1190) );
AND3_X1 U874 ( .A1(n1181), .A2(n1014), .A3(n1191), .ZN(n1167) );
AND3_X1 U875 ( .A1(n1174), .A2(n1175), .A3(n1024), .ZN(n1191) );
XNOR2_X1 U876 ( .A(G101), .B(n1161), .ZN(G3) );
NAND3_X1 U877 ( .A1(n1159), .A2(n999), .A3(n997), .ZN(n1161) );
XNOR2_X1 U878 ( .A(G125), .B(n1063), .ZN(G27) );
NAND3_X1 U879 ( .A1(n1023), .A2(n1176), .A3(n1000), .ZN(n1063) );
AND3_X1 U880 ( .A1(n1181), .A2(n1024), .A3(n1013), .ZN(n1176) );
AND2_X1 U881 ( .A1(n1030), .A2(n1188), .ZN(n1181) );
NAND2_X1 U882 ( .A1(n1192), .A2(n1031), .ZN(n1188) );
NAND4_X1 U883 ( .A1(n1193), .A2(G953), .A3(n1194), .A4(n1195), .ZN(n1192) );
XNOR2_X1 U884 ( .A(KEYINPUT57), .B(n1151), .ZN(n1194) );
INV_X1 U885 ( .A(n1049), .ZN(n1193) );
XOR2_X1 U886 ( .A(G900), .B(KEYINPUT27), .Z(n1049) );
XNOR2_X1 U887 ( .A(G122), .B(n1160), .ZN(G24) );
NAND4_X1 U888 ( .A1(n1164), .A2(n1007), .A3(n1182), .A4(n1183), .ZN(n1160) );
NOR2_X1 U889 ( .A1(n1175), .A2(n1024), .ZN(n1007) );
XNOR2_X1 U890 ( .A(G119), .B(n1196), .ZN(G21) );
NAND4_X1 U891 ( .A1(n1197), .A2(n1000), .A3(n1163), .A4(n1030), .ZN(n1196) );
AND3_X1 U892 ( .A1(n1024), .A2(n1175), .A3(n999), .ZN(n1163) );
XOR2_X1 U893 ( .A(n1198), .B(KEYINPUT28), .Z(n1197) );
XOR2_X1 U894 ( .A(G116), .B(n1157), .Z(G18) );
AND3_X1 U895 ( .A1(n997), .A2(n1014), .A3(n1164), .ZN(n1157) );
XOR2_X1 U896 ( .A(G113), .B(n1156), .Z(G15) );
AND3_X1 U897 ( .A1(n997), .A2(n1013), .A3(n1164), .ZN(n1156) );
AND3_X1 U898 ( .A1(n1030), .A2(n1198), .A3(n1000), .ZN(n1164) );
AND2_X1 U899 ( .A1(n1199), .A2(n1019), .ZN(n1000) );
XOR2_X1 U900 ( .A(KEYINPUT14), .B(n1018), .Z(n1199) );
NOR2_X1 U901 ( .A1(n1182), .A2(n1033), .ZN(n1013) );
NOR2_X1 U902 ( .A1(n1024), .A2(n1023), .ZN(n997) );
XNOR2_X1 U903 ( .A(G110), .B(n1158), .ZN(G12) );
NAND4_X1 U904 ( .A1(n1023), .A2(n1159), .A3(n999), .A4(n1024), .ZN(n1158) );
XOR2_X1 U905 ( .A(n1200), .B(n1096), .Z(n1024) );
NAND2_X1 U906 ( .A1(G217), .A2(n1201), .ZN(n1096) );
NAND2_X1 U907 ( .A1(n1202), .A2(n1095), .ZN(n1200) );
XOR2_X1 U908 ( .A(n1203), .B(n1204), .Z(n1095) );
XNOR2_X1 U909 ( .A(n1205), .B(KEYINPUT0), .ZN(n1204) );
NAND2_X1 U910 ( .A1(KEYINPUT31), .A2(n1206), .ZN(n1205) );
XOR2_X1 U911 ( .A(n1207), .B(n1208), .Z(n1203) );
AND3_X1 U912 ( .A1(G221), .A2(n1002), .A3(G234), .ZN(n1208) );
NAND3_X1 U913 ( .A1(n1209), .A2(n1210), .A3(KEYINPUT18), .ZN(n1207) );
NAND2_X1 U914 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XNOR2_X1 U915 ( .A(n1213), .B(G119), .ZN(n1212) );
XNOR2_X1 U916 ( .A(n1214), .B(n1215), .ZN(n1211) );
XOR2_X1 U917 ( .A(KEYINPUT61), .B(KEYINPUT48), .Z(n1215) );
NAND2_X1 U918 ( .A1(n1216), .A2(n1214), .ZN(n1209) );
XNOR2_X1 U919 ( .A(n1217), .B(n1218), .ZN(n1214) );
XNOR2_X1 U920 ( .A(n1219), .B(n1138), .ZN(n1217) );
NAND2_X1 U921 ( .A1(KEYINPUT36), .A2(n1058), .ZN(n1219) );
XNOR2_X1 U922 ( .A(G119), .B(G128), .ZN(n1216) );
XNOR2_X1 U923 ( .A(G902), .B(KEYINPUT40), .ZN(n1202) );
NAND2_X1 U924 ( .A1(n1220), .A2(n1221), .ZN(n999) );
OR3_X1 U925 ( .A1(n1182), .A2(n1183), .A3(KEYINPUT9), .ZN(n1221) );
NAND2_X1 U926 ( .A1(KEYINPUT9), .A2(n1014), .ZN(n1220) );
AND2_X1 U927 ( .A1(n1033), .A2(n1182), .ZN(n1014) );
XNOR2_X1 U928 ( .A(n1037), .B(KEYINPUT16), .ZN(n1182) );
XOR2_X1 U929 ( .A(n1222), .B(n1101), .Z(n1037) );
INV_X1 U930 ( .A(G478), .ZN(n1101) );
NAND2_X1 U931 ( .A1(n1102), .A2(n1151), .ZN(n1222) );
XOR2_X1 U932 ( .A(n1223), .B(n1224), .Z(n1102) );
XNOR2_X1 U933 ( .A(n1225), .B(n1226), .ZN(n1224) );
XOR2_X1 U934 ( .A(KEYINPUT19), .B(G143), .Z(n1226) );
XNOR2_X1 U935 ( .A(G134), .B(G122), .ZN(n1225) );
XOR2_X1 U936 ( .A(n1227), .B(n1228), .Z(n1223) );
XOR2_X1 U937 ( .A(n1229), .B(n1230), .Z(n1228) );
AND3_X1 U938 ( .A1(n1231), .A2(G234), .A3(G217), .ZN(n1230) );
XNOR2_X1 U939 ( .A(KEYINPUT4), .B(G953), .ZN(n1231) );
NOR2_X1 U940 ( .A1(KEYINPUT15), .A2(n1232), .ZN(n1229) );
XNOR2_X1 U941 ( .A(G128), .B(KEYINPUT7), .ZN(n1232) );
XNOR2_X1 U942 ( .A(n1233), .B(n1234), .ZN(n1227) );
NOR2_X1 U943 ( .A1(G107), .A2(KEYINPUT17), .ZN(n1234) );
INV_X1 U944 ( .A(n1183), .ZN(n1033) );
XNOR2_X1 U945 ( .A(n1235), .B(G475), .ZN(n1183) );
NAND2_X1 U946 ( .A1(n1105), .A2(n1151), .ZN(n1235) );
XOR2_X1 U947 ( .A(n1236), .B(n1237), .Z(n1105) );
XOR2_X1 U948 ( .A(n1238), .B(n1239), .Z(n1237) );
XNOR2_X1 U949 ( .A(G131), .B(n1058), .ZN(n1239) );
INV_X1 U950 ( .A(G125), .ZN(n1058) );
NOR2_X1 U951 ( .A1(KEYINPUT26), .A2(n1240), .ZN(n1238) );
XOR2_X1 U952 ( .A(n1241), .B(n1242), .Z(n1240) );
NOR2_X1 U953 ( .A1(KEYINPUT56), .A2(n1243), .ZN(n1242) );
XNOR2_X1 U954 ( .A(KEYINPUT49), .B(n1244), .ZN(n1243) );
XNOR2_X1 U955 ( .A(G104), .B(G113), .ZN(n1241) );
XOR2_X1 U956 ( .A(n1245), .B(n1218), .Z(n1236) );
XNOR2_X1 U957 ( .A(G140), .B(n1246), .ZN(n1218) );
NAND2_X1 U958 ( .A1(n1247), .A2(n1248), .ZN(n1245) );
NAND4_X1 U959 ( .A1(G143), .A2(G214), .A3(n1249), .A4(n1002), .ZN(n1248) );
XOR2_X1 U960 ( .A(KEYINPUT22), .B(n1250), .Z(n1247) );
NOR2_X1 U961 ( .A1(n1251), .A2(G143), .ZN(n1250) );
AND3_X1 U962 ( .A1(G214), .A2(n1002), .A3(n1249), .ZN(n1251) );
AND3_X1 U963 ( .A1(n1174), .A2(n1198), .A3(n1030), .ZN(n1159) );
NOR2_X1 U964 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
INV_X1 U965 ( .A(n1189), .ZN(n1028) );
NAND2_X1 U966 ( .A1(G214), .A2(n1252), .ZN(n1189) );
XNOR2_X1 U967 ( .A(n1042), .B(n1040), .ZN(n1029) );
NAND2_X1 U968 ( .A1(G210), .A2(n1252), .ZN(n1040) );
NAND2_X1 U969 ( .A1(n1151), .A2(n1249), .ZN(n1252) );
NAND2_X1 U970 ( .A1(n1253), .A2(n1151), .ZN(n1042) );
XNOR2_X1 U971 ( .A(n1149), .B(n1146), .ZN(n1253) );
XOR2_X1 U972 ( .A(n1254), .B(n1255), .Z(n1146) );
INV_X1 U973 ( .A(n1086), .ZN(n1255) );
XNOR2_X1 U974 ( .A(n1256), .B(n1257), .ZN(n1086) );
XOR2_X1 U975 ( .A(G113), .B(n1258), .Z(n1257) );
XNOR2_X1 U976 ( .A(KEYINPUT43), .B(n1244), .ZN(n1258) );
INV_X1 U977 ( .A(G122), .ZN(n1244) );
XNOR2_X1 U978 ( .A(n1259), .B(n1138), .ZN(n1256) );
NAND2_X1 U979 ( .A1(KEYINPUT39), .A2(n1087), .ZN(n1254) );
XOR2_X1 U980 ( .A(n1260), .B(n1261), .Z(n1087) );
XNOR2_X1 U981 ( .A(KEYINPUT5), .B(n1262), .ZN(n1260) );
NOR2_X1 U982 ( .A1(KEYINPUT13), .A2(n1125), .ZN(n1262) );
XOR2_X1 U983 ( .A(n1263), .B(n1121), .Z(n1149) );
XNOR2_X1 U984 ( .A(G125), .B(n1264), .ZN(n1263) );
NOR2_X1 U985 ( .A1(G953), .A2(n1081), .ZN(n1264) );
INV_X1 U986 ( .A(G224), .ZN(n1081) );
NAND2_X1 U987 ( .A1(n1031), .A2(n1265), .ZN(n1198) );
NAND3_X1 U988 ( .A1(n1082), .A2(n1195), .A3(G902), .ZN(n1265) );
NOR2_X1 U989 ( .A1(n1002), .A2(G898), .ZN(n1082) );
NAND3_X1 U990 ( .A1(n1195), .A2(n1002), .A3(G952), .ZN(n1031) );
NAND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1195) );
NOR2_X1 U992 ( .A1(n1019), .A2(n1018), .ZN(n1174) );
AND2_X1 U993 ( .A1(G221), .A2(n1201), .ZN(n1018) );
NAND2_X1 U994 ( .A1(G234), .A2(n1151), .ZN(n1201) );
XNOR2_X1 U995 ( .A(n1038), .B(n1266), .ZN(n1019) );
NOR2_X1 U996 ( .A1(KEYINPUT63), .A2(n1039), .ZN(n1266) );
XOR2_X1 U997 ( .A(n1132), .B(KEYINPUT23), .Z(n1039) );
INV_X1 U998 ( .A(G469), .ZN(n1132) );
NAND2_X1 U999 ( .A1(n1267), .A2(n1151), .ZN(n1038) );
XOR2_X1 U1000 ( .A(n1268), .B(n1269), .Z(n1267) );
XNOR2_X1 U1001 ( .A(n1270), .B(n1129), .ZN(n1269) );
XNOR2_X1 U1002 ( .A(n1059), .B(n1271), .ZN(n1129) );
XNOR2_X1 U1003 ( .A(n1125), .B(n1261), .ZN(n1271) );
XNOR2_X1 U1004 ( .A(n1272), .B(G107), .ZN(n1261) );
INV_X1 U1005 ( .A(G104), .ZN(n1272) );
XOR2_X1 U1006 ( .A(n1273), .B(n1274), .Z(n1059) );
XNOR2_X1 U1007 ( .A(G143), .B(n1213), .ZN(n1274) );
INV_X1 U1008 ( .A(G128), .ZN(n1213) );
NAND2_X1 U1009 ( .A1(KEYINPUT11), .A2(n1246), .ZN(n1273) );
INV_X1 U1010 ( .A(G146), .ZN(n1246) );
NAND2_X1 U1011 ( .A1(KEYINPUT20), .A2(n1138), .ZN(n1270) );
INV_X1 U1012 ( .A(G110), .ZN(n1138) );
XOR2_X1 U1013 ( .A(n1275), .B(n1276), .Z(n1268) );
XNOR2_X1 U1014 ( .A(G140), .B(n1136), .ZN(n1276) );
AND2_X1 U1015 ( .A1(G227), .A2(n1002), .ZN(n1136) );
NAND2_X1 U1016 ( .A1(KEYINPUT35), .A2(n1060), .ZN(n1275) );
INV_X1 U1017 ( .A(n1175), .ZN(n1023) );
XOR2_X1 U1018 ( .A(n1277), .B(n1112), .Z(n1175) );
INV_X1 U1019 ( .A(G472), .ZN(n1112) );
NAND2_X1 U1020 ( .A1(n1278), .A2(n1151), .ZN(n1277) );
INV_X1 U1021 ( .A(G902), .ZN(n1151) );
XOR2_X1 U1022 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U1023 ( .A(n1060), .B(n1281), .Z(n1280) );
XNOR2_X1 U1024 ( .A(n1125), .B(n1124), .ZN(n1281) );
AND3_X1 U1025 ( .A1(n1249), .A2(n1002), .A3(G210), .ZN(n1124) );
INV_X1 U1026 ( .A(G953), .ZN(n1002) );
INV_X1 U1027 ( .A(G237), .ZN(n1249) );
INV_X1 U1028 ( .A(G101), .ZN(n1125) );
XOR2_X1 U1029 ( .A(G131), .B(n1282), .Z(n1060) );
XNOR2_X1 U1030 ( .A(n1206), .B(G134), .ZN(n1282) );
INV_X1 U1031 ( .A(G137), .ZN(n1206) );
XNOR2_X1 U1032 ( .A(n1119), .B(n1121), .ZN(n1279) );
XNOR2_X1 U1033 ( .A(n1283), .B(n1284), .ZN(n1121) );
NOR2_X1 U1034 ( .A1(KEYINPUT37), .A2(G143), .ZN(n1284) );
XNOR2_X1 U1035 ( .A(G146), .B(G128), .ZN(n1283) );
XNOR2_X1 U1036 ( .A(n1259), .B(n1285), .ZN(n1119) );
NOR2_X1 U1037 ( .A1(G113), .A2(KEYINPUT24), .ZN(n1285) );
XNOR2_X1 U1038 ( .A(G119), .B(n1233), .ZN(n1259) );
XOR2_X1 U1039 ( .A(G116), .B(KEYINPUT47), .Z(n1233) );
endmodule


