//Key = 1000011100011100111000110101100110110111111100000101001111011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268;

XNOR2_X1 U698 ( .A(G107), .B(n965), .ZN(G9) );
NAND4_X1 U699 ( .A1(n966), .A2(n967), .A3(n968), .A4(n969), .ZN(n965) );
XNOR2_X1 U700 ( .A(n970), .B(KEYINPUT12), .ZN(n966) );
NAND4_X1 U701 ( .A1(n971), .A2(n972), .A3(n973), .A4(n974), .ZN(G75) );
OR3_X1 U702 ( .A1(G953), .A2(KEYINPUT41), .A3(G952), .ZN(n974) );
NAND2_X1 U703 ( .A1(G952), .A2(n975), .ZN(n973) );
NAND4_X1 U704 ( .A1(n976), .A2(n977), .A3(n978), .A4(n979), .ZN(n975) );
NAND3_X1 U705 ( .A1(n980), .A2(n981), .A3(KEYINPUT39), .ZN(n978) );
NAND2_X1 U706 ( .A1(n982), .A2(n983), .ZN(n980) );
NAND4_X1 U707 ( .A1(n984), .A2(n985), .A3(n986), .A4(n987), .ZN(n983) );
NAND3_X1 U708 ( .A1(n988), .A2(n989), .A3(n990), .ZN(n987) );
NAND2_X1 U709 ( .A1(n991), .A2(n992), .ZN(n989) );
NAND2_X1 U710 ( .A1(n970), .A2(n993), .ZN(n988) );
INV_X1 U711 ( .A(KEYINPUT5), .ZN(n993) );
NAND4_X1 U712 ( .A1(n994), .A2(n995), .A3(n996), .A4(n969), .ZN(n986) );
NAND2_X1 U713 ( .A1(KEYINPUT5), .A2(n970), .ZN(n996) );
OR3_X1 U714 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n995) );
NAND2_X1 U715 ( .A1(n999), .A2(n991), .ZN(n994) );
XOR2_X1 U716 ( .A(KEYINPUT47), .B(KEYINPUT36), .Z(n999) );
NAND3_X1 U717 ( .A1(n969), .A2(n1000), .A3(n991), .ZN(n982) );
NAND2_X1 U718 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
NAND2_X1 U719 ( .A1(n985), .A2(n1003), .ZN(n1002) );
NAND2_X1 U720 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
OR2_X1 U721 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NAND2_X1 U722 ( .A1(n984), .A2(n1008), .ZN(n1001) );
NAND2_X1 U723 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
XOR2_X1 U724 ( .A(KEYINPUT38), .B(n967), .Z(n1009) );
NAND4_X1 U725 ( .A1(n1011), .A2(n985), .A3(n1012), .A4(n1013), .ZN(n972) );
NOR3_X1 U726 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NOR2_X1 U727 ( .A1(KEYINPUT59), .A2(n1017), .ZN(n1016) );
NOR2_X1 U728 ( .A1(n1018), .A2(n1019), .ZN(n1015) );
NAND3_X1 U729 ( .A1(n997), .A2(n1020), .A3(n1007), .ZN(n1014) );
NOR3_X1 U730 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1012) );
NOR2_X1 U731 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NOR2_X1 U732 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
XNOR2_X1 U733 ( .A(KEYINPUT9), .B(n1017), .ZN(n1027) );
INV_X1 U734 ( .A(KEYINPUT59), .ZN(n1026) );
AND3_X1 U735 ( .A1(n1024), .A2(n1017), .A3(KEYINPUT59), .ZN(n1022) );
XOR2_X1 U736 ( .A(KEYINPUT2), .B(n998), .Z(n1021) );
NAND2_X1 U737 ( .A1(KEYINPUT41), .A2(G953), .ZN(n971) );
NAND2_X1 U738 ( .A1(n1028), .A2(n1029), .ZN(G72) );
NAND2_X1 U739 ( .A1(n1030), .A2(n979), .ZN(n1029) );
XOR2_X1 U740 ( .A(n1031), .B(n1032), .Z(n1030) );
NAND2_X1 U741 ( .A1(KEYINPUT13), .A2(n1033), .ZN(n1032) );
NAND2_X1 U742 ( .A1(n1034), .A2(G953), .ZN(n1028) );
XOR2_X1 U743 ( .A(n1031), .B(n1035), .Z(n1034) );
NOR2_X1 U744 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U745 ( .A1(n1038), .A2(n1039), .ZN(n1031) );
NAND2_X1 U746 ( .A1(n1040), .A2(n1037), .ZN(n1039) );
XOR2_X1 U747 ( .A(n1041), .B(n1042), .Z(n1038) );
XNOR2_X1 U748 ( .A(n1043), .B(n1044), .ZN(n1041) );
NOR2_X1 U749 ( .A1(KEYINPUT46), .A2(n1045), .ZN(n1044) );
XOR2_X1 U750 ( .A(n1046), .B(n1047), .Z(G69) );
XOR2_X1 U751 ( .A(n1048), .B(n1049), .Z(n1047) );
NAND2_X1 U752 ( .A1(G953), .A2(n1050), .ZN(n1049) );
NAND2_X1 U753 ( .A1(G898), .A2(G224), .ZN(n1050) );
NAND2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1048) );
NAND2_X1 U755 ( .A1(n1040), .A2(n1053), .ZN(n1052) );
XOR2_X1 U756 ( .A(n1054), .B(n1055), .Z(n1051) );
NOR2_X1 U757 ( .A1(n976), .A2(G953), .ZN(n1046) );
NOR2_X1 U758 ( .A1(n1056), .A2(n1057), .ZN(G66) );
XNOR2_X1 U759 ( .A(n1058), .B(n1059), .ZN(n1057) );
NOR2_X1 U760 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U761 ( .A1(n1056), .A2(n1062), .ZN(G63) );
XNOR2_X1 U762 ( .A(n1063), .B(n1064), .ZN(n1062) );
AND2_X1 U763 ( .A1(G478), .A2(n1065), .ZN(n1063) );
NOR2_X1 U764 ( .A1(n1056), .A2(n1066), .ZN(G60) );
XNOR2_X1 U765 ( .A(n1067), .B(n1068), .ZN(n1066) );
NAND2_X1 U766 ( .A1(KEYINPUT31), .A2(n1069), .ZN(n1067) );
NAND2_X1 U767 ( .A1(n1065), .A2(G475), .ZN(n1069) );
XOR2_X1 U768 ( .A(G104), .B(n1070), .Z(G6) );
NOR2_X1 U769 ( .A1(n1056), .A2(n1071), .ZN(G57) );
XOR2_X1 U770 ( .A(n1072), .B(n1073), .Z(n1071) );
XOR2_X1 U771 ( .A(n1074), .B(n1075), .Z(n1072) );
NOR2_X1 U772 ( .A1(n1019), .A2(n1061), .ZN(n1075) );
NAND2_X1 U773 ( .A1(KEYINPUT7), .A2(n1076), .ZN(n1074) );
NOR2_X1 U774 ( .A1(n1056), .A2(n1077), .ZN(G54) );
XOR2_X1 U775 ( .A(n1078), .B(n1079), .Z(n1077) );
XOR2_X1 U776 ( .A(n1080), .B(n1081), .Z(n1079) );
XOR2_X1 U777 ( .A(n1082), .B(n1083), .Z(n1078) );
AND2_X1 U778 ( .A1(G469), .A2(n1065), .ZN(n1083) );
INV_X1 U779 ( .A(n1061), .ZN(n1065) );
XOR2_X1 U780 ( .A(n1084), .B(n1085), .Z(n1082) );
NOR2_X1 U781 ( .A1(KEYINPUT10), .A2(n1086), .ZN(n1085) );
XOR2_X1 U782 ( .A(n1087), .B(n1043), .Z(n1086) );
NAND2_X1 U783 ( .A1(KEYINPUT11), .A2(n1088), .ZN(n1087) );
NOR2_X1 U784 ( .A1(n1056), .A2(n1089), .ZN(G51) );
NOR2_X1 U785 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U786 ( .A(n1092), .B(KEYINPUT54), .Z(n1091) );
NAND2_X1 U787 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U788 ( .A(KEYINPUT16), .B(n1095), .Z(n1094) );
NOR2_X1 U789 ( .A1(n1096), .A2(n1061), .ZN(n1095) );
NOR3_X1 U790 ( .A1(n1061), .A2(n1093), .A3(n1096), .ZN(n1090) );
INV_X1 U791 ( .A(G210), .ZN(n1096) );
AND2_X1 U792 ( .A1(n1097), .A2(n1098), .ZN(n1093) );
NAND2_X1 U793 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U794 ( .A(KEYINPUT55), .B(n1101), .Z(n1099) );
NAND2_X1 U795 ( .A1(n1101), .A2(n1102), .ZN(n1097) );
INV_X1 U796 ( .A(n1100), .ZN(n1102) );
XNOR2_X1 U797 ( .A(n1103), .B(n1104), .ZN(n1101) );
XOR2_X1 U798 ( .A(G125), .B(n1105), .Z(n1104) );
NOR2_X1 U799 ( .A1(KEYINPUT45), .A2(n1106), .ZN(n1105) );
XOR2_X1 U800 ( .A(KEYINPUT57), .B(n1107), .Z(n1106) );
NAND2_X1 U801 ( .A1(G902), .A2(n1108), .ZN(n1061) );
NAND2_X1 U802 ( .A1(n976), .A2(n977), .ZN(n1108) );
INV_X1 U803 ( .A(n1033), .ZN(n977) );
NAND4_X1 U804 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1033) );
NOR4_X1 U805 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1112) );
INV_X1 U806 ( .A(n1117), .ZN(n1116) );
NOR3_X1 U807 ( .A1(n984), .A2(n1118), .A3(n1119), .ZN(n1114) );
INV_X1 U808 ( .A(KEYINPUT30), .ZN(n1119) );
NOR2_X1 U809 ( .A1(n1120), .A2(n1121), .ZN(n1113) );
NOR2_X1 U810 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
NOR2_X1 U811 ( .A1(KEYINPUT30), .A2(n1118), .ZN(n1122) );
NOR2_X1 U812 ( .A1(n1124), .A2(n1125), .ZN(n1111) );
INV_X1 U813 ( .A(n1126), .ZN(n1125) );
AND2_X1 U814 ( .A1(n1127), .A2(n1128), .ZN(n976) );
AND4_X1 U815 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1128) );
NOR4_X1 U816 ( .A1(n1133), .A2(n1070), .A3(n1134), .A4(n1135), .ZN(n1127) );
NOR3_X1 U817 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
INV_X1 U818 ( .A(n967), .ZN(n1137) );
XOR2_X1 U819 ( .A(KEYINPUT60), .B(n969), .Z(n1136) );
INV_X1 U820 ( .A(n990), .ZN(n969) );
NOR3_X1 U821 ( .A1(n1138), .A2(n990), .A3(n1010), .ZN(n1070) );
AND2_X1 U822 ( .A1(n1139), .A2(G953), .ZN(n1056) );
XNOR2_X1 U823 ( .A(G952), .B(KEYINPUT29), .ZN(n1139) );
XOR2_X1 U824 ( .A(n1140), .B(n1117), .Z(G48) );
NAND2_X1 U825 ( .A1(n1141), .A2(n1142), .ZN(n1117) );
XOR2_X1 U826 ( .A(G143), .B(n1115), .Z(G45) );
AND3_X1 U827 ( .A1(n1011), .A2(n1143), .A3(n1144), .ZN(n1115) );
NOR3_X1 U828 ( .A1(n1004), .A2(n1145), .A3(n1146), .ZN(n1144) );
XOR2_X1 U829 ( .A(n1147), .B(n1148), .Z(G42) );
NOR2_X1 U830 ( .A1(KEYINPUT33), .A2(n1149), .ZN(n1148) );
NOR2_X1 U831 ( .A1(n1121), .A2(n1118), .ZN(n1149) );
NAND2_X1 U832 ( .A1(n1150), .A2(n970), .ZN(n1118) );
XOR2_X1 U833 ( .A(n1084), .B(KEYINPUT3), .Z(n1147) );
XOR2_X1 U834 ( .A(G137), .B(n1151), .Z(G39) );
NOR3_X1 U835 ( .A1(n1121), .A2(KEYINPUT1), .A3(n1152), .ZN(n1151) );
XNOR2_X1 U836 ( .A(n1123), .B(KEYINPUT44), .ZN(n1152) );
AND3_X1 U837 ( .A1(n985), .A2(n1153), .A3(n1143), .ZN(n1123) );
XOR2_X1 U838 ( .A(n1124), .B(n1154), .Z(G36) );
NOR2_X1 U839 ( .A1(KEYINPUT50), .A2(n1155), .ZN(n1154) );
INV_X1 U840 ( .A(G134), .ZN(n1155) );
AND4_X1 U841 ( .A1(n1143), .A2(n984), .A3(n1011), .A4(n967), .ZN(n1124) );
XOR2_X1 U842 ( .A(n1156), .B(n1109), .Z(G33) );
NAND4_X1 U843 ( .A1(n1143), .A2(n984), .A3(n1011), .A4(n1142), .ZN(n1109) );
INV_X1 U844 ( .A(n1121), .ZN(n984) );
NAND2_X1 U845 ( .A1(n1157), .A2(n1007), .ZN(n1121) );
INV_X1 U846 ( .A(n1006), .ZN(n1157) );
XOR2_X1 U847 ( .A(n1158), .B(n1110), .Z(G30) );
NAND2_X1 U848 ( .A1(n1141), .A2(n967), .ZN(n1110) );
AND3_X1 U849 ( .A1(n1159), .A2(n1153), .A3(n1143), .ZN(n1141) );
AND3_X1 U850 ( .A1(n1160), .A2(n1161), .A3(n970), .ZN(n1143) );
XOR2_X1 U851 ( .A(G101), .B(n1134), .Z(G3) );
AND4_X1 U852 ( .A1(n1162), .A2(n985), .A3(n1011), .A4(n1161), .ZN(n1134) );
XOR2_X1 U853 ( .A(n1163), .B(n1126), .Z(G27) );
NAND3_X1 U854 ( .A1(n991), .A2(n1159), .A3(n1150), .ZN(n1126) );
AND4_X1 U855 ( .A1(n1142), .A2(n1164), .A3(n1153), .A4(n1160), .ZN(n1150) );
NAND2_X1 U856 ( .A1(n1165), .A2(n1166), .ZN(n1160) );
NAND2_X1 U857 ( .A1(n1167), .A2(n1037), .ZN(n1166) );
INV_X1 U858 ( .A(G900), .ZN(n1037) );
XOR2_X1 U859 ( .A(n1168), .B(n1169), .Z(G24) );
NOR2_X1 U860 ( .A1(n1133), .A2(KEYINPUT53), .ZN(n1169) );
AND3_X1 U861 ( .A1(n991), .A2(n968), .A3(n1170), .ZN(n1133) );
NOR3_X1 U862 ( .A1(n990), .A2(n1145), .A3(n1146), .ZN(n1170) );
XNOR2_X1 U863 ( .A(n1171), .B(KEYINPUT63), .ZN(n1146) );
NAND2_X1 U864 ( .A1(n1164), .A2(n1011), .ZN(n990) );
XOR2_X1 U865 ( .A(n1172), .B(n1173), .Z(G21) );
XOR2_X1 U866 ( .A(KEYINPUT23), .B(G119), .Z(n1173) );
NOR2_X1 U867 ( .A1(n1174), .A2(n1175), .ZN(n1172) );
NOR2_X1 U868 ( .A1(n1176), .A2(n1132), .ZN(n1175) );
NAND3_X1 U869 ( .A1(n985), .A2(n1153), .A3(n1177), .ZN(n1132) );
INV_X1 U870 ( .A(KEYINPUT42), .ZN(n1176) );
NOR4_X1 U871 ( .A1(KEYINPUT42), .A2(n1178), .A3(n1179), .A4(n992), .ZN(n1174) );
NAND2_X1 U872 ( .A1(n1153), .A2(n1161), .ZN(n992) );
NAND3_X1 U873 ( .A1(n1004), .A2(n1180), .A3(n985), .ZN(n1178) );
XOR2_X1 U874 ( .A(n1181), .B(n1131), .Z(G18) );
NAND3_X1 U875 ( .A1(n1011), .A2(n967), .A3(n1177), .ZN(n1131) );
NOR2_X1 U876 ( .A1(n1171), .A2(n1145), .ZN(n967) );
XNOR2_X1 U877 ( .A(G113), .B(n1130), .ZN(G15) );
NAND3_X1 U878 ( .A1(n1011), .A2(n1142), .A3(n1177), .ZN(n1130) );
AND3_X1 U879 ( .A1(n968), .A2(n1161), .A3(n991), .ZN(n1177) );
INV_X1 U880 ( .A(n1179), .ZN(n991) );
NAND2_X1 U881 ( .A1(n1182), .A2(n997), .ZN(n1179) );
INV_X1 U882 ( .A(n1010), .ZN(n1142) );
NAND2_X1 U883 ( .A1(n1145), .A2(n1171), .ZN(n1010) );
NAND2_X1 U884 ( .A1(n1183), .A2(n1184), .ZN(G12) );
NAND2_X1 U885 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U886 ( .A(n1187), .B(KEYINPUT62), .Z(n1183) );
OR2_X1 U887 ( .A1(n1186), .A2(n1185), .ZN(n1187) );
INV_X1 U888 ( .A(n1129), .ZN(n1185) );
NAND4_X1 U889 ( .A1(n1162), .A2(n985), .A3(n1164), .A4(n1153), .ZN(n1129) );
INV_X1 U890 ( .A(n1011), .ZN(n1153) );
XNOR2_X1 U891 ( .A(n1188), .B(n1060), .ZN(n1011) );
NAND2_X1 U892 ( .A1(G217), .A2(n1189), .ZN(n1060) );
NAND2_X1 U893 ( .A1(n1059), .A2(n1190), .ZN(n1188) );
XOR2_X1 U894 ( .A(n1191), .B(n1192), .Z(n1059) );
XOR2_X1 U895 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U896 ( .A(G137), .B(G119), .Z(n1194) );
XOR2_X1 U897 ( .A(KEYINPUT25), .B(KEYINPUT24), .Z(n1193) );
XOR2_X1 U898 ( .A(n1195), .B(n1196), .Z(n1191) );
XNOR2_X1 U899 ( .A(n1197), .B(n1198), .ZN(n1196) );
NAND2_X1 U900 ( .A1(G221), .A2(n1199), .ZN(n1197) );
XOR2_X1 U901 ( .A(n1200), .B(G110), .Z(n1195) );
NAND2_X1 U902 ( .A1(KEYINPUT40), .A2(n1042), .ZN(n1200) );
INV_X1 U903 ( .A(n1161), .ZN(n1164) );
NAND2_X1 U904 ( .A1(n1201), .A2(n1020), .ZN(n1161) );
NAND2_X1 U905 ( .A1(n1018), .A2(n1019), .ZN(n1020) );
NAND2_X1 U906 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XNOR2_X1 U907 ( .A(n1018), .B(KEYINPUT21), .ZN(n1203) );
AND2_X1 U908 ( .A1(n1204), .A2(n1190), .ZN(n1018) );
XNOR2_X1 U909 ( .A(n1073), .B(n1205), .ZN(n1204) );
XOR2_X1 U910 ( .A(KEYINPUT32), .B(n1076), .Z(n1205) );
XNOR2_X1 U911 ( .A(n1206), .B(n1207), .ZN(n1076) );
NOR2_X1 U912 ( .A1(KEYINPUT58), .A2(n1208), .ZN(n1207) );
XNOR2_X1 U913 ( .A(G113), .B(KEYINPUT20), .ZN(n1206) );
XNOR2_X1 U914 ( .A(n1209), .B(n1210), .ZN(n1073) );
XNOR2_X1 U915 ( .A(G101), .B(n1211), .ZN(n1210) );
NAND2_X1 U916 ( .A1(G210), .A2(n1212), .ZN(n1211) );
XOR2_X1 U917 ( .A(n1080), .B(n1107), .Z(n1209) );
XOR2_X1 U918 ( .A(n1019), .B(KEYINPUT35), .Z(n1202) );
INV_X1 U919 ( .A(G472), .ZN(n1019) );
NOR2_X1 U920 ( .A1(n1213), .A2(n1171), .ZN(n985) );
XNOR2_X1 U921 ( .A(n1214), .B(G475), .ZN(n1171) );
NAND2_X1 U922 ( .A1(n1190), .A2(n1068), .ZN(n1214) );
NAND2_X1 U923 ( .A1(n1215), .A2(n1216), .ZN(n1068) );
NAND2_X1 U924 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XOR2_X1 U925 ( .A(n1219), .B(KEYINPUT4), .Z(n1215) );
OR2_X1 U926 ( .A1(n1218), .A2(n1217), .ZN(n1219) );
XNOR2_X1 U927 ( .A(n1220), .B(n1221), .ZN(n1217) );
XOR2_X1 U928 ( .A(G131), .B(n1222), .Z(n1221) );
NOR2_X1 U929 ( .A1(KEYINPUT48), .A2(n1223), .ZN(n1222) );
XNOR2_X1 U930 ( .A(n1224), .B(n1042), .ZN(n1223) );
XOR2_X1 U931 ( .A(n1163), .B(n1084), .Z(n1042) );
NAND2_X1 U932 ( .A1(KEYINPUT28), .A2(n1140), .ZN(n1224) );
INV_X1 U933 ( .A(G146), .ZN(n1140) );
NAND2_X1 U934 ( .A1(KEYINPUT34), .A2(n1225), .ZN(n1220) );
XNOR2_X1 U935 ( .A(n1226), .B(n1227), .ZN(n1225) );
NAND2_X1 U936 ( .A1(G214), .A2(n1212), .ZN(n1226) );
NOR2_X1 U937 ( .A1(G953), .A2(G237), .ZN(n1212) );
XOR2_X1 U938 ( .A(G104), .B(n1228), .Z(n1218) );
XOR2_X1 U939 ( .A(G122), .B(G113), .Z(n1228) );
INV_X1 U940 ( .A(n1145), .ZN(n1213) );
XOR2_X1 U941 ( .A(n1229), .B(G478), .Z(n1145) );
NAND2_X1 U942 ( .A1(n1064), .A2(n1190), .ZN(n1229) );
XOR2_X1 U943 ( .A(n1230), .B(n1231), .Z(n1064) );
XOR2_X1 U944 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U945 ( .A(G128), .B(G107), .Z(n1233) );
XOR2_X1 U946 ( .A(KEYINPUT52), .B(G134), .Z(n1232) );
XOR2_X1 U947 ( .A(n1234), .B(n1227), .Z(n1230) );
XOR2_X1 U948 ( .A(n1235), .B(n1236), .Z(n1234) );
AND2_X1 U949 ( .A1(n1199), .A2(G217), .ZN(n1236) );
AND2_X1 U950 ( .A1(G234), .A2(n979), .ZN(n1199) );
NAND3_X1 U951 ( .A1(n1237), .A2(n1238), .A3(KEYINPUT27), .ZN(n1235) );
NAND2_X1 U952 ( .A1(KEYINPUT6), .A2(n1239), .ZN(n1238) );
XOR2_X1 U953 ( .A(n1181), .B(G122), .Z(n1239) );
INV_X1 U954 ( .A(G116), .ZN(n1181) );
OR3_X1 U955 ( .A1(n1168), .A2(G116), .A3(KEYINPUT6), .ZN(n1237) );
INV_X1 U956 ( .A(G122), .ZN(n1168) );
INV_X1 U957 ( .A(n1138), .ZN(n1162) );
NAND2_X1 U958 ( .A1(n968), .A2(n970), .ZN(n1138) );
AND2_X1 U959 ( .A1(n998), .A2(n997), .ZN(n970) );
NAND2_X1 U960 ( .A1(G221), .A2(n1189), .ZN(n997) );
NAND2_X1 U961 ( .A1(G234), .A2(n1240), .ZN(n1189) );
INV_X1 U962 ( .A(n1182), .ZN(n998) );
XOR2_X1 U963 ( .A(n1241), .B(G469), .Z(n1182) );
NAND2_X1 U964 ( .A1(n1242), .A2(n1190), .ZN(n1241) );
XOR2_X1 U965 ( .A(n1243), .B(n1081), .Z(n1242) );
XOR2_X1 U966 ( .A(G110), .B(n1244), .Z(n1081) );
NOR2_X1 U967 ( .A1(G953), .A2(n1036), .ZN(n1244) );
INV_X1 U968 ( .A(G227), .ZN(n1036) );
XNOR2_X1 U969 ( .A(n1245), .B(n1246), .ZN(n1243) );
NAND2_X1 U970 ( .A1(KEYINPUT56), .A2(n1084), .ZN(n1246) );
INV_X1 U971 ( .A(G140), .ZN(n1084) );
NAND2_X1 U972 ( .A1(KEYINPUT51), .A2(n1247), .ZN(n1245) );
XOR2_X1 U973 ( .A(n1248), .B(n1249), .Z(n1247) );
INV_X1 U974 ( .A(n1080), .ZN(n1249) );
XNOR2_X1 U975 ( .A(n1045), .B(KEYINPUT49), .ZN(n1080) );
XNOR2_X1 U976 ( .A(n1156), .B(n1250), .ZN(n1045) );
XOR2_X1 U977 ( .A(G137), .B(G134), .Z(n1250) );
INV_X1 U978 ( .A(G131), .ZN(n1156) );
NOR2_X1 U979 ( .A1(KEYINPUT26), .A2(n1251), .ZN(n1248) );
XOR2_X1 U980 ( .A(n1043), .B(n1088), .Z(n1251) );
XNOR2_X1 U981 ( .A(n1252), .B(n1198), .ZN(n1043) );
NAND2_X1 U982 ( .A1(n1253), .A2(KEYINPUT37), .ZN(n1252) );
XNOR2_X1 U983 ( .A(n1227), .B(KEYINPUT18), .ZN(n1253) );
AND2_X1 U984 ( .A1(n1159), .A2(n1180), .ZN(n968) );
NAND2_X1 U985 ( .A1(n1254), .A2(n1255), .ZN(n1180) );
NAND2_X1 U986 ( .A1(n1167), .A2(n1053), .ZN(n1255) );
INV_X1 U987 ( .A(G898), .ZN(n1053) );
AND3_X1 U988 ( .A1(n1040), .A2(n981), .A3(G902), .ZN(n1167) );
XOR2_X1 U989 ( .A(G953), .B(KEYINPUT14), .Z(n1040) );
XNOR2_X1 U990 ( .A(KEYINPUT43), .B(n1165), .ZN(n1254) );
NAND3_X1 U991 ( .A1(n981), .A2(n979), .A3(G952), .ZN(n1165) );
NAND2_X1 U992 ( .A1(G237), .A2(G234), .ZN(n981) );
INV_X1 U993 ( .A(n1004), .ZN(n1159) );
NAND2_X1 U994 ( .A1(n1256), .A2(n1006), .ZN(n1004) );
XNOR2_X1 U995 ( .A(n1017), .B(n1024), .ZN(n1006) );
AND2_X1 U996 ( .A1(n1257), .A2(n1258), .ZN(n1024) );
XOR2_X1 U997 ( .A(KEYINPUT19), .B(G210), .Z(n1257) );
NAND3_X1 U998 ( .A1(n1259), .A2(n1260), .A3(n1190), .ZN(n1017) );
XOR2_X1 U999 ( .A(G902), .B(KEYINPUT22), .Z(n1190) );
NAND2_X1 U1000 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XNOR2_X1 U1001 ( .A(n1263), .B(KEYINPUT15), .ZN(n1262) );
XOR2_X1 U1002 ( .A(n1163), .B(n1107), .Z(n1261) );
INV_X1 U1003 ( .A(G125), .ZN(n1163) );
NAND2_X1 U1004 ( .A1(n1264), .A2(n1263), .ZN(n1259) );
XOR2_X1 U1005 ( .A(n1100), .B(n1103), .Z(n1263) );
NAND2_X1 U1006 ( .A1(G224), .A2(n979), .ZN(n1103) );
INV_X1 U1007 ( .A(G953), .ZN(n979) );
XOR2_X1 U1008 ( .A(n1054), .B(n1265), .Z(n1100) );
NOR2_X1 U1009 ( .A1(KEYINPUT61), .A2(n1055), .ZN(n1265) );
XNOR2_X1 U1010 ( .A(G113), .B(n1208), .ZN(n1055) );
XNOR2_X1 U1011 ( .A(G119), .B(G116), .ZN(n1208) );
XOR2_X1 U1012 ( .A(n1088), .B(n1266), .Z(n1054) );
XOR2_X1 U1013 ( .A(G122), .B(G110), .Z(n1266) );
XNOR2_X1 U1014 ( .A(G101), .B(n1267), .ZN(n1088) );
XOR2_X1 U1015 ( .A(G107), .B(G104), .Z(n1267) );
XOR2_X1 U1016 ( .A(G125), .B(n1107), .Z(n1264) );
XOR2_X1 U1017 ( .A(n1198), .B(n1227), .Z(n1107) );
XOR2_X1 U1018 ( .A(G143), .B(KEYINPUT0), .Z(n1227) );
XNOR2_X1 U1019 ( .A(n1158), .B(G146), .ZN(n1198) );
INV_X1 U1020 ( .A(G128), .ZN(n1158) );
XOR2_X1 U1021 ( .A(n1007), .B(KEYINPUT8), .Z(n1256) );
NAND2_X1 U1022 ( .A1(G214), .A2(n1258), .ZN(n1007) );
NAND2_X1 U1023 ( .A1(n1268), .A2(n1240), .ZN(n1258) );
INV_X1 U1024 ( .A(G902), .ZN(n1240) );
INV_X1 U1025 ( .A(G237), .ZN(n1268) );
XOR2_X1 U1026 ( .A(G110), .B(KEYINPUT17), .Z(n1186) );
endmodule


