//Key = 0000111010010110101011010100000001001100100000000100000100101101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398;

XNOR2_X1 U747 ( .A(G107), .B(n1047), .ZN(G9) );
NOR2_X1 U748 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR4_X1 U749 ( .A1(n1050), .A2(n1051), .A3(G953), .A4(n1052), .ZN(n1049) );
NOR4_X1 U750 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1051) );
INV_X1 U751 ( .A(n1057), .ZN(n1054) );
NOR3_X1 U752 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1053) );
NOR3_X1 U753 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NOR3_X1 U754 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1058) );
NAND3_X1 U755 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1050) );
NAND2_X1 U756 ( .A1(n1062), .A2(n1070), .ZN(n1068) );
NAND2_X1 U757 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U758 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U759 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND3_X1 U760 ( .A1(n1057), .A2(n1077), .A3(n1078), .ZN(n1076) );
NAND2_X1 U761 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NAND2_X1 U762 ( .A1(n1081), .A2(n1082), .ZN(n1075) );
NAND2_X1 U763 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U764 ( .A1(n1057), .A2(n1085), .ZN(n1084) );
NAND2_X1 U765 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U766 ( .A1(n1088), .A2(n1061), .ZN(n1087) );
INV_X1 U767 ( .A(KEYINPUT28), .ZN(n1061) );
NAND2_X1 U768 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NAND2_X1 U769 ( .A1(n1078), .A2(n1091), .ZN(n1083) );
NAND2_X1 U770 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U771 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
INV_X1 U772 ( .A(KEYINPUT30), .ZN(n1095) );
NAND2_X1 U773 ( .A1(KEYINPUT30), .A2(n1096), .ZN(n1071) );
NAND4_X1 U774 ( .A1(n1073), .A2(n1094), .A3(n1081), .A4(n1078), .ZN(n1096) );
INV_X1 U775 ( .A(n1056), .ZN(n1073) );
NOR3_X1 U776 ( .A1(n1052), .A2(G953), .A3(G952), .ZN(n1048) );
AND4_X1 U777 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1052) );
NOR4_X1 U778 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1100) );
XOR2_X1 U779 ( .A(KEYINPUT9), .B(n1105), .Z(n1104) );
XOR2_X1 U780 ( .A(KEYINPUT22), .B(n1106), .Z(n1103) );
NOR2_X1 U781 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U782 ( .A1(G478), .A2(n1109), .ZN(n1108) );
XNOR2_X1 U783 ( .A(n1110), .B(KEYINPUT6), .ZN(n1109) );
NOR3_X1 U784 ( .A1(n1111), .A2(n1112), .A3(n1089), .ZN(n1099) );
NOR2_X1 U785 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR2_X1 U786 ( .A1(G902), .A2(n1115), .ZN(n1113) );
XNOR2_X1 U787 ( .A(KEYINPUT60), .B(n1116), .ZN(n1098) );
XOR2_X1 U788 ( .A(n1117), .B(n1118), .Z(G72) );
XOR2_X1 U789 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U790 ( .A1(G953), .A2(n1121), .ZN(n1120) );
NAND2_X1 U791 ( .A1(G900), .A2(G227), .ZN(n1121) );
NAND2_X1 U792 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
XOR2_X1 U793 ( .A(KEYINPUT33), .B(n1124), .Z(n1123) );
NOR2_X1 U794 ( .A1(G900), .A2(n1125), .ZN(n1124) );
XNOR2_X1 U795 ( .A(n1126), .B(n1127), .ZN(n1122) );
NOR2_X1 U796 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U797 ( .A(n1130), .B(KEYINPUT8), .Z(n1129) );
NAND2_X1 U798 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR2_X1 U799 ( .A1(n1131), .A2(n1132), .ZN(n1128) );
XNOR2_X1 U800 ( .A(KEYINPUT62), .B(n1133), .ZN(n1131) );
NOR2_X1 U801 ( .A1(n1067), .A2(G953), .ZN(n1117) );
XOR2_X1 U802 ( .A(n1134), .B(n1135), .Z(G69) );
NOR2_X1 U803 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XOR2_X1 U804 ( .A(n1138), .B(KEYINPUT37), .Z(n1137) );
NAND3_X1 U805 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1138) );
NAND2_X1 U806 ( .A1(KEYINPUT55), .A2(n1142), .ZN(n1140) );
NAND2_X1 U807 ( .A1(G953), .A2(n1143), .ZN(n1139) );
NOR3_X1 U808 ( .A1(n1069), .A2(n1144), .A3(n1145), .ZN(n1136) );
NOR2_X1 U809 ( .A1(G953), .A2(n1146), .ZN(n1145) );
NOR2_X1 U810 ( .A1(n1141), .A2(n1147), .ZN(n1146) );
NOR2_X1 U811 ( .A1(n1125), .A2(n1147), .ZN(n1144) );
INV_X1 U812 ( .A(KEYINPUT55), .ZN(n1147) );
NAND2_X1 U813 ( .A1(G953), .A2(n1148), .ZN(n1134) );
NAND2_X1 U814 ( .A1(G898), .A2(G224), .ZN(n1148) );
NOR2_X1 U815 ( .A1(n1149), .A2(n1150), .ZN(G66) );
XOR2_X1 U816 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U817 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
NOR2_X1 U818 ( .A1(n1149), .A2(n1155), .ZN(G63) );
NOR3_X1 U819 ( .A1(n1110), .A2(n1156), .A3(n1157), .ZN(n1155) );
NOR3_X1 U820 ( .A1(n1158), .A2(n1159), .A3(n1154), .ZN(n1157) );
NOR2_X1 U821 ( .A1(n1160), .A2(n1161), .ZN(n1156) );
NOR2_X1 U822 ( .A1(n1162), .A2(n1159), .ZN(n1160) );
NOR2_X1 U823 ( .A1(n1163), .A2(n1142), .ZN(n1162) );
NOR2_X1 U824 ( .A1(n1149), .A2(n1164), .ZN(G60) );
XNOR2_X1 U825 ( .A(n1165), .B(n1166), .ZN(n1164) );
AND2_X1 U826 ( .A1(G475), .A2(n1167), .ZN(n1166) );
XOR2_X1 U827 ( .A(n1168), .B(G104), .Z(G6) );
NAND2_X1 U828 ( .A1(KEYINPUT23), .A2(n1169), .ZN(n1168) );
NOR2_X1 U829 ( .A1(n1149), .A2(n1170), .ZN(G57) );
XOR2_X1 U830 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U831 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U832 ( .A1(KEYINPUT45), .A2(n1175), .ZN(n1174) );
AND2_X1 U833 ( .A1(G472), .A2(n1167), .ZN(n1173) );
XNOR2_X1 U834 ( .A(G101), .B(n1176), .ZN(n1171) );
NOR2_X1 U835 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XOR2_X1 U836 ( .A(n1179), .B(KEYINPUT49), .Z(n1178) );
NAND2_X1 U837 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NOR2_X1 U838 ( .A1(n1180), .A2(n1181), .ZN(n1177) );
NAND3_X1 U839 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1181) );
OR2_X1 U840 ( .A1(n1133), .A2(KEYINPUT63), .ZN(n1184) );
NAND3_X1 U841 ( .A1(KEYINPUT63), .A2(n1133), .A3(n1185), .ZN(n1183) );
NAND2_X1 U842 ( .A1(n1186), .A2(n1187), .ZN(n1182) );
NAND2_X1 U843 ( .A1(KEYINPUT63), .A2(n1188), .ZN(n1187) );
XNOR2_X1 U844 ( .A(KEYINPUT42), .B(n1189), .ZN(n1188) );
INV_X1 U845 ( .A(n1133), .ZN(n1189) );
NOR3_X1 U846 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(G54) );
AND3_X1 U847 ( .A1(KEYINPUT57), .A2(G953), .A3(G952), .ZN(n1192) );
NOR2_X1 U848 ( .A1(KEYINPUT57), .A2(n1193), .ZN(n1191) );
INV_X1 U849 ( .A(n1149), .ZN(n1193) );
XOR2_X1 U850 ( .A(n1194), .B(n1195), .Z(n1190) );
XNOR2_X1 U851 ( .A(n1196), .B(n1133), .ZN(n1195) );
NAND2_X1 U852 ( .A1(KEYINPUT21), .A2(n1197), .ZN(n1196) );
NAND2_X1 U853 ( .A1(n1167), .A2(G469), .ZN(n1197) );
INV_X1 U854 ( .A(n1154), .ZN(n1167) );
XOR2_X1 U855 ( .A(n1198), .B(n1199), .Z(n1194) );
XNOR2_X1 U856 ( .A(n1200), .B(n1201), .ZN(n1199) );
NOR2_X1 U857 ( .A1(KEYINPUT56), .A2(n1202), .ZN(n1200) );
XOR2_X1 U858 ( .A(n1203), .B(n1204), .Z(n1202) );
NOR2_X1 U859 ( .A1(n1205), .A2(n1206), .ZN(n1198) );
XOR2_X1 U860 ( .A(KEYINPUT17), .B(n1207), .Z(n1206) );
AND2_X1 U861 ( .A1(G140), .A2(n1208), .ZN(n1207) );
NOR2_X1 U862 ( .A1(G140), .A2(n1208), .ZN(n1205) );
NOR2_X1 U863 ( .A1(n1149), .A2(n1209), .ZN(G51) );
XOR2_X1 U864 ( .A(n1210), .B(n1115), .Z(n1209) );
NOR2_X1 U865 ( .A1(n1114), .A2(n1154), .ZN(n1210) );
NAND2_X1 U866 ( .A1(G902), .A2(n1211), .ZN(n1154) );
NAND2_X1 U867 ( .A1(n1069), .A2(n1067), .ZN(n1211) );
INV_X1 U868 ( .A(n1163), .ZN(n1067) );
NAND4_X1 U869 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1163) );
AND4_X1 U870 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1215) );
INV_X1 U871 ( .A(n1220), .ZN(n1218) );
OR3_X1 U872 ( .A1(n1221), .A2(n1222), .A3(n1079), .ZN(n1216) );
XNOR2_X1 U873 ( .A(n1223), .B(KEYINPUT29), .ZN(n1222) );
NOR3_X1 U874 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1214) );
NOR2_X1 U875 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NAND4_X1 U876 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1228) );
INV_X1 U877 ( .A(KEYINPUT1), .ZN(n1227) );
NOR2_X1 U878 ( .A1(KEYINPUT1), .A2(n1233), .ZN(n1225) );
NOR2_X1 U879 ( .A1(n1234), .A2(n1235), .ZN(n1224) );
XOR2_X1 U880 ( .A(n1236), .B(KEYINPUT53), .Z(n1234) );
NAND2_X1 U881 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XNOR2_X1 U882 ( .A(KEYINPUT47), .B(n1055), .ZN(n1238) );
INV_X1 U883 ( .A(n1221), .ZN(n1237) );
INV_X1 U884 ( .A(n1142), .ZN(n1069) );
NAND4_X1 U885 ( .A1(n1169), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1142) );
AND4_X1 U886 ( .A1(n1047), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1241) );
NAND3_X1 U887 ( .A1(n1057), .A2(n1245), .A3(n1246), .ZN(n1047) );
NAND2_X1 U888 ( .A1(n1081), .A2(n1247), .ZN(n1240) );
NAND2_X1 U889 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND3_X1 U890 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1249) );
OR2_X1 U891 ( .A1(n1253), .A2(n1245), .ZN(n1251) );
NAND2_X1 U892 ( .A1(n1254), .A2(n1253), .ZN(n1250) );
INV_X1 U893 ( .A(KEYINPUT5), .ZN(n1253) );
NAND3_X1 U894 ( .A1(n1255), .A2(n1256), .A3(n1088), .ZN(n1254) );
NAND2_X1 U895 ( .A1(n1094), .A2(n1245), .ZN(n1248) );
OR2_X1 U896 ( .A1(n1257), .A2(n1258), .ZN(n1239) );
NAND3_X1 U897 ( .A1(n1057), .A2(n1245), .A3(n1259), .ZN(n1169) );
NOR2_X1 U898 ( .A1(n1125), .A2(G952), .ZN(n1149) );
XOR2_X1 U899 ( .A(G146), .B(n1260), .Z(G48) );
NOR3_X1 U900 ( .A1(n1261), .A2(n1079), .A3(n1221), .ZN(n1260) );
XNOR2_X1 U901 ( .A(KEYINPUT61), .B(n1232), .ZN(n1261) );
NAND2_X1 U902 ( .A1(n1262), .A2(n1263), .ZN(G45) );
OR2_X1 U903 ( .A1(n1233), .A2(G143), .ZN(n1263) );
XOR2_X1 U904 ( .A(n1264), .B(KEYINPUT38), .Z(n1262) );
NAND2_X1 U905 ( .A1(G143), .A2(n1233), .ZN(n1264) );
NAND4_X1 U906 ( .A1(n1231), .A2(n1229), .A3(n1223), .A4(n1230), .ZN(n1233) );
XNOR2_X1 U907 ( .A(G140), .B(n1212), .ZN(G42) );
NAND3_X1 U908 ( .A1(n1265), .A2(n1088), .A3(n1062), .ZN(n1212) );
XOR2_X1 U909 ( .A(G137), .B(n1266), .Z(G39) );
NOR3_X1 U910 ( .A1(n1235), .A2(n1055), .A3(n1221), .ZN(n1266) );
INV_X1 U911 ( .A(n1081), .ZN(n1055) );
XNOR2_X1 U912 ( .A(G134), .B(n1213), .ZN(G36) );
NAND3_X1 U913 ( .A1(n1062), .A2(n1246), .A3(n1229), .ZN(n1213) );
XNOR2_X1 U914 ( .A(G131), .B(n1219), .ZN(G33) );
NAND3_X1 U915 ( .A1(n1062), .A2(n1259), .A3(n1229), .ZN(n1219) );
AND3_X1 U916 ( .A1(n1088), .A2(n1267), .A3(n1252), .ZN(n1229) );
INV_X1 U917 ( .A(n1235), .ZN(n1062) );
NAND2_X1 U918 ( .A1(n1268), .A2(n1269), .ZN(n1235) );
NAND2_X1 U919 ( .A1(n1270), .A2(n1271), .ZN(G30) );
NAND2_X1 U920 ( .A1(n1220), .A2(n1272), .ZN(n1271) );
XOR2_X1 U921 ( .A(n1273), .B(KEYINPUT44), .Z(n1270) );
OR2_X1 U922 ( .A1(n1272), .A2(n1220), .ZN(n1273) );
NOR3_X1 U923 ( .A1(n1080), .A2(n1232), .A3(n1221), .ZN(n1220) );
NAND4_X1 U924 ( .A1(n1088), .A2(n1274), .A3(n1102), .A4(n1267), .ZN(n1221) );
INV_X1 U925 ( .A(n1246), .ZN(n1080) );
XOR2_X1 U926 ( .A(G128), .B(KEYINPUT11), .Z(n1272) );
XNOR2_X1 U927 ( .A(G101), .B(n1275), .ZN(G3) );
NAND3_X1 U928 ( .A1(n1252), .A2(n1245), .A3(n1081), .ZN(n1275) );
NOR3_X1 U929 ( .A1(n1063), .A2(n1258), .A3(n1255), .ZN(n1245) );
INV_X1 U930 ( .A(n1088), .ZN(n1063) );
XNOR2_X1 U931 ( .A(G125), .B(n1217), .ZN(G27) );
NAND2_X1 U932 ( .A1(n1265), .A2(n1059), .ZN(n1217) );
AND3_X1 U933 ( .A1(n1259), .A2(n1267), .A3(n1094), .ZN(n1265) );
NAND2_X1 U934 ( .A1(n1056), .A2(n1276), .ZN(n1267) );
NAND4_X1 U935 ( .A1(G953), .A2(G902), .A3(n1277), .A4(n1278), .ZN(n1276) );
INV_X1 U936 ( .A(G900), .ZN(n1278) );
XOR2_X1 U937 ( .A(n1279), .B(n1280), .Z(G24) );
XNOR2_X1 U938 ( .A(KEYINPUT54), .B(n1281), .ZN(n1280) );
NOR2_X1 U939 ( .A1(n1257), .A2(n1282), .ZN(n1279) );
XNOR2_X1 U940 ( .A(KEYINPUT3), .B(n1256), .ZN(n1282) );
NAND4_X1 U941 ( .A1(n1059), .A2(n1057), .A3(n1231), .A4(n1230), .ZN(n1257) );
NOR2_X1 U942 ( .A1(n1102), .A2(n1274), .ZN(n1057) );
NAND2_X1 U943 ( .A1(n1283), .A2(n1284), .ZN(G21) );
NAND2_X1 U944 ( .A1(G119), .A2(n1244), .ZN(n1284) );
XOR2_X1 U945 ( .A(n1285), .B(KEYINPUT31), .Z(n1283) );
OR2_X1 U946 ( .A1(n1244), .A2(G119), .ZN(n1285) );
NAND3_X1 U947 ( .A1(n1081), .A2(n1059), .A3(n1286), .ZN(n1244) );
AND3_X1 U948 ( .A1(n1274), .A2(n1256), .A3(n1102), .ZN(n1286) );
XNOR2_X1 U949 ( .A(G116), .B(n1243), .ZN(G18) );
NAND4_X1 U950 ( .A1(n1059), .A2(n1252), .A3(n1246), .A4(n1256), .ZN(n1243) );
NOR2_X1 U951 ( .A1(n1287), .A2(n1230), .ZN(n1246) );
NOR2_X1 U952 ( .A1(n1066), .A2(n1232), .ZN(n1059) );
INV_X1 U953 ( .A(n1223), .ZN(n1232) );
XNOR2_X1 U954 ( .A(n1255), .B(KEYINPUT48), .ZN(n1223) );
XNOR2_X1 U955 ( .A(G113), .B(n1242), .ZN(G15) );
NAND3_X1 U956 ( .A1(n1078), .A2(n1252), .A3(n1288), .ZN(n1242) );
NOR3_X1 U957 ( .A1(n1079), .A2(n1258), .A3(n1255), .ZN(n1288) );
INV_X1 U958 ( .A(n1259), .ZN(n1079) );
NOR2_X1 U959 ( .A1(n1097), .A2(n1231), .ZN(n1259) );
INV_X1 U960 ( .A(n1230), .ZN(n1097) );
INV_X1 U961 ( .A(n1092), .ZN(n1252) );
NAND2_X1 U962 ( .A1(n1289), .A2(n1102), .ZN(n1092) );
XNOR2_X1 U963 ( .A(n1274), .B(KEYINPUT43), .ZN(n1289) );
INV_X1 U964 ( .A(n1066), .ZN(n1078) );
NAND2_X1 U965 ( .A1(n1090), .A2(n1290), .ZN(n1066) );
XNOR2_X1 U966 ( .A(KEYINPUT40), .B(n1291), .ZN(n1290) );
XNOR2_X1 U967 ( .A(G110), .B(n1292), .ZN(G12) );
NAND4_X1 U968 ( .A1(n1094), .A2(n1081), .A3(n1293), .A4(n1088), .ZN(n1292) );
NOR2_X1 U969 ( .A1(n1090), .A2(n1089), .ZN(n1088) );
INV_X1 U970 ( .A(n1291), .ZN(n1089) );
NAND2_X1 U971 ( .A1(G221), .A2(n1294), .ZN(n1291) );
INV_X1 U972 ( .A(n1101), .ZN(n1090) );
XNOR2_X1 U973 ( .A(n1295), .B(G469), .ZN(n1101) );
NAND2_X1 U974 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
XOR2_X1 U975 ( .A(n1298), .B(n1299), .Z(n1296) );
XOR2_X1 U976 ( .A(n1208), .B(n1300), .Z(n1299) );
NOR2_X1 U977 ( .A1(KEYINPUT39), .A2(n1201), .ZN(n1300) );
NAND2_X1 U978 ( .A1(G227), .A2(n1125), .ZN(n1201) );
XOR2_X1 U979 ( .A(n1301), .B(n1302), .Z(n1298) );
NOR2_X1 U980 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
XOR2_X1 U981 ( .A(n1305), .B(KEYINPUT14), .Z(n1304) );
NAND2_X1 U982 ( .A1(n1306), .A2(n1133), .ZN(n1305) );
NOR2_X1 U983 ( .A1(n1133), .A2(n1306), .ZN(n1303) );
XNOR2_X1 U984 ( .A(n1307), .B(n1203), .ZN(n1306) );
XOR2_X1 U985 ( .A(G101), .B(n1308), .Z(n1203) );
NOR2_X1 U986 ( .A1(KEYINPUT26), .A2(n1309), .ZN(n1308) );
XNOR2_X1 U987 ( .A(G104), .B(G107), .ZN(n1309) );
NAND2_X1 U988 ( .A1(KEYINPUT20), .A2(n1204), .ZN(n1307) );
XNOR2_X1 U989 ( .A(n1132), .B(KEYINPUT10), .ZN(n1204) );
NAND2_X1 U990 ( .A1(n1310), .A2(n1311), .ZN(n1132) );
NAND2_X1 U991 ( .A1(n1312), .A2(G128), .ZN(n1311) );
XNOR2_X1 U992 ( .A(G143), .B(n1313), .ZN(n1312) );
XOR2_X1 U993 ( .A(n1314), .B(KEYINPUT59), .Z(n1310) );
NAND2_X1 U994 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XNOR2_X1 U995 ( .A(n1317), .B(n1313), .ZN(n1315) );
NOR2_X1 U996 ( .A1(KEYINPUT19), .A2(G146), .ZN(n1313) );
XNOR2_X1 U997 ( .A(KEYINPUT16), .B(n1318), .ZN(n1301) );
NOR2_X1 U998 ( .A1(G140), .A2(KEYINPUT7), .ZN(n1318) );
NOR2_X1 U999 ( .A1(n1258), .A2(n1319), .ZN(n1293) );
XOR2_X1 U1000 ( .A(n1255), .B(KEYINPUT34), .Z(n1319) );
NAND2_X1 U1001 ( .A1(n1269), .A2(n1064), .ZN(n1255) );
INV_X1 U1002 ( .A(n1268), .ZN(n1064) );
NOR2_X1 U1003 ( .A1(n1320), .A2(n1105), .ZN(n1268) );
NOR3_X1 U1004 ( .A1(n1321), .A2(G902), .A3(n1115), .ZN(n1105) );
AND2_X1 U1005 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
OR2_X1 U1006 ( .A1(n1115), .A2(G902), .ZN(n1322) );
XNOR2_X1 U1007 ( .A(n1323), .B(n1324), .ZN(n1115) );
XNOR2_X1 U1008 ( .A(n1141), .B(n1186), .ZN(n1324) );
XOR2_X1 U1009 ( .A(n1325), .B(n1326), .Z(n1141) );
XNOR2_X1 U1010 ( .A(n1327), .B(n1328), .ZN(n1326) );
XOR2_X1 U1011 ( .A(n1329), .B(n1330), .Z(n1328) );
NAND2_X1 U1012 ( .A1(n1331), .A2(n1332), .ZN(n1329) );
NAND2_X1 U1013 ( .A1(n1208), .A2(G122), .ZN(n1332) );
XOR2_X1 U1014 ( .A(KEYINPUT36), .B(n1333), .Z(n1331) );
NOR2_X1 U1015 ( .A1(G122), .A2(n1208), .ZN(n1333) );
XOR2_X1 U1016 ( .A(n1334), .B(n1335), .Z(n1325) );
XNOR2_X1 U1017 ( .A(n1336), .B(G101), .ZN(n1335) );
INV_X1 U1018 ( .A(G107), .ZN(n1336) );
XNOR2_X1 U1019 ( .A(KEYINPUT50), .B(KEYINPUT4), .ZN(n1334) );
XNOR2_X1 U1020 ( .A(G125), .B(n1337), .ZN(n1323) );
AND2_X1 U1021 ( .A1(n1125), .A2(G224), .ZN(n1337) );
INV_X1 U1022 ( .A(n1114), .ZN(n1321) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1338), .ZN(n1114) );
XNOR2_X1 U1024 ( .A(n1112), .B(KEYINPUT52), .ZN(n1269) );
INV_X1 U1025 ( .A(n1065), .ZN(n1112) );
NAND2_X1 U1026 ( .A1(G214), .A2(n1338), .ZN(n1065) );
NAND2_X1 U1027 ( .A1(n1339), .A2(n1297), .ZN(n1338) );
INV_X1 U1028 ( .A(n1256), .ZN(n1258) );
NAND2_X1 U1029 ( .A1(n1056), .A2(n1340), .ZN(n1256) );
NAND4_X1 U1030 ( .A1(G953), .A2(G902), .A3(n1277), .A4(n1143), .ZN(n1340) );
INV_X1 U1031 ( .A(G898), .ZN(n1143) );
NAND3_X1 U1032 ( .A1(n1277), .A2(n1125), .A3(G952), .ZN(n1056) );
NAND2_X1 U1033 ( .A1(G237), .A2(G234), .ZN(n1277) );
NOR2_X1 U1034 ( .A1(n1230), .A2(n1231), .ZN(n1081) );
INV_X1 U1035 ( .A(n1287), .ZN(n1231) );
NAND2_X1 U1036 ( .A1(n1341), .A2(n1342), .ZN(n1287) );
NAND2_X1 U1037 ( .A1(KEYINPUT25), .A2(n1343), .ZN(n1342) );
NAND2_X1 U1038 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
NAND2_X1 U1039 ( .A1(n1346), .A2(n1159), .ZN(n1345) );
INV_X1 U1040 ( .A(n1107), .ZN(n1344) );
NOR2_X1 U1041 ( .A1(n1346), .A2(n1159), .ZN(n1107) );
INV_X1 U1042 ( .A(n1110), .ZN(n1346) );
NAND2_X1 U1043 ( .A1(n1347), .A2(n1348), .ZN(n1341) );
INV_X1 U1044 ( .A(KEYINPUT25), .ZN(n1348) );
XNOR2_X1 U1045 ( .A(n1159), .B(n1110), .ZN(n1347) );
NOR2_X1 U1046 ( .A1(n1161), .A2(G902), .ZN(n1110) );
INV_X1 U1047 ( .A(n1158), .ZN(n1161) );
XNOR2_X1 U1048 ( .A(n1349), .B(n1350), .ZN(n1158) );
NOR2_X1 U1049 ( .A1(KEYINPUT24), .A2(n1351), .ZN(n1350) );
XOR2_X1 U1050 ( .A(n1352), .B(n1353), .Z(n1351) );
XNOR2_X1 U1051 ( .A(n1316), .B(n1354), .ZN(n1353) );
XNOR2_X1 U1052 ( .A(n1317), .B(G134), .ZN(n1354) );
XNOR2_X1 U1053 ( .A(G107), .B(n1355), .ZN(n1352) );
XNOR2_X1 U1054 ( .A(n1281), .B(G116), .ZN(n1355) );
INV_X1 U1055 ( .A(G122), .ZN(n1281) );
NAND2_X1 U1056 ( .A1(G217), .A2(n1356), .ZN(n1349) );
INV_X1 U1057 ( .A(n1357), .ZN(n1356) );
INV_X1 U1058 ( .A(G478), .ZN(n1159) );
XNOR2_X1 U1059 ( .A(n1358), .B(G475), .ZN(n1230) );
NAND2_X1 U1060 ( .A1(n1165), .A2(n1297), .ZN(n1358) );
XNOR2_X1 U1061 ( .A(n1359), .B(n1360), .ZN(n1165) );
XNOR2_X1 U1062 ( .A(n1330), .B(n1361), .ZN(n1360) );
XOR2_X1 U1063 ( .A(n1362), .B(n1363), .Z(n1361) );
NOR4_X1 U1064 ( .A1(n1364), .A2(n1365), .A3(KEYINPUT51), .A4(n1366), .ZN(n1363) );
AND2_X1 U1065 ( .A1(n1367), .A2(KEYINPUT15), .ZN(n1366) );
NOR2_X1 U1066 ( .A1(n1368), .A2(n1317), .ZN(n1365) );
NOR2_X1 U1067 ( .A1(KEYINPUT0), .A2(n1367), .ZN(n1368) );
NOR4_X1 U1068 ( .A1(G143), .A2(n1367), .A3(KEYINPUT15), .A4(KEYINPUT0), .ZN(n1364) );
NAND3_X1 U1069 ( .A1(n1339), .A2(n1125), .A3(G214), .ZN(n1367) );
NAND2_X1 U1070 ( .A1(n1369), .A2(n1370), .ZN(n1362) );
XOR2_X1 U1071 ( .A(n1371), .B(KEYINPUT32), .Z(n1369) );
XOR2_X1 U1072 ( .A(G104), .B(G113), .Z(n1330) );
XNOR2_X1 U1073 ( .A(G122), .B(n1372), .ZN(n1359) );
XNOR2_X1 U1074 ( .A(G146), .B(n1373), .ZN(n1372) );
INV_X1 U1075 ( .A(G131), .ZN(n1373) );
NOR2_X1 U1076 ( .A1(n1102), .A2(n1116), .ZN(n1094) );
INV_X1 U1077 ( .A(n1274), .ZN(n1116) );
XOR2_X1 U1078 ( .A(n1374), .B(n1153), .Z(n1274) );
NAND2_X1 U1079 ( .A1(G217), .A2(n1294), .ZN(n1153) );
NAND2_X1 U1080 ( .A1(G234), .A2(n1297), .ZN(n1294) );
OR2_X1 U1081 ( .A1(n1152), .A2(G902), .ZN(n1374) );
XNOR2_X1 U1082 ( .A(n1375), .B(n1376), .ZN(n1152) );
XOR2_X1 U1083 ( .A(n1377), .B(n1378), .Z(n1376) );
XOR2_X1 U1084 ( .A(G146), .B(G137), .Z(n1378) );
XOR2_X1 U1085 ( .A(KEYINPUT46), .B(KEYINPUT35), .Z(n1377) );
XOR2_X1 U1086 ( .A(n1126), .B(n1379), .Z(n1375) );
XOR2_X1 U1087 ( .A(n1380), .B(n1381), .Z(n1379) );
NOR3_X1 U1088 ( .A1(n1382), .A2(KEYINPUT27), .A3(n1357), .ZN(n1381) );
NAND2_X1 U1089 ( .A1(G234), .A2(n1125), .ZN(n1357) );
INV_X1 U1090 ( .A(G221), .ZN(n1382) );
NOR2_X1 U1091 ( .A1(n1383), .A2(n1384), .ZN(n1380) );
XOR2_X1 U1092 ( .A(n1385), .B(KEYINPUT18), .Z(n1384) );
NAND2_X1 U1093 ( .A1(n1208), .A2(n1386), .ZN(n1385) );
XOR2_X1 U1094 ( .A(KEYINPUT12), .B(n1387), .Z(n1386) );
NOR2_X1 U1095 ( .A1(n1208), .A2(n1387), .ZN(n1383) );
XNOR2_X1 U1096 ( .A(n1388), .B(G119), .ZN(n1387) );
NAND2_X1 U1097 ( .A1(KEYINPUT58), .A2(n1316), .ZN(n1388) );
XNOR2_X1 U1098 ( .A(G110), .B(KEYINPUT41), .ZN(n1208) );
NAND2_X1 U1099 ( .A1(n1370), .A2(n1371), .ZN(n1126) );
NAND2_X1 U1100 ( .A1(G125), .A2(n1389), .ZN(n1371) );
OR2_X1 U1101 ( .A1(n1389), .A2(G125), .ZN(n1370) );
INV_X1 U1102 ( .A(G140), .ZN(n1389) );
XNOR2_X1 U1103 ( .A(n1390), .B(G472), .ZN(n1102) );
NAND2_X1 U1104 ( .A1(n1391), .A2(n1297), .ZN(n1390) );
INV_X1 U1105 ( .A(G902), .ZN(n1297) );
XNOR2_X1 U1106 ( .A(n1175), .B(n1392), .ZN(n1391) );
XOR2_X1 U1107 ( .A(G101), .B(n1393), .Z(n1392) );
NOR2_X1 U1108 ( .A1(KEYINPUT2), .A2(n1394), .ZN(n1393) );
XNOR2_X1 U1109 ( .A(n1180), .B(n1395), .ZN(n1394) );
XNOR2_X1 U1110 ( .A(n1133), .B(n1185), .ZN(n1395) );
INV_X1 U1111 ( .A(n1186), .ZN(n1185) );
XNOR2_X1 U1112 ( .A(n1396), .B(n1397), .ZN(n1186) );
XNOR2_X1 U1113 ( .A(G146), .B(n1316), .ZN(n1397) );
INV_X1 U1114 ( .A(G128), .ZN(n1316) );
NAND2_X1 U1115 ( .A1(KEYINPUT13), .A2(n1317), .ZN(n1396) );
INV_X1 U1116 ( .A(G143), .ZN(n1317) );
XOR2_X1 U1117 ( .A(G131), .B(n1398), .Z(n1133) );
XOR2_X1 U1118 ( .A(G137), .B(G134), .Z(n1398) );
XNOR2_X1 U1119 ( .A(G113), .B(n1327), .ZN(n1180) );
XOR2_X1 U1120 ( .A(G116), .B(G119), .Z(n1327) );
NAND3_X1 U1121 ( .A1(n1339), .A2(n1125), .A3(G210), .ZN(n1175) );
INV_X1 U1122 ( .A(G953), .ZN(n1125) );
INV_X1 U1123 ( .A(G237), .ZN(n1339) );
endmodule


