//Key = 1110101000011010000000001001010010101110100110110111010011000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373;

XOR2_X1 U757 ( .A(n1043), .B(n1044), .Z(G9) );
NOR2_X1 U758 ( .A1(G107), .A2(KEYINPUT33), .ZN(n1044) );
NOR2_X1 U759 ( .A1(n1045), .A2(n1046), .ZN(G75) );
XOR2_X1 U760 ( .A(n1047), .B(KEYINPUT44), .Z(n1046) );
NAND3_X1 U761 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
XOR2_X1 U762 ( .A(n1051), .B(KEYINPUT25), .Z(n1050) );
NOR4_X1 U763 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1048), .ZN(n1045) );
INV_X1 U764 ( .A(G952), .ZN(n1048) );
NOR2_X1 U765 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
AND3_X1 U766 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1055) );
NAND4_X1 U767 ( .A1(n1060), .A2(n1061), .A3(n1051), .A4(n1049), .ZN(n1052) );
NAND4_X1 U768 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1051) );
NOR3_X1 U769 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
XOR2_X1 U770 ( .A(n1069), .B(n1070), .Z(n1066) );
XOR2_X1 U771 ( .A(KEYINPUT50), .B(n1071), .Z(n1062) );
NAND4_X1 U772 ( .A1(n1072), .A2(n1059), .A3(n1073), .A4(n1074), .ZN(n1061) );
NAND2_X1 U773 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND3_X1 U774 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1076) );
NAND2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NAND3_X1 U776 ( .A1(n1082), .A2(n1083), .A3(n1063), .ZN(n1077) );
NAND2_X1 U777 ( .A1(n1084), .A2(n1085), .ZN(n1075) );
INV_X1 U778 ( .A(n1086), .ZN(n1072) );
NAND2_X1 U779 ( .A1(n1057), .A2(n1087), .ZN(n1060) );
NAND2_X1 U780 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U781 ( .A1(n1073), .A2(n1090), .ZN(n1089) );
NAND2_X1 U782 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U783 ( .A1(n1059), .A2(n1093), .ZN(n1088) );
NAND2_X1 U784 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U785 ( .A1(n1058), .A2(n1056), .ZN(n1095) );
INV_X1 U786 ( .A(KEYINPUT42), .ZN(n1056) );
NAND2_X1 U787 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NOR4_X1 U788 ( .A1(n1071), .A2(n1086), .A3(n1081), .A4(n1080), .ZN(n1057) );
NAND2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(G72) );
NAND2_X1 U790 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
INV_X1 U791 ( .A(n1102), .ZN(n1100) );
XOR2_X1 U792 ( .A(n1103), .B(KEYINPUT41), .Z(n1098) );
NAND2_X1 U793 ( .A1(n1104), .A2(n1102), .ZN(n1103) );
NAND2_X1 U794 ( .A1(G953), .A2(n1105), .ZN(n1102) );
XOR2_X1 U795 ( .A(KEYINPUT12), .B(n1106), .Z(n1105) );
NOR2_X1 U796 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U797 ( .A(n1101), .B(n1109), .ZN(n1104) );
NOR2_X1 U798 ( .A1(n1110), .A2(G953), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1111), .A2(n1112), .ZN(n1101) );
NAND2_X1 U800 ( .A1(G953), .A2(n1108), .ZN(n1112) );
XOR2_X1 U801 ( .A(n1113), .B(n1114), .Z(n1111) );
NOR2_X1 U802 ( .A1(KEYINPUT23), .A2(n1115), .ZN(n1114) );
XOR2_X1 U803 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U805 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U806 ( .A(KEYINPUT46), .B(n1122), .Z(n1120) );
NAND2_X1 U807 ( .A1(G131), .A2(n1123), .ZN(n1118) );
XNOR2_X1 U808 ( .A(n1122), .B(KEYINPUT34), .ZN(n1123) );
NAND2_X1 U809 ( .A1(KEYINPUT53), .A2(n1124), .ZN(n1116) );
NAND3_X1 U810 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(G69) );
NAND2_X1 U811 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U812 ( .A1(KEYINPUT60), .A2(n1130), .ZN(n1126) );
NAND2_X1 U813 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XNOR2_X1 U814 ( .A(n1133), .B(n1129), .ZN(n1131) );
NAND2_X1 U815 ( .A1(n1134), .A2(n1135), .ZN(n1125) );
INV_X1 U816 ( .A(KEYINPUT60), .ZN(n1135) );
NAND2_X1 U817 ( .A1(n1136), .A2(n1137), .ZN(n1134) );
OR3_X1 U818 ( .A1(n1129), .A2(n1128), .A3(n1133), .ZN(n1137) );
INV_X1 U819 ( .A(n1132), .ZN(n1128) );
NAND2_X1 U820 ( .A1(n1138), .A2(G953), .ZN(n1132) );
XOR2_X1 U821 ( .A(n1139), .B(KEYINPUT26), .Z(n1138) );
NAND2_X1 U822 ( .A1(G898), .A2(G224), .ZN(n1139) );
NAND2_X1 U823 ( .A1(n1133), .A2(n1129), .ZN(n1136) );
NAND2_X1 U824 ( .A1(n1140), .A2(n1141), .ZN(n1129) );
NAND2_X1 U825 ( .A1(G953), .A2(n1142), .ZN(n1141) );
XNOR2_X1 U826 ( .A(n1143), .B(n1144), .ZN(n1140) );
NAND2_X1 U827 ( .A1(KEYINPUT11), .A2(n1145), .ZN(n1143) );
NOR2_X1 U828 ( .A1(n1146), .A2(G953), .ZN(n1133) );
NOR2_X1 U829 ( .A1(n1147), .A2(n1148), .ZN(G66) );
XNOR2_X1 U830 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR2_X1 U831 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U832 ( .A1(n1147), .A2(n1153), .ZN(G63) );
XOR2_X1 U833 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U834 ( .A(KEYINPUT4), .B(n1156), .Z(n1155) );
NOR2_X1 U835 ( .A1(n1157), .A2(n1152), .ZN(n1156) );
XNOR2_X1 U836 ( .A(G478), .B(KEYINPUT52), .ZN(n1157) );
NOR3_X1 U837 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(G60) );
AND2_X1 U838 ( .A1(KEYINPUT24), .A2(n1147), .ZN(n1160) );
NOR3_X1 U839 ( .A1(KEYINPUT24), .A2(G953), .A3(G952), .ZN(n1159) );
XNOR2_X1 U840 ( .A(n1161), .B(n1162), .ZN(n1158) );
NOR2_X1 U841 ( .A1(n1163), .A2(n1152), .ZN(n1162) );
INV_X1 U842 ( .A(G475), .ZN(n1163) );
XOR2_X1 U843 ( .A(G104), .B(n1164), .Z(G6) );
NOR2_X1 U844 ( .A1(n1147), .A2(n1165), .ZN(G57) );
NOR2_X1 U845 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U846 ( .A(KEYINPUT17), .B(n1168), .Z(n1167) );
NOR2_X1 U847 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
AND2_X1 U848 ( .A1(n1170), .A2(n1169), .ZN(n1166) );
XNOR2_X1 U849 ( .A(n1171), .B(n1172), .ZN(n1170) );
NOR2_X1 U850 ( .A1(n1069), .A2(n1152), .ZN(n1172) );
NAND2_X1 U851 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
XOR2_X1 U852 ( .A(n1175), .B(KEYINPUT16), .Z(n1173) );
NOR2_X1 U853 ( .A1(n1147), .A2(n1176), .ZN(G54) );
NOR2_X1 U854 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR2_X1 U855 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NOR2_X1 U856 ( .A1(n1181), .A2(n1182), .ZN(n1177) );
XOR2_X1 U857 ( .A(KEYINPUT0), .B(n1180), .Z(n1182) );
XNOR2_X1 U858 ( .A(n1183), .B(n1184), .ZN(n1180) );
XOR2_X1 U859 ( .A(n1185), .B(n1186), .Z(n1184) );
XNOR2_X1 U860 ( .A(KEYINPUT13), .B(KEYINPUT10), .ZN(n1186) );
XOR2_X1 U861 ( .A(n1187), .B(n1188), .Z(n1183) );
XOR2_X1 U862 ( .A(n1189), .B(n1190), .Z(n1187) );
XOR2_X1 U863 ( .A(KEYINPUT2), .B(n1179), .Z(n1181) );
NOR2_X1 U864 ( .A1(n1152), .A2(n1191), .ZN(n1179) );
NOR2_X1 U865 ( .A1(n1147), .A2(n1192), .ZN(G51) );
XOR2_X1 U866 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U867 ( .A(n1195), .B(n1196), .Z(n1194) );
XNOR2_X1 U868 ( .A(KEYINPUT15), .B(n1197), .ZN(n1193) );
NOR3_X1 U869 ( .A1(n1152), .A2(KEYINPUT35), .A3(n1198), .ZN(n1197) );
NAND2_X1 U870 ( .A1(n1199), .A2(n1053), .ZN(n1152) );
NAND2_X1 U871 ( .A1(n1110), .A2(n1146), .ZN(n1053) );
AND4_X1 U872 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1146) );
AND4_X1 U873 ( .A1(n1043), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1203) );
OR3_X1 U874 ( .A1(n1207), .A2(n1092), .A3(n1081), .ZN(n1043) );
NOR2_X1 U875 ( .A1(n1164), .A2(n1208), .ZN(n1202) );
NOR3_X1 U876 ( .A1(n1068), .A2(n1207), .A3(n1083), .ZN(n1208) );
NOR3_X1 U877 ( .A1(n1081), .A2(n1207), .A3(n1091), .ZN(n1164) );
INV_X1 U878 ( .A(n1084), .ZN(n1081) );
AND2_X1 U879 ( .A1(n1209), .A2(n1210), .ZN(n1110) );
AND4_X1 U880 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1210) );
NOR4_X1 U881 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1209) );
NOR4_X1 U882 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1218) );
AND2_X1 U883 ( .A1(KEYINPUT37), .A2(n1223), .ZN(n1222) );
NOR3_X1 U884 ( .A1(KEYINPUT37), .A2(n1224), .A3(n1223), .ZN(n1221) );
NAND2_X1 U885 ( .A1(n1225), .A2(n1226), .ZN(n1219) );
NAND2_X1 U886 ( .A1(n1227), .A2(n1091), .ZN(n1226) );
INV_X1 U887 ( .A(n1228), .ZN(n1217) );
AND3_X1 U888 ( .A1(KEYINPUT30), .A2(n1092), .A3(n1229), .ZN(n1216) );
NOR2_X1 U889 ( .A1(KEYINPUT30), .A2(n1230), .ZN(n1215) );
XOR2_X1 U890 ( .A(n1231), .B(KEYINPUT49), .Z(n1199) );
NOR2_X1 U891 ( .A1(n1049), .A2(G952), .ZN(n1147) );
NAND3_X1 U892 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(G48) );
OR2_X1 U893 ( .A1(n1235), .A2(G146), .ZN(n1234) );
NAND2_X1 U894 ( .A1(KEYINPUT62), .A2(n1236), .ZN(n1233) );
NAND2_X1 U895 ( .A1(G146), .A2(n1237), .ZN(n1236) );
XNOR2_X1 U896 ( .A(KEYINPUT43), .B(n1235), .ZN(n1237) );
NAND2_X1 U897 ( .A1(n1238), .A2(n1239), .ZN(n1232) );
INV_X1 U898 ( .A(KEYINPUT62), .ZN(n1239) );
NAND2_X1 U899 ( .A1(n1240), .A2(n1241), .ZN(n1238) );
NAND3_X1 U900 ( .A1(KEYINPUT43), .A2(G146), .A3(n1235), .ZN(n1241) );
OR2_X1 U901 ( .A1(n1235), .A2(KEYINPUT43), .ZN(n1240) );
NAND3_X1 U902 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1235) );
NOR3_X1 U903 ( .A1(n1245), .A2(n1223), .A3(n1246), .ZN(n1244) );
XOR2_X1 U904 ( .A(n1247), .B(KEYINPUT63), .Z(n1246) );
XOR2_X1 U905 ( .A(G143), .B(n1248), .Z(G45) );
NOR2_X1 U906 ( .A1(KEYINPUT39), .A2(n1228), .ZN(n1248) );
NAND3_X1 U907 ( .A1(n1249), .A2(n1225), .A3(n1250), .ZN(n1228) );
NOR3_X1 U908 ( .A1(n1251), .A2(n1223), .A3(n1252), .ZN(n1250) );
XOR2_X1 U909 ( .A(n1185), .B(n1214), .Z(G42) );
NAND3_X1 U910 ( .A1(n1243), .A2(n1253), .A3(n1254), .ZN(n1214) );
XNOR2_X1 U911 ( .A(G137), .B(n1213), .ZN(G39) );
NAND3_X1 U912 ( .A1(n1059), .A2(n1254), .A3(n1242), .ZN(n1213) );
XOR2_X1 U913 ( .A(n1255), .B(n1230), .Z(G36) );
NAND2_X1 U914 ( .A1(n1229), .A2(n1224), .ZN(n1230) );
NAND2_X1 U915 ( .A1(n1256), .A2(G134), .ZN(n1255) );
XNOR2_X1 U916 ( .A(KEYINPUT7), .B(KEYINPUT58), .ZN(n1256) );
XOR2_X1 U917 ( .A(n1121), .B(n1212), .Z(G33) );
NAND2_X1 U918 ( .A1(n1229), .A2(n1243), .ZN(n1212) );
AND2_X1 U919 ( .A1(n1249), .A2(n1254), .ZN(n1229) );
NOR4_X1 U920 ( .A1(n1071), .A2(n1245), .A3(n1223), .A4(n1080), .ZN(n1254) );
INV_X1 U921 ( .A(n1063), .ZN(n1080) );
INV_X1 U922 ( .A(n1058), .ZN(n1245) );
XOR2_X1 U923 ( .A(G128), .B(n1257), .Z(G30) );
NOR4_X1 U924 ( .A1(KEYINPUT55), .A2(n1258), .A3(n1220), .A4(n1227), .ZN(n1257) );
NAND2_X1 U925 ( .A1(n1224), .A2(n1259), .ZN(n1227) );
XOR2_X1 U926 ( .A(G101), .B(n1260), .Z(G3) );
NOR3_X1 U927 ( .A1(n1068), .A2(n1261), .A3(n1207), .ZN(n1260) );
XOR2_X1 U928 ( .A(n1083), .B(KEYINPUT61), .Z(n1261) );
XNOR2_X1 U929 ( .A(G125), .B(n1211), .ZN(G27) );
NAND4_X1 U930 ( .A1(n1243), .A2(n1073), .A3(n1262), .A4(n1253), .ZN(n1211) );
NOR2_X1 U931 ( .A1(n1223), .A2(n1247), .ZN(n1262) );
INV_X1 U932 ( .A(n1259), .ZN(n1223) );
NAND2_X1 U933 ( .A1(n1086), .A2(n1263), .ZN(n1259) );
NAND2_X1 U934 ( .A1(n1264), .A2(n1108), .ZN(n1263) );
INV_X1 U935 ( .A(G900), .ZN(n1108) );
NAND2_X1 U936 ( .A1(n1265), .A2(n1266), .ZN(G24) );
NAND2_X1 U937 ( .A1(G122), .A2(n1200), .ZN(n1266) );
XOR2_X1 U938 ( .A(n1267), .B(KEYINPUT22), .Z(n1265) );
OR2_X1 U939 ( .A1(n1200), .A2(G122), .ZN(n1267) );
NAND4_X1 U940 ( .A1(n1268), .A2(n1084), .A3(n1269), .A4(n1270), .ZN(n1200) );
NOR2_X1 U941 ( .A1(n1271), .A2(n1272), .ZN(n1084) );
XOR2_X1 U942 ( .A(n1201), .B(n1273), .Z(G21) );
NAND2_X1 U943 ( .A1(KEYINPUT1), .A2(G119), .ZN(n1273) );
NAND3_X1 U944 ( .A1(n1242), .A2(n1059), .A3(n1268), .ZN(n1201) );
INV_X1 U945 ( .A(n1068), .ZN(n1059) );
INV_X1 U946 ( .A(n1220), .ZN(n1242) );
NAND2_X1 U947 ( .A1(n1272), .A2(n1271), .ZN(n1220) );
INV_X1 U948 ( .A(n1064), .ZN(n1272) );
XNOR2_X1 U949 ( .A(G116), .B(n1206), .ZN(G18) );
NAND3_X1 U950 ( .A1(n1249), .A2(n1224), .A3(n1268), .ZN(n1206) );
INV_X1 U951 ( .A(n1092), .ZN(n1224) );
NAND2_X1 U952 ( .A1(n1252), .A2(n1269), .ZN(n1092) );
INV_X1 U953 ( .A(n1251), .ZN(n1269) );
XOR2_X1 U954 ( .A(n1274), .B(n1205), .Z(G15) );
NAND3_X1 U955 ( .A1(n1249), .A2(n1243), .A3(n1268), .ZN(n1205) );
AND3_X1 U956 ( .A1(n1085), .A2(n1275), .A3(n1073), .ZN(n1268) );
INV_X1 U957 ( .A(n1067), .ZN(n1073) );
NAND2_X1 U958 ( .A1(n1097), .A2(n1276), .ZN(n1067) );
INV_X1 U959 ( .A(n1091), .ZN(n1243) );
NAND2_X1 U960 ( .A1(n1251), .A2(n1270), .ZN(n1091) );
INV_X1 U961 ( .A(n1252), .ZN(n1270) );
INV_X1 U962 ( .A(n1083), .ZN(n1249) );
NAND2_X1 U963 ( .A1(n1064), .A2(n1271), .ZN(n1083) );
XNOR2_X1 U964 ( .A(G110), .B(n1204), .ZN(G12) );
OR3_X1 U965 ( .A1(n1082), .A2(n1207), .A3(n1068), .ZN(n1204) );
NAND2_X1 U966 ( .A1(n1251), .A2(n1252), .ZN(n1068) );
XOR2_X1 U967 ( .A(n1277), .B(G475), .Z(n1252) );
NAND2_X1 U968 ( .A1(n1161), .A2(n1231), .ZN(n1277) );
XNOR2_X1 U969 ( .A(n1278), .B(n1279), .ZN(n1161) );
XOR2_X1 U970 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U971 ( .A(n1282), .B(n1283), .Z(n1281) );
NAND2_X1 U972 ( .A1(G214), .A2(n1284), .ZN(n1282) );
XNOR2_X1 U973 ( .A(n1285), .B(n1286), .ZN(n1280) );
NOR2_X1 U974 ( .A1(KEYINPUT19), .A2(n1287), .ZN(n1286) );
NOR2_X1 U975 ( .A1(G122), .A2(KEYINPUT21), .ZN(n1285) );
XOR2_X1 U976 ( .A(n1288), .B(n1289), .Z(n1278) );
XOR2_X1 U977 ( .A(G143), .B(G131), .Z(n1289) );
XOR2_X1 U978 ( .A(G104), .B(n1274), .Z(n1288) );
XOR2_X1 U979 ( .A(n1290), .B(G478), .Z(n1251) );
NAND2_X1 U980 ( .A1(n1154), .A2(n1231), .ZN(n1290) );
XOR2_X1 U981 ( .A(n1291), .B(n1292), .Z(n1154) );
XOR2_X1 U982 ( .A(G116), .B(n1293), .Z(n1292) );
XOR2_X1 U983 ( .A(G134), .B(G122), .Z(n1293) );
XOR2_X1 U984 ( .A(n1294), .B(n1295), .Z(n1291) );
AND2_X1 U985 ( .A1(G217), .A2(n1296), .ZN(n1295) );
XNOR2_X1 U986 ( .A(n1297), .B(n1298), .ZN(n1294) );
NAND2_X1 U987 ( .A1(KEYINPUT51), .A2(G107), .ZN(n1298) );
NAND2_X1 U988 ( .A1(KEYINPUT40), .A2(n1299), .ZN(n1297) );
NAND2_X1 U989 ( .A1(n1225), .A2(n1275), .ZN(n1207) );
NAND2_X1 U990 ( .A1(n1086), .A2(n1300), .ZN(n1275) );
NAND2_X1 U991 ( .A1(n1264), .A2(n1142), .ZN(n1300) );
INV_X1 U992 ( .A(G898), .ZN(n1142) );
AND3_X1 U993 ( .A1(n1301), .A2(n1302), .A3(G953), .ZN(n1264) );
XOR2_X1 U994 ( .A(KEYINPUT45), .B(G902), .Z(n1301) );
NAND3_X1 U995 ( .A1(n1302), .A2(n1049), .A3(G952), .ZN(n1086) );
NAND2_X1 U996 ( .A1(G237), .A2(G234), .ZN(n1302) );
INV_X1 U997 ( .A(n1258), .ZN(n1225) );
NAND2_X1 U998 ( .A1(n1085), .A2(n1058), .ZN(n1258) );
NOR2_X1 U999 ( .A1(n1097), .A2(n1096), .ZN(n1058) );
INV_X1 U1000 ( .A(n1276), .ZN(n1096) );
NAND2_X1 U1001 ( .A1(G221), .A2(n1303), .ZN(n1276) );
XNOR2_X1 U1002 ( .A(n1304), .B(n1191), .ZN(n1097) );
INV_X1 U1003 ( .A(G469), .ZN(n1191) );
NAND2_X1 U1004 ( .A1(n1305), .A2(n1231), .ZN(n1304) );
XOR2_X1 U1005 ( .A(n1189), .B(n1306), .Z(n1305) );
XNOR2_X1 U1006 ( .A(n1307), .B(n1308), .ZN(n1306) );
NAND2_X1 U1007 ( .A1(KEYINPUT38), .A2(n1185), .ZN(n1308) );
INV_X1 U1008 ( .A(G140), .ZN(n1185) );
NAND3_X1 U1009 ( .A1(n1309), .A2(n1310), .A3(KEYINPUT6), .ZN(n1307) );
NAND2_X1 U1010 ( .A1(n1188), .A2(n1311), .ZN(n1310) );
NAND2_X1 U1011 ( .A1(KEYINPUT29), .A2(n1312), .ZN(n1311) );
NAND2_X1 U1012 ( .A1(n1190), .A2(n1313), .ZN(n1312) );
INV_X1 U1013 ( .A(n1314), .ZN(n1188) );
NAND2_X1 U1014 ( .A1(n1315), .A2(n1316), .ZN(n1309) );
NAND2_X1 U1015 ( .A1(n1313), .A2(n1317), .ZN(n1316) );
NAND2_X1 U1016 ( .A1(n1314), .A2(KEYINPUT29), .ZN(n1317) );
XOR2_X1 U1017 ( .A(n1124), .B(KEYINPUT31), .Z(n1314) );
XOR2_X1 U1018 ( .A(n1299), .B(n1318), .Z(n1124) );
XNOR2_X1 U1019 ( .A(n1319), .B(KEYINPUT56), .ZN(n1318) );
NAND2_X1 U1020 ( .A1(KEYINPUT27), .A2(n1320), .ZN(n1319) );
XOR2_X1 U1021 ( .A(n1321), .B(G143), .Z(n1299) );
INV_X1 U1022 ( .A(G128), .ZN(n1321) );
INV_X1 U1023 ( .A(KEYINPUT5), .ZN(n1313) );
XOR2_X1 U1024 ( .A(n1322), .B(n1323), .Z(n1189) );
XOR2_X1 U1025 ( .A(G110), .B(n1324), .Z(n1323) );
NOR2_X1 U1026 ( .A1(G953), .A2(n1107), .ZN(n1324) );
INV_X1 U1027 ( .A(G227), .ZN(n1107) );
INV_X1 U1028 ( .A(n1247), .ZN(n1085) );
NAND2_X1 U1029 ( .A1(n1071), .A2(n1063), .ZN(n1247) );
NAND2_X1 U1030 ( .A1(G214), .A2(n1325), .ZN(n1063) );
INV_X1 U1031 ( .A(n1079), .ZN(n1071) );
XNOR2_X1 U1032 ( .A(n1326), .B(n1198), .ZN(n1079) );
NAND2_X1 U1033 ( .A1(G210), .A2(n1325), .ZN(n1198) );
NAND2_X1 U1034 ( .A1(n1327), .A2(n1231), .ZN(n1325) );
INV_X1 U1035 ( .A(G237), .ZN(n1327) );
NAND3_X1 U1036 ( .A1(n1328), .A2(n1231), .A3(n1329), .ZN(n1326) );
XOR2_X1 U1037 ( .A(n1330), .B(KEYINPUT3), .Z(n1329) );
OR2_X1 U1038 ( .A1(n1196), .A2(n1195), .ZN(n1330) );
NAND2_X1 U1039 ( .A1(n1195), .A2(n1196), .ZN(n1328) );
XNOR2_X1 U1040 ( .A(n1331), .B(n1332), .ZN(n1196) );
XNOR2_X1 U1041 ( .A(G125), .B(n1333), .ZN(n1331) );
AND2_X1 U1042 ( .A1(n1049), .A2(G224), .ZN(n1333) );
XNOR2_X1 U1043 ( .A(n1145), .B(n1334), .ZN(n1195) );
NOR2_X1 U1044 ( .A1(KEYINPUT28), .A2(n1144), .ZN(n1334) );
XOR2_X1 U1045 ( .A(G110), .B(G122), .Z(n1144) );
XNOR2_X1 U1046 ( .A(n1335), .B(n1336), .ZN(n1145) );
NOR2_X1 U1047 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
AND3_X1 U1048 ( .A1(KEYINPUT18), .A2(n1339), .A3(G116), .ZN(n1338) );
NOR2_X1 U1049 ( .A1(KEYINPUT18), .A2(n1340), .ZN(n1337) );
XOR2_X1 U1050 ( .A(n1274), .B(n1190), .Z(n1335) );
INV_X1 U1051 ( .A(n1315), .ZN(n1190) );
XOR2_X1 U1052 ( .A(n1341), .B(n1342), .Z(n1315) );
XOR2_X1 U1053 ( .A(KEYINPUT36), .B(G107), .Z(n1342) );
XNOR2_X1 U1054 ( .A(G101), .B(G104), .ZN(n1341) );
INV_X1 U1055 ( .A(n1253), .ZN(n1082) );
NOR2_X1 U1056 ( .A1(n1271), .A2(n1064), .ZN(n1253) );
XNOR2_X1 U1057 ( .A(n1343), .B(n1151), .ZN(n1064) );
NAND2_X1 U1058 ( .A1(G217), .A2(n1303), .ZN(n1151) );
NAND2_X1 U1059 ( .A1(G234), .A2(n1231), .ZN(n1303) );
NAND2_X1 U1060 ( .A1(n1149), .A2(n1231), .ZN(n1343) );
XNOR2_X1 U1061 ( .A(n1344), .B(n1345), .ZN(n1149) );
XOR2_X1 U1062 ( .A(n1346), .B(n1347), .Z(n1345) );
XOR2_X1 U1063 ( .A(G128), .B(G110), .Z(n1347) );
NOR2_X1 U1064 ( .A1(KEYINPUT9), .A2(n1348), .ZN(n1346) );
XOR2_X1 U1065 ( .A(n1349), .B(n1287), .Z(n1348) );
XOR2_X1 U1066 ( .A(n1320), .B(KEYINPUT14), .Z(n1287) );
NAND2_X1 U1067 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
NAND2_X1 U1068 ( .A1(KEYINPUT20), .A2(n1113), .ZN(n1351) );
INV_X1 U1069 ( .A(n1283), .ZN(n1113) );
NAND2_X1 U1070 ( .A1(KEYINPUT32), .A2(n1283), .ZN(n1350) );
XOR2_X1 U1071 ( .A(G125), .B(G140), .Z(n1283) );
XOR2_X1 U1072 ( .A(n1352), .B(n1353), .Z(n1344) );
XOR2_X1 U1073 ( .A(n1354), .B(n1355), .Z(n1353) );
NAND2_X1 U1074 ( .A1(KEYINPUT57), .A2(n1339), .ZN(n1355) );
INV_X1 U1075 ( .A(G119), .ZN(n1339) );
NAND2_X1 U1076 ( .A1(G221), .A2(n1296), .ZN(n1354) );
AND2_X1 U1077 ( .A1(G234), .A2(n1049), .ZN(n1296) );
INV_X1 U1078 ( .A(G953), .ZN(n1049) );
NAND2_X1 U1079 ( .A1(n1356), .A2(n1357), .ZN(n1271) );
NAND2_X1 U1080 ( .A1(n1358), .A2(n1069), .ZN(n1357) );
XOR2_X1 U1081 ( .A(n1359), .B(KEYINPUT54), .Z(n1356) );
OR2_X1 U1082 ( .A1(n1069), .A2(n1358), .ZN(n1359) );
XNOR2_X1 U1083 ( .A(n1070), .B(KEYINPUT48), .ZN(n1358) );
NAND2_X1 U1084 ( .A1(n1360), .A2(n1231), .ZN(n1070) );
INV_X1 U1085 ( .A(G902), .ZN(n1231) );
XNOR2_X1 U1086 ( .A(n1361), .B(n1169), .ZN(n1360) );
XOR2_X1 U1087 ( .A(n1362), .B(G101), .Z(n1169) );
NAND2_X1 U1088 ( .A1(G210), .A2(n1284), .ZN(n1362) );
NOR2_X1 U1089 ( .A1(G953), .A2(G237), .ZN(n1284) );
XOR2_X1 U1090 ( .A(n1363), .B(KEYINPUT47), .Z(n1361) );
NAND2_X1 U1091 ( .A1(n1174), .A2(n1175), .ZN(n1363) );
NAND2_X1 U1092 ( .A1(n1364), .A2(n1365), .ZN(n1175) );
XOR2_X1 U1093 ( .A(G113), .B(n1340), .Z(n1365) );
XOR2_X1 U1094 ( .A(n1322), .B(n1332), .Z(n1364) );
INV_X1 U1095 ( .A(n1366), .ZN(n1332) );
NAND2_X1 U1096 ( .A1(n1367), .A2(n1368), .ZN(n1174) );
XOR2_X1 U1097 ( .A(n1322), .B(n1366), .Z(n1368) );
XOR2_X1 U1098 ( .A(n1369), .B(G128), .Z(n1366) );
NAND2_X1 U1099 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
NAND2_X1 U1100 ( .A1(G143), .A2(n1320), .ZN(n1371) );
XOR2_X1 U1101 ( .A(n1372), .B(KEYINPUT8), .Z(n1370) );
OR2_X1 U1102 ( .A1(n1320), .A2(G143), .ZN(n1372) );
INV_X1 U1103 ( .A(G146), .ZN(n1320) );
XOR2_X1 U1104 ( .A(n1122), .B(n1121), .Z(n1322) );
INV_X1 U1105 ( .A(G131), .ZN(n1121) );
XOR2_X1 U1106 ( .A(G134), .B(n1373), .Z(n1122) );
INV_X1 U1107 ( .A(n1352), .ZN(n1373) );
XNOR2_X1 U1108 ( .A(G137), .B(KEYINPUT59), .ZN(n1352) );
XOR2_X1 U1109 ( .A(n1274), .B(n1340), .Z(n1367) );
XOR2_X1 U1110 ( .A(G116), .B(G119), .Z(n1340) );
INV_X1 U1111 ( .A(G113), .ZN(n1274) );
INV_X1 U1112 ( .A(G472), .ZN(n1069) );
endmodule


