//Key = 1000111010011011110110000110111001011100111101010011100000101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362;

XOR2_X1 U760 ( .A(n1040), .B(n1041), .Z(G9) );
NOR2_X1 U761 ( .A1(n1042), .A2(n1043), .ZN(G75) );
NOR4_X1 U762 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
XOR2_X1 U763 ( .A(KEYINPUT54), .B(n1048), .Z(n1047) );
NOR4_X1 U764 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
INV_X1 U765 ( .A(n1053), .ZN(n1051) );
NAND2_X1 U766 ( .A1(n1054), .A2(n1055), .ZN(n1049) );
XOR2_X1 U767 ( .A(KEYINPUT22), .B(n1056), .Z(n1045) );
NOR3_X1 U768 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
NOR2_X1 U769 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR3_X1 U770 ( .A1(n1050), .A2(n1062), .A3(n1063), .ZN(n1061) );
NOR2_X1 U771 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U772 ( .A1(n1066), .A2(n1052), .ZN(n1065) );
XNOR2_X1 U773 ( .A(n1067), .B(KEYINPUT39), .ZN(n1066) );
NOR3_X1 U774 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1064) );
NOR3_X1 U775 ( .A1(n1052), .A2(n1071), .A3(n1070), .ZN(n1060) );
NOR2_X1 U776 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U777 ( .A1(n1063), .A2(n1074), .ZN(n1073) );
NOR3_X1 U778 ( .A1(n1050), .A2(n1075), .A3(n1076), .ZN(n1072) );
NAND3_X1 U779 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1044) );
NAND3_X1 U780 ( .A1(n1080), .A2(n1081), .A3(n1054), .ZN(n1079) );
INV_X1 U781 ( .A(n1057), .ZN(n1054) );
NAND2_X1 U782 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND3_X1 U783 ( .A1(n1084), .A2(n1053), .A3(n1085), .ZN(n1083) );
NAND2_X1 U784 ( .A1(n1086), .A2(n1087), .ZN(n1082) );
NAND2_X1 U785 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U786 ( .A1(n1085), .A2(n1090), .ZN(n1089) );
NAND2_X1 U787 ( .A1(n1053), .A2(n1091), .ZN(n1088) );
NOR3_X1 U788 ( .A1(n1092), .A2(G953), .A3(G952), .ZN(n1042) );
INV_X1 U789 ( .A(n1077), .ZN(n1092) );
NAND4_X1 U790 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1077) );
NOR4_X1 U791 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
XOR2_X1 U792 ( .A(KEYINPUT1), .B(n1076), .Z(n1100) );
XNOR2_X1 U793 ( .A(G469), .B(n1101), .ZN(n1099) );
XOR2_X1 U794 ( .A(KEYINPUT5), .B(n1102), .Z(n1098) );
NOR2_X1 U795 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U796 ( .A(KEYINPUT2), .B(n1105), .ZN(n1104) );
INV_X1 U797 ( .A(n1106), .ZN(n1103) );
NOR3_X1 U798 ( .A1(n1107), .A2(n1108), .A3(n1067), .ZN(n1095) );
INV_X1 U799 ( .A(n1068), .ZN(n1108) );
NOR2_X1 U800 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
AND2_X1 U801 ( .A1(n1111), .A2(KEYINPUT63), .ZN(n1110) );
NAND2_X1 U802 ( .A1(n1112), .A2(KEYINPUT63), .ZN(n1094) );
INV_X1 U803 ( .A(n1113), .ZN(n1112) );
XOR2_X1 U804 ( .A(n1114), .B(n1115), .Z(n1093) );
NAND2_X1 U805 ( .A1(KEYINPUT8), .A2(n1116), .ZN(n1115) );
XOR2_X1 U806 ( .A(n1117), .B(n1118), .Z(G72) );
NAND2_X1 U807 ( .A1(G953), .A2(n1119), .ZN(n1118) );
NAND2_X1 U808 ( .A1(G900), .A2(G227), .ZN(n1119) );
NAND2_X1 U809 ( .A1(KEYINPUT0), .A2(n1120), .ZN(n1117) );
XOR2_X1 U810 ( .A(n1121), .B(n1122), .Z(n1120) );
NAND2_X1 U811 ( .A1(n1078), .A2(n1123), .ZN(n1122) );
NAND3_X1 U812 ( .A1(n1124), .A2(n1125), .A3(KEYINPUT58), .ZN(n1121) );
NAND2_X1 U813 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U814 ( .A(n1128), .B(n1129), .Z(n1124) );
XOR2_X1 U815 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U816 ( .A1(KEYINPUT33), .A2(n1132), .ZN(n1130) );
XOR2_X1 U817 ( .A(n1133), .B(n1134), .Z(n1128) );
XNOR2_X1 U818 ( .A(G131), .B(n1135), .ZN(n1134) );
NOR2_X1 U819 ( .A1(G134), .A2(KEYINPUT44), .ZN(n1135) );
NAND2_X1 U820 ( .A1(KEYINPUT52), .A2(n1136), .ZN(n1133) );
XOR2_X1 U821 ( .A(n1137), .B(n1138), .Z(G69) );
NOR2_X1 U822 ( .A1(n1139), .A2(n1078), .ZN(n1138) );
NOR2_X1 U823 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U824 ( .A1(n1142), .A2(n1143), .ZN(n1137) );
NAND2_X1 U825 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U826 ( .A(KEYINPUT29), .B(n1146), .Z(n1142) );
NOR2_X1 U827 ( .A1(n1144), .A2(n1147), .ZN(n1146) );
XOR2_X1 U828 ( .A(n1145), .B(KEYINPUT32), .Z(n1147) );
NAND2_X1 U829 ( .A1(n1148), .A2(n1149), .ZN(n1145) );
NAND2_X1 U830 ( .A1(n1126), .A2(n1141), .ZN(n1149) );
AND2_X1 U831 ( .A1(n1150), .A2(n1078), .ZN(n1144) );
NAND2_X1 U832 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U833 ( .A1(n1153), .A2(n1154), .ZN(G66) );
XNOR2_X1 U834 ( .A(n1155), .B(n1156), .ZN(n1154) );
AND3_X1 U835 ( .A1(n1157), .A2(n1158), .A3(G217), .ZN(n1155) );
NOR2_X1 U836 ( .A1(n1153), .A2(n1159), .ZN(G63) );
XOR2_X1 U837 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U838 ( .A1(n1114), .A2(n1162), .ZN(n1161) );
INV_X1 U839 ( .A(G478), .ZN(n1114) );
NAND2_X1 U840 ( .A1(KEYINPUT36), .A2(n1163), .ZN(n1160) );
NOR3_X1 U841 ( .A1(n1153), .A2(n1164), .A3(n1165), .ZN(G60) );
AND4_X1 U842 ( .A1(n1166), .A2(KEYINPUT51), .A3(G475), .A4(n1157), .ZN(n1165) );
NOR2_X1 U843 ( .A1(n1166), .A2(n1167), .ZN(n1164) );
NOR3_X1 U844 ( .A1(n1162), .A2(n1168), .A3(n1169), .ZN(n1167) );
INV_X1 U845 ( .A(G475), .ZN(n1169) );
NOR2_X1 U846 ( .A1(KEYINPUT51), .A2(n1170), .ZN(n1168) );
NOR2_X1 U847 ( .A1(KEYINPUT27), .A2(n1171), .ZN(n1166) );
INV_X1 U848 ( .A(n1170), .ZN(n1171) );
XNOR2_X1 U849 ( .A(G104), .B(n1172), .ZN(G6) );
NOR2_X1 U850 ( .A1(n1153), .A2(n1173), .ZN(G57) );
XOR2_X1 U851 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U852 ( .A(n1176), .B(n1177), .ZN(n1175) );
NAND2_X1 U853 ( .A1(n1178), .A2(n1179), .ZN(n1176) );
NAND2_X1 U854 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U855 ( .A(n1182), .B(n1183), .Z(n1178) );
AND2_X1 U856 ( .A1(G472), .A2(n1157), .ZN(n1183) );
OR2_X1 U857 ( .A1(n1181), .A2(n1180), .ZN(n1182) );
XOR2_X1 U858 ( .A(n1184), .B(n1185), .Z(n1180) );
XNOR2_X1 U859 ( .A(n1186), .B(n1187), .ZN(n1185) );
INV_X1 U860 ( .A(KEYINPUT43), .ZN(n1181) );
XNOR2_X1 U861 ( .A(G101), .B(KEYINPUT20), .ZN(n1174) );
NOR2_X1 U862 ( .A1(n1153), .A2(n1188), .ZN(G54) );
XOR2_X1 U863 ( .A(n1189), .B(n1190), .Z(n1188) );
XNOR2_X1 U864 ( .A(n1191), .B(n1186), .ZN(n1190) );
AND2_X1 U865 ( .A1(G469), .A2(n1157), .ZN(n1191) );
INV_X1 U866 ( .A(n1162), .ZN(n1157) );
XOR2_X1 U867 ( .A(n1192), .B(n1193), .Z(n1189) );
XOR2_X1 U868 ( .A(n1194), .B(KEYINPUT24), .Z(n1193) );
NAND3_X1 U869 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1194) );
OR2_X1 U870 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NAND3_X1 U871 ( .A1(n1198), .A2(n1199), .A3(KEYINPUT14), .ZN(n1196) );
NOR2_X1 U872 ( .A1(KEYINPUT38), .A2(n1200), .ZN(n1198) );
NAND2_X1 U873 ( .A1(n1200), .A2(n1201), .ZN(n1195) );
INV_X1 U874 ( .A(KEYINPUT14), .ZN(n1201) );
XNOR2_X1 U875 ( .A(n1202), .B(KEYINPUT42), .ZN(n1200) );
NAND2_X1 U876 ( .A1(n1203), .A2(n1204), .ZN(n1192) );
NAND2_X1 U877 ( .A1(n1205), .A2(n1132), .ZN(n1204) );
XOR2_X1 U878 ( .A(KEYINPUT17), .B(n1206), .Z(n1203) );
NOR2_X1 U879 ( .A1(n1132), .A2(n1205), .ZN(n1206) );
NOR2_X1 U880 ( .A1(n1153), .A2(n1207), .ZN(G51) );
XOR2_X1 U881 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U882 ( .A(n1210), .B(n1148), .Z(n1209) );
NOR2_X1 U883 ( .A1(n1111), .A2(n1162), .ZN(n1210) );
NAND2_X1 U884 ( .A1(G902), .A2(n1046), .ZN(n1162) );
NAND3_X1 U885 ( .A1(n1211), .A2(n1151), .A3(n1212), .ZN(n1046) );
XNOR2_X1 U886 ( .A(n1152), .B(KEYINPUT28), .ZN(n1212) );
AND4_X1 U887 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1152) );
AND4_X1 U888 ( .A1(n1217), .A2(n1172), .A3(n1218), .A4(n1041), .ZN(n1151) );
NAND3_X1 U889 ( .A1(n1219), .A2(n1080), .A3(n1220), .ZN(n1041) );
NAND3_X1 U890 ( .A1(n1220), .A2(n1080), .A3(n1084), .ZN(n1172) );
NAND3_X1 U891 ( .A1(n1086), .A2(n1220), .A3(n1055), .ZN(n1217) );
INV_X1 U892 ( .A(n1123), .ZN(n1211) );
NAND4_X1 U893 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1123) );
AND4_X1 U894 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1224) );
NAND2_X1 U895 ( .A1(n1229), .A2(n1230), .ZN(n1223) );
NAND2_X1 U896 ( .A1(n1231), .A2(n1074), .ZN(n1230) );
XOR2_X1 U897 ( .A(KEYINPUT11), .B(n1084), .Z(n1231) );
INV_X1 U898 ( .A(n1232), .ZN(n1229) );
XOR2_X1 U899 ( .A(n1233), .B(n1234), .Z(n1208) );
XOR2_X1 U900 ( .A(KEYINPUT59), .B(n1235), .Z(n1234) );
NOR2_X1 U901 ( .A1(KEYINPUT49), .A2(n1236), .ZN(n1233) );
XNOR2_X1 U902 ( .A(n1187), .B(G125), .ZN(n1236) );
NOR2_X1 U903 ( .A1(n1078), .A2(G952), .ZN(n1153) );
XNOR2_X1 U904 ( .A(G146), .B(n1221), .ZN(G48) );
NAND2_X1 U905 ( .A1(n1237), .A2(n1084), .ZN(n1221) );
XOR2_X1 U906 ( .A(n1238), .B(n1222), .Z(G45) );
NAND4_X1 U907 ( .A1(n1091), .A2(n1090), .A3(n1055), .A4(n1239), .ZN(n1222) );
NOR3_X1 U908 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1239) );
XNOR2_X1 U909 ( .A(G140), .B(n1228), .ZN(G42) );
NAND4_X1 U910 ( .A1(n1085), .A2(n1243), .A3(n1244), .A4(n1084), .ZN(n1228) );
XNOR2_X1 U911 ( .A(G137), .B(n1227), .ZN(G39) );
NAND4_X1 U912 ( .A1(n1086), .A2(n1085), .A3(n1243), .A4(n1076), .ZN(n1227) );
XOR2_X1 U913 ( .A(G134), .B(n1245), .Z(G36) );
NOR2_X1 U914 ( .A1(n1074), .A2(n1232), .ZN(n1245) );
XOR2_X1 U915 ( .A(G131), .B(n1246), .Z(G33) );
NOR2_X1 U916 ( .A1(n1247), .A2(n1232), .ZN(n1246) );
NAND4_X1 U917 ( .A1(n1055), .A2(n1085), .A3(n1090), .A4(n1248), .ZN(n1232) );
INV_X1 U918 ( .A(n1052), .ZN(n1085) );
NAND2_X1 U919 ( .A1(n1249), .A2(n1068), .ZN(n1052) );
XOR2_X1 U920 ( .A(n1069), .B(KEYINPUT60), .Z(n1249) );
XOR2_X1 U921 ( .A(n1250), .B(n1226), .Z(G30) );
NAND2_X1 U922 ( .A1(n1237), .A2(n1219), .ZN(n1226) );
AND3_X1 U923 ( .A1(n1091), .A2(n1076), .A3(n1243), .ZN(n1237) );
AND3_X1 U924 ( .A1(n1248), .A2(n1251), .A3(n1090), .ZN(n1243) );
XNOR2_X1 U925 ( .A(G101), .B(n1252), .ZN(G3) );
NAND3_X1 U926 ( .A1(n1086), .A2(n1220), .A3(n1253), .ZN(n1252) );
XNOR2_X1 U927 ( .A(n1055), .B(KEYINPUT26), .ZN(n1253) );
XNOR2_X1 U928 ( .A(G125), .B(n1225), .ZN(G27) );
NAND4_X1 U929 ( .A1(n1244), .A2(n1053), .A3(n1084), .A4(n1254), .ZN(n1225) );
NOR3_X1 U930 ( .A1(n1255), .A2(n1075), .A3(n1241), .ZN(n1254) );
INV_X1 U931 ( .A(n1248), .ZN(n1241) );
NAND2_X1 U932 ( .A1(n1057), .A2(n1256), .ZN(n1248) );
NAND4_X1 U933 ( .A1(G902), .A2(n1126), .A3(n1257), .A4(n1127), .ZN(n1256) );
INV_X1 U934 ( .A(G900), .ZN(n1127) );
XNOR2_X1 U935 ( .A(G122), .B(n1213), .ZN(G24) );
NAND4_X1 U936 ( .A1(n1258), .A2(n1080), .A3(n1097), .A4(n1259), .ZN(n1213) );
INV_X1 U937 ( .A(n1063), .ZN(n1080) );
NAND2_X1 U938 ( .A1(n1075), .A2(n1244), .ZN(n1063) );
INV_X1 U939 ( .A(n1251), .ZN(n1075) );
XNOR2_X1 U940 ( .A(G119), .B(n1214), .ZN(G21) );
NAND4_X1 U941 ( .A1(n1258), .A2(n1086), .A3(n1076), .A4(n1251), .ZN(n1214) );
INV_X1 U942 ( .A(n1244), .ZN(n1076) );
XNOR2_X1 U943 ( .A(G116), .B(n1215), .ZN(G18) );
NAND3_X1 U944 ( .A1(n1055), .A2(n1219), .A3(n1258), .ZN(n1215) );
INV_X1 U945 ( .A(n1074), .ZN(n1219) );
NAND2_X1 U946 ( .A1(n1240), .A2(n1259), .ZN(n1074) );
INV_X1 U947 ( .A(n1242), .ZN(n1259) );
XOR2_X1 U948 ( .A(n1260), .B(n1261), .Z(G15) );
NAND2_X1 U949 ( .A1(KEYINPUT47), .A2(n1262), .ZN(n1261) );
INV_X1 U950 ( .A(n1216), .ZN(n1262) );
NAND3_X1 U951 ( .A1(n1055), .A2(n1084), .A3(n1258), .ZN(n1216) );
AND3_X1 U952 ( .A1(n1091), .A2(n1263), .A3(n1053), .ZN(n1258) );
NOR2_X1 U953 ( .A1(n1070), .A2(n1059), .ZN(n1053) );
INV_X1 U954 ( .A(n1247), .ZN(n1084) );
NAND2_X1 U955 ( .A1(n1242), .A2(n1097), .ZN(n1247) );
INV_X1 U956 ( .A(n1240), .ZN(n1097) );
NOR2_X1 U957 ( .A1(n1251), .A2(n1244), .ZN(n1055) );
XOR2_X1 U958 ( .A(n1264), .B(n1218), .Z(G12) );
NAND4_X1 U959 ( .A1(n1086), .A2(n1220), .A3(n1244), .A4(n1251), .ZN(n1218) );
NAND2_X1 U960 ( .A1(n1106), .A2(n1105), .ZN(n1251) );
NAND3_X1 U961 ( .A1(n1265), .A2(n1266), .A3(n1156), .ZN(n1105) );
NAND2_X1 U962 ( .A1(G217), .A2(n1158), .ZN(n1265) );
NAND3_X1 U963 ( .A1(n1267), .A2(n1158), .A3(G217), .ZN(n1106) );
NAND2_X1 U964 ( .A1(n1156), .A2(n1266), .ZN(n1267) );
XOR2_X1 U965 ( .A(n1268), .B(n1269), .Z(n1156) );
XOR2_X1 U966 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U967 ( .A(n1272), .B(n1273), .Z(n1271) );
NAND2_X1 U968 ( .A1(KEYINPUT50), .A2(G119), .ZN(n1273) );
NAND2_X1 U969 ( .A1(n1274), .A2(G221), .ZN(n1272) );
XOR2_X1 U970 ( .A(n1275), .B(n1276), .Z(n1268) );
NOR2_X1 U971 ( .A1(KEYINPUT46), .A2(n1277), .ZN(n1276) );
XOR2_X1 U972 ( .A(n1264), .B(G128), .Z(n1275) );
XOR2_X1 U973 ( .A(n1278), .B(G472), .Z(n1244) );
NAND2_X1 U974 ( .A1(n1279), .A2(n1266), .ZN(n1278) );
XOR2_X1 U975 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U976 ( .A(n1187), .B(n1282), .ZN(n1281) );
NOR2_X1 U977 ( .A1(KEYINPUT10), .A2(n1184), .ZN(n1282) );
XNOR2_X1 U978 ( .A(n1283), .B(n1284), .ZN(n1184) );
NAND2_X1 U979 ( .A1(KEYINPUT4), .A2(n1260), .ZN(n1283) );
INV_X1 U980 ( .A(G113), .ZN(n1260) );
XOR2_X1 U981 ( .A(n1285), .B(n1286), .Z(n1280) );
NOR2_X1 U982 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XOR2_X1 U983 ( .A(n1289), .B(KEYINPUT25), .Z(n1288) );
NAND2_X1 U984 ( .A1(G101), .A2(n1290), .ZN(n1289) );
NOR2_X1 U985 ( .A1(G101), .A2(n1290), .ZN(n1287) );
XNOR2_X1 U986 ( .A(KEYINPUT55), .B(n1177), .ZN(n1290) );
NAND2_X1 U987 ( .A1(n1291), .A2(G210), .ZN(n1177) );
NAND2_X1 U988 ( .A1(KEYINPUT45), .A2(n1186), .ZN(n1285) );
AND3_X1 U989 ( .A1(n1090), .A2(n1263), .A3(n1091), .ZN(n1220) );
INV_X1 U990 ( .A(n1255), .ZN(n1091) );
NAND2_X1 U991 ( .A1(n1068), .A2(n1069), .ZN(n1255) );
NAND2_X1 U992 ( .A1(n1292), .A2(n1113), .ZN(n1069) );
NAND2_X1 U993 ( .A1(n1109), .A2(n1111), .ZN(n1113) );
OR2_X1 U994 ( .A1(n1111), .A2(n1109), .ZN(n1292) );
AND2_X1 U995 ( .A1(n1293), .A2(n1266), .ZN(n1109) );
XOR2_X1 U996 ( .A(n1294), .B(n1148), .Z(n1293) );
XNOR2_X1 U997 ( .A(n1295), .B(n1296), .ZN(n1148) );
XOR2_X1 U998 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U999 ( .A(n1299), .B(n1300), .Z(n1298) );
NOR2_X1 U1000 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
XOR2_X1 U1001 ( .A(n1303), .B(KEYINPUT35), .Z(n1302) );
NAND2_X1 U1002 ( .A1(G113), .A2(n1284), .ZN(n1303) );
NOR2_X1 U1003 ( .A1(G113), .A2(n1284), .ZN(n1301) );
XOR2_X1 U1004 ( .A(G116), .B(G119), .Z(n1284) );
NAND2_X1 U1005 ( .A1(KEYINPUT30), .A2(n1264), .ZN(n1299) );
NAND2_X1 U1006 ( .A1(n1304), .A2(n1305), .ZN(n1297) );
OR2_X1 U1007 ( .A1(n1306), .A2(KEYINPUT31), .ZN(n1305) );
NAND3_X1 U1008 ( .A1(G104), .A2(n1040), .A3(KEYINPUT31), .ZN(n1304) );
XNOR2_X1 U1009 ( .A(G101), .B(n1307), .ZN(n1295) );
XOR2_X1 U1010 ( .A(KEYINPUT34), .B(G122), .Z(n1307) );
NOR2_X1 U1011 ( .A1(KEYINPUT9), .A2(n1308), .ZN(n1294) );
XOR2_X1 U1012 ( .A(n1309), .B(n1310), .Z(n1308) );
NOR2_X1 U1013 ( .A1(KEYINPUT18), .A2(n1187), .ZN(n1310) );
XNOR2_X1 U1014 ( .A(n1250), .B(n1311), .ZN(n1187) );
XOR2_X1 U1015 ( .A(G146), .B(G143), .Z(n1311) );
XNOR2_X1 U1016 ( .A(G125), .B(n1235), .ZN(n1309) );
NOR2_X1 U1017 ( .A1(n1140), .A2(G953), .ZN(n1235) );
INV_X1 U1018 ( .A(G224), .ZN(n1140) );
NAND2_X1 U1019 ( .A1(G210), .A2(n1312), .ZN(n1111) );
NAND2_X1 U1020 ( .A1(G214), .A2(n1312), .ZN(n1068) );
NAND2_X1 U1021 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
INV_X1 U1022 ( .A(G237), .ZN(n1314) );
NAND2_X1 U1023 ( .A1(n1057), .A2(n1315), .ZN(n1263) );
NAND4_X1 U1024 ( .A1(n1316), .A2(n1126), .A3(n1257), .A4(n1141), .ZN(n1315) );
INV_X1 U1025 ( .A(G898), .ZN(n1141) );
XOR2_X1 U1026 ( .A(G953), .B(KEYINPUT13), .Z(n1126) );
XOR2_X1 U1027 ( .A(n1266), .B(KEYINPUT16), .Z(n1316) );
NAND3_X1 U1028 ( .A1(n1257), .A2(n1078), .A3(G952), .ZN(n1057) );
NAND2_X1 U1029 ( .A1(G237), .A2(G234), .ZN(n1257) );
NOR2_X1 U1030 ( .A1(n1070), .A2(n1317), .ZN(n1090) );
INV_X1 U1031 ( .A(n1059), .ZN(n1317) );
XOR2_X1 U1032 ( .A(n1101), .B(n1318), .Z(n1059) );
NOR2_X1 U1033 ( .A1(G469), .A2(KEYINPUT48), .ZN(n1318) );
NAND2_X1 U1034 ( .A1(n1319), .A2(n1266), .ZN(n1101) );
XOR2_X1 U1035 ( .A(n1320), .B(n1321), .Z(n1319) );
XNOR2_X1 U1036 ( .A(n1132), .B(n1322), .ZN(n1321) );
XNOR2_X1 U1037 ( .A(n1199), .B(KEYINPUT23), .ZN(n1322) );
AND2_X1 U1038 ( .A1(G227), .A2(n1078), .ZN(n1199) );
AND2_X1 U1039 ( .A1(n1323), .A2(n1324), .ZN(n1132) );
NAND2_X1 U1040 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NAND2_X1 U1041 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
NAND2_X1 U1042 ( .A1(KEYINPUT15), .A2(n1250), .ZN(n1328) );
INV_X1 U1043 ( .A(KEYINPUT53), .ZN(n1327) );
NAND2_X1 U1044 ( .A1(G128), .A2(n1329), .ZN(n1323) );
NAND2_X1 U1045 ( .A1(KEYINPUT15), .A2(n1330), .ZN(n1329) );
OR2_X1 U1046 ( .A1(n1325), .A2(KEYINPUT53), .ZN(n1330) );
XNOR2_X1 U1047 ( .A(n1331), .B(n1332), .ZN(n1325) );
XOR2_X1 U1048 ( .A(KEYINPUT62), .B(G146), .Z(n1332) );
NAND2_X1 U1049 ( .A1(KEYINPUT19), .A2(n1333), .ZN(n1331) );
XOR2_X1 U1050 ( .A(KEYINPUT3), .B(G143), .Z(n1333) );
XOR2_X1 U1051 ( .A(n1205), .B(n1334), .Z(n1320) );
XNOR2_X1 U1052 ( .A(n1186), .B(n1202), .ZN(n1334) );
XNOR2_X1 U1053 ( .A(n1264), .B(n1335), .ZN(n1202) );
XOR2_X1 U1054 ( .A(n1336), .B(G131), .Z(n1186) );
NAND2_X1 U1055 ( .A1(KEYINPUT37), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1056 ( .A(n1270), .B(n1338), .Z(n1337) );
XOR2_X1 U1057 ( .A(KEYINPUT7), .B(G134), .Z(n1338) );
INV_X1 U1058 ( .A(n1131), .ZN(n1270) );
XNOR2_X1 U1059 ( .A(G137), .B(KEYINPUT40), .ZN(n1131) );
XNOR2_X1 U1060 ( .A(G101), .B(n1306), .ZN(n1205) );
XOR2_X1 U1061 ( .A(G104), .B(G107), .Z(n1306) );
XOR2_X1 U1062 ( .A(n1067), .B(KEYINPUT56), .Z(n1070) );
AND2_X1 U1063 ( .A1(G221), .A2(n1158), .ZN(n1067) );
NAND2_X1 U1064 ( .A1(G234), .A2(n1313), .ZN(n1158) );
XOR2_X1 U1065 ( .A(n1266), .B(KEYINPUT61), .Z(n1313) );
INV_X1 U1066 ( .A(n1050), .ZN(n1086) );
NAND2_X1 U1067 ( .A1(n1242), .A2(n1240), .ZN(n1050) );
XOR2_X1 U1068 ( .A(n1339), .B(G475), .Z(n1240) );
NAND2_X1 U1069 ( .A1(n1170), .A2(n1266), .ZN(n1339) );
XOR2_X1 U1070 ( .A(n1340), .B(n1341), .Z(n1170) );
XOR2_X1 U1071 ( .A(G122), .B(G113), .Z(n1341) );
XOR2_X1 U1072 ( .A(n1342), .B(G104), .Z(n1340) );
NAND3_X1 U1073 ( .A1(n1343), .A2(n1344), .A3(KEYINPUT41), .ZN(n1342) );
NAND2_X1 U1074 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
NAND2_X1 U1075 ( .A1(KEYINPUT12), .A2(n1347), .ZN(n1346) );
OR2_X1 U1076 ( .A1(n1277), .A2(KEYINPUT21), .ZN(n1347) );
NAND2_X1 U1077 ( .A1(n1277), .A2(n1348), .ZN(n1343) );
NAND2_X1 U1078 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1079 ( .A1(KEYINPUT12), .A2(n1351), .ZN(n1350) );
INV_X1 U1080 ( .A(n1345), .ZN(n1351) );
XOR2_X1 U1081 ( .A(n1352), .B(n1353), .Z(n1345) );
XOR2_X1 U1082 ( .A(G143), .B(G131), .Z(n1353) );
NAND2_X1 U1083 ( .A1(n1291), .A2(G214), .ZN(n1352) );
NOR2_X1 U1084 ( .A1(G953), .A2(G237), .ZN(n1291) );
INV_X1 U1085 ( .A(KEYINPUT21), .ZN(n1349) );
XNOR2_X1 U1086 ( .A(n1136), .B(G146), .ZN(n1277) );
XNOR2_X1 U1087 ( .A(G125), .B(n1335), .ZN(n1136) );
XOR2_X1 U1088 ( .A(G140), .B(KEYINPUT6), .Z(n1335) );
XOR2_X1 U1089 ( .A(n1116), .B(G478), .Z(n1242) );
NAND2_X1 U1090 ( .A1(n1163), .A2(n1266), .ZN(n1116) );
INV_X1 U1091 ( .A(G902), .ZN(n1266) );
XOR2_X1 U1092 ( .A(n1354), .B(n1355), .Z(n1163) );
XOR2_X1 U1093 ( .A(G116), .B(n1356), .Z(n1355) );
XOR2_X1 U1094 ( .A(G134), .B(G122), .Z(n1356) );
XOR2_X1 U1095 ( .A(n1357), .B(n1358), .Z(n1354) );
XOR2_X1 U1096 ( .A(n1040), .B(n1359), .Z(n1358) );
NAND2_X1 U1097 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NAND2_X1 U1098 ( .A1(G128), .A2(n1238), .ZN(n1361) );
INV_X1 U1099 ( .A(G143), .ZN(n1238) );
XOR2_X1 U1100 ( .A(n1362), .B(KEYINPUT57), .Z(n1360) );
NAND2_X1 U1101 ( .A1(G143), .A2(n1250), .ZN(n1362) );
INV_X1 U1102 ( .A(G128), .ZN(n1250) );
INV_X1 U1103 ( .A(G107), .ZN(n1040) );
NAND2_X1 U1104 ( .A1(G217), .A2(n1274), .ZN(n1357) );
AND2_X1 U1105 ( .A1(G234), .A2(n1078), .ZN(n1274) );
INV_X1 U1106 ( .A(G953), .ZN(n1078) );
INV_X1 U1107 ( .A(G110), .ZN(n1264) );
endmodule


