//Key = 1001110101100111110011011101011100110001110111001010000000100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395;

XNOR2_X1 U760 ( .A(n1063), .B(n1064), .ZN(G9) );
NOR2_X1 U761 ( .A1(KEYINPUT53), .A2(n1065), .ZN(n1064) );
NOR2_X1 U762 ( .A1(n1066), .A2(n1067), .ZN(G75) );
XOR2_X1 U763 ( .A(KEYINPUT47), .B(n1068), .Z(n1067) );
NOR4_X1 U764 ( .A1(G953), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1068) );
XOR2_X1 U765 ( .A(KEYINPUT48), .B(n1072), .Z(n1071) );
NOR2_X1 U766 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR4_X1 U767 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
INV_X1 U768 ( .A(n1079), .ZN(n1077) );
NOR2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(n1075) );
NOR2_X1 U770 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U771 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NOR2_X1 U772 ( .A1(n1086), .A2(n1087), .ZN(n1080) );
NOR3_X1 U773 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1086) );
NOR3_X1 U774 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
INV_X1 U775 ( .A(KEYINPUT41), .ZN(n1091) );
NOR2_X1 U776 ( .A1(KEYINPUT41), .A2(n1083), .ZN(n1089) );
NOR4_X1 U777 ( .A1(n1094), .A2(n1087), .A3(n1083), .A4(n1078), .ZN(n1073) );
INV_X1 U778 ( .A(n1095), .ZN(n1087) );
NOR2_X1 U779 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
AND2_X1 U780 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR3_X1 U781 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1096) );
NOR3_X1 U782 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
NOR2_X1 U783 ( .A1(n1099), .A2(n1106), .ZN(n1101) );
NOR3_X1 U784 ( .A1(n1069), .A2(G953), .A3(G952), .ZN(n1066) );
AND4_X1 U785 ( .A1(n1107), .A2(n1108), .A3(n1109), .A4(n1110), .ZN(n1069) );
NOR4_X1 U786 ( .A1(n1103), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1110) );
XOR2_X1 U787 ( .A(n1114), .B(n1115), .Z(n1112) );
NAND2_X1 U788 ( .A1(KEYINPUT30), .A2(n1116), .ZN(n1114) );
NOR3_X1 U789 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1111) );
NOR2_X1 U790 ( .A1(KEYINPUT61), .A2(n1120), .ZN(n1119) );
NOR4_X1 U791 ( .A1(n1121), .A2(n1122), .A3(KEYINPUT42), .A4(G469), .ZN(n1118) );
INV_X1 U792 ( .A(KEYINPUT61), .ZN(n1122) );
NOR2_X1 U793 ( .A1(n1123), .A2(n1124), .ZN(n1117) );
INV_X1 U794 ( .A(G469), .ZN(n1124) );
NOR2_X1 U795 ( .A1(KEYINPUT42), .A2(n1121), .ZN(n1123) );
XNOR2_X1 U796 ( .A(n1125), .B(G478), .ZN(n1109) );
XNOR2_X1 U797 ( .A(n1126), .B(KEYINPUT8), .ZN(n1107) );
XOR2_X1 U798 ( .A(n1127), .B(n1128), .Z(G72) );
NOR2_X1 U799 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR3_X1 U800 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1130) );
NOR2_X1 U801 ( .A1(G953), .A2(n1134), .ZN(n1129) );
NOR2_X1 U802 ( .A1(n1135), .A2(n1136), .ZN(n1127) );
XOR2_X1 U803 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U804 ( .A(G134), .B(n1139), .Z(n1138) );
XNOR2_X1 U805 ( .A(n1140), .B(G137), .ZN(n1139) );
XOR2_X1 U806 ( .A(n1141), .B(n1142), .Z(n1137) );
XNOR2_X1 U807 ( .A(G131), .B(n1143), .ZN(n1142) );
NOR2_X1 U808 ( .A1(n1131), .A2(n1144), .ZN(n1135) );
XNOR2_X1 U809 ( .A(KEYINPUT37), .B(n1133), .ZN(n1144) );
INV_X1 U810 ( .A(G900), .ZN(n1133) );
XOR2_X1 U811 ( .A(n1145), .B(n1146), .Z(G69) );
XOR2_X1 U812 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U813 ( .A1(n1149), .A2(n1131), .ZN(n1148) );
NOR2_X1 U814 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND2_X1 U815 ( .A1(n1152), .A2(n1153), .ZN(n1147) );
NAND2_X1 U816 ( .A1(G953), .A2(n1151), .ZN(n1153) );
XOR2_X1 U817 ( .A(n1154), .B(n1155), .Z(n1152) );
XNOR2_X1 U818 ( .A(n1156), .B(n1157), .ZN(n1155) );
XNOR2_X1 U819 ( .A(KEYINPUT5), .B(n1158), .ZN(n1154) );
NOR2_X1 U820 ( .A1(KEYINPUT52), .A2(n1159), .ZN(n1158) );
NAND2_X1 U821 ( .A1(n1131), .A2(n1160), .ZN(n1145) );
NOR2_X1 U822 ( .A1(n1161), .A2(n1162), .ZN(G66) );
NOR3_X1 U823 ( .A1(n1115), .A2(n1163), .A3(n1164), .ZN(n1162) );
NOR3_X1 U824 ( .A1(n1165), .A2(n1116), .A3(n1166), .ZN(n1164) );
INV_X1 U825 ( .A(n1167), .ZN(n1166) );
NOR2_X1 U826 ( .A1(n1168), .A2(n1169), .ZN(n1163) );
NOR2_X1 U827 ( .A1(n1170), .A2(n1116), .ZN(n1168) );
NOR2_X1 U828 ( .A1(n1161), .A2(n1171), .ZN(G63) );
NOR3_X1 U829 ( .A1(n1125), .A2(n1172), .A3(n1173), .ZN(n1171) );
NOR3_X1 U830 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1173) );
AND2_X1 U831 ( .A1(n1174), .A2(n1175), .ZN(n1172) );
NAND3_X1 U832 ( .A1(G478), .A2(n1070), .A3(KEYINPUT34), .ZN(n1174) );
NOR2_X1 U833 ( .A1(n1161), .A2(n1177), .ZN(G60) );
XNOR2_X1 U834 ( .A(n1178), .B(n1179), .ZN(n1177) );
NAND2_X1 U835 ( .A1(n1167), .A2(G475), .ZN(n1178) );
XNOR2_X1 U836 ( .A(G104), .B(n1180), .ZN(G6) );
NOR2_X1 U837 ( .A1(n1161), .A2(n1181), .ZN(G57) );
XNOR2_X1 U838 ( .A(n1182), .B(n1183), .ZN(n1181) );
NOR3_X1 U839 ( .A1(n1184), .A2(n1176), .A3(n1185), .ZN(n1183) );
XNOR2_X1 U840 ( .A(KEYINPUT46), .B(n1070), .ZN(n1184) );
INV_X1 U841 ( .A(n1170), .ZN(n1070) );
NOR2_X1 U842 ( .A1(n1161), .A2(n1186), .ZN(G54) );
XNOR2_X1 U843 ( .A(n1187), .B(n1188), .ZN(n1186) );
NAND2_X1 U844 ( .A1(n1167), .A2(G469), .ZN(n1187) );
NOR2_X1 U845 ( .A1(n1131), .A2(G952), .ZN(n1161) );
NOR2_X1 U846 ( .A1(n1189), .A2(n1190), .ZN(G51) );
XOR2_X1 U847 ( .A(n1191), .B(n1192), .Z(n1190) );
NAND2_X1 U848 ( .A1(n1167), .A2(n1193), .ZN(n1192) );
NOR2_X1 U849 ( .A1(n1176), .A2(n1170), .ZN(n1167) );
NOR2_X1 U850 ( .A1(n1160), .A2(n1134), .ZN(n1170) );
NAND4_X1 U851 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1134) );
NOR4_X1 U852 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
AND4_X1 U853 ( .A1(n1113), .A2(n1202), .A3(n1085), .A4(n1203), .ZN(n1200) );
NOR3_X1 U854 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1199) );
NOR2_X1 U855 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
INV_X1 U856 ( .A(KEYINPUT26), .ZN(n1208) );
AND4_X1 U857 ( .A1(n1078), .A2(n1209), .A3(n1098), .A4(n1108), .ZN(n1207) );
NOR2_X1 U858 ( .A1(KEYINPUT26), .A2(n1210), .ZN(n1205) );
INV_X1 U859 ( .A(n1211), .ZN(n1204) );
NOR3_X1 U860 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1196) );
NOR2_X1 U861 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND4_X1 U862 ( .A1(n1217), .A2(n1105), .A3(n1079), .A4(n1218), .ZN(n1216) );
INV_X1 U863 ( .A(KEYINPUT22), .ZN(n1215) );
NOR2_X1 U864 ( .A1(KEYINPUT22), .A2(n1219), .ZN(n1213) );
INV_X1 U865 ( .A(n1220), .ZN(n1212) );
NAND4_X1 U866 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1160) );
AND4_X1 U867 ( .A1(n1065), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1224) );
NAND3_X1 U868 ( .A1(n1104), .A2(n1095), .A3(n1228), .ZN(n1065) );
AND2_X1 U869 ( .A1(n1229), .A2(n1180), .ZN(n1223) );
NAND3_X1 U870 ( .A1(n1228), .A2(n1095), .A3(n1105), .ZN(n1180) );
NAND3_X1 U871 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1222) );
XNOR2_X1 U872 ( .A(KEYINPUT51), .B(n1076), .ZN(n1231) );
NAND4_X1 U873 ( .A1(n1104), .A2(n1233), .A3(n1079), .A4(n1234), .ZN(n1221) );
NOR2_X1 U874 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XOR2_X1 U875 ( .A(KEYINPUT29), .B(n1088), .Z(n1236) );
NAND2_X1 U876 ( .A1(n1237), .A2(n1238), .ZN(n1191) );
NAND2_X1 U877 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
XOR2_X1 U878 ( .A(n1241), .B(KEYINPUT19), .Z(n1237) );
OR2_X1 U879 ( .A1(n1240), .A2(n1239), .ZN(n1241) );
XNOR2_X1 U880 ( .A(n1242), .B(KEYINPUT16), .ZN(n1240) );
NOR2_X1 U881 ( .A1(G952), .A2(n1243), .ZN(n1189) );
XNOR2_X1 U882 ( .A(G953), .B(KEYINPUT18), .ZN(n1243) );
XNOR2_X1 U883 ( .A(G146), .B(n1220), .ZN(G48) );
NAND3_X1 U884 ( .A1(n1232), .A2(n1105), .A3(n1203), .ZN(n1220) );
XNOR2_X1 U885 ( .A(G143), .B(n1244), .ZN(G45) );
NAND4_X1 U886 ( .A1(n1245), .A2(n1203), .A3(n1202), .A4(n1113), .ZN(n1244) );
XNOR2_X1 U887 ( .A(n1085), .B(KEYINPUT4), .ZN(n1245) );
XNOR2_X1 U888 ( .A(G140), .B(n1246), .ZN(G42) );
NAND2_X1 U889 ( .A1(n1211), .A2(n1210), .ZN(n1246) );
XNOR2_X1 U890 ( .A(G137), .B(n1194), .ZN(G39) );
NAND2_X1 U891 ( .A1(n1247), .A2(n1210), .ZN(n1194) );
XOR2_X1 U892 ( .A(G134), .B(n1198), .Z(G36) );
AND3_X1 U893 ( .A1(n1085), .A2(n1104), .A3(n1210), .ZN(n1198) );
XNOR2_X1 U894 ( .A(G131), .B(n1195), .ZN(G33) );
NAND3_X1 U895 ( .A1(n1105), .A2(n1085), .A3(n1210), .ZN(n1195) );
AND3_X1 U896 ( .A1(n1098), .A2(n1248), .A3(n1108), .ZN(n1210) );
INV_X1 U897 ( .A(n1083), .ZN(n1108) );
NAND2_X1 U898 ( .A1(n1249), .A2(n1093), .ZN(n1083) );
INV_X1 U899 ( .A(n1092), .ZN(n1249) );
INV_X1 U900 ( .A(n1250), .ZN(n1105) );
XNOR2_X1 U901 ( .A(n1201), .B(n1251), .ZN(G30) );
XOR2_X1 U902 ( .A(KEYINPUT50), .B(G128), .Z(n1251) );
AND3_X1 U903 ( .A1(n1232), .A2(n1104), .A3(n1203), .ZN(n1201) );
AND2_X1 U904 ( .A1(n1217), .A2(n1098), .ZN(n1203) );
INV_X1 U905 ( .A(n1252), .ZN(n1104) );
NAND3_X1 U906 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(G3) );
OR2_X1 U907 ( .A1(n1256), .A2(n1229), .ZN(n1255) );
NAND3_X1 U908 ( .A1(n1229), .A2(n1256), .A3(G101), .ZN(n1254) );
NAND2_X1 U909 ( .A1(n1257), .A2(n1258), .ZN(n1253) );
NAND2_X1 U910 ( .A1(n1259), .A2(n1256), .ZN(n1257) );
INV_X1 U911 ( .A(KEYINPUT28), .ZN(n1256) );
XNOR2_X1 U912 ( .A(KEYINPUT25), .B(n1229), .ZN(n1259) );
NAND3_X1 U913 ( .A1(n1099), .A2(n1228), .A3(n1085), .ZN(n1229) );
XOR2_X1 U914 ( .A(n1219), .B(n1260), .Z(G27) );
XNOR2_X1 U915 ( .A(KEYINPUT45), .B(n1261), .ZN(n1260) );
NAND3_X1 U916 ( .A1(n1211), .A2(n1079), .A3(n1217), .ZN(n1219) );
AND2_X1 U917 ( .A1(n1088), .A2(n1248), .ZN(n1217) );
NAND2_X1 U918 ( .A1(n1078), .A2(n1209), .ZN(n1248) );
NAND4_X1 U919 ( .A1(n1262), .A2(G953), .A3(G902), .A4(n1263), .ZN(n1209) );
XNOR2_X1 U920 ( .A(G900), .B(KEYINPUT37), .ZN(n1262) );
NOR2_X1 U921 ( .A1(n1250), .A2(n1218), .ZN(n1211) );
XNOR2_X1 U922 ( .A(G122), .B(n1227), .ZN(G24) );
NAND4_X1 U923 ( .A1(n1202), .A2(n1230), .A3(n1095), .A4(n1113), .ZN(n1227) );
NAND2_X1 U924 ( .A1(n1264), .A2(n1265), .ZN(n1095) );
OR3_X1 U925 ( .A1(n1266), .A2(n1126), .A3(KEYINPUT55), .ZN(n1265) );
NAND2_X1 U926 ( .A1(KEYINPUT55), .A2(n1084), .ZN(n1264) );
XNOR2_X1 U927 ( .A(G119), .B(n1267), .ZN(G21) );
NAND2_X1 U928 ( .A1(n1247), .A2(n1230), .ZN(n1267) );
AND2_X1 U929 ( .A1(n1232), .A2(n1099), .ZN(n1247) );
AND2_X1 U930 ( .A1(n1126), .A2(n1266), .ZN(n1232) );
XOR2_X1 U931 ( .A(G116), .B(n1268), .Z(G18) );
NOR2_X1 U932 ( .A1(n1252), .A2(n1269), .ZN(n1268) );
NAND2_X1 U933 ( .A1(n1202), .A2(n1270), .ZN(n1252) );
XOR2_X1 U934 ( .A(n1271), .B(KEYINPUT17), .Z(n1202) );
XNOR2_X1 U935 ( .A(G113), .B(n1226), .ZN(G15) );
OR2_X1 U936 ( .A1(n1250), .A2(n1269), .ZN(n1226) );
NAND2_X1 U937 ( .A1(n1230), .A2(n1085), .ZN(n1269) );
INV_X1 U938 ( .A(n1235), .ZN(n1085) );
NAND2_X1 U939 ( .A1(n1272), .A2(n1126), .ZN(n1235) );
XNOR2_X1 U940 ( .A(KEYINPUT55), .B(n1266), .ZN(n1272) );
AND3_X1 U941 ( .A1(n1088), .A2(n1233), .A3(n1079), .ZN(n1230) );
NOR2_X1 U942 ( .A1(n1100), .A2(n1103), .ZN(n1079) );
INV_X1 U943 ( .A(n1106), .ZN(n1103) );
NAND2_X1 U944 ( .A1(n1271), .A2(n1113), .ZN(n1250) );
XNOR2_X1 U945 ( .A(G110), .B(n1225), .ZN(G12) );
NAND3_X1 U946 ( .A1(n1228), .A2(n1084), .A3(n1099), .ZN(n1225) );
INV_X1 U947 ( .A(n1076), .ZN(n1099) );
NAND2_X1 U948 ( .A1(n1270), .A2(n1271), .ZN(n1076) );
XOR2_X1 U949 ( .A(n1273), .B(n1274), .Z(n1271) );
NOR2_X1 U950 ( .A1(G478), .A2(KEYINPUT6), .ZN(n1274) );
XNOR2_X1 U951 ( .A(n1125), .B(KEYINPUT10), .ZN(n1273) );
AND2_X1 U952 ( .A1(n1175), .A2(n1176), .ZN(n1125) );
XOR2_X1 U953 ( .A(n1275), .B(n1276), .Z(n1175) );
XOR2_X1 U954 ( .A(G134), .B(n1277), .Z(n1276) );
XNOR2_X1 U955 ( .A(KEYINPUT43), .B(n1278), .ZN(n1277) );
XOR2_X1 U956 ( .A(n1279), .B(n1280), .Z(n1275) );
XNOR2_X1 U957 ( .A(G128), .B(n1281), .ZN(n1280) );
NAND2_X1 U958 ( .A1(G217), .A2(n1282), .ZN(n1281) );
INV_X1 U959 ( .A(n1283), .ZN(n1282) );
NAND3_X1 U960 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1279) );
NAND2_X1 U961 ( .A1(KEYINPUT1), .A2(G107), .ZN(n1286) );
OR3_X1 U962 ( .A1(G107), .A2(KEYINPUT1), .A3(n1287), .ZN(n1285) );
NAND2_X1 U963 ( .A1(n1287), .A2(n1288), .ZN(n1284) );
NAND2_X1 U964 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
INV_X1 U965 ( .A(KEYINPUT1), .ZN(n1290) );
XNOR2_X1 U966 ( .A(KEYINPUT13), .B(n1063), .ZN(n1289) );
XOR2_X1 U967 ( .A(n1291), .B(n1292), .Z(n1287) );
NOR2_X1 U968 ( .A1(KEYINPUT63), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U969 ( .A(G116), .B(KEYINPUT9), .ZN(n1291) );
INV_X1 U970 ( .A(n1113), .ZN(n1270) );
XNOR2_X1 U971 ( .A(n1294), .B(G475), .ZN(n1113) );
NAND2_X1 U972 ( .A1(n1295), .A2(n1176), .ZN(n1294) );
XNOR2_X1 U973 ( .A(KEYINPUT39), .B(n1296), .ZN(n1295) );
INV_X1 U974 ( .A(n1179), .ZN(n1296) );
XNOR2_X1 U975 ( .A(n1297), .B(n1298), .ZN(n1179) );
XOR2_X1 U976 ( .A(KEYINPUT3), .B(G104), .Z(n1298) );
XOR2_X1 U977 ( .A(n1299), .B(n1300), .Z(n1297) );
NOR2_X1 U978 ( .A1(KEYINPUT56), .A2(n1301), .ZN(n1300) );
XOR2_X1 U979 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U980 ( .A(n1304), .B(n1305), .Z(n1303) );
NOR2_X1 U981 ( .A1(KEYINPUT32), .A2(n1306), .ZN(n1305) );
NOR2_X1 U982 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
XOR2_X1 U983 ( .A(KEYINPUT60), .B(n1309), .Z(n1308) );
NOR2_X1 U984 ( .A1(G125), .A2(n1310), .ZN(n1309) );
NOR2_X1 U985 ( .A1(n1311), .A2(n1261), .ZN(n1307) );
INV_X1 U986 ( .A(G125), .ZN(n1261) );
INV_X1 U987 ( .A(n1310), .ZN(n1311) );
NAND2_X1 U988 ( .A1(n1312), .A2(G214), .ZN(n1304) );
XNOR2_X1 U989 ( .A(G131), .B(n1313), .ZN(n1302) );
XNOR2_X1 U990 ( .A(n1314), .B(G143), .ZN(n1313) );
NAND3_X1 U991 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n1299) );
OR2_X1 U992 ( .A1(G122), .A2(KEYINPUT20), .ZN(n1317) );
NAND3_X1 U993 ( .A1(KEYINPUT20), .A2(G122), .A3(n1318), .ZN(n1316) );
INV_X1 U994 ( .A(G113), .ZN(n1318) );
NAND2_X1 U995 ( .A1(G113), .A2(n1319), .ZN(n1315) );
NAND2_X1 U996 ( .A1(n1320), .A2(KEYINPUT20), .ZN(n1319) );
XNOR2_X1 U997 ( .A(G122), .B(KEYINPUT0), .ZN(n1320) );
INV_X1 U998 ( .A(n1218), .ZN(n1084) );
NAND2_X1 U999 ( .A1(n1321), .A2(n1266), .ZN(n1218) );
NAND3_X1 U1000 ( .A1(n1322), .A2(n1323), .A3(n1324), .ZN(n1266) );
NAND2_X1 U1001 ( .A1(n1115), .A2(n1325), .ZN(n1324) );
OR3_X1 U1002 ( .A1(n1325), .A2(n1115), .A3(n1116), .ZN(n1323) );
INV_X1 U1003 ( .A(KEYINPUT7), .ZN(n1325) );
NAND2_X1 U1004 ( .A1(n1326), .A2(n1116), .ZN(n1322) );
NAND2_X1 U1005 ( .A1(G217), .A2(n1327), .ZN(n1116) );
NAND2_X1 U1006 ( .A1(n1328), .A2(KEYINPUT7), .ZN(n1326) );
XNOR2_X1 U1007 ( .A(n1115), .B(KEYINPUT12), .ZN(n1328) );
NOR2_X1 U1008 ( .A1(n1169), .A2(G902), .ZN(n1115) );
INV_X1 U1009 ( .A(n1165), .ZN(n1169) );
XNOR2_X1 U1010 ( .A(n1329), .B(n1330), .ZN(n1165) );
XNOR2_X1 U1011 ( .A(n1310), .B(n1331), .ZN(n1330) );
XOR2_X1 U1012 ( .A(n1332), .B(n1333), .Z(n1331) );
NOR3_X1 U1013 ( .A1(n1334), .A2(KEYINPUT57), .A3(n1335), .ZN(n1333) );
NOR3_X1 U1014 ( .A1(n1336), .A2(n1337), .A3(n1283), .ZN(n1335) );
XOR2_X1 U1015 ( .A(KEYINPUT24), .B(G137), .Z(n1336) );
NOR2_X1 U1016 ( .A1(n1338), .A2(G137), .ZN(n1334) );
NOR2_X1 U1017 ( .A1(n1337), .A2(n1283), .ZN(n1338) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1131), .ZN(n1283) );
INV_X1 U1019 ( .A(G221), .ZN(n1337) );
NAND3_X1 U1020 ( .A1(n1339), .A2(n1340), .A3(n1341), .ZN(n1332) );
NAND2_X1 U1021 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
INV_X1 U1022 ( .A(KEYINPUT21), .ZN(n1343) );
NAND3_X1 U1023 ( .A1(KEYINPUT21), .A2(n1344), .A3(G110), .ZN(n1340) );
OR2_X1 U1024 ( .A1(n1344), .A2(G110), .ZN(n1339) );
NOR2_X1 U1025 ( .A1(n1345), .A2(n1342), .ZN(n1344) );
XOR2_X1 U1026 ( .A(G119), .B(G128), .Z(n1342) );
INV_X1 U1027 ( .A(KEYINPUT40), .ZN(n1345) );
XOR2_X1 U1028 ( .A(G140), .B(KEYINPUT58), .Z(n1310) );
XOR2_X1 U1029 ( .A(n1346), .B(n1347), .Z(n1329) );
XNOR2_X1 U1030 ( .A(n1314), .B(G125), .ZN(n1347) );
INV_X1 U1031 ( .A(G146), .ZN(n1314) );
XNOR2_X1 U1032 ( .A(KEYINPUT44), .B(KEYINPUT35), .ZN(n1346) );
INV_X1 U1033 ( .A(n1126), .ZN(n1321) );
XOR2_X1 U1034 ( .A(n1348), .B(n1185), .Z(n1126) );
INV_X1 U1035 ( .A(G472), .ZN(n1185) );
NAND2_X1 U1036 ( .A1(n1349), .A2(n1176), .ZN(n1348) );
XNOR2_X1 U1037 ( .A(KEYINPUT33), .B(n1350), .ZN(n1349) );
INV_X1 U1038 ( .A(n1182), .ZN(n1350) );
XNOR2_X1 U1039 ( .A(n1351), .B(n1352), .ZN(n1182) );
XNOR2_X1 U1040 ( .A(n1258), .B(n1353), .ZN(n1352) );
XNOR2_X1 U1041 ( .A(n1278), .B(G113), .ZN(n1353) );
XOR2_X1 U1042 ( .A(n1354), .B(n1355), .Z(n1351) );
XOR2_X1 U1043 ( .A(n1356), .B(n1357), .Z(n1354) );
AND2_X1 U1044 ( .A1(G210), .A2(n1312), .ZN(n1357) );
NOR2_X1 U1045 ( .A1(G953), .A2(G237), .ZN(n1312) );
AND3_X1 U1046 ( .A1(n1098), .A2(n1233), .A3(n1088), .ZN(n1228) );
AND2_X1 U1047 ( .A1(n1092), .A2(n1093), .ZN(n1088) );
NAND2_X1 U1048 ( .A1(G214), .A2(n1358), .ZN(n1093) );
XNOR2_X1 U1049 ( .A(n1359), .B(n1193), .ZN(n1092) );
AND2_X1 U1050 ( .A1(G210), .A2(n1358), .ZN(n1193) );
NAND2_X1 U1051 ( .A1(n1360), .A2(n1361), .ZN(n1358) );
INV_X1 U1052 ( .A(G237), .ZN(n1361) );
NAND2_X1 U1053 ( .A1(n1362), .A2(n1176), .ZN(n1359) );
XNOR2_X1 U1054 ( .A(n1239), .B(n1363), .ZN(n1362) );
XOR2_X1 U1055 ( .A(n1242), .B(KEYINPUT54), .Z(n1363) );
XOR2_X1 U1056 ( .A(n1141), .B(n1364), .Z(n1242) );
XNOR2_X1 U1057 ( .A(n1278), .B(n1365), .ZN(n1364) );
NOR2_X1 U1058 ( .A1(G953), .A2(n1150), .ZN(n1365) );
INV_X1 U1059 ( .A(G224), .ZN(n1150) );
INV_X1 U1060 ( .A(G143), .ZN(n1278) );
XNOR2_X1 U1061 ( .A(G125), .B(n1366), .ZN(n1141) );
XOR2_X1 U1062 ( .A(n1367), .B(n1159), .Z(n1239) );
NAND2_X1 U1063 ( .A1(n1368), .A2(n1369), .ZN(n1159) );
NAND2_X1 U1064 ( .A1(n1370), .A2(G107), .ZN(n1369) );
NAND2_X1 U1065 ( .A1(n1371), .A2(n1063), .ZN(n1368) );
XNOR2_X1 U1066 ( .A(n1370), .B(KEYINPUT59), .ZN(n1371) );
XNOR2_X1 U1067 ( .A(n1157), .B(n1372), .ZN(n1367) );
NOR2_X1 U1068 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
NOR2_X1 U1069 ( .A1(KEYINPUT15), .A2(n1375), .ZN(n1374) );
NOR2_X1 U1070 ( .A1(KEYINPUT36), .A2(n1156), .ZN(n1373) );
INV_X1 U1071 ( .A(n1375), .ZN(n1156) );
XOR2_X1 U1072 ( .A(G110), .B(n1376), .Z(n1375) );
XNOR2_X1 U1073 ( .A(KEYINPUT14), .B(n1293), .ZN(n1376) );
INV_X1 U1074 ( .A(G122), .ZN(n1293) );
XOR2_X1 U1075 ( .A(G113), .B(n1377), .Z(n1157) );
NOR2_X1 U1076 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
AND3_X1 U1077 ( .A1(KEYINPUT11), .A2(n1380), .A3(G116), .ZN(n1379) );
NOR2_X1 U1078 ( .A1(KEYINPUT11), .A2(n1355), .ZN(n1378) );
XNOR2_X1 U1079 ( .A(G116), .B(n1380), .ZN(n1355) );
INV_X1 U1080 ( .A(G119), .ZN(n1380) );
NAND2_X1 U1081 ( .A1(n1078), .A2(n1381), .ZN(n1233) );
NAND4_X1 U1082 ( .A1(G953), .A2(G902), .A3(n1263), .A4(n1151), .ZN(n1381) );
INV_X1 U1083 ( .A(G898), .ZN(n1151) );
NAND3_X1 U1084 ( .A1(n1263), .A2(n1131), .A3(G952), .ZN(n1078) );
INV_X1 U1085 ( .A(G953), .ZN(n1131) );
NAND2_X1 U1086 ( .A1(G237), .A2(G234), .ZN(n1263) );
AND2_X1 U1087 ( .A1(n1100), .A2(n1106), .ZN(n1098) );
NAND2_X1 U1088 ( .A1(n1382), .A2(G221), .ZN(n1106) );
XOR2_X1 U1089 ( .A(n1327), .B(KEYINPUT49), .Z(n1382) );
NAND2_X1 U1090 ( .A1(G234), .A2(n1360), .ZN(n1327) );
XNOR2_X1 U1091 ( .A(n1176), .B(KEYINPUT31), .ZN(n1360) );
XOR2_X1 U1092 ( .A(n1121), .B(G469), .Z(n1100) );
INV_X1 U1093 ( .A(n1120), .ZN(n1121) );
NAND2_X1 U1094 ( .A1(n1383), .A2(n1176), .ZN(n1120) );
INV_X1 U1095 ( .A(G902), .ZN(n1176) );
XNOR2_X1 U1096 ( .A(KEYINPUT62), .B(n1384), .ZN(n1383) );
INV_X1 U1097 ( .A(n1188), .ZN(n1384) );
XNOR2_X1 U1098 ( .A(n1385), .B(n1386), .ZN(n1188) );
XOR2_X1 U1099 ( .A(n1387), .B(n1388), .Z(n1386) );
XNOR2_X1 U1100 ( .A(n1063), .B(n1389), .ZN(n1388) );
NOR2_X1 U1101 ( .A1(G953), .A2(n1132), .ZN(n1389) );
INV_X1 U1102 ( .A(G227), .ZN(n1132) );
INV_X1 U1103 ( .A(G107), .ZN(n1063) );
XNOR2_X1 U1104 ( .A(n1140), .B(G110), .ZN(n1387) );
INV_X1 U1105 ( .A(G140), .ZN(n1140) );
XNOR2_X1 U1106 ( .A(n1390), .B(n1143), .ZN(n1385) );
XNOR2_X1 U1107 ( .A(KEYINPUT38), .B(n1391), .ZN(n1143) );
NOR2_X1 U1108 ( .A1(KEYINPUT2), .A2(n1392), .ZN(n1391) );
XNOR2_X1 U1109 ( .A(G143), .B(KEYINPUT23), .ZN(n1392) );
XOR2_X1 U1110 ( .A(n1356), .B(n1370), .Z(n1390) );
XNOR2_X1 U1111 ( .A(G104), .B(n1258), .ZN(n1370) );
INV_X1 U1112 ( .A(G101), .ZN(n1258) );
XOR2_X1 U1113 ( .A(n1393), .B(n1394), .Z(n1356) );
XOR2_X1 U1114 ( .A(G137), .B(G131), .Z(n1394) );
XOR2_X1 U1115 ( .A(n1395), .B(n1366), .Z(n1393) );
XOR2_X1 U1116 ( .A(G128), .B(G146), .Z(n1366) );
NAND2_X1 U1117 ( .A1(KEYINPUT27), .A2(G134), .ZN(n1395) );
endmodule


