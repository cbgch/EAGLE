//Key = 0111110101010110010110101111100010110000111001010011001000010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361;

XNOR2_X1 U744 ( .A(G107), .B(n1039), .ZN(G9) );
NOR2_X1 U745 ( .A1(n1040), .A2(n1041), .ZN(G75) );
NOR4_X1 U746 ( .A1(n1042), .A2(n1043), .A3(G953), .A4(n1044), .ZN(n1041) );
NOR4_X1 U747 ( .A1(KEYINPUT62), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
NOR3_X1 U748 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1045) );
NAND3_X1 U749 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1042) );
NAND3_X1 U750 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1052) );
NAND2_X1 U751 ( .A1(n1057), .A2(n1058), .ZN(n1054) );
NAND2_X1 U752 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U753 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U754 ( .A1(n1063), .A2(n1064), .ZN(n1057) );
NAND2_X1 U755 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND3_X1 U756 ( .A1(n1067), .A2(n1068), .A3(KEYINPUT62), .ZN(n1066) );
NAND2_X1 U757 ( .A1(KEYINPUT25), .A2(n1069), .ZN(n1065) );
NAND3_X1 U758 ( .A1(n1070), .A2(n1071), .A3(n1063), .ZN(n1051) );
NAND2_X1 U759 ( .A1(n1049), .A2(n1072), .ZN(n1071) );
OR3_X1 U760 ( .A1(n1073), .A2(KEYINPUT25), .A3(n1050), .ZN(n1072) );
NAND2_X1 U761 ( .A1(n1074), .A2(n1055), .ZN(n1070) );
NAND2_X1 U762 ( .A1(n1059), .A2(n1075), .ZN(n1074) );
NAND2_X1 U763 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND3_X1 U764 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
OR2_X1 U765 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NAND3_X1 U766 ( .A1(n1083), .A2(n1084), .A3(n1081), .ZN(n1078) );
OR2_X1 U767 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR3_X1 U768 ( .A1(n1044), .A2(G953), .A3(G952), .ZN(n1040) );
AND4_X1 U769 ( .A1(n1087), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1044) );
NOR4_X1 U770 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1090) );
XOR2_X1 U771 ( .A(n1095), .B(n1096), .Z(n1094) );
XNOR2_X1 U772 ( .A(G469), .B(n1097), .ZN(n1093) );
NAND2_X1 U773 ( .A1(n1098), .A2(KEYINPUT17), .ZN(n1097) );
XOR2_X1 U774 ( .A(n1099), .B(KEYINPUT32), .Z(n1098) );
XOR2_X1 U775 ( .A(n1100), .B(n1101), .Z(n1091) );
NOR2_X1 U776 ( .A1(n1102), .A2(KEYINPUT38), .ZN(n1101) );
AND3_X1 U777 ( .A1(n1103), .A2(n1046), .A3(n1085), .ZN(n1089) );
NAND3_X1 U778 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1087) );
NAND2_X1 U779 ( .A1(KEYINPUT16), .A2(n1107), .ZN(n1106) );
NAND3_X1 U780 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1105) );
INV_X1 U781 ( .A(KEYINPUT16), .ZN(n1109) );
OR2_X1 U782 ( .A1(n1110), .A2(n1108), .ZN(n1104) );
NOR2_X1 U783 ( .A1(n1111), .A2(n1107), .ZN(n1108) );
INV_X1 U784 ( .A(KEYINPUT28), .ZN(n1111) );
XNOR2_X1 U785 ( .A(n1112), .B(KEYINPUT47), .ZN(n1110) );
XOR2_X1 U786 ( .A(n1113), .B(n1114), .Z(G72) );
NAND2_X1 U787 ( .A1(G953), .A2(n1115), .ZN(n1114) );
NAND2_X1 U788 ( .A1(G900), .A2(G227), .ZN(n1115) );
NAND4_X1 U789 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1113) );
NAND3_X1 U790 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
NAND2_X1 U791 ( .A1(G953), .A2(n1123), .ZN(n1118) );
NAND2_X1 U792 ( .A1(G900), .A2(n1120), .ZN(n1123) );
OR2_X1 U793 ( .A1(n1121), .A2(n1120), .ZN(n1117) );
XOR2_X1 U794 ( .A(n1124), .B(n1125), .Z(n1120) );
XOR2_X1 U795 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U796 ( .A1(n1128), .A2(KEYINPUT35), .ZN(n1127) );
XNOR2_X1 U797 ( .A(n1129), .B(KEYINPUT12), .ZN(n1128) );
XOR2_X1 U798 ( .A(n1130), .B(n1131), .Z(n1124) );
NOR3_X1 U799 ( .A1(n1132), .A2(KEYINPUT49), .A3(n1133), .ZN(n1131) );
XOR2_X1 U800 ( .A(KEYINPUT33), .B(n1134), .Z(n1132) );
NOR2_X1 U801 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U802 ( .A(KEYINPUT21), .B(KEYINPUT1), .Z(n1116) );
XOR2_X1 U803 ( .A(n1137), .B(n1138), .Z(G69) );
NOR2_X1 U804 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U805 ( .A(KEYINPUT23), .B(n1141), .Z(n1140) );
NOR2_X1 U806 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
AND2_X1 U807 ( .A1(n1143), .A2(n1142), .ZN(n1139) );
AND2_X1 U808 ( .A1(n1144), .A2(n1145), .ZN(n1142) );
XOR2_X1 U809 ( .A(KEYINPUT2), .B(G953), .Z(n1144) );
NAND2_X1 U810 ( .A1(n1146), .A2(n1147), .ZN(n1143) );
NAND2_X1 U811 ( .A1(G953), .A2(n1148), .ZN(n1147) );
XNOR2_X1 U812 ( .A(n1149), .B(n1150), .ZN(n1146) );
XOR2_X1 U813 ( .A(n1151), .B(KEYINPUT54), .Z(n1150) );
NAND3_X1 U814 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
NAND2_X1 U815 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
OR3_X1 U816 ( .A1(n1156), .A2(n1155), .A3(n1157), .ZN(n1153) );
INV_X1 U817 ( .A(KEYINPUT19), .ZN(n1156) );
NAND2_X1 U818 ( .A1(n1157), .A2(n1158), .ZN(n1152) );
NAND2_X1 U819 ( .A1(n1159), .A2(KEYINPUT19), .ZN(n1158) );
XNOR2_X1 U820 ( .A(n1155), .B(KEYINPUT43), .ZN(n1159) );
NAND2_X1 U821 ( .A1(G953), .A2(n1160), .ZN(n1137) );
NAND2_X1 U822 ( .A1(G898), .A2(G224), .ZN(n1160) );
NOR2_X1 U823 ( .A1(n1161), .A2(n1162), .ZN(G66) );
XOR2_X1 U824 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U825 ( .A1(KEYINPUT57), .A2(n1165), .ZN(n1164) );
AND2_X1 U826 ( .A1(n1102), .A2(n1166), .ZN(n1163) );
NOR2_X1 U827 ( .A1(n1161), .A2(n1167), .ZN(G63) );
NOR3_X1 U828 ( .A1(n1107), .A2(n1168), .A3(n1169), .ZN(n1167) );
AND3_X1 U829 ( .A1(n1170), .A2(G478), .A3(n1166), .ZN(n1169) );
NOR2_X1 U830 ( .A1(n1171), .A2(n1170), .ZN(n1168) );
NOR2_X1 U831 ( .A1(n1053), .A2(n1112), .ZN(n1171) );
INV_X1 U832 ( .A(G478), .ZN(n1112) );
NOR2_X1 U833 ( .A1(n1161), .A2(n1172), .ZN(G60) );
XOR2_X1 U834 ( .A(n1173), .B(n1174), .Z(n1172) );
NAND2_X1 U835 ( .A1(n1166), .A2(G475), .ZN(n1173) );
XOR2_X1 U836 ( .A(G104), .B(n1175), .Z(G6) );
NOR2_X1 U837 ( .A1(n1161), .A2(n1176), .ZN(G57) );
NOR2_X1 U838 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XOR2_X1 U839 ( .A(n1179), .B(KEYINPUT14), .Z(n1178) );
NAND2_X1 U840 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NOR2_X1 U841 ( .A1(n1180), .A2(n1181), .ZN(n1177) );
XNOR2_X1 U842 ( .A(n1182), .B(n1183), .ZN(n1181) );
XOR2_X1 U843 ( .A(n1184), .B(n1185), .Z(n1183) );
XOR2_X1 U844 ( .A(n1186), .B(n1187), .Z(n1182) );
XOR2_X1 U845 ( .A(KEYINPUT30), .B(n1188), .Z(n1187) );
INV_X1 U846 ( .A(n1189), .ZN(n1188) );
NAND2_X1 U847 ( .A1(n1166), .A2(G472), .ZN(n1186) );
NOR2_X1 U848 ( .A1(n1161), .A2(n1190), .ZN(G54) );
XOR2_X1 U849 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U850 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR3_X1 U851 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1194) );
NOR2_X1 U852 ( .A1(n1198), .A2(n1130), .ZN(n1197) );
AND3_X1 U853 ( .A1(n1130), .A2(n1198), .A3(KEYINPUT40), .ZN(n1196) );
NOR2_X1 U854 ( .A1(KEYINPUT46), .A2(n1199), .ZN(n1198) );
NOR2_X1 U855 ( .A1(KEYINPUT40), .A2(n1200), .ZN(n1195) );
NAND3_X1 U856 ( .A1(n1166), .A2(G469), .A3(KEYINPUT41), .ZN(n1193) );
XOR2_X1 U857 ( .A(n1189), .B(n1201), .Z(n1191) );
NOR2_X1 U858 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XOR2_X1 U859 ( .A(KEYINPUT53), .B(n1204), .Z(n1203) );
NOR2_X1 U860 ( .A1(n1161), .A2(n1205), .ZN(G51) );
XOR2_X1 U861 ( .A(n1206), .B(n1207), .Z(n1205) );
XNOR2_X1 U862 ( .A(n1208), .B(KEYINPUT48), .ZN(n1207) );
NAND2_X1 U863 ( .A1(KEYINPUT4), .A2(G125), .ZN(n1208) );
XOR2_X1 U864 ( .A(n1209), .B(n1210), .Z(n1206) );
NAND2_X1 U865 ( .A1(n1166), .A2(n1211), .ZN(n1209) );
NOR2_X1 U866 ( .A1(n1212), .A2(n1053), .ZN(n1166) );
NOR2_X1 U867 ( .A1(n1145), .A2(n1121), .ZN(n1053) );
NAND4_X1 U868 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1121) );
AND4_X1 U869 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1216) );
NAND2_X1 U870 ( .A1(n1059), .A2(n1221), .ZN(n1213) );
NAND2_X1 U871 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
XOR2_X1 U872 ( .A(n1224), .B(KEYINPUT58), .Z(n1222) );
NAND2_X1 U873 ( .A1(n1225), .A2(n1226), .ZN(n1145) );
AND4_X1 U874 ( .A1(n1227), .A2(n1039), .A3(n1228), .A4(n1229), .ZN(n1226) );
NAND3_X1 U875 ( .A1(n1081), .A2(n1230), .A3(n1231), .ZN(n1039) );
NOR4_X1 U876 ( .A1(n1232), .A2(n1233), .A3(n1175), .A4(n1234), .ZN(n1225) );
NOR3_X1 U877 ( .A1(n1076), .A2(n1235), .A3(n1062), .ZN(n1234) );
AND3_X1 U878 ( .A1(n1081), .A2(n1230), .A3(n1236), .ZN(n1175) );
NOR2_X1 U879 ( .A1(n1122), .A2(G952), .ZN(n1161) );
XNOR2_X1 U880 ( .A(G146), .B(n1214), .ZN(G48) );
NAND4_X1 U881 ( .A1(n1237), .A2(n1238), .A3(n1236), .A4(n1069), .ZN(n1214) );
XOR2_X1 U882 ( .A(n1239), .B(n1240), .Z(G45) );
NAND2_X1 U883 ( .A1(KEYINPUT24), .A2(n1241), .ZN(n1240) );
INV_X1 U884 ( .A(n1215), .ZN(n1241) );
NAND4_X1 U885 ( .A1(n1242), .A2(n1069), .A3(n1243), .A4(n1244), .ZN(n1215) );
XOR2_X1 U886 ( .A(n1245), .B(n1246), .Z(G42) );
NAND2_X1 U887 ( .A1(n1247), .A2(n1059), .ZN(n1246) );
XOR2_X1 U888 ( .A(n1223), .B(KEYINPUT7), .Z(n1247) );
NAND2_X1 U889 ( .A1(n1237), .A2(n1248), .ZN(n1223) );
XOR2_X1 U890 ( .A(n1136), .B(n1249), .Z(G39) );
NAND2_X1 U891 ( .A1(n1250), .A2(n1059), .ZN(n1249) );
XOR2_X1 U892 ( .A(n1224), .B(KEYINPUT22), .Z(n1250) );
NAND3_X1 U893 ( .A1(n1238), .A2(n1063), .A3(n1237), .ZN(n1224) );
XOR2_X1 U894 ( .A(G134), .B(n1251), .Z(G36) );
NOR2_X1 U895 ( .A1(KEYINPUT6), .A2(n1220), .ZN(n1251) );
NAND3_X1 U896 ( .A1(n1242), .A2(n1231), .A3(n1059), .ZN(n1220) );
XNOR2_X1 U897 ( .A(n1219), .B(n1252), .ZN(G33) );
NOR2_X1 U898 ( .A1(KEYINPUT52), .A2(n1126), .ZN(n1252) );
NAND3_X1 U899 ( .A1(n1242), .A2(n1236), .A3(n1059), .ZN(n1219) );
NOR2_X1 U900 ( .A1(n1047), .A2(n1068), .ZN(n1059) );
INV_X1 U901 ( .A(n1046), .ZN(n1068) );
AND2_X1 U902 ( .A1(n1237), .A2(n1253), .ZN(n1242) );
NOR2_X1 U903 ( .A1(n1083), .A2(n1254), .ZN(n1237) );
INV_X1 U904 ( .A(n1255), .ZN(n1254) );
XOR2_X1 U905 ( .A(n1256), .B(KEYINPUT39), .Z(n1083) );
XOR2_X1 U906 ( .A(n1257), .B(n1218), .Z(G30) );
NAND4_X1 U907 ( .A1(n1069), .A2(n1255), .A3(n1258), .A4(n1259), .ZN(n1218) );
AND2_X1 U908 ( .A1(n1231), .A2(n1238), .ZN(n1259) );
INV_X1 U909 ( .A(n1256), .ZN(n1258) );
XOR2_X1 U910 ( .A(G101), .B(n1233), .Z(G3) );
AND3_X1 U911 ( .A1(n1063), .A2(n1260), .A3(n1253), .ZN(n1233) );
XOR2_X1 U912 ( .A(n1261), .B(n1217), .Z(G27) );
NAND4_X1 U913 ( .A1(n1248), .A2(n1082), .A3(n1069), .A4(n1255), .ZN(n1217) );
NAND2_X1 U914 ( .A1(n1262), .A2(n1263), .ZN(n1255) );
OR4_X1 U915 ( .A1(n1122), .A2(n1212), .A3(n1049), .A4(G900), .ZN(n1263) );
INV_X1 U916 ( .A(n1055), .ZN(n1049) );
NOR3_X1 U917 ( .A1(n1092), .A2(n1081), .A3(n1061), .ZN(n1248) );
INV_X1 U918 ( .A(n1080), .ZN(n1092) );
XOR2_X1 U919 ( .A(G122), .B(n1264), .Z(G24) );
NOR2_X1 U920 ( .A1(KEYINPUT55), .A2(n1227), .ZN(n1264) );
NAND4_X1 U921 ( .A1(n1056), .A2(n1265), .A3(n1243), .A4(n1244), .ZN(n1227) );
INV_X1 U922 ( .A(n1050), .ZN(n1056) );
NAND3_X1 U923 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1050) );
XOR2_X1 U924 ( .A(G119), .B(n1232), .Z(G21) );
AND4_X1 U925 ( .A1(n1238), .A2(n1063), .A3(n1082), .A4(n1265), .ZN(n1232) );
NOR2_X1 U926 ( .A1(n1080), .A2(n1081), .ZN(n1238) );
XNOR2_X1 U927 ( .A(G116), .B(n1266), .ZN(G18) );
NAND4_X1 U928 ( .A1(n1267), .A2(n1268), .A3(n1231), .A4(n1269), .ZN(n1266) );
INV_X1 U929 ( .A(n1062), .ZN(n1231) );
NAND2_X1 U930 ( .A1(n1270), .A2(n1243), .ZN(n1062) );
XOR2_X1 U931 ( .A(n1073), .B(KEYINPUT13), .Z(n1267) );
NAND2_X1 U932 ( .A1(n1271), .A2(n1272), .ZN(G15) );
NAND2_X1 U933 ( .A1(G113), .A2(n1229), .ZN(n1272) );
XOR2_X1 U934 ( .A(KEYINPUT42), .B(n1273), .Z(n1271) );
NOR2_X1 U935 ( .A1(G113), .A2(n1229), .ZN(n1273) );
NAND3_X1 U936 ( .A1(n1268), .A2(n1265), .A3(n1236), .ZN(n1229) );
INV_X1 U937 ( .A(n1061), .ZN(n1236) );
NAND2_X1 U938 ( .A1(n1274), .A2(n1244), .ZN(n1061) );
INV_X1 U939 ( .A(n1235), .ZN(n1265) );
INV_X1 U940 ( .A(n1076), .ZN(n1268) );
NAND2_X1 U941 ( .A1(n1253), .A2(n1082), .ZN(n1076) );
NOR2_X1 U942 ( .A1(n1086), .A2(n1275), .ZN(n1082) );
INV_X1 U943 ( .A(n1085), .ZN(n1275) );
NOR2_X1 U944 ( .A1(n1276), .A2(n1080), .ZN(n1253) );
XOR2_X1 U945 ( .A(n1277), .B(n1228), .Z(G12) );
NAND3_X1 U946 ( .A1(n1230), .A2(n1276), .A3(n1063), .ZN(n1228) );
INV_X1 U947 ( .A(n1048), .ZN(n1063) );
NAND2_X1 U948 ( .A1(n1274), .A2(n1270), .ZN(n1048) );
XOR2_X1 U949 ( .A(n1244), .B(KEYINPUT59), .Z(n1270) );
NAND3_X1 U950 ( .A1(n1278), .A2(n1279), .A3(n1103), .ZN(n1244) );
NAND3_X1 U951 ( .A1(n1280), .A2(n1212), .A3(n1174), .ZN(n1103) );
NAND2_X1 U952 ( .A1(KEYINPUT37), .A2(n1280), .ZN(n1279) );
INV_X1 U953 ( .A(G475), .ZN(n1280) );
OR2_X1 U954 ( .A1(n1088), .A2(KEYINPUT37), .ZN(n1278) );
NAND2_X1 U955 ( .A1(G475), .A2(n1281), .ZN(n1088) );
NAND2_X1 U956 ( .A1(n1174), .A2(n1212), .ZN(n1281) );
XOR2_X1 U957 ( .A(n1282), .B(n1283), .Z(n1174) );
XOR2_X1 U958 ( .A(n1284), .B(n1285), .Z(n1283) );
XOR2_X1 U959 ( .A(G113), .B(G104), .Z(n1285) );
XOR2_X1 U960 ( .A(KEYINPUT27), .B(G131), .Z(n1284) );
XOR2_X1 U961 ( .A(n1286), .B(n1287), .Z(n1282) );
XOR2_X1 U962 ( .A(n1288), .B(n1289), .Z(n1286) );
NAND3_X1 U963 ( .A1(G214), .A2(n1290), .A3(KEYINPUT61), .ZN(n1288) );
INV_X1 U964 ( .A(n1243), .ZN(n1274) );
XOR2_X1 U965 ( .A(n1107), .B(G478), .Z(n1243) );
NOR2_X1 U966 ( .A1(n1170), .A2(G902), .ZN(n1107) );
XOR2_X1 U967 ( .A(n1291), .B(n1292), .Z(n1170) );
XNOR2_X1 U968 ( .A(n1287), .B(n1293), .ZN(n1292) );
XOR2_X1 U969 ( .A(n1294), .B(n1295), .Z(n1293) );
AND3_X1 U970 ( .A1(G234), .A2(n1122), .A3(G217), .ZN(n1295) );
NAND2_X1 U971 ( .A1(KEYINPUT63), .A2(G107), .ZN(n1294) );
XOR2_X1 U972 ( .A(G122), .B(G143), .Z(n1287) );
XNOR2_X1 U973 ( .A(G116), .B(n1296), .ZN(n1291) );
XOR2_X1 U974 ( .A(G134), .B(G128), .Z(n1296) );
INV_X1 U975 ( .A(n1081), .ZN(n1276) );
XOR2_X1 U976 ( .A(n1100), .B(n1102), .Z(n1081) );
AND2_X1 U977 ( .A1(G217), .A2(n1297), .ZN(n1102) );
NAND2_X1 U978 ( .A1(n1165), .A2(n1212), .ZN(n1100) );
XOR2_X1 U979 ( .A(n1298), .B(n1299), .Z(n1165) );
NOR2_X1 U980 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
XOR2_X1 U981 ( .A(n1302), .B(KEYINPUT51), .Z(n1301) );
NAND2_X1 U982 ( .A1(n1303), .A2(n1289), .ZN(n1302) );
NOR2_X1 U983 ( .A1(n1289), .A2(n1303), .ZN(n1300) );
XOR2_X1 U984 ( .A(n1277), .B(n1304), .Z(n1303) );
NAND3_X1 U985 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1304) );
OR2_X1 U986 ( .A1(n1308), .A2(G119), .ZN(n1307) );
NAND3_X1 U987 ( .A1(G119), .A2(n1308), .A3(n1257), .ZN(n1306) );
NAND2_X1 U988 ( .A1(G128), .A2(n1309), .ZN(n1305) );
NAND2_X1 U989 ( .A1(n1310), .A2(n1308), .ZN(n1309) );
INV_X1 U990 ( .A(KEYINPUT60), .ZN(n1308) );
XOR2_X1 U991 ( .A(KEYINPUT8), .B(G119), .Z(n1310) );
XOR2_X1 U992 ( .A(n1311), .B(n1312), .Z(n1289) );
XOR2_X1 U993 ( .A(KEYINPUT26), .B(n1129), .Z(n1312) );
XNOR2_X1 U994 ( .A(n1261), .B(G140), .ZN(n1129) );
INV_X1 U995 ( .A(G125), .ZN(n1261) );
XOR2_X1 U996 ( .A(n1136), .B(n1313), .Z(n1298) );
AND3_X1 U997 ( .A1(G221), .A2(n1122), .A3(G234), .ZN(n1313) );
AND2_X1 U998 ( .A1(n1260), .A2(n1080), .ZN(n1230) );
XOR2_X1 U999 ( .A(n1314), .B(G472), .Z(n1080) );
NAND2_X1 U1000 ( .A1(n1315), .A2(n1212), .ZN(n1314) );
XOR2_X1 U1001 ( .A(n1316), .B(n1317), .Z(n1315) );
XNOR2_X1 U1002 ( .A(n1185), .B(n1180), .ZN(n1317) );
XOR2_X1 U1003 ( .A(n1318), .B(G101), .Z(n1180) );
NAND2_X1 U1004 ( .A1(G210), .A2(n1290), .ZN(n1318) );
NOR2_X1 U1005 ( .A1(G953), .A2(G237), .ZN(n1290) );
XNOR2_X1 U1006 ( .A(G116), .B(n1319), .ZN(n1185) );
XOR2_X1 U1007 ( .A(n1189), .B(n1320), .Z(n1316) );
NOR2_X1 U1008 ( .A1(KEYINPUT29), .A2(n1184), .ZN(n1320) );
NOR2_X1 U1009 ( .A1(n1235), .A2(n1256), .ZN(n1260) );
NAND2_X1 U1010 ( .A1(n1086), .A2(n1085), .ZN(n1256) );
NAND2_X1 U1011 ( .A1(G221), .A2(n1297), .ZN(n1085) );
NAND2_X1 U1012 ( .A1(G234), .A2(n1212), .ZN(n1297) );
NAND2_X1 U1013 ( .A1(n1321), .A2(n1322), .ZN(n1086) );
NAND2_X1 U1014 ( .A1(G469), .A2(n1099), .ZN(n1322) );
XOR2_X1 U1015 ( .A(n1323), .B(KEYINPUT15), .Z(n1321) );
OR2_X1 U1016 ( .A1(n1099), .A2(G469), .ZN(n1323) );
NAND2_X1 U1017 ( .A1(n1324), .A2(n1212), .ZN(n1099) );
XOR2_X1 U1018 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1019 ( .A(n1130), .B(n1200), .Z(n1326) );
INV_X1 U1020 ( .A(n1199), .ZN(n1200) );
XNOR2_X1 U1021 ( .A(G101), .B(n1327), .ZN(n1199) );
XOR2_X1 U1022 ( .A(n1328), .B(G128), .Z(n1130) );
NAND3_X1 U1023 ( .A1(n1329), .A2(n1330), .A3(KEYINPUT20), .ZN(n1328) );
NAND2_X1 U1024 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
INV_X1 U1025 ( .A(KEYINPUT31), .ZN(n1332) );
XOR2_X1 U1026 ( .A(G143), .B(n1311), .Z(n1331) );
NAND3_X1 U1027 ( .A1(G143), .A2(n1311), .A3(KEYINPUT31), .ZN(n1329) );
XOR2_X1 U1028 ( .A(n1189), .B(n1333), .Z(n1325) );
NOR2_X1 U1029 ( .A1(n1202), .A2(n1204), .ZN(n1333) );
AND2_X1 U1030 ( .A1(n1334), .A2(n1335), .ZN(n1204) );
NAND2_X1 U1031 ( .A1(G227), .A2(n1122), .ZN(n1335) );
XOR2_X1 U1032 ( .A(G140), .B(G110), .Z(n1334) );
AND3_X1 U1033 ( .A1(G227), .A2(n1122), .A3(n1336), .ZN(n1202) );
XOR2_X1 U1034 ( .A(n1245), .B(G110), .Z(n1336) );
INV_X1 U1035 ( .A(G140), .ZN(n1245) );
NAND3_X1 U1036 ( .A1(n1337), .A2(n1338), .A3(n1339), .ZN(n1189) );
NAND2_X1 U1037 ( .A1(n1133), .A2(n1340), .ZN(n1339) );
AND2_X1 U1038 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
INV_X1 U1039 ( .A(G137), .ZN(n1136) );
OR3_X1 U1040 ( .A1(n1340), .A2(n1135), .A3(G137), .ZN(n1338) );
NAND2_X1 U1041 ( .A1(n1341), .A2(G137), .ZN(n1337) );
XOR2_X1 U1042 ( .A(n1340), .B(n1135), .Z(n1341) );
XOR2_X1 U1043 ( .A(G134), .B(KEYINPUT44), .Z(n1135) );
XOR2_X1 U1044 ( .A(n1126), .B(KEYINPUT10), .Z(n1340) );
INV_X1 U1045 ( .A(G131), .ZN(n1126) );
NAND2_X1 U1046 ( .A1(n1069), .A2(n1269), .ZN(n1235) );
NAND2_X1 U1047 ( .A1(n1342), .A2(n1262), .ZN(n1269) );
NAND3_X1 U1048 ( .A1(n1055), .A2(n1122), .A3(n1343), .ZN(n1262) );
XOR2_X1 U1049 ( .A(KEYINPUT36), .B(G952), .Z(n1343) );
INV_X1 U1050 ( .A(G953), .ZN(n1122) );
NAND4_X1 U1051 ( .A1(G953), .A2(G902), .A3(n1055), .A4(n1148), .ZN(n1342) );
INV_X1 U1052 ( .A(G898), .ZN(n1148) );
NAND2_X1 U1053 ( .A1(G237), .A2(G234), .ZN(n1055) );
INV_X1 U1054 ( .A(n1073), .ZN(n1069) );
NAND2_X1 U1055 ( .A1(n1047), .A2(n1046), .ZN(n1073) );
NAND2_X1 U1056 ( .A1(G214), .A2(n1344), .ZN(n1046) );
INV_X1 U1057 ( .A(n1067), .ZN(n1047) );
XOR2_X1 U1058 ( .A(n1345), .B(n1211), .Z(n1067) );
INV_X1 U1059 ( .A(n1095), .ZN(n1211) );
NAND2_X1 U1060 ( .A1(G210), .A2(n1344), .ZN(n1095) );
NAND2_X1 U1061 ( .A1(n1212), .A2(n1346), .ZN(n1344) );
INV_X1 U1062 ( .A(G237), .ZN(n1346) );
NAND2_X1 U1063 ( .A1(KEYINPUT34), .A2(n1347), .ZN(n1345) );
INV_X1 U1064 ( .A(n1096), .ZN(n1347) );
NAND2_X1 U1065 ( .A1(n1348), .A2(n1212), .ZN(n1096) );
INV_X1 U1066 ( .A(G902), .ZN(n1212) );
XOR2_X1 U1067 ( .A(G125), .B(n1210), .Z(n1348) );
XNOR2_X1 U1068 ( .A(n1349), .B(n1350), .ZN(n1210) );
XNOR2_X1 U1069 ( .A(n1184), .B(n1155), .ZN(n1350) );
XOR2_X1 U1070 ( .A(n1327), .B(n1351), .Z(n1155) );
NOR2_X1 U1071 ( .A1(G101), .A2(KEYINPUT56), .ZN(n1351) );
XOR2_X1 U1072 ( .A(G104), .B(G107), .Z(n1327) );
XOR2_X1 U1073 ( .A(n1352), .B(n1311), .Z(n1184) );
XOR2_X1 U1074 ( .A(G146), .B(KEYINPUT45), .Z(n1311) );
XNOR2_X1 U1075 ( .A(n1353), .B(n1354), .ZN(n1352) );
NAND2_X1 U1076 ( .A1(KEYINPUT5), .A2(n1257), .ZN(n1354) );
INV_X1 U1077 ( .A(G128), .ZN(n1257) );
NAND2_X1 U1078 ( .A1(KEYINPUT11), .A2(n1239), .ZN(n1353) );
INV_X1 U1079 ( .A(G143), .ZN(n1239) );
XOR2_X1 U1080 ( .A(n1355), .B(n1356), .Z(n1349) );
NOR2_X1 U1081 ( .A1(KEYINPUT0), .A2(n1149), .ZN(n1356) );
XOR2_X1 U1082 ( .A(G122), .B(G110), .Z(n1149) );
XOR2_X1 U1083 ( .A(n1357), .B(n1358), .Z(n1355) );
NOR2_X1 U1084 ( .A1(G953), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1085 ( .A(KEYINPUT9), .B(G224), .Z(n1359) );
NAND2_X1 U1086 ( .A1(KEYINPUT3), .A2(n1157), .ZN(n1357) );
XOR2_X1 U1087 ( .A(n1360), .B(n1319), .Z(n1157) );
XOR2_X1 U1088 ( .A(G113), .B(G119), .Z(n1319) );
XNOR2_X1 U1089 ( .A(KEYINPUT50), .B(n1361), .ZN(n1360) );
NOR2_X1 U1090 ( .A1(G116), .A2(KEYINPUT18), .ZN(n1361) );
INV_X1 U1091 ( .A(G110), .ZN(n1277) );
endmodule


