//Key = 0101100110011010100110011111011101101010101010001110101101000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417, n1418, n1419, n1420, n1421, n1422;

XOR2_X1 U778 ( .A(G107), .B(n1077), .Z(G9) );
NOR2_X1 U779 ( .A1(n1078), .A2(n1079), .ZN(G75) );
NOR4_X1 U780 ( .A1(n1080), .A2(n1081), .A3(G953), .A4(n1082), .ZN(n1079) );
NOR3_X1 U781 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1081) );
NOR2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
INV_X1 U783 ( .A(n1088), .ZN(n1083) );
NAND3_X1 U784 ( .A1(n1089), .A2(n1090), .A3(KEYINPUT16), .ZN(n1080) );
NAND2_X1 U785 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U786 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U787 ( .A1(n1088), .A2(n1095), .ZN(n1094) );
NAND2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR3_X1 U789 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1088) );
NAND3_X1 U790 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1093) );
NAND2_X1 U791 ( .A1(n1104), .A2(n1100), .ZN(n1102) );
NAND2_X1 U792 ( .A1(KEYINPUT10), .A2(n1105), .ZN(n1104) );
NAND4_X1 U793 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1101) );
INV_X1 U794 ( .A(n1100), .ZN(n1109) );
NAND2_X1 U795 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NAND2_X1 U796 ( .A1(n1112), .A2(n1113), .ZN(n1107) );
NAND2_X1 U797 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XNOR2_X1 U799 ( .A(KEYINPUT35), .B(n1118), .ZN(n1117) );
NAND2_X1 U800 ( .A1(n1105), .A2(n1119), .ZN(n1106) );
INV_X1 U801 ( .A(KEYINPUT10), .ZN(n1119) );
NOR3_X1 U802 ( .A1(n1120), .A2(n1099), .A3(n1121), .ZN(n1105) );
INV_X1 U803 ( .A(n1122), .ZN(n1089) );
NOR3_X1 U804 ( .A1(n1082), .A2(G953), .A3(G952), .ZN(n1078) );
AND4_X1 U805 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n1082) );
NOR4_X1 U806 ( .A1(n1127), .A2(n1116), .A3(n1128), .A4(n1129), .ZN(n1126) );
NOR2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U808 ( .A1(G469), .A2(n1132), .ZN(n1128) );
NOR2_X1 U809 ( .A1(n1133), .A2(n1130), .ZN(n1132) );
INV_X1 U810 ( .A(KEYINPUT23), .ZN(n1130) );
NOR2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(n1125) );
INV_X1 U812 ( .A(n1091), .ZN(n1135) );
XOR2_X1 U813 ( .A(n1136), .B(G475), .Z(n1134) );
NAND2_X1 U814 ( .A1(KEYINPUT50), .A2(n1137), .ZN(n1136) );
XOR2_X1 U815 ( .A(n1138), .B(n1139), .Z(n1124) );
XNOR2_X1 U816 ( .A(KEYINPUT5), .B(n1140), .ZN(n1139) );
NAND2_X1 U817 ( .A1(KEYINPUT61), .A2(n1141), .ZN(n1138) );
XNOR2_X1 U818 ( .A(n1142), .B(n1143), .ZN(n1123) );
NAND2_X1 U819 ( .A1(n1144), .A2(n1145), .ZN(G72) );
NAND2_X1 U820 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND2_X1 U821 ( .A1(G953), .A2(n1148), .ZN(n1147) );
NAND3_X1 U822 ( .A1(G953), .A2(n1149), .A3(n1150), .ZN(n1144) );
INV_X1 U823 ( .A(n1146), .ZN(n1150) );
XNOR2_X1 U824 ( .A(n1151), .B(n1152), .ZN(n1146) );
NOR2_X1 U825 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U826 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U827 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U828 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
OR2_X1 U829 ( .A1(n1161), .A2(KEYINPUT51), .ZN(n1160) );
NAND3_X1 U830 ( .A1(G134), .A2(n1162), .A3(KEYINPUT51), .ZN(n1159) );
XNOR2_X1 U831 ( .A(n1163), .B(n1164), .ZN(n1155) );
XNOR2_X1 U832 ( .A(G131), .B(KEYINPUT54), .ZN(n1163) );
NOR2_X1 U833 ( .A1(G900), .A2(n1165), .ZN(n1153) );
NAND3_X1 U834 ( .A1(n1166), .A2(n1165), .A3(KEYINPUT31), .ZN(n1151) );
NAND2_X1 U835 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND2_X1 U836 ( .A1(G900), .A2(G227), .ZN(n1149) );
NAND3_X1 U837 ( .A1(n1169), .A2(n1170), .A3(n1171), .ZN(G69) );
OR2_X1 U838 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NAND2_X1 U839 ( .A1(n1174), .A2(n1175), .ZN(n1170) );
INV_X1 U840 ( .A(KEYINPUT14), .ZN(n1175) );
NAND2_X1 U841 ( .A1(n1173), .A2(n1176), .ZN(n1174) );
XNOR2_X1 U842 ( .A(KEYINPUT44), .B(n1172), .ZN(n1176) );
NAND2_X1 U843 ( .A1(KEYINPUT14), .A2(n1177), .ZN(n1169) );
NAND2_X1 U844 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND3_X1 U845 ( .A1(KEYINPUT44), .A2(n1173), .A3(n1172), .ZN(n1179) );
XOR2_X1 U846 ( .A(n1180), .B(n1181), .Z(n1173) );
NOR2_X1 U847 ( .A1(G953), .A2(n1182), .ZN(n1181) );
NOR2_X1 U848 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XNOR2_X1 U849 ( .A(KEYINPUT59), .B(n1185), .ZN(n1184) );
NAND2_X1 U850 ( .A1(KEYINPUT8), .A2(n1186), .ZN(n1180) );
NAND2_X1 U851 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND2_X1 U852 ( .A1(G953), .A2(n1189), .ZN(n1188) );
XOR2_X1 U853 ( .A(n1190), .B(n1191), .Z(n1187) );
XOR2_X1 U854 ( .A(KEYINPUT17), .B(KEYINPUT13), .Z(n1191) );
XOR2_X1 U855 ( .A(n1192), .B(n1193), .Z(n1190) );
OR2_X1 U856 ( .A1(n1172), .A2(KEYINPUT44), .ZN(n1178) );
NAND2_X1 U857 ( .A1(G953), .A2(n1194), .ZN(n1172) );
NAND2_X1 U858 ( .A1(G898), .A2(G224), .ZN(n1194) );
NOR2_X1 U859 ( .A1(n1195), .A2(n1196), .ZN(G66) );
XOR2_X1 U860 ( .A(n1197), .B(n1198), .Z(n1196) );
NOR2_X1 U861 ( .A1(n1199), .A2(n1200), .ZN(n1197) );
NOR2_X1 U862 ( .A1(n1201), .A2(n1202), .ZN(G63) );
XOR2_X1 U863 ( .A(KEYINPUT22), .B(n1195), .Z(n1202) );
XOR2_X1 U864 ( .A(n1203), .B(n1204), .Z(n1201) );
NOR2_X1 U865 ( .A1(n1140), .A2(n1200), .ZN(n1203) );
NOR2_X1 U866 ( .A1(n1195), .A2(n1205), .ZN(G60) );
XNOR2_X1 U867 ( .A(n1206), .B(n1207), .ZN(n1205) );
NOR2_X1 U868 ( .A1(n1208), .A2(n1200), .ZN(n1207) );
XNOR2_X1 U869 ( .A(G475), .B(KEYINPUT18), .ZN(n1208) );
XNOR2_X1 U870 ( .A(n1209), .B(n1210), .ZN(G6) );
NOR2_X1 U871 ( .A1(n1195), .A2(n1211), .ZN(G57) );
XNOR2_X1 U872 ( .A(n1212), .B(n1213), .ZN(n1211) );
NOR2_X1 U873 ( .A1(n1214), .A2(n1200), .ZN(n1213) );
NOR3_X1 U874 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(G54) );
AND2_X1 U875 ( .A1(KEYINPUT19), .A2(n1195), .ZN(n1217) );
NOR3_X1 U876 ( .A1(KEYINPUT19), .A2(G953), .A3(G952), .ZN(n1216) );
XOR2_X1 U877 ( .A(n1218), .B(n1219), .Z(n1215) );
XOR2_X1 U878 ( .A(n1220), .B(n1221), .Z(n1219) );
NAND2_X1 U879 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
NAND2_X1 U880 ( .A1(G140), .A2(n1224), .ZN(n1223) );
XOR2_X1 U881 ( .A(KEYINPUT49), .B(n1225), .Z(n1222) );
NOR2_X1 U882 ( .A1(G140), .A2(n1224), .ZN(n1225) );
XOR2_X1 U883 ( .A(KEYINPUT45), .B(n1226), .Z(n1218) );
NOR2_X1 U884 ( .A1(n1227), .A2(n1200), .ZN(n1226) );
NOR2_X1 U885 ( .A1(n1195), .A2(n1228), .ZN(G51) );
XOR2_X1 U886 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U887 ( .A(n1231), .B(n1232), .Z(n1230) );
NOR2_X1 U888 ( .A1(n1143), .A2(n1200), .ZN(n1231) );
NAND2_X1 U889 ( .A1(G902), .A2(n1122), .ZN(n1200) );
NAND4_X1 U890 ( .A1(n1233), .A2(n1167), .A3(n1234), .A4(n1185), .ZN(n1122) );
NAND2_X1 U891 ( .A1(n1235), .A2(n1110), .ZN(n1185) );
INV_X1 U892 ( .A(n1183), .ZN(n1234) );
NAND4_X1 U893 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1183) );
NOR4_X1 U894 ( .A1(n1240), .A2(n1241), .A3(n1077), .A4(n1210), .ZN(n1239) );
NOR3_X1 U895 ( .A1(n1242), .A2(n1243), .A3(n1096), .ZN(n1210) );
NOR3_X1 U896 ( .A1(n1243), .A2(n1097), .A3(n1242), .ZN(n1077) );
INV_X1 U897 ( .A(n1244), .ZN(n1241) );
OR2_X1 U898 ( .A1(n1245), .A2(n1096), .ZN(n1238) );
NAND4_X1 U899 ( .A1(n1112), .A2(n1091), .A3(n1246), .A4(n1247), .ZN(n1237) );
NOR3_X1 U900 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1247) );
XNOR2_X1 U901 ( .A(n1251), .B(KEYINPUT34), .ZN(n1246) );
NAND2_X1 U902 ( .A1(n1251), .A2(n1252), .ZN(n1236) );
XNOR2_X1 U903 ( .A(KEYINPUT0), .B(n1253), .ZN(n1252) );
AND4_X1 U904 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1167) );
AND4_X1 U905 ( .A1(n1258), .A2(n1259), .A3(n1260), .A4(n1261), .ZN(n1257) );
NAND4_X1 U906 ( .A1(n1262), .A2(n1110), .A3(n1263), .A4(n1264), .ZN(n1256) );
NOR2_X1 U907 ( .A1(n1265), .A2(n1114), .ZN(n1263) );
XOR2_X1 U908 ( .A(n1266), .B(KEYINPUT7), .Z(n1265) );
NAND3_X1 U909 ( .A1(n1267), .A2(n1266), .A3(n1268), .ZN(n1254) );
XNOR2_X1 U910 ( .A(n1110), .B(KEYINPUT11), .ZN(n1268) );
XOR2_X1 U911 ( .A(n1168), .B(KEYINPUT28), .Z(n1233) );
NOR2_X1 U912 ( .A1(n1165), .A2(G952), .ZN(n1195) );
XNOR2_X1 U913 ( .A(G146), .B(n1255), .ZN(G48) );
NAND4_X1 U914 ( .A1(n1262), .A2(n1269), .A3(n1270), .A4(n1251), .ZN(n1255) );
XNOR2_X1 U915 ( .A(G143), .B(n1261), .ZN(G45) );
NAND3_X1 U916 ( .A1(n1086), .A2(n1269), .A3(n1271), .ZN(n1261) );
NOR3_X1 U917 ( .A1(n1114), .A2(n1250), .A3(n1248), .ZN(n1271) );
XOR2_X1 U918 ( .A(n1272), .B(G140), .Z(G42) );
NAND2_X1 U919 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND3_X1 U920 ( .A1(n1275), .A2(n1099), .A3(n1276), .ZN(n1274) );
OR2_X1 U921 ( .A1(n1168), .A2(n1276), .ZN(n1273) );
INV_X1 U922 ( .A(KEYINPUT12), .ZN(n1276) );
NAND2_X1 U923 ( .A1(n1275), .A2(n1111), .ZN(n1168) );
AND3_X1 U924 ( .A1(n1087), .A2(n1270), .A3(n1269), .ZN(n1275) );
XNOR2_X1 U925 ( .A(n1162), .B(n1277), .ZN(G39) );
AND2_X1 U926 ( .A1(n1269), .A2(n1267), .ZN(n1277) );
NOR3_X1 U927 ( .A1(n1085), .A2(n1099), .A3(n1278), .ZN(n1267) );
INV_X1 U928 ( .A(n1111), .ZN(n1099) );
XOR2_X1 U929 ( .A(n1260), .B(n1279), .Z(G36) );
NAND2_X1 U930 ( .A1(KEYINPUT24), .A2(G134), .ZN(n1279) );
NAND2_X1 U931 ( .A1(n1280), .A2(n1264), .ZN(n1260) );
XNOR2_X1 U932 ( .A(n1281), .B(n1282), .ZN(G33) );
NAND2_X1 U933 ( .A1(KEYINPUT29), .A2(n1259), .ZN(n1281) );
NAND2_X1 U934 ( .A1(n1280), .A2(n1270), .ZN(n1259) );
AND3_X1 U935 ( .A1(n1269), .A2(n1111), .A3(n1086), .ZN(n1280) );
NAND2_X1 U936 ( .A1(n1283), .A2(n1284), .ZN(n1111) );
OR3_X1 U937 ( .A1(n1118), .A2(n1116), .A3(KEYINPUT35), .ZN(n1284) );
INV_X1 U938 ( .A(n1285), .ZN(n1116) );
NAND2_X1 U939 ( .A1(KEYINPUT35), .A2(n1251), .ZN(n1283) );
INV_X1 U940 ( .A(n1286), .ZN(n1269) );
XOR2_X1 U941 ( .A(n1287), .B(n1288), .Z(G30) );
NOR4_X1 U942 ( .A1(n1114), .A2(n1097), .A3(n1286), .A4(n1278), .ZN(n1288) );
NAND2_X1 U943 ( .A1(n1110), .A2(n1266), .ZN(n1286) );
XNOR2_X1 U944 ( .A(G128), .B(KEYINPUT3), .ZN(n1287) );
XOR2_X1 U945 ( .A(n1289), .B(n1290), .Z(G3) );
NOR2_X1 U946 ( .A1(n1114), .A2(n1253), .ZN(n1290) );
NAND4_X1 U947 ( .A1(n1086), .A2(n1103), .A3(n1110), .A4(n1291), .ZN(n1253) );
NAND2_X1 U948 ( .A1(n1292), .A2(KEYINPUT36), .ZN(n1289) );
XNOR2_X1 U949 ( .A(G101), .B(KEYINPUT2), .ZN(n1292) );
XNOR2_X1 U950 ( .A(G125), .B(n1258), .ZN(G27) );
NAND4_X1 U951 ( .A1(n1087), .A2(n1270), .A3(n1293), .A4(n1112), .ZN(n1258) );
AND2_X1 U952 ( .A1(n1266), .A2(n1251), .ZN(n1293) );
INV_X1 U953 ( .A(n1114), .ZN(n1251) );
NAND2_X1 U954 ( .A1(n1100), .A2(n1294), .ZN(n1266) );
NAND2_X1 U955 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
INV_X1 U956 ( .A(G900), .ZN(n1296) );
INV_X1 U957 ( .A(n1096), .ZN(n1270) );
XOR2_X1 U958 ( .A(n1297), .B(n1298), .Z(G24) );
NOR2_X1 U959 ( .A1(KEYINPUT46), .A2(n1299), .ZN(n1298) );
NOR4_X1 U960 ( .A1(n1250), .A2(n1248), .A3(n1242), .A4(n1098), .ZN(n1297) );
INV_X1 U961 ( .A(n1112), .ZN(n1098) );
NAND2_X1 U962 ( .A1(n1300), .A2(n1091), .ZN(n1242) );
NOR2_X1 U963 ( .A1(n1301), .A2(n1302), .ZN(n1091) );
XNOR2_X1 U964 ( .A(G119), .B(n1244), .ZN(G21) );
NAND4_X1 U965 ( .A1(n1262), .A2(n1103), .A3(n1112), .A4(n1300), .ZN(n1244) );
INV_X1 U966 ( .A(n1278), .ZN(n1262) );
NAND2_X1 U967 ( .A1(n1302), .A2(n1301), .ZN(n1278) );
XNOR2_X1 U968 ( .A(n1303), .B(n1240), .ZN(G18) );
NOR2_X1 U969 ( .A1(n1245), .A2(n1097), .ZN(n1240) );
INV_X1 U970 ( .A(n1264), .ZN(n1097) );
NOR2_X1 U971 ( .A1(n1304), .A2(n1248), .ZN(n1264) );
XNOR2_X1 U972 ( .A(n1305), .B(n1306), .ZN(G15) );
NOR3_X1 U973 ( .A1(n1245), .A2(KEYINPUT6), .A3(n1096), .ZN(n1306) );
NAND2_X1 U974 ( .A1(n1248), .A2(n1304), .ZN(n1096) );
NAND3_X1 U975 ( .A1(n1112), .A2(n1300), .A3(n1086), .ZN(n1245) );
AND2_X1 U976 ( .A1(n1307), .A2(n1302), .ZN(n1086) );
NOR2_X1 U977 ( .A1(n1121), .A2(n1308), .ZN(n1112) );
NAND2_X1 U978 ( .A1(n1309), .A2(n1310), .ZN(G12) );
NAND2_X1 U979 ( .A1(G110), .A2(n1311), .ZN(n1310) );
XOR2_X1 U980 ( .A(KEYINPUT4), .B(n1312), .Z(n1309) );
NOR2_X1 U981 ( .A1(G110), .A2(n1311), .ZN(n1312) );
NAND2_X1 U982 ( .A1(n1235), .A2(n1313), .ZN(n1311) );
XNOR2_X1 U983 ( .A(KEYINPUT41), .B(n1243), .ZN(n1313) );
INV_X1 U984 ( .A(n1110), .ZN(n1243) );
NOR2_X1 U985 ( .A1(n1308), .A2(n1314), .ZN(n1110) );
INV_X1 U986 ( .A(n1121), .ZN(n1314) );
NAND2_X1 U987 ( .A1(n1131), .A2(n1315), .ZN(n1121) );
NAND2_X1 U988 ( .A1(n1133), .A2(n1227), .ZN(n1315) );
INV_X1 U989 ( .A(G469), .ZN(n1227) );
INV_X1 U990 ( .A(n1316), .ZN(n1133) );
NAND2_X1 U991 ( .A1(G469), .A2(n1316), .ZN(n1131) );
NAND2_X1 U992 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
XOR2_X1 U993 ( .A(n1319), .B(n1221), .Z(n1317) );
XOR2_X1 U994 ( .A(n1320), .B(n1321), .Z(n1221) );
XOR2_X1 U995 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U996 ( .A(KEYINPUT1), .B(n1209), .ZN(n1323) );
INV_X1 U997 ( .A(G104), .ZN(n1209) );
NOR2_X1 U998 ( .A1(G953), .A2(n1148), .ZN(n1322) );
INV_X1 U999 ( .A(G227), .ZN(n1148) );
XNOR2_X1 U1000 ( .A(n1324), .B(n1157), .ZN(n1320) );
NAND2_X1 U1001 ( .A1(n1325), .A2(n1326), .ZN(n1157) );
NAND2_X1 U1002 ( .A1(n1327), .A2(G146), .ZN(n1326) );
NAND2_X1 U1003 ( .A1(n1328), .A2(n1329), .ZN(n1325) );
XNOR2_X1 U1004 ( .A(n1327), .B(KEYINPUT21), .ZN(n1328) );
XNOR2_X1 U1005 ( .A(n1330), .B(n1331), .ZN(n1324) );
NAND2_X1 U1006 ( .A1(KEYINPUT26), .A2(n1332), .ZN(n1319) );
XNOR2_X1 U1007 ( .A(G140), .B(n1224), .ZN(n1332) );
XOR2_X1 U1008 ( .A(n1127), .B(KEYINPUT58), .Z(n1308) );
INV_X1 U1009 ( .A(n1120), .ZN(n1127) );
NAND2_X1 U1010 ( .A1(G221), .A2(n1333), .ZN(n1120) );
NAND2_X1 U1011 ( .A1(G234), .A2(n1318), .ZN(n1333) );
AND3_X1 U1012 ( .A1(n1103), .A2(n1300), .A3(n1087), .ZN(n1235) );
NOR2_X1 U1013 ( .A1(n1302), .A2(n1307), .ZN(n1087) );
INV_X1 U1014 ( .A(n1301), .ZN(n1307) );
NAND3_X1 U1015 ( .A1(n1334), .A2(n1335), .A3(n1336), .ZN(n1301) );
NAND2_X1 U1016 ( .A1(n1337), .A2(n1198), .ZN(n1336) );
OR3_X1 U1017 ( .A1(n1198), .A2(n1337), .A3(G902), .ZN(n1335) );
NOR2_X1 U1018 ( .A1(n1199), .A2(G234), .ZN(n1337) );
INV_X1 U1019 ( .A(G217), .ZN(n1199) );
XNOR2_X1 U1020 ( .A(n1338), .B(n1339), .ZN(n1198) );
XNOR2_X1 U1021 ( .A(n1224), .B(n1340), .ZN(n1339) );
XNOR2_X1 U1022 ( .A(n1341), .B(n1342), .ZN(n1340) );
NOR4_X1 U1023 ( .A1(n1343), .A2(n1344), .A3(KEYINPUT62), .A4(n1345), .ZN(n1342) );
NOR2_X1 U1024 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
AND2_X1 U1025 ( .A1(n1348), .A2(KEYINPUT30), .ZN(n1346) );
NOR2_X1 U1026 ( .A1(KEYINPUT57), .A2(n1348), .ZN(n1344) );
AND4_X1 U1027 ( .A1(n1348), .A2(KEYINPUT57), .A3(n1347), .A4(KEYINPUT30), .ZN(n1343) );
NAND2_X1 U1028 ( .A1(KEYINPUT48), .A2(n1164), .ZN(n1341) );
XNOR2_X1 U1029 ( .A(G125), .B(G140), .ZN(n1164) );
XOR2_X1 U1030 ( .A(n1349), .B(n1350), .Z(n1338) );
XNOR2_X1 U1031 ( .A(n1329), .B(G137), .ZN(n1350) );
NAND3_X1 U1032 ( .A1(n1351), .A2(n1165), .A3(G234), .ZN(n1349) );
XOR2_X1 U1033 ( .A(KEYINPUT56), .B(G221), .Z(n1351) );
NAND2_X1 U1034 ( .A1(G217), .A2(G902), .ZN(n1334) );
XOR2_X1 U1035 ( .A(n1352), .B(n1214), .Z(n1302) );
INV_X1 U1036 ( .A(G472), .ZN(n1214) );
NAND2_X1 U1037 ( .A1(n1212), .A2(n1318), .ZN(n1352) );
XNOR2_X1 U1038 ( .A(n1353), .B(n1354), .ZN(n1212) );
XNOR2_X1 U1039 ( .A(n1355), .B(n1356), .ZN(n1354) );
XNOR2_X1 U1040 ( .A(n1331), .B(n1357), .ZN(n1353) );
XOR2_X1 U1041 ( .A(n1358), .B(n1359), .Z(n1357) );
NAND2_X1 U1042 ( .A1(n1360), .A2(G210), .ZN(n1359) );
NAND2_X1 U1043 ( .A1(n1361), .A2(n1362), .ZN(n1358) );
XOR2_X1 U1044 ( .A(n1363), .B(KEYINPUT60), .Z(n1361) );
XNOR2_X1 U1045 ( .A(n1282), .B(n1161), .ZN(n1331) );
XNOR2_X1 U1046 ( .A(G134), .B(n1162), .ZN(n1161) );
INV_X1 U1047 ( .A(G137), .ZN(n1162) );
NOR2_X1 U1048 ( .A1(n1114), .A2(n1249), .ZN(n1300) );
INV_X1 U1049 ( .A(n1291), .ZN(n1249) );
NAND2_X1 U1050 ( .A1(n1364), .A2(n1100), .ZN(n1291) );
NAND3_X1 U1051 ( .A1(n1365), .A2(n1165), .A3(G952), .ZN(n1100) );
NAND2_X1 U1052 ( .A1(n1295), .A2(n1189), .ZN(n1364) );
INV_X1 U1053 ( .A(G898), .ZN(n1189) );
AND3_X1 U1054 ( .A1(n1366), .A2(n1365), .A3(G953), .ZN(n1295) );
NAND2_X1 U1055 ( .A1(G237), .A2(G234), .ZN(n1365) );
XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n1318), .ZN(n1366) );
NAND2_X1 U1057 ( .A1(n1118), .A2(n1285), .ZN(n1114) );
NAND2_X1 U1058 ( .A1(G214), .A2(n1367), .ZN(n1285) );
NAND2_X1 U1059 ( .A1(n1368), .A2(n1369), .ZN(n1118) );
NAND2_X1 U1060 ( .A1(n1370), .A2(n1142), .ZN(n1369) );
XOR2_X1 U1061 ( .A(KEYINPUT63), .B(n1371), .Z(n1368) );
NOR2_X1 U1062 ( .A1(n1370), .A2(n1142), .ZN(n1371) );
NAND2_X1 U1063 ( .A1(n1372), .A2(n1318), .ZN(n1142) );
XOR2_X1 U1064 ( .A(n1373), .B(n1232), .Z(n1372) );
XOR2_X1 U1065 ( .A(n1193), .B(n1374), .Z(n1232) );
XNOR2_X1 U1066 ( .A(n1375), .B(KEYINPUT33), .ZN(n1374) );
NAND2_X1 U1067 ( .A1(KEYINPUT52), .A2(n1192), .ZN(n1375) );
XOR2_X1 U1068 ( .A(n1376), .B(n1330), .Z(n1192) );
XNOR2_X1 U1069 ( .A(G107), .B(n1377), .ZN(n1330) );
INV_X1 U1070 ( .A(n1355), .ZN(n1377) );
XOR2_X1 U1071 ( .A(G101), .B(KEYINPUT25), .Z(n1355) );
XOR2_X1 U1072 ( .A(n1378), .B(n1379), .Z(n1376) );
NOR2_X1 U1073 ( .A1(G104), .A2(KEYINPUT32), .ZN(n1379) );
NAND2_X1 U1074 ( .A1(n1380), .A2(n1363), .ZN(n1378) );
NAND2_X1 U1075 ( .A1(n1381), .A2(n1305), .ZN(n1363) );
INV_X1 U1076 ( .A(G113), .ZN(n1305) );
XNOR2_X1 U1077 ( .A(G116), .B(G119), .ZN(n1381) );
XOR2_X1 U1078 ( .A(n1362), .B(KEYINPUT15), .Z(n1380) );
NAND2_X1 U1079 ( .A1(G113), .A2(n1382), .ZN(n1362) );
XNOR2_X1 U1080 ( .A(n1348), .B(G116), .ZN(n1382) );
INV_X1 U1081 ( .A(G119), .ZN(n1348) );
XNOR2_X1 U1082 ( .A(G122), .B(n1224), .ZN(n1193) );
XNOR2_X1 U1083 ( .A(G110), .B(KEYINPUT39), .ZN(n1224) );
NOR2_X1 U1084 ( .A1(KEYINPUT43), .A2(n1229), .ZN(n1373) );
XNOR2_X1 U1085 ( .A(n1356), .B(n1383), .ZN(n1229) );
XOR2_X1 U1086 ( .A(G125), .B(n1384), .Z(n1383) );
AND2_X1 U1087 ( .A1(n1165), .A2(G224), .ZN(n1384) );
XOR2_X1 U1088 ( .A(n1385), .B(n1386), .Z(n1356) );
XNOR2_X1 U1089 ( .A(n1329), .B(G143), .ZN(n1386) );
NAND2_X1 U1090 ( .A1(KEYINPUT27), .A2(n1347), .ZN(n1385) );
INV_X1 U1091 ( .A(G128), .ZN(n1347) );
INV_X1 U1092 ( .A(n1143), .ZN(n1370) );
NAND2_X1 U1093 ( .A1(G210), .A2(n1367), .ZN(n1143) );
NAND2_X1 U1094 ( .A1(n1387), .A2(n1318), .ZN(n1367) );
INV_X1 U1095 ( .A(G237), .ZN(n1387) );
INV_X1 U1096 ( .A(n1085), .ZN(n1103) );
NAND2_X1 U1097 ( .A1(n1248), .A2(n1250), .ZN(n1085) );
INV_X1 U1098 ( .A(n1304), .ZN(n1250) );
XNOR2_X1 U1099 ( .A(n1137), .B(G475), .ZN(n1304) );
NAND2_X1 U1100 ( .A1(n1388), .A2(n1206), .ZN(n1137) );
XNOR2_X1 U1101 ( .A(n1389), .B(n1390), .ZN(n1206) );
XOR2_X1 U1102 ( .A(n1391), .B(n1392), .Z(n1390) );
XOR2_X1 U1103 ( .A(n1393), .B(n1394), .Z(n1392) );
NOR2_X1 U1104 ( .A1(KEYINPUT37), .A2(n1282), .ZN(n1394) );
INV_X1 U1105 ( .A(G131), .ZN(n1282) );
NAND2_X1 U1106 ( .A1(n1395), .A2(n1396), .ZN(n1393) );
NAND3_X1 U1107 ( .A1(G125), .A2(n1397), .A3(n1398), .ZN(n1396) );
XNOR2_X1 U1108 ( .A(G146), .B(n1399), .ZN(n1398) );
NOR2_X1 U1109 ( .A1(G140), .A2(n1400), .ZN(n1399) );
INV_X1 U1110 ( .A(KEYINPUT38), .ZN(n1400) );
NAND2_X1 U1111 ( .A1(n1401), .A2(n1402), .ZN(n1395) );
NAND2_X1 U1112 ( .A1(G125), .A2(n1397), .ZN(n1402) );
INV_X1 U1113 ( .A(KEYINPUT9), .ZN(n1397) );
XNOR2_X1 U1114 ( .A(n1403), .B(n1329), .ZN(n1401) );
INV_X1 U1115 ( .A(G146), .ZN(n1329) );
NAND2_X1 U1116 ( .A1(KEYINPUT38), .A2(G140), .ZN(n1403) );
NAND2_X1 U1117 ( .A1(n1360), .A2(G214), .ZN(n1391) );
NOR2_X1 U1118 ( .A1(G953), .A2(G237), .ZN(n1360) );
XOR2_X1 U1119 ( .A(n1404), .B(n1405), .Z(n1389) );
XNOR2_X1 U1120 ( .A(n1406), .B(G122), .ZN(n1405) );
XNOR2_X1 U1121 ( .A(G104), .B(G113), .ZN(n1404) );
XNOR2_X1 U1122 ( .A(KEYINPUT42), .B(n1318), .ZN(n1388) );
INV_X1 U1123 ( .A(G902), .ZN(n1318) );
XOR2_X1 U1124 ( .A(n1141), .B(n1140), .Z(n1248) );
INV_X1 U1125 ( .A(G478), .ZN(n1140) );
NOR2_X1 U1126 ( .A1(n1204), .A2(G902), .ZN(n1141) );
XNOR2_X1 U1127 ( .A(n1407), .B(n1408), .ZN(n1204) );
XOR2_X1 U1128 ( .A(n1409), .B(n1327), .Z(n1408) );
XNOR2_X1 U1129 ( .A(G128), .B(n1406), .ZN(n1327) );
INV_X1 U1130 ( .A(G143), .ZN(n1406) );
AND3_X1 U1131 ( .A1(G217), .A2(n1165), .A3(G234), .ZN(n1409) );
INV_X1 U1132 ( .A(G953), .ZN(n1165) );
XOR2_X1 U1133 ( .A(n1410), .B(G134), .Z(n1407) );
NAND3_X1 U1134 ( .A1(n1411), .A2(n1412), .A3(KEYINPUT55), .ZN(n1410) );
NAND2_X1 U1135 ( .A1(n1413), .A2(n1414), .ZN(n1412) );
NAND2_X1 U1136 ( .A1(n1415), .A2(n1416), .ZN(n1413) );
NAND2_X1 U1137 ( .A1(n1417), .A2(n1299), .ZN(n1416) );
NAND2_X1 U1138 ( .A1(G107), .A2(G122), .ZN(n1415) );
NAND2_X1 U1139 ( .A1(n1418), .A2(n1419), .ZN(n1411) );
NAND2_X1 U1140 ( .A1(n1420), .A2(n1421), .ZN(n1419) );
NAND2_X1 U1141 ( .A1(G107), .A2(n1299), .ZN(n1421) );
INV_X1 U1142 ( .A(G122), .ZN(n1299) );
NAND2_X1 U1143 ( .A1(n1417), .A2(G122), .ZN(n1420) );
XNOR2_X1 U1144 ( .A(n1422), .B(G107), .ZN(n1417) );
XNOR2_X1 U1145 ( .A(KEYINPUT47), .B(KEYINPUT20), .ZN(n1422) );
INV_X1 U1146 ( .A(n1414), .ZN(n1418) );
NAND2_X1 U1147 ( .A1(KEYINPUT40), .A2(n1303), .ZN(n1414) );
INV_X1 U1148 ( .A(G116), .ZN(n1303) );
endmodule


