//Key = 1101001011101001110101101100100010011000011110000010001101100101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
n1480, n1481;

XOR2_X1 U805 ( .A(n1120), .B(n1121), .Z(G9) );
NOR2_X1 U806 ( .A1(n1122), .A2(n1123), .ZN(G75) );
NOR3_X1 U807 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
XOR2_X1 U808 ( .A(n1127), .B(KEYINPUT7), .Z(n1125) );
NAND3_X1 U809 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1124) );
NAND3_X1 U810 ( .A1(n1131), .A2(n1132), .A3(KEYINPUT6), .ZN(n1128) );
NAND2_X1 U811 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
NAND3_X1 U812 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1134) );
NAND2_X1 U813 ( .A1(n1138), .A2(n1139), .ZN(n1135) );
NAND4_X1 U814 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1139) );
INV_X1 U815 ( .A(KEYINPUT0), .ZN(n1143) );
NAND2_X1 U816 ( .A1(n1144), .A2(n1145), .ZN(n1138) );
NAND2_X1 U817 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND2_X1 U818 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND2_X1 U819 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND2_X1 U820 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U821 ( .A1(n1140), .A2(n1154), .ZN(n1146) );
NAND2_X1 U822 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND2_X1 U823 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND3_X1 U824 ( .A1(n1140), .A2(n1142), .A3(n1148), .ZN(n1133) );
NAND3_X1 U825 ( .A1(n1159), .A2(n1160), .A3(n1148), .ZN(n1142) );
NAND2_X1 U826 ( .A1(n1161), .A2(n1136), .ZN(n1160) );
NAND2_X1 U827 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND3_X1 U828 ( .A1(n1137), .A2(n1141), .A3(KEYINPUT0), .ZN(n1163) );
NAND2_X1 U829 ( .A1(n1144), .A2(n1164), .ZN(n1162) );
OR2_X1 U830 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NAND3_X1 U831 ( .A1(n1137), .A2(n1167), .A3(n1168), .ZN(n1159) );
AND3_X1 U832 ( .A1(n1130), .A2(n1169), .A3(n1129), .ZN(n1122) );
NAND4_X1 U833 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1129) );
NOR4_X1 U834 ( .A1(n1174), .A2(n1141), .A3(n1175), .A4(n1176), .ZN(n1173) );
XOR2_X1 U835 ( .A(n1177), .B(G478), .Z(n1175) );
NAND2_X1 U836 ( .A1(KEYINPUT21), .A2(n1178), .ZN(n1177) );
NAND3_X1 U837 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1174) );
XOR2_X1 U838 ( .A(n1182), .B(n1183), .Z(n1181) );
OR3_X1 U839 ( .A1(n1184), .A2(n1185), .A3(KEYINPUT39), .ZN(n1180) );
NAND2_X1 U840 ( .A1(KEYINPUT39), .A2(n1185), .ZN(n1179) );
NOR3_X1 U841 ( .A1(n1157), .A2(n1186), .A3(n1168), .ZN(n1172) );
NAND2_X1 U842 ( .A1(G475), .A2(n1187), .ZN(n1171) );
XOR2_X1 U843 ( .A(KEYINPUT55), .B(n1188), .Z(n1170) );
INV_X1 U844 ( .A(G952), .ZN(n1169) );
XOR2_X1 U845 ( .A(n1189), .B(n1190), .Z(G72) );
NOR2_X1 U846 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U847 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U848 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U849 ( .A(G131), .B(n1197), .Z(n1196) );
XOR2_X1 U850 ( .A(n1198), .B(n1199), .Z(n1193) );
NAND2_X1 U851 ( .A1(KEYINPUT41), .A2(n1200), .ZN(n1198) );
NAND2_X1 U852 ( .A1(n1201), .A2(n1202), .ZN(n1189) );
NAND2_X1 U853 ( .A1(KEYINPUT15), .A2(n1203), .ZN(n1202) );
NAND2_X1 U854 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NAND2_X1 U855 ( .A1(n1206), .A2(G953), .ZN(n1205) );
XNOR2_X1 U856 ( .A(G227), .B(KEYINPUT30), .ZN(n1206) );
INV_X1 U857 ( .A(n1191), .ZN(n1204) );
NAND2_X1 U858 ( .A1(n1126), .A2(n1207), .ZN(n1201) );
XOR2_X1 U859 ( .A(n1208), .B(n1209), .Z(G69) );
NOR2_X1 U860 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NOR3_X1 U861 ( .A1(n1212), .A2(n1213), .A3(n1207), .ZN(n1211) );
NOR2_X1 U862 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
INV_X1 U863 ( .A(n1216), .ZN(n1212) );
NOR2_X1 U864 ( .A1(n1217), .A2(n1216), .ZN(n1210) );
NAND3_X1 U865 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1216) );
XOR2_X1 U866 ( .A(n1221), .B(KEYINPUT29), .Z(n1220) );
OR2_X1 U867 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NAND2_X1 U868 ( .A1(n1222), .A2(n1223), .ZN(n1219) );
XNOR2_X1 U869 ( .A(n1224), .B(n1225), .ZN(n1222) );
XNOR2_X1 U870 ( .A(KEYINPUT26), .B(n1226), .ZN(n1224) );
NOR2_X1 U871 ( .A1(KEYINPUT40), .A2(n1227), .ZN(n1226) );
NAND2_X1 U872 ( .A1(G953), .A2(n1215), .ZN(n1218) );
NOR2_X1 U873 ( .A1(G224), .A2(n1207), .ZN(n1217) );
NAND2_X1 U874 ( .A1(n1207), .A2(n1127), .ZN(n1208) );
NOR3_X1 U875 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(G66) );
NOR2_X1 U876 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XOR2_X1 U877 ( .A(n1233), .B(KEYINPUT56), .Z(n1232) );
NOR2_X1 U878 ( .A1(n1234), .A2(n1235), .ZN(n1229) );
XNOR2_X1 U879 ( .A(KEYINPUT4), .B(n1233), .ZN(n1235) );
NAND2_X1 U880 ( .A1(n1236), .A2(n1237), .ZN(n1233) );
INV_X1 U881 ( .A(n1184), .ZN(n1237) );
INV_X1 U882 ( .A(n1231), .ZN(n1234) );
NOR2_X1 U883 ( .A1(n1228), .A2(n1238), .ZN(G63) );
XOR2_X1 U884 ( .A(n1239), .B(n1240), .Z(n1238) );
NAND2_X1 U885 ( .A1(n1236), .A2(G478), .ZN(n1240) );
NAND2_X1 U886 ( .A1(KEYINPUT1), .A2(n1241), .ZN(n1239) );
NOR2_X1 U887 ( .A1(n1228), .A2(n1242), .ZN(G60) );
XOR2_X1 U888 ( .A(n1243), .B(n1244), .Z(n1242) );
NAND2_X1 U889 ( .A1(n1236), .A2(G475), .ZN(n1243) );
XOR2_X1 U890 ( .A(n1245), .B(n1246), .Z(G6) );
NAND2_X1 U891 ( .A1(n1165), .A2(n1247), .ZN(n1246) );
NOR2_X1 U892 ( .A1(n1228), .A2(n1248), .ZN(G57) );
XOR2_X1 U893 ( .A(n1249), .B(n1250), .Z(n1248) );
XOR2_X1 U894 ( .A(n1251), .B(n1252), .Z(n1250) );
NAND2_X1 U895 ( .A1(KEYINPUT12), .A2(n1253), .ZN(n1251) );
XOR2_X1 U896 ( .A(n1254), .B(n1255), .Z(n1249) );
NOR3_X1 U897 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1255) );
AND2_X1 U898 ( .A1(n1259), .A2(KEYINPUT2), .ZN(n1258) );
AND3_X1 U899 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1257) );
INV_X1 U900 ( .A(KEYINPUT2), .ZN(n1260) );
NOR2_X1 U901 ( .A1(n1262), .A2(n1261), .ZN(n1256) );
NOR2_X1 U902 ( .A1(KEYINPUT62), .A2(n1259), .ZN(n1262) );
NAND2_X1 U903 ( .A1(n1236), .A2(G472), .ZN(n1254) );
NOR2_X1 U904 ( .A1(n1228), .A2(n1263), .ZN(G54) );
XOR2_X1 U905 ( .A(n1264), .B(n1265), .Z(n1263) );
NAND2_X1 U906 ( .A1(n1236), .A2(G469), .ZN(n1265) );
NAND2_X1 U907 ( .A1(n1266), .A2(n1267), .ZN(n1264) );
NAND2_X1 U908 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XOR2_X1 U909 ( .A(n1195), .B(n1270), .Z(n1269) );
XOR2_X1 U910 ( .A(n1271), .B(n1272), .Z(n1268) );
XOR2_X1 U911 ( .A(n1273), .B(KEYINPUT47), .Z(n1266) );
NAND2_X1 U912 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XNOR2_X1 U913 ( .A(n1271), .B(n1272), .ZN(n1275) );
XOR2_X1 U914 ( .A(G110), .B(n1276), .Z(n1272) );
NAND2_X1 U915 ( .A1(KEYINPUT36), .A2(n1277), .ZN(n1271) );
XOR2_X1 U916 ( .A(n1270), .B(n1278), .Z(n1274) );
INV_X1 U917 ( .A(n1195), .ZN(n1278) );
NOR2_X1 U918 ( .A1(n1228), .A2(n1279), .ZN(G51) );
XOR2_X1 U919 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U920 ( .A(n1282), .B(n1283), .Z(n1281) );
XOR2_X1 U921 ( .A(n1284), .B(n1285), .Z(n1280) );
XOR2_X1 U922 ( .A(KEYINPUT3), .B(n1286), .Z(n1285) );
NAND2_X1 U923 ( .A1(n1236), .A2(n1183), .ZN(n1284) );
AND2_X1 U924 ( .A1(G902), .A2(n1287), .ZN(n1236) );
OR2_X1 U925 ( .A1(n1126), .A2(n1127), .ZN(n1287) );
NAND4_X1 U926 ( .A1(n1288), .A2(n1289), .A3(n1290), .A4(n1291), .ZN(n1127) );
NOR4_X1 U927 ( .A1(n1292), .A2(n1293), .A3(n1294), .A4(n1295), .ZN(n1291) );
INV_X1 U928 ( .A(n1296), .ZN(n1295) );
INV_X1 U929 ( .A(n1121), .ZN(n1294) );
NAND2_X1 U930 ( .A1(n1166), .A2(n1247), .ZN(n1121) );
AND2_X1 U931 ( .A1(n1140), .A2(n1297), .ZN(n1247) );
NOR2_X1 U932 ( .A1(n1298), .A2(n1299), .ZN(n1290) );
AND4_X1 U933 ( .A1(n1300), .A2(n1140), .A3(n1165), .A4(n1301), .ZN(n1299) );
XOR2_X1 U934 ( .A(KEYINPUT52), .B(n1302), .Z(n1301) );
NAND4_X1 U935 ( .A1(n1303), .A2(n1304), .A3(n1305), .A4(n1306), .ZN(n1126) );
NOR4_X1 U936 ( .A1(n1307), .A2(n1308), .A3(n1309), .A4(n1310), .ZN(n1306) );
INV_X1 U937 ( .A(n1311), .ZN(n1310) );
INV_X1 U938 ( .A(n1312), .ZN(n1308) );
NAND2_X1 U939 ( .A1(n1313), .A2(n1314), .ZN(n1305) );
NAND2_X1 U940 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XNOR2_X1 U941 ( .A(n1317), .B(KEYINPUT53), .ZN(n1315) );
NAND2_X1 U942 ( .A1(n1148), .A2(n1318), .ZN(n1304) );
XOR2_X1 U943 ( .A(KEYINPUT46), .B(n1319), .Z(n1318) );
NAND2_X1 U944 ( .A1(n1320), .A2(n1321), .ZN(n1303) );
NOR2_X1 U945 ( .A1(n1207), .A2(G952), .ZN(n1228) );
XOR2_X1 U946 ( .A(n1322), .B(n1311), .Z(G48) );
NAND3_X1 U947 ( .A1(n1300), .A2(n1176), .A3(n1323), .ZN(n1311) );
XOR2_X1 U948 ( .A(n1324), .B(n1325), .Z(G45) );
NAND2_X1 U949 ( .A1(n1317), .A2(n1313), .ZN(n1325) );
AND3_X1 U950 ( .A1(n1326), .A2(n1327), .A3(n1328), .ZN(n1317) );
XOR2_X1 U951 ( .A(G140), .B(n1309), .Z(G42) );
AND3_X1 U952 ( .A1(n1148), .A2(n1141), .A3(n1329), .ZN(n1309) );
XOR2_X1 U953 ( .A(n1330), .B(n1312), .Z(G39) );
NAND4_X1 U954 ( .A1(n1148), .A2(n1141), .A3(n1331), .A4(n1332), .ZN(n1312) );
NOR3_X1 U955 ( .A1(n1152), .A2(n1168), .A3(n1333), .ZN(n1332) );
XOR2_X1 U956 ( .A(n1307), .B(n1334), .Z(G36) );
NOR2_X1 U957 ( .A1(KEYINPUT37), .A2(n1335), .ZN(n1334) );
AND3_X1 U958 ( .A1(n1148), .A2(n1166), .A3(n1328), .ZN(n1307) );
XNOR2_X1 U959 ( .A(G131), .B(n1336), .ZN(G33) );
NAND2_X1 U960 ( .A1(n1319), .A2(n1148), .ZN(n1336) );
AND2_X1 U961 ( .A1(n1158), .A2(n1337), .ZN(n1148) );
AND2_X1 U962 ( .A1(n1165), .A2(n1328), .ZN(n1319) );
NOR4_X1 U963 ( .A1(n1150), .A2(n1167), .A3(n1333), .A4(n1168), .ZN(n1328) );
XOR2_X1 U964 ( .A(n1338), .B(G128), .Z(G30) );
NAND2_X1 U965 ( .A1(KEYINPUT50), .A2(n1339), .ZN(n1338) );
NAND2_X1 U966 ( .A1(n1340), .A2(n1320), .ZN(n1339) );
AND4_X1 U967 ( .A1(n1166), .A2(n1300), .A3(n1176), .A4(n1153), .ZN(n1320) );
XOR2_X1 U968 ( .A(n1321), .B(KEYINPUT5), .Z(n1340) );
NAND3_X1 U969 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(G3) );
NAND2_X1 U970 ( .A1(G101), .A2(n1344), .ZN(n1343) );
NAND2_X1 U971 ( .A1(KEYINPUT20), .A2(n1345), .ZN(n1342) );
NAND2_X1 U972 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
XOR2_X1 U973 ( .A(KEYINPUT18), .B(n1298), .Z(n1346) );
INV_X1 U974 ( .A(n1344), .ZN(n1298) );
NAND2_X1 U975 ( .A1(n1348), .A2(n1349), .ZN(n1341) );
INV_X1 U976 ( .A(KEYINPUT20), .ZN(n1349) );
NAND2_X1 U977 ( .A1(n1350), .A2(n1351), .ZN(n1348) );
OR3_X1 U978 ( .A1(n1344), .A2(G101), .A3(KEYINPUT18), .ZN(n1351) );
NAND2_X1 U979 ( .A1(KEYINPUT18), .A2(n1344), .ZN(n1350) );
NAND3_X1 U980 ( .A1(n1352), .A2(n1297), .A3(n1137), .ZN(n1344) );
XOR2_X1 U981 ( .A(n1200), .B(n1353), .Z(G27) );
NAND2_X1 U982 ( .A1(n1354), .A2(n1313), .ZN(n1353) );
XOR2_X1 U983 ( .A(n1316), .B(KEYINPUT9), .Z(n1354) );
NAND2_X1 U984 ( .A1(n1329), .A2(n1144), .ZN(n1316) );
AND3_X1 U985 ( .A1(n1152), .A2(n1136), .A3(n1323), .ZN(n1329) );
NOR3_X1 U986 ( .A1(n1333), .A2(n1355), .A3(n1356), .ZN(n1323) );
INV_X1 U987 ( .A(n1321), .ZN(n1333) );
NAND2_X1 U988 ( .A1(n1357), .A2(n1358), .ZN(n1321) );
NAND3_X1 U989 ( .A1(G902), .A2(n1132), .A3(n1191), .ZN(n1358) );
NOR2_X1 U990 ( .A1(G900), .A2(n1207), .ZN(n1191) );
XNOR2_X1 U991 ( .A(G122), .B(n1288), .ZN(G24) );
NAND4_X1 U992 ( .A1(n1359), .A2(n1140), .A3(n1326), .A4(n1327), .ZN(n1288) );
NOR2_X1 U993 ( .A1(n1153), .A2(n1176), .ZN(n1140) );
XNOR2_X1 U994 ( .A(n1360), .B(n1289), .ZN(G21) );
NAND3_X1 U995 ( .A1(n1331), .A2(n1176), .A3(n1359), .ZN(n1289) );
XOR2_X1 U996 ( .A(n1361), .B(KEYINPUT58), .Z(n1360) );
XOR2_X1 U997 ( .A(G116), .B(n1293), .Z(G18) );
AND3_X1 U998 ( .A1(n1352), .A2(n1166), .A3(n1359), .ZN(n1293) );
NOR2_X1 U999 ( .A1(n1327), .A2(n1362), .ZN(n1166) );
XOR2_X1 U1000 ( .A(G113), .B(n1292), .Z(G15) );
AND3_X1 U1001 ( .A1(n1165), .A2(n1352), .A3(n1359), .ZN(n1292) );
AND4_X1 U1002 ( .A1(n1313), .A2(n1144), .A3(n1302), .A4(n1136), .ZN(n1359) );
XOR2_X1 U1003 ( .A(n1141), .B(KEYINPUT22), .Z(n1144) );
INV_X1 U1004 ( .A(n1167), .ZN(n1141) );
INV_X1 U1005 ( .A(n1150), .ZN(n1352) );
NAND2_X1 U1006 ( .A1(n1355), .A2(n1176), .ZN(n1150) );
INV_X1 U1007 ( .A(n1152), .ZN(n1176) );
INV_X1 U1008 ( .A(n1356), .ZN(n1165) );
NAND2_X1 U1009 ( .A1(n1362), .A2(n1327), .ZN(n1356) );
XOR2_X1 U1010 ( .A(G110), .B(n1363), .Z(G12) );
NOR2_X1 U1011 ( .A1(KEYINPUT11), .A2(n1296), .ZN(n1363) );
NAND3_X1 U1012 ( .A1(n1152), .A2(n1297), .A3(n1331), .ZN(n1296) );
AND2_X1 U1013 ( .A1(n1137), .A2(n1153), .ZN(n1331) );
INV_X1 U1014 ( .A(n1355), .ZN(n1153) );
NOR2_X1 U1015 ( .A1(n1186), .A2(n1364), .ZN(n1355) );
NOR2_X1 U1016 ( .A1(n1184), .A2(n1185), .ZN(n1364) );
AND2_X1 U1017 ( .A1(n1185), .A2(n1184), .ZN(n1186) );
NAND2_X1 U1018 ( .A1(G217), .A2(n1365), .ZN(n1184) );
NOR2_X1 U1019 ( .A1(n1231), .A2(G902), .ZN(n1185) );
XOR2_X1 U1020 ( .A(n1366), .B(n1367), .Z(n1231) );
XOR2_X1 U1021 ( .A(n1368), .B(n1369), .Z(n1367) );
NOR2_X1 U1022 ( .A1(KEYINPUT51), .A2(n1370), .ZN(n1369) );
XOR2_X1 U1023 ( .A(n1200), .B(n1371), .Z(n1370) );
XOR2_X1 U1024 ( .A(G146), .B(G140), .Z(n1371) );
NOR2_X1 U1025 ( .A1(n1372), .A2(n1373), .ZN(n1368) );
NOR2_X1 U1026 ( .A1(n1374), .A2(G137), .ZN(n1373) );
NOR2_X1 U1027 ( .A1(n1375), .A2(n1376), .ZN(n1374) );
NOR3_X1 U1028 ( .A1(n1376), .A2(n1377), .A3(n1375), .ZN(n1372) );
XOR2_X1 U1029 ( .A(n1330), .B(KEYINPUT45), .Z(n1377) );
INV_X1 U1030 ( .A(G221), .ZN(n1376) );
XNOR2_X1 U1031 ( .A(G110), .B(n1378), .ZN(n1366) );
XOR2_X1 U1032 ( .A(G128), .B(G119), .Z(n1378) );
NOR2_X1 U1033 ( .A1(n1326), .A2(n1327), .ZN(n1137) );
NAND2_X1 U1034 ( .A1(n1379), .A2(n1380), .ZN(n1327) );
NAND2_X1 U1035 ( .A1(G475), .A2(n1381), .ZN(n1380) );
NAND2_X1 U1036 ( .A1(KEYINPUT19), .A2(n1382), .ZN(n1381) );
INV_X1 U1037 ( .A(n1187), .ZN(n1382) );
NAND2_X1 U1038 ( .A1(n1188), .A2(KEYINPUT19), .ZN(n1379) );
NOR2_X1 U1039 ( .A1(n1187), .A2(G475), .ZN(n1188) );
NAND2_X1 U1040 ( .A1(n1244), .A2(n1383), .ZN(n1187) );
XNOR2_X1 U1041 ( .A(n1384), .B(n1385), .ZN(n1244) );
XOR2_X1 U1042 ( .A(n1386), .B(n1387), .Z(n1385) );
XNOR2_X1 U1043 ( .A(n1388), .B(n1389), .ZN(n1387) );
NOR4_X1 U1044 ( .A1(KEYINPUT27), .A2(G953), .A3(G237), .A4(n1390), .ZN(n1389) );
INV_X1 U1045 ( .A(G214), .ZN(n1390) );
NAND2_X1 U1046 ( .A1(n1391), .A2(KEYINPUT43), .ZN(n1388) );
XOR2_X1 U1047 ( .A(n1245), .B(n1392), .Z(n1391) );
XOR2_X1 U1048 ( .A(G122), .B(G113), .Z(n1392) );
NOR3_X1 U1049 ( .A1(n1393), .A2(n1394), .A3(n1395), .ZN(n1386) );
NOR2_X1 U1050 ( .A1(KEYINPUT8), .A2(n1197), .ZN(n1395) );
NOR3_X1 U1051 ( .A1(G140), .A2(n1200), .A3(n1396), .ZN(n1394) );
INV_X1 U1052 ( .A(G125), .ZN(n1200) );
NOR2_X1 U1053 ( .A1(G125), .A2(n1397), .ZN(n1393) );
NOR2_X1 U1054 ( .A1(n1396), .A2(n1398), .ZN(n1397) );
XOR2_X1 U1055 ( .A(KEYINPUT48), .B(G140), .Z(n1398) );
INV_X1 U1056 ( .A(KEYINPUT8), .ZN(n1396) );
XNOR2_X1 U1057 ( .A(G131), .B(n1399), .ZN(n1384) );
XOR2_X1 U1058 ( .A(G146), .B(G143), .Z(n1399) );
INV_X1 U1059 ( .A(n1362), .ZN(n1326) );
XOR2_X1 U1060 ( .A(n1178), .B(G478), .Z(n1362) );
OR2_X1 U1061 ( .A1(n1241), .A2(G902), .ZN(n1178) );
XOR2_X1 U1062 ( .A(n1400), .B(n1401), .Z(n1241) );
XOR2_X1 U1063 ( .A(n1402), .B(n1403), .Z(n1401) );
XOR2_X1 U1064 ( .A(n1404), .B(G107), .Z(n1403) );
NAND2_X1 U1065 ( .A1(G217), .A2(n1405), .ZN(n1404) );
INV_X1 U1066 ( .A(n1375), .ZN(n1405) );
NAND2_X1 U1067 ( .A1(G234), .A2(n1207), .ZN(n1375) );
NAND2_X1 U1068 ( .A1(n1406), .A2(KEYINPUT35), .ZN(n1402) );
XOR2_X1 U1069 ( .A(n1324), .B(n1407), .Z(n1406) );
NOR2_X1 U1070 ( .A1(G128), .A2(KEYINPUT33), .ZN(n1407) );
XOR2_X1 U1071 ( .A(n1408), .B(n1409), .Z(n1400) );
XOR2_X1 U1072 ( .A(G134), .B(G122), .Z(n1409) );
AND2_X1 U1073 ( .A1(n1300), .A2(n1302), .ZN(n1297) );
NAND2_X1 U1074 ( .A1(n1357), .A2(n1410), .ZN(n1302) );
NAND4_X1 U1075 ( .A1(G953), .A2(G902), .A3(n1132), .A4(n1215), .ZN(n1410) );
INV_X1 U1076 ( .A(G898), .ZN(n1215) );
NAND3_X1 U1077 ( .A1(n1130), .A2(n1132), .A3(G952), .ZN(n1357) );
NAND2_X1 U1078 ( .A1(G237), .A2(G234), .ZN(n1132) );
XNOR2_X1 U1079 ( .A(n1207), .B(KEYINPUT32), .ZN(n1130) );
NOR3_X1 U1080 ( .A1(n1167), .A2(n1168), .A3(n1155), .ZN(n1300) );
INV_X1 U1081 ( .A(n1313), .ZN(n1155) );
NOR2_X1 U1082 ( .A1(n1158), .A2(n1157), .ZN(n1313) );
INV_X1 U1083 ( .A(n1337), .ZN(n1157) );
NAND2_X1 U1084 ( .A1(G214), .A2(n1411), .ZN(n1337) );
XNOR2_X1 U1085 ( .A(n1412), .B(n1183), .ZN(n1158) );
AND2_X1 U1086 ( .A1(G210), .A2(n1411), .ZN(n1183) );
NAND2_X1 U1087 ( .A1(n1413), .A2(n1383), .ZN(n1411) );
NAND2_X1 U1088 ( .A1(KEYINPUT42), .A2(n1182), .ZN(n1412) );
NAND2_X1 U1089 ( .A1(n1414), .A2(n1383), .ZN(n1182) );
XOR2_X1 U1090 ( .A(n1415), .B(n1416), .Z(n1414) );
NOR2_X1 U1091 ( .A1(KEYINPUT14), .A2(n1283), .ZN(n1416) );
XNOR2_X1 U1092 ( .A(n1417), .B(n1223), .ZN(n1283) );
XNOR2_X1 U1093 ( .A(G110), .B(n1418), .ZN(n1223) );
XOR2_X1 U1094 ( .A(KEYINPUT54), .B(G122), .Z(n1418) );
XOR2_X1 U1095 ( .A(n1419), .B(n1227), .Z(n1417) );
AND2_X1 U1096 ( .A1(n1420), .A2(n1421), .ZN(n1227) );
NAND2_X1 U1097 ( .A1(n1422), .A2(n1423), .ZN(n1421) );
XOR2_X1 U1098 ( .A(KEYINPUT25), .B(n1424), .Z(n1420) );
NOR2_X1 U1099 ( .A1(n1422), .A2(n1423), .ZN(n1424) );
INV_X1 U1100 ( .A(n1425), .ZN(n1423) );
AND2_X1 U1101 ( .A1(n1426), .A2(n1427), .ZN(n1422) );
NAND2_X1 U1102 ( .A1(n1428), .A2(n1245), .ZN(n1427) );
NAND2_X1 U1103 ( .A1(KEYINPUT24), .A2(n1429), .ZN(n1428) );
NAND2_X1 U1104 ( .A1(KEYINPUT28), .A2(n1120), .ZN(n1429) );
INV_X1 U1105 ( .A(G107), .ZN(n1120) );
NAND2_X1 U1106 ( .A1(G107), .A2(n1430), .ZN(n1426) );
NAND2_X1 U1107 ( .A1(KEYINPUT28), .A2(n1431), .ZN(n1430) );
NAND2_X1 U1108 ( .A1(KEYINPUT24), .A2(G104), .ZN(n1431) );
NAND2_X1 U1109 ( .A1(KEYINPUT16), .A2(n1225), .ZN(n1419) );
AND2_X1 U1110 ( .A1(n1432), .A2(n1433), .ZN(n1225) );
NAND2_X1 U1111 ( .A1(n1434), .A2(n1435), .ZN(n1433) );
INV_X1 U1112 ( .A(G113), .ZN(n1435) );
XOR2_X1 U1113 ( .A(G116), .B(n1436), .Z(n1434) );
NAND2_X1 U1114 ( .A1(G113), .A2(n1437), .ZN(n1432) );
XOR2_X1 U1115 ( .A(n1408), .B(n1436), .Z(n1437) );
NOR2_X1 U1116 ( .A1(G119), .A2(KEYINPUT38), .ZN(n1436) );
INV_X1 U1117 ( .A(G116), .ZN(n1408) );
XNOR2_X1 U1118 ( .A(n1286), .B(n1438), .ZN(n1415) );
NOR2_X1 U1119 ( .A1(KEYINPUT23), .A2(n1282), .ZN(n1438) );
XOR2_X1 U1120 ( .A(n1261), .B(G125), .Z(n1282) );
NOR2_X1 U1121 ( .A1(n1214), .A2(G953), .ZN(n1286) );
INV_X1 U1122 ( .A(G224), .ZN(n1214) );
INV_X1 U1123 ( .A(n1136), .ZN(n1168) );
NAND2_X1 U1124 ( .A1(G221), .A2(n1365), .ZN(n1136) );
NAND2_X1 U1125 ( .A1(G234), .A2(n1383), .ZN(n1365) );
XOR2_X1 U1126 ( .A(n1439), .B(G469), .Z(n1167) );
NAND2_X1 U1127 ( .A1(n1440), .A2(n1383), .ZN(n1439) );
XOR2_X1 U1128 ( .A(n1441), .B(n1442), .Z(n1440) );
XNOR2_X1 U1129 ( .A(n1270), .B(n1277), .ZN(n1442) );
XNOR2_X1 U1130 ( .A(n1197), .B(KEYINPUT63), .ZN(n1277) );
INV_X1 U1131 ( .A(G140), .ZN(n1197) );
XOR2_X1 U1132 ( .A(n1443), .B(n1444), .Z(n1270) );
XOR2_X1 U1133 ( .A(n1259), .B(n1445), .Z(n1444) );
NAND2_X1 U1134 ( .A1(KEYINPUT44), .A2(n1425), .ZN(n1445) );
XOR2_X1 U1135 ( .A(n1347), .B(KEYINPUT13), .Z(n1425) );
INV_X1 U1136 ( .A(G101), .ZN(n1347) );
XOR2_X1 U1137 ( .A(n1245), .B(G107), .Z(n1443) );
INV_X1 U1138 ( .A(G104), .ZN(n1245) );
XOR2_X1 U1139 ( .A(n1446), .B(n1447), .Z(n1441) );
XNOR2_X1 U1140 ( .A(G110), .B(n1448), .ZN(n1447) );
NOR2_X1 U1141 ( .A1(KEYINPUT49), .A2(n1195), .ZN(n1448) );
NAND3_X1 U1142 ( .A1(n1449), .A2(n1450), .A3(n1451), .ZN(n1195) );
NAND2_X1 U1143 ( .A1(G143), .A2(n1452), .ZN(n1450) );
XOR2_X1 U1144 ( .A(n1453), .B(n1454), .Z(n1452) );
NAND2_X1 U1145 ( .A1(n1455), .A2(n1324), .ZN(n1449) );
NAND2_X1 U1146 ( .A1(n1456), .A2(n1457), .ZN(n1455) );
NAND2_X1 U1147 ( .A1(n1454), .A2(n1453), .ZN(n1457) );
NOR2_X1 U1148 ( .A1(KEYINPUT59), .A2(G146), .ZN(n1454) );
NAND2_X1 U1149 ( .A1(KEYINPUT59), .A2(G128), .ZN(n1456) );
NAND2_X1 U1150 ( .A1(KEYINPUT57), .A2(n1276), .ZN(n1446) );
AND2_X1 U1151 ( .A1(G227), .A2(n1207), .ZN(n1276) );
XOR2_X1 U1152 ( .A(n1458), .B(G472), .Z(n1152) );
NAND2_X1 U1153 ( .A1(n1459), .A2(n1383), .ZN(n1458) );
INV_X1 U1154 ( .A(G902), .ZN(n1383) );
XNOR2_X1 U1155 ( .A(n1460), .B(n1253), .ZN(n1459) );
XNOR2_X1 U1156 ( .A(n1461), .B(G101), .ZN(n1253) );
NAND3_X1 U1157 ( .A1(n1413), .A2(n1207), .A3(G210), .ZN(n1461) );
INV_X1 U1158 ( .A(G953), .ZN(n1207) );
INV_X1 U1159 ( .A(G237), .ZN(n1413) );
NAND2_X1 U1160 ( .A1(n1462), .A2(n1463), .ZN(n1460) );
XOR2_X1 U1161 ( .A(KEYINPUT31), .B(KEYINPUT10), .Z(n1463) );
XOR2_X1 U1162 ( .A(n1464), .B(n1465), .Z(n1462) );
INV_X1 U1163 ( .A(n1252), .ZN(n1465) );
XOR2_X1 U1164 ( .A(n1466), .B(n1467), .Z(n1252) );
XOR2_X1 U1165 ( .A(G116), .B(G113), .Z(n1467) );
NAND2_X1 U1166 ( .A1(KEYINPUT61), .A2(n1361), .ZN(n1466) );
INV_X1 U1167 ( .A(G119), .ZN(n1361) );
XNOR2_X1 U1168 ( .A(n1259), .B(n1261), .ZN(n1464) );
NAND3_X1 U1169 ( .A1(n1468), .A2(n1469), .A3(n1451), .ZN(n1261) );
NAND3_X1 U1170 ( .A1(G146), .A2(n1324), .A3(G128), .ZN(n1451) );
INV_X1 U1171 ( .A(G143), .ZN(n1324) );
NAND2_X1 U1172 ( .A1(n1470), .A2(n1453), .ZN(n1469) );
INV_X1 U1173 ( .A(G128), .ZN(n1453) );
XOR2_X1 U1174 ( .A(G143), .B(n1471), .Z(n1470) );
NOR2_X1 U1175 ( .A1(G146), .A2(KEYINPUT60), .ZN(n1471) );
NAND3_X1 U1176 ( .A1(n1472), .A2(n1322), .A3(G128), .ZN(n1468) );
INV_X1 U1177 ( .A(G146), .ZN(n1322) );
XOR2_X1 U1178 ( .A(KEYINPUT60), .B(G143), .Z(n1472) );
NAND3_X1 U1179 ( .A1(n1473), .A2(n1474), .A3(n1475), .ZN(n1259) );
OR2_X1 U1180 ( .A1(n1199), .A2(G131), .ZN(n1475) );
NAND2_X1 U1181 ( .A1(KEYINPUT34), .A2(n1476), .ZN(n1474) );
NAND2_X1 U1182 ( .A1(n1477), .A2(G131), .ZN(n1476) );
XNOR2_X1 U1183 ( .A(KEYINPUT17), .B(n1199), .ZN(n1477) );
NAND2_X1 U1184 ( .A1(n1478), .A2(n1479), .ZN(n1473) );
INV_X1 U1185 ( .A(KEYINPUT34), .ZN(n1479) );
NAND2_X1 U1186 ( .A1(n1480), .A2(n1481), .ZN(n1478) );
OR2_X1 U1187 ( .A1(n1199), .A2(KEYINPUT17), .ZN(n1481) );
NAND3_X1 U1188 ( .A1(G131), .A2(n1199), .A3(KEYINPUT17), .ZN(n1480) );
XOR2_X1 U1189 ( .A(n1335), .B(n1330), .Z(n1199) );
INV_X1 U1190 ( .A(G137), .ZN(n1330) );
INV_X1 U1191 ( .A(G134), .ZN(n1335) );
endmodule


