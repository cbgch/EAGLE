//Key = 0011100001111111110001001010000000101110011110111111101011010110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305;

XOR2_X1 U722 ( .A(G107), .B(n996), .Z(G9) );
NOR2_X1 U723 ( .A1(n997), .A2(n998), .ZN(G75) );
NOR4_X1 U724 ( .A1(n999), .A2(n1000), .A3(G953), .A4(n1001), .ZN(n998) );
NOR3_X1 U725 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(n1000) );
NOR2_X1 U726 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
NOR2_X1 U727 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NOR2_X1 U728 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U729 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NOR2_X1 U730 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
NOR3_X1 U731 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1013) );
NOR2_X1 U732 ( .A1(n1018), .A2(n1019), .ZN(n1009) );
NOR2_X1 U733 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR3_X1 U734 ( .A1(n1012), .A2(n1022), .A3(n1019), .ZN(n1005) );
NOR2_X1 U735 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR2_X1 U736 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NAND2_X1 U737 ( .A1(n1027), .A2(n1028), .ZN(n999) );
NAND4_X1 U738 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1028) );
NOR2_X1 U739 ( .A1(n1012), .A2(n1002), .ZN(n1032) );
NAND2_X1 U740 ( .A1(n1033), .A2(n1034), .ZN(n1030) );
XOR2_X1 U741 ( .A(KEYINPUT24), .B(n1035), .Z(n1033) );
NOR2_X1 U742 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR3_X1 U743 ( .A1(n1001), .A2(G953), .A3(G952), .ZN(n997) );
AND4_X1 U744 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1001) );
NOR4_X1 U745 ( .A1(n1019), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1041) );
XOR2_X1 U746 ( .A(n1045), .B(n1046), .Z(n1044) );
XNOR2_X1 U747 ( .A(G472), .B(KEYINPUT18), .ZN(n1046) );
XNOR2_X1 U748 ( .A(n1047), .B(n1048), .ZN(n1043) );
INV_X1 U749 ( .A(n1031), .ZN(n1019) );
NOR2_X1 U750 ( .A1(n1049), .A2(n1050), .ZN(n1040) );
NAND2_X1 U751 ( .A1(n1051), .A2(n1052), .ZN(n1039) );
XNOR2_X1 U752 ( .A(n1053), .B(n1054), .ZN(n1038) );
XOR2_X1 U753 ( .A(n1055), .B(KEYINPUT14), .Z(n1054) );
XOR2_X1 U754 ( .A(n1056), .B(n1057), .Z(G72) );
NOR2_X1 U755 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U756 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND2_X1 U757 ( .A1(n1062), .A2(n1063), .ZN(n1056) );
NAND2_X1 U758 ( .A1(n1064), .A2(n1059), .ZN(n1063) );
XOR2_X1 U759 ( .A(n1065), .B(n1066), .Z(n1064) );
NAND3_X1 U760 ( .A1(G900), .A2(n1066), .A3(G953), .ZN(n1062) );
XOR2_X1 U761 ( .A(n1067), .B(n1068), .Z(n1066) );
XNOR2_X1 U762 ( .A(n1069), .B(G131), .ZN(n1068) );
XNOR2_X1 U763 ( .A(n1070), .B(n1071), .ZN(n1067) );
XOR2_X1 U764 ( .A(n1072), .B(n1073), .Z(G69) );
XOR2_X1 U765 ( .A(n1074), .B(n1075), .Z(n1073) );
NOR2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XNOR2_X1 U767 ( .A(G953), .B(KEYINPUT47), .ZN(n1077) );
INV_X1 U768 ( .A(n1078), .ZN(n1076) );
NOR2_X1 U769 ( .A1(n1079), .A2(n1080), .ZN(n1074) );
XOR2_X1 U770 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND2_X1 U771 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U772 ( .A1(KEYINPUT41), .A2(n1085), .ZN(n1084) );
OR3_X1 U773 ( .A1(n1086), .A2(n1087), .A3(KEYINPUT41), .ZN(n1083) );
NAND2_X1 U774 ( .A1(n1088), .A2(n1089), .ZN(n1081) );
XOR2_X1 U775 ( .A(KEYINPUT27), .B(KEYINPUT21), .Z(n1089) );
NOR2_X1 U776 ( .A1(n1090), .A2(n1059), .ZN(n1079) );
XNOR2_X1 U777 ( .A(G898), .B(KEYINPUT11), .ZN(n1090) );
NOR2_X1 U778 ( .A1(n1091), .A2(n1059), .ZN(n1072) );
NOR2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR2_X1 U780 ( .A1(n1094), .A2(n1095), .ZN(G66) );
XOR2_X1 U781 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U782 ( .A1(n1098), .A2(G217), .ZN(n1096) );
NOR2_X1 U783 ( .A1(n1094), .A2(n1099), .ZN(G63) );
XOR2_X1 U784 ( .A(n1100), .B(n1101), .Z(n1099) );
NAND2_X1 U785 ( .A1(n1098), .A2(G478), .ZN(n1100) );
NOR2_X1 U786 ( .A1(n1094), .A2(n1102), .ZN(G60) );
XOR2_X1 U787 ( .A(n1103), .B(n1104), .Z(n1102) );
NAND2_X1 U788 ( .A1(n1105), .A2(n1098), .ZN(n1103) );
XNOR2_X1 U789 ( .A(G475), .B(KEYINPUT61), .ZN(n1105) );
XOR2_X1 U790 ( .A(n1106), .B(n1107), .Z(G6) );
XNOR2_X1 U791 ( .A(G104), .B(KEYINPUT20), .ZN(n1107) );
NAND3_X1 U792 ( .A1(n1108), .A2(n1109), .A3(n1021), .ZN(n1106) );
XNOR2_X1 U793 ( .A(KEYINPUT55), .B(n1008), .ZN(n1109) );
INV_X1 U794 ( .A(n1029), .ZN(n1008) );
NOR2_X1 U795 ( .A1(n1094), .A2(n1110), .ZN(G57) );
XOR2_X1 U796 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U797 ( .A(n1113), .B(n1114), .Z(n1111) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U799 ( .A(KEYINPUT29), .B(n1117), .Z(n1116) );
NOR2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
AND2_X1 U801 ( .A1(n1119), .A2(n1118), .ZN(n1115) );
NAND2_X1 U802 ( .A1(n1098), .A2(G472), .ZN(n1113) );
NOR2_X1 U803 ( .A1(n1094), .A2(n1120), .ZN(G54) );
XOR2_X1 U804 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U805 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U806 ( .A1(n1098), .A2(G469), .ZN(n1123) );
XNOR2_X1 U807 ( .A(n1125), .B(KEYINPUT13), .ZN(n1121) );
NAND2_X1 U808 ( .A1(KEYINPUT46), .A2(n1126), .ZN(n1125) );
NOR2_X1 U809 ( .A1(n1094), .A2(n1127), .ZN(G51) );
XOR2_X1 U810 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U811 ( .A(n1130), .B(n1131), .Z(n1128) );
NOR2_X1 U812 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XOR2_X1 U813 ( .A(KEYINPUT30), .B(n1134), .Z(n1133) );
NOR4_X1 U814 ( .A1(G953), .A2(n1135), .A3(n1136), .A4(n1092), .ZN(n1134) );
NOR2_X1 U815 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
NOR2_X1 U816 ( .A1(G953), .A2(n1092), .ZN(n1138) );
INV_X1 U817 ( .A(G224), .ZN(n1092) );
NOR2_X1 U818 ( .A1(n1135), .A2(n1136), .ZN(n1137) );
NOR2_X1 U819 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
NAND2_X1 U820 ( .A1(n1098), .A2(n1053), .ZN(n1130) );
INV_X1 U821 ( .A(n1141), .ZN(n1053) );
NOR2_X1 U822 ( .A1(n1142), .A2(n1027), .ZN(n1098) );
NOR2_X1 U823 ( .A1(n1078), .A2(n1065), .ZN(n1027) );
NAND4_X1 U824 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1065) );
NOR4_X1 U825 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1146) );
NAND2_X1 U826 ( .A1(n1151), .A2(n1152), .ZN(n1145) );
NAND2_X1 U827 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND4_X1 U828 ( .A1(n1155), .A2(n1014), .A3(n1021), .A4(n1024), .ZN(n1154) );
XNOR2_X1 U829 ( .A(n1156), .B(KEYINPUT39), .ZN(n1155) );
XNOR2_X1 U830 ( .A(KEYINPUT26), .B(n1157), .ZN(n1153) );
NAND4_X1 U831 ( .A1(n1158), .A2(n1020), .A3(n1159), .A4(n1160), .ZN(n1143) );
NAND4_X1 U832 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1078) );
NOR4_X1 U833 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n996), .ZN(n1164) );
AND3_X1 U834 ( .A1(n1020), .A2(n1029), .A3(n1108), .ZN(n996) );
NAND2_X1 U835 ( .A1(n1021), .A2(n1168), .ZN(n1163) );
NAND2_X1 U836 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND2_X1 U837 ( .A1(n1108), .A2(n1029), .ZN(n1170) );
NAND2_X1 U838 ( .A1(n1171), .A2(n1024), .ZN(n1169) );
AND2_X1 U839 ( .A1(n1172), .A2(G953), .ZN(n1094) );
XNOR2_X1 U840 ( .A(G952), .B(KEYINPUT28), .ZN(n1172) );
XNOR2_X1 U841 ( .A(G146), .B(n1144), .ZN(G48) );
NAND3_X1 U842 ( .A1(n1173), .A2(n1160), .A3(n1174), .ZN(n1144) );
XNOR2_X1 U843 ( .A(n1175), .B(n1150), .ZN(G45) );
AND4_X1 U844 ( .A1(n1176), .A2(n1177), .A3(n1173), .A4(n1042), .ZN(n1150) );
XOR2_X1 U845 ( .A(n1178), .B(n1179), .Z(G42) );
NOR2_X1 U846 ( .A1(n1004), .A2(n1157), .ZN(n1179) );
NAND2_X1 U847 ( .A1(n1174), .A2(n1180), .ZN(n1157) );
AND4_X1 U848 ( .A1(n1014), .A2(n1021), .A3(n1181), .A4(n1182), .ZN(n1174) );
NAND2_X1 U849 ( .A1(KEYINPUT17), .A2(n1183), .ZN(n1178) );
XOR2_X1 U850 ( .A(G137), .B(n1149), .Z(G39) );
AND4_X1 U851 ( .A1(n1014), .A2(n1151), .A3(n1184), .A4(n1185), .ZN(n1149) );
NOR2_X1 U852 ( .A1(n1156), .A2(n1186), .ZN(n1184) );
XNOR2_X1 U853 ( .A(n1069), .B(n1148), .ZN(G36) );
AND3_X1 U854 ( .A1(n1177), .A2(n1020), .A3(n1151), .ZN(n1148) );
INV_X1 U855 ( .A(n1187), .ZN(n1177) );
XNOR2_X1 U856 ( .A(n1188), .B(n1189), .ZN(G33) );
NOR3_X1 U857 ( .A1(n1190), .A2(n1187), .A3(n1004), .ZN(n1189) );
INV_X1 U858 ( .A(n1151), .ZN(n1004) );
NOR2_X1 U859 ( .A1(n1036), .A2(n1050), .ZN(n1151) );
NAND3_X1 U860 ( .A1(n1024), .A2(n1181), .A3(n1014), .ZN(n1187) );
XNOR2_X1 U861 ( .A(n1159), .B(KEYINPUT51), .ZN(n1014) );
XOR2_X1 U862 ( .A(KEYINPUT50), .B(n1021), .Z(n1190) );
XOR2_X1 U863 ( .A(n1191), .B(n1192), .Z(G30) );
NAND2_X1 U864 ( .A1(KEYINPUT34), .A2(G128), .ZN(n1192) );
NAND4_X1 U865 ( .A1(n1020), .A2(n1159), .A3(n1193), .A4(n1194), .ZN(n1191) );
NOR3_X1 U866 ( .A1(n1186), .A2(n1025), .A3(n1156), .ZN(n1194) );
XNOR2_X1 U867 ( .A(n1173), .B(KEYINPUT56), .ZN(n1193) );
XNOR2_X1 U868 ( .A(G101), .B(n1161), .ZN(G3) );
NAND3_X1 U869 ( .A1(n1195), .A2(n1108), .A3(n1024), .ZN(n1161) );
INV_X1 U870 ( .A(n1012), .ZN(n1195) );
XNOR2_X1 U871 ( .A(n1147), .B(n1196), .ZN(G27) );
XNOR2_X1 U872 ( .A(G125), .B(KEYINPUT7), .ZN(n1196) );
AND4_X1 U873 ( .A1(n1158), .A2(n1021), .A3(n1031), .A4(n1180), .ZN(n1147) );
NOR3_X1 U874 ( .A1(n1156), .A2(n1025), .A3(n1034), .ZN(n1158) );
INV_X1 U875 ( .A(n1173), .ZN(n1034) );
INV_X1 U876 ( .A(n1181), .ZN(n1156) );
NAND2_X1 U877 ( .A1(n1197), .A2(n1002), .ZN(n1181) );
NAND4_X1 U878 ( .A1(G953), .A2(G902), .A3(n1198), .A4(n1061), .ZN(n1197) );
INV_X1 U879 ( .A(G900), .ZN(n1061) );
NAND2_X1 U880 ( .A1(n1199), .A2(n1200), .ZN(G24) );
OR2_X1 U881 ( .A1(n1162), .A2(G122), .ZN(n1200) );
XOR2_X1 U882 ( .A(n1201), .B(KEYINPUT8), .Z(n1199) );
NAND2_X1 U883 ( .A1(G122), .A2(n1162), .ZN(n1201) );
NAND4_X1 U884 ( .A1(n1171), .A2(n1029), .A3(n1176), .A4(n1042), .ZN(n1162) );
INV_X1 U885 ( .A(n1202), .ZN(n1176) );
NOR2_X1 U886 ( .A1(n1182), .A2(n1026), .ZN(n1029) );
INV_X1 U887 ( .A(n1180), .ZN(n1026) );
XOR2_X1 U888 ( .A(G119), .B(n1167), .Z(G21) );
AND3_X1 U889 ( .A1(n1185), .A2(n1160), .A3(n1171), .ZN(n1167) );
XNOR2_X1 U890 ( .A(G116), .B(n1203), .ZN(G18) );
NAND2_X1 U891 ( .A1(KEYINPUT37), .A2(n1166), .ZN(n1203) );
AND3_X1 U892 ( .A1(n1024), .A2(n1020), .A3(n1171), .ZN(n1166) );
NOR2_X1 U893 ( .A1(n1042), .A2(n1202), .ZN(n1020) );
XNOR2_X1 U894 ( .A(G113), .B(n1204), .ZN(G15) );
NAND4_X1 U895 ( .A1(n1205), .A2(KEYINPUT42), .A3(n1021), .A4(n1171), .ZN(n1204) );
AND2_X1 U896 ( .A1(n1031), .A2(n1206), .ZN(n1171) );
NOR2_X1 U897 ( .A1(n1015), .A2(n1207), .ZN(n1031) );
NOR2_X1 U898 ( .A1(n1017), .A2(n1016), .ZN(n1207) );
INV_X1 U899 ( .A(n1208), .ZN(n1016) );
INV_X1 U900 ( .A(G221), .ZN(n1017) );
AND2_X1 U901 ( .A1(n1209), .A2(n1042), .ZN(n1021) );
XNOR2_X1 U902 ( .A(n1202), .B(KEYINPUT10), .ZN(n1209) );
XNOR2_X1 U903 ( .A(n1024), .B(KEYINPUT49), .ZN(n1205) );
NOR2_X1 U904 ( .A1(n1182), .A2(n1186), .ZN(n1024) );
INV_X1 U905 ( .A(n1160), .ZN(n1186) );
XOR2_X1 U906 ( .A(n1180), .B(KEYINPUT62), .Z(n1160) );
INV_X1 U907 ( .A(n1025), .ZN(n1182) );
XOR2_X1 U908 ( .A(G110), .B(n1165), .Z(G12) );
AND3_X1 U909 ( .A1(n1108), .A2(n1180), .A3(n1185), .ZN(n1165) );
NOR2_X1 U910 ( .A1(n1012), .A2(n1025), .ZN(n1185) );
NOR2_X1 U911 ( .A1(n1210), .A2(n1049), .ZN(n1025) );
NOR2_X1 U912 ( .A1(n1052), .A2(n1051), .ZN(n1049) );
AND2_X1 U913 ( .A1(n1211), .A2(n1052), .ZN(n1210) );
NAND2_X1 U914 ( .A1(n1212), .A2(n1097), .ZN(n1052) );
XNOR2_X1 U915 ( .A(n1213), .B(n1214), .ZN(n1097) );
XOR2_X1 U916 ( .A(G110), .B(n1215), .Z(n1214) );
XOR2_X1 U917 ( .A(KEYINPUT2), .B(G119), .Z(n1215) );
XOR2_X1 U918 ( .A(n1216), .B(n1071), .Z(n1213) );
XNOR2_X1 U919 ( .A(n1139), .B(n1217), .ZN(n1071) );
XNOR2_X1 U920 ( .A(n1183), .B(G137), .ZN(n1217) );
XOR2_X1 U921 ( .A(n1218), .B(n1219), .Z(n1216) );
NOR2_X1 U922 ( .A1(n1220), .A2(KEYINPUT63), .ZN(n1219) );
AND3_X1 U923 ( .A1(G221), .A2(n1059), .A3(G234), .ZN(n1220) );
XOR2_X1 U924 ( .A(KEYINPUT58), .B(n1051), .Z(n1211) );
AND2_X1 U925 ( .A1(G217), .A2(n1221), .ZN(n1051) );
XNOR2_X1 U926 ( .A(KEYINPUT57), .B(n1208), .ZN(n1221) );
NAND2_X1 U927 ( .A1(n1222), .A2(n1202), .ZN(n1012) );
XNOR2_X1 U928 ( .A(n1223), .B(n1048), .ZN(n1202) );
AND2_X1 U929 ( .A1(n1101), .A2(n1212), .ZN(n1048) );
XOR2_X1 U930 ( .A(n1224), .B(n1225), .Z(n1101) );
NOR2_X1 U931 ( .A1(KEYINPUT40), .A2(n1226), .ZN(n1225) );
XOR2_X1 U932 ( .A(n1227), .B(n1228), .Z(n1226) );
XOR2_X1 U933 ( .A(G116), .B(n1229), .Z(n1228) );
XNOR2_X1 U934 ( .A(n1069), .B(G122), .ZN(n1229) );
INV_X1 U935 ( .A(G134), .ZN(n1069) );
XOR2_X1 U936 ( .A(n1230), .B(G107), .Z(n1227) );
NAND3_X1 U937 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1230) );
NAND2_X1 U938 ( .A1(G143), .A2(n1234), .ZN(n1233) );
INV_X1 U939 ( .A(G128), .ZN(n1234) );
NAND2_X1 U940 ( .A1(n1235), .A2(n1236), .ZN(n1232) );
INV_X1 U941 ( .A(KEYINPUT12), .ZN(n1236) );
NAND2_X1 U942 ( .A1(n1237), .A2(n1175), .ZN(n1235) );
XNOR2_X1 U943 ( .A(KEYINPUT52), .B(G128), .ZN(n1237) );
NAND2_X1 U944 ( .A1(KEYINPUT12), .A2(n1238), .ZN(n1231) );
NAND2_X1 U945 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
OR2_X1 U946 ( .A1(G128), .A2(KEYINPUT52), .ZN(n1240) );
NAND3_X1 U947 ( .A1(G128), .A2(n1175), .A3(KEYINPUT52), .ZN(n1239) );
NAND3_X1 U948 ( .A1(n1241), .A2(n1059), .A3(G217), .ZN(n1224) );
XOR2_X1 U949 ( .A(KEYINPUT1), .B(G234), .Z(n1241) );
NAND2_X1 U950 ( .A1(KEYINPUT43), .A2(n1047), .ZN(n1223) );
INV_X1 U951 ( .A(G478), .ZN(n1047) );
XOR2_X1 U952 ( .A(KEYINPUT3), .B(n1042), .Z(n1222) );
XNOR2_X1 U953 ( .A(n1242), .B(G475), .ZN(n1042) );
NAND2_X1 U954 ( .A1(n1104), .A2(n1212), .ZN(n1242) );
XOR2_X1 U955 ( .A(n1243), .B(n1244), .Z(n1104) );
XOR2_X1 U956 ( .A(n1245), .B(n1246), .Z(n1244) );
XOR2_X1 U957 ( .A(G122), .B(G104), .Z(n1246) );
NOR2_X1 U958 ( .A1(KEYINPUT31), .A2(n1247), .ZN(n1245) );
XOR2_X1 U959 ( .A(n1248), .B(n1249), .Z(n1247) );
XOR2_X1 U960 ( .A(n1250), .B(n1251), .Z(n1249) );
NAND2_X1 U961 ( .A1(KEYINPUT4), .A2(G125), .ZN(n1250) );
XNOR2_X1 U962 ( .A(G140), .B(n1252), .ZN(n1248) );
XOR2_X1 U963 ( .A(KEYINPUT2), .B(KEYINPUT0), .Z(n1252) );
XOR2_X1 U964 ( .A(n1253), .B(n1254), .Z(n1243) );
NAND3_X1 U965 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1253) );
NAND2_X1 U966 ( .A1(KEYINPUT23), .A2(n1258), .ZN(n1257) );
NAND3_X1 U967 ( .A1(n1259), .A2(n1260), .A3(n1188), .ZN(n1256) );
INV_X1 U968 ( .A(KEYINPUT23), .ZN(n1260) );
OR2_X1 U969 ( .A1(n1188), .A2(n1259), .ZN(n1255) );
NOR2_X1 U970 ( .A1(KEYINPUT60), .A2(n1258), .ZN(n1259) );
XNOR2_X1 U971 ( .A(n1261), .B(G143), .ZN(n1258) );
NAND2_X1 U972 ( .A1(n1262), .A2(G214), .ZN(n1261) );
XNOR2_X1 U973 ( .A(n1045), .B(n1263), .ZN(n1180) );
NOR2_X1 U974 ( .A1(G472), .A2(KEYINPUT19), .ZN(n1263) );
NAND2_X1 U975 ( .A1(n1264), .A2(n1212), .ZN(n1045) );
XOR2_X1 U976 ( .A(n1265), .B(n1266), .Z(n1264) );
XNOR2_X1 U977 ( .A(KEYINPUT45), .B(n1118), .ZN(n1266) );
XOR2_X1 U978 ( .A(n1267), .B(n1254), .Z(n1118) );
XNOR2_X1 U979 ( .A(G116), .B(G119), .ZN(n1267) );
XNOR2_X1 U980 ( .A(n1119), .B(n1112), .ZN(n1265) );
XNOR2_X1 U981 ( .A(n1268), .B(G101), .ZN(n1112) );
NAND2_X1 U982 ( .A1(n1262), .A2(G210), .ZN(n1268) );
NOR2_X1 U983 ( .A1(G953), .A2(G237), .ZN(n1262) );
XNOR2_X1 U984 ( .A(n1269), .B(KEYINPUT59), .ZN(n1119) );
AND2_X1 U985 ( .A1(n1206), .A2(n1159), .ZN(n1108) );
AND2_X1 U986 ( .A1(n1015), .A2(n1270), .ZN(n1159) );
NAND2_X1 U987 ( .A1(G221), .A2(n1208), .ZN(n1270) );
NAND2_X1 U988 ( .A1(G234), .A2(n1142), .ZN(n1208) );
XNOR2_X1 U989 ( .A(n1271), .B(G469), .ZN(n1015) );
NAND2_X1 U990 ( .A1(n1272), .A2(n1212), .ZN(n1271) );
XNOR2_X1 U991 ( .A(n1124), .B(n1126), .ZN(n1272) );
XOR2_X1 U992 ( .A(n1273), .B(n1274), .Z(n1124) );
XNOR2_X1 U993 ( .A(n1183), .B(G110), .ZN(n1274) );
INV_X1 U994 ( .A(G140), .ZN(n1183) );
XOR2_X1 U995 ( .A(n1269), .B(n1275), .Z(n1273) );
NOR2_X1 U996 ( .A1(G953), .A2(n1060), .ZN(n1275) );
INV_X1 U997 ( .A(G227), .ZN(n1060) );
XNOR2_X1 U998 ( .A(n1276), .B(n1277), .ZN(n1269) );
INV_X1 U999 ( .A(n1070), .ZN(n1277) );
NAND2_X1 U1000 ( .A1(n1278), .A2(n1279), .ZN(n1276) );
NAND2_X1 U1001 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U1002 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U1003 ( .A1(KEYINPUT44), .A2(G131), .ZN(n1283) );
INV_X1 U1004 ( .A(KEYINPUT35), .ZN(n1282) );
NAND2_X1 U1005 ( .A1(n1284), .A2(n1188), .ZN(n1278) );
INV_X1 U1006 ( .A(G131), .ZN(n1188) );
NAND2_X1 U1007 ( .A1(KEYINPUT44), .A2(n1285), .ZN(n1284) );
OR2_X1 U1008 ( .A1(n1280), .A2(KEYINPUT35), .ZN(n1285) );
XNOR2_X1 U1009 ( .A(G134), .B(n1286), .ZN(n1280) );
XOR2_X1 U1010 ( .A(KEYINPUT6), .B(G137), .Z(n1286) );
AND2_X1 U1011 ( .A1(n1173), .A2(n1287), .ZN(n1206) );
NAND2_X1 U1012 ( .A1(n1002), .A2(n1288), .ZN(n1287) );
NAND4_X1 U1013 ( .A1(G953), .A2(G902), .A3(n1198), .A4(n1093), .ZN(n1288) );
INV_X1 U1014 ( .A(G898), .ZN(n1093) );
NAND3_X1 U1015 ( .A1(n1198), .A2(n1059), .A3(G952), .ZN(n1002) );
NAND2_X1 U1016 ( .A1(G234), .A2(G237), .ZN(n1198) );
NOR2_X1 U1017 ( .A1(n1289), .A2(n1050), .ZN(n1173) );
INV_X1 U1018 ( .A(n1037), .ZN(n1050) );
NAND2_X1 U1019 ( .A1(G214), .A2(n1290), .ZN(n1037) );
INV_X1 U1020 ( .A(n1036), .ZN(n1289) );
XNOR2_X1 U1021 ( .A(n1055), .B(n1291), .ZN(n1036) );
NOR2_X1 U1022 ( .A1(KEYINPUT33), .A2(n1141), .ZN(n1291) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1290), .ZN(n1141) );
NAND2_X1 U1024 ( .A1(n1292), .A2(n1142), .ZN(n1290) );
INV_X1 U1025 ( .A(G902), .ZN(n1142) );
XOR2_X1 U1026 ( .A(KEYINPUT9), .B(G237), .Z(n1292) );
NAND2_X1 U1027 ( .A1(n1293), .A2(n1212), .ZN(n1055) );
XNOR2_X1 U1028 ( .A(G902), .B(KEYINPUT22), .ZN(n1212) );
XOR2_X1 U1029 ( .A(n1294), .B(n1295), .Z(n1293) );
NOR2_X1 U1030 ( .A1(KEYINPUT53), .A2(n1129), .ZN(n1295) );
XOR2_X1 U1031 ( .A(n1085), .B(n1088), .Z(n1129) );
XOR2_X1 U1032 ( .A(n1296), .B(G110), .Z(n1088) );
NAND2_X1 U1033 ( .A1(KEYINPUT36), .A2(G122), .ZN(n1296) );
XOR2_X1 U1034 ( .A(n1086), .B(n1087), .Z(n1085) );
XNOR2_X1 U1035 ( .A(n1126), .B(KEYINPUT16), .ZN(n1087) );
XNOR2_X1 U1036 ( .A(G101), .B(n1297), .ZN(n1126) );
XOR2_X1 U1037 ( .A(G107), .B(G104), .Z(n1297) );
XOR2_X1 U1038 ( .A(n1298), .B(n1299), .Z(n1086) );
XOR2_X1 U1039 ( .A(n1300), .B(n1254), .Z(n1299) );
XOR2_X1 U1040 ( .A(G113), .B(KEYINPUT38), .Z(n1254) );
NOR2_X1 U1041 ( .A1(G119), .A2(KEYINPUT32), .ZN(n1300) );
XNOR2_X1 U1042 ( .A(G116), .B(KEYINPUT25), .ZN(n1298) );
XOR2_X1 U1043 ( .A(n1301), .B(n1302), .Z(n1294) );
NOR2_X1 U1044 ( .A1(n1135), .A2(n1303), .ZN(n1302) );
NOR2_X1 U1045 ( .A1(n1140), .A2(n1304), .ZN(n1303) );
XNOR2_X1 U1046 ( .A(n1305), .B(n1139), .ZN(n1304) );
XNOR2_X1 U1047 ( .A(KEYINPUT48), .B(KEYINPUT15), .ZN(n1305) );
AND2_X1 U1048 ( .A1(n1140), .A2(n1139), .ZN(n1135) );
INV_X1 U1049 ( .A(G125), .ZN(n1139) );
XNOR2_X1 U1050 ( .A(n1070), .B(KEYINPUT59), .ZN(n1140) );
XOR2_X1 U1051 ( .A(n1218), .B(n1175), .Z(n1070) );
INV_X1 U1052 ( .A(G143), .ZN(n1175) );
XNOR2_X1 U1053 ( .A(G128), .B(n1251), .ZN(n1218) );
XOR2_X1 U1054 ( .A(G146), .B(KEYINPUT5), .Z(n1251) );
NAND3_X1 U1055 ( .A1(G224), .A2(n1059), .A3(KEYINPUT54), .ZN(n1301) );
INV_X1 U1056 ( .A(G953), .ZN(n1059) );
endmodule


