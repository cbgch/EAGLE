//Key = 1110111111110110110110010110101000100011011001000110011101000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
n1461, n1462, n1463, n1464, n1465, n1466, n1467;

XNOR2_X1 U800 ( .A(n1111), .B(n1112), .ZN(G9) );
NAND2_X1 U801 ( .A1(KEYINPUT39), .A2(G107), .ZN(n1112) );
NOR2_X1 U802 ( .A1(n1113), .A2(n1114), .ZN(G75) );
NOR3_X1 U803 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
NOR2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NOR2_X1 U805 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
NOR3_X1 U806 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1121) );
NOR2_X1 U807 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR2_X1 U808 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
NOR2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR2_X1 U811 ( .A1(n1133), .A2(n1134), .ZN(n1129) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NOR3_X1 U813 ( .A1(n1132), .A2(n1137), .A3(n1134), .ZN(n1125) );
NOR2_X1 U814 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR2_X1 U815 ( .A1(n1131), .A2(n1140), .ZN(n1138) );
NOR3_X1 U816 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1131) );
NOR4_X1 U817 ( .A1(n1144), .A2(n1134), .A3(n1128), .A4(n1132), .ZN(n1120) );
INV_X1 U818 ( .A(n1145), .ZN(n1128) );
NOR2_X1 U819 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
NOR2_X1 U820 ( .A1(n1122), .A2(n1148), .ZN(n1146) );
NOR2_X1 U821 ( .A1(G952), .A2(n1117), .ZN(n1113) );
NAND2_X1 U822 ( .A1(n1149), .A2(n1150), .ZN(n1117) );
NAND4_X1 U823 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
NOR4_X1 U824 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1154) );
AND3_X1 U825 ( .A1(KEYINPUT25), .A2(n1159), .A3(G478), .ZN(n1158) );
NOR2_X1 U826 ( .A1(KEYINPUT25), .A2(G478), .ZN(n1157) );
XOR2_X1 U827 ( .A(n1160), .B(n1161), .Z(n1156) );
NAND3_X1 U828 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1155) );
XOR2_X1 U829 ( .A(KEYINPUT45), .B(n1165), .Z(n1163) );
NOR3_X1 U830 ( .A1(n1166), .A2(n1123), .A3(n1167), .ZN(n1153) );
NAND2_X1 U831 ( .A1(n1168), .A2(n1169), .ZN(n1151) );
XOR2_X1 U832 ( .A(n1170), .B(n1171), .Z(G72) );
NOR2_X1 U833 ( .A1(n1172), .A2(n1149), .ZN(n1171) );
AND2_X1 U834 ( .A1(G227), .A2(G900), .ZN(n1172) );
NAND2_X1 U835 ( .A1(n1173), .A2(n1174), .ZN(n1170) );
NAND2_X1 U836 ( .A1(n1175), .A2(n1149), .ZN(n1174) );
XOR2_X1 U837 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U838 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
OR3_X1 U839 ( .A1(n1176), .A2(n1180), .A3(n1149), .ZN(n1173) );
NAND2_X1 U840 ( .A1(n1181), .A2(n1182), .ZN(n1176) );
NAND3_X1 U841 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1182) );
XOR2_X1 U842 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U843 ( .A1(G125), .A2(n1188), .ZN(n1187) );
NAND2_X1 U844 ( .A1(n1189), .A2(n1190), .ZN(n1181) );
NAND2_X1 U845 ( .A1(n1183), .A2(n1184), .ZN(n1190) );
INV_X1 U846 ( .A(KEYINPUT24), .ZN(n1184) );
XOR2_X1 U847 ( .A(n1186), .B(n1191), .Z(n1189) );
NOR2_X1 U848 ( .A1(n1192), .A2(n1188), .ZN(n1191) );
INV_X1 U849 ( .A(KEYINPUT8), .ZN(n1188) );
NAND2_X1 U850 ( .A1(n1193), .A2(n1194), .ZN(n1186) );
NAND2_X1 U851 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XOR2_X1 U852 ( .A(KEYINPUT4), .B(n1197), .Z(n1193) );
NOR2_X1 U853 ( .A1(n1195), .A2(n1196), .ZN(n1197) );
XOR2_X1 U854 ( .A(n1198), .B(n1199), .Z(n1196) );
OR2_X1 U855 ( .A1(G131), .A2(KEYINPUT18), .ZN(n1199) );
NAND2_X1 U856 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
NAND2_X1 U857 ( .A1(G134), .A2(n1202), .ZN(n1201) );
XOR2_X1 U858 ( .A(KEYINPUT19), .B(n1203), .Z(n1200) );
NOR2_X1 U859 ( .A1(G134), .A2(n1202), .ZN(n1203) );
NAND2_X1 U860 ( .A1(n1204), .A2(n1205), .ZN(G69) );
NAND2_X1 U861 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U862 ( .A1(n1208), .A2(n1209), .ZN(n1206) );
INV_X1 U863 ( .A(n1210), .ZN(n1208) );
NAND2_X1 U864 ( .A1(n1211), .A2(n1209), .ZN(n1204) );
NAND2_X1 U865 ( .A1(G953), .A2(n1212), .ZN(n1209) );
INV_X1 U866 ( .A(n1207), .ZN(n1211) );
NAND2_X1 U867 ( .A1(n1213), .A2(n1214), .ZN(n1207) );
XOR2_X1 U868 ( .A(n1215), .B(n1216), .Z(n1214) );
NOR3_X1 U869 ( .A1(n1217), .A2(n1210), .A3(n1218), .ZN(n1216) );
NOR2_X1 U870 ( .A1(n1219), .A2(n1220), .ZN(n1217) );
INV_X1 U871 ( .A(n1221), .ZN(n1220) );
XNOR2_X1 U872 ( .A(n1222), .B(KEYINPUT40), .ZN(n1219) );
NOR2_X1 U873 ( .A1(G953), .A2(n1223), .ZN(n1215) );
NOR3_X1 U874 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1223) );
XOR2_X1 U875 ( .A(n1227), .B(KEYINPUT34), .Z(n1226) );
XOR2_X1 U876 ( .A(KEYINPUT52), .B(KEYINPUT2), .Z(n1213) );
NOR2_X1 U877 ( .A1(n1228), .A2(n1229), .ZN(G66) );
XNOR2_X1 U878 ( .A(n1230), .B(n1231), .ZN(n1229) );
NOR2_X1 U879 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
INV_X1 U880 ( .A(G217), .ZN(n1232) );
NOR2_X1 U881 ( .A1(n1228), .A2(n1234), .ZN(G63) );
XNOR2_X1 U882 ( .A(n1235), .B(n1236), .ZN(n1234) );
NOR2_X1 U883 ( .A1(n1237), .A2(n1233), .ZN(n1236) );
NOR2_X1 U884 ( .A1(n1228), .A2(n1238), .ZN(G60) );
XOR2_X1 U885 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U886 ( .A(KEYINPUT7), .B(n1241), .Z(n1240) );
NOR2_X1 U887 ( .A1(n1242), .A2(n1233), .ZN(n1241) );
INV_X1 U888 ( .A(G475), .ZN(n1242) );
XOR2_X1 U889 ( .A(G104), .B(n1243), .Z(G6) );
NOR2_X1 U890 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
NOR2_X1 U891 ( .A1(n1228), .A2(n1246), .ZN(G57) );
XOR2_X1 U892 ( .A(n1247), .B(n1248), .Z(n1246) );
XNOR2_X1 U893 ( .A(n1249), .B(n1250), .ZN(n1248) );
NAND2_X1 U894 ( .A1(KEYINPUT57), .A2(n1251), .ZN(n1249) );
XOR2_X1 U895 ( .A(n1252), .B(n1253), .Z(n1247) );
NOR2_X1 U896 ( .A1(KEYINPUT56), .A2(n1254), .ZN(n1253) );
NAND3_X1 U897 ( .A1(n1255), .A2(n1256), .A3(G472), .ZN(n1252) );
NAND2_X1 U898 ( .A1(KEYINPUT17), .A2(n1233), .ZN(n1256) );
NAND2_X1 U899 ( .A1(n1257), .A2(n1258), .ZN(n1255) );
INV_X1 U900 ( .A(KEYINPUT17), .ZN(n1258) );
NAND2_X1 U901 ( .A1(n1259), .A2(G902), .ZN(n1257) );
NOR3_X1 U902 ( .A1(n1228), .A2(n1260), .A3(n1261), .ZN(G54) );
NOR2_X1 U903 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XOR2_X1 U904 ( .A(n1264), .B(n1265), .Z(n1263) );
OR2_X1 U905 ( .A1(n1266), .A2(KEYINPUT12), .ZN(n1264) );
NOR2_X1 U906 ( .A1(n1267), .A2(n1268), .ZN(n1260) );
XOR2_X1 U907 ( .A(n1269), .B(n1265), .Z(n1268) );
XNOR2_X1 U908 ( .A(n1270), .B(n1271), .ZN(n1265) );
XOR2_X1 U909 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U910 ( .A(KEYINPUT30), .B(n1274), .Z(n1273) );
NOR2_X1 U911 ( .A1(n1160), .A2(n1233), .ZN(n1272) );
XOR2_X1 U912 ( .A(n1195), .B(n1254), .Z(n1270) );
NAND2_X1 U913 ( .A1(n1266), .A2(n1275), .ZN(n1269) );
INV_X1 U914 ( .A(KEYINPUT12), .ZN(n1275) );
XNOR2_X1 U915 ( .A(n1276), .B(n1277), .ZN(n1266) );
NOR2_X1 U916 ( .A1(KEYINPUT51), .A2(n1183), .ZN(n1277) );
INV_X1 U917 ( .A(n1262), .ZN(n1267) );
NOR2_X1 U918 ( .A1(n1228), .A2(n1278), .ZN(G51) );
XOR2_X1 U919 ( .A(n1279), .B(n1280), .Z(n1278) );
NOR2_X1 U920 ( .A1(n1281), .A2(n1233), .ZN(n1280) );
NAND2_X1 U921 ( .A1(G902), .A2(n1115), .ZN(n1233) );
INV_X1 U922 ( .A(n1259), .ZN(n1115) );
NOR4_X1 U923 ( .A1(n1282), .A2(n1179), .A3(n1283), .A4(n1224), .ZN(n1259) );
NAND4_X1 U924 ( .A1(n1284), .A2(n1285), .A3(n1286), .A4(n1287), .ZN(n1224) );
NOR3_X1 U925 ( .A1(n1111), .A2(n1288), .A3(n1289), .ZN(n1287) );
INV_X1 U926 ( .A(n1290), .ZN(n1288) );
AND3_X1 U927 ( .A1(n1135), .A2(n1291), .A3(n1292), .ZN(n1111) );
NAND2_X1 U928 ( .A1(n1293), .A2(n1139), .ZN(n1286) );
XOR2_X1 U929 ( .A(n1245), .B(KEYINPUT6), .Z(n1293) );
NAND4_X1 U930 ( .A1(n1136), .A2(n1291), .A3(n1147), .A4(n1294), .ZN(n1245) );
NAND2_X1 U931 ( .A1(n1227), .A2(n1295), .ZN(n1283) );
XOR2_X1 U932 ( .A(n1225), .B(KEYINPUT50), .Z(n1295) );
INV_X1 U933 ( .A(n1296), .ZN(n1225) );
NAND4_X1 U934 ( .A1(n1297), .A2(n1298), .A3(n1299), .A4(n1300), .ZN(n1179) );
NAND3_X1 U935 ( .A1(n1136), .A2(n1301), .A3(n1142), .ZN(n1297) );
XNOR2_X1 U936 ( .A(n1178), .B(KEYINPUT9), .ZN(n1282) );
NAND4_X1 U937 ( .A1(n1302), .A2(n1303), .A3(n1304), .A4(n1305), .ZN(n1178) );
NAND3_X1 U938 ( .A1(n1306), .A2(n1135), .A3(n1307), .ZN(n1302) );
NOR2_X1 U939 ( .A1(n1308), .A2(n1309), .ZN(n1279) );
XOR2_X1 U940 ( .A(n1310), .B(KEYINPUT20), .Z(n1309) );
NAND2_X1 U941 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NOR2_X1 U942 ( .A1(n1311), .A2(n1312), .ZN(n1308) );
XOR2_X1 U943 ( .A(n1313), .B(KEYINPUT36), .Z(n1311) );
NOR2_X1 U944 ( .A1(n1149), .A2(G952), .ZN(n1228) );
XOR2_X1 U945 ( .A(n1314), .B(n1298), .Z(G48) );
NAND3_X1 U946 ( .A1(n1307), .A2(n1306), .A3(n1136), .ZN(n1298) );
XNOR2_X1 U947 ( .A(G143), .B(n1299), .ZN(G45) );
NAND4_X1 U948 ( .A1(n1141), .A2(n1307), .A3(n1315), .A4(n1316), .ZN(n1299) );
XOR2_X1 U949 ( .A(n1183), .B(n1317), .Z(G42) );
NAND3_X1 U950 ( .A1(n1301), .A2(n1318), .A3(n1136), .ZN(n1317) );
XOR2_X1 U951 ( .A(KEYINPUT48), .B(n1142), .Z(n1318) );
XOR2_X1 U952 ( .A(n1202), .B(n1300), .Z(G39) );
NAND3_X1 U953 ( .A1(n1306), .A2(n1301), .A3(n1319), .ZN(n1300) );
XOR2_X1 U954 ( .A(n1303), .B(n1320), .Z(G36) );
NAND2_X1 U955 ( .A1(KEYINPUT11), .A2(G134), .ZN(n1320) );
NAND3_X1 U956 ( .A1(n1301), .A2(n1135), .A3(n1141), .ZN(n1303) );
XOR2_X1 U957 ( .A(n1321), .B(n1304), .Z(G33) );
NAND3_X1 U958 ( .A1(n1141), .A2(n1301), .A3(n1136), .ZN(n1304) );
AND3_X1 U959 ( .A1(n1147), .A2(n1322), .A3(n1145), .ZN(n1301) );
NOR2_X1 U960 ( .A1(n1140), .A2(n1143), .ZN(n1145) );
INV_X1 U961 ( .A(n1152), .ZN(n1143) );
XOR2_X1 U962 ( .A(n1323), .B(n1324), .Z(G30) );
NAND3_X1 U963 ( .A1(n1307), .A2(n1135), .A3(n1325), .ZN(n1324) );
XNOR2_X1 U964 ( .A(n1306), .B(KEYINPUT13), .ZN(n1325) );
AND3_X1 U965 ( .A1(n1139), .A2(n1322), .A3(n1147), .ZN(n1307) );
XOR2_X1 U966 ( .A(n1326), .B(n1227), .Z(G3) );
NAND3_X1 U967 ( .A1(n1319), .A2(n1292), .A3(n1141), .ZN(n1227) );
XOR2_X1 U968 ( .A(n1192), .B(n1305), .Z(G27) );
NAND4_X1 U969 ( .A1(n1322), .A2(n1148), .A3(n1327), .A4(n1328), .ZN(n1305) );
AND3_X1 U970 ( .A1(n1142), .A2(n1139), .A3(n1136), .ZN(n1328) );
NAND2_X1 U971 ( .A1(n1119), .A2(n1329), .ZN(n1322) );
NAND4_X1 U972 ( .A1(G902), .A2(G953), .A3(n1330), .A4(n1180), .ZN(n1329) );
INV_X1 U973 ( .A(G900), .ZN(n1180) );
XNOR2_X1 U974 ( .A(G122), .B(n1284), .ZN(G24) );
NAND4_X1 U975 ( .A1(n1331), .A2(n1291), .A3(n1315), .A4(n1316), .ZN(n1284) );
INV_X1 U976 ( .A(n1134), .ZN(n1291) );
NAND2_X1 U977 ( .A1(n1332), .A2(n1333), .ZN(n1134) );
XOR2_X1 U978 ( .A(n1334), .B(KEYINPUT44), .Z(n1332) );
XOR2_X1 U979 ( .A(n1335), .B(n1285), .Z(G21) );
NAND3_X1 U980 ( .A1(n1319), .A2(n1306), .A3(n1331), .ZN(n1285) );
NOR2_X1 U981 ( .A1(n1334), .A2(n1333), .ZN(n1306) );
XOR2_X1 U982 ( .A(G116), .B(n1289), .Z(G18) );
AND3_X1 U983 ( .A1(n1141), .A2(n1135), .A3(n1331), .ZN(n1289) );
NOR2_X1 U984 ( .A1(n1315), .A2(n1336), .ZN(n1135) );
INV_X1 U985 ( .A(n1162), .ZN(n1315) );
XOR2_X1 U986 ( .A(n1337), .B(G113), .Z(G15) );
NAND2_X1 U987 ( .A1(KEYINPUT16), .A2(n1296), .ZN(n1337) );
NAND3_X1 U988 ( .A1(n1136), .A2(n1141), .A3(n1331), .ZN(n1296) );
AND4_X1 U989 ( .A1(n1139), .A2(n1327), .A3(n1294), .A4(n1148), .ZN(n1331) );
NOR2_X1 U990 ( .A1(n1165), .A2(n1334), .ZN(n1141) );
NOR2_X1 U991 ( .A1(n1316), .A2(n1162), .ZN(n1136) );
INV_X1 U992 ( .A(n1336), .ZN(n1316) );
XOR2_X1 U993 ( .A(n1276), .B(n1290), .Z(G12) );
NAND3_X1 U994 ( .A1(n1319), .A2(n1292), .A3(n1142), .ZN(n1290) );
AND2_X1 U995 ( .A1(n1334), .A2(n1165), .ZN(n1142) );
INV_X1 U996 ( .A(n1333), .ZN(n1165) );
XOR2_X1 U997 ( .A(n1338), .B(n1339), .Z(n1333) );
NOR2_X1 U998 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
XOR2_X1 U999 ( .A(KEYINPUT5), .B(G217), .Z(n1341) );
INV_X1 U1000 ( .A(n1342), .ZN(n1340) );
NAND2_X1 U1001 ( .A1(n1230), .A2(n1343), .ZN(n1338) );
XNOR2_X1 U1002 ( .A(n1344), .B(n1345), .ZN(n1230) );
XOR2_X1 U1003 ( .A(n1346), .B(n1347), .Z(n1345) );
NAND3_X1 U1004 ( .A1(G234), .A2(n1149), .A3(G221), .ZN(n1347) );
NAND3_X1 U1005 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1346) );
NAND2_X1 U1006 ( .A1(G128), .A2(n1351), .ZN(n1350) );
NAND3_X1 U1007 ( .A1(n1352), .A2(n1323), .A3(KEYINPUT14), .ZN(n1349) );
INV_X1 U1008 ( .A(n1351), .ZN(n1352) );
NAND2_X1 U1009 ( .A1(KEYINPUT63), .A2(n1335), .ZN(n1351) );
OR2_X1 U1010 ( .A1(n1335), .A2(KEYINPUT14), .ZN(n1348) );
INV_X1 U1011 ( .A(G119), .ZN(n1335) );
XOR2_X1 U1012 ( .A(n1353), .B(n1354), .Z(n1344) );
XOR2_X1 U1013 ( .A(G137), .B(G110), .Z(n1354) );
NAND2_X1 U1014 ( .A1(n1355), .A2(KEYINPUT61), .ZN(n1353) );
XOR2_X1 U1015 ( .A(n1356), .B(n1357), .Z(n1355) );
XOR2_X1 U1016 ( .A(G146), .B(G140), .Z(n1357) );
NAND2_X1 U1017 ( .A1(KEYINPUT28), .A2(n1358), .ZN(n1356) );
XOR2_X1 U1018 ( .A(KEYINPUT0), .B(G125), .Z(n1358) );
XOR2_X1 U1019 ( .A(n1164), .B(KEYINPUT46), .Z(n1334) );
XOR2_X1 U1020 ( .A(n1359), .B(G472), .Z(n1164) );
NAND2_X1 U1021 ( .A1(n1360), .A2(n1343), .ZN(n1359) );
XOR2_X1 U1022 ( .A(n1361), .B(n1362), .Z(n1360) );
XOR2_X1 U1023 ( .A(KEYINPUT41), .B(n1254), .Z(n1362) );
XOR2_X1 U1024 ( .A(n1250), .B(n1251), .Z(n1361) );
AND2_X1 U1025 ( .A1(n1363), .A2(n1364), .ZN(n1251) );
NAND2_X1 U1026 ( .A1(n1365), .A2(n1326), .ZN(n1364) );
NAND2_X1 U1027 ( .A1(n1366), .A2(G210), .ZN(n1365) );
NAND3_X1 U1028 ( .A1(n1366), .A2(G210), .A3(G101), .ZN(n1363) );
NAND2_X1 U1029 ( .A1(n1367), .A2(n1368), .ZN(n1250) );
NAND2_X1 U1030 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
INV_X1 U1031 ( .A(G113), .ZN(n1370) );
XOR2_X1 U1032 ( .A(n1371), .B(KEYINPUT58), .Z(n1369) );
NAND2_X1 U1033 ( .A1(n1372), .A2(G113), .ZN(n1367) );
XOR2_X1 U1034 ( .A(KEYINPUT32), .B(n1373), .Z(n1372) );
INV_X1 U1035 ( .A(n1371), .ZN(n1373) );
XOR2_X1 U1036 ( .A(n1374), .B(n1375), .Z(n1371) );
XOR2_X1 U1037 ( .A(n1376), .B(G119), .Z(n1374) );
INV_X1 U1038 ( .A(G116), .ZN(n1376) );
AND3_X1 U1039 ( .A1(n1139), .A2(n1294), .A3(n1147), .ZN(n1292) );
NOR2_X1 U1040 ( .A1(n1327), .A2(n1123), .ZN(n1147) );
INV_X1 U1041 ( .A(n1148), .ZN(n1123) );
NAND2_X1 U1042 ( .A1(G221), .A2(n1342), .ZN(n1148) );
NAND2_X1 U1043 ( .A1(G234), .A2(n1343), .ZN(n1342) );
INV_X1 U1044 ( .A(n1122), .ZN(n1327) );
XOR2_X1 U1045 ( .A(n1160), .B(n1377), .Z(n1122) );
NOR2_X1 U1046 ( .A1(n1378), .A2(KEYINPUT35), .ZN(n1377) );
INV_X1 U1047 ( .A(n1161), .ZN(n1378) );
NAND2_X1 U1048 ( .A1(n1379), .A2(n1343), .ZN(n1161) );
XOR2_X1 U1049 ( .A(n1380), .B(n1381), .Z(n1379) );
XOR2_X1 U1050 ( .A(n1382), .B(n1262), .Z(n1381) );
NAND2_X1 U1051 ( .A1(G227), .A2(n1149), .ZN(n1262) );
NAND2_X1 U1052 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
NAND2_X1 U1053 ( .A1(n1385), .A2(n1254), .ZN(n1384) );
XOR2_X1 U1054 ( .A(KEYINPUT26), .B(n1386), .Z(n1383) );
NOR2_X1 U1055 ( .A1(n1385), .A2(n1254), .ZN(n1386) );
XNOR2_X1 U1056 ( .A(n1387), .B(n1388), .ZN(n1254) );
XOR2_X1 U1057 ( .A(G131), .B(n1389), .Z(n1388) );
NOR2_X1 U1058 ( .A1(G134), .A2(KEYINPUT31), .ZN(n1389) );
XOR2_X1 U1059 ( .A(n1202), .B(KEYINPUT37), .Z(n1387) );
INV_X1 U1060 ( .A(G137), .ZN(n1202) );
XNOR2_X1 U1061 ( .A(n1390), .B(n1274), .ZN(n1385) );
AND2_X1 U1062 ( .A1(n1391), .A2(n1392), .ZN(n1274) );
NAND2_X1 U1063 ( .A1(G101), .A2(n1393), .ZN(n1392) );
XOR2_X1 U1064 ( .A(KEYINPUT54), .B(n1394), .Z(n1391) );
NOR2_X1 U1065 ( .A1(n1395), .A2(n1393), .ZN(n1394) );
XOR2_X1 U1066 ( .A(G104), .B(n1396), .Z(n1393) );
XOR2_X1 U1067 ( .A(KEYINPUT15), .B(G107), .Z(n1396) );
XOR2_X1 U1068 ( .A(n1326), .B(KEYINPUT1), .Z(n1395) );
INV_X1 U1069 ( .A(G101), .ZN(n1326) );
NAND2_X1 U1070 ( .A1(KEYINPUT62), .A2(n1397), .ZN(n1390) );
INV_X1 U1071 ( .A(n1195), .ZN(n1397) );
XOR2_X1 U1072 ( .A(n1398), .B(n1399), .Z(n1195) );
XOR2_X1 U1073 ( .A(KEYINPUT53), .B(KEYINPUT3), .Z(n1399) );
XOR2_X1 U1074 ( .A(n1314), .B(n1400), .Z(n1398) );
XOR2_X1 U1075 ( .A(G110), .B(n1401), .Z(n1380) );
XOR2_X1 U1076 ( .A(KEYINPUT59), .B(G140), .Z(n1401) );
INV_X1 U1077 ( .A(G469), .ZN(n1160) );
NAND2_X1 U1078 ( .A1(n1119), .A2(n1402), .ZN(n1294) );
NAND3_X1 U1079 ( .A1(n1210), .A2(n1330), .A3(G902), .ZN(n1402) );
NOR2_X1 U1080 ( .A1(G898), .A2(n1149), .ZN(n1210) );
NAND3_X1 U1081 ( .A1(n1330), .A2(n1149), .A3(G952), .ZN(n1119) );
NAND2_X1 U1082 ( .A1(G237), .A2(G234), .ZN(n1330) );
INV_X1 U1083 ( .A(n1244), .ZN(n1139) );
NAND2_X1 U1084 ( .A1(n1152), .A2(n1140), .ZN(n1244) );
NAND3_X1 U1085 ( .A1(n1403), .A2(n1404), .A3(n1405), .ZN(n1140) );
INV_X1 U1086 ( .A(n1167), .ZN(n1405) );
NOR2_X1 U1087 ( .A1(n1169), .A2(n1168), .ZN(n1167) );
OR2_X1 U1088 ( .A1(n1168), .A2(KEYINPUT49), .ZN(n1404) );
NAND3_X1 U1089 ( .A1(n1168), .A2(n1169), .A3(KEYINPUT49), .ZN(n1403) );
NAND2_X1 U1090 ( .A1(n1406), .A2(n1343), .ZN(n1169) );
XOR2_X1 U1091 ( .A(n1312), .B(n1407), .Z(n1406) );
INV_X1 U1092 ( .A(n1313), .ZN(n1407) );
XOR2_X1 U1093 ( .A(n1408), .B(n1375), .Z(n1313) );
XOR2_X1 U1094 ( .A(n1400), .B(n1409), .Z(n1375) );
NOR2_X1 U1095 ( .A1(G146), .A2(KEYINPUT60), .ZN(n1409) );
XOR2_X1 U1096 ( .A(G128), .B(G143), .Z(n1400) );
XOR2_X1 U1097 ( .A(n1192), .B(n1410), .Z(n1408) );
NOR2_X1 U1098 ( .A1(G953), .A2(n1212), .ZN(n1410) );
INV_X1 U1099 ( .A(G224), .ZN(n1212) );
NAND2_X1 U1100 ( .A1(n1411), .A2(n1412), .ZN(n1312) );
NAND2_X1 U1101 ( .A1(n1413), .A2(n1414), .ZN(n1412) );
INV_X1 U1102 ( .A(KEYINPUT38), .ZN(n1414) );
NAND2_X1 U1103 ( .A1(n1415), .A2(n1416), .ZN(n1413) );
NAND2_X1 U1104 ( .A1(n1221), .A2(n1222), .ZN(n1416) );
INV_X1 U1105 ( .A(n1218), .ZN(n1415) );
NOR2_X1 U1106 ( .A1(n1222), .A2(n1221), .ZN(n1218) );
NAND2_X1 U1107 ( .A1(KEYINPUT38), .A2(n1417), .ZN(n1411) );
XOR2_X1 U1108 ( .A(n1222), .B(n1221), .Z(n1417) );
XOR2_X1 U1109 ( .A(n1276), .B(G122), .Z(n1221) );
XNOR2_X1 U1110 ( .A(n1418), .B(n1419), .ZN(n1222) );
XOR2_X1 U1111 ( .A(n1420), .B(n1421), .Z(n1419) );
NOR2_X1 U1112 ( .A1(G116), .A2(KEYINPUT21), .ZN(n1420) );
XOR2_X1 U1113 ( .A(n1422), .B(n1423), .Z(n1418) );
XOR2_X1 U1114 ( .A(G119), .B(G101), .Z(n1423) );
NAND2_X1 U1115 ( .A1(KEYINPUT23), .A2(n1424), .ZN(n1422) );
INV_X1 U1116 ( .A(n1281), .ZN(n1168) );
NAND2_X1 U1117 ( .A1(G210), .A2(n1425), .ZN(n1281) );
NAND2_X1 U1118 ( .A1(G214), .A2(n1425), .ZN(n1152) );
NAND2_X1 U1119 ( .A1(n1426), .A2(n1343), .ZN(n1425) );
INV_X1 U1120 ( .A(G237), .ZN(n1426) );
INV_X1 U1121 ( .A(n1132), .ZN(n1319) );
NAND2_X1 U1122 ( .A1(n1336), .A2(n1162), .ZN(n1132) );
XOR2_X1 U1123 ( .A(n1427), .B(G475), .Z(n1162) );
NAND2_X1 U1124 ( .A1(n1239), .A2(n1343), .ZN(n1427) );
XOR2_X1 U1125 ( .A(n1428), .B(n1429), .Z(n1239) );
XNOR2_X1 U1126 ( .A(n1430), .B(n1421), .ZN(n1429) );
XOR2_X1 U1127 ( .A(G104), .B(G113), .Z(n1421) );
NAND3_X1 U1128 ( .A1(n1431), .A2(n1432), .A3(n1433), .ZN(n1430) );
NAND2_X1 U1129 ( .A1(n1434), .A2(n1435), .ZN(n1433) );
NAND2_X1 U1130 ( .A1(KEYINPUT55), .A2(n1436), .ZN(n1435) );
XOR2_X1 U1131 ( .A(KEYINPUT10), .B(G131), .Z(n1436) );
NAND3_X1 U1132 ( .A1(KEYINPUT55), .A2(n1437), .A3(n1321), .ZN(n1432) );
INV_X1 U1133 ( .A(n1434), .ZN(n1437) );
XOR2_X1 U1134 ( .A(n1438), .B(G143), .Z(n1434) );
NAND2_X1 U1135 ( .A1(n1366), .A2(G214), .ZN(n1438) );
NOR2_X1 U1136 ( .A1(G953), .A2(G237), .ZN(n1366) );
OR2_X1 U1137 ( .A1(n1321), .A2(KEYINPUT55), .ZN(n1431) );
INV_X1 U1138 ( .A(G131), .ZN(n1321) );
XOR2_X1 U1139 ( .A(n1439), .B(G122), .Z(n1428) );
NAND3_X1 U1140 ( .A1(n1440), .A2(n1441), .A3(n1442), .ZN(n1439) );
NAND2_X1 U1141 ( .A1(G146), .A2(n1443), .ZN(n1442) );
NAND2_X1 U1142 ( .A1(KEYINPUT33), .A2(n1444), .ZN(n1441) );
NAND2_X1 U1143 ( .A1(n1445), .A2(n1314), .ZN(n1444) );
INV_X1 U1144 ( .A(G146), .ZN(n1314) );
XNOR2_X1 U1145 ( .A(KEYINPUT43), .B(n1443), .ZN(n1445) );
NAND2_X1 U1146 ( .A1(n1446), .A2(n1447), .ZN(n1440) );
INV_X1 U1147 ( .A(KEYINPUT33), .ZN(n1447) );
NAND2_X1 U1148 ( .A1(n1448), .A2(n1449), .ZN(n1446) );
OR3_X1 U1149 ( .A1(n1443), .A2(G146), .A3(KEYINPUT43), .ZN(n1449) );
NAND2_X1 U1150 ( .A1(KEYINPUT43), .A2(n1443), .ZN(n1448) );
XOR2_X1 U1151 ( .A(n1192), .B(n1183), .Z(n1443) );
INV_X1 U1152 ( .A(G140), .ZN(n1183) );
INV_X1 U1153 ( .A(G125), .ZN(n1192) );
NOR2_X1 U1154 ( .A1(n1166), .A2(n1450), .ZN(n1336) );
AND2_X1 U1155 ( .A1(n1451), .A2(n1452), .ZN(n1450) );
XOR2_X1 U1156 ( .A(n1159), .B(KEYINPUT22), .Z(n1452) );
XOR2_X1 U1157 ( .A(n1237), .B(KEYINPUT42), .Z(n1451) );
INV_X1 U1158 ( .A(G478), .ZN(n1237) );
NOR2_X1 U1159 ( .A1(n1159), .A2(G478), .ZN(n1166) );
NAND2_X1 U1160 ( .A1(n1343), .A2(n1235), .ZN(n1159) );
NAND2_X1 U1161 ( .A1(n1453), .A2(n1454), .ZN(n1235) );
NAND4_X1 U1162 ( .A1(n1455), .A2(G217), .A3(n1456), .A4(G234), .ZN(n1454) );
NOR2_X1 U1163 ( .A1(G953), .A2(n1457), .ZN(n1456) );
NAND2_X1 U1164 ( .A1(n1458), .A2(n1459), .ZN(n1453) );
NAND3_X1 U1165 ( .A1(G234), .A2(n1149), .A3(G217), .ZN(n1459) );
INV_X1 U1166 ( .A(G953), .ZN(n1149) );
NAND2_X1 U1167 ( .A1(n1455), .A2(n1460), .ZN(n1458) );
INV_X1 U1168 ( .A(n1457), .ZN(n1460) );
NOR2_X1 U1169 ( .A1(n1461), .A2(n1462), .ZN(n1457) );
XOR2_X1 U1170 ( .A(n1463), .B(KEYINPUT27), .Z(n1455) );
NAND2_X1 U1171 ( .A1(n1462), .A2(n1461), .ZN(n1463) );
XNOR2_X1 U1172 ( .A(n1424), .B(n1464), .ZN(n1461) );
XOR2_X1 U1173 ( .A(G122), .B(G116), .Z(n1464) );
INV_X1 U1174 ( .A(G107), .ZN(n1424) );
XNOR2_X1 U1175 ( .A(n1465), .B(n1466), .ZN(n1462) );
NOR2_X1 U1176 ( .A1(KEYINPUT29), .A2(n1467), .ZN(n1466) );
XOR2_X1 U1177 ( .A(KEYINPUT47), .B(G143), .Z(n1467) );
XOR2_X1 U1178 ( .A(n1323), .B(G134), .Z(n1465) );
INV_X1 U1179 ( .A(G128), .ZN(n1323) );
INV_X1 U1180 ( .A(G902), .ZN(n1343) );
INV_X1 U1181 ( .A(G110), .ZN(n1276) );
endmodule


