//Key = 0111111100000100011111111000010111001010011001100011001001000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368;

XNOR2_X1 U747 ( .A(G107), .B(n1031), .ZN(G9) );
NOR2_X1 U748 ( .A1(n1032), .A2(n1033), .ZN(G75) );
XOR2_X1 U749 ( .A(KEYINPUT34), .B(n1034), .Z(n1033) );
NOR2_X1 U750 ( .A1(G952), .A2(n1035), .ZN(n1034) );
NOR4_X1 U751 ( .A1(n1036), .A2(n1037), .A3(n1035), .A4(n1038), .ZN(n1032) );
NAND2_X1 U752 ( .A1(n1039), .A2(n1040), .ZN(n1035) );
NAND4_X1 U753 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1040) );
NOR4_X1 U754 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1044) );
NOR2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
INV_X1 U756 ( .A(KEYINPUT24), .ZN(n1049) );
NOR2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1047) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1046) );
AND3_X1 U759 ( .A1(KEYINPUT24), .A2(n1055), .A3(n1056), .ZN(n1053) );
INV_X1 U760 ( .A(n1057), .ZN(n1045) );
NOR2_X1 U761 ( .A1(n1058), .A2(n1059), .ZN(n1043) );
XNOR2_X1 U762 ( .A(G472), .B(n1060), .ZN(n1042) );
NOR2_X1 U763 ( .A1(KEYINPUT48), .A2(n1061), .ZN(n1060) );
XNOR2_X1 U764 ( .A(n1062), .B(KEYINPUT37), .ZN(n1041) );
NOR2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(n1036) );
NOR2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR3_X1 U767 ( .A1(n1059), .A2(n1067), .A3(n1068), .ZN(n1066) );
NOR2_X1 U768 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR3_X1 U769 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1070) );
NOR2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U772 ( .A1(n1078), .A2(n1058), .ZN(n1069) );
NOR2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U774 ( .A1(n1081), .A2(n1073), .ZN(n1079) );
NOR4_X1 U775 ( .A1(n1082), .A2(n1073), .A3(n1071), .A4(n1058), .ZN(n1065) );
NOR2_X1 U776 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U777 ( .A1(n1085), .A2(n1068), .ZN(n1084) );
INV_X1 U778 ( .A(n1086), .ZN(n1068) );
NOR2_X1 U779 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR2_X1 U780 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR2_X1 U781 ( .A1(n1091), .A2(n1059), .ZN(n1083) );
NOR2_X1 U782 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
INV_X1 U783 ( .A(n1094), .ZN(n1063) );
XOR2_X1 U784 ( .A(n1095), .B(n1096), .Z(G72) );
XOR2_X1 U785 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U786 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U787 ( .A(G953), .B(KEYINPUT42), .ZN(n1100) );
NOR2_X1 U788 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
XNOR2_X1 U789 ( .A(KEYINPUT30), .B(n1103), .ZN(n1102) );
NOR2_X1 U790 ( .A1(n1104), .A2(n1105), .ZN(n1097) );
XOR2_X1 U791 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U792 ( .A(n1108), .B(n1109), .Z(n1107) );
XNOR2_X1 U793 ( .A(n1110), .B(KEYINPUT27), .ZN(n1109) );
NAND2_X1 U794 ( .A1(KEYINPUT1), .A2(n1111), .ZN(n1110) );
INV_X1 U795 ( .A(G134), .ZN(n1111) );
XOR2_X1 U796 ( .A(n1112), .B(n1113), .Z(n1106) );
NOR2_X1 U797 ( .A1(G900), .A2(n1114), .ZN(n1104) );
XNOR2_X1 U798 ( .A(KEYINPUT54), .B(n1039), .ZN(n1114) );
NOR2_X1 U799 ( .A1(n1115), .A2(n1039), .ZN(n1095) );
NOR2_X1 U800 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U801 ( .A(n1118), .B(n1119), .Z(G69) );
NOR2_X1 U802 ( .A1(n1120), .A2(n1039), .ZN(n1119) );
AND2_X1 U803 ( .A1(G224), .A2(G898), .ZN(n1120) );
NOR2_X1 U804 ( .A1(KEYINPUT11), .A2(n1121), .ZN(n1118) );
XOR2_X1 U805 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U806 ( .A1(n1124), .A2(G953), .ZN(n1123) );
NAND3_X1 U807 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1122) );
XOR2_X1 U808 ( .A(n1128), .B(KEYINPUT16), .Z(n1127) );
NAND2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
OR2_X1 U810 ( .A1(n1130), .A2(n1129), .ZN(n1126) );
NAND2_X1 U811 ( .A1(G953), .A2(n1131), .ZN(n1125) );
NOR2_X1 U812 ( .A1(n1132), .A2(n1133), .ZN(G66) );
XNOR2_X1 U813 ( .A(n1134), .B(n1056), .ZN(n1133) );
NOR2_X1 U814 ( .A1(n1054), .A2(n1135), .ZN(n1134) );
NOR2_X1 U815 ( .A1(n1136), .A2(n1137), .ZN(G63) );
XOR2_X1 U816 ( .A(KEYINPUT14), .B(n1132), .Z(n1137) );
XOR2_X1 U817 ( .A(n1138), .B(n1139), .Z(n1136) );
NAND3_X1 U818 ( .A1(n1140), .A2(G478), .A3(KEYINPUT4), .ZN(n1138) );
NOR2_X1 U819 ( .A1(n1132), .A2(n1141), .ZN(G60) );
XOR2_X1 U820 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U821 ( .A(KEYINPUT56), .B(n1144), .Z(n1143) );
NOR2_X1 U822 ( .A1(n1052), .A2(n1135), .ZN(n1144) );
XOR2_X1 U823 ( .A(G104), .B(n1145), .Z(G6) );
NOR2_X1 U824 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NOR2_X1 U825 ( .A1(KEYINPUT52), .A2(n1148), .ZN(n1147) );
NOR2_X1 U826 ( .A1(KEYINPUT31), .A2(n1149), .ZN(n1146) );
NOR2_X1 U827 ( .A1(n1132), .A2(n1150), .ZN(G57) );
XNOR2_X1 U828 ( .A(n1151), .B(n1152), .ZN(n1150) );
XOR2_X1 U829 ( .A(KEYINPUT49), .B(n1153), .Z(n1152) );
NOR2_X1 U830 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XOR2_X1 U831 ( .A(KEYINPUT44), .B(n1156), .Z(n1155) );
NOR3_X1 U832 ( .A1(n1135), .A2(n1157), .A3(n1158), .ZN(n1156) );
XNOR2_X1 U833 ( .A(n1159), .B(n1160), .ZN(n1158) );
NOR2_X1 U834 ( .A1(n1161), .A2(n1162), .ZN(n1154) );
XOR2_X1 U835 ( .A(n1160), .B(n1159), .Z(n1162) );
NOR2_X1 U836 ( .A1(n1157), .A2(n1135), .ZN(n1161) );
XNOR2_X1 U837 ( .A(KEYINPUT55), .B(G472), .ZN(n1157) );
NOR2_X1 U838 ( .A1(n1132), .A2(n1163), .ZN(G54) );
XOR2_X1 U839 ( .A(n1164), .B(n1165), .Z(n1163) );
XNOR2_X1 U840 ( .A(n1166), .B(n1167), .ZN(n1165) );
AND2_X1 U841 ( .A1(G469), .A2(n1140), .ZN(n1166) );
INV_X1 U842 ( .A(n1135), .ZN(n1140) );
XOR2_X1 U843 ( .A(n1168), .B(n1169), .Z(n1164) );
NOR2_X1 U844 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U845 ( .A(KEYINPUT15), .B(n1172), .Z(n1171) );
AND2_X1 U846 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NOR2_X1 U847 ( .A1(n1174), .A2(n1173), .ZN(n1170) );
XOR2_X1 U848 ( .A(n1175), .B(n1176), .Z(n1173) );
NAND2_X1 U849 ( .A1(KEYINPUT21), .A2(n1177), .ZN(n1175) );
XNOR2_X1 U850 ( .A(KEYINPUT12), .B(n1178), .ZN(n1168) );
NOR2_X1 U851 ( .A1(KEYINPUT58), .A2(n1179), .ZN(n1178) );
INV_X1 U852 ( .A(n1180), .ZN(n1179) );
NOR2_X1 U853 ( .A1(n1132), .A2(n1181), .ZN(G51) );
XOR2_X1 U854 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U855 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U856 ( .A1(n1186), .A2(n1135), .ZN(n1184) );
NAND2_X1 U857 ( .A1(n1187), .A2(n1037), .ZN(n1135) );
NAND3_X1 U858 ( .A1(n1188), .A2(n1103), .A3(n1124), .ZN(n1037) );
AND4_X1 U859 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1124) );
NOR4_X1 U860 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
INV_X1 U861 ( .A(n1031), .ZN(n1195) );
NAND3_X1 U862 ( .A1(n1092), .A2(n1197), .A3(n1088), .ZN(n1031) );
NOR2_X1 U863 ( .A1(n1148), .A2(n1198), .ZN(n1191) );
NOR2_X1 U864 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
INV_X1 U865 ( .A(n1149), .ZN(n1148) );
NAND3_X1 U866 ( .A1(n1088), .A2(n1197), .A3(n1093), .ZN(n1149) );
INV_X1 U867 ( .A(n1101), .ZN(n1188) );
NAND3_X1 U868 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1101) );
AND3_X1 U869 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1203) );
NAND3_X1 U870 ( .A1(n1207), .A2(n1086), .A3(n1208), .ZN(n1202) );
NAND2_X1 U871 ( .A1(n1075), .A2(n1209), .ZN(n1201) );
NAND3_X1 U872 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1209) );
XNOR2_X1 U873 ( .A(n1213), .B(KEYINPUT39), .ZN(n1212) );
XNOR2_X1 U874 ( .A(KEYINPUT0), .B(n1055), .ZN(n1187) );
XNOR2_X1 U875 ( .A(n1214), .B(n1215), .ZN(n1182) );
NOR2_X1 U876 ( .A1(KEYINPUT9), .A2(n1216), .ZN(n1215) );
XNOR2_X1 U877 ( .A(n1217), .B(G125), .ZN(n1216) );
AND2_X1 U878 ( .A1(n1218), .A2(n1038), .ZN(n1132) );
XNOR2_X1 U879 ( .A(KEYINPUT8), .B(n1039), .ZN(n1218) );
XNOR2_X1 U880 ( .A(G146), .B(n1219), .ZN(G48) );
NAND2_X1 U881 ( .A1(n1220), .A2(n1075), .ZN(n1219) );
XOR2_X1 U882 ( .A(n1210), .B(KEYINPUT32), .Z(n1220) );
NAND2_X1 U883 ( .A1(n1221), .A2(n1093), .ZN(n1210) );
NAND3_X1 U884 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(G45) );
NAND3_X1 U885 ( .A1(n1075), .A2(n1225), .A3(n1213), .ZN(n1224) );
NAND2_X1 U886 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
NAND2_X1 U887 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND3_X1 U888 ( .A1(G143), .A2(n1230), .A3(n1226), .ZN(n1223) );
INV_X1 U889 ( .A(KEYINPUT28), .ZN(n1226) );
NAND3_X1 U890 ( .A1(n1075), .A2(n1229), .A3(n1213), .ZN(n1230) );
AND4_X1 U891 ( .A1(n1080), .A2(n1231), .A3(n1232), .A4(n1088), .ZN(n1213) );
NOR2_X1 U892 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
INV_X1 U893 ( .A(n1062), .ZN(n1234) );
INV_X1 U894 ( .A(KEYINPUT59), .ZN(n1229) );
NAND2_X1 U895 ( .A1(KEYINPUT28), .A2(n1228), .ZN(n1222) );
NAND2_X1 U896 ( .A1(n1235), .A2(n1236), .ZN(G42) );
NAND2_X1 U897 ( .A1(n1237), .A2(n1204), .ZN(n1236) );
NAND2_X1 U898 ( .A1(n1176), .A2(n1238), .ZN(n1237) );
NAND2_X1 U899 ( .A1(KEYINPUT17), .A2(n1239), .ZN(n1238) );
INV_X1 U900 ( .A(KEYINPUT33), .ZN(n1239) );
NAND3_X1 U901 ( .A1(n1240), .A2(n1241), .A3(KEYINPUT33), .ZN(n1235) );
OR2_X1 U902 ( .A1(G140), .A2(KEYINPUT17), .ZN(n1241) );
NAND2_X1 U903 ( .A1(KEYINPUT17), .A2(n1242), .ZN(n1240) );
OR2_X1 U904 ( .A1(n1204), .A2(G140), .ZN(n1242) );
NAND2_X1 U905 ( .A1(n1243), .A2(n1207), .ZN(n1204) );
XNOR2_X1 U906 ( .A(G137), .B(n1244), .ZN(G39) );
NAND3_X1 U907 ( .A1(n1208), .A2(n1207), .A3(n1245), .ZN(n1244) );
XNOR2_X1 U908 ( .A(KEYINPUT45), .B(n1086), .ZN(n1245) );
XNOR2_X1 U909 ( .A(G134), .B(n1103), .ZN(G36) );
NAND3_X1 U910 ( .A1(n1207), .A2(n1092), .A3(n1080), .ZN(n1103) );
XNOR2_X1 U911 ( .A(G131), .B(n1205), .ZN(G33) );
NAND3_X1 U912 ( .A1(n1080), .A2(n1207), .A3(n1093), .ZN(n1205) );
AND3_X1 U913 ( .A1(n1246), .A2(n1088), .A3(n1231), .ZN(n1207) );
INV_X1 U914 ( .A(n1058), .ZN(n1246) );
NAND2_X1 U915 ( .A1(n1247), .A2(n1077), .ZN(n1058) );
INV_X1 U916 ( .A(n1076), .ZN(n1247) );
XNOR2_X1 U917 ( .A(G128), .B(n1248), .ZN(G30) );
NAND2_X1 U918 ( .A1(n1249), .A2(n1075), .ZN(n1248) );
XOR2_X1 U919 ( .A(n1211), .B(KEYINPUT51), .Z(n1249) );
NAND2_X1 U920 ( .A1(n1221), .A2(n1092), .ZN(n1211) );
AND3_X1 U921 ( .A1(n1231), .A2(n1088), .A3(n1208), .ZN(n1221) );
XOR2_X1 U922 ( .A(G101), .B(n1250), .Z(G3) );
NOR3_X1 U923 ( .A1(n1200), .A2(KEYINPUT62), .A3(n1199), .ZN(n1250) );
INV_X1 U924 ( .A(n1080), .ZN(n1199) );
XNOR2_X1 U925 ( .A(G125), .B(n1206), .ZN(G27) );
NAND4_X1 U926 ( .A1(n1243), .A2(n1231), .A3(n1251), .A4(n1075), .ZN(n1206) );
AND3_X1 U927 ( .A1(n1252), .A2(n1253), .A3(n1094), .ZN(n1231) );
NAND2_X1 U928 ( .A1(G953), .A2(n1254), .ZN(n1252) );
NAND2_X1 U929 ( .A1(G902), .A2(n1117), .ZN(n1254) );
INV_X1 U930 ( .A(G900), .ZN(n1117) );
AND3_X1 U931 ( .A1(n1255), .A2(n1071), .A3(n1093), .ZN(n1243) );
XNOR2_X1 U932 ( .A(G122), .B(n1189), .ZN(G24) );
NAND4_X1 U933 ( .A1(n1251), .A2(n1197), .A3(n1062), .A4(n1256), .ZN(n1189) );
AND3_X1 U934 ( .A1(n1257), .A2(n1255), .A3(n1081), .ZN(n1197) );
XNOR2_X1 U935 ( .A(G119), .B(n1190), .ZN(G21) );
NAND4_X1 U936 ( .A1(n1208), .A2(n1251), .A3(n1257), .A4(n1086), .ZN(n1190) );
AND2_X1 U937 ( .A1(n1258), .A2(n1071), .ZN(n1208) );
XNOR2_X1 U938 ( .A(KEYINPUT38), .B(n1073), .ZN(n1258) );
XNOR2_X1 U939 ( .A(n1259), .B(n1196), .ZN(G18) );
AND4_X1 U940 ( .A1(n1080), .A2(n1251), .A3(n1092), .A4(n1257), .ZN(n1196) );
AND2_X1 U941 ( .A1(n1260), .A2(n1062), .ZN(n1092) );
XNOR2_X1 U942 ( .A(KEYINPUT40), .B(n1256), .ZN(n1260) );
NAND2_X1 U943 ( .A1(n1261), .A2(n1262), .ZN(G15) );
OR2_X1 U944 ( .A1(n1263), .A2(G113), .ZN(n1262) );
NAND2_X1 U945 ( .A1(G113), .A2(n1264), .ZN(n1261) );
NAND2_X1 U946 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NAND2_X1 U947 ( .A1(n1194), .A2(n1267), .ZN(n1266) );
INV_X1 U948 ( .A(KEYINPUT3), .ZN(n1267) );
NAND2_X1 U949 ( .A1(KEYINPUT3), .A2(n1263), .ZN(n1265) );
NAND2_X1 U950 ( .A1(KEYINPUT63), .A2(n1194), .ZN(n1263) );
AND4_X1 U951 ( .A1(n1093), .A2(n1080), .A3(n1251), .A4(n1257), .ZN(n1194) );
INV_X1 U952 ( .A(n1059), .ZN(n1251) );
NAND2_X1 U953 ( .A1(n1268), .A2(n1090), .ZN(n1059) );
INV_X1 U954 ( .A(n1089), .ZN(n1268) );
NOR2_X1 U955 ( .A1(n1255), .A2(n1071), .ZN(n1080) );
XNOR2_X1 U956 ( .A(n1177), .B(n1193), .ZN(G12) );
NOR3_X1 U957 ( .A1(n1073), .A2(n1081), .A3(n1200), .ZN(n1193) );
NAND3_X1 U958 ( .A1(n1257), .A2(n1086), .A3(n1088), .ZN(n1200) );
AND2_X1 U959 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U960 ( .A1(G221), .A2(n1269), .ZN(n1090) );
XNOR2_X1 U961 ( .A(n1270), .B(G469), .ZN(n1089) );
NAND2_X1 U962 ( .A1(n1271), .A2(n1055), .ZN(n1270) );
XOR2_X1 U963 ( .A(n1272), .B(n1273), .Z(n1271) );
XNOR2_X1 U964 ( .A(n1177), .B(n1174), .ZN(n1273) );
NOR2_X1 U965 ( .A1(n1116), .A2(G953), .ZN(n1174) );
INV_X1 U966 ( .A(G227), .ZN(n1116) );
XNOR2_X1 U967 ( .A(n1274), .B(n1275), .ZN(n1272) );
NAND2_X1 U968 ( .A1(KEYINPUT50), .A2(n1176), .ZN(n1275) );
NAND3_X1 U969 ( .A1(n1276), .A2(n1277), .A3(KEYINPUT57), .ZN(n1274) );
NAND2_X1 U970 ( .A1(n1167), .A2(n1180), .ZN(n1277) );
XOR2_X1 U971 ( .A(KEYINPUT22), .B(n1278), .Z(n1276) );
NOR2_X1 U972 ( .A1(n1167), .A2(n1180), .ZN(n1278) );
XNOR2_X1 U973 ( .A(n1112), .B(n1279), .ZN(n1180) );
XOR2_X1 U974 ( .A(G104), .B(n1280), .Z(n1279) );
NAND2_X1 U975 ( .A1(n1281), .A2(n1282), .ZN(n1112) );
NAND2_X1 U976 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
INV_X1 U977 ( .A(G146), .ZN(n1284) );
XOR2_X1 U978 ( .A(KEYINPUT7), .B(n1285), .Z(n1283) );
NAND2_X1 U979 ( .A1(n1285), .A2(G146), .ZN(n1281) );
NAND2_X1 U980 ( .A1(n1286), .A2(n1287), .ZN(n1086) );
OR3_X1 U981 ( .A1(n1256), .A2(n1062), .A3(KEYINPUT40), .ZN(n1287) );
NAND2_X1 U982 ( .A1(KEYINPUT40), .A2(n1093), .ZN(n1286) );
NOR2_X1 U983 ( .A1(n1062), .A2(n1233), .ZN(n1093) );
INV_X1 U984 ( .A(n1256), .ZN(n1233) );
NAND3_X1 U985 ( .A1(n1288), .A2(n1289), .A3(n1057), .ZN(n1256) );
NAND2_X1 U986 ( .A1(n1051), .A2(n1052), .ZN(n1057) );
OR3_X1 U987 ( .A1(n1052), .A2(n1051), .A3(KEYINPUT25), .ZN(n1289) );
NOR2_X1 U988 ( .A1(n1142), .A2(G902), .ZN(n1051) );
XOR2_X1 U989 ( .A(n1290), .B(n1291), .Z(n1142) );
XOR2_X1 U990 ( .A(n1292), .B(n1293), .Z(n1291) );
XNOR2_X1 U991 ( .A(G131), .B(G122), .ZN(n1293) );
NAND2_X1 U992 ( .A1(G214), .A2(n1294), .ZN(n1292) );
XNOR2_X1 U993 ( .A(n1113), .B(n1295), .ZN(n1290) );
XOR2_X1 U994 ( .A(n1296), .B(n1297), .Z(n1295) );
NAND2_X1 U995 ( .A1(KEYINPUT25), .A2(n1052), .ZN(n1288) );
INV_X1 U996 ( .A(G475), .ZN(n1052) );
XNOR2_X1 U997 ( .A(n1298), .B(G478), .ZN(n1062) );
NAND2_X1 U998 ( .A1(n1139), .A2(n1055), .ZN(n1298) );
XNOR2_X1 U999 ( .A(n1299), .B(n1300), .ZN(n1139) );
AND2_X1 U1000 ( .A1(n1301), .A2(G217), .ZN(n1300) );
NAND2_X1 U1001 ( .A1(n1302), .A2(n1303), .ZN(n1299) );
NAND2_X1 U1002 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND2_X1 U1003 ( .A1(KEYINPUT19), .A2(n1306), .ZN(n1305) );
NAND2_X1 U1004 ( .A1(KEYINPUT13), .A2(n1307), .ZN(n1306) );
NAND2_X1 U1005 ( .A1(n1308), .A2(n1309), .ZN(n1302) );
NAND2_X1 U1006 ( .A1(KEYINPUT13), .A2(n1310), .ZN(n1309) );
NAND2_X1 U1007 ( .A1(n1311), .A2(KEYINPUT19), .ZN(n1310) );
INV_X1 U1008 ( .A(n1304), .ZN(n1311) );
XOR2_X1 U1009 ( .A(G134), .B(n1285), .Z(n1304) );
XNOR2_X1 U1010 ( .A(n1312), .B(G143), .ZN(n1285) );
INV_X1 U1011 ( .A(n1307), .ZN(n1308) );
XNOR2_X1 U1012 ( .A(n1313), .B(n1314), .ZN(n1307) );
XOR2_X1 U1013 ( .A(KEYINPUT47), .B(G122), .Z(n1314) );
XNOR2_X1 U1014 ( .A(G107), .B(G116), .ZN(n1313) );
AND4_X1 U1015 ( .A1(n1075), .A2(n1094), .A3(n1315), .A4(n1253), .ZN(n1257) );
NAND2_X1 U1016 ( .A1(n1038), .A2(n1039), .ZN(n1253) );
INV_X1 U1017 ( .A(G952), .ZN(n1038) );
NAND2_X1 U1018 ( .A1(G953), .A2(n1316), .ZN(n1315) );
NAND2_X1 U1019 ( .A1(G902), .A2(n1131), .ZN(n1316) );
INV_X1 U1020 ( .A(G898), .ZN(n1131) );
NAND2_X1 U1021 ( .A1(G237), .A2(n1317), .ZN(n1094) );
AND2_X1 U1022 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U1023 ( .A1(G214), .A2(n1318), .ZN(n1077) );
XOR2_X1 U1024 ( .A(n1319), .B(n1186), .Z(n1076) );
NAND2_X1 U1025 ( .A1(G210), .A2(n1318), .ZN(n1186) );
NAND2_X1 U1026 ( .A1(n1320), .A2(n1055), .ZN(n1318) );
INV_X1 U1027 ( .A(G237), .ZN(n1320) );
NAND2_X1 U1028 ( .A1(n1321), .A2(n1055), .ZN(n1319) );
XOR2_X1 U1029 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1030 ( .A(n1185), .B(KEYINPUT2), .ZN(n1323) );
XOR2_X1 U1031 ( .A(n1129), .B(n1130), .Z(n1185) );
XNOR2_X1 U1032 ( .A(n1177), .B(n1324), .ZN(n1130) );
XOR2_X1 U1033 ( .A(KEYINPUT6), .B(G122), .Z(n1324) );
XNOR2_X1 U1034 ( .A(n1325), .B(n1326), .ZN(n1129) );
XNOR2_X1 U1035 ( .A(n1259), .B(n1327), .ZN(n1326) );
XNOR2_X1 U1036 ( .A(n1280), .B(n1297), .ZN(n1325) );
XOR2_X1 U1037 ( .A(G104), .B(G113), .Z(n1297) );
XOR2_X1 U1038 ( .A(G101), .B(n1328), .Z(n1280) );
XNOR2_X1 U1039 ( .A(KEYINPUT18), .B(n1329), .ZN(n1328) );
INV_X1 U1040 ( .A(G107), .ZN(n1329) );
NAND2_X1 U1041 ( .A1(n1330), .A2(n1331), .ZN(n1322) );
NAND2_X1 U1042 ( .A1(n1332), .A2(n1214), .ZN(n1331) );
NAND2_X1 U1043 ( .A1(n1333), .A2(n1334), .ZN(n1330) );
INV_X1 U1044 ( .A(n1214), .ZN(n1334) );
NAND2_X1 U1045 ( .A1(G224), .A2(n1039), .ZN(n1214) );
XOR2_X1 U1046 ( .A(KEYINPUT20), .B(n1332), .Z(n1333) );
AND2_X1 U1047 ( .A1(n1335), .A2(n1336), .ZN(n1332) );
NAND2_X1 U1048 ( .A1(n1217), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1049 ( .A(n1338), .B(KEYINPUT26), .Z(n1335) );
NAND2_X1 U1050 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
XNOR2_X1 U1051 ( .A(KEYINPUT60), .B(n1337), .ZN(n1340) );
INV_X1 U1052 ( .A(G125), .ZN(n1337) );
INV_X1 U1053 ( .A(n1071), .ZN(n1081) );
NAND2_X1 U1054 ( .A1(n1341), .A2(n1050), .ZN(n1071) );
NAND3_X1 U1055 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1050) );
NAND2_X1 U1056 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NAND2_X1 U1057 ( .A1(n1056), .A2(n1055), .ZN(n1343) );
XOR2_X1 U1058 ( .A(n1344), .B(n1345), .Z(n1056) );
XOR2_X1 U1059 ( .A(n1346), .B(n1347), .Z(n1345) );
XNOR2_X1 U1060 ( .A(n1348), .B(n1349), .ZN(n1347) );
NAND2_X1 U1061 ( .A1(KEYINPUT46), .A2(n1312), .ZN(n1349) );
INV_X1 U1062 ( .A(G128), .ZN(n1312) );
NAND2_X1 U1063 ( .A1(n1350), .A2(KEYINPUT23), .ZN(n1348) );
XNOR2_X1 U1064 ( .A(G110), .B(KEYINPUT61), .ZN(n1350) );
XNOR2_X1 U1065 ( .A(G137), .B(G146), .ZN(n1346) );
XOR2_X1 U1066 ( .A(n1351), .B(n1113), .Z(n1344) );
XNOR2_X1 U1067 ( .A(G125), .B(n1176), .ZN(n1113) );
INV_X1 U1068 ( .A(G140), .ZN(n1176) );
XNOR2_X1 U1069 ( .A(n1352), .B(n1353), .ZN(n1351) );
NAND2_X1 U1070 ( .A1(n1301), .A2(G221), .ZN(n1352) );
AND2_X1 U1071 ( .A1(G234), .A2(n1039), .ZN(n1301) );
INV_X1 U1072 ( .A(G953), .ZN(n1039) );
INV_X1 U1073 ( .A(n1054), .ZN(n1342) );
NAND2_X1 U1074 ( .A1(G217), .A2(n1269), .ZN(n1054) );
NAND2_X1 U1075 ( .A1(n1317), .A2(n1055), .ZN(n1269) );
XNOR2_X1 U1076 ( .A(G234), .B(KEYINPUT29), .ZN(n1317) );
INV_X1 U1077 ( .A(n1255), .ZN(n1073) );
XOR2_X1 U1078 ( .A(G472), .B(n1354), .Z(n1255) );
NOR2_X1 U1079 ( .A1(n1355), .A2(KEYINPUT53), .ZN(n1354) );
INV_X1 U1080 ( .A(n1061), .ZN(n1355) );
NAND2_X1 U1081 ( .A1(n1356), .A2(n1055), .ZN(n1061) );
INV_X1 U1082 ( .A(G902), .ZN(n1055) );
XNOR2_X1 U1083 ( .A(n1357), .B(n1358), .ZN(n1356) );
XNOR2_X1 U1084 ( .A(n1359), .B(n1160), .ZN(n1358) );
XNOR2_X1 U1085 ( .A(n1360), .B(G113), .ZN(n1160) );
NAND3_X1 U1086 ( .A1(n1361), .A2(n1362), .A3(n1363), .ZN(n1360) );
OR2_X1 U1087 ( .A1(n1259), .A2(n1364), .ZN(n1363) );
NAND3_X1 U1088 ( .A1(n1364), .A2(n1259), .A3(KEYINPUT41), .ZN(n1362) );
INV_X1 U1089 ( .A(G116), .ZN(n1259) );
NOR2_X1 U1090 ( .A1(KEYINPUT35), .A2(n1353), .ZN(n1364) );
INV_X1 U1091 ( .A(n1327), .ZN(n1353) );
OR2_X1 U1092 ( .A1(n1327), .A2(KEYINPUT41), .ZN(n1361) );
XOR2_X1 U1093 ( .A(G119), .B(KEYINPUT5), .Z(n1327) );
NAND2_X1 U1094 ( .A1(KEYINPUT36), .A2(n1159), .ZN(n1359) );
XOR2_X1 U1095 ( .A(n1167), .B(n1339), .Z(n1159) );
INV_X1 U1096 ( .A(n1217), .ZN(n1339) );
XOR2_X1 U1097 ( .A(G128), .B(n1296), .Z(n1217) );
XNOR2_X1 U1098 ( .A(n1228), .B(G146), .ZN(n1296) );
INV_X1 U1099 ( .A(G143), .ZN(n1228) );
XOR2_X1 U1100 ( .A(n1365), .B(n1366), .Z(n1167) );
XOR2_X1 U1101 ( .A(KEYINPUT43), .B(KEYINPUT10), .Z(n1366) );
XNOR2_X1 U1102 ( .A(G134), .B(n1108), .ZN(n1365) );
XNOR2_X1 U1103 ( .A(n1367), .B(G137), .ZN(n1108) );
INV_X1 U1104 ( .A(G131), .ZN(n1367) );
INV_X1 U1105 ( .A(n1151), .ZN(n1357) );
XNOR2_X1 U1106 ( .A(n1368), .B(G101), .ZN(n1151) );
NAND2_X1 U1107 ( .A1(G210), .A2(n1294), .ZN(n1368) );
NOR2_X1 U1108 ( .A1(G953), .A2(G237), .ZN(n1294) );
INV_X1 U1109 ( .A(G110), .ZN(n1177) );
endmodule


