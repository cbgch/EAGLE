//Key = 1111000011101100101001011011100010101011001001111101010000000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256;

XOR2_X1 U693 ( .A(G107), .B(n958), .Z(G9) );
NOR2_X1 U694 ( .A1(n959), .A2(n960), .ZN(G75) );
NOR3_X1 U695 ( .A1(n961), .A2(n962), .A3(n963), .ZN(n960) );
XOR2_X1 U696 ( .A(KEYINPUT63), .B(n964), .Z(n963) );
NAND3_X1 U697 ( .A1(n965), .A2(n966), .A3(n967), .ZN(n961) );
NAND2_X1 U698 ( .A1(n968), .A2(n969), .ZN(n967) );
NAND2_X1 U699 ( .A1(n970), .A2(n971), .ZN(n968) );
NAND3_X1 U700 ( .A1(n972), .A2(n973), .A3(n974), .ZN(n971) );
NAND2_X1 U701 ( .A1(n975), .A2(n976), .ZN(n973) );
NAND2_X1 U702 ( .A1(n977), .A2(n978), .ZN(n976) );
NAND2_X1 U703 ( .A1(n979), .A2(n980), .ZN(n978) );
NAND2_X1 U704 ( .A1(n981), .A2(n982), .ZN(n975) );
NAND2_X1 U705 ( .A1(n983), .A2(n984), .ZN(n982) );
NAND2_X1 U706 ( .A1(n985), .A2(n986), .ZN(n984) );
NAND3_X1 U707 ( .A1(n977), .A2(n987), .A3(n981), .ZN(n970) );
NAND2_X1 U708 ( .A1(n988), .A2(n989), .ZN(n987) );
NAND2_X1 U709 ( .A1(n974), .A2(n990), .ZN(n989) );
NAND2_X1 U710 ( .A1(n991), .A2(n992), .ZN(n990) );
NAND2_X1 U711 ( .A1(n972), .A2(n993), .ZN(n988) );
NAND2_X1 U712 ( .A1(n994), .A2(n995), .ZN(n993) );
NAND2_X1 U713 ( .A1(n996), .A2(n997), .ZN(n995) );
AND3_X1 U714 ( .A1(n965), .A2(n966), .A3(n998), .ZN(n959) );
NAND4_X1 U715 ( .A1(n996), .A2(n977), .A3(n999), .A4(n1000), .ZN(n965) );
NOR4_X1 U716 ( .A1(n997), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(n1000) );
XOR2_X1 U717 ( .A(n1004), .B(n1005), .Z(n1002) );
NAND2_X1 U718 ( .A1(KEYINPUT47), .A2(n1006), .ZN(n1004) );
XOR2_X1 U719 ( .A(n1007), .B(n1008), .Z(n1001) );
NOR2_X1 U720 ( .A1(n1009), .A2(KEYINPUT5), .ZN(n1008) );
XNOR2_X1 U721 ( .A(n1010), .B(n1011), .ZN(n999) );
XOR2_X1 U722 ( .A(n1012), .B(n1013), .Z(G72) );
XOR2_X1 U723 ( .A(n1014), .B(n1015), .Z(n1013) );
NOR2_X1 U724 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
XOR2_X1 U725 ( .A(n1018), .B(n1019), .Z(n1017) );
XOR2_X1 U726 ( .A(n1020), .B(n1021), .Z(n1019) );
XNOR2_X1 U727 ( .A(G143), .B(n1022), .ZN(n1021) );
NOR2_X1 U728 ( .A1(G131), .A2(KEYINPUT22), .ZN(n1022) );
XOR2_X1 U729 ( .A(n1023), .B(n1024), .Z(n1018) );
NOR2_X1 U730 ( .A1(G900), .A2(n966), .ZN(n1016) );
NAND2_X1 U731 ( .A1(n966), .A2(n962), .ZN(n1014) );
NAND2_X1 U732 ( .A1(G953), .A2(n1025), .ZN(n1012) );
NAND2_X1 U733 ( .A1(G900), .A2(G227), .ZN(n1025) );
XOR2_X1 U734 ( .A(n1026), .B(n1027), .Z(G69) );
XOR2_X1 U735 ( .A(n1028), .B(n1029), .Z(n1027) );
NOR2_X1 U736 ( .A1(n964), .A2(n1030), .ZN(n1029) );
XNOR2_X1 U737 ( .A(G953), .B(KEYINPUT0), .ZN(n1030) );
NAND2_X1 U738 ( .A1(G953), .A2(n1031), .ZN(n1028) );
NAND2_X1 U739 ( .A1(G898), .A2(G224), .ZN(n1031) );
NAND2_X1 U740 ( .A1(n1032), .A2(n1033), .ZN(n1026) );
NAND2_X1 U741 ( .A1(G953), .A2(n1034), .ZN(n1033) );
NOR2_X1 U742 ( .A1(n1035), .A2(n1036), .ZN(G66) );
XOR2_X1 U743 ( .A(n1037), .B(n1038), .Z(n1036) );
NOR2_X1 U744 ( .A1(KEYINPUT6), .A2(n1039), .ZN(n1038) );
XOR2_X1 U745 ( .A(n1040), .B(n1041), .Z(n1039) );
NAND2_X1 U746 ( .A1(n1042), .A2(n1009), .ZN(n1037) );
NOR2_X1 U747 ( .A1(n1035), .A2(n1043), .ZN(G63) );
XOR2_X1 U748 ( .A(n1044), .B(n1045), .Z(n1043) );
NAND3_X1 U749 ( .A1(G478), .A2(n1042), .A3(KEYINPUT53), .ZN(n1044) );
NOR2_X1 U750 ( .A1(n1035), .A2(n1046), .ZN(G60) );
XNOR2_X1 U751 ( .A(n1047), .B(n1048), .ZN(n1046) );
NOR2_X1 U752 ( .A1(n1011), .A2(n1049), .ZN(n1048) );
XNOR2_X1 U753 ( .A(G104), .B(n1050), .ZN(G6) );
NOR2_X1 U754 ( .A1(n1035), .A2(n1051), .ZN(G57) );
XOR2_X1 U755 ( .A(n1052), .B(n1053), .Z(n1051) );
XNOR2_X1 U756 ( .A(n1054), .B(n1055), .ZN(n1053) );
NOR2_X1 U757 ( .A1(KEYINPUT44), .A2(n1056), .ZN(n1055) );
XOR2_X1 U758 ( .A(n1057), .B(n1058), .Z(n1056) );
XOR2_X1 U759 ( .A(n1059), .B(n1060), .Z(n1058) );
NOR2_X1 U760 ( .A1(KEYINPUT31), .A2(n1061), .ZN(n1060) );
AND2_X1 U761 ( .A1(G472), .A2(n1042), .ZN(n1059) );
NOR2_X1 U762 ( .A1(n1035), .A2(n1062), .ZN(G54) );
XOR2_X1 U763 ( .A(n1063), .B(n1064), .Z(n1062) );
XOR2_X1 U764 ( .A(n1065), .B(n1066), .Z(n1064) );
XNOR2_X1 U765 ( .A(n1067), .B(n1068), .ZN(n1063) );
AND2_X1 U766 ( .A1(G469), .A2(n1042), .ZN(n1068) );
INV_X1 U767 ( .A(n1049), .ZN(n1042) );
NOR2_X1 U768 ( .A1(n1035), .A2(n1069), .ZN(G51) );
XOR2_X1 U769 ( .A(n1070), .B(n1071), .Z(n1069) );
NOR2_X1 U770 ( .A1(n1072), .A2(n1049), .ZN(n1071) );
NAND2_X1 U771 ( .A1(G902), .A2(n1073), .ZN(n1049) );
NAND2_X1 U772 ( .A1(n1074), .A2(n964), .ZN(n1073) );
AND4_X1 U773 ( .A1(n1050), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n964) );
NOR4_X1 U774 ( .A1(n1078), .A2(n958), .A3(n1079), .A4(n1080), .ZN(n1077) );
NOR3_X1 U775 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1079) );
XNOR2_X1 U776 ( .A(KEYINPUT48), .B(n991), .ZN(n1081) );
AND3_X1 U777 ( .A1(n972), .A2(n1084), .A3(n1085), .ZN(n958) );
NOR2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1076) );
NAND3_X1 U779 ( .A1(n1085), .A2(n972), .A3(n1088), .ZN(n1050) );
INV_X1 U780 ( .A(n1082), .ZN(n1085) );
INV_X1 U781 ( .A(n962), .ZN(n1074) );
NAND4_X1 U782 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n962) );
AND4_X1 U783 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1092) );
NAND2_X1 U784 ( .A1(n1097), .A2(n974), .ZN(n1091) );
NAND3_X1 U785 ( .A1(n1088), .A2(n1098), .A3(n1099), .ZN(n1090) );
NAND2_X1 U786 ( .A1(n1100), .A2(n1101), .ZN(n1089) );
NAND2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND3_X1 U788 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1070) );
NAND2_X1 U789 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
INV_X1 U790 ( .A(KEYINPUT16), .ZN(n1108) );
NAND3_X1 U791 ( .A1(KEYINPUT16), .A2(n1109), .A3(n1110), .ZN(n1105) );
OR2_X1 U792 ( .A1(n1110), .A2(n1109), .ZN(n1104) );
NOR2_X1 U793 ( .A1(KEYINPUT14), .A2(n1107), .ZN(n1109) );
XOR2_X1 U794 ( .A(n1111), .B(n1112), .Z(n1107) );
XOR2_X1 U795 ( .A(G125), .B(n1113), .Z(n1111) );
INV_X1 U796 ( .A(n1032), .ZN(n1110) );
NOR2_X1 U797 ( .A1(n966), .A2(G952), .ZN(n1035) );
XNOR2_X1 U798 ( .A(G146), .B(n1114), .ZN(G48) );
NAND2_X1 U799 ( .A1(n1115), .A2(n1100), .ZN(n1114) );
XOR2_X1 U800 ( .A(n1103), .B(KEYINPUT3), .Z(n1115) );
NAND3_X1 U801 ( .A1(n1088), .A2(n1116), .A3(n1117), .ZN(n1103) );
XOR2_X1 U802 ( .A(n1118), .B(n1119), .Z(G45) );
XOR2_X1 U803 ( .A(KEYINPUT60), .B(G143), .Z(n1119) );
NOR2_X1 U804 ( .A1(n1120), .A2(n994), .ZN(n1118) );
INV_X1 U805 ( .A(n1100), .ZN(n994) );
XOR2_X1 U806 ( .A(n1102), .B(KEYINPUT19), .Z(n1120) );
NAND4_X1 U807 ( .A1(n1117), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1102) );
XNOR2_X1 U808 ( .A(G140), .B(n1124), .ZN(G42) );
NAND4_X1 U809 ( .A1(KEYINPUT38), .A2(n1099), .A3(n1088), .A4(n1098), .ZN(n1124) );
XNOR2_X1 U810 ( .A(G137), .B(n1096), .ZN(G39) );
NAND3_X1 U811 ( .A1(n1099), .A2(n1116), .A3(n981), .ZN(n1096) );
NAND2_X1 U812 ( .A1(n1125), .A2(n1126), .ZN(G36) );
NAND3_X1 U813 ( .A1(KEYINPUT51), .A2(G134), .A3(n1127), .ZN(n1126) );
NAND2_X1 U814 ( .A1(n1128), .A2(n1129), .ZN(n1125) );
NAND2_X1 U815 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U816 ( .A1(G134), .A2(n1132), .ZN(n1131) );
INV_X1 U817 ( .A(KEYINPUT46), .ZN(n1132) );
NAND2_X1 U818 ( .A1(KEYINPUT46), .A2(n1133), .ZN(n1130) );
NAND2_X1 U819 ( .A1(KEYINPUT51), .A2(G134), .ZN(n1133) );
INV_X1 U820 ( .A(n1127), .ZN(n1128) );
NAND2_X1 U821 ( .A1(n974), .A2(n1134), .ZN(n1127) );
XOR2_X1 U822 ( .A(KEYINPUT41), .B(n1097), .Z(n1134) );
AND3_X1 U823 ( .A1(n1121), .A2(n1084), .A3(n1117), .ZN(n1097) );
INV_X1 U824 ( .A(n980), .ZN(n1084) );
XNOR2_X1 U825 ( .A(G131), .B(n1095), .ZN(G33) );
NAND3_X1 U826 ( .A1(n1121), .A2(n1088), .A3(n1099), .ZN(n1095) );
AND2_X1 U827 ( .A1(n1117), .A2(n974), .ZN(n1099) );
NOR2_X1 U828 ( .A1(n1135), .A2(n1136), .ZN(n974) );
INV_X1 U829 ( .A(n996), .ZN(n1135) );
NOR2_X1 U830 ( .A1(n1137), .A2(n983), .ZN(n1117) );
NAND2_X1 U831 ( .A1(n1138), .A2(n1139), .ZN(G30) );
NAND2_X1 U832 ( .A1(G128), .A2(n1094), .ZN(n1139) );
XOR2_X1 U833 ( .A(n1140), .B(KEYINPUT15), .Z(n1138) );
OR2_X1 U834 ( .A1(n1094), .A2(G128), .ZN(n1140) );
NAND4_X1 U835 ( .A1(n1100), .A2(n1116), .A3(n1141), .A4(n1142), .ZN(n1094) );
NOR2_X1 U836 ( .A1(n980), .A2(n1137), .ZN(n1142) );
XNOR2_X1 U837 ( .A(G101), .B(n1143), .ZN(G3) );
NOR2_X1 U838 ( .A1(n1144), .A2(KEYINPUT25), .ZN(n1143) );
NOR3_X1 U839 ( .A1(n1083), .A2(n1082), .A3(n991), .ZN(n1144) );
XOR2_X1 U840 ( .A(G125), .B(n1145), .Z(G27) );
NOR2_X1 U841 ( .A1(KEYINPUT57), .A2(n1093), .ZN(n1145) );
NAND4_X1 U842 ( .A1(n977), .A2(n1100), .A3(n1098), .A4(n1146), .ZN(n1093) );
NOR2_X1 U843 ( .A1(n1137), .A2(n979), .ZN(n1146) );
NAND3_X1 U844 ( .A1(n1147), .A2(n1148), .A3(n969), .ZN(n1137) );
NAND2_X1 U845 ( .A1(G953), .A2(n1149), .ZN(n1147) );
OR2_X1 U846 ( .A1(n1150), .A2(G900), .ZN(n1149) );
INV_X1 U847 ( .A(n992), .ZN(n1098) );
XOR2_X1 U848 ( .A(G122), .B(n1078), .Z(G24) );
AND4_X1 U849 ( .A1(n977), .A2(n972), .A3(n1151), .A4(n1122), .ZN(n1078) );
NOR2_X1 U850 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NOR2_X1 U851 ( .A1(n1003), .A2(n1154), .ZN(n972) );
XNOR2_X1 U852 ( .A(n1155), .B(n1075), .ZN(G21) );
NAND4_X1 U853 ( .A1(n981), .A2(n977), .A3(n1156), .A4(n1116), .ZN(n1075) );
NAND2_X1 U854 ( .A1(n1157), .A2(n1158), .ZN(n1116) );
OR2_X1 U855 ( .A1(n991), .A2(KEYINPUT10), .ZN(n1158) );
NAND3_X1 U856 ( .A1(n1154), .A2(n1003), .A3(KEYINPUT10), .ZN(n1157) );
XNOR2_X1 U857 ( .A(G119), .B(KEYINPUT24), .ZN(n1155) );
XOR2_X1 U858 ( .A(n1159), .B(n1087), .Z(G18) );
NOR4_X1 U859 ( .A1(n991), .A2(n1160), .A3(n980), .A4(n1152), .ZN(n1087) );
NAND2_X1 U860 ( .A1(n1122), .A2(n1161), .ZN(n980) );
XNOR2_X1 U861 ( .A(KEYINPUT54), .B(n1123), .ZN(n1161) );
XNOR2_X1 U862 ( .A(G116), .B(KEYINPUT49), .ZN(n1159) );
XOR2_X1 U863 ( .A(n1162), .B(G113), .Z(G15) );
NAND2_X1 U864 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NAND2_X1 U865 ( .A1(n1080), .A2(n1165), .ZN(n1164) );
INV_X1 U866 ( .A(KEYINPUT40), .ZN(n1165) );
AND2_X1 U867 ( .A1(n1166), .A2(n977), .ZN(n1080) );
INV_X1 U868 ( .A(n1160), .ZN(n977) );
NAND3_X1 U869 ( .A1(n1166), .A2(n1160), .A3(KEYINPUT40), .ZN(n1163) );
NAND2_X1 U870 ( .A1(n986), .A2(n1167), .ZN(n1160) );
NOR3_X1 U871 ( .A1(n979), .A2(n1152), .A3(n991), .ZN(n1166) );
INV_X1 U872 ( .A(n1121), .ZN(n991) );
NOR2_X1 U873 ( .A1(n1154), .A2(n1168), .ZN(n1121) );
INV_X1 U874 ( .A(n1088), .ZN(n979) );
NOR2_X1 U875 ( .A1(n1153), .A2(n1122), .ZN(n1088) );
XNOR2_X1 U876 ( .A(n1169), .B(n1086), .ZN(G12) );
NOR3_X1 U877 ( .A1(n992), .A2(n1082), .A3(n1083), .ZN(n1086) );
INV_X1 U878 ( .A(n981), .ZN(n1083) );
NOR2_X1 U879 ( .A1(n1123), .A2(n1122), .ZN(n981) );
XOR2_X1 U880 ( .A(n1170), .B(n1005), .Z(n1122) );
AND2_X1 U881 ( .A1(n1045), .A2(n1171), .ZN(n1005) );
XOR2_X1 U882 ( .A(n1172), .B(n1173), .Z(n1045) );
XOR2_X1 U883 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U884 ( .A(n1176), .B(n1177), .Z(n1172) );
AND2_X1 U885 ( .A1(G217), .A2(n1178), .ZN(n1177) );
XOR2_X1 U886 ( .A(n1179), .B(G134), .Z(n1176) );
NAND2_X1 U887 ( .A1(KEYINPUT26), .A2(n1180), .ZN(n1179) );
NAND2_X1 U888 ( .A1(KEYINPUT45), .A2(n1006), .ZN(n1170) );
INV_X1 U889 ( .A(G478), .ZN(n1006) );
INV_X1 U890 ( .A(n1153), .ZN(n1123) );
XOR2_X1 U891 ( .A(n1181), .B(n1010), .Z(n1153) );
NAND2_X1 U892 ( .A1(n1171), .A2(n1047), .ZN(n1010) );
XNOR2_X1 U893 ( .A(n1182), .B(n1183), .ZN(n1047) );
XOR2_X1 U894 ( .A(n1184), .B(n1185), .Z(n1183) );
NAND2_X1 U895 ( .A1(KEYINPUT42), .A2(n1186), .ZN(n1185) );
XOR2_X1 U896 ( .A(n1187), .B(n1188), .Z(n1186) );
XNOR2_X1 U897 ( .A(G131), .B(G143), .ZN(n1188) );
NAND2_X1 U898 ( .A1(n1189), .A2(G214), .ZN(n1187) );
NAND2_X1 U899 ( .A1(n1190), .A2(KEYINPUT61), .ZN(n1184) );
XOR2_X1 U900 ( .A(n1191), .B(n1192), .Z(n1190) );
NAND2_X1 U901 ( .A1(KEYINPUT34), .A2(G122), .ZN(n1191) );
XOR2_X1 U902 ( .A(n1193), .B(n1194), .Z(n1182) );
NOR2_X1 U903 ( .A1(KEYINPUT56), .A2(n1195), .ZN(n1194) );
XOR2_X1 U904 ( .A(n1020), .B(KEYINPUT30), .Z(n1195) );
XNOR2_X1 U905 ( .A(G104), .B(G146), .ZN(n1193) );
NAND2_X1 U906 ( .A1(KEYINPUT23), .A2(n1011), .ZN(n1181) );
INV_X1 U907 ( .A(G475), .ZN(n1011) );
NAND2_X1 U908 ( .A1(n1156), .A2(n1141), .ZN(n1082) );
XOR2_X1 U909 ( .A(n983), .B(KEYINPUT32), .Z(n1141) );
OR2_X1 U910 ( .A1(n986), .A2(n985), .ZN(n983) );
INV_X1 U911 ( .A(n1167), .ZN(n985) );
NAND2_X1 U912 ( .A1(G221), .A2(n1196), .ZN(n1167) );
XOR2_X1 U913 ( .A(n1197), .B(G469), .Z(n986) );
NAND2_X1 U914 ( .A1(n1171), .A2(n1198), .ZN(n1197) );
XNOR2_X1 U915 ( .A(n1199), .B(n1200), .ZN(n1198) );
XNOR2_X1 U916 ( .A(n1201), .B(n1202), .ZN(n1200) );
NOR2_X1 U917 ( .A1(KEYINPUT29), .A2(n1203), .ZN(n1202) );
XOR2_X1 U918 ( .A(n1204), .B(n1065), .Z(n1203) );
XNOR2_X1 U919 ( .A(n1205), .B(G140), .ZN(n1065) );
NAND2_X1 U920 ( .A1(G227), .A2(n1206), .ZN(n1205) );
XNOR2_X1 U921 ( .A(KEYINPUT18), .B(n966), .ZN(n1206) );
XNOR2_X1 U922 ( .A(G110), .B(KEYINPUT11), .ZN(n1204) );
INV_X1 U923 ( .A(G104), .ZN(n1201) );
INV_X1 U924 ( .A(n1067), .ZN(n1199) );
XNOR2_X1 U925 ( .A(n1207), .B(n1208), .ZN(n1067) );
XOR2_X1 U926 ( .A(n1209), .B(n1023), .Z(n1208) );
XOR2_X1 U927 ( .A(n1210), .B(KEYINPUT17), .Z(n1023) );
XNOR2_X1 U928 ( .A(G101), .B(n1175), .ZN(n1207) );
XOR2_X1 U929 ( .A(G107), .B(G143), .Z(n1175) );
INV_X1 U930 ( .A(n1152), .ZN(n1156) );
NAND4_X1 U931 ( .A1(n1100), .A2(n969), .A3(n1211), .A4(n1148), .ZN(n1152) );
NAND2_X1 U932 ( .A1(n998), .A2(n966), .ZN(n1148) );
INV_X1 U933 ( .A(G952), .ZN(n998) );
NAND2_X1 U934 ( .A1(G953), .A2(n1212), .ZN(n1211) );
NAND2_X1 U935 ( .A1(G902), .A2(n1034), .ZN(n1212) );
INV_X1 U936 ( .A(G898), .ZN(n1034) );
NAND2_X1 U937 ( .A1(G237), .A2(n1213), .ZN(n969) );
XOR2_X1 U938 ( .A(KEYINPUT62), .B(G234), .Z(n1213) );
NOR2_X1 U939 ( .A1(n1136), .A2(n996), .ZN(n1100) );
XNOR2_X1 U940 ( .A(n1214), .B(n1072), .ZN(n996) );
NAND2_X1 U941 ( .A1(G210), .A2(n1215), .ZN(n1072) );
NAND2_X1 U942 ( .A1(n1171), .A2(n1216), .ZN(n1214) );
XNOR2_X1 U943 ( .A(n1217), .B(n1032), .ZN(n1216) );
XNOR2_X1 U944 ( .A(n1218), .B(n1219), .ZN(n1032) );
XOR2_X1 U945 ( .A(n1220), .B(n1221), .Z(n1219) );
XNOR2_X1 U946 ( .A(n1222), .B(n1223), .ZN(n1221) );
NAND2_X1 U947 ( .A1(KEYINPUT8), .A2(n1224), .ZN(n1223) );
NAND2_X1 U948 ( .A1(KEYINPUT21), .A2(n1054), .ZN(n1222) );
XNOR2_X1 U949 ( .A(G107), .B(KEYINPUT7), .ZN(n1220) );
XNOR2_X1 U950 ( .A(n1066), .B(n1225), .ZN(n1218) );
XOR2_X1 U951 ( .A(n1174), .B(n1226), .Z(n1225) );
XNOR2_X1 U952 ( .A(n1227), .B(G122), .ZN(n1174) );
INV_X1 U953 ( .A(G116), .ZN(n1227) );
XNOR2_X1 U954 ( .A(G104), .B(n1169), .ZN(n1066) );
NAND2_X1 U955 ( .A1(n1228), .A2(n1229), .ZN(n1217) );
NAND2_X1 U956 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U957 ( .A(n1113), .B(KEYINPUT37), .Z(n1230) );
XOR2_X1 U958 ( .A(KEYINPUT39), .B(n1232), .Z(n1228) );
NOR2_X1 U959 ( .A1(n1231), .A2(n1113), .ZN(n1232) );
NAND2_X1 U960 ( .A1(G224), .A2(n966), .ZN(n1113) );
XNOR2_X1 U961 ( .A(G125), .B(n1233), .ZN(n1231) );
NOR2_X1 U962 ( .A1(KEYINPUT33), .A2(n1112), .ZN(n1233) );
XOR2_X1 U963 ( .A(n997), .B(KEYINPUT50), .Z(n1136) );
AND2_X1 U964 ( .A1(G214), .A2(n1215), .ZN(n997) );
OR2_X1 U965 ( .A1(G902), .A2(G237), .ZN(n1215) );
NAND2_X1 U966 ( .A1(n1168), .A2(n1154), .ZN(n992) );
XNOR2_X1 U967 ( .A(n1007), .B(n1009), .ZN(n1154) );
AND2_X1 U968 ( .A1(G217), .A2(n1196), .ZN(n1009) );
NAND2_X1 U969 ( .A1(G234), .A2(n1150), .ZN(n1196) );
INV_X1 U970 ( .A(G902), .ZN(n1150) );
NAND2_X1 U971 ( .A1(n1234), .A2(n1171), .ZN(n1007) );
XNOR2_X1 U972 ( .A(n1040), .B(n1041), .ZN(n1234) );
NAND2_X1 U973 ( .A1(n1235), .A2(KEYINPUT9), .ZN(n1041) );
XOR2_X1 U974 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U975 ( .A(KEYINPUT12), .B(G137), .Z(n1237) );
NAND2_X1 U976 ( .A1(n1178), .A2(G221), .ZN(n1236) );
AND2_X1 U977 ( .A1(G234), .A2(n966), .ZN(n1178) );
INV_X1 U978 ( .A(G953), .ZN(n966) );
NAND2_X1 U979 ( .A1(n1238), .A2(n1239), .ZN(n1040) );
NAND2_X1 U980 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
XOR2_X1 U981 ( .A(KEYINPUT27), .B(n1242), .Z(n1238) );
NOR2_X1 U982 ( .A1(n1240), .A2(n1243), .ZN(n1242) );
XNOR2_X1 U983 ( .A(n1241), .B(KEYINPUT2), .ZN(n1243) );
XNOR2_X1 U984 ( .A(n1020), .B(n1244), .ZN(n1241) );
NOR2_X1 U985 ( .A1(G146), .A2(KEYINPUT55), .ZN(n1244) );
XNOR2_X1 U986 ( .A(G140), .B(G125), .ZN(n1020) );
XOR2_X1 U987 ( .A(n1180), .B(n1245), .Z(n1240) );
XNOR2_X1 U988 ( .A(n1246), .B(n1247), .ZN(n1245) );
NOR2_X1 U989 ( .A1(KEYINPUT35), .A2(n1248), .ZN(n1247) );
XNOR2_X1 U990 ( .A(G119), .B(KEYINPUT28), .ZN(n1248) );
NAND2_X1 U991 ( .A1(KEYINPUT1), .A2(G110), .ZN(n1246) );
INV_X1 U992 ( .A(n1003), .ZN(n1168) );
XNOR2_X1 U993 ( .A(n1249), .B(G472), .ZN(n1003) );
NAND2_X1 U994 ( .A1(n1171), .A2(n1250), .ZN(n1249) );
XOR2_X1 U995 ( .A(n1251), .B(n1252), .Z(n1250) );
XOR2_X1 U996 ( .A(n1057), .B(n1061), .Z(n1252) );
XOR2_X1 U997 ( .A(n1209), .B(n1112), .Z(n1061) );
XOR2_X1 U998 ( .A(n1210), .B(n1253), .Z(n1112) );
NOR2_X1 U999 ( .A1(G143), .A2(KEYINPUT52), .ZN(n1253) );
XOR2_X1 U1000 ( .A(G146), .B(n1180), .Z(n1210) );
XNOR2_X1 U1001 ( .A(G128), .B(KEYINPUT59), .ZN(n1180) );
XNOR2_X1 U1002 ( .A(G131), .B(n1024), .ZN(n1209) );
XOR2_X1 U1003 ( .A(G137), .B(G134), .Z(n1024) );
XNOR2_X1 U1004 ( .A(n1254), .B(n1224), .ZN(n1057) );
XOR2_X1 U1005 ( .A(n1192), .B(KEYINPUT36), .Z(n1224) );
XOR2_X1 U1006 ( .A(G113), .B(KEYINPUT13), .Z(n1192) );
XNOR2_X1 U1007 ( .A(G116), .B(n1226), .ZN(n1254) );
XOR2_X1 U1008 ( .A(G119), .B(KEYINPUT4), .Z(n1226) );
XOR2_X1 U1009 ( .A(n1255), .B(n1256), .Z(n1251) );
XNOR2_X1 U1010 ( .A(KEYINPUT43), .B(n1054), .ZN(n1256) );
INV_X1 U1011 ( .A(G101), .ZN(n1054) );
NOR2_X1 U1012 ( .A1(n1052), .A2(KEYINPUT58), .ZN(n1255) );
AND2_X1 U1013 ( .A1(n1189), .A2(G210), .ZN(n1052) );
NOR2_X1 U1014 ( .A1(G953), .A2(G237), .ZN(n1189) );
XNOR2_X1 U1015 ( .A(G902), .B(KEYINPUT20), .ZN(n1171) );
INV_X1 U1016 ( .A(G110), .ZN(n1169) );
endmodule


