//Key = 0101010001111111001001111000001100111110111011101110101100100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306;

XOR2_X1 U715 ( .A(n989), .B(n990), .Z(G9) );
NAND2_X1 U716 ( .A1(KEYINPUT31), .A2(G107), .ZN(n990) );
NOR2_X1 U717 ( .A1(n991), .A2(n992), .ZN(G75) );
NOR3_X1 U718 ( .A1(n993), .A2(n994), .A3(n995), .ZN(n992) );
NAND3_X1 U719 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n993) );
NAND2_X1 U720 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND2_X1 U721 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
NAND3_X1 U722 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1002) );
NAND2_X1 U723 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NAND3_X1 U724 ( .A1(n1008), .A2(n1009), .A3(KEYINPUT28), .ZN(n1007) );
NAND2_X1 U725 ( .A1(n1010), .A2(n1011), .ZN(n1006) );
OR2_X1 U726 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND2_X1 U727 ( .A1(n1014), .A2(n1015), .ZN(n1001) );
NAND2_X1 U728 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND3_X1 U729 ( .A1(n1003), .A2(n1018), .A3(n1010), .ZN(n1017) );
NAND2_X1 U730 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND2_X1 U731 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U732 ( .A1(n1005), .A2(n1009), .ZN(n1016) );
NAND4_X1 U733 ( .A1(n1014), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1009) );
NAND2_X1 U734 ( .A1(n1010), .A2(n1026), .ZN(n1025) );
NAND2_X1 U735 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U736 ( .A1(KEYINPUT12), .A2(n1029), .ZN(n1028) );
OR3_X1 U737 ( .A1(n1030), .A2(KEYINPUT12), .A3(n1010), .ZN(n1024) );
NAND2_X1 U738 ( .A1(n1003), .A2(n1031), .ZN(n1023) );
NAND2_X1 U739 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
OR2_X1 U740 ( .A1(n1034), .A2(KEYINPUT28), .ZN(n1033) );
NAND2_X1 U741 ( .A1(n1035), .A2(n1036), .ZN(n1032) );
INV_X1 U742 ( .A(n1037), .ZN(n999) );
AND3_X1 U743 ( .A1(n996), .A2(n997), .A3(n1038), .ZN(n991) );
NAND3_X1 U744 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n996) );
NOR3_X1 U745 ( .A1(n1042), .A2(n1021), .A3(n1035), .ZN(n1041) );
XOR2_X1 U746 ( .A(n1043), .B(n1044), .Z(n1042) );
XOR2_X1 U747 ( .A(KEYINPUT51), .B(KEYINPUT33), .Z(n1044) );
XOR2_X1 U748 ( .A(n1036), .B(KEYINPUT22), .Z(n1043) );
XOR2_X1 U749 ( .A(n1045), .B(n1046), .Z(n1040) );
NAND2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
XOR2_X1 U751 ( .A(KEYINPUT30), .B(n1049), .Z(n1048) );
XNOR2_X1 U752 ( .A(KEYINPUT49), .B(KEYINPUT18), .ZN(n1047) );
XOR2_X1 U753 ( .A(KEYINPUT47), .B(n1050), .Z(n1039) );
AND4_X1 U754 ( .A1(n1051), .A2(n1052), .A3(n1014), .A4(n1053), .ZN(n1050) );
XNOR2_X1 U755 ( .A(KEYINPUT58), .B(n1054), .ZN(n1053) );
NOR2_X1 U756 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
INV_X1 U757 ( .A(n1057), .ZN(n1055) );
XOR2_X1 U758 ( .A(n1058), .B(n1059), .Z(G72) );
XOR2_X1 U759 ( .A(n1060), .B(n1061), .Z(n1059) );
NOR2_X1 U760 ( .A1(n1062), .A2(n997), .ZN(n1061) );
AND2_X1 U761 ( .A1(G227), .A2(G900), .ZN(n1062) );
NAND2_X1 U762 ( .A1(n1063), .A2(n1064), .ZN(n1060) );
NAND2_X1 U763 ( .A1(G953), .A2(n1065), .ZN(n1064) );
XOR2_X1 U764 ( .A(n1066), .B(n1067), .Z(n1063) );
XOR2_X1 U765 ( .A(n1068), .B(n1069), .Z(n1067) );
XOR2_X1 U766 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND2_X1 U767 ( .A1(KEYINPUT55), .A2(n1072), .ZN(n1070) );
INV_X1 U768 ( .A(G134), .ZN(n1072) );
XOR2_X1 U769 ( .A(n1073), .B(n1074), .Z(n1066) );
XOR2_X1 U770 ( .A(n1075), .B(G125), .Z(n1074) );
NAND2_X1 U771 ( .A1(KEYINPUT15), .A2(n1076), .ZN(n1075) );
XNOR2_X1 U772 ( .A(G131), .B(KEYINPUT57), .ZN(n1073) );
NAND2_X1 U773 ( .A1(n997), .A2(n994), .ZN(n1058) );
XOR2_X1 U774 ( .A(n1077), .B(n1078), .Z(G69) );
XOR2_X1 U775 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U776 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U777 ( .A1(G898), .A2(n997), .ZN(n1081) );
NOR2_X1 U778 ( .A1(G953), .A2(n1083), .ZN(n1079) );
XOR2_X1 U779 ( .A(KEYINPUT32), .B(n1084), .Z(n1083) );
NOR2_X1 U780 ( .A1(n1085), .A2(n997), .ZN(n1077) );
AND2_X1 U781 ( .A1(G224), .A2(G898), .ZN(n1085) );
NOR2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(G66) );
XOR2_X1 U783 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U784 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR2_X1 U785 ( .A1(n1086), .A2(n1092), .ZN(G63) );
XOR2_X1 U786 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U787 ( .A1(KEYINPUT6), .A2(n1095), .ZN(n1094) );
XOR2_X1 U788 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U789 ( .A1(n1090), .A2(G478), .ZN(n1093) );
NOR2_X1 U790 ( .A1(n1086), .A2(n1098), .ZN(G60) );
XOR2_X1 U791 ( .A(n1099), .B(n1100), .Z(n1098) );
NAND2_X1 U792 ( .A1(n1090), .A2(G475), .ZN(n1099) );
XOR2_X1 U793 ( .A(n1101), .B(n1102), .Z(G6) );
NAND2_X1 U794 ( .A1(n1012), .A2(n1103), .ZN(n1102) );
NOR2_X1 U795 ( .A1(n1086), .A2(n1104), .ZN(G57) );
XOR2_X1 U796 ( .A(n1105), .B(n1106), .Z(n1104) );
XNOR2_X1 U797 ( .A(n1107), .B(n1108), .ZN(n1106) );
XOR2_X1 U798 ( .A(n1109), .B(n1110), .Z(n1105) );
XOR2_X1 U799 ( .A(n1111), .B(KEYINPUT62), .Z(n1110) );
NAND2_X1 U800 ( .A1(n1090), .A2(G472), .ZN(n1111) );
NAND2_X1 U801 ( .A1(KEYINPUT3), .A2(n1112), .ZN(n1109) );
NOR2_X1 U802 ( .A1(n1086), .A2(n1113), .ZN(G54) );
XOR2_X1 U803 ( .A(n1114), .B(n1115), .Z(n1113) );
XNOR2_X1 U804 ( .A(n1107), .B(n1116), .ZN(n1115) );
XOR2_X1 U805 ( .A(n1117), .B(n1118), .Z(n1114) );
NOR2_X1 U806 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
NOR2_X1 U809 ( .A1(KEYINPUT56), .A2(n1125), .ZN(n1123) );
NOR2_X1 U810 ( .A1(n1126), .A2(n1127), .ZN(n1119) );
NOR2_X1 U811 ( .A1(n1128), .A2(KEYINPUT56), .ZN(n1126) );
NOR2_X1 U812 ( .A1(n1068), .A2(n1124), .ZN(n1128) );
INV_X1 U813 ( .A(KEYINPUT10), .ZN(n1124) );
INV_X1 U814 ( .A(n1122), .ZN(n1068) );
NAND2_X1 U815 ( .A1(n1090), .A2(G469), .ZN(n1117) );
INV_X1 U816 ( .A(n1129), .ZN(n1090) );
NOR2_X1 U817 ( .A1(n1086), .A2(n1130), .ZN(G51) );
XOR2_X1 U818 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U819 ( .A(n1133), .B(n1134), .ZN(n1131) );
NOR2_X1 U820 ( .A1(KEYINPUT0), .A2(n1135), .ZN(n1134) );
NOR3_X1 U821 ( .A1(n1129), .A2(KEYINPUT7), .A3(n1136), .ZN(n1133) );
NAND2_X1 U822 ( .A1(G902), .A2(n1137), .ZN(n1129) );
NAND2_X1 U823 ( .A1(n1084), .A2(n1138), .ZN(n1137) );
XNOR2_X1 U824 ( .A(KEYINPUT20), .B(n994), .ZN(n1138) );
NAND4_X1 U825 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n994) );
AND4_X1 U826 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1142) );
NAND3_X1 U827 ( .A1(n1029), .A2(n1147), .A3(n1012), .ZN(n1141) );
NAND3_X1 U828 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1147) );
NAND2_X1 U829 ( .A1(KEYINPUT38), .A2(n1151), .ZN(n1150) );
NAND2_X1 U830 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
NAND2_X1 U831 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NAND3_X1 U832 ( .A1(n1034), .A2(n1156), .A3(n1005), .ZN(n1155) );
INV_X1 U833 ( .A(KEYINPUT38), .ZN(n1156) );
NAND2_X1 U834 ( .A1(KEYINPUT52), .A2(n1157), .ZN(n1154) );
INV_X1 U835 ( .A(n1158), .ZN(n1157) );
OR3_X1 U836 ( .A1(n1158), .A2(KEYINPUT52), .A3(n1153), .ZN(n1148) );
INV_X1 U837 ( .A(n995), .ZN(n1084) );
NAND4_X1 U838 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n995) );
AND4_X1 U839 ( .A1(n989), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1162) );
NAND2_X1 U840 ( .A1(n1013), .A2(n1103), .ZN(n989) );
AND2_X1 U841 ( .A1(n1166), .A2(n1003), .ZN(n1103) );
NOR3_X1 U842 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1161) );
NOR2_X1 U843 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
INV_X1 U844 ( .A(KEYINPUT5), .ZN(n1170) );
NOR3_X1 U845 ( .A1(KEYINPUT5), .A2(n1172), .A3(n1019), .ZN(n1168) );
AND3_X1 U846 ( .A1(n1173), .A2(n1013), .A3(n1174), .ZN(n1167) );
NAND4_X1 U847 ( .A1(n1012), .A2(n1003), .A3(n1175), .A4(n1176), .ZN(n1159) );
OR2_X1 U848 ( .A1(n1177), .A2(n1166), .ZN(n1176) );
NAND2_X1 U849 ( .A1(n1178), .A2(n1177), .ZN(n1175) );
INV_X1 U850 ( .A(KEYINPUT35), .ZN(n1177) );
NAND3_X1 U851 ( .A1(n1179), .A2(n1008), .A3(n1180), .ZN(n1178) );
AND2_X1 U852 ( .A1(n1181), .A2(n1038), .ZN(n1086) );
INV_X1 U853 ( .A(G952), .ZN(n1038) );
XOR2_X1 U854 ( .A(n997), .B(KEYINPUT45), .Z(n1181) );
XOR2_X1 U855 ( .A(n1182), .B(n1139), .Z(G48) );
NAND3_X1 U856 ( .A1(n1012), .A2(n1183), .A3(n1184), .ZN(n1139) );
XOR2_X1 U857 ( .A(n1140), .B(n1185), .Z(G45) );
NOR2_X1 U858 ( .A1(G143), .A2(KEYINPUT27), .ZN(n1185) );
NAND4_X1 U859 ( .A1(n1184), .A2(n1173), .A3(n1186), .A4(n1187), .ZN(n1140) );
XOR2_X1 U860 ( .A(n1076), .B(n1188), .Z(G42) );
NAND3_X1 U861 ( .A1(n1012), .A2(n1029), .A3(n1151), .ZN(n1188) );
INV_X1 U862 ( .A(G140), .ZN(n1076) );
XNOR2_X1 U863 ( .A(G137), .B(n1189), .ZN(G39) );
NOR2_X1 U864 ( .A1(n1190), .A2(KEYINPUT26), .ZN(n1189) );
INV_X1 U865 ( .A(n1146), .ZN(n1190) );
NAND3_X1 U866 ( .A1(n1183), .A2(n1014), .A3(n1151), .ZN(n1146) );
XOR2_X1 U867 ( .A(n1145), .B(n1191), .Z(G36) );
NAND2_X1 U868 ( .A1(KEYINPUT37), .A2(G134), .ZN(n1191) );
NAND3_X1 U869 ( .A1(n1173), .A2(n1013), .A3(n1151), .ZN(n1145) );
XNOR2_X1 U870 ( .A(G131), .B(n1144), .ZN(G33) );
NAND3_X1 U871 ( .A1(n1012), .A2(n1173), .A3(n1151), .ZN(n1144) );
AND3_X1 U872 ( .A1(n1008), .A2(n1153), .A3(n1005), .ZN(n1151) );
NOR2_X1 U873 ( .A1(n1192), .A2(n1021), .ZN(n1005) );
INV_X1 U874 ( .A(n1022), .ZN(n1192) );
XNOR2_X1 U875 ( .A(G128), .B(n1143), .ZN(G30) );
NAND3_X1 U876 ( .A1(n1183), .A2(n1013), .A3(n1184), .ZN(n1143) );
NOR3_X1 U877 ( .A1(n1034), .A2(n1193), .A3(n1019), .ZN(n1184) );
XOR2_X1 U878 ( .A(n1160), .B(n1194), .Z(G3) );
NAND2_X1 U879 ( .A1(KEYINPUT61), .A2(G101), .ZN(n1194) );
NAND3_X1 U880 ( .A1(n1014), .A2(n1166), .A3(n1173), .ZN(n1160) );
XOR2_X1 U881 ( .A(n1195), .B(n1196), .Z(G27) );
NOR2_X1 U882 ( .A1(KEYINPUT25), .A2(n1197), .ZN(n1196) );
NOR4_X1 U883 ( .A1(n1193), .A2(n1030), .A3(n1158), .A4(n1198), .ZN(n1195) );
INV_X1 U884 ( .A(n1029), .ZN(n1030) );
INV_X1 U885 ( .A(n1153), .ZN(n1193) );
NAND2_X1 U886 ( .A1(n1037), .A2(n1199), .ZN(n1153) );
NAND4_X1 U887 ( .A1(G902), .A2(G953), .A3(n1200), .A4(n1065), .ZN(n1199) );
INV_X1 U888 ( .A(G900), .ZN(n1065) );
XNOR2_X1 U889 ( .A(G122), .B(n1165), .ZN(G24) );
NAND4_X1 U890 ( .A1(n1174), .A2(n1003), .A3(n1186), .A4(n1187), .ZN(n1165) );
NOR2_X1 U891 ( .A1(n1201), .A2(n1202), .ZN(n1003) );
XNOR2_X1 U892 ( .A(G119), .B(n1164), .ZN(G21) );
NAND3_X1 U893 ( .A1(n1183), .A2(n1014), .A3(n1174), .ZN(n1164) );
AND2_X1 U894 ( .A1(n1202), .A2(n1201), .ZN(n1183) );
XOR2_X1 U895 ( .A(n1203), .B(n1204), .Z(G18) );
NAND3_X1 U896 ( .A1(n1174), .A2(n1013), .A3(n1205), .ZN(n1204) );
XOR2_X1 U897 ( .A(n1027), .B(KEYINPUT14), .Z(n1205) );
NOR2_X1 U898 ( .A1(n1187), .A2(n1206), .ZN(n1013) );
NOR2_X1 U899 ( .A1(n1158), .A2(n1180), .ZN(n1174) );
NAND2_X1 U900 ( .A1(n1010), .A2(n1179), .ZN(n1158) );
XOR2_X1 U901 ( .A(n1171), .B(n1207), .Z(G15) );
NAND2_X1 U902 ( .A1(KEYINPUT46), .A2(G113), .ZN(n1207) );
NAND2_X1 U903 ( .A1(n1172), .A2(n1179), .ZN(n1171) );
AND4_X1 U904 ( .A1(n1012), .A2(n1173), .A3(n1010), .A4(n1208), .ZN(n1172) );
NOR2_X1 U905 ( .A1(n1209), .A2(n1035), .ZN(n1010) );
INV_X1 U906 ( .A(n1036), .ZN(n1209) );
INV_X1 U907 ( .A(n1027), .ZN(n1173) );
NAND2_X1 U908 ( .A1(n1210), .A2(n1201), .ZN(n1027) );
INV_X1 U909 ( .A(n1198), .ZN(n1012) );
NAND2_X1 U910 ( .A1(n1206), .A2(n1187), .ZN(n1198) );
XOR2_X1 U911 ( .A(n1211), .B(n1163), .Z(G12) );
NAND3_X1 U912 ( .A1(n1014), .A2(n1166), .A3(n1029), .ZN(n1163) );
NOR2_X1 U913 ( .A1(n1201), .A2(n1210), .ZN(n1029) );
INV_X1 U914 ( .A(n1202), .ZN(n1210) );
NAND2_X1 U915 ( .A1(n1212), .A2(n1051), .ZN(n1202) );
NAND3_X1 U916 ( .A1(n1213), .A2(n1214), .A3(n1089), .ZN(n1051) );
XOR2_X1 U917 ( .A(n1052), .B(KEYINPUT39), .Z(n1212) );
NAND2_X1 U918 ( .A1(n1091), .A2(n1215), .ZN(n1052) );
NAND2_X1 U919 ( .A1(n1089), .A2(n1214), .ZN(n1215) );
XOR2_X1 U920 ( .A(n1216), .B(n1071), .Z(n1089) );
XOR2_X1 U921 ( .A(n1217), .B(n1218), .Z(n1216) );
NOR2_X1 U922 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
INV_X1 U923 ( .A(G221), .ZN(n1220) );
NAND2_X1 U924 ( .A1(n1221), .A2(n1222), .ZN(n1217) );
NAND2_X1 U925 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XOR2_X1 U926 ( .A(G146), .B(n1225), .Z(n1224) );
XOR2_X1 U927 ( .A(n1226), .B(G110), .Z(n1223) );
XOR2_X1 U928 ( .A(n1227), .B(KEYINPUT4), .Z(n1221) );
NAND2_X1 U929 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
XOR2_X1 U930 ( .A(n1211), .B(n1226), .Z(n1229) );
NAND2_X1 U931 ( .A1(KEYINPUT23), .A2(n1230), .ZN(n1226) );
XOR2_X1 U932 ( .A(G128), .B(G119), .Z(n1230) );
XOR2_X1 U933 ( .A(n1182), .B(n1225), .Z(n1228) );
INV_X1 U934 ( .A(n1213), .ZN(n1091) );
NAND2_X1 U935 ( .A1(G217), .A2(n1231), .ZN(n1213) );
NAND2_X1 U936 ( .A1(n1232), .A2(n1057), .ZN(n1201) );
NAND2_X1 U937 ( .A1(G472), .A2(n1233), .ZN(n1057) );
NAND2_X1 U938 ( .A1(n1234), .A2(n1214), .ZN(n1233) );
XOR2_X1 U939 ( .A(n1235), .B(n1108), .Z(n1234) );
XOR2_X1 U940 ( .A(KEYINPUT41), .B(n1056), .Z(n1232) );
NOR3_X1 U941 ( .A1(G472), .A2(G902), .A3(n1236), .ZN(n1056) );
XNOR2_X1 U942 ( .A(n1235), .B(n1108), .ZN(n1236) );
XOR2_X1 U943 ( .A(n1237), .B(n1238), .Z(n1108) );
XOR2_X1 U944 ( .A(n1239), .B(n1240), .Z(n1238) );
NAND2_X1 U945 ( .A1(KEYINPUT40), .A2(n1241), .ZN(n1240) );
NAND3_X1 U946 ( .A1(n1242), .A2(n997), .A3(n1243), .ZN(n1239) );
XOR2_X1 U947 ( .A(n1136), .B(KEYINPUT11), .Z(n1243) );
INV_X1 U948 ( .A(G210), .ZN(n1136) );
INV_X1 U949 ( .A(G237), .ZN(n1242) );
XNOR2_X1 U950 ( .A(G113), .B(G101), .ZN(n1237) );
XNOR2_X1 U951 ( .A(n1244), .B(n1112), .ZN(n1235) );
NAND2_X1 U952 ( .A1(KEYINPUT9), .A2(n1107), .ZN(n1244) );
NOR3_X1 U953 ( .A1(n1034), .A2(n1180), .A3(n1019), .ZN(n1166) );
INV_X1 U954 ( .A(n1179), .ZN(n1019) );
NOR2_X1 U955 ( .A1(n1022), .A2(n1021), .ZN(n1179) );
AND2_X1 U956 ( .A1(G214), .A2(n1245), .ZN(n1021) );
XOR2_X1 U957 ( .A(n1046), .B(n1049), .Z(n1022) );
AND2_X1 U958 ( .A1(G210), .A2(n1245), .ZN(n1049) );
NAND2_X1 U959 ( .A1(n1246), .A2(n1214), .ZN(n1245) );
XOR2_X1 U960 ( .A(KEYINPUT21), .B(G237), .Z(n1246) );
NAND2_X1 U961 ( .A1(n1247), .A2(n1214), .ZN(n1046) );
XNOR2_X1 U962 ( .A(n1135), .B(n1132), .ZN(n1247) );
XNOR2_X1 U963 ( .A(n1082), .B(KEYINPUT24), .ZN(n1132) );
XOR2_X1 U964 ( .A(n1248), .B(n1249), .Z(n1082) );
XOR2_X1 U965 ( .A(G101), .B(n1250), .Z(n1249) );
XOR2_X1 U966 ( .A(KEYINPUT1), .B(G110), .Z(n1250) );
XOR2_X1 U967 ( .A(n1251), .B(n1252), .Z(n1248) );
XOR2_X1 U968 ( .A(n1253), .B(n1241), .Z(n1251) );
XOR2_X1 U969 ( .A(G116), .B(G119), .Z(n1241) );
NAND3_X1 U970 ( .A1(n1254), .A2(n1255), .A3(KEYINPUT42), .ZN(n1253) );
NAND2_X1 U971 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
INV_X1 U972 ( .A(KEYINPUT63), .ZN(n1257) );
XOR2_X1 U973 ( .A(n1101), .B(G107), .Z(n1256) );
NAND3_X1 U974 ( .A1(G107), .A2(n1101), .A3(KEYINPUT63), .ZN(n1254) );
XOR2_X1 U975 ( .A(n1258), .B(n1259), .Z(n1135) );
XOR2_X1 U976 ( .A(n1197), .B(n1112), .Z(n1259) );
NAND2_X1 U977 ( .A1(n1260), .A2(n1261), .ZN(n1112) );
NAND2_X1 U978 ( .A1(G128), .A2(n1262), .ZN(n1261) );
XOR2_X1 U979 ( .A(KEYINPUT54), .B(n1263), .Z(n1260) );
NOR2_X1 U980 ( .A1(G128), .A2(n1262), .ZN(n1263) );
XOR2_X1 U981 ( .A(n1264), .B(n1265), .Z(n1262) );
XOR2_X1 U982 ( .A(G143), .B(KEYINPUT48), .Z(n1265) );
AND2_X1 U983 ( .A1(KEYINPUT50), .A2(n1182), .ZN(n1264) );
NAND2_X1 U984 ( .A1(G224), .A2(n997), .ZN(n1258) );
INV_X1 U985 ( .A(n1208), .ZN(n1180) );
NAND2_X1 U986 ( .A1(n1037), .A2(n1266), .ZN(n1208) );
NAND4_X1 U987 ( .A1(G902), .A2(n1267), .A3(n1200), .A4(n1268), .ZN(n1266) );
INV_X1 U988 ( .A(G898), .ZN(n1268) );
XOR2_X1 U989 ( .A(KEYINPUT8), .B(G953), .Z(n1267) );
NAND3_X1 U990 ( .A1(n1200), .A2(n997), .A3(G952), .ZN(n1037) );
NAND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1200) );
INV_X1 U992 ( .A(n1008), .ZN(n1034) );
NOR2_X1 U993 ( .A1(n1036), .A2(n1035), .ZN(n1008) );
AND2_X1 U994 ( .A1(G221), .A2(n1231), .ZN(n1035) );
NAND2_X1 U995 ( .A1(G234), .A2(n1214), .ZN(n1231) );
XOR2_X1 U996 ( .A(n1269), .B(G469), .Z(n1036) );
NAND2_X1 U997 ( .A1(n1270), .A2(n1214), .ZN(n1269) );
XOR2_X1 U998 ( .A(n1271), .B(n1116), .Z(n1270) );
XNOR2_X1 U999 ( .A(n1272), .B(n1273), .ZN(n1116) );
XOR2_X1 U1000 ( .A(G140), .B(G110), .Z(n1273) );
NAND2_X1 U1001 ( .A1(G227), .A2(n997), .ZN(n1272) );
NOR2_X1 U1002 ( .A1(KEYINPUT2), .A2(n1274), .ZN(n1271) );
XOR2_X1 U1003 ( .A(n1122), .B(n1275), .Z(n1274) );
XOR2_X1 U1004 ( .A(n1107), .B(n1125), .Z(n1275) );
INV_X1 U1005 ( .A(n1127), .ZN(n1125) );
XOR2_X1 U1006 ( .A(n1276), .B(n1277), .Z(n1127) );
XOR2_X1 U1007 ( .A(G101), .B(n1278), .Z(n1277) );
NOR2_X1 U1008 ( .A1(G107), .A2(KEYINPUT19), .ZN(n1278) );
XOR2_X1 U1009 ( .A(n1101), .B(KEYINPUT13), .Z(n1276) );
INV_X1 U1010 ( .A(G104), .ZN(n1101) );
XNOR2_X1 U1011 ( .A(n1279), .B(n1280), .ZN(n1107) );
NOR2_X1 U1012 ( .A1(KEYINPUT43), .A2(n1281), .ZN(n1280) );
XOR2_X1 U1013 ( .A(n1282), .B(n1283), .Z(n1281) );
XOR2_X1 U1014 ( .A(KEYINPUT16), .B(G134), .Z(n1283) );
INV_X1 U1015 ( .A(n1071), .ZN(n1282) );
XNOR2_X1 U1016 ( .A(G137), .B(KEYINPUT44), .ZN(n1071) );
XNOR2_X1 U1017 ( .A(G131), .B(KEYINPUT59), .ZN(n1279) );
XOR2_X1 U1018 ( .A(n1182), .B(n1284), .Z(n1122) );
INV_X1 U1019 ( .A(G146), .ZN(n1182) );
NOR2_X1 U1020 ( .A1(n1186), .A2(n1187), .ZN(n1014) );
XNOR2_X1 U1021 ( .A(n1285), .B(G475), .ZN(n1187) );
NAND2_X1 U1022 ( .A1(n1100), .A2(n1214), .ZN(n1285) );
XOR2_X1 U1023 ( .A(n1252), .B(n1286), .Z(n1100) );
XOR2_X1 U1024 ( .A(G104), .B(n1287), .Z(n1286) );
NOR2_X1 U1025 ( .A1(KEYINPUT53), .A2(n1288), .ZN(n1287) );
XOR2_X1 U1026 ( .A(n1289), .B(n1290), .Z(n1288) );
XOR2_X1 U1027 ( .A(G131), .B(n1291), .Z(n1290) );
NOR2_X1 U1028 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NOR2_X1 U1029 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
INV_X1 U1030 ( .A(n1225), .ZN(n1295) );
XOR2_X1 U1031 ( .A(KEYINPUT60), .B(n1296), .Z(n1294) );
NOR2_X1 U1032 ( .A1(n1225), .A2(n1297), .ZN(n1292) );
XOR2_X1 U1033 ( .A(KEYINPUT36), .B(n1296), .Z(n1297) );
NOR4_X1 U1034 ( .A1(G237), .A2(n1298), .A3(KEYINPUT29), .A4(G953), .ZN(n1296) );
INV_X1 U1035 ( .A(G214), .ZN(n1298) );
XNOR2_X1 U1036 ( .A(n1197), .B(G140), .ZN(n1225) );
INV_X1 U1037 ( .A(G125), .ZN(n1197) );
XOR2_X1 U1038 ( .A(G146), .B(G143), .Z(n1289) );
XOR2_X1 U1039 ( .A(G113), .B(G122), .Z(n1252) );
INV_X1 U1040 ( .A(n1206), .ZN(n1186) );
XOR2_X1 U1041 ( .A(n1299), .B(G478), .Z(n1206) );
NAND2_X1 U1042 ( .A1(n1300), .A2(n1214), .ZN(n1299) );
INV_X1 U1043 ( .A(G902), .ZN(n1214) );
XNOR2_X1 U1044 ( .A(n1096), .B(n1097), .ZN(n1300) );
XNOR2_X1 U1045 ( .A(n1301), .B(n1302), .ZN(n1097) );
XOR2_X1 U1046 ( .A(KEYINPUT17), .B(G134), .Z(n1302) );
XOR2_X1 U1047 ( .A(n1203), .B(G122), .Z(n1301) );
INV_X1 U1048 ( .A(G116), .ZN(n1203) );
XOR2_X1 U1049 ( .A(n1303), .B(n1304), .Z(n1096) );
NOR2_X1 U1050 ( .A1(n1219), .A2(n1305), .ZN(n1304) );
INV_X1 U1051 ( .A(G217), .ZN(n1305) );
NAND2_X1 U1052 ( .A1(G234), .A2(n997), .ZN(n1219) );
INV_X1 U1053 ( .A(G953), .ZN(n997) );
XOR2_X1 U1054 ( .A(n1306), .B(G107), .Z(n1303) );
NAND2_X1 U1055 ( .A1(KEYINPUT34), .A2(n1284), .ZN(n1306) );
XOR2_X1 U1056 ( .A(G128), .B(G143), .Z(n1284) );
INV_X1 U1057 ( .A(G110), .ZN(n1211) );
endmodule


