//Key = 1000100010011100111101110000000000111110100000111101001110111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327;

XOR2_X1 U723 ( .A(n1006), .B(n1007), .Z(G9) );
NOR2_X1 U724 ( .A1(n1008), .A2(n1009), .ZN(G75) );
NOR4_X1 U725 ( .A1(n1010), .A2(n1011), .A3(G953), .A4(n1012), .ZN(n1009) );
NOR4_X1 U726 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1011) );
NOR4_X1 U727 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1014) );
NOR2_X1 U728 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
XOR2_X1 U729 ( .A(n1023), .B(KEYINPUT31), .Z(n1021) );
NOR3_X1 U730 ( .A1(n1023), .A2(KEYINPUT28), .A3(n1024), .ZN(n1019) );
NOR2_X1 U731 ( .A1(n1025), .A2(n1026), .ZN(n1018) );
NOR3_X1 U732 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1025) );
NOR3_X1 U733 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
INV_X1 U734 ( .A(KEYINPUT22), .ZN(n1030) );
NOR2_X1 U735 ( .A1(KEYINPUT60), .A2(n1023), .ZN(n1027) );
NOR2_X1 U736 ( .A1(n1033), .A2(n1034), .ZN(n1013) );
NOR4_X1 U737 ( .A1(KEYINPUT22), .A2(n1026), .A3(n1031), .A4(n1032), .ZN(n1034) );
INV_X1 U738 ( .A(n1035), .ZN(n1026) );
NAND2_X1 U739 ( .A1(n1036), .A2(n1037), .ZN(n1010) );
NAND2_X1 U740 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U741 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND3_X1 U742 ( .A1(n1035), .A2(n1042), .A3(n1033), .ZN(n1041) );
NAND2_X1 U743 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U744 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U745 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U746 ( .A1(n1049), .A2(n1050), .ZN(n1043) );
NAND2_X1 U747 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND3_X1 U748 ( .A1(n1053), .A2(n1054), .A3(KEYINPUT60), .ZN(n1052) );
INV_X1 U749 ( .A(n1055), .ZN(n1051) );
NAND2_X1 U750 ( .A1(KEYINPUT28), .A2(n1056), .ZN(n1040) );
NAND4_X1 U751 ( .A1(n1033), .A2(n1057), .A3(n1045), .A4(n1049), .ZN(n1056) );
INV_X1 U752 ( .A(n1017), .ZN(n1033) );
NOR3_X1 U753 ( .A1(n1012), .A2(G953), .A3(G952), .ZN(n1008) );
AND4_X1 U754 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1012) );
NOR3_X1 U755 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
XOR2_X1 U756 ( .A(n1065), .B(KEYINPUT40), .Z(n1064) );
NOR2_X1 U757 ( .A1(G472), .A2(n1066), .ZN(n1063) );
NAND3_X1 U758 ( .A1(n1067), .A2(n1031), .A3(n1068), .ZN(n1062) );
NOR3_X1 U759 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1060) );
NOR2_X1 U760 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XNOR2_X1 U761 ( .A(n1074), .B(KEYINPUT26), .ZN(n1073) );
NOR2_X1 U762 ( .A1(n1074), .A2(n1075), .ZN(n1070) );
XOR2_X1 U763 ( .A(n1076), .B(n1077), .Z(n1069) );
NAND2_X1 U764 ( .A1(KEYINPUT58), .A2(n1078), .ZN(n1077) );
XOR2_X1 U765 ( .A(n1079), .B(G469), .Z(n1058) );
XOR2_X1 U766 ( .A(n1080), .B(n1081), .Z(G72) );
NOR3_X1 U767 ( .A1(n1082), .A2(KEYINPUT33), .A3(n1083), .ZN(n1081) );
NOR2_X1 U768 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U769 ( .A1(n1086), .A2(n1087), .ZN(n1080) );
NAND2_X1 U770 ( .A1(n1088), .A2(n1082), .ZN(n1087) );
XOR2_X1 U771 ( .A(n1089), .B(n1090), .Z(n1088) );
NAND3_X1 U772 ( .A1(n1090), .A2(G900), .A3(G953), .ZN(n1086) );
AND2_X1 U773 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U774 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U775 ( .A(KEYINPUT13), .B(n1095), .Z(n1091) );
NOR2_X1 U776 ( .A1(n1093), .A2(n1094), .ZN(n1095) );
XNOR2_X1 U777 ( .A(n1096), .B(n1097), .ZN(n1094) );
XOR2_X1 U778 ( .A(KEYINPUT52), .B(KEYINPUT42), .Z(n1097) );
XOR2_X1 U779 ( .A(n1098), .B(n1099), .Z(n1096) );
XOR2_X1 U780 ( .A(n1100), .B(n1101), .Z(G69) );
NAND4_X1 U781 ( .A1(KEYINPUT46), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1101) );
NAND3_X1 U782 ( .A1(n1105), .A2(n1106), .A3(n1082), .ZN(n1104) );
NAND2_X1 U783 ( .A1(G953), .A2(n1107), .ZN(n1103) );
NAND2_X1 U784 ( .A1(G898), .A2(n1105), .ZN(n1107) );
OR2_X1 U785 ( .A1(n1106), .A2(n1105), .ZN(n1102) );
NAND2_X1 U786 ( .A1(n1108), .A2(G953), .ZN(n1100) );
XOR2_X1 U787 ( .A(n1109), .B(KEYINPUT6), .Z(n1108) );
NAND2_X1 U788 ( .A1(G898), .A2(G224), .ZN(n1109) );
NOR2_X1 U789 ( .A1(n1110), .A2(n1111), .ZN(G66) );
NOR3_X1 U790 ( .A1(n1074), .A2(n1112), .A3(n1113), .ZN(n1111) );
AND3_X1 U791 ( .A1(n1114), .A2(n1072), .A3(n1115), .ZN(n1113) );
NOR2_X1 U792 ( .A1(n1116), .A2(n1114), .ZN(n1112) );
NOR2_X1 U793 ( .A1(n1036), .A2(n1075), .ZN(n1116) );
NOR2_X1 U794 ( .A1(n1110), .A2(n1117), .ZN(G63) );
XOR2_X1 U795 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND2_X1 U796 ( .A1(n1115), .A2(G478), .ZN(n1118) );
NOR2_X1 U797 ( .A1(n1110), .A2(n1120), .ZN(G60) );
XOR2_X1 U798 ( .A(n1121), .B(n1122), .Z(n1120) );
NAND2_X1 U799 ( .A1(n1115), .A2(G475), .ZN(n1121) );
XOR2_X1 U800 ( .A(G104), .B(n1123), .Z(G6) );
NOR2_X1 U801 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U802 ( .A(n1126), .B(KEYINPUT32), .Z(n1124) );
NOR2_X1 U803 ( .A1(n1110), .A2(n1127), .ZN(G57) );
XOR2_X1 U804 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U805 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U806 ( .A1(n1132), .A2(KEYINPUT1), .ZN(n1131) );
AND2_X1 U807 ( .A1(G472), .A2(n1115), .ZN(n1132) );
NOR2_X1 U808 ( .A1(n1133), .A2(n1134), .ZN(n1130) );
XOR2_X1 U809 ( .A(n1135), .B(KEYINPUT0), .Z(n1134) );
NAND2_X1 U810 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XNOR2_X1 U811 ( .A(n1138), .B(KEYINPUT23), .ZN(n1136) );
NOR2_X1 U812 ( .A1(n1137), .A2(n1138), .ZN(n1133) );
XOR2_X1 U813 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U814 ( .A1(n1110), .A2(n1141), .ZN(G54) );
XOR2_X1 U815 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U816 ( .A(KEYINPUT15), .B(n1144), .Z(n1143) );
NOR3_X1 U817 ( .A1(n1145), .A2(KEYINPUT27), .A3(n1146), .ZN(n1144) );
XOR2_X1 U818 ( .A(n1147), .B(KEYINPUT59), .Z(n1145) );
NAND2_X1 U819 ( .A1(n1148), .A2(n1099), .ZN(n1147) );
XOR2_X1 U820 ( .A(n1149), .B(n1150), .Z(n1142) );
NAND2_X1 U821 ( .A1(n1115), .A2(G469), .ZN(n1149) );
NOR2_X1 U822 ( .A1(n1110), .A2(n1151), .ZN(G51) );
XOR2_X1 U823 ( .A(n1152), .B(n1153), .Z(n1151) );
XNOR2_X1 U824 ( .A(n1140), .B(n1154), .ZN(n1153) );
XOR2_X1 U825 ( .A(n1155), .B(n1156), .Z(n1152) );
XNOR2_X1 U826 ( .A(KEYINPUT41), .B(n1157), .ZN(n1156) );
NOR2_X1 U827 ( .A1(G125), .A2(KEYINPUT7), .ZN(n1157) );
NAND2_X1 U828 ( .A1(n1115), .A2(n1078), .ZN(n1155) );
NOR2_X1 U829 ( .A1(n1158), .A2(n1036), .ZN(n1115) );
NOR2_X1 U830 ( .A1(n1106), .A2(n1089), .ZN(n1036) );
NAND4_X1 U831 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1089) );
AND4_X1 U832 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1162) );
NAND2_X1 U833 ( .A1(n1038), .A2(n1167), .ZN(n1161) );
NAND2_X1 U834 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XOR2_X1 U835 ( .A(KEYINPUT36), .B(n1170), .Z(n1168) );
NOR2_X1 U836 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XOR2_X1 U837 ( .A(KEYINPUT45), .B(n1015), .Z(n1171) );
INV_X1 U838 ( .A(n1049), .ZN(n1015) );
NAND2_X1 U839 ( .A1(n1173), .A2(n1174), .ZN(n1159) );
NAND4_X1 U840 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1106) );
AND4_X1 U841 ( .A1(n1179), .A2(n1180), .A3(n1007), .A4(n1181), .ZN(n1178) );
NAND4_X1 U842 ( .A1(n1182), .A2(n1055), .A3(n1183), .A4(n1035), .ZN(n1007) );
NOR2_X1 U843 ( .A1(n1184), .A2(n1185), .ZN(n1177) );
NOR2_X1 U844 ( .A1(n1186), .A2(n1126), .ZN(n1185) );
XOR2_X1 U845 ( .A(n1125), .B(KEYINPUT61), .Z(n1186) );
NAND4_X1 U846 ( .A1(n1187), .A2(n1055), .A3(n1035), .A4(n1188), .ZN(n1125) );
NOR2_X1 U847 ( .A1(n1082), .A2(G952), .ZN(n1110) );
XNOR2_X1 U848 ( .A(G146), .B(n1160), .ZN(G48) );
NAND3_X1 U849 ( .A1(n1187), .A2(n1028), .A3(n1189), .ZN(n1160) );
XNOR2_X1 U850 ( .A(G143), .B(n1166), .ZN(G45) );
NAND3_X1 U851 ( .A1(n1190), .A2(n1028), .A3(n1191), .ZN(n1166) );
XNOR2_X1 U852 ( .A(G140), .B(n1165), .ZN(G42) );
NAND4_X1 U853 ( .A1(n1038), .A2(n1192), .A3(n1193), .A4(n1187), .ZN(n1165) );
XNOR2_X1 U854 ( .A(G137), .B(n1194), .ZN(G39) );
NAND3_X1 U855 ( .A1(n1189), .A2(n1049), .A3(n1038), .ZN(n1194) );
XNOR2_X1 U856 ( .A(G134), .B(n1164), .ZN(G36) );
NAND3_X1 U857 ( .A1(n1191), .A2(n1183), .A3(n1038), .ZN(n1164) );
XOR2_X1 U858 ( .A(n1195), .B(n1196), .Z(G33) );
NAND2_X1 U859 ( .A1(n1197), .A2(n1038), .ZN(n1196) );
INV_X1 U860 ( .A(n1023), .ZN(n1038) );
NAND2_X1 U861 ( .A1(n1198), .A2(n1031), .ZN(n1023) );
XOR2_X1 U862 ( .A(n1169), .B(KEYINPUT38), .Z(n1197) );
NAND2_X1 U863 ( .A1(n1191), .A2(n1187), .ZN(n1169) );
AND2_X1 U864 ( .A1(n1192), .A2(n1057), .ZN(n1191) );
NAND2_X1 U865 ( .A1(n1199), .A2(n1200), .ZN(G30) );
NAND2_X1 U866 ( .A1(G128), .A2(n1201), .ZN(n1200) );
NAND2_X1 U867 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NAND2_X1 U868 ( .A1(KEYINPUT57), .A2(n1204), .ZN(n1203) );
NAND3_X1 U869 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1199) );
INV_X1 U870 ( .A(KEYINPUT57), .ZN(n1207) );
NAND2_X1 U871 ( .A1(n1163), .A2(n1204), .ZN(n1206) );
INV_X1 U872 ( .A(KEYINPUT44), .ZN(n1204) );
NAND2_X1 U873 ( .A1(n1202), .A2(n1208), .ZN(n1205) );
OR2_X1 U874 ( .A1(G128), .A2(KEYINPUT44), .ZN(n1208) );
INV_X1 U875 ( .A(n1163), .ZN(n1202) );
NAND3_X1 U876 ( .A1(n1183), .A2(n1028), .A3(n1189), .ZN(n1163) );
INV_X1 U877 ( .A(n1172), .ZN(n1189) );
NAND3_X1 U878 ( .A1(n1209), .A2(n1210), .A3(n1192), .ZN(n1172) );
AND2_X1 U879 ( .A1(n1055), .A2(n1174), .ZN(n1192) );
XNOR2_X1 U880 ( .A(n1184), .B(n1211), .ZN(G3) );
XNOR2_X1 U881 ( .A(G101), .B(KEYINPUT14), .ZN(n1211) );
AND4_X1 U882 ( .A1(n1057), .A2(n1182), .A3(n1055), .A4(n1049), .ZN(n1184) );
XOR2_X1 U883 ( .A(n1212), .B(n1213), .Z(G27) );
NAND2_X1 U884 ( .A1(KEYINPUT47), .A2(G125), .ZN(n1213) );
NAND2_X1 U885 ( .A1(n1173), .A2(n1214), .ZN(n1212) );
XNOR2_X1 U886 ( .A(KEYINPUT51), .B(n1174), .ZN(n1214) );
NAND2_X1 U887 ( .A1(n1017), .A2(n1215), .ZN(n1174) );
NAND4_X1 U888 ( .A1(G953), .A2(G902), .A3(n1216), .A4(n1085), .ZN(n1215) );
INV_X1 U889 ( .A(G900), .ZN(n1085) );
NOR4_X1 U890 ( .A1(n1016), .A2(n1022), .A3(n1047), .A4(n1126), .ZN(n1173) );
INV_X1 U891 ( .A(n1193), .ZN(n1022) );
XNOR2_X1 U892 ( .A(G122), .B(n1175), .ZN(G24) );
NAND3_X1 U893 ( .A1(n1217), .A2(n1035), .A3(n1190), .ZN(n1175) );
AND2_X1 U894 ( .A1(n1218), .A2(n1219), .ZN(n1190) );
XOR2_X1 U895 ( .A(n1059), .B(KEYINPUT49), .Z(n1218) );
NOR2_X1 U896 ( .A1(n1220), .A2(n1210), .ZN(n1035) );
XNOR2_X1 U897 ( .A(G119), .B(n1176), .ZN(G21) );
NAND4_X1 U898 ( .A1(n1217), .A2(n1049), .A3(n1209), .A4(n1210), .ZN(n1176) );
XNOR2_X1 U899 ( .A(G116), .B(n1180), .ZN(G18) );
NAND3_X1 U900 ( .A1(n1217), .A2(n1183), .A3(n1057), .ZN(n1180) );
INV_X1 U901 ( .A(n1048), .ZN(n1183) );
NAND2_X1 U902 ( .A1(n1059), .A2(n1219), .ZN(n1048) );
XOR2_X1 U903 ( .A(G113), .B(n1221), .Z(G15) );
NOR2_X1 U904 ( .A1(KEYINPUT43), .A2(n1181), .ZN(n1221) );
NAND3_X1 U905 ( .A1(n1217), .A2(n1187), .A3(n1057), .ZN(n1181) );
INV_X1 U906 ( .A(n1024), .ZN(n1057) );
NAND2_X1 U907 ( .A1(n1222), .A2(n1209), .ZN(n1024) );
XNOR2_X1 U908 ( .A(n1220), .B(KEYINPUT17), .ZN(n1209) );
AND2_X1 U909 ( .A1(n1045), .A2(n1182), .ZN(n1217) );
INV_X1 U910 ( .A(n1016), .ZN(n1045) );
NAND2_X1 U911 ( .A1(n1054), .A2(n1067), .ZN(n1016) );
XNOR2_X1 U912 ( .A(G110), .B(n1179), .ZN(G12) );
NAND4_X1 U913 ( .A1(n1193), .A2(n1182), .A3(n1055), .A4(n1049), .ZN(n1179) );
NAND2_X1 U914 ( .A1(n1223), .A2(n1224), .ZN(n1049) );
OR2_X1 U915 ( .A1(n1047), .A2(KEYINPUT19), .ZN(n1224) );
INV_X1 U916 ( .A(n1187), .ZN(n1047) );
NOR2_X1 U917 ( .A1(n1219), .A2(n1059), .ZN(n1187) );
INV_X1 U918 ( .A(n1065), .ZN(n1219) );
NAND3_X1 U919 ( .A1(n1059), .A2(n1065), .A3(KEYINPUT19), .ZN(n1223) );
XOR2_X1 U920 ( .A(n1225), .B(G478), .Z(n1065) );
NAND2_X1 U921 ( .A1(n1119), .A2(n1158), .ZN(n1225) );
XOR2_X1 U922 ( .A(n1226), .B(n1227), .Z(n1119) );
XOR2_X1 U923 ( .A(n1228), .B(n1229), .Z(n1227) );
NOR2_X1 U924 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U925 ( .A(n1232), .B(KEYINPUT56), .Z(n1231) );
NAND2_X1 U926 ( .A1(n1233), .A2(n1006), .ZN(n1232) );
NOR2_X1 U927 ( .A1(n1006), .A2(n1233), .ZN(n1230) );
XOR2_X1 U928 ( .A(KEYINPUT8), .B(n1234), .Z(n1233) );
INV_X1 U929 ( .A(G107), .ZN(n1006) );
NOR2_X1 U930 ( .A1(KEYINPUT9), .A2(n1235), .ZN(n1228) );
XOR2_X1 U931 ( .A(n1236), .B(n1237), .Z(n1235) );
NAND2_X1 U932 ( .A1(KEYINPUT35), .A2(n1238), .ZN(n1236) );
XOR2_X1 U933 ( .A(G143), .B(G128), .Z(n1238) );
NAND2_X1 U934 ( .A1(G217), .A2(n1239), .ZN(n1226) );
XOR2_X1 U935 ( .A(n1240), .B(G475), .Z(n1059) );
NAND2_X1 U936 ( .A1(n1122), .A2(n1158), .ZN(n1240) );
XOR2_X1 U937 ( .A(n1241), .B(n1242), .Z(n1122) );
XOR2_X1 U938 ( .A(n1243), .B(n1244), .Z(n1242) );
XNOR2_X1 U939 ( .A(n1245), .B(n1093), .ZN(n1244) );
XNOR2_X1 U940 ( .A(G125), .B(G140), .ZN(n1093) );
XOR2_X1 U941 ( .A(n1246), .B(n1247), .Z(n1243) );
NOR2_X1 U942 ( .A1(KEYINPUT39), .A2(n1248), .ZN(n1247) );
XOR2_X1 U943 ( .A(KEYINPUT50), .B(G113), .Z(n1248) );
NAND2_X1 U944 ( .A1(n1249), .A2(G214), .ZN(n1246) );
XOR2_X1 U945 ( .A(n1250), .B(n1251), .Z(n1241) );
XOR2_X1 U946 ( .A(KEYINPUT20), .B(G131), .Z(n1251) );
XOR2_X1 U947 ( .A(G122), .B(n1252), .Z(n1250) );
NOR2_X1 U948 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
INV_X1 U949 ( .A(n1067), .ZN(n1053) );
NAND2_X1 U950 ( .A1(G221), .A2(n1253), .ZN(n1067) );
XOR2_X1 U951 ( .A(n1254), .B(n1079), .Z(n1054) );
NAND3_X1 U952 ( .A1(n1255), .A2(n1158), .A3(n1256), .ZN(n1079) );
NAND3_X1 U953 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1256) );
NAND2_X1 U954 ( .A1(n1150), .A2(n1260), .ZN(n1258) );
NAND2_X1 U955 ( .A1(n1148), .A2(n1261), .ZN(n1260) );
OR2_X1 U956 ( .A1(n1150), .A2(n1146), .ZN(n1257) );
NOR2_X1 U957 ( .A1(n1099), .A2(n1148), .ZN(n1146) );
INV_X1 U958 ( .A(n1261), .ZN(n1099) );
NAND2_X1 U959 ( .A1(n1262), .A2(n1263), .ZN(n1255) );
NAND2_X1 U960 ( .A1(n1261), .A2(n1259), .ZN(n1263) );
INV_X1 U961 ( .A(KEYINPUT53), .ZN(n1259) );
XNOR2_X1 U962 ( .A(G128), .B(n1264), .ZN(n1261) );
NOR2_X1 U963 ( .A1(KEYINPUT29), .A2(n1245), .ZN(n1264) );
XOR2_X1 U964 ( .A(n1148), .B(n1150), .Z(n1262) );
XNOR2_X1 U965 ( .A(n1265), .B(n1266), .ZN(n1150) );
XOR2_X1 U966 ( .A(G140), .B(G110), .Z(n1266) );
XOR2_X1 U967 ( .A(n1139), .B(n1267), .Z(n1265) );
NOR2_X1 U968 ( .A1(G953), .A2(n1084), .ZN(n1267) );
INV_X1 U969 ( .A(G227), .ZN(n1084) );
AND3_X1 U970 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1148) );
NAND2_X1 U971 ( .A1(KEYINPUT11), .A2(n1271), .ZN(n1254) );
INV_X1 U972 ( .A(G469), .ZN(n1271) );
AND2_X1 U973 ( .A1(n1028), .A2(n1188), .ZN(n1182) );
NAND2_X1 U974 ( .A1(n1017), .A2(n1272), .ZN(n1188) );
NAND4_X1 U975 ( .A1(G953), .A2(G902), .A3(n1216), .A4(n1273), .ZN(n1272) );
INV_X1 U976 ( .A(G898), .ZN(n1273) );
NAND3_X1 U977 ( .A1(n1216), .A2(n1082), .A3(G952), .ZN(n1017) );
NAND2_X1 U978 ( .A1(G237), .A2(G234), .ZN(n1216) );
INV_X1 U979 ( .A(n1126), .ZN(n1028) );
NAND2_X1 U980 ( .A1(n1032), .A2(n1031), .ZN(n1126) );
NAND2_X1 U981 ( .A1(G214), .A2(n1274), .ZN(n1031) );
INV_X1 U982 ( .A(n1198), .ZN(n1032) );
XOR2_X1 U983 ( .A(n1076), .B(n1275), .Z(n1198) );
XOR2_X1 U984 ( .A(KEYINPUT25), .B(n1078), .Z(n1275) );
AND2_X1 U985 ( .A1(G210), .A2(n1274), .ZN(n1078) );
NAND2_X1 U986 ( .A1(n1276), .A2(n1158), .ZN(n1274) );
INV_X1 U987 ( .A(G237), .ZN(n1276) );
NAND2_X1 U988 ( .A1(n1277), .A2(n1158), .ZN(n1076) );
XOR2_X1 U989 ( .A(n1278), .B(n1279), .Z(n1277) );
XNOR2_X1 U990 ( .A(n1280), .B(n1154), .ZN(n1279) );
XNOR2_X1 U991 ( .A(n1105), .B(n1281), .ZN(n1154) );
AND2_X1 U992 ( .A1(n1082), .A2(G224), .ZN(n1281) );
XOR2_X1 U993 ( .A(n1282), .B(n1283), .Z(n1105) );
XOR2_X1 U994 ( .A(n1284), .B(n1285), .Z(n1283) );
NAND4_X1 U995 ( .A1(n1268), .A2(n1269), .A3(n1286), .A4(n1287), .ZN(n1285) );
OR2_X1 U996 ( .A1(n1270), .A2(KEYINPUT24), .ZN(n1287) );
OR2_X1 U997 ( .A1(n1288), .A2(G107), .ZN(n1270) );
NAND2_X1 U998 ( .A1(n1288), .A2(KEYINPUT24), .ZN(n1286) );
XOR2_X1 U999 ( .A(n1252), .B(n1289), .Z(n1288) );
NAND3_X1 U1000 ( .A1(n1289), .A2(G104), .A3(G107), .ZN(n1269) );
NAND3_X1 U1001 ( .A1(n1290), .A2(n1252), .A3(G107), .ZN(n1268) );
INV_X1 U1002 ( .A(G104), .ZN(n1252) );
XNOR2_X1 U1003 ( .A(n1234), .B(n1291), .ZN(n1282) );
XOR2_X1 U1004 ( .A(G116), .B(G122), .Z(n1234) );
NAND2_X1 U1005 ( .A1(KEYINPUT16), .A2(n1292), .ZN(n1280) );
XNOR2_X1 U1006 ( .A(n1140), .B(n1293), .ZN(n1292) );
XOR2_X1 U1007 ( .A(KEYINPUT62), .B(G125), .Z(n1293) );
XOR2_X1 U1008 ( .A(KEYINPUT34), .B(KEYINPUT18), .Z(n1278) );
NOR2_X1 U1009 ( .A1(n1220), .A2(n1222), .ZN(n1193) );
INV_X1 U1010 ( .A(n1210), .ZN(n1222) );
XOR2_X1 U1011 ( .A(n1074), .B(n1072), .Z(n1210) );
INV_X1 U1012 ( .A(n1075), .ZN(n1072) );
NAND2_X1 U1013 ( .A1(G217), .A2(n1253), .ZN(n1075) );
NAND2_X1 U1014 ( .A1(G234), .A2(n1158), .ZN(n1253) );
NOR2_X1 U1015 ( .A1(n1114), .A2(G902), .ZN(n1074) );
XOR2_X1 U1016 ( .A(n1294), .B(n1295), .Z(n1114) );
XOR2_X1 U1017 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U1018 ( .A(G137), .B(G128), .Z(n1297) );
XOR2_X1 U1019 ( .A(KEYINPUT20), .B(G146), .Z(n1296) );
XOR2_X1 U1020 ( .A(n1298), .B(n1291), .Z(n1294) );
XOR2_X1 U1021 ( .A(G110), .B(G119), .Z(n1291) );
XOR2_X1 U1022 ( .A(n1299), .B(n1300), .Z(n1298) );
AND2_X1 U1023 ( .A1(G221), .A2(n1239), .ZN(n1300) );
AND2_X1 U1024 ( .A1(G234), .A2(n1082), .ZN(n1239) );
INV_X1 U1025 ( .A(G953), .ZN(n1082) );
NAND2_X1 U1026 ( .A1(n1301), .A2(KEYINPUT21), .ZN(n1299) );
XNOR2_X1 U1027 ( .A(G140), .B(n1302), .ZN(n1301) );
NOR2_X1 U1028 ( .A1(G125), .A2(KEYINPUT5), .ZN(n1302) );
NAND2_X1 U1029 ( .A1(n1303), .A2(n1304), .ZN(n1220) );
NAND2_X1 U1030 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND2_X1 U1031 ( .A1(KEYINPUT48), .A2(G472), .ZN(n1306) );
INV_X1 U1032 ( .A(n1066), .ZN(n1305) );
NAND2_X1 U1033 ( .A1(n1307), .A2(KEYINPUT48), .ZN(n1303) );
INV_X1 U1034 ( .A(n1068), .ZN(n1307) );
NAND2_X1 U1035 ( .A1(G472), .A2(n1066), .ZN(n1068) );
NAND2_X1 U1036 ( .A1(n1308), .A2(n1158), .ZN(n1066) );
INV_X1 U1037 ( .A(G902), .ZN(n1158) );
XOR2_X1 U1038 ( .A(n1309), .B(n1128), .Z(n1308) );
AND2_X1 U1039 ( .A1(n1310), .A2(n1311), .ZN(n1128) );
NAND2_X1 U1040 ( .A1(n1289), .A2(n1312), .ZN(n1311) );
NAND2_X1 U1041 ( .A1(n1249), .A2(G210), .ZN(n1312) );
NAND3_X1 U1042 ( .A1(n1249), .A2(G210), .A3(n1290), .ZN(n1310) );
INV_X1 U1043 ( .A(n1289), .ZN(n1290) );
XNOR2_X1 U1044 ( .A(G101), .B(KEYINPUT2), .ZN(n1289) );
NOR2_X1 U1045 ( .A1(G953), .A2(G237), .ZN(n1249) );
NAND3_X1 U1046 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1309) );
NAND2_X1 U1047 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
OR3_X1 U1048 ( .A1(n1317), .A2(n1316), .A3(KEYINPUT63), .ZN(n1314) );
INV_X1 U1049 ( .A(n1137), .ZN(n1316) );
XOR2_X1 U1050 ( .A(n1318), .B(n1319), .Z(n1137) );
XOR2_X1 U1051 ( .A(KEYINPUT3), .B(G119), .Z(n1319) );
XOR2_X1 U1052 ( .A(n1320), .B(G116), .Z(n1318) );
NAND2_X1 U1053 ( .A1(KEYINPUT12), .A2(n1284), .ZN(n1320) );
INV_X1 U1054 ( .A(G113), .ZN(n1284) );
NAND2_X1 U1055 ( .A1(KEYINPUT55), .A2(n1321), .ZN(n1317) );
INV_X1 U1056 ( .A(n1322), .ZN(n1321) );
NAND2_X1 U1057 ( .A1(KEYINPUT63), .A2(n1322), .ZN(n1313) );
XOR2_X1 U1058 ( .A(n1323), .B(n1324), .Z(n1322) );
INV_X1 U1059 ( .A(n1139), .ZN(n1324) );
XOR2_X1 U1060 ( .A(n1098), .B(KEYINPUT30), .Z(n1139) );
XOR2_X1 U1061 ( .A(n1325), .B(n1326), .Z(n1098) );
XOR2_X1 U1062 ( .A(KEYINPUT54), .B(G137), .Z(n1326) );
XOR2_X1 U1063 ( .A(n1195), .B(n1237), .Z(n1325) );
XOR2_X1 U1064 ( .A(G134), .B(KEYINPUT4), .Z(n1237) );
INV_X1 U1065 ( .A(G131), .ZN(n1195) );
NAND2_X1 U1066 ( .A1(KEYINPUT37), .A2(n1140), .ZN(n1323) );
XNOR2_X1 U1067 ( .A(n1327), .B(n1245), .ZN(n1140) );
XNOR2_X1 U1068 ( .A(G143), .B(G146), .ZN(n1245) );
XNOR2_X1 U1069 ( .A(G128), .B(KEYINPUT10), .ZN(n1327) );
endmodule


