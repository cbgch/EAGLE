//Key = 0011001100101011100011101100011100010110101110000010110111110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408;

XOR2_X1 U775 ( .A(n1082), .B(n1083), .Z(G9) );
AND3_X1 U776 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1083) );
NAND2_X1 U777 ( .A1(KEYINPUT6), .A2(n1087), .ZN(n1082) );
NOR2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(G75) );
NOR3_X1 U779 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
NOR2_X1 U780 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NOR2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NOR2_X1 U782 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR3_X1 U783 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1097) );
NOR2_X1 U784 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR2_X1 U785 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NOR3_X1 U786 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1100) );
XNOR2_X1 U787 ( .A(KEYINPUT25), .B(n1109), .ZN(n1106) );
NOR2_X1 U788 ( .A1(n1110), .A2(n1109), .ZN(n1099) );
NOR4_X1 U789 ( .A1(n1111), .A2(n1109), .A3(n1103), .A4(n1112), .ZN(n1095) );
NOR2_X1 U790 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR2_X1 U791 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NAND3_X1 U792 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1090) );
NAND3_X1 U793 ( .A1(n1084), .A2(n1120), .A3(n1121), .ZN(n1119) );
NAND2_X1 U794 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
NAND3_X1 U795 ( .A1(n1124), .A2(n1125), .A3(n1085), .ZN(n1123) );
NAND2_X1 U796 ( .A1(KEYINPUT24), .A2(n1098), .ZN(n1125) );
INV_X1 U797 ( .A(n1126), .ZN(n1098) );
NAND2_X1 U798 ( .A1(n1127), .A2(n1128), .ZN(n1124) );
INV_X1 U799 ( .A(KEYINPUT24), .ZN(n1128) );
NAND2_X1 U800 ( .A1(n1129), .A2(n1112), .ZN(n1127) );
NAND2_X1 U801 ( .A1(n1126), .A2(n1130), .ZN(n1122) );
NOR2_X1 U802 ( .A1(n1112), .A2(n1131), .ZN(n1126) );
NOR3_X1 U803 ( .A1(n1132), .A2(G953), .A3(G952), .ZN(n1088) );
INV_X1 U804 ( .A(n1117), .ZN(n1132) );
NAND4_X1 U805 ( .A1(n1133), .A2(n1134), .A3(n1121), .A4(n1135), .ZN(n1117) );
NOR4_X1 U806 ( .A1(n1136), .A2(n1137), .A3(n1131), .A4(n1138), .ZN(n1135) );
XNOR2_X1 U807 ( .A(G472), .B(n1139), .ZN(n1138) );
INV_X1 U808 ( .A(n1129), .ZN(n1131) );
NOR2_X1 U809 ( .A1(G478), .A2(n1140), .ZN(n1137) );
XNOR2_X1 U810 ( .A(n1141), .B(KEYINPUT49), .ZN(n1140) );
NOR2_X1 U811 ( .A1(n1141), .A2(n1142), .ZN(n1136) );
INV_X1 U812 ( .A(G478), .ZN(n1142) );
XOR2_X1 U813 ( .A(n1143), .B(n1144), .Z(n1134) );
NOR2_X1 U814 ( .A1(KEYINPUT45), .A2(n1145), .ZN(n1144) );
XOR2_X1 U815 ( .A(KEYINPUT57), .B(n1146), .Z(n1133) );
NAND2_X1 U816 ( .A1(n1147), .A2(n1148), .ZN(G72) );
NAND3_X1 U817 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1148) );
XNOR2_X1 U818 ( .A(n1152), .B(n1153), .ZN(n1151) );
NAND3_X1 U819 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1147) );
XOR2_X1 U820 ( .A(n1153), .B(n1152), .Z(n1156) );
NAND2_X1 U821 ( .A1(n1157), .A2(n1158), .ZN(n1152) );
XNOR2_X1 U822 ( .A(KEYINPUT12), .B(n1118), .ZN(n1157) );
NAND2_X1 U823 ( .A1(n1159), .A2(n1160), .ZN(n1153) );
NAND2_X1 U824 ( .A1(G953), .A2(n1161), .ZN(n1160) );
XOR2_X1 U825 ( .A(n1162), .B(n1163), .Z(n1159) );
XNOR2_X1 U826 ( .A(n1164), .B(n1165), .ZN(n1163) );
NOR2_X1 U827 ( .A1(KEYINPUT4), .A2(n1166), .ZN(n1165) );
NAND2_X1 U828 ( .A1(n1167), .A2(KEYINPUT58), .ZN(n1164) );
XNOR2_X1 U829 ( .A(n1168), .B(n1169), .ZN(n1167) );
NAND2_X1 U830 ( .A1(KEYINPUT22), .A2(n1170), .ZN(n1168) );
XNOR2_X1 U831 ( .A(n1171), .B(n1172), .ZN(n1170) );
XOR2_X1 U832 ( .A(KEYINPUT23), .B(G140), .Z(n1162) );
OR2_X1 U833 ( .A1(n1149), .A2(KEYINPUT56), .ZN(n1155) );
NAND3_X1 U834 ( .A1(n1149), .A2(n1150), .A3(KEYINPUT56), .ZN(n1154) );
INV_X1 U835 ( .A(KEYINPUT60), .ZN(n1150) );
AND2_X1 U836 ( .A1(G953), .A2(n1173), .ZN(n1149) );
NAND2_X1 U837 ( .A1(G900), .A2(G227), .ZN(n1173) );
XOR2_X1 U838 ( .A(n1174), .B(n1175), .Z(G69) );
XOR2_X1 U839 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U840 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND2_X1 U841 ( .A1(n1180), .A2(n1118), .ZN(n1176) );
NAND3_X1 U842 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
XNOR2_X1 U843 ( .A(KEYINPUT17), .B(n1184), .ZN(n1183) );
INV_X1 U844 ( .A(n1185), .ZN(n1182) );
NAND2_X1 U845 ( .A1(G953), .A2(n1186), .ZN(n1174) );
NAND2_X1 U846 ( .A1(G898), .A2(G224), .ZN(n1186) );
NOR2_X1 U847 ( .A1(n1187), .A2(n1188), .ZN(G66) );
XOR2_X1 U848 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U849 ( .A1(n1191), .A2(n1192), .ZN(n1189) );
NOR2_X1 U850 ( .A1(n1187), .A2(n1193), .ZN(G63) );
NOR3_X1 U851 ( .A1(n1141), .A2(n1194), .A3(n1195), .ZN(n1193) );
AND3_X1 U852 ( .A1(n1196), .A2(G478), .A3(n1197), .ZN(n1195) );
NOR2_X1 U853 ( .A1(n1198), .A2(n1196), .ZN(n1194) );
AND2_X1 U854 ( .A1(n1092), .A2(G478), .ZN(n1198) );
NOR2_X1 U855 ( .A1(n1187), .A2(n1199), .ZN(G60) );
NOR3_X1 U856 ( .A1(n1143), .A2(n1200), .A3(n1201), .ZN(n1199) );
AND3_X1 U857 ( .A1(n1202), .A2(G475), .A3(n1197), .ZN(n1201) );
NOR2_X1 U858 ( .A1(n1203), .A2(n1202), .ZN(n1200) );
AND2_X1 U859 ( .A1(n1092), .A2(G475), .ZN(n1203) );
XOR2_X1 U860 ( .A(n1204), .B(n1205), .Z(G6) );
NOR2_X1 U861 ( .A1(KEYINPUT8), .A2(n1206), .ZN(n1205) );
NOR2_X1 U862 ( .A1(n1187), .A2(n1207), .ZN(G57) );
XOR2_X1 U863 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U864 ( .A(n1210), .B(KEYINPUT36), .Z(n1208) );
NAND2_X1 U865 ( .A1(n1197), .A2(G472), .ZN(n1210) );
NOR2_X1 U866 ( .A1(n1187), .A2(n1211), .ZN(G54) );
XOR2_X1 U867 ( .A(n1212), .B(n1213), .Z(n1211) );
XOR2_X1 U868 ( .A(n1214), .B(n1215), .Z(n1213) );
NOR2_X1 U869 ( .A1(KEYINPUT39), .A2(n1216), .ZN(n1215) );
AND2_X1 U870 ( .A1(G469), .A2(n1197), .ZN(n1214) );
INV_X1 U871 ( .A(n1192), .ZN(n1197) );
NOR2_X1 U872 ( .A1(n1187), .A2(n1217), .ZN(G51) );
XOR2_X1 U873 ( .A(n1218), .B(n1219), .Z(n1217) );
XNOR2_X1 U874 ( .A(n1220), .B(n1221), .ZN(n1219) );
NOR2_X1 U875 ( .A1(n1222), .A2(n1192), .ZN(n1220) );
NAND2_X1 U876 ( .A1(G902), .A2(n1092), .ZN(n1192) );
NAND3_X1 U877 ( .A1(n1181), .A2(n1223), .A3(n1224), .ZN(n1092) );
INV_X1 U878 ( .A(n1158), .ZN(n1224) );
NAND4_X1 U879 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1158) );
AND4_X1 U880 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1228) );
NAND2_X1 U881 ( .A1(n1114), .A2(n1233), .ZN(n1227) );
NAND2_X1 U882 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND4_X1 U883 ( .A1(n1105), .A2(n1130), .A3(n1121), .A4(n1236), .ZN(n1235) );
XOR2_X1 U884 ( .A(n1237), .B(KEYINPUT5), .Z(n1234) );
NAND2_X1 U885 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
INV_X1 U886 ( .A(n1240), .ZN(n1239) );
XOR2_X1 U887 ( .A(n1236), .B(KEYINPUT27), .Z(n1238) );
NAND3_X1 U888 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1225) );
XOR2_X1 U889 ( .A(KEYINPUT51), .B(n1244), .Z(n1223) );
NOR2_X1 U890 ( .A1(n1184), .A2(n1185), .ZN(n1244) );
NAND3_X1 U891 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1185) );
NAND4_X1 U892 ( .A1(n1130), .A2(n1104), .A3(n1248), .A4(n1249), .ZN(n1247) );
NAND2_X1 U893 ( .A1(KEYINPUT52), .A2(n1250), .ZN(n1249) );
NAND2_X1 U894 ( .A1(n1251), .A2(n1252), .ZN(n1248) );
INV_X1 U895 ( .A(KEYINPUT52), .ZN(n1252) );
NAND3_X1 U896 ( .A1(n1253), .A2(n1254), .A3(n1121), .ZN(n1251) );
NAND2_X1 U897 ( .A1(n1255), .A2(n1256), .ZN(n1184) );
OR4_X1 U898 ( .A1(n1109), .A2(n1257), .A3(n1250), .A4(KEYINPUT35), .ZN(n1256) );
INV_X1 U899 ( .A(n1084), .ZN(n1109) );
NAND2_X1 U900 ( .A1(n1258), .A2(KEYINPUT35), .ZN(n1255) );
AND4_X1 U901 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1181) );
NOR2_X1 U902 ( .A1(n1263), .A2(n1204), .ZN(n1262) );
AND3_X1 U903 ( .A1(n1084), .A2(n1086), .A3(n1130), .ZN(n1204) );
NAND4_X1 U904 ( .A1(n1264), .A2(n1085), .A3(n1265), .A4(n1266), .ZN(n1261) );
OR2_X1 U905 ( .A1(n1086), .A2(KEYINPUT18), .ZN(n1266) );
NAND2_X1 U906 ( .A1(KEYINPUT18), .A2(n1267), .ZN(n1265) );
NAND2_X1 U907 ( .A1(n1268), .A2(n1254), .ZN(n1267) );
XNOR2_X1 U908 ( .A(n1084), .B(KEYINPUT20), .ZN(n1264) );
NAND3_X1 U909 ( .A1(n1114), .A2(n1269), .A3(n1270), .ZN(n1260) );
INV_X1 U910 ( .A(KEYINPUT37), .ZN(n1270) );
NAND3_X1 U911 ( .A1(n1104), .A2(n1268), .A3(n1243), .ZN(n1269) );
NAND4_X1 U912 ( .A1(n1104), .A2(n1086), .A3(n1243), .A4(KEYINPUT37), .ZN(n1259) );
NOR2_X1 U913 ( .A1(n1271), .A2(n1272), .ZN(n1218) );
NOR2_X1 U914 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XOR2_X1 U915 ( .A(KEYINPUT30), .B(n1275), .Z(n1273) );
NOR2_X1 U916 ( .A1(n1276), .A2(n1277), .ZN(n1271) );
XOR2_X1 U917 ( .A(KEYINPUT1), .B(n1275), .Z(n1277) );
INV_X1 U918 ( .A(n1274), .ZN(n1276) );
XOR2_X1 U919 ( .A(n1278), .B(n1166), .Z(n1274) );
INV_X1 U920 ( .A(G125), .ZN(n1166) );
NOR2_X1 U921 ( .A1(n1118), .A2(G952), .ZN(n1187) );
XNOR2_X1 U922 ( .A(n1279), .B(n1280), .ZN(G48) );
NOR2_X1 U923 ( .A1(n1281), .A2(n1240), .ZN(n1280) );
NAND3_X1 U924 ( .A1(n1242), .A2(n1282), .A3(n1130), .ZN(n1240) );
XNOR2_X1 U925 ( .A(G143), .B(n1226), .ZN(G45) );
NAND4_X1 U926 ( .A1(n1257), .A2(n1104), .A3(n1283), .A4(n1282), .ZN(n1226) );
XNOR2_X1 U927 ( .A(G140), .B(n1232), .ZN(G42) );
NAND3_X1 U928 ( .A1(n1241), .A2(n1130), .A3(n1105), .ZN(n1232) );
XNOR2_X1 U929 ( .A(G137), .B(n1284), .ZN(G39) );
NAND3_X1 U930 ( .A1(n1243), .A2(n1241), .A3(n1285), .ZN(n1284) );
XNOR2_X1 U931 ( .A(n1242), .B(KEYINPUT31), .ZN(n1285) );
XNOR2_X1 U932 ( .A(G134), .B(n1231), .ZN(G36) );
NAND3_X1 U933 ( .A1(n1104), .A2(n1085), .A3(n1241), .ZN(n1231) );
XNOR2_X1 U934 ( .A(G131), .B(n1230), .ZN(G33) );
NAND3_X1 U935 ( .A1(n1130), .A2(n1104), .A3(n1241), .ZN(n1230) );
AND3_X1 U936 ( .A1(n1282), .A2(n1236), .A3(n1129), .ZN(n1241) );
NOR2_X1 U937 ( .A1(n1115), .A2(n1286), .ZN(n1129) );
INV_X1 U938 ( .A(n1116), .ZN(n1286) );
XNOR2_X1 U939 ( .A(G128), .B(n1229), .ZN(G30) );
NAND4_X1 U940 ( .A1(n1242), .A2(n1283), .A3(n1287), .A4(n1085), .ZN(n1229) );
NAND2_X1 U941 ( .A1(n1288), .A2(n1289), .ZN(G3) );
NAND2_X1 U942 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
XOR2_X1 U943 ( .A(KEYINPUT14), .B(n1292), .Z(n1288) );
NOR2_X1 U944 ( .A1(n1290), .A2(n1291), .ZN(n1292) );
AND3_X1 U945 ( .A1(n1086), .A2(n1293), .A3(n1104), .ZN(n1290) );
XNOR2_X1 U946 ( .A(KEYINPUT9), .B(n1094), .ZN(n1293) );
XNOR2_X1 U947 ( .A(G125), .B(n1294), .ZN(G27) );
NAND4_X1 U948 ( .A1(n1105), .A2(n1130), .A3(n1283), .A4(n1295), .ZN(n1294) );
XNOR2_X1 U949 ( .A(KEYINPUT54), .B(n1103), .ZN(n1295) );
INV_X1 U950 ( .A(n1121), .ZN(n1103) );
INV_X1 U951 ( .A(n1281), .ZN(n1283) );
NAND2_X1 U952 ( .A1(n1114), .A2(n1236), .ZN(n1281) );
NAND2_X1 U953 ( .A1(n1112), .A2(n1296), .ZN(n1236) );
NAND4_X1 U954 ( .A1(G902), .A2(G953), .A3(n1297), .A4(n1161), .ZN(n1296) );
INV_X1 U955 ( .A(G900), .ZN(n1161) );
XNOR2_X1 U956 ( .A(n1258), .B(n1298), .ZN(G24) );
NOR2_X1 U957 ( .A1(G122), .A2(KEYINPUT46), .ZN(n1298) );
AND3_X1 U958 ( .A1(n1257), .A2(n1084), .A3(n1299), .ZN(n1258) );
NOR2_X1 U959 ( .A1(n1300), .A2(n1301), .ZN(n1084) );
NOR2_X1 U960 ( .A1(n1302), .A2(n1303), .ZN(n1257) );
XNOR2_X1 U961 ( .A(G119), .B(n1245), .ZN(G21) );
NAND3_X1 U962 ( .A1(n1243), .A2(n1242), .A3(n1299), .ZN(n1245) );
AND2_X1 U963 ( .A1(n1301), .A2(n1300), .ZN(n1242) );
NAND2_X1 U964 ( .A1(n1304), .A2(n1305), .ZN(G18) );
NAND2_X1 U965 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XOR2_X1 U966 ( .A(KEYINPUT43), .B(n1308), .Z(n1304) );
NOR2_X1 U967 ( .A1(n1306), .A2(n1307), .ZN(n1308) );
INV_X1 U968 ( .A(n1246), .ZN(n1306) );
NAND3_X1 U969 ( .A1(n1104), .A2(n1085), .A3(n1299), .ZN(n1246) );
NOR2_X1 U970 ( .A1(n1303), .A2(n1309), .ZN(n1085) );
XNOR2_X1 U971 ( .A(G113), .B(n1310), .ZN(G15) );
NAND3_X1 U972 ( .A1(n1130), .A2(n1104), .A3(n1299), .ZN(n1310) );
INV_X1 U973 ( .A(n1250), .ZN(n1299) );
NAND3_X1 U974 ( .A1(n1114), .A2(n1253), .A3(n1121), .ZN(n1250) );
NOR2_X1 U975 ( .A1(n1108), .A2(n1311), .ZN(n1121) );
INV_X1 U976 ( .A(n1107), .ZN(n1311) );
NOR2_X1 U977 ( .A1(n1301), .A2(n1312), .ZN(n1104) );
AND2_X1 U978 ( .A1(n1313), .A2(n1303), .ZN(n1130) );
XNOR2_X1 U979 ( .A(n1309), .B(KEYINPUT16), .ZN(n1313) );
INV_X1 U980 ( .A(n1302), .ZN(n1309) );
XOR2_X1 U981 ( .A(G110), .B(n1263), .Z(G12) );
AND3_X1 U982 ( .A1(n1105), .A2(n1086), .A3(n1243), .ZN(n1263) );
INV_X1 U983 ( .A(n1094), .ZN(n1243) );
NAND2_X1 U984 ( .A1(n1303), .A2(n1302), .ZN(n1094) );
NAND2_X1 U985 ( .A1(n1314), .A2(n1315), .ZN(n1302) );
NAND2_X1 U986 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
NAND2_X1 U987 ( .A1(KEYINPUT3), .A2(n1318), .ZN(n1317) );
OR2_X1 U988 ( .A1(n1143), .A2(KEYINPUT11), .ZN(n1318) );
NAND2_X1 U989 ( .A1(n1143), .A2(n1319), .ZN(n1314) );
NAND2_X1 U990 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NAND2_X1 U991 ( .A1(n1145), .A2(KEYINPUT3), .ZN(n1321) );
INV_X1 U992 ( .A(n1316), .ZN(n1145) );
XOR2_X1 U993 ( .A(G475), .B(KEYINPUT29), .Z(n1316) );
INV_X1 U994 ( .A(KEYINPUT11), .ZN(n1320) );
NOR2_X1 U995 ( .A1(n1202), .A2(G902), .ZN(n1143) );
XOR2_X1 U996 ( .A(n1322), .B(n1323), .Z(n1202) );
XOR2_X1 U997 ( .A(G113), .B(n1324), .Z(n1323) );
XNOR2_X1 U998 ( .A(G131), .B(n1325), .ZN(n1324) );
XOR2_X1 U999 ( .A(n1326), .B(n1327), .Z(n1322) );
XNOR2_X1 U1000 ( .A(n1328), .B(n1329), .ZN(n1326) );
NAND2_X1 U1001 ( .A1(KEYINPUT15), .A2(n1206), .ZN(n1329) );
INV_X1 U1002 ( .A(G104), .ZN(n1206) );
NAND2_X1 U1003 ( .A1(n1330), .A2(KEYINPUT2), .ZN(n1328) );
XNOR2_X1 U1004 ( .A(G143), .B(n1331), .ZN(n1330) );
AND3_X1 U1005 ( .A1(G214), .A2(n1118), .A3(n1332), .ZN(n1331) );
XNOR2_X1 U1006 ( .A(n1141), .B(G478), .ZN(n1303) );
NOR2_X1 U1007 ( .A1(n1196), .A2(G902), .ZN(n1141) );
XOR2_X1 U1008 ( .A(n1333), .B(n1334), .Z(n1196) );
XOR2_X1 U1009 ( .A(n1335), .B(n1336), .Z(n1334) );
XNOR2_X1 U1010 ( .A(G128), .B(n1307), .ZN(n1336) );
XNOR2_X1 U1011 ( .A(n1337), .B(G134), .ZN(n1335) );
XOR2_X1 U1012 ( .A(n1338), .B(n1339), .Z(n1333) );
XNOR2_X1 U1013 ( .A(n1340), .B(n1341), .ZN(n1339) );
NOR2_X1 U1014 ( .A1(G122), .A2(KEYINPUT34), .ZN(n1341) );
NAND2_X1 U1015 ( .A1(KEYINPUT63), .A2(n1087), .ZN(n1340) );
INV_X1 U1016 ( .A(G107), .ZN(n1087) );
NAND2_X1 U1017 ( .A1(n1342), .A2(G217), .ZN(n1338) );
AND2_X1 U1018 ( .A1(n1114), .A2(n1268), .ZN(n1086) );
AND2_X1 U1019 ( .A1(n1287), .A2(n1253), .ZN(n1268) );
NAND2_X1 U1020 ( .A1(n1112), .A2(n1343), .ZN(n1253) );
NAND3_X1 U1021 ( .A1(n1178), .A2(n1297), .A3(G902), .ZN(n1343) );
NOR2_X1 U1022 ( .A1(n1118), .A2(G898), .ZN(n1178) );
NAND3_X1 U1023 ( .A1(n1297), .A2(n1118), .A3(G952), .ZN(n1112) );
NAND2_X1 U1024 ( .A1(G237), .A2(G234), .ZN(n1297) );
XNOR2_X1 U1025 ( .A(n1282), .B(KEYINPUT55), .ZN(n1287) );
INV_X1 U1026 ( .A(n1110), .ZN(n1282) );
NAND2_X1 U1027 ( .A1(n1108), .A2(n1107), .ZN(n1110) );
NAND2_X1 U1028 ( .A1(G221), .A2(n1344), .ZN(n1107) );
XNOR2_X1 U1029 ( .A(n1345), .B(G469), .ZN(n1108) );
NAND2_X1 U1030 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
XOR2_X1 U1031 ( .A(n1216), .B(n1348), .Z(n1346) );
XNOR2_X1 U1032 ( .A(n1349), .B(KEYINPUT53), .ZN(n1348) );
NAND2_X1 U1033 ( .A1(n1350), .A2(KEYINPUT21), .ZN(n1349) );
XNOR2_X1 U1034 ( .A(n1212), .B(KEYINPUT47), .ZN(n1350) );
XOR2_X1 U1035 ( .A(n1351), .B(n1352), .Z(n1212) );
XOR2_X1 U1036 ( .A(G140), .B(n1353), .Z(n1352) );
AND2_X1 U1037 ( .A1(n1118), .A2(G227), .ZN(n1353) );
XNOR2_X1 U1038 ( .A(n1354), .B(n1355), .ZN(n1216) );
XNOR2_X1 U1039 ( .A(n1356), .B(n1357), .ZN(n1355) );
XOR2_X1 U1040 ( .A(n1169), .B(n1358), .Z(n1354) );
XOR2_X1 U1041 ( .A(KEYINPUT59), .B(KEYINPUT40), .Z(n1358) );
NAND2_X1 U1042 ( .A1(n1359), .A2(n1360), .ZN(n1169) );
OR2_X1 U1043 ( .A1(n1361), .A2(G128), .ZN(n1360) );
XOR2_X1 U1044 ( .A(n1362), .B(KEYINPUT41), .Z(n1359) );
NAND2_X1 U1045 ( .A1(G128), .A2(n1361), .ZN(n1362) );
XNOR2_X1 U1046 ( .A(G146), .B(n1337), .ZN(n1361) );
INV_X1 U1047 ( .A(G143), .ZN(n1337) );
INV_X1 U1048 ( .A(n1254), .ZN(n1114) );
NAND2_X1 U1049 ( .A1(n1115), .A2(n1116), .ZN(n1254) );
NAND2_X1 U1050 ( .A1(G214), .A2(n1363), .ZN(n1116) );
XOR2_X1 U1051 ( .A(n1364), .B(n1222), .Z(n1115) );
NAND2_X1 U1052 ( .A1(G210), .A2(n1363), .ZN(n1222) );
NAND2_X1 U1053 ( .A1(n1332), .A2(n1347), .ZN(n1363) );
NAND2_X1 U1054 ( .A1(n1365), .A2(n1347), .ZN(n1364) );
XOR2_X1 U1055 ( .A(n1366), .B(KEYINPUT61), .Z(n1365) );
NAND2_X1 U1056 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
NAND2_X1 U1057 ( .A1(n1221), .A2(n1369), .ZN(n1368) );
NAND2_X1 U1058 ( .A1(KEYINPUT38), .A2(n1370), .ZN(n1369) );
OR2_X1 U1059 ( .A1(n1371), .A2(KEYINPUT19), .ZN(n1370) );
INV_X1 U1060 ( .A(n1179), .ZN(n1221) );
NAND2_X1 U1061 ( .A1(n1371), .A2(n1372), .ZN(n1367) );
NAND2_X1 U1062 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
NAND2_X1 U1063 ( .A1(KEYINPUT38), .A2(n1179), .ZN(n1374) );
XNOR2_X1 U1064 ( .A(n1375), .B(n1376), .ZN(n1179) );
XOR2_X1 U1065 ( .A(n1377), .B(n1378), .Z(n1376) );
XOR2_X1 U1066 ( .A(n1379), .B(G113), .Z(n1378) );
NAND2_X1 U1067 ( .A1(KEYINPUT44), .A2(n1291), .ZN(n1379) );
NAND2_X1 U1068 ( .A1(KEYINPUT42), .A2(n1325), .ZN(n1377) );
INV_X1 U1069 ( .A(G122), .ZN(n1325) );
XNOR2_X1 U1070 ( .A(n1380), .B(n1381), .ZN(n1375) );
XOR2_X1 U1071 ( .A(n1357), .B(n1351), .Z(n1381) );
XOR2_X1 U1072 ( .A(G104), .B(G107), .Z(n1357) );
INV_X1 U1073 ( .A(KEYINPUT19), .ZN(n1373) );
XOR2_X1 U1074 ( .A(n1382), .B(n1383), .Z(n1371) );
NOR2_X1 U1075 ( .A1(KEYINPUT33), .A2(n1278), .ZN(n1383) );
XNOR2_X1 U1076 ( .A(G125), .B(n1275), .ZN(n1382) );
AND2_X1 U1077 ( .A1(G224), .A2(n1118), .ZN(n1275) );
AND2_X1 U1078 ( .A1(n1312), .A2(n1301), .ZN(n1105) );
XOR2_X1 U1079 ( .A(n1146), .B(KEYINPUT26), .Z(n1301) );
XOR2_X1 U1080 ( .A(n1384), .B(n1191), .Z(n1146) );
NAND2_X1 U1081 ( .A1(G217), .A2(n1344), .ZN(n1191) );
NAND2_X1 U1082 ( .A1(G234), .A2(n1347), .ZN(n1344) );
OR2_X1 U1083 ( .A1(n1190), .A2(G902), .ZN(n1384) );
XNOR2_X1 U1084 ( .A(n1385), .B(n1386), .ZN(n1190) );
XNOR2_X1 U1085 ( .A(n1327), .B(n1387), .ZN(n1386) );
XOR2_X1 U1086 ( .A(n1388), .B(n1389), .Z(n1387) );
NOR2_X1 U1087 ( .A1(n1351), .A2(n1390), .ZN(n1389) );
XOR2_X1 U1088 ( .A(KEYINPUT28), .B(KEYINPUT13), .Z(n1390) );
XOR2_X1 U1089 ( .A(G110), .B(KEYINPUT32), .Z(n1351) );
NAND2_X1 U1090 ( .A1(G221), .A2(n1342), .ZN(n1388) );
AND2_X1 U1091 ( .A1(G234), .A2(n1118), .ZN(n1342) );
XOR2_X1 U1092 ( .A(G125), .B(n1391), .Z(n1327) );
XNOR2_X1 U1093 ( .A(n1279), .B(G140), .ZN(n1391) );
XNOR2_X1 U1094 ( .A(G119), .B(n1392), .ZN(n1385) );
XNOR2_X1 U1095 ( .A(n1171), .B(G128), .ZN(n1392) );
INV_X1 U1096 ( .A(n1300), .ZN(n1312) );
XOR2_X1 U1097 ( .A(n1393), .B(n1139), .Z(n1300) );
NAND2_X1 U1098 ( .A1(n1394), .A2(n1347), .ZN(n1139) );
INV_X1 U1099 ( .A(G902), .ZN(n1347) );
XNOR2_X1 U1100 ( .A(n1209), .B(KEYINPUT7), .ZN(n1394) );
XNOR2_X1 U1101 ( .A(n1395), .B(n1396), .ZN(n1209) );
XOR2_X1 U1102 ( .A(n1356), .B(n1397), .Z(n1396) );
XOR2_X1 U1103 ( .A(n1398), .B(n1399), .Z(n1397) );
NOR2_X1 U1104 ( .A1(G113), .A2(KEYINPUT48), .ZN(n1399) );
NAND3_X1 U1105 ( .A1(n1332), .A2(n1118), .A3(G210), .ZN(n1398) );
INV_X1 U1106 ( .A(G953), .ZN(n1118) );
INV_X1 U1107 ( .A(G237), .ZN(n1332) );
XOR2_X1 U1108 ( .A(n1400), .B(n1401), .Z(n1356) );
XNOR2_X1 U1109 ( .A(KEYINPUT0), .B(n1291), .ZN(n1401) );
INV_X1 U1110 ( .A(G101), .ZN(n1291) );
NAND2_X1 U1111 ( .A1(n1402), .A2(n1403), .ZN(n1400) );
NAND2_X1 U1112 ( .A1(n1172), .A2(G137), .ZN(n1403) );
NAND2_X1 U1113 ( .A1(n1404), .A2(n1171), .ZN(n1402) );
INV_X1 U1114 ( .A(G137), .ZN(n1171) );
XNOR2_X1 U1115 ( .A(n1172), .B(KEYINPUT62), .ZN(n1404) );
XOR2_X1 U1116 ( .A(G131), .B(G134), .Z(n1172) );
XNOR2_X1 U1117 ( .A(n1278), .B(n1380), .ZN(n1395) );
XNOR2_X1 U1118 ( .A(G119), .B(n1307), .ZN(n1380) );
INV_X1 U1119 ( .A(G116), .ZN(n1307) );
XNOR2_X1 U1120 ( .A(n1405), .B(G128), .ZN(n1278) );
NAND2_X1 U1121 ( .A1(n1406), .A2(n1407), .ZN(n1405) );
NAND2_X1 U1122 ( .A1(G143), .A2(n1279), .ZN(n1407) );
XOR2_X1 U1123 ( .A(KEYINPUT10), .B(n1408), .Z(n1406) );
NOR2_X1 U1124 ( .A1(G143), .A2(n1279), .ZN(n1408) );
INV_X1 U1125 ( .A(G146), .ZN(n1279) );
NAND2_X1 U1126 ( .A1(KEYINPUT50), .A2(G472), .ZN(n1393) );
endmodule


