//Key = 0100101100110001101101010110101011111001100110100111110101111111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312;

NAND2_X1 U723 ( .A1(n1004), .A2(n1005), .ZN(G9) );
NAND3_X1 U724 ( .A1(KEYINPUT35), .A2(n1006), .A3(n1007), .ZN(n1005) );
INV_X1 U725 ( .A(G107), .ZN(n1007) );
NAND2_X1 U726 ( .A1(G107), .A2(n1008), .ZN(n1004) );
NAND2_X1 U727 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND2_X1 U728 ( .A1(n1006), .A2(n1011), .ZN(n1010) );
INV_X1 U729 ( .A(KEYINPUT26), .ZN(n1011) );
NAND2_X1 U730 ( .A1(KEYINPUT26), .A2(n1012), .ZN(n1009) );
NAND2_X1 U731 ( .A1(KEYINPUT35), .A2(n1006), .ZN(n1012) );
AND3_X1 U732 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1006) );
XOR2_X1 U733 ( .A(KEYINPUT8), .B(n1016), .Z(n1014) );
NOR2_X1 U734 ( .A1(n1017), .A2(n1018), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
INV_X1 U736 ( .A(G952), .ZN(n1021) );
NAND4_X1 U737 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1019) );
NAND4_X1 U738 ( .A1(n1027), .A2(n1016), .A3(n1028), .A4(n1029), .ZN(n1024) );
NAND2_X1 U739 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND3_X1 U740 ( .A1(n1015), .A2(n1032), .A3(n1033), .ZN(n1031) );
NAND3_X1 U741 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1030) );
OR2_X1 U742 ( .A1(n1032), .A2(n1033), .ZN(n1035) );
NAND3_X1 U743 ( .A1(n1037), .A2(n1038), .A3(n1032), .ZN(n1034) );
NAND2_X1 U744 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U745 ( .A1(n1033), .A2(n1041), .ZN(n1023) );
NAND2_X1 U746 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND4_X1 U747 ( .A1(n1044), .A2(n1045), .A3(n1027), .A4(n1046), .ZN(n1043) );
NOR2_X1 U748 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U749 ( .A1(n1049), .A2(n1050), .ZN(n1045) );
NAND3_X1 U750 ( .A1(n1051), .A2(n1052), .A3(n1028), .ZN(n1044) );
INV_X1 U751 ( .A(n1049), .ZN(n1028) );
XOR2_X1 U752 ( .A(KEYINPUT7), .B(n1053), .Z(n1051) );
XOR2_X1 U753 ( .A(KEYINPUT57), .B(n1054), .Z(n1042) );
AND3_X1 U754 ( .A1(n1027), .A2(n1016), .A3(n1055), .ZN(n1054) );
INV_X1 U755 ( .A(n1056), .ZN(n1027) );
NOR3_X1 U756 ( .A1(n1057), .A2(G953), .A3(n1058), .ZN(n1017) );
INV_X1 U757 ( .A(n1025), .ZN(n1058) );
NAND4_X1 U758 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1025) );
NOR4_X1 U759 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1062) );
XOR2_X1 U760 ( .A(n1067), .B(n1068), .Z(n1066) );
XOR2_X1 U761 ( .A(n1069), .B(n1070), .Z(n1065) );
XNOR2_X1 U762 ( .A(n1071), .B(n1072), .ZN(n1064) );
NOR2_X1 U763 ( .A1(KEYINPUT14), .A2(n1073), .ZN(n1072) );
NOR2_X1 U764 ( .A1(n1039), .A2(n1047), .ZN(n1061) );
XOR2_X1 U765 ( .A(n1074), .B(n1075), .Z(n1060) );
NAND2_X1 U766 ( .A1(KEYINPUT18), .A2(n1076), .ZN(n1075) );
XOR2_X1 U767 ( .A(KEYINPUT21), .B(n1077), .Z(n1059) );
XOR2_X1 U768 ( .A(KEYINPUT2), .B(G952), .Z(n1057) );
XOR2_X1 U769 ( .A(n1078), .B(n1079), .Z(G72) );
NOR2_X1 U770 ( .A1(n1080), .A2(n1026), .ZN(n1079) );
NOR2_X1 U771 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XNOR2_X1 U772 ( .A(G227), .B(KEYINPUT5), .ZN(n1081) );
NAND2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(n1078) );
NAND2_X1 U774 ( .A1(n1085), .A2(n1026), .ZN(n1084) );
XOR2_X1 U775 ( .A(n1086), .B(n1022), .Z(n1085) );
NAND3_X1 U776 ( .A1(n1086), .A2(n1087), .A3(G953), .ZN(n1083) );
NOR2_X1 U777 ( .A1(KEYINPUT9), .A2(n1088), .ZN(n1086) );
XNOR2_X1 U778 ( .A(n1089), .B(n1090), .ZN(n1088) );
NOR2_X1 U779 ( .A1(KEYINPUT37), .A2(n1091), .ZN(n1090) );
XOR2_X1 U780 ( .A(n1092), .B(n1093), .Z(n1091) );
NOR2_X1 U781 ( .A1(KEYINPUT31), .A2(n1094), .ZN(n1093) );
NAND2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
NAND2_X1 U783 ( .A1(G131), .A2(n1097), .ZN(n1096) );
XOR2_X1 U784 ( .A(KEYINPUT46), .B(n1098), .Z(n1095) );
NOR2_X1 U785 ( .A1(G131), .A2(n1097), .ZN(n1098) );
XOR2_X1 U786 ( .A(n1099), .B(n1100), .Z(G69) );
XOR2_X1 U787 ( .A(n1101), .B(n1102), .Z(n1100) );
NAND2_X1 U788 ( .A1(KEYINPUT32), .A2(n1103), .ZN(n1102) );
NAND2_X1 U789 ( .A1(G953), .A2(n1104), .ZN(n1103) );
NAND2_X1 U790 ( .A1(n1105), .A2(G224), .ZN(n1104) );
XOR2_X1 U791 ( .A(n1106), .B(KEYINPUT52), .Z(n1105) );
NAND2_X1 U792 ( .A1(n1107), .A2(n1108), .ZN(n1101) );
NAND2_X1 U793 ( .A1(n1109), .A2(n1106), .ZN(n1108) );
XOR2_X1 U794 ( .A(n1026), .B(KEYINPUT61), .Z(n1109) );
XOR2_X1 U795 ( .A(n1110), .B(n1111), .Z(n1107) );
XNOR2_X1 U796 ( .A(n1112), .B(n1113), .ZN(n1111) );
XOR2_X1 U797 ( .A(n1114), .B(n1115), .Z(n1110) );
XOR2_X1 U798 ( .A(KEYINPUT58), .B(KEYINPUT29), .Z(n1115) );
NAND2_X1 U799 ( .A1(n1116), .A2(KEYINPUT25), .ZN(n1114) );
XOR2_X1 U800 ( .A(n1117), .B(KEYINPUT1), .Z(n1116) );
NAND2_X1 U801 ( .A1(n1026), .A2(n1020), .ZN(n1099) );
NOR2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(G66) );
NOR3_X1 U803 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
NOR3_X1 U804 ( .A1(n1123), .A2(n1068), .A3(n1124), .ZN(n1122) );
NOR2_X1 U805 ( .A1(n1125), .A2(n1126), .ZN(n1121) );
INV_X1 U806 ( .A(n1123), .ZN(n1126) );
NOR2_X1 U807 ( .A1(n1127), .A2(n1068), .ZN(n1125) );
NOR2_X1 U808 ( .A1(n1022), .A2(n1020), .ZN(n1127) );
NOR2_X1 U809 ( .A1(n1118), .A2(n1128), .ZN(G63) );
XOR2_X1 U810 ( .A(n1129), .B(n1130), .Z(n1128) );
AND2_X1 U811 ( .A1(G478), .A2(n1131), .ZN(n1129) );
NOR2_X1 U812 ( .A1(n1132), .A2(n1133), .ZN(G60) );
XNOR2_X1 U813 ( .A(n1118), .B(KEYINPUT4), .ZN(n1133) );
XNOR2_X1 U814 ( .A(n1134), .B(n1135), .ZN(n1132) );
AND2_X1 U815 ( .A1(G475), .A2(n1131), .ZN(n1135) );
XOR2_X1 U816 ( .A(G104), .B(n1136), .Z(G6) );
NOR2_X1 U817 ( .A1(n1118), .A2(n1137), .ZN(G57) );
XOR2_X1 U818 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U819 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U820 ( .A(KEYINPUT15), .B(n1142), .Z(n1141) );
NOR2_X1 U821 ( .A1(KEYINPUT42), .A2(n1143), .ZN(n1140) );
XOR2_X1 U822 ( .A(n1144), .B(n1145), .Z(n1138) );
XOR2_X1 U823 ( .A(n1146), .B(n1094), .Z(n1144) );
NAND3_X1 U824 ( .A1(n1131), .A2(G472), .A3(KEYINPUT50), .ZN(n1146) );
INV_X1 U825 ( .A(n1124), .ZN(n1131) );
NOR2_X1 U826 ( .A1(n1118), .A2(n1147), .ZN(G54) );
XOR2_X1 U827 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U828 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U829 ( .A1(n1073), .A2(n1124), .ZN(n1151) );
INV_X1 U830 ( .A(G469), .ZN(n1073) );
XNOR2_X1 U831 ( .A(KEYINPUT62), .B(n1152), .ZN(n1148) );
NOR2_X1 U832 ( .A1(KEYINPUT20), .A2(n1153), .ZN(n1152) );
XOR2_X1 U833 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U834 ( .A(G140), .B(n1156), .Z(n1155) );
NAND2_X1 U835 ( .A1(KEYINPUT30), .A2(n1157), .ZN(n1154) );
NOR2_X1 U836 ( .A1(n1118), .A2(n1158), .ZN(G51) );
XOR2_X1 U837 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U838 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U839 ( .A1(n1074), .A2(n1124), .ZN(n1162) );
NAND2_X1 U840 ( .A1(G902), .A2(n1163), .ZN(n1124) );
OR2_X1 U841 ( .A1(n1020), .A2(n1022), .ZN(n1163) );
NAND2_X1 U842 ( .A1(n1164), .A2(n1165), .ZN(n1022) );
AND4_X1 U843 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
OR2_X1 U844 ( .A1(n1170), .A2(n1171), .ZN(n1168) );
NOR2_X1 U845 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
NOR2_X1 U846 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NOR3_X1 U847 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1172) );
NAND3_X1 U848 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1176) );
NOR4_X1 U849 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1164) );
NOR2_X1 U850 ( .A1(n1186), .A2(n1180), .ZN(n1185) );
INV_X1 U851 ( .A(KEYINPUT43), .ZN(n1180) );
NAND4_X1 U852 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1020) );
NOR4_X1 U853 ( .A1(n1191), .A2(n1136), .A3(n1192), .A4(n1193), .ZN(n1190) );
INV_X1 U854 ( .A(n1194), .ZN(n1193) );
NOR4_X1 U855 ( .A1(n1195), .A2(n1196), .A3(n1048), .A4(n1052), .ZN(n1192) );
NOR2_X1 U856 ( .A1(KEYINPUT40), .A2(n1197), .ZN(n1196) );
NOR3_X1 U857 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1197) );
NOR2_X1 U858 ( .A1(n1013), .A2(n1201), .ZN(n1195) );
INV_X1 U859 ( .A(KEYINPUT40), .ZN(n1201) );
AND3_X1 U860 ( .A1(n1013), .A2(n1016), .A3(n1202), .ZN(n1136) );
NOR2_X1 U861 ( .A1(n1203), .A2(n1204), .ZN(n1189) );
NAND3_X1 U862 ( .A1(n1013), .A2(n1016), .A3(n1015), .ZN(n1187) );
XOR2_X1 U863 ( .A(n1205), .B(G125), .Z(n1159) );
NAND2_X1 U864 ( .A1(KEYINPUT53), .A2(n1206), .ZN(n1205) );
NOR2_X1 U865 ( .A1(n1026), .A2(G952), .ZN(n1118) );
XNOR2_X1 U866 ( .A(G146), .B(n1186), .ZN(G48) );
NAND2_X1 U867 ( .A1(n1207), .A2(n1202), .ZN(n1186) );
INV_X1 U868 ( .A(n1171), .ZN(n1202) );
XNOR2_X1 U869 ( .A(G143), .B(n1167), .ZN(G45) );
NAND4_X1 U870 ( .A1(n1181), .A2(n1208), .A3(n1209), .A4(n1053), .ZN(n1167) );
NOR2_X1 U871 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U872 ( .A(n1212), .B(n1166), .Z(G42) );
OR3_X1 U873 ( .A1(n1052), .A2(n1171), .A3(n1175), .ZN(n1166) );
XOR2_X1 U874 ( .A(G137), .B(n1184), .Z(G39) );
NOR3_X1 U875 ( .A1(n1177), .A2(n1048), .A3(n1175), .ZN(n1184) );
XOR2_X1 U876 ( .A(G134), .B(n1183), .Z(G36) );
NOR3_X1 U877 ( .A1(n1174), .A2(n1213), .A3(n1175), .ZN(n1183) );
INV_X1 U878 ( .A(n1015), .ZN(n1213) );
XOR2_X1 U879 ( .A(G131), .B(n1214), .Z(G33) );
NOR4_X1 U880 ( .A1(KEYINPUT38), .A2(n1174), .A3(n1171), .A4(n1175), .ZN(n1214) );
NAND2_X1 U881 ( .A1(n1208), .A2(n1033), .ZN(n1175) );
NOR2_X1 U882 ( .A1(n1215), .A2(n1039), .ZN(n1033) );
INV_X1 U883 ( .A(n1040), .ZN(n1215) );
XOR2_X1 U884 ( .A(G128), .B(n1182), .Z(G30) );
AND2_X1 U885 ( .A1(n1207), .A2(n1015), .ZN(n1182) );
AND3_X1 U886 ( .A1(n1181), .A2(n1216), .A3(n1208), .ZN(n1207) );
AND2_X1 U887 ( .A1(n1179), .A2(n1178), .ZN(n1208) );
XOR2_X1 U888 ( .A(G101), .B(n1191), .Z(G3) );
AND3_X1 U889 ( .A1(n1053), .A2(n1013), .A3(n1036), .ZN(n1191) );
XOR2_X1 U890 ( .A(n1217), .B(n1169), .Z(G27) );
NAND4_X1 U891 ( .A1(n1181), .A2(n1055), .A3(n1218), .A4(n1178), .ZN(n1169) );
NAND2_X1 U892 ( .A1(n1056), .A2(n1219), .ZN(n1178) );
NAND4_X1 U893 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1221), .ZN(n1219) );
INV_X1 U894 ( .A(n1087), .ZN(n1220) );
XOR2_X1 U895 ( .A(n1082), .B(KEYINPUT28), .Z(n1087) );
INV_X1 U896 ( .A(G900), .ZN(n1082) );
XNOR2_X1 U897 ( .A(n1222), .B(n1188), .ZN(G24) );
NAND4_X1 U898 ( .A1(n1223), .A2(n1016), .A3(n1077), .A4(n1063), .ZN(n1188) );
INV_X1 U899 ( .A(n1211), .ZN(n1077) );
INV_X1 U900 ( .A(n1050), .ZN(n1016) );
NAND2_X1 U901 ( .A1(n1224), .A2(n1225), .ZN(n1050) );
NAND2_X1 U902 ( .A1(KEYINPUT51), .A2(n1226), .ZN(n1222) );
INV_X1 U903 ( .A(G122), .ZN(n1226) );
NAND2_X1 U904 ( .A1(n1227), .A2(n1228), .ZN(G21) );
NAND2_X1 U905 ( .A1(G119), .A2(n1229), .ZN(n1228) );
XOR2_X1 U906 ( .A(n1230), .B(KEYINPUT12), .Z(n1227) );
NAND2_X1 U907 ( .A1(n1204), .A2(n1231), .ZN(n1230) );
INV_X1 U908 ( .A(n1229), .ZN(n1204) );
NAND3_X1 U909 ( .A1(n1223), .A2(n1036), .A3(n1216), .ZN(n1229) );
INV_X1 U910 ( .A(n1177), .ZN(n1216) );
NAND2_X1 U911 ( .A1(n1232), .A2(n1233), .ZN(n1177) );
XOR2_X1 U912 ( .A(G116), .B(n1203), .Z(G18) );
AND3_X1 U913 ( .A1(n1053), .A2(n1015), .A3(n1223), .ZN(n1203) );
NOR4_X1 U914 ( .A1(n1037), .A2(n1049), .A3(n1047), .A4(n1200), .ZN(n1223) );
INV_X1 U915 ( .A(n1234), .ZN(n1200) );
INV_X1 U916 ( .A(n1181), .ZN(n1037) );
XNOR2_X1 U917 ( .A(n1199), .B(KEYINPUT44), .ZN(n1181) );
NOR2_X1 U918 ( .A1(n1063), .A2(n1211), .ZN(n1015) );
XOR2_X1 U919 ( .A(n1235), .B(n1194), .Z(G15) );
NAND4_X1 U920 ( .A1(n1055), .A2(n1053), .A3(n1199), .A4(n1234), .ZN(n1194) );
INV_X1 U921 ( .A(n1174), .ZN(n1053) );
NAND2_X1 U922 ( .A1(n1224), .A2(n1233), .ZN(n1174) );
NOR3_X1 U923 ( .A1(n1049), .A2(n1047), .A3(n1171), .ZN(n1055) );
NAND2_X1 U924 ( .A1(n1211), .A2(n1063), .ZN(n1171) );
INV_X1 U925 ( .A(n1210), .ZN(n1063) );
INV_X1 U926 ( .A(n1032), .ZN(n1047) );
XOR2_X1 U927 ( .A(n1157), .B(n1236), .Z(G12) );
NAND3_X1 U928 ( .A1(n1036), .A2(n1013), .A3(n1218), .ZN(n1236) );
INV_X1 U929 ( .A(n1052), .ZN(n1218) );
NAND2_X1 U930 ( .A1(n1232), .A2(n1225), .ZN(n1052) );
XOR2_X1 U931 ( .A(n1233), .B(KEYINPUT39), .Z(n1225) );
XNOR2_X1 U932 ( .A(n1237), .B(n1238), .ZN(n1233) );
XNOR2_X1 U933 ( .A(KEYINPUT23), .B(n1070), .ZN(n1238) );
NAND2_X1 U934 ( .A1(n1239), .A2(n1240), .ZN(n1070) );
XOR2_X1 U935 ( .A(n1241), .B(n1242), .Z(n1239) );
XNOR2_X1 U936 ( .A(n1143), .B(n1145), .ZN(n1242) );
XOR2_X1 U937 ( .A(G101), .B(n1243), .Z(n1145) );
NOR3_X1 U938 ( .A1(n1244), .A2(G237), .A3(n1245), .ZN(n1243) );
INV_X1 U939 ( .A(G210), .ZN(n1245) );
XOR2_X1 U940 ( .A(KEYINPUT27), .B(G953), .Z(n1244) );
XOR2_X1 U941 ( .A(n1142), .B(n1246), .Z(n1241) );
NOR2_X1 U942 ( .A1(KEYINPUT41), .A2(n1094), .ZN(n1246) );
AND2_X1 U943 ( .A1(n1247), .A2(n1248), .ZN(n1142) );
NAND2_X1 U944 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
XOR2_X1 U945 ( .A(KEYINPUT33), .B(n1251), .Z(n1247) );
NOR2_X1 U946 ( .A1(n1249), .A2(n1250), .ZN(n1251) );
XOR2_X1 U947 ( .A(KEYINPUT6), .B(n1252), .Z(n1250) );
NAND2_X1 U948 ( .A1(KEYINPUT19), .A2(n1069), .ZN(n1237) );
INV_X1 U949 ( .A(G472), .ZN(n1069) );
XNOR2_X1 U950 ( .A(n1224), .B(KEYINPUT54), .ZN(n1232) );
XNOR2_X1 U951 ( .A(n1068), .B(n1253), .ZN(n1224) );
NOR2_X1 U952 ( .A1(KEYINPUT56), .A2(n1254), .ZN(n1253) );
XOR2_X1 U953 ( .A(KEYINPUT45), .B(n1120), .Z(n1254) );
INV_X1 U954 ( .A(n1067), .ZN(n1120) );
NAND2_X1 U955 ( .A1(n1123), .A2(n1240), .ZN(n1067) );
XOR2_X1 U956 ( .A(n1255), .B(n1256), .Z(n1123) );
XOR2_X1 U957 ( .A(n1257), .B(n1258), .Z(n1256) );
XOR2_X1 U958 ( .A(n1259), .B(n1260), .Z(n1258) );
NOR2_X1 U959 ( .A1(KEYINPUT17), .A2(n1261), .ZN(n1260) );
XOR2_X1 U960 ( .A(G110), .B(n1262), .Z(n1261) );
XOR2_X1 U961 ( .A(G128), .B(G119), .Z(n1262) );
NAND2_X1 U962 ( .A1(G221), .A2(n1263), .ZN(n1259) );
XNOR2_X1 U963 ( .A(G137), .B(n1264), .ZN(n1255) );
XOR2_X1 U964 ( .A(KEYINPUT47), .B(G146), .Z(n1264) );
NAND2_X1 U965 ( .A1(G217), .A2(n1265), .ZN(n1068) );
AND3_X1 U966 ( .A1(n1179), .A2(n1234), .A3(n1199), .ZN(n1013) );
NOR2_X1 U967 ( .A1(n1040), .A2(n1039), .ZN(n1199) );
AND2_X1 U968 ( .A1(G214), .A2(n1266), .ZN(n1039) );
XNOR2_X1 U969 ( .A(n1076), .B(n1074), .ZN(n1040) );
NAND2_X1 U970 ( .A1(G210), .A2(n1266), .ZN(n1074) );
NAND2_X1 U971 ( .A1(n1240), .A2(n1267), .ZN(n1266) );
NAND2_X1 U972 ( .A1(n1268), .A2(n1240), .ZN(n1076) );
XOR2_X1 U973 ( .A(n1161), .B(n1269), .Z(n1268) );
XOR2_X1 U974 ( .A(n1217), .B(n1094), .Z(n1269) );
INV_X1 U975 ( .A(n1206), .ZN(n1094) );
XOR2_X1 U976 ( .A(n1270), .B(n1271), .Z(n1161) );
AND2_X1 U977 ( .A1(n1026), .A2(G224), .ZN(n1271) );
NAND2_X1 U978 ( .A1(n1272), .A2(n1273), .ZN(n1270) );
NAND2_X1 U979 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XOR2_X1 U980 ( .A(KEYINPUT48), .B(n1112), .Z(n1275) );
XOR2_X1 U981 ( .A(n1113), .B(n1276), .Z(n1274) );
INV_X1 U982 ( .A(n1117), .ZN(n1276) );
NAND2_X1 U983 ( .A1(n1277), .A2(n1278), .ZN(n1272) );
XOR2_X1 U984 ( .A(n1113), .B(n1117), .Z(n1278) );
XOR2_X1 U985 ( .A(n1249), .B(n1252), .Z(n1117) );
XNOR2_X1 U986 ( .A(G116), .B(n1231), .ZN(n1252) );
INV_X1 U987 ( .A(G119), .ZN(n1231) );
XOR2_X1 U988 ( .A(n1235), .B(KEYINPUT13), .Z(n1249) );
XOR2_X1 U989 ( .A(n1279), .B(KEYINPUT10), .Z(n1113) );
XOR2_X1 U990 ( .A(KEYINPUT59), .B(n1112), .Z(n1277) );
XNOR2_X1 U991 ( .A(n1157), .B(G122), .ZN(n1112) );
NAND2_X1 U992 ( .A1(n1056), .A2(n1280), .ZN(n1234) );
NAND4_X1 U993 ( .A1(G953), .A2(G902), .A3(n1221), .A4(n1106), .ZN(n1280) );
INV_X1 U994 ( .A(G898), .ZN(n1106) );
NAND3_X1 U995 ( .A1(n1221), .A2(n1026), .A3(G952), .ZN(n1056) );
NAND2_X1 U996 ( .A1(G237), .A2(n1281), .ZN(n1221) );
INV_X1 U997 ( .A(n1198), .ZN(n1179) );
NAND2_X1 U998 ( .A1(n1049), .A2(n1032), .ZN(n1198) );
NAND2_X1 U999 ( .A1(G221), .A2(n1265), .ZN(n1032) );
NAND2_X1 U1000 ( .A1(n1281), .A2(n1240), .ZN(n1265) );
XOR2_X1 U1001 ( .A(G234), .B(KEYINPUT24), .Z(n1281) );
XOR2_X1 U1002 ( .A(n1071), .B(n1282), .Z(n1049) );
XOR2_X1 U1003 ( .A(KEYINPUT16), .B(G469), .Z(n1282) );
NAND2_X1 U1004 ( .A1(n1283), .A2(n1240), .ZN(n1071) );
XOR2_X1 U1005 ( .A(n1150), .B(n1284), .Z(n1283) );
NOR2_X1 U1006 ( .A1(KEYINPUT0), .A2(n1285), .ZN(n1284) );
XOR2_X1 U1007 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U1008 ( .A(n1157), .B(n1156), .Z(n1287) );
AND2_X1 U1009 ( .A1(G227), .A2(n1026), .ZN(n1156) );
NAND2_X1 U1010 ( .A1(KEYINPUT55), .A2(n1212), .ZN(n1286) );
INV_X1 U1011 ( .A(G140), .ZN(n1212) );
XOR2_X1 U1012 ( .A(n1279), .B(n1288), .Z(n1150) );
XOR2_X1 U1013 ( .A(n1206), .B(n1143), .Z(n1288) );
XOR2_X1 U1014 ( .A(n1289), .B(n1097), .Z(n1143) );
XOR2_X1 U1015 ( .A(G134), .B(G137), .Z(n1097) );
XOR2_X1 U1016 ( .A(n1290), .B(KEYINPUT34), .Z(n1289) );
XNOR2_X1 U1017 ( .A(G128), .B(n1291), .ZN(n1206) );
XNOR2_X1 U1018 ( .A(G101), .B(n1292), .ZN(n1279) );
XOR2_X1 U1019 ( .A(G107), .B(G104), .Z(n1292) );
INV_X1 U1020 ( .A(n1048), .ZN(n1036) );
NAND2_X1 U1021 ( .A1(n1211), .A2(n1210), .ZN(n1048) );
XOR2_X1 U1022 ( .A(n1293), .B(G475), .Z(n1210) );
NAND2_X1 U1023 ( .A1(n1134), .A2(n1240), .ZN(n1293) );
INV_X1 U1024 ( .A(G902), .ZN(n1240) );
XNOR2_X1 U1025 ( .A(n1294), .B(n1295), .ZN(n1134) );
XOR2_X1 U1026 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U1027 ( .A(n1298), .B(n1299), .Z(n1297) );
NOR2_X1 U1028 ( .A1(KEYINPUT3), .A2(n1300), .ZN(n1299) );
XOR2_X1 U1029 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1030 ( .A(G122), .B(G104), .Z(n1302) );
NAND2_X1 U1031 ( .A1(n1303), .A2(n1235), .ZN(n1301) );
INV_X1 U1032 ( .A(G113), .ZN(n1235) );
XNOR2_X1 U1033 ( .A(KEYINPUT63), .B(KEYINPUT60), .ZN(n1303) );
NAND3_X1 U1034 ( .A1(n1267), .A2(n1026), .A3(G214), .ZN(n1298) );
INV_X1 U1035 ( .A(G237), .ZN(n1267) );
NAND2_X1 U1036 ( .A1(KEYINPUT49), .A2(n1290), .ZN(n1296) );
INV_X1 U1037 ( .A(G131), .ZN(n1290) );
XOR2_X1 U1038 ( .A(n1257), .B(n1291), .Z(n1294) );
XOR2_X1 U1039 ( .A(G143), .B(G146), .Z(n1291) );
XOR2_X1 U1040 ( .A(n1304), .B(n1089), .Z(n1257) );
XNOR2_X1 U1041 ( .A(n1217), .B(G140), .ZN(n1089) );
INV_X1 U1042 ( .A(G125), .ZN(n1217) );
XNOR2_X1 U1043 ( .A(KEYINPUT36), .B(KEYINPUT11), .ZN(n1304) );
XOR2_X1 U1044 ( .A(n1305), .B(G478), .Z(n1211) );
OR2_X1 U1045 ( .A1(n1130), .A2(G902), .ZN(n1305) );
XNOR2_X1 U1046 ( .A(n1306), .B(n1307), .ZN(n1130) );
XOR2_X1 U1047 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U1048 ( .A(G122), .B(G116), .Z(n1309) );
XOR2_X1 U1049 ( .A(G143), .B(G134), .Z(n1308) );
XOR2_X1 U1050 ( .A(n1310), .B(n1311), .Z(n1306) );
NOR2_X1 U1051 ( .A1(G128), .A2(KEYINPUT22), .ZN(n1311) );
XOR2_X1 U1052 ( .A(n1312), .B(G107), .Z(n1310) );
NAND2_X1 U1053 ( .A1(G217), .A2(n1263), .ZN(n1312) );
AND2_X1 U1054 ( .A1(G234), .A2(n1026), .ZN(n1263) );
INV_X1 U1055 ( .A(G953), .ZN(n1026) );
INV_X1 U1056 ( .A(G110), .ZN(n1157) );
endmodule


