//Key = 1010101111100010110000110000010000100001000010100101110001000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352;

NAND2_X1 U752 ( .A1(n1041), .A2(n1042), .ZN(G9) );
OR2_X1 U753 ( .A1(n1043), .A2(G107), .ZN(n1042) );
XOR2_X1 U754 ( .A(n1044), .B(KEYINPUT1), .Z(n1041) );
NAND2_X1 U755 ( .A1(G107), .A2(n1043), .ZN(n1044) );
NAND2_X1 U756 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
XOR2_X1 U757 ( .A(n1047), .B(KEYINPUT6), .Z(n1045) );
NOR2_X1 U758 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR3_X1 U759 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
NAND3_X1 U760 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1050) );
NAND2_X1 U761 ( .A1(n1056), .A2(n1057), .ZN(n1053) );
NAND2_X1 U762 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND4_X1 U763 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1059) );
NAND2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
OR2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(n1064) );
NAND2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
OR2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
INV_X1 U770 ( .A(n1076), .ZN(n1072) );
NAND3_X1 U771 ( .A1(n1066), .A2(n1077), .A3(n1070), .ZN(n1058) );
NAND2_X1 U772 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND3_X1 U773 ( .A1(n1080), .A2(n1081), .A3(n1060), .ZN(n1079) );
NAND2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND3_X1 U775 ( .A1(n1084), .A2(n1085), .A3(n1063), .ZN(n1080) );
INV_X1 U776 ( .A(n1086), .ZN(n1085) );
NAND2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1084) );
NAND2_X1 U778 ( .A1(n1046), .A2(n1061), .ZN(n1078) );
INV_X1 U779 ( .A(n1089), .ZN(n1056) );
AND3_X1 U780 ( .A1(n1055), .A2(n1090), .A3(n1054), .ZN(n1048) );
NAND4_X1 U781 ( .A1(n1060), .A2(n1087), .A3(n1091), .A4(n1092), .ZN(n1054) );
NOR3_X1 U782 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
XNOR2_X1 U783 ( .A(G469), .B(n1096), .ZN(n1095) );
XNOR2_X1 U784 ( .A(KEYINPUT20), .B(n1074), .ZN(n1094) );
NAND3_X1 U785 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1093) );
XNOR2_X1 U786 ( .A(n1100), .B(G475), .ZN(n1099) );
OR2_X1 U787 ( .A1(n1101), .A2(KEYINPUT51), .ZN(n1098) );
NAND3_X1 U788 ( .A1(n1101), .A2(n1102), .A3(KEYINPUT51), .ZN(n1097) );
NOR3_X1 U789 ( .A1(n1103), .A2(n1104), .A3(n1082), .ZN(n1091) );
XOR2_X1 U790 ( .A(n1105), .B(KEYINPUT43), .Z(n1103) );
NAND2_X1 U791 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U792 ( .A1(G478), .A2(n1108), .ZN(n1106) );
XOR2_X1 U793 ( .A(n1109), .B(n1110), .Z(G72) );
XOR2_X1 U794 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U795 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XNOR2_X1 U796 ( .A(KEYINPUT26), .B(n1115), .ZN(n1114) );
INV_X1 U797 ( .A(n1051), .ZN(n1113) );
NAND2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1111) );
NAND2_X1 U799 ( .A1(G953), .A2(n1118), .ZN(n1117) );
XOR2_X1 U800 ( .A(n1119), .B(n1120), .Z(n1116) );
XNOR2_X1 U801 ( .A(n1121), .B(n1122), .ZN(n1120) );
XNOR2_X1 U802 ( .A(n1123), .B(n1124), .ZN(n1119) );
NAND2_X1 U803 ( .A1(G953), .A2(n1125), .ZN(n1109) );
NAND2_X1 U804 ( .A1(G900), .A2(G227), .ZN(n1125) );
XOR2_X1 U805 ( .A(n1126), .B(n1127), .Z(G69) );
XOR2_X1 U806 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XNOR2_X1 U808 ( .A(G953), .B(KEYINPUT57), .ZN(n1131) );
XNOR2_X1 U809 ( .A(n1132), .B(KEYINPUT29), .ZN(n1130) );
NAND3_X1 U810 ( .A1(n1133), .A2(n1134), .A3(KEYINPUT2), .ZN(n1128) );
NAND2_X1 U811 ( .A1(G953), .A2(n1135), .ZN(n1134) );
XOR2_X1 U812 ( .A(n1136), .B(n1137), .Z(n1133) );
NAND2_X1 U813 ( .A1(G953), .A2(n1138), .ZN(n1126) );
NAND2_X1 U814 ( .A1(G898), .A2(G224), .ZN(n1138) );
NOR2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(G66) );
XOR2_X1 U816 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U817 ( .A(KEYINPUT27), .B(n1143), .Z(n1142) );
NOR2_X1 U818 ( .A1(n1102), .A2(n1144), .ZN(n1143) );
NOR2_X1 U819 ( .A1(n1139), .A2(n1145), .ZN(G63) );
XOR2_X1 U820 ( .A(n1146), .B(n1147), .Z(n1145) );
XNOR2_X1 U821 ( .A(KEYINPUT13), .B(n1148), .ZN(n1147) );
NOR2_X1 U822 ( .A1(n1149), .A2(n1144), .ZN(n1146) );
INV_X1 U823 ( .A(G478), .ZN(n1149) );
NOR2_X1 U824 ( .A1(n1139), .A2(n1150), .ZN(G60) );
XOR2_X1 U825 ( .A(n1151), .B(n1152), .Z(n1150) );
AND2_X1 U826 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U827 ( .A1(n1155), .A2(n1144), .ZN(n1151) );
XOR2_X1 U828 ( .A(n1156), .B(n1157), .Z(G6) );
XOR2_X1 U829 ( .A(KEYINPUT38), .B(G104), .Z(n1157) );
NAND2_X1 U830 ( .A1(n1158), .A2(n1159), .ZN(n1156) );
NAND4_X1 U831 ( .A1(n1061), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1159) );
INV_X1 U832 ( .A(KEYINPUT12), .ZN(n1162) );
NAND4_X1 U833 ( .A1(n1160), .A2(n1083), .A3(n1161), .A4(KEYINPUT12), .ZN(n1158) );
NOR2_X1 U834 ( .A1(n1163), .A2(n1164), .ZN(n1161) );
INV_X1 U835 ( .A(n1061), .ZN(n1083) );
NOR2_X1 U836 ( .A1(n1139), .A2(n1165), .ZN(G57) );
XOR2_X1 U837 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U839 ( .A(n1170), .B(n1171), .Z(n1166) );
NOR2_X1 U840 ( .A1(n1172), .A2(n1144), .ZN(n1171) );
NOR2_X1 U841 ( .A1(n1139), .A2(n1173), .ZN(G54) );
XOR2_X1 U842 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U843 ( .A(n1176), .B(n1177), .ZN(n1175) );
XOR2_X1 U844 ( .A(n1178), .B(n1179), .Z(n1177) );
NOR3_X1 U845 ( .A1(n1144), .A2(KEYINPUT37), .A3(n1180), .ZN(n1178) );
XOR2_X1 U846 ( .A(n1181), .B(n1182), .Z(n1174) );
XOR2_X1 U847 ( .A(KEYINPUT62), .B(KEYINPUT40), .Z(n1182) );
XOR2_X1 U848 ( .A(n1183), .B(n1184), .Z(n1181) );
NOR2_X1 U849 ( .A1(KEYINPUT32), .A2(n1185), .ZN(n1184) );
XOR2_X1 U850 ( .A(n1186), .B(n1187), .Z(n1185) );
XNOR2_X1 U851 ( .A(G101), .B(n1188), .ZN(n1187) );
NAND2_X1 U852 ( .A1(KEYINPUT53), .A2(n1123), .ZN(n1186) );
NOR2_X1 U853 ( .A1(n1139), .A2(n1189), .ZN(G51) );
XOR2_X1 U854 ( .A(n1190), .B(n1191), .Z(n1189) );
XOR2_X1 U855 ( .A(n1192), .B(n1193), .Z(n1191) );
NOR2_X1 U856 ( .A1(n1194), .A2(n1144), .ZN(n1192) );
NAND2_X1 U857 ( .A1(G902), .A2(n1195), .ZN(n1144) );
NAND2_X1 U858 ( .A1(n1132), .A2(n1196), .ZN(n1195) );
XNOR2_X1 U859 ( .A(KEYINPUT36), .B(n1051), .ZN(n1196) );
NAND4_X1 U860 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1051) );
NOR4_X1 U861 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
AND2_X1 U862 ( .A1(n1205), .A2(n1206), .ZN(n1199) );
NAND3_X1 U863 ( .A1(n1207), .A2(n1069), .A3(n1208), .ZN(n1197) );
INV_X1 U864 ( .A(n1052), .ZN(n1132) );
NAND4_X1 U865 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1052) );
AND3_X1 U866 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1212) );
NAND2_X1 U867 ( .A1(n1046), .A2(n1216), .ZN(n1211) );
NAND3_X1 U868 ( .A1(n1217), .A2(n1047), .A3(n1218), .ZN(n1216) );
XOR2_X1 U869 ( .A(n1219), .B(KEYINPUT50), .Z(n1218) );
NAND3_X1 U870 ( .A1(n1061), .A2(n1160), .A3(n1069), .ZN(n1047) );
NAND3_X1 U871 ( .A1(n1061), .A2(n1160), .A3(n1068), .ZN(n1217) );
NAND4_X1 U872 ( .A1(n1068), .A2(n1086), .A3(n1220), .A4(n1221), .ZN(n1209) );
OR2_X1 U873 ( .A1(n1222), .A2(KEYINPUT47), .ZN(n1221) );
NAND2_X1 U874 ( .A1(KEYINPUT47), .A2(n1223), .ZN(n1220) );
NAND3_X1 U875 ( .A1(n1224), .A2(n1163), .A3(n1066), .ZN(n1223) );
XNOR2_X1 U876 ( .A(KEYINPUT18), .B(n1225), .ZN(n1190) );
NOR2_X1 U877 ( .A1(G125), .A2(KEYINPUT19), .ZN(n1225) );
AND2_X1 U878 ( .A1(n1226), .A2(n1090), .ZN(n1139) );
INV_X1 U879 ( .A(G952), .ZN(n1090) );
XNOR2_X1 U880 ( .A(G953), .B(KEYINPUT8), .ZN(n1226) );
XOR2_X1 U881 ( .A(G146), .B(n1204), .Z(G48) );
AND3_X1 U882 ( .A1(n1068), .A2(n1207), .A3(n1208), .ZN(n1204) );
XNOR2_X1 U883 ( .A(G143), .B(n1198), .ZN(G45) );
NAND4_X1 U884 ( .A1(n1208), .A2(n1086), .A3(n1227), .A4(n1228), .ZN(n1198) );
XOR2_X1 U885 ( .A(G140), .B(n1203), .Z(G42) );
AND4_X1 U886 ( .A1(n1229), .A2(n1068), .A3(n1087), .A4(n1088), .ZN(n1203) );
NAND2_X1 U887 ( .A1(n1230), .A2(n1231), .ZN(G39) );
OR2_X1 U888 ( .A1(n1206), .A2(G137), .ZN(n1231) );
XOR2_X1 U889 ( .A(n1232), .B(KEYINPUT42), .Z(n1230) );
NAND2_X1 U890 ( .A1(G137), .A2(n1206), .ZN(n1232) );
NAND3_X1 U891 ( .A1(n1207), .A2(n1070), .A3(n1229), .ZN(n1206) );
XOR2_X1 U892 ( .A(G134), .B(n1202), .Z(G36) );
AND3_X1 U893 ( .A1(n1086), .A2(n1069), .A3(n1229), .ZN(n1202) );
XOR2_X1 U894 ( .A(G131), .B(n1201), .Z(G33) );
AND3_X1 U895 ( .A1(n1068), .A2(n1086), .A3(n1229), .ZN(n1201) );
AND4_X1 U896 ( .A1(n1060), .A2(n1076), .A3(n1063), .A4(n1233), .ZN(n1229) );
XNOR2_X1 U897 ( .A(G128), .B(n1234), .ZN(G30) );
NAND3_X1 U898 ( .A1(n1069), .A2(n1235), .A3(n1208), .ZN(n1234) );
AND3_X1 U899 ( .A1(n1076), .A2(n1233), .A3(n1046), .ZN(n1208) );
XOR2_X1 U900 ( .A(KEYINPUT15), .B(n1207), .Z(n1235) );
XNOR2_X1 U901 ( .A(n1236), .B(n1237), .ZN(G3) );
NOR2_X1 U902 ( .A1(n1163), .A2(n1219), .ZN(n1237) );
NAND2_X1 U903 ( .A1(n1086), .A2(n1238), .ZN(n1219) );
XNOR2_X1 U904 ( .A(G125), .B(n1205), .ZN(G27) );
NAND4_X1 U905 ( .A1(n1068), .A2(n1239), .A3(n1066), .A4(n1233), .ZN(n1205) );
NAND2_X1 U906 ( .A1(n1240), .A2(n1089), .ZN(n1233) );
NAND4_X1 U907 ( .A1(G953), .A2(G902), .A3(n1241), .A4(n1118), .ZN(n1240) );
INV_X1 U908 ( .A(G900), .ZN(n1118) );
XOR2_X1 U909 ( .A(n1210), .B(n1242), .Z(G24) );
NOR2_X1 U910 ( .A1(KEYINPUT3), .A2(n1243), .ZN(n1242) );
XOR2_X1 U911 ( .A(KEYINPUT11), .B(G122), .Z(n1243) );
NAND4_X1 U912 ( .A1(n1222), .A2(n1061), .A3(n1227), .A4(n1228), .ZN(n1210) );
NOR2_X1 U913 ( .A1(n1088), .A2(n1244), .ZN(n1061) );
XNOR2_X1 U914 ( .A(G119), .B(n1213), .ZN(G21) );
NAND3_X1 U915 ( .A1(n1222), .A2(n1070), .A3(n1207), .ZN(n1213) );
NOR2_X1 U916 ( .A1(n1087), .A2(n1245), .ZN(n1207) );
XNOR2_X1 U917 ( .A(G116), .B(n1215), .ZN(G18) );
NAND3_X1 U918 ( .A1(n1222), .A2(n1069), .A3(n1086), .ZN(n1215) );
NOR2_X1 U919 ( .A1(n1227), .A2(n1246), .ZN(n1069) );
XNOR2_X1 U920 ( .A(G113), .B(n1247), .ZN(G15) );
NAND4_X1 U921 ( .A1(KEYINPUT46), .A2(n1068), .A3(n1086), .A4(n1222), .ZN(n1247) );
AND3_X1 U922 ( .A1(n1066), .A2(n1224), .A3(n1046), .ZN(n1222) );
NOR2_X1 U923 ( .A1(n1088), .A2(n1087), .ZN(n1086) );
INV_X1 U924 ( .A(n1244), .ZN(n1087) );
INV_X1 U925 ( .A(n1245), .ZN(n1088) );
INV_X1 U926 ( .A(n1164), .ZN(n1068) );
NAND2_X1 U927 ( .A1(n1246), .A2(n1227), .ZN(n1164) );
INV_X1 U928 ( .A(n1228), .ZN(n1246) );
XNOR2_X1 U929 ( .A(G110), .B(n1214), .ZN(G12) );
NAND2_X1 U930 ( .A1(n1239), .A2(n1238), .ZN(n1214) );
AND2_X1 U931 ( .A1(n1070), .A2(n1160), .ZN(n1238) );
AND2_X1 U932 ( .A1(n1076), .A2(n1224), .ZN(n1160) );
NAND2_X1 U933 ( .A1(n1089), .A2(n1248), .ZN(n1224) );
NAND4_X1 U934 ( .A1(G953), .A2(G902), .A3(n1241), .A4(n1135), .ZN(n1248) );
INV_X1 U935 ( .A(G898), .ZN(n1135) );
NAND3_X1 U936 ( .A1(n1055), .A2(n1241), .A3(G952), .ZN(n1089) );
NAND2_X1 U937 ( .A1(G237), .A2(G234), .ZN(n1241) );
XOR2_X1 U938 ( .A(n1115), .B(KEYINPUT54), .Z(n1055) );
NAND2_X1 U939 ( .A1(n1249), .A2(n1250), .ZN(n1076) );
NAND2_X1 U940 ( .A1(n1066), .A2(n1251), .ZN(n1250) );
INV_X1 U941 ( .A(KEYINPUT49), .ZN(n1251) );
NOR2_X1 U942 ( .A1(n1075), .A2(n1252), .ZN(n1066) );
INV_X1 U943 ( .A(n1074), .ZN(n1252) );
NAND3_X1 U944 ( .A1(n1075), .A2(n1074), .A3(KEYINPUT49), .ZN(n1249) );
NAND2_X1 U945 ( .A1(G221), .A2(n1253), .ZN(n1074) );
XNOR2_X1 U946 ( .A(n1096), .B(n1254), .ZN(n1075) );
NOR2_X1 U947 ( .A1(KEYINPUT48), .A2(n1180), .ZN(n1254) );
INV_X1 U948 ( .A(G469), .ZN(n1180) );
NAND2_X1 U949 ( .A1(n1255), .A2(n1256), .ZN(n1096) );
XOR2_X1 U950 ( .A(n1257), .B(n1258), .Z(n1255) );
XNOR2_X1 U951 ( .A(n1188), .B(n1259), .ZN(n1258) );
XOR2_X1 U952 ( .A(KEYINPUT40), .B(n1260), .Z(n1259) );
NOR2_X1 U953 ( .A1(KEYINPUT21), .A2(n1183), .ZN(n1260) );
NAND2_X1 U954 ( .A1(G227), .A2(n1115), .ZN(n1183) );
NAND2_X1 U955 ( .A1(n1261), .A2(n1262), .ZN(n1188) );
NAND2_X1 U956 ( .A1(G104), .A2(n1263), .ZN(n1262) );
XOR2_X1 U957 ( .A(KEYINPUT9), .B(n1264), .Z(n1261) );
NOR2_X1 U958 ( .A1(G104), .A2(n1263), .ZN(n1264) );
XOR2_X1 U959 ( .A(n1265), .B(n1168), .Z(n1257) );
XNOR2_X1 U960 ( .A(n1122), .B(G101), .ZN(n1168) );
XOR2_X1 U961 ( .A(n1123), .B(n1179), .Z(n1265) );
XOR2_X1 U962 ( .A(G110), .B(n1121), .Z(n1179) );
XNOR2_X1 U963 ( .A(n1266), .B(n1267), .ZN(n1123) );
XNOR2_X1 U964 ( .A(KEYINPUT39), .B(n1268), .ZN(n1267) );
NOR2_X1 U965 ( .A1(n1228), .A2(n1227), .ZN(n1070) );
NAND2_X1 U966 ( .A1(n1269), .A2(n1270), .ZN(n1227) );
NAND2_X1 U967 ( .A1(n1100), .A2(n1155), .ZN(n1270) );
XOR2_X1 U968 ( .A(KEYINPUT63), .B(n1271), .Z(n1269) );
NOR2_X1 U969 ( .A1(n1100), .A2(n1155), .ZN(n1271) );
INV_X1 U970 ( .A(G475), .ZN(n1155) );
AND2_X1 U971 ( .A1(n1256), .A2(n1272), .ZN(n1100) );
NAND2_X1 U972 ( .A1(n1153), .A2(n1154), .ZN(n1272) );
NAND2_X1 U973 ( .A1(n1273), .A2(n1274), .ZN(n1154) );
XNOR2_X1 U974 ( .A(n1275), .B(n1276), .ZN(n1274) );
XOR2_X1 U975 ( .A(KEYINPUT30), .B(n1277), .Z(n1273) );
NAND2_X1 U976 ( .A1(n1278), .A2(n1279), .ZN(n1153) );
XNOR2_X1 U977 ( .A(n1280), .B(n1276), .ZN(n1279) );
XNOR2_X1 U978 ( .A(n1281), .B(n1282), .ZN(n1276) );
NOR2_X1 U979 ( .A1(KEYINPUT59), .A2(n1124), .ZN(n1282) );
NAND2_X1 U980 ( .A1(KEYINPUT22), .A2(n1283), .ZN(n1281) );
XOR2_X1 U981 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U982 ( .A(n1286), .B(G131), .ZN(n1285) );
INV_X1 U983 ( .A(G143), .ZN(n1286) );
AND3_X1 U984 ( .A1(G214), .A2(n1115), .A3(n1287), .ZN(n1284) );
XNOR2_X1 U985 ( .A(n1277), .B(KEYINPUT25), .ZN(n1278) );
XNOR2_X1 U986 ( .A(n1288), .B(n1289), .ZN(n1277) );
XOR2_X1 U987 ( .A(KEYINPUT34), .B(G122), .Z(n1289) );
XNOR2_X1 U988 ( .A(G104), .B(n1290), .ZN(n1288) );
NOR2_X1 U989 ( .A1(KEYINPUT58), .A2(n1291), .ZN(n1290) );
NAND3_X1 U990 ( .A1(n1292), .A2(n1293), .A3(n1107), .ZN(n1228) );
OR2_X1 U991 ( .A1(n1108), .A2(G478), .ZN(n1107) );
OR2_X1 U992 ( .A1(G478), .A2(KEYINPUT16), .ZN(n1293) );
NAND3_X1 U993 ( .A1(G478), .A2(n1108), .A3(KEYINPUT16), .ZN(n1292) );
NAND2_X1 U994 ( .A1(n1256), .A2(n1148), .ZN(n1108) );
NAND2_X1 U995 ( .A1(n1294), .A2(n1295), .ZN(n1148) );
NAND4_X1 U996 ( .A1(G234), .A2(G217), .A3(n1296), .A4(n1115), .ZN(n1295) );
NAND2_X1 U997 ( .A1(n1297), .A2(n1298), .ZN(n1294) );
NAND3_X1 U998 ( .A1(G217), .A2(n1115), .A3(G234), .ZN(n1298) );
XOR2_X1 U999 ( .A(KEYINPUT23), .B(n1296), .Z(n1297) );
AND2_X1 U1000 ( .A1(n1299), .A2(n1300), .ZN(n1296) );
NAND2_X1 U1001 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U1002 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND3_X1 U1003 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(n1299) );
INV_X1 U1004 ( .A(n1301), .ZN(n1305) );
XNOR2_X1 U1005 ( .A(n1306), .B(n1307), .ZN(n1301) );
XNOR2_X1 U1006 ( .A(G134), .B(n1268), .ZN(n1307) );
NAND2_X1 U1007 ( .A1(KEYINPUT10), .A2(G143), .ZN(n1306) );
NAND2_X1 U1008 ( .A1(n1308), .A2(n1309), .ZN(n1304) );
XNOR2_X1 U1009 ( .A(KEYINPUT28), .B(n1263), .ZN(n1309) );
XNOR2_X1 U1010 ( .A(G122), .B(n1310), .ZN(n1308) );
INV_X1 U1011 ( .A(G116), .ZN(n1310) );
XNOR2_X1 U1012 ( .A(n1311), .B(KEYINPUT7), .ZN(n1303) );
NAND2_X1 U1013 ( .A1(n1312), .A2(n1263), .ZN(n1311) );
INV_X1 U1014 ( .A(G107), .ZN(n1263) );
XNOR2_X1 U1015 ( .A(G116), .B(G122), .ZN(n1312) );
NOR3_X1 U1016 ( .A1(n1244), .A2(n1245), .A3(n1163), .ZN(n1239) );
INV_X1 U1017 ( .A(n1046), .ZN(n1163) );
NOR2_X1 U1018 ( .A1(n1060), .A2(n1082), .ZN(n1046) );
INV_X1 U1019 ( .A(n1063), .ZN(n1082) );
NAND2_X1 U1020 ( .A1(n1313), .A2(n1314), .ZN(n1063) );
XOR2_X1 U1021 ( .A(KEYINPUT45), .B(G214), .Z(n1313) );
XNOR2_X1 U1022 ( .A(n1315), .B(n1194), .ZN(n1060) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1314), .ZN(n1194) );
NAND2_X1 U1024 ( .A1(n1316), .A2(n1287), .ZN(n1314) );
NAND2_X1 U1025 ( .A1(n1317), .A2(n1256), .ZN(n1315) );
XOR2_X1 U1026 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1027 ( .A(KEYINPUT44), .B(n1320), .Z(n1319) );
XOR2_X1 U1028 ( .A(KEYINPUT56), .B(KEYINPUT52), .Z(n1320) );
XNOR2_X1 U1029 ( .A(n1193), .B(G125), .ZN(n1318) );
XNOR2_X1 U1030 ( .A(n1321), .B(n1322), .ZN(n1193) );
XOR2_X1 U1031 ( .A(n1323), .B(n1324), .Z(n1322) );
NAND2_X1 U1032 ( .A1(G224), .A2(n1115), .ZN(n1324) );
NAND2_X1 U1033 ( .A1(KEYINPUT61), .A2(n1136), .ZN(n1323) );
XNOR2_X1 U1034 ( .A(n1325), .B(KEYINPUT35), .ZN(n1136) );
XOR2_X1 U1035 ( .A(n1137), .B(n1326), .Z(n1321) );
XOR2_X1 U1036 ( .A(n1327), .B(n1328), .Z(n1137) );
XNOR2_X1 U1037 ( .A(n1236), .B(n1329), .ZN(n1328) );
NOR2_X1 U1038 ( .A1(KEYINPUT55), .A2(n1330), .ZN(n1329) );
XNOR2_X1 U1039 ( .A(G104), .B(G107), .ZN(n1330) );
XNOR2_X1 U1040 ( .A(G110), .B(G122), .ZN(n1327) );
NOR2_X1 U1041 ( .A1(n1104), .A2(n1331), .ZN(n1245) );
AND2_X1 U1042 ( .A1(n1101), .A2(n1102), .ZN(n1331) );
NOR2_X1 U1043 ( .A1(n1102), .A2(n1101), .ZN(n1104) );
NOR2_X1 U1044 ( .A1(n1141), .A2(G902), .ZN(n1101) );
XOR2_X1 U1045 ( .A(n1332), .B(n1333), .Z(n1141) );
XNOR2_X1 U1046 ( .A(n1124), .B(n1334), .ZN(n1333) );
NOR2_X1 U1047 ( .A1(KEYINPUT24), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1048 ( .A(G110), .B(n1336), .Z(n1335) );
XNOR2_X1 U1049 ( .A(n1268), .B(G119), .ZN(n1336) );
INV_X1 U1050 ( .A(G125), .ZN(n1124) );
XNOR2_X1 U1051 ( .A(n1337), .B(n1275), .ZN(n1332) );
INV_X1 U1052 ( .A(n1280), .ZN(n1275) );
XOR2_X1 U1053 ( .A(n1121), .B(n1338), .Z(n1280) );
XOR2_X1 U1054 ( .A(G140), .B(KEYINPUT14), .Z(n1121) );
NAND2_X1 U1055 ( .A1(KEYINPUT0), .A2(n1339), .ZN(n1337) );
XOR2_X1 U1056 ( .A(G137), .B(n1340), .Z(n1339) );
AND3_X1 U1057 ( .A1(G221), .A2(n1115), .A3(G234), .ZN(n1340) );
NAND2_X1 U1058 ( .A1(G217), .A2(n1253), .ZN(n1102) );
NAND2_X1 U1059 ( .A1(G234), .A2(n1316), .ZN(n1253) );
XNOR2_X1 U1060 ( .A(G902), .B(KEYINPUT41), .ZN(n1316) );
XOR2_X1 U1061 ( .A(n1341), .B(n1172), .Z(n1244) );
INV_X1 U1062 ( .A(G472), .ZN(n1172) );
NAND2_X1 U1063 ( .A1(n1342), .A2(n1256), .ZN(n1341) );
INV_X1 U1064 ( .A(G902), .ZN(n1256) );
XOR2_X1 U1065 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1066 ( .A(n1170), .B(n1345), .ZN(n1344) );
NOR2_X1 U1067 ( .A1(KEYINPUT33), .A2(n1346), .ZN(n1345) );
XNOR2_X1 U1068 ( .A(n1169), .B(n1347), .ZN(n1346) );
XNOR2_X1 U1069 ( .A(KEYINPUT60), .B(n1122), .ZN(n1347) );
INV_X1 U1070 ( .A(n1176), .ZN(n1122) );
XOR2_X1 U1071 ( .A(G131), .B(n1348), .Z(n1176) );
XOR2_X1 U1072 ( .A(G137), .B(G134), .Z(n1348) );
XNOR2_X1 U1073 ( .A(n1326), .B(n1349), .ZN(n1169) );
INV_X1 U1074 ( .A(n1325), .ZN(n1349) );
XOR2_X1 U1075 ( .A(n1350), .B(n1291), .Z(n1325) );
XNOR2_X1 U1076 ( .A(G113), .B(KEYINPUT4), .ZN(n1291) );
XNOR2_X1 U1077 ( .A(G119), .B(G116), .ZN(n1350) );
XOR2_X1 U1078 ( .A(n1351), .B(n1352), .Z(n1326) );
INV_X1 U1079 ( .A(n1266), .ZN(n1352) );
XOR2_X1 U1080 ( .A(G143), .B(n1338), .Z(n1266) );
XOR2_X1 U1081 ( .A(G146), .B(KEYINPUT5), .Z(n1338) );
NAND2_X1 U1082 ( .A1(KEYINPUT17), .A2(n1268), .ZN(n1351) );
INV_X1 U1083 ( .A(G128), .ZN(n1268) );
NAND3_X1 U1084 ( .A1(n1287), .A2(n1115), .A3(G210), .ZN(n1170) );
INV_X1 U1085 ( .A(G953), .ZN(n1115) );
INV_X1 U1086 ( .A(G237), .ZN(n1287) );
XNOR2_X1 U1087 ( .A(KEYINPUT31), .B(n1236), .ZN(n1343) );
INV_X1 U1088 ( .A(G101), .ZN(n1236) );
endmodule


