//Key = 1111001011001010100001111100001001110111100100000001110111100101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
n1448;

XOR2_X1 U777 ( .A(G107), .B(n1088), .Z(G9) );
AND2_X1 U778 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(G75) );
NOR2_X1 U780 ( .A1(G952), .A2(n1093), .ZN(n1092) );
NOR3_X1 U781 ( .A1(n1094), .A2(n1093), .A3(n1095), .ZN(n1091) );
NAND2_X1 U782 ( .A1(n1096), .A2(n1097), .ZN(n1093) );
NAND4_X1 U783 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
NOR4_X1 U784 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1101) );
NAND3_X1 U785 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1102) );
NAND2_X1 U786 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U787 ( .A(KEYINPUT62), .B(G469), .Z(n1109) );
NOR3_X1 U788 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1100) );
NOR2_X1 U789 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
XOR2_X1 U790 ( .A(n1116), .B(KEYINPUT47), .Z(n1099) );
NAND2_X1 U791 ( .A1(n1114), .A2(n1115), .ZN(n1116) );
INV_X1 U792 ( .A(n1117), .ZN(n1114) );
XNOR2_X1 U793 ( .A(n1118), .B(KEYINPUT31), .ZN(n1098) );
NAND3_X1 U794 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1094) );
XOR2_X1 U795 ( .A(KEYINPUT3), .B(n1122), .Z(n1121) );
NOR2_X1 U796 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U797 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NOR2_X1 U798 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U799 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
NOR2_X1 U800 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR2_X1 U801 ( .A1(n1133), .A2(n1134), .ZN(n1129) );
NOR2_X1 U802 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NOR2_X1 U803 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U804 ( .A1(n1139), .A2(n1140), .ZN(n1135) );
NOR3_X1 U805 ( .A1(n1141), .A2(n1132), .A3(n1134), .ZN(n1125) );
NAND3_X1 U806 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1120) );
NAND2_X1 U807 ( .A1(n1145), .A2(n1146), .ZN(n1143) );
OR3_X1 U808 ( .A1(n1147), .A2(n1106), .A3(n1132), .ZN(n1146) );
INV_X1 U809 ( .A(n1148), .ZN(n1132) );
NAND2_X1 U810 ( .A1(n1149), .A2(n1150), .ZN(n1145) );
NAND2_X1 U811 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NAND3_X1 U812 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1152) );
NAND2_X1 U813 ( .A1(n1156), .A2(n1157), .ZN(n1151) );
NAND4_X1 U814 ( .A1(n1144), .A2(n1149), .A3(n1148), .A4(n1090), .ZN(n1119) );
INV_X1 U815 ( .A(n1124), .ZN(n1144) );
XOR2_X1 U816 ( .A(n1158), .B(n1159), .Z(G72) );
XOR2_X1 U817 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U818 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U819 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U820 ( .A(n1166), .B(n1167), .Z(n1165) );
XNOR2_X1 U821 ( .A(n1168), .B(n1169), .ZN(n1166) );
XNOR2_X1 U822 ( .A(G131), .B(n1170), .ZN(n1164) );
XOR2_X1 U823 ( .A(KEYINPUT12), .B(G137), .Z(n1170) );
NOR2_X1 U824 ( .A1(G900), .A2(n1096), .ZN(n1162) );
NOR2_X1 U825 ( .A1(n1171), .A2(G953), .ZN(n1160) );
NOR2_X1 U826 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XNOR2_X1 U827 ( .A(KEYINPUT11), .B(n1174), .ZN(n1173) );
NOR2_X1 U828 ( .A1(n1175), .A2(n1096), .ZN(n1158) );
NOR2_X1 U829 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U830 ( .A(n1178), .B(n1179), .Z(G69) );
NAND2_X1 U831 ( .A1(n1096), .A2(n1180), .ZN(n1179) );
NAND2_X1 U832 ( .A1(n1181), .A2(n1182), .ZN(n1178) );
NAND3_X1 U833 ( .A1(n1183), .A2(n1184), .A3(G898), .ZN(n1182) );
NAND2_X1 U834 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND2_X1 U835 ( .A1(G953), .A2(n1187), .ZN(n1185) );
NAND2_X1 U836 ( .A1(G224), .A2(n1187), .ZN(n1183) );
OR2_X1 U837 ( .A1(n1187), .A2(G953), .ZN(n1181) );
XNOR2_X1 U838 ( .A(n1188), .B(KEYINPUT50), .ZN(n1187) );
NAND2_X1 U839 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U840 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U841 ( .A(n1193), .B(KEYINPUT46), .Z(n1189) );
NAND2_X1 U842 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
INV_X1 U843 ( .A(n1191), .ZN(n1195) );
XNOR2_X1 U844 ( .A(n1196), .B(n1197), .ZN(n1191) );
XNOR2_X1 U845 ( .A(G122), .B(KEYINPUT58), .ZN(n1196) );
XNOR2_X1 U846 ( .A(n1192), .B(KEYINPUT26), .ZN(n1194) );
XOR2_X1 U847 ( .A(n1198), .B(n1199), .Z(n1192) );
NOR2_X1 U848 ( .A1(KEYINPUT10), .A2(n1200), .ZN(n1199) );
XNOR2_X1 U849 ( .A(n1201), .B(n1202), .ZN(n1200) );
NOR2_X1 U850 ( .A1(n1203), .A2(n1204), .ZN(G66) );
XNOR2_X1 U851 ( .A(n1205), .B(n1206), .ZN(n1204) );
NAND2_X1 U852 ( .A1(n1207), .A2(n1208), .ZN(n1205) );
XNOR2_X1 U853 ( .A(G217), .B(KEYINPUT40), .ZN(n1207) );
NOR2_X1 U854 ( .A1(n1209), .A2(n1210), .ZN(G63) );
XNOR2_X1 U855 ( .A(n1211), .B(n1212), .ZN(n1210) );
XNOR2_X1 U856 ( .A(KEYINPUT22), .B(n1213), .ZN(n1211) );
NOR3_X1 U857 ( .A1(n1214), .A2(KEYINPUT49), .A3(n1215), .ZN(n1213) );
NOR2_X1 U858 ( .A1(n1216), .A2(n1217), .ZN(n1209) );
XNOR2_X1 U859 ( .A(G953), .B(KEYINPUT44), .ZN(n1217) );
XNOR2_X1 U860 ( .A(KEYINPUT21), .B(G952), .ZN(n1216) );
NOR2_X1 U861 ( .A1(n1203), .A2(n1218), .ZN(G60) );
NOR2_X1 U862 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
XOR2_X1 U863 ( .A(KEYINPUT7), .B(n1221), .Z(n1220) );
NOR2_X1 U864 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
AND2_X1 U865 ( .A1(n1223), .A2(n1222), .ZN(n1219) );
NAND2_X1 U866 ( .A1(n1208), .A2(G475), .ZN(n1223) );
XNOR2_X1 U867 ( .A(G104), .B(n1224), .ZN(G6) );
NOR2_X1 U868 ( .A1(n1203), .A2(n1225), .ZN(G57) );
NOR2_X1 U869 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
XOR2_X1 U870 ( .A(KEYINPUT17), .B(n1228), .Z(n1227) );
NOR2_X1 U871 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
AND2_X1 U872 ( .A1(n1230), .A2(n1229), .ZN(n1226) );
INV_X1 U873 ( .A(n1231), .ZN(n1229) );
XNOR2_X1 U874 ( .A(n1232), .B(n1233), .ZN(n1230) );
NOR3_X1 U875 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
NAND3_X1 U876 ( .A1(n1208), .A2(G472), .A3(KEYINPUT35), .ZN(n1232) );
NOR2_X1 U877 ( .A1(n1203), .A2(n1237), .ZN(G54) );
XOR2_X1 U878 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U879 ( .A(n1240), .B(n1241), .Z(n1239) );
NAND2_X1 U880 ( .A1(n1208), .A2(G469), .ZN(n1240) );
INV_X1 U881 ( .A(n1214), .ZN(n1208) );
NOR2_X1 U882 ( .A1(n1242), .A2(n1243), .ZN(n1238) );
NOR2_X1 U883 ( .A1(KEYINPUT29), .A2(n1244), .ZN(n1243) );
AND2_X1 U884 ( .A1(KEYINPUT48), .A2(n1244), .ZN(n1242) );
NOR2_X1 U885 ( .A1(n1203), .A2(n1245), .ZN(G51) );
XOR2_X1 U886 ( .A(n1246), .B(n1247), .Z(n1245) );
OR2_X1 U887 ( .A1(n1214), .A2(n1115), .ZN(n1247) );
NAND2_X1 U888 ( .A1(G902), .A2(n1095), .ZN(n1214) );
OR3_X1 U889 ( .A1(n1180), .A2(n1248), .A3(n1172), .ZN(n1095) );
NAND4_X1 U890 ( .A1(n1249), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1172) );
NOR3_X1 U891 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1252) );
NOR3_X1 U892 ( .A1(n1256), .A2(n1134), .A3(n1128), .ZN(n1255) );
NAND3_X1 U893 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1256) );
NAND2_X1 U894 ( .A1(KEYINPUT51), .A2(n1260), .ZN(n1258) );
NAND2_X1 U895 ( .A1(n1261), .A2(n1262), .ZN(n1257) );
INV_X1 U896 ( .A(KEYINPUT51), .ZN(n1262) );
NAND2_X1 U897 ( .A1(n1263), .A2(n1139), .ZN(n1261) );
NOR2_X1 U898 ( .A1(n1264), .A2(n1131), .ZN(n1254) );
NOR2_X1 U899 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NOR2_X1 U900 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NOR3_X1 U901 ( .A1(n1260), .A2(n1269), .A3(n1270), .ZN(n1265) );
XNOR2_X1 U902 ( .A(n1259), .B(KEYINPUT5), .ZN(n1269) );
NAND3_X1 U903 ( .A1(n1156), .A2(n1271), .A3(n1272), .ZN(n1251) );
XNOR2_X1 U904 ( .A(KEYINPUT15), .B(n1134), .ZN(n1271) );
NAND4_X1 U905 ( .A1(n1273), .A2(n1224), .A3(n1274), .A4(n1275), .ZN(n1180) );
NAND2_X1 U906 ( .A1(n1276), .A2(n1089), .ZN(n1224) );
NOR3_X1 U907 ( .A1(n1140), .A2(n1139), .A3(n1277), .ZN(n1089) );
NAND2_X1 U908 ( .A1(n1278), .A2(n1279), .ZN(n1273) );
NAND2_X1 U909 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U910 ( .A1(n1090), .A2(n1282), .ZN(n1281) );
NAND2_X1 U911 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NAND2_X1 U912 ( .A1(n1154), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U913 ( .A(KEYINPUT32), .B(n1139), .ZN(n1285) );
NAND2_X1 U914 ( .A1(n1286), .A2(n1157), .ZN(n1283) );
NAND2_X1 U915 ( .A1(n1142), .A2(n1287), .ZN(n1280) );
NAND2_X1 U916 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U917 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NAND2_X1 U918 ( .A1(n1292), .A2(n1138), .ZN(n1291) );
NAND2_X1 U919 ( .A1(n1259), .A2(n1157), .ZN(n1288) );
NAND2_X1 U920 ( .A1(n1293), .A2(n1294), .ZN(n1246) );
NAND2_X1 U921 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
XOR2_X1 U922 ( .A(KEYINPUT0), .B(n1297), .Z(n1293) );
NOR2_X1 U923 ( .A1(n1296), .A2(n1295), .ZN(n1297) );
XOR2_X1 U924 ( .A(n1298), .B(n1299), .Z(n1295) );
XOR2_X1 U925 ( .A(n1300), .B(n1301), .Z(n1299) );
NOR2_X1 U926 ( .A1(G125), .A2(KEYINPUT13), .ZN(n1301) );
AND2_X1 U927 ( .A1(G953), .A2(n1302), .ZN(n1203) );
XOR2_X1 U928 ( .A(KEYINPUT21), .B(G952), .Z(n1302) );
XNOR2_X1 U929 ( .A(n1303), .B(n1304), .ZN(G48) );
NOR3_X1 U930 ( .A1(n1268), .A2(n1305), .A3(n1267), .ZN(n1304) );
XNOR2_X1 U931 ( .A(n1306), .B(KEYINPUT19), .ZN(n1305) );
XNOR2_X1 U932 ( .A(G143), .B(n1249), .ZN(G45) );
NAND3_X1 U933 ( .A1(n1286), .A2(n1307), .A3(n1308), .ZN(n1249) );
NOR3_X1 U934 ( .A1(n1131), .A2(n1309), .A3(n1310), .ZN(n1308) );
XOR2_X1 U935 ( .A(n1311), .B(n1312), .Z(G42) );
XNOR2_X1 U936 ( .A(G140), .B(KEYINPUT60), .ZN(n1312) );
NAND2_X1 U937 ( .A1(n1313), .A2(n1156), .ZN(n1311) );
XOR2_X1 U938 ( .A(G137), .B(n1314), .Z(G39) );
NOR3_X1 U939 ( .A1(n1315), .A2(n1134), .A3(n1128), .ZN(n1314) );
XNOR2_X1 U940 ( .A(G134), .B(n1250), .ZN(G36) );
NAND4_X1 U941 ( .A1(n1286), .A2(n1307), .A3(n1149), .A4(n1090), .ZN(n1250) );
INV_X1 U942 ( .A(n1134), .ZN(n1149) );
XOR2_X1 U943 ( .A(G131), .B(n1253), .Z(G33) );
AND2_X1 U944 ( .A1(n1286), .A2(n1313), .ZN(n1253) );
NOR2_X1 U945 ( .A1(n1268), .A2(n1134), .ZN(n1313) );
NAND2_X1 U946 ( .A1(n1316), .A2(n1106), .ZN(n1134) );
INV_X1 U947 ( .A(n1272), .ZN(n1268) );
NOR2_X1 U948 ( .A1(n1141), .A2(n1260), .ZN(n1272) );
XOR2_X1 U949 ( .A(G128), .B(n1317), .Z(G30) );
NOR3_X1 U950 ( .A1(n1315), .A2(n1131), .A3(n1270), .ZN(n1317) );
INV_X1 U951 ( .A(n1090), .ZN(n1270) );
NAND2_X1 U952 ( .A1(n1307), .A2(n1259), .ZN(n1315) );
INV_X1 U953 ( .A(n1260), .ZN(n1307) );
NAND2_X1 U954 ( .A1(n1290), .A2(n1263), .ZN(n1260) );
XOR2_X1 U955 ( .A(n1318), .B(n1319), .Z(G3) );
XOR2_X1 U956 ( .A(KEYINPUT30), .B(G101), .Z(n1319) );
NAND3_X1 U957 ( .A1(n1320), .A2(n1142), .A3(n1321), .ZN(n1318) );
XNOR2_X1 U958 ( .A(n1290), .B(KEYINPUT43), .ZN(n1321) );
XNOR2_X1 U959 ( .A(n1248), .B(n1322), .ZN(G27) );
NOR2_X1 U960 ( .A1(G125), .A2(KEYINPUT54), .ZN(n1322) );
INV_X1 U961 ( .A(n1174), .ZN(n1248) );
NAND4_X1 U962 ( .A1(n1306), .A2(n1263), .A3(n1157), .A4(n1323), .ZN(n1174) );
NOR2_X1 U963 ( .A1(n1292), .A2(n1141), .ZN(n1323) );
INV_X1 U964 ( .A(n1276), .ZN(n1141) );
NAND2_X1 U965 ( .A1(n1124), .A2(n1324), .ZN(n1263) );
NAND4_X1 U966 ( .A1(G953), .A2(G902), .A3(n1325), .A4(n1177), .ZN(n1324) );
INV_X1 U967 ( .A(G900), .ZN(n1177) );
NAND2_X1 U968 ( .A1(n1326), .A2(n1327), .ZN(G24) );
NAND2_X1 U969 ( .A1(G122), .A2(n1274), .ZN(n1327) );
XOR2_X1 U970 ( .A(KEYINPUT6), .B(n1328), .Z(n1326) );
NOR2_X1 U971 ( .A1(G122), .A2(n1274), .ZN(n1328) );
NAND4_X1 U972 ( .A1(n1148), .A2(n1278), .A3(n1113), .A4(n1329), .ZN(n1274) );
NOR2_X1 U973 ( .A1(n1137), .A2(n1140), .ZN(n1148) );
INV_X1 U974 ( .A(n1154), .ZN(n1140) );
NOR2_X1 U975 ( .A1(n1111), .A2(n1118), .ZN(n1154) );
NAND2_X1 U976 ( .A1(n1330), .A2(n1331), .ZN(G21) );
NAND2_X1 U977 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
XOR2_X1 U978 ( .A(KEYINPUT25), .B(n1334), .Z(n1330) );
NOR2_X1 U979 ( .A1(n1332), .A2(n1333), .ZN(n1334) );
INV_X1 U980 ( .A(G119), .ZN(n1333) );
AND4_X1 U981 ( .A1(n1142), .A2(n1157), .A3(n1278), .A4(n1335), .ZN(n1332) );
XNOR2_X1 U982 ( .A(KEYINPUT27), .B(n1267), .ZN(n1335) );
INV_X1 U983 ( .A(n1259), .ZN(n1267) );
NOR2_X1 U984 ( .A1(n1336), .A2(n1337), .ZN(n1259) );
INV_X1 U985 ( .A(n1277), .ZN(n1278) );
XNOR2_X1 U986 ( .A(G116), .B(n1338), .ZN(G18) );
NAND3_X1 U987 ( .A1(n1320), .A2(n1157), .A3(n1339), .ZN(n1338) );
XNOR2_X1 U988 ( .A(n1090), .B(KEYINPUT23), .ZN(n1339) );
NOR2_X1 U989 ( .A1(n1113), .A2(n1309), .ZN(n1090) );
XOR2_X1 U990 ( .A(n1275), .B(n1340), .Z(G15) );
NAND2_X1 U991 ( .A1(n1341), .A2(KEYINPUT33), .ZN(n1340) );
XNOR2_X1 U992 ( .A(G113), .B(KEYINPUT34), .ZN(n1341) );
NAND3_X1 U993 ( .A1(n1276), .A2(n1157), .A3(n1320), .ZN(n1275) );
NOR2_X1 U994 ( .A1(n1138), .A2(n1277), .ZN(n1320) );
INV_X1 U995 ( .A(n1286), .ZN(n1138) );
NOR2_X1 U996 ( .A1(n1111), .A2(n1336), .ZN(n1286) );
INV_X1 U997 ( .A(n1118), .ZN(n1336) );
INV_X1 U998 ( .A(n1137), .ZN(n1157) );
NAND2_X1 U999 ( .A1(n1153), .A2(n1107), .ZN(n1137) );
NOR2_X1 U1000 ( .A1(n1329), .A2(n1310), .ZN(n1276) );
INV_X1 U1001 ( .A(n1309), .ZN(n1329) );
NAND2_X1 U1002 ( .A1(n1342), .A2(n1343), .ZN(G12) );
OR2_X1 U1003 ( .A1(n1344), .A2(G110), .ZN(n1343) );
NAND2_X1 U1004 ( .A1(G110), .A2(n1345), .ZN(n1342) );
NAND2_X1 U1005 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
NAND2_X1 U1006 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
INV_X1 U1007 ( .A(KEYINPUT39), .ZN(n1349) );
NAND2_X1 U1008 ( .A1(KEYINPUT39), .A2(n1344), .ZN(n1346) );
NAND2_X1 U1009 ( .A1(KEYINPUT8), .A2(n1348), .ZN(n1344) );
AND4_X1 U1010 ( .A1(n1350), .A2(n1351), .A3(n1142), .A4(n1352), .ZN(n1348) );
NOR2_X1 U1011 ( .A1(n1139), .A2(n1292), .ZN(n1352) );
INV_X1 U1012 ( .A(n1156), .ZN(n1292) );
NOR2_X1 U1013 ( .A1(n1118), .A2(n1337), .ZN(n1156) );
INV_X1 U1014 ( .A(n1111), .ZN(n1337) );
NAND3_X1 U1015 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1111) );
NAND2_X1 U1016 ( .A1(n1356), .A2(n1206), .ZN(n1355) );
OR3_X1 U1017 ( .A1(n1206), .A2(n1356), .A3(G902), .ZN(n1354) );
NOR2_X1 U1018 ( .A1(n1357), .A2(G234), .ZN(n1356) );
INV_X1 U1019 ( .A(G217), .ZN(n1357) );
XOR2_X1 U1020 ( .A(n1358), .B(n1359), .Z(n1206) );
XOR2_X1 U1021 ( .A(n1360), .B(n1361), .Z(n1359) );
XNOR2_X1 U1022 ( .A(G119), .B(G137), .ZN(n1361) );
NAND2_X1 U1023 ( .A1(KEYINPUT55), .A2(n1362), .ZN(n1360) );
XOR2_X1 U1024 ( .A(n1363), .B(n1364), .Z(n1358) );
XOR2_X1 U1025 ( .A(n1365), .B(n1366), .Z(n1364) );
NAND3_X1 U1026 ( .A1(n1367), .A2(n1096), .A3(G221), .ZN(n1365) );
NAND2_X1 U1027 ( .A1(G902), .A2(G217), .ZN(n1353) );
XNOR2_X1 U1028 ( .A(n1368), .B(G472), .ZN(n1118) );
NAND2_X1 U1029 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
XOR2_X1 U1030 ( .A(n1371), .B(n1372), .Z(n1370) );
NAND2_X1 U1031 ( .A1(KEYINPUT14), .A2(n1231), .ZN(n1372) );
XNOR2_X1 U1032 ( .A(n1373), .B(G101), .ZN(n1231) );
NAND2_X1 U1033 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
XNOR2_X1 U1034 ( .A(G210), .B(KEYINPUT16), .ZN(n1374) );
NAND3_X1 U1035 ( .A1(n1376), .A2(n1377), .A3(n1378), .ZN(n1371) );
INV_X1 U1036 ( .A(n1236), .ZN(n1378) );
NOR3_X1 U1037 ( .A1(n1298), .A2(n1379), .A3(n1380), .ZN(n1236) );
NAND2_X1 U1038 ( .A1(n1381), .A2(n1382), .ZN(n1377) );
INV_X1 U1039 ( .A(KEYINPUT41), .ZN(n1382) );
OR2_X1 U1040 ( .A1(n1235), .A2(n1234), .ZN(n1381) );
NOR3_X1 U1041 ( .A1(n1198), .A2(n1383), .A3(n1298), .ZN(n1234) );
AND2_X1 U1042 ( .A1(n1384), .A2(n1298), .ZN(n1235) );
XNOR2_X1 U1043 ( .A(n1198), .B(n1380), .ZN(n1384) );
NAND2_X1 U1044 ( .A1(n1385), .A2(KEYINPUT41), .ZN(n1376) );
XNOR2_X1 U1045 ( .A(n1386), .B(n1198), .ZN(n1385) );
NAND2_X1 U1046 ( .A1(n1298), .A2(n1380), .ZN(n1386) );
XNOR2_X1 U1047 ( .A(G902), .B(KEYINPUT28), .ZN(n1369) );
INV_X1 U1048 ( .A(n1290), .ZN(n1139) );
NOR2_X1 U1049 ( .A1(n1155), .A2(n1153), .ZN(n1290) );
NOR2_X1 U1050 ( .A1(n1387), .A2(n1103), .ZN(n1153) );
NOR2_X1 U1051 ( .A1(n1110), .A2(G469), .ZN(n1103) );
AND2_X1 U1052 ( .A1(n1388), .A2(n1110), .ZN(n1387) );
NAND2_X1 U1053 ( .A1(n1389), .A2(n1390), .ZN(n1110) );
XOR2_X1 U1054 ( .A(n1241), .B(n1244), .Z(n1389) );
XNOR2_X1 U1055 ( .A(n1391), .B(n1202), .ZN(n1244) );
XNOR2_X1 U1056 ( .A(n1392), .B(n1393), .ZN(n1391) );
INV_X1 U1057 ( .A(n1168), .ZN(n1393) );
XOR2_X1 U1058 ( .A(G146), .B(n1394), .Z(n1168) );
NAND2_X1 U1059 ( .A1(KEYINPUT9), .A2(n1201), .ZN(n1392) );
INV_X1 U1060 ( .A(G104), .ZN(n1201) );
XOR2_X1 U1061 ( .A(n1395), .B(n1396), .Z(n1241) );
XNOR2_X1 U1062 ( .A(n1383), .B(n1397), .ZN(n1396) );
INV_X1 U1063 ( .A(n1380), .ZN(n1383) );
XNOR2_X1 U1064 ( .A(n1398), .B(G131), .ZN(n1380) );
NAND2_X1 U1065 ( .A1(n1399), .A2(n1400), .ZN(n1398) );
NAND2_X1 U1066 ( .A1(G137), .A2(n1401), .ZN(n1400) );
XOR2_X1 U1067 ( .A(n1402), .B(KEYINPUT42), .Z(n1399) );
OR2_X1 U1068 ( .A1(n1401), .A2(G137), .ZN(n1402) );
XNOR2_X1 U1069 ( .A(G110), .B(n1403), .ZN(n1395) );
NOR2_X1 U1070 ( .A1(G953), .A2(n1176), .ZN(n1403) );
INV_X1 U1071 ( .A(G227), .ZN(n1176) );
XNOR2_X1 U1072 ( .A(G469), .B(KEYINPUT37), .ZN(n1388) );
INV_X1 U1073 ( .A(n1107), .ZN(n1155) );
NAND2_X1 U1074 ( .A1(G221), .A2(n1404), .ZN(n1107) );
NAND2_X1 U1075 ( .A1(G234), .A2(n1390), .ZN(n1404) );
INV_X1 U1076 ( .A(n1128), .ZN(n1142) );
NAND2_X1 U1077 ( .A1(n1309), .A2(n1405), .ZN(n1128) );
XNOR2_X1 U1078 ( .A(KEYINPUT57), .B(n1310), .ZN(n1405) );
INV_X1 U1079 ( .A(n1113), .ZN(n1310) );
XNOR2_X1 U1080 ( .A(n1406), .B(G475), .ZN(n1113) );
NAND2_X1 U1081 ( .A1(n1222), .A2(n1390), .ZN(n1406) );
XNOR2_X1 U1082 ( .A(n1407), .B(n1408), .ZN(n1222) );
XOR2_X1 U1083 ( .A(n1409), .B(n1410), .Z(n1408) );
XOR2_X1 U1084 ( .A(n1411), .B(G131), .Z(n1410) );
NAND2_X1 U1085 ( .A1(G214), .A2(n1375), .ZN(n1411) );
NOR2_X1 U1086 ( .A1(G953), .A2(G237), .ZN(n1375) );
XNOR2_X1 U1087 ( .A(G143), .B(KEYINPUT2), .ZN(n1409) );
XOR2_X1 U1088 ( .A(n1412), .B(n1413), .Z(n1407) );
XOR2_X1 U1089 ( .A(n1363), .B(n1414), .Z(n1412) );
XNOR2_X1 U1090 ( .A(n1167), .B(G146), .ZN(n1363) );
XOR2_X1 U1091 ( .A(G125), .B(n1397), .Z(n1167) );
XOR2_X1 U1092 ( .A(G140), .B(KEYINPUT36), .Z(n1397) );
NOR2_X1 U1093 ( .A1(n1415), .A2(n1105), .ZN(n1309) );
AND3_X1 U1094 ( .A1(n1215), .A2(n1390), .A3(n1212), .ZN(n1105) );
INV_X1 U1095 ( .A(G478), .ZN(n1215) );
XOR2_X1 U1096 ( .A(n1104), .B(KEYINPUT4), .Z(n1415) );
AND2_X1 U1097 ( .A1(G478), .A2(n1416), .ZN(n1104) );
NAND2_X1 U1098 ( .A1(n1212), .A2(n1390), .ZN(n1416) );
XOR2_X1 U1099 ( .A(n1417), .B(n1418), .Z(n1212) );
XOR2_X1 U1100 ( .A(G107), .B(n1419), .Z(n1418) );
XNOR2_X1 U1101 ( .A(n1420), .B(G116), .ZN(n1419) );
XNOR2_X1 U1102 ( .A(n1421), .B(n1401), .ZN(n1417) );
INV_X1 U1103 ( .A(n1169), .ZN(n1401) );
XOR2_X1 U1104 ( .A(G134), .B(KEYINPUT18), .Z(n1169) );
XOR2_X1 U1105 ( .A(n1422), .B(n1423), .Z(n1421) );
AND3_X1 U1106 ( .A1(G217), .A2(n1096), .A3(n1367), .ZN(n1423) );
XNOR2_X1 U1107 ( .A(G234), .B(KEYINPUT38), .ZN(n1367) );
NAND2_X1 U1108 ( .A1(n1424), .A2(n1425), .ZN(n1422) );
NAND2_X1 U1109 ( .A1(n1366), .A2(n1426), .ZN(n1425) );
XOR2_X1 U1110 ( .A(n1427), .B(KEYINPUT45), .Z(n1424) );
OR2_X1 U1111 ( .A1(n1426), .A2(n1366), .ZN(n1427) );
INV_X1 U1112 ( .A(G143), .ZN(n1426) );
NAND2_X1 U1113 ( .A1(KEYINPUT63), .A2(n1277), .ZN(n1351) );
NAND2_X1 U1114 ( .A1(n1306), .A2(n1428), .ZN(n1277) );
INV_X1 U1115 ( .A(n1131), .ZN(n1306) );
NAND2_X1 U1116 ( .A1(n1429), .A2(n1430), .ZN(n1350) );
INV_X1 U1117 ( .A(KEYINPUT63), .ZN(n1430) );
NAND2_X1 U1118 ( .A1(n1131), .A2(n1428), .ZN(n1429) );
NAND2_X1 U1119 ( .A1(n1431), .A2(n1124), .ZN(n1428) );
NAND3_X1 U1120 ( .A1(n1325), .A2(n1096), .A3(G952), .ZN(n1124) );
INV_X1 U1121 ( .A(G953), .ZN(n1096) );
NAND4_X1 U1122 ( .A1(G953), .A2(G902), .A3(n1325), .A4(n1432), .ZN(n1431) );
INV_X1 U1123 ( .A(G898), .ZN(n1432) );
NAND2_X1 U1124 ( .A1(G237), .A2(G234), .ZN(n1325) );
NAND2_X1 U1125 ( .A1(n1147), .A2(n1106), .ZN(n1131) );
NAND2_X1 U1126 ( .A1(G214), .A2(n1433), .ZN(n1106) );
INV_X1 U1127 ( .A(n1316), .ZN(n1147) );
XOR2_X1 U1128 ( .A(n1115), .B(n1434), .Z(n1316) );
NOR2_X1 U1129 ( .A1(KEYINPUT20), .A2(n1117), .ZN(n1434) );
NAND3_X1 U1130 ( .A1(n1435), .A2(n1390), .A3(n1436), .ZN(n1117) );
XOR2_X1 U1131 ( .A(KEYINPUT24), .B(n1437), .Z(n1436) );
NOR2_X1 U1132 ( .A1(n1438), .A2(n1296), .ZN(n1437) );
NAND2_X1 U1133 ( .A1(n1438), .A2(n1296), .ZN(n1435) );
XNOR2_X1 U1134 ( .A(n1439), .B(n1440), .ZN(n1296) );
XNOR2_X1 U1135 ( .A(n1202), .B(n1379), .ZN(n1440) );
INV_X1 U1136 ( .A(n1198), .ZN(n1379) );
XNOR2_X1 U1137 ( .A(n1441), .B(n1414), .ZN(n1198) );
XOR2_X1 U1138 ( .A(G113), .B(KEYINPUT53), .Z(n1414) );
XNOR2_X1 U1139 ( .A(G116), .B(G119), .ZN(n1441) );
XOR2_X1 U1140 ( .A(G101), .B(G107), .Z(n1202) );
XNOR2_X1 U1141 ( .A(n1413), .B(n1197), .ZN(n1439) );
XNOR2_X1 U1142 ( .A(n1362), .B(KEYINPUT59), .ZN(n1197) );
INV_X1 U1143 ( .A(G110), .ZN(n1362) );
XNOR2_X1 U1144 ( .A(G104), .B(n1420), .ZN(n1413) );
INV_X1 U1145 ( .A(G122), .ZN(n1420) );
XOR2_X1 U1146 ( .A(n1298), .B(n1442), .Z(n1438) );
XOR2_X1 U1147 ( .A(n1443), .B(n1444), .Z(n1442) );
NAND2_X1 U1148 ( .A1(KEYINPUT1), .A2(n1300), .ZN(n1444) );
NOR2_X1 U1149 ( .A1(n1186), .A2(G953), .ZN(n1300) );
INV_X1 U1150 ( .A(G224), .ZN(n1186) );
NAND2_X1 U1151 ( .A1(KEYINPUT52), .A2(G125), .ZN(n1443) );
NAND2_X1 U1152 ( .A1(n1445), .A2(n1446), .ZN(n1298) );
OR2_X1 U1153 ( .A1(n1303), .A2(n1394), .ZN(n1446) );
NAND2_X1 U1154 ( .A1(n1447), .A2(n1303), .ZN(n1445) );
INV_X1 U1155 ( .A(G146), .ZN(n1303) );
XNOR2_X1 U1156 ( .A(n1394), .B(KEYINPUT61), .ZN(n1447) );
XNOR2_X1 U1157 ( .A(G143), .B(n1366), .ZN(n1394) );
XNOR2_X1 U1158 ( .A(G128), .B(KEYINPUT56), .ZN(n1366) );
NAND2_X1 U1159 ( .A1(G210), .A2(n1433), .ZN(n1115) );
NAND2_X1 U1160 ( .A1(n1448), .A2(n1390), .ZN(n1433) );
INV_X1 U1161 ( .A(G902), .ZN(n1390) );
INV_X1 U1162 ( .A(G237), .ZN(n1448) );
endmodule


