//Key = 1000100011101001111010111010001110001110100011001001011110010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374;

XNOR2_X1 U774 ( .A(G107), .B(n1050), .ZN(G9) );
NAND3_X1 U775 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1050) );
NOR2_X1 U776 ( .A1(n1054), .A2(n1055), .ZN(G75) );
NOR4_X1 U777 ( .A1(n1056), .A2(n1057), .A3(G953), .A4(n1058), .ZN(n1055) );
NOR2_X1 U778 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U779 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR3_X1 U780 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
NOR2_X1 U781 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U782 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U783 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U784 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U785 ( .A(KEYINPUT17), .B(n1074), .Z(n1073) );
NOR2_X1 U786 ( .A1(n1075), .A2(n1076), .ZN(n1066) );
XNOR2_X1 U787 ( .A(KEYINPUT50), .B(n1077), .ZN(n1075) );
NOR3_X1 U788 ( .A1(n1069), .A2(n1078), .A3(n1079), .ZN(n1061) );
NOR2_X1 U789 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR2_X1 U790 ( .A1(n1082), .A2(n1063), .ZN(n1081) );
NOR2_X1 U791 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U792 ( .A1(n1085), .A2(n1065), .ZN(n1080) );
NOR2_X1 U793 ( .A1(n1053), .A2(n1086), .ZN(n1085) );
NAND3_X1 U794 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1056) );
XOR2_X1 U795 ( .A(n1090), .B(KEYINPUT57), .Z(n1089) );
NAND4_X1 U796 ( .A1(n1077), .A2(n1091), .A3(n1051), .A4(n1092), .ZN(n1090) );
NOR3_X1 U797 ( .A1(n1093), .A2(n1063), .A3(n1060), .ZN(n1092) );
NOR3_X1 U798 ( .A1(n1058), .A2(G953), .A3(G952), .ZN(n1054) );
AND4_X1 U799 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1058) );
NOR4_X1 U800 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
XOR2_X1 U801 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U802 ( .A1(G475), .A2(KEYINPUT46), .ZN(n1103) );
XNOR2_X1 U803 ( .A(n1104), .B(n1105), .ZN(n1100) );
NAND2_X1 U804 ( .A1(KEYINPUT18), .A2(n1106), .ZN(n1104) );
INV_X1 U805 ( .A(G469), .ZN(n1106) );
NOR2_X1 U806 ( .A1(n1107), .A2(n1108), .ZN(n1096) );
XOR2_X1 U807 ( .A(n1109), .B(n1110), .Z(n1094) );
NOR2_X1 U808 ( .A1(KEYINPUT13), .A2(n1111), .ZN(n1110) );
XOR2_X1 U809 ( .A(n1112), .B(n1113), .Z(G72) );
NOR2_X1 U810 ( .A1(KEYINPUT33), .A2(n1114), .ZN(n1113) );
XOR2_X1 U811 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U812 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U813 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U814 ( .A(n1121), .B(n1122), .Z(n1120) );
NAND2_X1 U815 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
INV_X1 U816 ( .A(n1125), .ZN(n1124) );
XOR2_X1 U817 ( .A(KEYINPUT56), .B(n1126), .Z(n1123) );
NOR2_X1 U818 ( .A1(G134), .A2(n1127), .ZN(n1126) );
NAND3_X1 U819 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1121) );
NAND2_X1 U820 ( .A1(KEYINPUT49), .A2(n1131), .ZN(n1129) );
OR2_X1 U821 ( .A1(n1132), .A2(KEYINPUT49), .ZN(n1128) );
XNOR2_X1 U822 ( .A(G131), .B(n1133), .ZN(n1119) );
NOR2_X1 U823 ( .A1(KEYINPUT43), .A2(n1134), .ZN(n1133) );
NOR2_X1 U824 ( .A1(G900), .A2(n1135), .ZN(n1117) );
NAND2_X1 U825 ( .A1(n1135), .A2(n1136), .ZN(n1115) );
NOR2_X1 U826 ( .A1(n1137), .A2(n1135), .ZN(n1112) );
XOR2_X1 U827 ( .A(n1138), .B(KEYINPUT45), .Z(n1137) );
NAND2_X1 U828 ( .A1(G900), .A2(G227), .ZN(n1138) );
XOR2_X1 U829 ( .A(n1139), .B(n1140), .Z(G69) );
NOR2_X1 U830 ( .A1(n1141), .A2(n1135), .ZN(n1140) );
AND2_X1 U831 ( .A1(G224), .A2(G898), .ZN(n1141) );
NOR2_X1 U832 ( .A1(KEYINPUT62), .A2(n1142), .ZN(n1139) );
XOR2_X1 U833 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR3_X1 U834 ( .A1(n1145), .A2(KEYINPUT60), .A3(n1146), .ZN(n1144) );
XOR2_X1 U835 ( .A(n1147), .B(n1148), .Z(n1145) );
NAND2_X1 U836 ( .A1(n1135), .A2(n1149), .ZN(n1143) );
NOR2_X1 U837 ( .A1(n1150), .A2(n1151), .ZN(G66) );
XNOR2_X1 U838 ( .A(n1152), .B(n1153), .ZN(n1151) );
XOR2_X1 U839 ( .A(n1154), .B(KEYINPUT16), .Z(n1153) );
NAND2_X1 U840 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U841 ( .A1(n1150), .A2(n1157), .ZN(G63) );
XOR2_X1 U842 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND2_X1 U843 ( .A1(n1155), .A2(n1160), .ZN(n1158) );
XOR2_X1 U844 ( .A(KEYINPUT41), .B(G478), .Z(n1160) );
NOR3_X1 U845 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(G60) );
NOR3_X1 U846 ( .A1(n1164), .A2(G953), .A3(G952), .ZN(n1163) );
AND2_X1 U847 ( .A1(n1164), .A2(n1150), .ZN(n1162) );
INV_X1 U848 ( .A(KEYINPUT7), .ZN(n1164) );
NOR2_X1 U849 ( .A1(n1165), .A2(n1166), .ZN(n1161) );
XOR2_X1 U850 ( .A(n1167), .B(KEYINPUT20), .Z(n1166) );
NAND2_X1 U851 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U852 ( .A1(n1168), .A2(n1169), .ZN(n1165) );
AND2_X1 U853 ( .A1(n1155), .A2(G475), .ZN(n1168) );
XOR2_X1 U854 ( .A(n1170), .B(n1171), .Z(G6) );
XNOR2_X1 U855 ( .A(KEYINPUT30), .B(n1172), .ZN(n1171) );
NOR2_X1 U856 ( .A1(n1150), .A2(n1173), .ZN(G57) );
XOR2_X1 U857 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U858 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U859 ( .A(n1178), .B(n1179), .Z(n1177) );
NAND2_X1 U860 ( .A1(KEYINPUT12), .A2(n1180), .ZN(n1179) );
NAND2_X1 U861 ( .A1(n1155), .A2(G472), .ZN(n1178) );
XOR2_X1 U862 ( .A(n1181), .B(n1182), .Z(n1174) );
XNOR2_X1 U863 ( .A(KEYINPUT27), .B(n1183), .ZN(n1182) );
NOR2_X1 U864 ( .A1(n1150), .A2(n1184), .ZN(G54) );
XOR2_X1 U865 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U866 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U867 ( .A(n1189), .B(n1190), .Z(n1187) );
NAND2_X1 U868 ( .A1(n1155), .A2(G469), .ZN(n1189) );
XOR2_X1 U869 ( .A(n1191), .B(n1192), .Z(n1185) );
XOR2_X1 U870 ( .A(G110), .B(n1193), .Z(n1192) );
XNOR2_X1 U871 ( .A(G140), .B(KEYINPUT58), .ZN(n1191) );
NOR2_X1 U872 ( .A1(n1150), .A2(n1194), .ZN(G51) );
XOR2_X1 U873 ( .A(n1195), .B(n1196), .Z(n1194) );
XNOR2_X1 U874 ( .A(n1197), .B(n1198), .ZN(n1196) );
XOR2_X1 U875 ( .A(n1199), .B(n1200), .Z(n1195) );
XNOR2_X1 U876 ( .A(n1201), .B(n1202), .ZN(n1200) );
NAND2_X1 U877 ( .A1(n1155), .A2(n1203), .ZN(n1199) );
AND2_X1 U878 ( .A1(G902), .A2(n1204), .ZN(n1155) );
NAND2_X1 U879 ( .A1(n1205), .A2(n1088), .ZN(n1204) );
INV_X1 U880 ( .A(n1136), .ZN(n1088) );
NAND4_X1 U881 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1136) );
NOR4_X1 U882 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1209) );
INV_X1 U883 ( .A(n1214), .ZN(n1213) );
NOR2_X1 U884 ( .A1(n1215), .A2(n1216), .ZN(n1208) );
NOR2_X1 U885 ( .A1(KEYINPUT39), .A2(n1217), .ZN(n1216) );
INV_X1 U886 ( .A(n1218), .ZN(n1215) );
NAND2_X1 U887 ( .A1(n1219), .A2(n1220), .ZN(n1207) );
NAND3_X1 U888 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1220) );
OR3_X1 U889 ( .A1(n1224), .A2(KEYINPUT2), .A3(n1225), .ZN(n1223) );
NAND4_X1 U890 ( .A1(n1084), .A2(n1226), .A3(n1086), .A4(n1227), .ZN(n1222) );
AND2_X1 U891 ( .A1(KEYINPUT39), .A2(n1079), .ZN(n1227) );
NAND4_X1 U892 ( .A1(n1228), .A2(n1083), .A3(n1229), .A4(n1230), .ZN(n1221) );
NAND4_X1 U893 ( .A1(n1231), .A2(n1053), .A3(KEYINPUT2), .A4(n1076), .ZN(n1206) );
XNOR2_X1 U894 ( .A(n1087), .B(KEYINPUT15), .ZN(n1205) );
INV_X1 U895 ( .A(n1149), .ZN(n1087) );
NAND2_X1 U896 ( .A1(n1232), .A2(n1233), .ZN(n1149) );
AND4_X1 U897 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1233) );
AND4_X1 U898 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1170), .ZN(n1232) );
NAND3_X1 U899 ( .A1(n1051), .A2(n1052), .A3(n1086), .ZN(n1170) );
OR3_X1 U900 ( .A1(n1241), .A2(n1242), .A3(n1224), .ZN(n1240) );
NAND3_X1 U901 ( .A1(n1243), .A2(n1244), .A3(n1245), .ZN(n1241) );
XNOR2_X1 U902 ( .A(KEYINPUT47), .B(n1076), .ZN(n1245) );
XNOR2_X1 U903 ( .A(KEYINPUT19), .B(n1065), .ZN(n1243) );
NOR2_X1 U904 ( .A1(n1135), .A2(G952), .ZN(n1150) );
XOR2_X1 U905 ( .A(G146), .B(n1212), .Z(G48) );
AND3_X1 U906 ( .A1(n1086), .A2(n1219), .A3(n1231), .ZN(n1212) );
INV_X1 U907 ( .A(n1225), .ZN(n1231) );
XNOR2_X1 U908 ( .A(G143), .B(n1246), .ZN(G45) );
NAND4_X1 U909 ( .A1(n1219), .A2(n1247), .A3(n1083), .A4(n1248), .ZN(n1246) );
NOR3_X1 U910 ( .A1(n1095), .A2(n1249), .A3(n1250), .ZN(n1248) );
XNOR2_X1 U911 ( .A(KEYINPUT1), .B(n1242), .ZN(n1247) );
XNOR2_X1 U912 ( .A(G140), .B(n1218), .ZN(G42) );
NAND4_X1 U913 ( .A1(n1228), .A2(n1251), .A3(n1086), .A4(n1084), .ZN(n1218) );
XNOR2_X1 U914 ( .A(n1127), .B(n1211), .ZN(G39) );
NOR3_X1 U915 ( .A1(n1069), .A2(n1063), .A3(n1225), .ZN(n1211) );
INV_X1 U916 ( .A(n1252), .ZN(n1063) );
XNOR2_X1 U917 ( .A(G134), .B(n1214), .ZN(G36) );
NAND4_X1 U918 ( .A1(n1228), .A2(n1251), .A3(n1083), .A4(n1053), .ZN(n1214) );
XNOR2_X1 U919 ( .A(n1210), .B(n1253), .ZN(G33) );
NAND2_X1 U920 ( .A1(KEYINPUT54), .A2(G131), .ZN(n1253) );
AND4_X1 U921 ( .A1(n1228), .A2(n1251), .A3(n1083), .A4(n1086), .ZN(n1210) );
INV_X1 U922 ( .A(n1069), .ZN(n1251) );
NAND2_X1 U923 ( .A1(n1091), .A2(n1093), .ZN(n1069) );
XOR2_X1 U924 ( .A(G128), .B(n1254), .Z(G30) );
NOR3_X1 U925 ( .A1(n1225), .A2(n1076), .A3(n1224), .ZN(n1254) );
INV_X1 U926 ( .A(n1053), .ZN(n1224) );
INV_X1 U927 ( .A(n1219), .ZN(n1076) );
NAND3_X1 U928 ( .A1(n1108), .A2(n1255), .A3(n1228), .ZN(n1225) );
NOR2_X1 U929 ( .A1(n1242), .A2(n1249), .ZN(n1228) );
XNOR2_X1 U930 ( .A(G101), .B(n1239), .ZN(G3) );
NAND3_X1 U931 ( .A1(n1252), .A2(n1052), .A3(n1083), .ZN(n1239) );
XOR2_X1 U932 ( .A(n1217), .B(n1256), .Z(G27) );
NAND2_X1 U933 ( .A1(KEYINPUT32), .A2(G125), .ZN(n1256) );
NAND4_X1 U934 ( .A1(n1086), .A2(n1084), .A3(n1257), .A4(n1219), .ZN(n1217) );
NOR2_X1 U935 ( .A1(n1249), .A2(n1079), .ZN(n1257) );
INV_X1 U936 ( .A(n1077), .ZN(n1079) );
INV_X1 U937 ( .A(n1226), .ZN(n1249) );
NAND2_X1 U938 ( .A1(n1060), .A2(n1258), .ZN(n1226) );
NAND4_X1 U939 ( .A1(G902), .A2(G953), .A3(n1259), .A4(n1260), .ZN(n1258) );
INV_X1 U940 ( .A(G900), .ZN(n1260) );
XNOR2_X1 U941 ( .A(G122), .B(n1238), .ZN(G24) );
NAND4_X1 U942 ( .A1(n1261), .A2(n1051), .A3(n1229), .A4(n1230), .ZN(n1238) );
INV_X1 U943 ( .A(n1065), .ZN(n1051) );
NAND2_X1 U944 ( .A1(n1262), .A2(n1263), .ZN(n1065) );
XNOR2_X1 U945 ( .A(G119), .B(n1237), .ZN(G21) );
NAND4_X1 U946 ( .A1(n1261), .A2(n1252), .A3(n1108), .A4(n1255), .ZN(n1237) );
XNOR2_X1 U947 ( .A(G116), .B(n1236), .ZN(G18) );
NAND3_X1 U948 ( .A1(n1261), .A2(n1053), .A3(n1083), .ZN(n1236) );
NOR2_X1 U949 ( .A1(n1230), .A2(n1095), .ZN(n1053) );
INV_X1 U950 ( .A(n1229), .ZN(n1095) );
XNOR2_X1 U951 ( .A(G113), .B(n1235), .ZN(G15) );
NAND3_X1 U952 ( .A1(n1261), .A2(n1086), .A3(n1083), .ZN(n1235) );
AND2_X1 U953 ( .A1(n1263), .A2(n1255), .ZN(n1083) );
INV_X1 U954 ( .A(n1108), .ZN(n1263) );
NOR2_X1 U955 ( .A1(n1229), .A2(n1250), .ZN(n1086) );
INV_X1 U956 ( .A(n1230), .ZN(n1250) );
AND3_X1 U957 ( .A1(n1077), .A2(n1244), .A3(n1219), .ZN(n1261) );
NAND2_X1 U958 ( .A1(n1264), .A2(n1265), .ZN(n1077) );
OR2_X1 U959 ( .A1(n1242), .A2(KEYINPUT17), .ZN(n1265) );
INV_X1 U960 ( .A(n1070), .ZN(n1242) );
NAND3_X1 U961 ( .A1(n1074), .A2(n1072), .A3(KEYINPUT17), .ZN(n1264) );
XNOR2_X1 U962 ( .A(G110), .B(n1234), .ZN(G12) );
NAND3_X1 U963 ( .A1(n1084), .A2(n1052), .A3(n1252), .ZN(n1234) );
NOR2_X1 U964 ( .A1(n1229), .A2(n1230), .ZN(n1252) );
XNOR2_X1 U965 ( .A(n1102), .B(G475), .ZN(n1230) );
OR2_X1 U966 ( .A1(n1169), .A2(G902), .ZN(n1102) );
XOR2_X1 U967 ( .A(n1266), .B(n1267), .Z(n1169) );
XOR2_X1 U968 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U969 ( .A(n1270), .B(n1271), .Z(n1269) );
AND3_X1 U970 ( .A1(G214), .A2(n1135), .A3(n1272), .ZN(n1271) );
NAND2_X1 U971 ( .A1(n1273), .A2(n1274), .ZN(n1270) );
NAND3_X1 U972 ( .A1(n1130), .A2(n1132), .A3(n1275), .ZN(n1274) );
XNOR2_X1 U973 ( .A(n1276), .B(n1172), .ZN(n1275) );
INV_X1 U974 ( .A(n1277), .ZN(n1130) );
NAND2_X1 U975 ( .A1(n1278), .A2(n1279), .ZN(n1273) );
XNOR2_X1 U976 ( .A(G104), .B(n1276), .ZN(n1279) );
NAND2_X1 U977 ( .A1(n1280), .A2(KEYINPUT22), .ZN(n1276) );
XOR2_X1 U978 ( .A(n1281), .B(G113), .Z(n1280) );
NAND2_X1 U979 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
INV_X1 U980 ( .A(G122), .ZN(n1283) );
XNOR2_X1 U981 ( .A(KEYINPUT37), .B(KEYINPUT24), .ZN(n1282) );
XNOR2_X1 U982 ( .A(G140), .B(G125), .ZN(n1278) );
NAND2_X1 U983 ( .A1(KEYINPUT31), .A2(n1284), .ZN(n1268) );
XNOR2_X1 U984 ( .A(G143), .B(n1285), .ZN(n1266) );
XOR2_X1 U985 ( .A(KEYINPUT21), .B(G146), .Z(n1285) );
XNOR2_X1 U986 ( .A(n1286), .B(G478), .ZN(n1229) );
NAND2_X1 U987 ( .A1(n1159), .A2(n1287), .ZN(n1286) );
XNOR2_X1 U988 ( .A(n1288), .B(n1289), .ZN(n1159) );
XOR2_X1 U989 ( .A(n1290), .B(n1291), .Z(n1289) );
XNOR2_X1 U990 ( .A(n1292), .B(n1293), .ZN(n1291) );
INV_X1 U991 ( .A(G107), .ZN(n1293) );
NAND2_X1 U992 ( .A1(KEYINPUT51), .A2(G143), .ZN(n1292) );
NAND2_X1 U993 ( .A1(G217), .A2(n1294), .ZN(n1290) );
XOR2_X1 U994 ( .A(n1295), .B(n1296), .Z(n1288) );
XNOR2_X1 U995 ( .A(n1297), .B(G128), .ZN(n1296) );
XNOR2_X1 U996 ( .A(G116), .B(G122), .ZN(n1295) );
AND3_X1 U997 ( .A1(n1070), .A2(n1244), .A3(n1219), .ZN(n1052) );
NOR2_X1 U998 ( .A1(n1091), .A2(n1098), .ZN(n1219) );
INV_X1 U999 ( .A(n1093), .ZN(n1098) );
NAND2_X1 U1000 ( .A1(G214), .A2(n1298), .ZN(n1093) );
XOR2_X1 U1001 ( .A(n1107), .B(KEYINPUT59), .Z(n1091) );
XNOR2_X1 U1002 ( .A(n1299), .B(n1203), .ZN(n1107) );
AND2_X1 U1003 ( .A1(G210), .A2(n1298), .ZN(n1203) );
NAND2_X1 U1004 ( .A1(n1272), .A2(n1287), .ZN(n1298) );
NAND2_X1 U1005 ( .A1(n1300), .A2(n1287), .ZN(n1299) );
XOR2_X1 U1006 ( .A(n1301), .B(n1302), .Z(n1300) );
XNOR2_X1 U1007 ( .A(n1303), .B(n1304), .ZN(n1302) );
NAND2_X1 U1008 ( .A1(KEYINPUT23), .A2(n1202), .ZN(n1304) );
AND2_X1 U1009 ( .A1(G224), .A2(n1135), .ZN(n1202) );
NAND2_X1 U1010 ( .A1(KEYINPUT48), .A2(n1198), .ZN(n1303) );
XOR2_X1 U1011 ( .A(n1305), .B(n1148), .Z(n1198) );
XOR2_X1 U1012 ( .A(G110), .B(n1306), .Z(n1148) );
NOR2_X1 U1013 ( .A1(G122), .A2(KEYINPUT5), .ZN(n1306) );
NAND2_X1 U1014 ( .A1(KEYINPUT9), .A2(n1147), .ZN(n1305) );
XOR2_X1 U1015 ( .A(n1307), .B(n1308), .Z(n1147) );
XNOR2_X1 U1016 ( .A(n1309), .B(n1183), .ZN(n1307) );
NAND2_X1 U1017 ( .A1(KEYINPUT8), .A2(n1310), .ZN(n1309) );
XOR2_X1 U1018 ( .A(n1311), .B(KEYINPUT10), .Z(n1301) );
NAND2_X1 U1019 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NAND2_X1 U1020 ( .A1(n1197), .A2(n1314), .ZN(n1313) );
NAND2_X1 U1021 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND2_X1 U1022 ( .A1(G125), .A2(n1317), .ZN(n1316) );
INV_X1 U1023 ( .A(KEYINPUT61), .ZN(n1315) );
NAND2_X1 U1024 ( .A1(n1318), .A2(n1201), .ZN(n1312) );
NAND2_X1 U1025 ( .A1(n1317), .A2(n1319), .ZN(n1318) );
OR2_X1 U1026 ( .A1(n1197), .A2(KEYINPUT61), .ZN(n1319) );
INV_X1 U1027 ( .A(KEYINPUT42), .ZN(n1317) );
NAND2_X1 U1028 ( .A1(n1060), .A2(n1320), .ZN(n1244) );
NAND3_X1 U1029 ( .A1(n1146), .A2(n1259), .A3(G902), .ZN(n1320) );
NOR2_X1 U1030 ( .A1(n1135), .A2(G898), .ZN(n1146) );
NAND3_X1 U1031 ( .A1(n1259), .A2(n1135), .A3(G952), .ZN(n1060) );
NAND2_X1 U1032 ( .A1(G237), .A2(G234), .ZN(n1259) );
NOR2_X1 U1033 ( .A1(n1074), .A2(n1099), .ZN(n1070) );
INV_X1 U1034 ( .A(n1072), .ZN(n1099) );
NAND2_X1 U1035 ( .A1(G221), .A2(n1321), .ZN(n1072) );
XNOR2_X1 U1036 ( .A(n1105), .B(n1322), .ZN(n1074) );
NOR2_X1 U1037 ( .A1(KEYINPUT6), .A2(n1323), .ZN(n1322) );
XNOR2_X1 U1038 ( .A(G469), .B(KEYINPUT63), .ZN(n1323) );
NAND2_X1 U1039 ( .A1(n1324), .A2(n1287), .ZN(n1105) );
XOR2_X1 U1040 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1041 ( .A(n1327), .B(n1188), .Z(n1326) );
NAND2_X1 U1042 ( .A1(KEYINPUT40), .A2(n1193), .ZN(n1327) );
AND2_X1 U1043 ( .A1(G227), .A2(n1135), .ZN(n1193) );
XOR2_X1 U1044 ( .A(n1328), .B(n1329), .Z(n1325) );
NOR2_X1 U1045 ( .A1(G110), .A2(KEYINPUT34), .ZN(n1329) );
XNOR2_X1 U1046 ( .A(n1330), .B(n1131), .ZN(n1328) );
INV_X1 U1047 ( .A(G140), .ZN(n1131) );
NAND2_X1 U1048 ( .A1(KEYINPUT36), .A2(n1190), .ZN(n1330) );
XNOR2_X1 U1049 ( .A(n1331), .B(n1134), .ZN(n1190) );
XNOR2_X1 U1050 ( .A(n1332), .B(n1333), .ZN(n1134) );
XOR2_X1 U1051 ( .A(G146), .B(n1334), .Z(n1333) );
NOR2_X1 U1052 ( .A1(G143), .A2(KEYINPUT35), .ZN(n1334) );
NAND2_X1 U1053 ( .A1(KEYINPUT44), .A2(G128), .ZN(n1332) );
NAND3_X1 U1054 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1331) );
OR2_X1 U1055 ( .A1(n1183), .A2(n1338), .ZN(n1337) );
NAND3_X1 U1056 ( .A1(n1338), .A2(n1183), .A3(KEYINPUT55), .ZN(n1336) );
INV_X1 U1057 ( .A(G101), .ZN(n1183) );
NOR2_X1 U1058 ( .A1(KEYINPUT11), .A2(n1339), .ZN(n1338) );
INV_X1 U1059 ( .A(n1310), .ZN(n1339) );
OR2_X1 U1060 ( .A1(n1310), .A2(KEYINPUT55), .ZN(n1335) );
XNOR2_X1 U1061 ( .A(G107), .B(n1172), .ZN(n1310) );
INV_X1 U1062 ( .A(G104), .ZN(n1172) );
AND2_X1 U1063 ( .A1(n1262), .A2(n1108), .ZN(n1084) );
XNOR2_X1 U1064 ( .A(n1340), .B(n1156), .ZN(n1108) );
AND2_X1 U1065 ( .A1(G217), .A2(n1321), .ZN(n1156) );
NAND2_X1 U1066 ( .A1(G234), .A2(n1287), .ZN(n1321) );
NAND2_X1 U1067 ( .A1(n1152), .A2(n1287), .ZN(n1340) );
XNOR2_X1 U1068 ( .A(n1341), .B(n1342), .ZN(n1152) );
XOR2_X1 U1069 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1070 ( .A(n1345), .B(n1346), .Z(n1344) );
NAND2_X1 U1071 ( .A1(G221), .A2(n1294), .ZN(n1345) );
AND2_X1 U1072 ( .A1(G234), .A2(n1135), .ZN(n1294) );
XOR2_X1 U1073 ( .A(n1347), .B(n1348), .Z(n1343) );
NOR2_X1 U1074 ( .A1(G110), .A2(KEYINPUT52), .ZN(n1348) );
NAND3_X1 U1075 ( .A1(n1349), .A2(n1350), .A3(n1132), .ZN(n1347) );
NAND2_X1 U1076 ( .A1(G140), .A2(G125), .ZN(n1132) );
OR2_X1 U1077 ( .A1(n1201), .A2(KEYINPUT38), .ZN(n1350) );
INV_X1 U1078 ( .A(G125), .ZN(n1201) );
NAND2_X1 U1079 ( .A1(n1277), .A2(KEYINPUT38), .ZN(n1349) );
NOR2_X1 U1080 ( .A1(G125), .A2(G140), .ZN(n1277) );
XOR2_X1 U1081 ( .A(n1351), .B(n1352), .Z(n1341) );
XOR2_X1 U1082 ( .A(KEYINPUT53), .B(KEYINPUT21), .Z(n1352) );
XNOR2_X1 U1083 ( .A(G119), .B(G137), .ZN(n1351) );
XNOR2_X1 U1084 ( .A(n1255), .B(KEYINPUT29), .ZN(n1262) );
XOR2_X1 U1085 ( .A(n1109), .B(n1111), .Z(n1255) );
INV_X1 U1086 ( .A(G472), .ZN(n1111) );
NAND3_X1 U1087 ( .A1(n1353), .A2(n1354), .A3(n1287), .ZN(n1109) );
INV_X1 U1088 ( .A(G902), .ZN(n1287) );
NAND2_X1 U1089 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
INV_X1 U1090 ( .A(KEYINPUT3), .ZN(n1356) );
XOR2_X1 U1091 ( .A(n1357), .B(n1358), .Z(n1355) );
NOR2_X1 U1092 ( .A1(KEYINPUT14), .A2(n1359), .ZN(n1357) );
NAND3_X1 U1093 ( .A1(n1360), .A2(n1361), .A3(KEYINPUT3), .ZN(n1353) );
INV_X1 U1094 ( .A(n1359), .ZN(n1361) );
NAND3_X1 U1095 ( .A1(n1362), .A2(n1363), .A3(n1364), .ZN(n1359) );
NAND2_X1 U1096 ( .A1(G101), .A2(n1365), .ZN(n1364) );
OR3_X1 U1097 ( .A1(n1365), .A2(G101), .A3(KEYINPUT25), .ZN(n1363) );
NAND2_X1 U1098 ( .A1(KEYINPUT4), .A2(n1366), .ZN(n1365) );
INV_X1 U1099 ( .A(n1181), .ZN(n1366) );
NAND2_X1 U1100 ( .A1(KEYINPUT25), .A2(n1181), .ZN(n1362) );
NAND3_X1 U1101 ( .A1(n1272), .A2(n1135), .A3(G210), .ZN(n1181) );
INV_X1 U1102 ( .A(G953), .ZN(n1135) );
INV_X1 U1103 ( .A(G237), .ZN(n1272) );
XOR2_X1 U1104 ( .A(KEYINPUT14), .B(n1358), .Z(n1360) );
XOR2_X1 U1105 ( .A(n1176), .B(n1180), .Z(n1358) );
NAND2_X1 U1106 ( .A1(n1367), .A2(n1368), .ZN(n1180) );
NAND3_X1 U1107 ( .A1(G113), .A2(n1369), .A3(n1370), .ZN(n1368) );
INV_X1 U1108 ( .A(KEYINPUT26), .ZN(n1370) );
NAND2_X1 U1109 ( .A1(n1308), .A2(KEYINPUT26), .ZN(n1367) );
XOR2_X1 U1110 ( .A(G113), .B(n1369), .Z(n1308) );
XOR2_X1 U1111 ( .A(G116), .B(G119), .Z(n1369) );
XNOR2_X1 U1112 ( .A(n1197), .B(n1188), .ZN(n1176) );
XNOR2_X1 U1113 ( .A(n1284), .B(n1371), .ZN(n1188) );
NOR2_X1 U1114 ( .A1(n1125), .A2(n1372), .ZN(n1371) );
XOR2_X1 U1115 ( .A(n1373), .B(KEYINPUT0), .Z(n1372) );
NAND2_X1 U1116 ( .A1(n1374), .A2(n1297), .ZN(n1373) );
XNOR2_X1 U1117 ( .A(KEYINPUT28), .B(n1127), .ZN(n1374) );
INV_X1 U1118 ( .A(G137), .ZN(n1127) );
NOR2_X1 U1119 ( .A1(n1297), .A2(G137), .ZN(n1125) );
INV_X1 U1120 ( .A(G134), .ZN(n1297) );
INV_X1 U1121 ( .A(G131), .ZN(n1284) );
XOR2_X1 U1122 ( .A(G143), .B(n1346), .Z(n1197) );
XOR2_X1 U1123 ( .A(G128), .B(G146), .Z(n1346) );
endmodule


