//Key = 0001111010110000110000001000000100100010111110101000011101000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
n1425, n1426, n1427, n1428, n1429, n1430, n1431;

XOR2_X1 U780 ( .A(n1085), .B(n1086), .Z(G9) );
XOR2_X1 U781 ( .A(KEYINPUT48), .B(G107), .Z(n1086) );
NOR2_X1 U782 ( .A1(n1087), .A2(n1088), .ZN(G75) );
XOR2_X1 U783 ( .A(n1089), .B(KEYINPUT44), .Z(n1088) );
NAND3_X1 U784 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
NOR3_X1 U785 ( .A1(n1093), .A2(n1090), .A3(n1094), .ZN(n1087) );
INV_X1 U786 ( .A(G952), .ZN(n1090) );
NAND3_X1 U787 ( .A1(n1095), .A2(n1091), .A3(n1096), .ZN(n1093) );
XNOR2_X1 U788 ( .A(KEYINPUT40), .B(n1092), .ZN(n1096) );
NAND4_X1 U789 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1092) );
NOR4_X1 U790 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1100) );
NOR2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1102) );
INV_X1 U792 ( .A(KEYINPUT51), .ZN(n1106) );
NOR3_X1 U793 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1105) );
NOR2_X1 U794 ( .A1(KEYINPUT51), .A2(n1110), .ZN(n1101) );
XOR2_X1 U795 ( .A(KEYINPUT53), .B(n1111), .Z(n1098) );
NAND2_X1 U796 ( .A1(n1112), .A2(n1113), .ZN(n1095) );
NAND2_X1 U797 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND4_X1 U798 ( .A1(n1099), .A2(n1116), .A3(n1097), .A4(n1117), .ZN(n1115) );
NAND2_X1 U799 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U800 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U801 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U802 ( .A1(n1109), .A2(n1124), .ZN(n1123) );
NAND2_X1 U803 ( .A1(n1110), .A2(n1125), .ZN(n1118) );
NAND2_X1 U804 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
OR2_X1 U805 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U806 ( .A(KEYINPUT16), .B(n1130), .Z(n1126) );
NAND3_X1 U807 ( .A1(n1110), .A2(n1131), .A3(n1120), .ZN(n1114) );
NAND2_X1 U808 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NAND3_X1 U809 ( .A1(n1134), .A2(n1135), .A3(n1097), .ZN(n1133) );
NAND2_X1 U810 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND3_X1 U811 ( .A1(n1138), .A2(n1139), .A3(n1099), .ZN(n1134) );
NAND2_X1 U812 ( .A1(n1116), .A2(n1140), .ZN(n1132) );
INV_X1 U813 ( .A(n1141), .ZN(n1112) );
XOR2_X1 U814 ( .A(n1142), .B(n1143), .Z(G72) );
XOR2_X1 U815 ( .A(n1144), .B(n1145), .Z(n1143) );
NAND2_X1 U816 ( .A1(G953), .A2(n1146), .ZN(n1145) );
NAND2_X1 U817 ( .A1(G900), .A2(G227), .ZN(n1146) );
NAND2_X1 U818 ( .A1(n1147), .A2(n1148), .ZN(n1144) );
NAND2_X1 U819 ( .A1(G953), .A2(n1149), .ZN(n1148) );
XOR2_X1 U820 ( .A(n1150), .B(n1151), .Z(n1147) );
XOR2_X1 U821 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U822 ( .A(n1154), .B(n1155), .Z(n1150) );
XNOR2_X1 U823 ( .A(KEYINPUT52), .B(n1156), .ZN(n1155) );
NOR2_X1 U824 ( .A1(KEYINPUT23), .A2(n1157), .ZN(n1156) );
NOR2_X1 U825 ( .A1(n1158), .A2(G953), .ZN(n1142) );
NAND2_X1 U826 ( .A1(n1159), .A2(n1160), .ZN(G69) );
NAND2_X1 U827 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U828 ( .A1(G953), .A2(n1163), .ZN(n1161) );
NAND2_X1 U829 ( .A1(G898), .A2(G224), .ZN(n1163) );
NAND2_X1 U830 ( .A1(n1164), .A2(n1165), .ZN(n1159) );
NAND2_X1 U831 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
OR2_X1 U832 ( .A1(n1091), .A2(G224), .ZN(n1167) );
INV_X1 U833 ( .A(n1168), .ZN(n1166) );
INV_X1 U834 ( .A(n1162), .ZN(n1164) );
NAND2_X1 U835 ( .A1(n1169), .A2(n1170), .ZN(n1162) );
NAND2_X1 U836 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XOR2_X1 U837 ( .A(KEYINPUT38), .B(n1173), .Z(n1169) );
NOR3_X1 U838 ( .A1(n1172), .A2(n1168), .A3(n1171), .ZN(n1173) );
AND2_X1 U839 ( .A1(n1091), .A2(n1174), .ZN(n1171) );
NAND2_X1 U840 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND2_X1 U841 ( .A1(n1177), .A2(n1178), .ZN(n1172) );
NAND2_X1 U842 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NAND2_X1 U843 ( .A1(n1181), .A2(n1182), .ZN(n1177) );
XOR2_X1 U844 ( .A(n1180), .B(n1183), .Z(n1182) );
XOR2_X1 U845 ( .A(KEYINPUT26), .B(KEYINPUT17), .Z(n1183) );
NAND2_X1 U846 ( .A1(n1184), .A2(n1185), .ZN(n1180) );
XOR2_X1 U847 ( .A(n1186), .B(KEYINPUT33), .Z(n1184) );
NOR2_X1 U848 ( .A1(n1187), .A2(n1188), .ZN(G66) );
XNOR2_X1 U849 ( .A(n1189), .B(n1190), .ZN(n1188) );
NOR2_X1 U850 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NOR2_X1 U851 ( .A1(n1187), .A2(n1193), .ZN(G63) );
XNOR2_X1 U852 ( .A(n1194), .B(n1195), .ZN(n1193) );
NOR2_X1 U853 ( .A1(n1192), .A2(n1196), .ZN(n1195) );
XOR2_X1 U854 ( .A(KEYINPUT34), .B(G478), .Z(n1196) );
NOR2_X1 U855 ( .A1(n1187), .A2(n1197), .ZN(G60) );
NOR2_X1 U856 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U857 ( .A(n1200), .B(n1201), .Z(n1199) );
NOR2_X1 U858 ( .A1(n1202), .A2(n1192), .ZN(n1201) );
INV_X1 U859 ( .A(G475), .ZN(n1202) );
AND2_X1 U860 ( .A1(n1203), .A2(KEYINPUT4), .ZN(n1200) );
NOR2_X1 U861 ( .A1(KEYINPUT4), .A2(n1203), .ZN(n1198) );
NAND2_X1 U862 ( .A1(n1204), .A2(n1205), .ZN(G6) );
OR2_X1 U863 ( .A1(n1206), .A2(G104), .ZN(n1205) );
XOR2_X1 U864 ( .A(n1207), .B(KEYINPUT20), .Z(n1204) );
NAND2_X1 U865 ( .A1(G104), .A2(n1206), .ZN(n1207) );
NOR2_X1 U866 ( .A1(n1187), .A2(n1208), .ZN(G57) );
XOR2_X1 U867 ( .A(n1209), .B(n1210), .Z(n1208) );
XOR2_X1 U868 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U869 ( .A(n1213), .B(n1214), .Z(n1209) );
NOR2_X1 U870 ( .A1(n1215), .A2(n1192), .ZN(n1214) );
INV_X1 U871 ( .A(G472), .ZN(n1215) );
NAND3_X1 U872 ( .A1(n1216), .A2(n1217), .A3(KEYINPUT57), .ZN(n1213) );
NAND2_X1 U873 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
INV_X1 U874 ( .A(KEYINPUT29), .ZN(n1219) );
XOR2_X1 U875 ( .A(G101), .B(n1220), .Z(n1218) );
NAND3_X1 U876 ( .A1(n1220), .A2(G101), .A3(KEYINPUT29), .ZN(n1216) );
NOR2_X1 U877 ( .A1(n1187), .A2(n1221), .ZN(G54) );
XOR2_X1 U878 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR2_X1 U879 ( .A1(KEYINPUT63), .A2(n1224), .ZN(n1223) );
XOR2_X1 U880 ( .A(n1225), .B(n1226), .Z(n1224) );
XOR2_X1 U881 ( .A(n1227), .B(n1211), .Z(n1226) );
XOR2_X1 U882 ( .A(n1228), .B(n1229), .Z(n1225) );
NOR2_X1 U883 ( .A1(KEYINPUT35), .A2(n1230), .ZN(n1229) );
XOR2_X1 U884 ( .A(n1231), .B(n1153), .Z(n1230) );
OR2_X1 U885 ( .A1(n1192), .A2(n1107), .ZN(n1222) );
INV_X1 U886 ( .A(G469), .ZN(n1107) );
NOR2_X1 U887 ( .A1(n1187), .A2(n1232), .ZN(G51) );
XOR2_X1 U888 ( .A(n1233), .B(n1234), .Z(n1232) );
XOR2_X1 U889 ( .A(n1235), .B(n1236), .Z(n1234) );
XOR2_X1 U890 ( .A(n1237), .B(n1238), .Z(n1236) );
NOR2_X1 U891 ( .A1(n1239), .A2(n1192), .ZN(n1237) );
NAND2_X1 U892 ( .A1(G902), .A2(n1094), .ZN(n1192) );
NAND3_X1 U893 ( .A1(n1175), .A2(n1240), .A3(n1158), .ZN(n1094) );
AND4_X1 U894 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1158) );
NOR4_X1 U895 ( .A1(n1245), .A2(n1246), .A3(n1247), .A4(n1248), .ZN(n1244) );
NOR3_X1 U896 ( .A1(n1249), .A2(n1138), .A3(n1250), .ZN(n1248) );
XOR2_X1 U897 ( .A(KEYINPUT10), .B(n1130), .Z(n1249) );
INV_X1 U898 ( .A(n1251), .ZN(n1247) );
NOR2_X1 U899 ( .A1(n1252), .A2(n1253), .ZN(n1243) );
XNOR2_X1 U900 ( .A(KEYINPUT43), .B(n1176), .ZN(n1240) );
AND4_X1 U901 ( .A1(n1206), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1175) );
AND4_X1 U902 ( .A1(n1257), .A2(n1085), .A3(n1258), .A4(n1259), .ZN(n1256) );
NAND3_X1 U903 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1085) );
NAND4_X1 U904 ( .A1(n1263), .A2(n1264), .A3(n1265), .A4(n1266), .ZN(n1255) );
NOR2_X1 U905 ( .A1(n1138), .A2(n1267), .ZN(n1266) );
XOR2_X1 U906 ( .A(KEYINPUT36), .B(n1130), .Z(n1265) );
XOR2_X1 U907 ( .A(KEYINPUT58), .B(n1140), .Z(n1263) );
NAND3_X1 U908 ( .A1(n1268), .A2(n1264), .A3(n1269), .ZN(n1254) );
XOR2_X1 U909 ( .A(KEYINPUT37), .B(n1130), .Z(n1268) );
NAND3_X1 U910 ( .A1(n1262), .A2(n1260), .A3(n1270), .ZN(n1206) );
XOR2_X1 U911 ( .A(n1271), .B(n1272), .Z(n1233) );
NOR2_X1 U912 ( .A1(KEYINPUT56), .A2(n1273), .ZN(n1272) );
XOR2_X1 U913 ( .A(n1274), .B(KEYINPUT54), .Z(n1271) );
NOR2_X1 U914 ( .A1(n1091), .A2(G952), .ZN(n1187) );
XOR2_X1 U915 ( .A(n1275), .B(n1276), .Z(G48) );
NAND3_X1 U916 ( .A1(n1270), .A2(n1130), .A3(n1277), .ZN(n1276) );
NAND2_X1 U917 ( .A1(KEYINPUT8), .A2(G146), .ZN(n1275) );
XOR2_X1 U918 ( .A(n1278), .B(n1251), .Z(G45) );
NAND3_X1 U919 ( .A1(n1279), .A2(n1130), .A3(n1280), .ZN(n1251) );
NOR3_X1 U920 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1280) );
XOR2_X1 U921 ( .A(G140), .B(n1246), .Z(G42) );
AND3_X1 U922 ( .A1(n1284), .A2(n1262), .A3(n1120), .ZN(n1246) );
XOR2_X1 U923 ( .A(G137), .B(n1245), .Z(G39) );
NOR3_X1 U924 ( .A1(n1103), .A2(n1250), .A3(n1137), .ZN(n1245) );
XNOR2_X1 U925 ( .A(G134), .B(n1241), .ZN(G36) );
NAND4_X1 U926 ( .A1(n1279), .A2(n1120), .A3(n1261), .A4(n1285), .ZN(n1241) );
XNOR2_X1 U927 ( .A(n1242), .B(n1286), .ZN(G33) );
NOR2_X1 U928 ( .A1(KEYINPUT28), .A2(n1157), .ZN(n1286) );
NAND4_X1 U929 ( .A1(n1279), .A2(n1120), .A3(n1270), .A4(n1285), .ZN(n1242) );
INV_X1 U930 ( .A(n1138), .ZN(n1270) );
INV_X1 U931 ( .A(n1103), .ZN(n1120) );
NAND2_X1 U932 ( .A1(n1287), .A2(n1129), .ZN(n1103) );
INV_X1 U933 ( .A(n1128), .ZN(n1287) );
XOR2_X1 U934 ( .A(G128), .B(n1253), .Z(G30) );
AND3_X1 U935 ( .A1(n1261), .A2(n1130), .A3(n1277), .ZN(n1253) );
INV_X1 U936 ( .A(n1250), .ZN(n1277) );
NAND4_X1 U937 ( .A1(n1262), .A2(n1288), .A3(n1136), .A4(n1285), .ZN(n1250) );
INV_X1 U938 ( .A(n1139), .ZN(n1261) );
XNOR2_X1 U939 ( .A(G101), .B(n1289), .ZN(G3) );
NAND2_X1 U940 ( .A1(n1269), .A2(n1290), .ZN(n1289) );
AND2_X1 U941 ( .A1(n1116), .A2(n1279), .ZN(n1269) );
AND2_X1 U942 ( .A1(n1140), .A2(n1262), .ZN(n1279) );
INV_X1 U943 ( .A(n1137), .ZN(n1116) );
XOR2_X1 U944 ( .A(G125), .B(n1252), .Z(G27) );
AND3_X1 U945 ( .A1(n1284), .A2(n1130), .A3(n1110), .ZN(n1252) );
NOR4_X1 U946 ( .A1(n1288), .A2(n1138), .A3(n1099), .A4(n1282), .ZN(n1284) );
INV_X1 U947 ( .A(n1285), .ZN(n1282) );
NAND2_X1 U948 ( .A1(n1141), .A2(n1291), .ZN(n1285) );
NAND4_X1 U949 ( .A1(G902), .A2(G953), .A3(n1292), .A4(n1149), .ZN(n1291) );
INV_X1 U950 ( .A(G900), .ZN(n1149) );
XOR2_X1 U951 ( .A(n1293), .B(n1259), .Z(G24) );
NAND4_X1 U952 ( .A1(n1110), .A2(n1260), .A3(n1111), .A4(n1104), .ZN(n1259) );
AND3_X1 U953 ( .A1(n1099), .A2(n1097), .A3(n1290), .ZN(n1260) );
XNOR2_X1 U954 ( .A(G119), .B(n1176), .ZN(G21) );
NAND4_X1 U955 ( .A1(n1288), .A2(n1136), .A3(n1290), .A4(n1294), .ZN(n1176) );
NOR2_X1 U956 ( .A1(n1267), .A2(n1137), .ZN(n1294) );
INV_X1 U957 ( .A(n1097), .ZN(n1288) );
XOR2_X1 U958 ( .A(n1295), .B(n1258), .Z(G18) );
OR2_X1 U959 ( .A1(n1296), .A2(n1139), .ZN(n1258) );
NAND2_X1 U960 ( .A1(n1283), .A2(n1111), .ZN(n1139) );
INV_X1 U961 ( .A(n1281), .ZN(n1111) );
XOR2_X1 U962 ( .A(G113), .B(n1297), .Z(G15) );
NOR2_X1 U963 ( .A1(n1138), .A2(n1296), .ZN(n1297) );
NAND3_X1 U964 ( .A1(n1110), .A2(n1290), .A3(n1140), .ZN(n1296) );
NOR2_X1 U965 ( .A1(n1136), .A2(n1097), .ZN(n1140) );
INV_X1 U966 ( .A(n1267), .ZN(n1110) );
NAND2_X1 U967 ( .A1(n1124), .A2(n1298), .ZN(n1267) );
NAND2_X1 U968 ( .A1(n1281), .A2(n1104), .ZN(n1138) );
INV_X1 U969 ( .A(n1283), .ZN(n1104) );
XNOR2_X1 U970 ( .A(G110), .B(n1257), .ZN(G12) );
NAND4_X1 U971 ( .A1(n1097), .A2(n1136), .A3(n1290), .A4(n1299), .ZN(n1257) );
NOR2_X1 U972 ( .A1(n1122), .A2(n1137), .ZN(n1299) );
NAND2_X1 U973 ( .A1(n1281), .A2(n1283), .ZN(n1137) );
XOR2_X1 U974 ( .A(n1300), .B(G475), .Z(n1283) );
NAND2_X1 U975 ( .A1(n1203), .A2(n1301), .ZN(n1300) );
XNOR2_X1 U976 ( .A(n1302), .B(n1303), .ZN(n1203) );
NOR2_X1 U977 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
XOR2_X1 U978 ( .A(n1306), .B(KEYINPUT41), .Z(n1305) );
NAND2_X1 U979 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NOR2_X1 U980 ( .A1(n1307), .A2(n1308), .ZN(n1304) );
INV_X1 U981 ( .A(G104), .ZN(n1308) );
AND2_X1 U982 ( .A1(n1309), .A2(n1310), .ZN(n1307) );
NAND2_X1 U983 ( .A1(G122), .A2(n1311), .ZN(n1310) );
XOR2_X1 U984 ( .A(n1312), .B(KEYINPUT30), .Z(n1309) );
NAND2_X1 U985 ( .A1(G113), .A2(n1293), .ZN(n1312) );
NAND2_X1 U986 ( .A1(n1313), .A2(n1314), .ZN(n1302) );
OR2_X1 U987 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XOR2_X1 U988 ( .A(n1317), .B(KEYINPUT61), .Z(n1313) );
NAND2_X1 U989 ( .A1(n1316), .A2(n1315), .ZN(n1317) );
NAND3_X1 U990 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1315) );
NAND2_X1 U991 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
OR3_X1 U992 ( .A1(n1321), .A2(n1322), .A3(KEYINPUT2), .ZN(n1319) );
OR2_X1 U993 ( .A1(n1323), .A2(KEYINPUT12), .ZN(n1321) );
NOR2_X1 U994 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
AND2_X1 U995 ( .A1(n1154), .A2(KEYINPUT42), .ZN(n1325) );
NAND3_X1 U996 ( .A1(n1326), .A2(n1327), .A3(KEYINPUT2), .ZN(n1318) );
INV_X1 U997 ( .A(n1324), .ZN(n1327) );
NOR2_X1 U998 ( .A1(n1328), .A2(KEYINPUT42), .ZN(n1324) );
NAND2_X1 U999 ( .A1(KEYINPUT42), .A2(n1154), .ZN(n1326) );
NAND2_X1 U1000 ( .A1(n1329), .A2(n1330), .ZN(n1154) );
OR2_X1 U1001 ( .A1(n1331), .A2(G125), .ZN(n1330) );
XNOR2_X1 U1002 ( .A(n1332), .B(n1333), .ZN(n1316) );
XOR2_X1 U1003 ( .A(G143), .B(G131), .Z(n1333) );
NAND3_X1 U1004 ( .A1(n1334), .A2(n1091), .A3(G214), .ZN(n1332) );
INV_X1 U1005 ( .A(G237), .ZN(n1334) );
XOR2_X1 U1006 ( .A(n1335), .B(G478), .Z(n1281) );
NAND2_X1 U1007 ( .A1(n1194), .A2(n1301), .ZN(n1335) );
XNOR2_X1 U1008 ( .A(n1336), .B(n1337), .ZN(n1194) );
XOR2_X1 U1009 ( .A(n1338), .B(n1339), .Z(n1337) );
XOR2_X1 U1010 ( .A(G128), .B(G122), .Z(n1339) );
XOR2_X1 U1011 ( .A(G143), .B(G134), .Z(n1338) );
XOR2_X1 U1012 ( .A(n1340), .B(n1341), .Z(n1336) );
XNOR2_X1 U1013 ( .A(n1295), .B(G107), .ZN(n1341) );
NAND2_X1 U1014 ( .A1(n1342), .A2(G217), .ZN(n1340) );
INV_X1 U1015 ( .A(n1262), .ZN(n1122) );
NOR2_X1 U1016 ( .A1(n1124), .A2(n1109), .ZN(n1262) );
INV_X1 U1017 ( .A(n1298), .ZN(n1109) );
NAND2_X1 U1018 ( .A1(G221), .A2(n1343), .ZN(n1298) );
XNOR2_X1 U1019 ( .A(n1108), .B(G469), .ZN(n1124) );
AND3_X1 U1020 ( .A1(n1344), .A2(n1345), .A3(n1301), .ZN(n1108) );
NAND2_X1 U1021 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
XOR2_X1 U1022 ( .A(KEYINPUT19), .B(n1348), .Z(n1346) );
NAND2_X1 U1023 ( .A1(n1349), .A2(n1350), .ZN(n1344) );
INV_X1 U1024 ( .A(n1347), .ZN(n1350) );
XOR2_X1 U1025 ( .A(n1351), .B(n1211), .Z(n1347) );
XOR2_X1 U1026 ( .A(n1352), .B(KEYINPUT49), .Z(n1351) );
NAND3_X1 U1027 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1352) );
NAND2_X1 U1028 ( .A1(n1231), .A2(n1356), .ZN(n1355) );
NAND2_X1 U1029 ( .A1(n1357), .A2(n1358), .ZN(n1354) );
INV_X1 U1030 ( .A(KEYINPUT3), .ZN(n1358) );
NAND2_X1 U1031 ( .A1(n1153), .A2(n1359), .ZN(n1357) );
XOR2_X1 U1032 ( .A(KEYINPUT47), .B(n1360), .Z(n1359) );
INV_X1 U1033 ( .A(n1231), .ZN(n1360) );
NAND2_X1 U1034 ( .A1(KEYINPUT3), .A2(n1361), .ZN(n1353) );
NAND2_X1 U1035 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
NAND2_X1 U1036 ( .A1(KEYINPUT47), .A2(n1231), .ZN(n1363) );
OR3_X1 U1037 ( .A1(n1356), .A2(KEYINPUT47), .A3(n1231), .ZN(n1362) );
INV_X1 U1038 ( .A(n1153), .ZN(n1356) );
XOR2_X1 U1039 ( .A(n1364), .B(G128), .Z(n1153) );
NAND3_X1 U1040 ( .A1(n1365), .A2(n1366), .A3(n1367), .ZN(n1364) );
NAND2_X1 U1041 ( .A1(G143), .A2(n1322), .ZN(n1367) );
NAND2_X1 U1042 ( .A1(KEYINPUT0), .A2(n1368), .ZN(n1366) );
NAND2_X1 U1043 ( .A1(n1369), .A2(n1278), .ZN(n1368) );
XOR2_X1 U1044 ( .A(KEYINPUT9), .B(G146), .Z(n1369) );
NAND2_X1 U1045 ( .A1(n1370), .A2(n1371), .ZN(n1365) );
INV_X1 U1046 ( .A(KEYINPUT0), .ZN(n1371) );
NAND2_X1 U1047 ( .A1(n1372), .A2(n1373), .ZN(n1370) );
NAND2_X1 U1048 ( .A1(KEYINPUT9), .A2(n1322), .ZN(n1373) );
OR3_X1 U1049 ( .A1(G143), .A2(KEYINPUT9), .A3(n1322), .ZN(n1372) );
INV_X1 U1050 ( .A(G146), .ZN(n1322) );
XOR2_X1 U1051 ( .A(KEYINPUT46), .B(n1348), .Z(n1349) );
XNOR2_X1 U1052 ( .A(n1228), .B(n1374), .ZN(n1348) );
NOR2_X1 U1053 ( .A1(KEYINPUT59), .A2(n1227), .ZN(n1374) );
XOR2_X1 U1054 ( .A(G110), .B(n1331), .Z(n1227) );
NAND2_X1 U1055 ( .A1(G227), .A2(n1091), .ZN(n1228) );
AND2_X1 U1056 ( .A1(n1130), .A2(n1264), .ZN(n1290) );
NAND2_X1 U1057 ( .A1(n1141), .A2(n1375), .ZN(n1264) );
NAND3_X1 U1058 ( .A1(n1168), .A2(n1292), .A3(G902), .ZN(n1375) );
NOR2_X1 U1059 ( .A1(n1091), .A2(G898), .ZN(n1168) );
NAND3_X1 U1060 ( .A1(n1292), .A2(n1091), .A3(n1376), .ZN(n1141) );
XOR2_X1 U1061 ( .A(KEYINPUT32), .B(G952), .Z(n1376) );
NAND2_X1 U1062 ( .A1(G237), .A2(G234), .ZN(n1292) );
AND2_X1 U1063 ( .A1(n1377), .A2(n1128), .ZN(n1130) );
XNOR2_X1 U1064 ( .A(n1378), .B(n1379), .ZN(n1128) );
NOR2_X1 U1065 ( .A1(n1380), .A2(n1239), .ZN(n1379) );
XOR2_X1 U1066 ( .A(n1381), .B(KEYINPUT55), .Z(n1380) );
NAND3_X1 U1067 ( .A1(n1382), .A2(n1301), .A3(n1383), .ZN(n1378) );
XOR2_X1 U1068 ( .A(KEYINPUT24), .B(n1384), .Z(n1383) );
NOR2_X1 U1069 ( .A1(n1385), .A2(n1235), .ZN(n1384) );
NAND2_X1 U1070 ( .A1(n1385), .A2(n1235), .ZN(n1382) );
NAND2_X1 U1071 ( .A1(n1386), .A2(n1387), .ZN(n1235) );
NAND2_X1 U1072 ( .A1(n1179), .A2(n1388), .ZN(n1387) );
NAND2_X1 U1073 ( .A1(n1185), .A2(n1186), .ZN(n1388) );
OR2_X1 U1074 ( .A1(n1389), .A2(n1231), .ZN(n1186) );
NAND2_X1 U1075 ( .A1(n1389), .A2(n1231), .ZN(n1185) );
NAND2_X1 U1076 ( .A1(n1390), .A2(n1181), .ZN(n1386) );
INV_X1 U1077 ( .A(n1179), .ZN(n1181) );
XOR2_X1 U1078 ( .A(n1391), .B(n1392), .Z(n1179) );
XOR2_X1 U1079 ( .A(KEYINPUT7), .B(G110), .Z(n1392) );
NAND2_X1 U1080 ( .A1(KEYINPUT5), .A2(n1293), .ZN(n1391) );
INV_X1 U1081 ( .A(G122), .ZN(n1293) );
XOR2_X1 U1082 ( .A(n1231), .B(n1389), .Z(n1390) );
XOR2_X1 U1083 ( .A(n1393), .B(n1394), .Z(n1389) );
XNOR2_X1 U1084 ( .A(n1295), .B(n1395), .ZN(n1394) );
NOR2_X1 U1085 ( .A1(KEYINPUT14), .A2(n1311), .ZN(n1395) );
INV_X1 U1086 ( .A(G113), .ZN(n1311) );
XNOR2_X1 U1087 ( .A(G119), .B(KEYINPUT21), .ZN(n1393) );
XNOR2_X1 U1088 ( .A(G101), .B(n1396), .ZN(n1231) );
XOR2_X1 U1089 ( .A(G107), .B(G104), .Z(n1396) );
XNOR2_X1 U1090 ( .A(n1238), .B(n1397), .ZN(n1385) );
XOR2_X1 U1091 ( .A(n1274), .B(n1273), .Z(n1397) );
NAND2_X1 U1092 ( .A1(G224), .A2(n1091), .ZN(n1274) );
XNOR2_X1 U1093 ( .A(n1328), .B(KEYINPUT62), .ZN(n1238) );
INV_X1 U1094 ( .A(G125), .ZN(n1328) );
XOR2_X1 U1095 ( .A(n1129), .B(KEYINPUT27), .Z(n1377) );
NAND2_X1 U1096 ( .A1(G214), .A2(n1381), .ZN(n1129) );
NAND2_X1 U1097 ( .A1(n1398), .A2(n1301), .ZN(n1381) );
XOR2_X1 U1098 ( .A(KEYINPUT31), .B(G237), .Z(n1398) );
INV_X1 U1099 ( .A(n1099), .ZN(n1136) );
XNOR2_X1 U1100 ( .A(n1399), .B(n1191), .ZN(n1099) );
NAND2_X1 U1101 ( .A1(G217), .A2(n1343), .ZN(n1191) );
NAND2_X1 U1102 ( .A1(G234), .A2(n1301), .ZN(n1343) );
NAND2_X1 U1103 ( .A1(n1189), .A2(n1301), .ZN(n1399) );
XNOR2_X1 U1104 ( .A(n1400), .B(n1401), .ZN(n1189) );
XNOR2_X1 U1105 ( .A(n1402), .B(n1403), .ZN(n1401) );
XOR2_X1 U1106 ( .A(n1404), .B(n1405), .Z(n1403) );
NOR2_X1 U1107 ( .A1(KEYINPUT45), .A2(n1406), .ZN(n1405) );
NAND3_X1 U1108 ( .A1(n1407), .A2(n1408), .A3(n1329), .ZN(n1404) );
NAND2_X1 U1109 ( .A1(G125), .A2(n1331), .ZN(n1329) );
OR3_X1 U1110 ( .A1(n1331), .A2(G125), .A3(KEYINPUT50), .ZN(n1408) );
XNOR2_X1 U1111 ( .A(G140), .B(KEYINPUT11), .ZN(n1331) );
NAND2_X1 U1112 ( .A1(KEYINPUT50), .A2(G125), .ZN(n1407) );
XOR2_X1 U1113 ( .A(n1409), .B(n1410), .Z(n1400) );
XOR2_X1 U1114 ( .A(G146), .B(G119), .Z(n1410) );
XOR2_X1 U1115 ( .A(n1411), .B(G110), .Z(n1409) );
NAND2_X1 U1116 ( .A1(n1342), .A2(G221), .ZN(n1411) );
AND2_X1 U1117 ( .A1(G234), .A2(n1091), .ZN(n1342) );
INV_X1 U1118 ( .A(G953), .ZN(n1091) );
XOR2_X1 U1119 ( .A(n1412), .B(G472), .Z(n1097) );
NAND2_X1 U1120 ( .A1(n1413), .A2(n1301), .ZN(n1412) );
INV_X1 U1121 ( .A(G902), .ZN(n1301) );
XOR2_X1 U1122 ( .A(n1414), .B(n1415), .Z(n1413) );
XOR2_X1 U1123 ( .A(n1416), .B(n1220), .Z(n1415) );
NOR3_X1 U1124 ( .A1(G237), .A2(G953), .A3(n1239), .ZN(n1220) );
INV_X1 U1125 ( .A(G210), .ZN(n1239) );
NAND2_X1 U1126 ( .A1(n1417), .A2(n1418), .ZN(n1416) );
NAND2_X1 U1127 ( .A1(n1212), .A2(n1419), .ZN(n1418) );
NAND2_X1 U1128 ( .A1(n1211), .A2(n1420), .ZN(n1417) );
XNOR2_X1 U1129 ( .A(n1212), .B(KEYINPUT1), .ZN(n1420) );
XNOR2_X1 U1130 ( .A(n1273), .B(n1421), .ZN(n1212) );
XOR2_X1 U1131 ( .A(G113), .B(n1422), .Z(n1421) );
NOR2_X1 U1132 ( .A1(KEYINPUT13), .A2(n1423), .ZN(n1422) );
NOR3_X1 U1133 ( .A1(n1424), .A2(n1425), .A3(n1426), .ZN(n1423) );
AND2_X1 U1134 ( .A1(n1427), .A2(G119), .ZN(n1426) );
NOR3_X1 U1135 ( .A1(G119), .A2(KEYINPUT15), .A3(n1427), .ZN(n1425) );
NAND2_X1 U1136 ( .A1(KEYINPUT6), .A2(n1295), .ZN(n1427) );
INV_X1 U1137 ( .A(G116), .ZN(n1295) );
AND2_X1 U1138 ( .A1(G116), .A2(KEYINPUT15), .ZN(n1424) );
XOR2_X1 U1139 ( .A(n1406), .B(n1428), .Z(n1273) );
NOR2_X1 U1140 ( .A1(KEYINPUT22), .A2(n1429), .ZN(n1428) );
XOR2_X1 U1141 ( .A(n1278), .B(G146), .Z(n1429) );
INV_X1 U1142 ( .A(G143), .ZN(n1278) );
INV_X1 U1143 ( .A(G128), .ZN(n1406) );
INV_X1 U1144 ( .A(n1419), .ZN(n1211) );
XOR2_X1 U1145 ( .A(n1157), .B(n1430), .Z(n1419) );
NOR2_X1 U1146 ( .A1(KEYINPUT39), .A2(n1152), .ZN(n1430) );
XNOR2_X1 U1147 ( .A(G134), .B(n1402), .ZN(n1152) );
XOR2_X1 U1148 ( .A(G137), .B(KEYINPUT25), .Z(n1402) );
INV_X1 U1149 ( .A(G131), .ZN(n1157) );
XOR2_X1 U1150 ( .A(n1431), .B(G101), .Z(n1414) );
XNOR2_X1 U1151 ( .A(KEYINPUT60), .B(KEYINPUT18), .ZN(n1431) );
endmodule


