//Key = 0101110110000100010101111001100101111010101110101111011101011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350;

XNOR2_X1 U738 ( .A(G107), .B(n1020), .ZN(G9) );
NAND4_X1 U739 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(G75) );
NAND4_X1 U740 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1023) );
NOR3_X1 U741 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
XNOR2_X1 U742 ( .A(n1032), .B(n1033), .ZN(n1031) );
NAND2_X1 U743 ( .A1(KEYINPUT36), .A2(n1034), .ZN(n1033) );
NAND3_X1 U744 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1029) );
XNOR2_X1 U745 ( .A(G478), .B(n1038), .ZN(n1037) );
NAND2_X1 U746 ( .A1(KEYINPUT56), .A2(n1039), .ZN(n1036) );
OR3_X1 U747 ( .A1(n1040), .A2(KEYINPUT56), .A3(n1039), .ZN(n1035) );
NOR3_X1 U748 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1027) );
XNOR2_X1 U749 ( .A(G469), .B(n1044), .ZN(n1026) );
NAND2_X1 U750 ( .A1(KEYINPUT4), .A2(n1045), .ZN(n1044) );
XNOR2_X1 U751 ( .A(n1046), .B(n1047), .ZN(n1025) );
NOR2_X1 U752 ( .A1(KEYINPUT2), .A2(n1048), .ZN(n1047) );
XNOR2_X1 U753 ( .A(n1049), .B(KEYINPUT35), .ZN(n1048) );
NAND2_X1 U754 ( .A1(n1050), .A2(n1051), .ZN(n1022) );
NAND2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND4_X1 U756 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1053) );
NAND2_X1 U757 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NAND2_X1 U758 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1058) );
NAND2_X1 U761 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U762 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND3_X1 U763 ( .A1(n1060), .A2(n1070), .A3(n1064), .ZN(n1052) );
NAND3_X1 U764 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1070) );
NAND2_X1 U765 ( .A1(n1055), .A2(n1074), .ZN(n1073) );
NAND3_X1 U766 ( .A1(n1075), .A2(n1076), .A3(n1054), .ZN(n1071) );
NAND2_X1 U767 ( .A1(n1043), .A2(n1077), .ZN(n1076) );
NAND2_X1 U768 ( .A1(n1078), .A2(n1057), .ZN(n1075) );
NAND2_X1 U769 ( .A1(n1041), .A2(n1079), .ZN(n1078) );
INV_X1 U770 ( .A(n1080), .ZN(n1050) );
XOR2_X1 U771 ( .A(n1081), .B(n1082), .Z(G72) );
NOR2_X1 U772 ( .A1(n1083), .A2(n1024), .ZN(n1082) );
AND2_X1 U773 ( .A1(G227), .A2(G900), .ZN(n1083) );
NAND2_X1 U774 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
NAND2_X1 U775 ( .A1(n1086), .A2(n1024), .ZN(n1085) );
XOR2_X1 U776 ( .A(n1087), .B(n1088), .Z(n1086) );
NAND3_X1 U777 ( .A1(G900), .A2(n1088), .A3(G953), .ZN(n1084) );
XNOR2_X1 U778 ( .A(n1089), .B(n1090), .ZN(n1088) );
XNOR2_X1 U779 ( .A(KEYINPUT52), .B(n1091), .ZN(n1089) );
NOR3_X1 U780 ( .A1(KEYINPUT20), .A2(n1092), .A3(n1093), .ZN(n1091) );
NOR2_X1 U781 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NOR2_X1 U782 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U783 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U784 ( .A1(n1100), .A2(n1101), .ZN(n1096) );
NOR2_X1 U785 ( .A1(G128), .A2(n1102), .ZN(n1092) );
NOR2_X1 U786 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U787 ( .A1(n1101), .A2(n1099), .ZN(n1104) );
XOR2_X1 U788 ( .A(n1105), .B(KEYINPUT18), .Z(n1099) );
NOR2_X1 U789 ( .A1(n1098), .A2(n1100), .ZN(n1103) );
XNOR2_X1 U790 ( .A(n1105), .B(KEYINPUT63), .ZN(n1100) );
XOR2_X1 U791 ( .A(n1106), .B(G131), .Z(n1105) );
NAND2_X1 U792 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U793 ( .A1(G137), .A2(n1109), .ZN(n1108) );
XOR2_X1 U794 ( .A(KEYINPUT62), .B(n1110), .Z(n1107) );
NOR2_X1 U795 ( .A1(G137), .A2(n1109), .ZN(n1110) );
XOR2_X1 U796 ( .A(KEYINPUT61), .B(G134), .Z(n1109) );
NAND2_X1 U797 ( .A1(n1111), .A2(n1112), .ZN(G69) );
NAND2_X1 U798 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND2_X1 U799 ( .A1(G953), .A2(n1115), .ZN(n1113) );
NAND2_X1 U800 ( .A1(G898), .A2(G224), .ZN(n1115) );
NAND2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1111) );
NAND2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U803 ( .A1(G953), .A2(n1120), .ZN(n1119) );
INV_X1 U804 ( .A(n1121), .ZN(n1118) );
INV_X1 U805 ( .A(n1114), .ZN(n1116) );
NAND2_X1 U806 ( .A1(n1122), .A2(n1123), .ZN(n1114) );
NAND3_X1 U807 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
NAND2_X1 U808 ( .A1(G953), .A2(n1127), .ZN(n1125) );
NAND2_X1 U809 ( .A1(n1128), .A2(n1024), .ZN(n1124) );
NAND2_X1 U810 ( .A1(n1129), .A2(n1127), .ZN(n1128) );
XOR2_X1 U811 ( .A(KEYINPUT49), .B(n1130), .Z(n1122) );
NOR3_X1 U812 ( .A1(n1129), .A2(n1121), .A3(n1131), .ZN(n1130) );
AND2_X1 U813 ( .A1(n1127), .A2(n1126), .ZN(n1131) );
INV_X1 U814 ( .A(KEYINPUT41), .ZN(n1127) );
XNOR2_X1 U815 ( .A(n1132), .B(n1133), .ZN(n1129) );
XOR2_X1 U816 ( .A(KEYINPUT42), .B(KEYINPUT32), .Z(n1133) );
XNOR2_X1 U817 ( .A(n1134), .B(n1135), .ZN(n1132) );
NOR2_X1 U818 ( .A1(n1136), .A2(n1137), .ZN(G66) );
NOR3_X1 U819 ( .A1(n1032), .A2(n1138), .A3(n1139), .ZN(n1137) );
AND3_X1 U820 ( .A1(n1140), .A2(n1034), .A3(n1141), .ZN(n1139) );
INV_X1 U821 ( .A(n1142), .ZN(n1034) );
NOR2_X1 U822 ( .A1(n1143), .A2(n1140), .ZN(n1138) );
NOR2_X1 U823 ( .A1(n1021), .A2(n1142), .ZN(n1143) );
NOR2_X1 U824 ( .A1(n1136), .A2(n1144), .ZN(G63) );
NOR3_X1 U825 ( .A1(n1038), .A2(n1145), .A3(n1146), .ZN(n1144) );
NOR3_X1 U826 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1146) );
NOR2_X1 U827 ( .A1(n1150), .A2(n1151), .ZN(n1145) );
NOR2_X1 U828 ( .A1(n1021), .A2(n1148), .ZN(n1150) );
XOR2_X1 U829 ( .A(G478), .B(KEYINPUT57), .Z(n1148) );
NOR2_X1 U830 ( .A1(n1136), .A2(n1152), .ZN(G60) );
NOR3_X1 U831 ( .A1(n1049), .A2(n1153), .A3(n1154), .ZN(n1152) );
AND3_X1 U832 ( .A1(n1155), .A2(G475), .A3(n1141), .ZN(n1154) );
NOR2_X1 U833 ( .A1(n1156), .A2(n1155), .ZN(n1153) );
NOR2_X1 U834 ( .A1(n1021), .A2(n1046), .ZN(n1156) );
XNOR2_X1 U835 ( .A(G104), .B(n1157), .ZN(G6) );
NAND3_X1 U836 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1157) );
XOR2_X1 U837 ( .A(KEYINPUT47), .B(n1060), .Z(n1159) );
NOR3_X1 U838 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(G57) );
AND3_X1 U839 ( .A1(KEYINPUT11), .A2(G953), .A3(G952), .ZN(n1163) );
NOR2_X1 U840 ( .A1(KEYINPUT11), .A2(n1164), .ZN(n1162) );
INV_X1 U841 ( .A(n1136), .ZN(n1164) );
NOR3_X1 U842 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1161) );
NOR2_X1 U843 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
INV_X1 U844 ( .A(n1170), .ZN(n1169) );
NOR2_X1 U845 ( .A1(KEYINPUT26), .A2(n1171), .ZN(n1168) );
XOR2_X1 U846 ( .A(KEYINPUT58), .B(n1172), .Z(n1171) );
NOR3_X1 U847 ( .A1(n1170), .A2(KEYINPUT26), .A3(n1172), .ZN(n1166) );
XNOR2_X1 U848 ( .A(n1173), .B(n1174), .ZN(n1170) );
NAND2_X1 U849 ( .A1(KEYINPUT17), .A2(n1175), .ZN(n1173) );
AND2_X1 U850 ( .A1(n1172), .A2(KEYINPUT26), .ZN(n1165) );
AND2_X1 U851 ( .A1(n1176), .A2(n1177), .ZN(n1172) );
NAND2_X1 U852 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND2_X1 U853 ( .A1(n1141), .A2(G472), .ZN(n1179) );
INV_X1 U854 ( .A(n1180), .ZN(n1178) );
NAND3_X1 U855 ( .A1(n1141), .A2(G472), .A3(n1180), .ZN(n1176) );
XNOR2_X1 U856 ( .A(n1181), .B(n1182), .ZN(n1180) );
XOR2_X1 U857 ( .A(KEYINPUT15), .B(n1183), .Z(n1182) );
NOR2_X1 U858 ( .A1(n1136), .A2(n1184), .ZN(G54) );
XOR2_X1 U859 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U860 ( .A(n1187), .B(n1188), .Z(n1186) );
NOR2_X1 U861 ( .A1(n1189), .A2(n1149), .ZN(n1188) );
NAND2_X1 U862 ( .A1(KEYINPUT55), .A2(n1190), .ZN(n1187) );
XNOR2_X1 U863 ( .A(G140), .B(n1191), .ZN(n1190) );
NAND2_X1 U864 ( .A1(KEYINPUT8), .A2(n1192), .ZN(n1191) );
XOR2_X1 U865 ( .A(n1193), .B(n1194), .Z(n1185) );
NOR2_X1 U866 ( .A1(KEYINPUT14), .A2(n1195), .ZN(n1194) );
XOR2_X1 U867 ( .A(n1196), .B(n1197), .Z(n1195) );
NAND2_X1 U868 ( .A1(KEYINPUT50), .A2(n1198), .ZN(n1196) );
NOR2_X1 U869 ( .A1(n1136), .A2(n1199), .ZN(G51) );
NOR2_X1 U870 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U871 ( .A(n1202), .B(KEYINPUT28), .Z(n1201) );
NAND2_X1 U872 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NOR2_X1 U873 ( .A1(n1203), .A2(n1204), .ZN(n1200) );
NOR2_X1 U874 ( .A1(n1149), .A2(n1039), .ZN(n1203) );
INV_X1 U875 ( .A(n1141), .ZN(n1149) );
NOR2_X1 U876 ( .A1(n1205), .A2(n1021), .ZN(n1141) );
NOR2_X1 U877 ( .A1(n1126), .A2(n1087), .ZN(n1021) );
NAND4_X1 U878 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1087) );
NOR3_X1 U879 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1209) );
AND4_X1 U880 ( .A1(n1213), .A2(KEYINPUT45), .A3(n1160), .A4(n1214), .ZN(n1212) );
NOR2_X1 U881 ( .A1(n1215), .A2(n1213), .ZN(n1211) );
NOR3_X1 U882 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
NOR2_X1 U883 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NOR2_X1 U884 ( .A1(n1221), .A2(n1222), .ZN(n1219) );
NOR2_X1 U885 ( .A1(KEYINPUT45), .A2(n1062), .ZN(n1221) );
INV_X1 U886 ( .A(n1160), .ZN(n1062) );
NOR2_X1 U887 ( .A1(n1077), .A2(n1223), .ZN(n1216) );
NOR2_X1 U888 ( .A1(n1072), .A2(n1223), .ZN(n1210) );
NAND4_X1 U889 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1126) );
AND4_X1 U890 ( .A1(n1020), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1227) );
NAND3_X1 U891 ( .A1(n1158), .A2(n1222), .A3(n1060), .ZN(n1020) );
NAND2_X1 U892 ( .A1(n1074), .A2(n1231), .ZN(n1226) );
NAND2_X1 U893 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NAND3_X1 U894 ( .A1(n1234), .A2(n1222), .A3(n1235), .ZN(n1233) );
NAND3_X1 U895 ( .A1(n1060), .A2(n1158), .A3(n1160), .ZN(n1224) );
NOR2_X1 U896 ( .A1(n1024), .A2(G952), .ZN(n1136) );
XNOR2_X1 U897 ( .A(G146), .B(n1236), .ZN(G48) );
NAND2_X1 U898 ( .A1(n1237), .A2(n1160), .ZN(n1236) );
XOR2_X1 U899 ( .A(n1238), .B(n1239), .Z(G45) );
NAND2_X1 U900 ( .A1(KEYINPUT51), .A2(G143), .ZN(n1239) );
NAND2_X1 U901 ( .A1(n1240), .A2(n1074), .ZN(n1238) );
XNOR2_X1 U902 ( .A(n1217), .B(KEYINPUT33), .ZN(n1240) );
AND4_X1 U903 ( .A1(n1241), .A2(n1235), .A3(n1242), .A4(n1243), .ZN(n1217) );
NOR2_X1 U904 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
NAND2_X1 U905 ( .A1(n1246), .A2(n1247), .ZN(G42) );
NAND4_X1 U906 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1247) );
NAND2_X1 U907 ( .A1(KEYINPUT10), .A2(n1252), .ZN(n1251) );
NAND2_X1 U908 ( .A1(KEYINPUT43), .A2(G140), .ZN(n1250) );
INV_X1 U909 ( .A(n1072), .ZN(n1249) );
INV_X1 U910 ( .A(n1223), .ZN(n1248) );
NAND3_X1 U911 ( .A1(G140), .A2(n1253), .A3(KEYINPUT43), .ZN(n1246) );
OR3_X1 U912 ( .A1(n1072), .A2(KEYINPUT10), .A3(n1223), .ZN(n1253) );
XOR2_X1 U913 ( .A(n1208), .B(n1254), .Z(G39) );
NAND2_X1 U914 ( .A1(KEYINPUT38), .A2(G137), .ZN(n1254) );
NAND4_X1 U915 ( .A1(n1214), .A2(n1054), .A3(n1064), .A4(n1057), .ZN(n1208) );
INV_X1 U916 ( .A(n1220), .ZN(n1214) );
XNOR2_X1 U917 ( .A(G134), .B(n1206), .ZN(G36) );
NAND2_X1 U918 ( .A1(n1255), .A2(n1222), .ZN(n1206) );
XOR2_X1 U919 ( .A(n1207), .B(n1256), .Z(G33) );
NAND2_X1 U920 ( .A1(KEYINPUT21), .A2(G131), .ZN(n1256) );
NAND2_X1 U921 ( .A1(n1255), .A2(n1160), .ZN(n1207) );
NOR3_X1 U922 ( .A1(n1066), .A2(n1244), .A3(n1072), .ZN(n1255) );
NAND3_X1 U923 ( .A1(n1243), .A2(n1057), .A3(n1054), .ZN(n1072) );
INV_X1 U924 ( .A(n1257), .ZN(n1244) );
INV_X1 U925 ( .A(n1235), .ZN(n1066) );
XNOR2_X1 U926 ( .A(G128), .B(n1258), .ZN(G30) );
NAND3_X1 U927 ( .A1(n1237), .A2(n1222), .A3(KEYINPUT48), .ZN(n1258) );
INV_X1 U928 ( .A(n1063), .ZN(n1222) );
NOR2_X1 U929 ( .A1(n1220), .A2(n1213), .ZN(n1237) );
NAND4_X1 U930 ( .A1(n1243), .A2(n1030), .A3(n1257), .A4(n1069), .ZN(n1220) );
XNOR2_X1 U931 ( .A(G101), .B(n1225), .ZN(G3) );
NAND3_X1 U932 ( .A1(n1064), .A2(n1158), .A3(n1235), .ZN(n1225) );
XNOR2_X1 U933 ( .A(n1259), .B(n1260), .ZN(G27) );
NOR3_X1 U934 ( .A1(n1223), .A2(n1261), .A3(n1213), .ZN(n1260) );
XNOR2_X1 U935 ( .A(n1055), .B(KEYINPUT12), .ZN(n1261) );
NAND4_X1 U936 ( .A1(n1068), .A2(n1160), .A3(n1257), .A4(n1069), .ZN(n1223) );
NAND2_X1 U937 ( .A1(n1080), .A2(n1262), .ZN(n1257) );
NAND4_X1 U938 ( .A1(G953), .A2(G902), .A3(n1263), .A4(n1264), .ZN(n1262) );
INV_X1 U939 ( .A(G900), .ZN(n1264) );
XNOR2_X1 U940 ( .A(G122), .B(n1265), .ZN(G24) );
NAND2_X1 U941 ( .A1(n1266), .A2(n1074), .ZN(n1265) );
XOR2_X1 U942 ( .A(n1232), .B(KEYINPUT40), .Z(n1266) );
NAND4_X1 U943 ( .A1(n1234), .A2(n1060), .A3(n1241), .A4(n1267), .ZN(n1232) );
NOR2_X1 U944 ( .A1(n1069), .A2(n1030), .ZN(n1060) );
XOR2_X1 U945 ( .A(n1230), .B(n1268), .Z(G21) );
XNOR2_X1 U946 ( .A(KEYINPUT19), .B(n1269), .ZN(n1268) );
NAND3_X1 U947 ( .A1(n1234), .A2(n1064), .A3(n1270), .ZN(n1230) );
AND3_X1 U948 ( .A1(n1074), .A2(n1069), .A3(n1030), .ZN(n1270) );
XNOR2_X1 U949 ( .A(G116), .B(n1271), .ZN(G18) );
NAND4_X1 U950 ( .A1(KEYINPUT27), .A2(n1235), .A3(n1272), .A4(n1234), .ZN(n1271) );
NOR2_X1 U951 ( .A1(n1213), .A2(n1063), .ZN(n1272) );
NAND2_X1 U952 ( .A1(n1241), .A2(n1245), .ZN(n1063) );
XOR2_X1 U953 ( .A(G113), .B(n1273), .Z(G15) );
NOR2_X1 U954 ( .A1(KEYINPUT37), .A2(n1229), .ZN(n1273) );
NAND4_X1 U955 ( .A1(n1160), .A2(n1235), .A3(n1234), .A4(n1274), .ZN(n1229) );
AND2_X1 U956 ( .A1(n1055), .A2(n1275), .ZN(n1234) );
INV_X1 U957 ( .A(n1077), .ZN(n1055) );
NAND2_X1 U958 ( .A1(n1079), .A2(n1276), .ZN(n1077) );
NOR2_X1 U959 ( .A1(n1069), .A2(n1068), .ZN(n1235) );
NOR2_X1 U960 ( .A1(n1245), .A2(n1241), .ZN(n1160) );
INV_X1 U961 ( .A(n1267), .ZN(n1245) );
XNOR2_X1 U962 ( .A(G110), .B(n1228), .ZN(G12) );
NAND4_X1 U963 ( .A1(n1064), .A2(n1158), .A3(n1068), .A4(n1069), .ZN(n1228) );
NAND2_X1 U964 ( .A1(n1277), .A2(n1278), .ZN(n1069) );
NAND2_X1 U965 ( .A1(n1032), .A2(n1279), .ZN(n1278) );
XOR2_X1 U966 ( .A(KEYINPUT1), .B(n1280), .Z(n1277) );
NOR2_X1 U967 ( .A1(n1032), .A2(n1279), .ZN(n1280) );
XNOR2_X1 U968 ( .A(KEYINPUT7), .B(n1142), .ZN(n1279) );
NAND2_X1 U969 ( .A1(G217), .A2(n1281), .ZN(n1142) );
NOR2_X1 U970 ( .A1(n1140), .A2(G902), .ZN(n1032) );
XOR2_X1 U971 ( .A(n1282), .B(n1283), .Z(n1140) );
XOR2_X1 U972 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U973 ( .A(n1286), .B(n1287), .ZN(n1285) );
NAND2_X1 U974 ( .A1(KEYINPUT31), .A2(n1192), .ZN(n1287) );
INV_X1 U975 ( .A(G110), .ZN(n1192) );
NAND2_X1 U976 ( .A1(KEYINPUT23), .A2(G128), .ZN(n1286) );
XOR2_X1 U977 ( .A(n1288), .B(n1289), .Z(n1284) );
AND3_X1 U978 ( .A1(G234), .A2(n1024), .A3(G221), .ZN(n1289) );
NAND2_X1 U979 ( .A1(KEYINPUT13), .A2(n1259), .ZN(n1288) );
XOR2_X1 U980 ( .A(n1290), .B(n1291), .Z(n1282) );
XNOR2_X1 U981 ( .A(G146), .B(n1252), .ZN(n1291) );
XNOR2_X1 U982 ( .A(G119), .B(G137), .ZN(n1290) );
INV_X1 U983 ( .A(n1030), .ZN(n1068) );
XNOR2_X1 U984 ( .A(n1292), .B(G472), .ZN(n1030) );
NAND2_X1 U985 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U986 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U987 ( .A(n1297), .B(n1181), .Z(n1296) );
XOR2_X1 U988 ( .A(n1298), .B(n1198), .Z(n1181) );
XOR2_X1 U989 ( .A(n1299), .B(KEYINPUT22), .Z(n1298) );
NAND2_X1 U990 ( .A1(KEYINPUT54), .A2(n1183), .ZN(n1297) );
XNOR2_X1 U991 ( .A(n1175), .B(n1174), .ZN(n1295) );
AND3_X1 U992 ( .A1(n1300), .A2(n1024), .A3(G210), .ZN(n1174) );
XNOR2_X1 U993 ( .A(KEYINPUT53), .B(n1205), .ZN(n1293) );
AND3_X1 U994 ( .A1(n1274), .A2(n1275), .A3(n1243), .ZN(n1158) );
NOR2_X1 U995 ( .A1(n1079), .A2(n1041), .ZN(n1243) );
INV_X1 U996 ( .A(n1276), .ZN(n1041) );
NAND2_X1 U997 ( .A1(G221), .A2(n1281), .ZN(n1276) );
NAND2_X1 U998 ( .A1(G234), .A2(n1205), .ZN(n1281) );
XNOR2_X1 U999 ( .A(n1045), .B(n1189), .ZN(n1079) );
INV_X1 U1000 ( .A(G469), .ZN(n1189) );
NAND2_X1 U1001 ( .A1(n1301), .A2(n1205), .ZN(n1045) );
XOR2_X1 U1002 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U1003 ( .A(n1197), .B(n1198), .ZN(n1303) );
XNOR2_X1 U1004 ( .A(n1304), .B(G131), .ZN(n1198) );
NAND2_X1 U1005 ( .A1(KEYINPUT3), .A2(n1305), .ZN(n1304) );
XOR2_X1 U1006 ( .A(G137), .B(G134), .Z(n1305) );
XOR2_X1 U1007 ( .A(n1306), .B(n1307), .Z(n1197) );
XNOR2_X1 U1008 ( .A(n1175), .B(n1308), .ZN(n1307) );
INV_X1 U1009 ( .A(G101), .ZN(n1175) );
XOR2_X1 U1010 ( .A(n1193), .B(n1309), .Z(n1302) );
XNOR2_X1 U1011 ( .A(n1252), .B(G110), .ZN(n1309) );
INV_X1 U1012 ( .A(G140), .ZN(n1252) );
NAND2_X1 U1013 ( .A1(G227), .A2(n1024), .ZN(n1193) );
NAND2_X1 U1014 ( .A1(n1080), .A2(n1310), .ZN(n1275) );
NAND3_X1 U1015 ( .A1(G902), .A2(n1263), .A3(n1121), .ZN(n1310) );
NOR2_X1 U1016 ( .A1(n1024), .A2(G898), .ZN(n1121) );
NAND3_X1 U1017 ( .A1(n1263), .A2(n1024), .A3(G952), .ZN(n1080) );
NAND2_X1 U1018 ( .A1(G237), .A2(G234), .ZN(n1263) );
XNOR2_X1 U1019 ( .A(n1213), .B(KEYINPUT16), .ZN(n1274) );
INV_X1 U1020 ( .A(n1074), .ZN(n1213) );
NOR2_X1 U1021 ( .A1(n1054), .A2(n1043), .ZN(n1074) );
INV_X1 U1022 ( .A(n1057), .ZN(n1043) );
NAND2_X1 U1023 ( .A1(G214), .A2(n1311), .ZN(n1057) );
NOR2_X1 U1024 ( .A1(n1042), .A2(n1312), .ZN(n1054) );
NOR2_X1 U1025 ( .A1(n1039), .A2(n1040), .ZN(n1312) );
AND2_X1 U1026 ( .A1(n1040), .A2(n1039), .ZN(n1042) );
NAND2_X1 U1027 ( .A1(G210), .A2(n1311), .ZN(n1039) );
NAND2_X1 U1028 ( .A1(n1300), .A2(n1205), .ZN(n1311) );
INV_X1 U1029 ( .A(G902), .ZN(n1205) );
NOR2_X1 U1030 ( .A1(n1204), .A2(G902), .ZN(n1040) );
XOR2_X1 U1031 ( .A(n1313), .B(n1314), .Z(n1204) );
XOR2_X1 U1032 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1033 ( .A(n1259), .B(n1317), .ZN(n1316) );
NOR2_X1 U1034 ( .A1(G953), .A2(n1120), .ZN(n1317) );
INV_X1 U1035 ( .A(G224), .ZN(n1120) );
XOR2_X1 U1036 ( .A(KEYINPUT6), .B(KEYINPUT29), .Z(n1315) );
XOR2_X1 U1037 ( .A(n1318), .B(n1183), .Z(n1313) );
XNOR2_X1 U1038 ( .A(n1319), .B(n1098), .ZN(n1183) );
NAND2_X1 U1039 ( .A1(KEYINPUT46), .A2(n1094), .ZN(n1319) );
XNOR2_X1 U1040 ( .A(n1320), .B(n1321), .ZN(n1318) );
INV_X1 U1041 ( .A(n1134), .ZN(n1321) );
XNOR2_X1 U1042 ( .A(n1299), .B(n1322), .ZN(n1134) );
XNOR2_X1 U1043 ( .A(G110), .B(n1323), .ZN(n1322) );
NAND2_X1 U1044 ( .A1(KEYINPUT34), .A2(n1324), .ZN(n1323) );
XNOR2_X1 U1045 ( .A(G113), .B(n1325), .ZN(n1299) );
XNOR2_X1 U1046 ( .A(n1269), .B(G116), .ZN(n1325) );
INV_X1 U1047 ( .A(G119), .ZN(n1269) );
NAND2_X1 U1048 ( .A1(KEYINPUT5), .A2(n1135), .ZN(n1320) );
XNOR2_X1 U1049 ( .A(n1326), .B(G101), .ZN(n1135) );
NAND3_X1 U1050 ( .A1(n1327), .A2(n1328), .A3(KEYINPUT44), .ZN(n1326) );
NAND2_X1 U1051 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XNOR2_X1 U1052 ( .A(G104), .B(G107), .ZN(n1329) );
OR3_X1 U1053 ( .A1(n1331), .A2(G107), .A3(n1330), .ZN(n1327) );
INV_X1 U1054 ( .A(KEYINPUT9), .ZN(n1330) );
NOR2_X1 U1055 ( .A1(n1267), .A2(n1241), .ZN(n1064) );
XNOR2_X1 U1056 ( .A(n1038), .B(n1332), .ZN(n1241) );
NOR2_X1 U1057 ( .A1(G478), .A2(KEYINPUT39), .ZN(n1332) );
NOR2_X1 U1058 ( .A1(n1151), .A2(G902), .ZN(n1038) );
INV_X1 U1059 ( .A(n1147), .ZN(n1151) );
XNOR2_X1 U1060 ( .A(n1333), .B(n1334), .ZN(n1147) );
AND3_X1 U1061 ( .A1(G217), .A2(n1024), .A3(G234), .ZN(n1334) );
NAND2_X1 U1062 ( .A1(n1335), .A2(KEYINPUT24), .ZN(n1333) );
XOR2_X1 U1063 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1064 ( .A(n1338), .B(n1306), .Z(n1337) );
XNOR2_X1 U1065 ( .A(G107), .B(n1094), .ZN(n1306) );
INV_X1 U1066 ( .A(G128), .ZN(n1094) );
NOR2_X1 U1067 ( .A1(G143), .A2(KEYINPUT25), .ZN(n1338) );
XNOR2_X1 U1068 ( .A(G116), .B(n1339), .ZN(n1336) );
XNOR2_X1 U1069 ( .A(G134), .B(n1324), .ZN(n1339) );
XOR2_X1 U1070 ( .A(n1049), .B(n1340), .Z(n1267) );
XNOR2_X1 U1071 ( .A(KEYINPUT0), .B(n1046), .ZN(n1340) );
INV_X1 U1072 ( .A(G475), .ZN(n1046) );
NOR2_X1 U1073 ( .A1(n1155), .A2(G902), .ZN(n1049) );
XOR2_X1 U1074 ( .A(n1341), .B(n1342), .Z(n1155) );
XOR2_X1 U1075 ( .A(n1308), .B(n1343), .Z(n1342) );
XOR2_X1 U1076 ( .A(n1344), .B(n1090), .Z(n1343) );
XNOR2_X1 U1077 ( .A(n1259), .B(G140), .ZN(n1090) );
INV_X1 U1078 ( .A(G125), .ZN(n1259) );
AND3_X1 U1079 ( .A1(G214), .A2(n1024), .A3(n1300), .ZN(n1344) );
INV_X1 U1080 ( .A(G237), .ZN(n1300) );
INV_X1 U1081 ( .A(G953), .ZN(n1024) );
XNOR2_X1 U1082 ( .A(n1331), .B(n1098), .ZN(n1308) );
INV_X1 U1083 ( .A(n1101), .ZN(n1098) );
XNOR2_X1 U1084 ( .A(G143), .B(G146), .ZN(n1101) );
INV_X1 U1085 ( .A(G104), .ZN(n1331) );
XOR2_X1 U1086 ( .A(n1345), .B(n1346), .Z(n1341) );
XOR2_X1 U1087 ( .A(KEYINPUT60), .B(KEYINPUT30), .Z(n1346) );
XOR2_X1 U1088 ( .A(n1347), .B(G131), .Z(n1345) );
NAND2_X1 U1089 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
NAND2_X1 U1090 ( .A1(G113), .A2(n1324), .ZN(n1349) );
XOR2_X1 U1091 ( .A(KEYINPUT59), .B(n1350), .Z(n1348) );
NOR2_X1 U1092 ( .A1(G113), .A2(n1324), .ZN(n1350) );
INV_X1 U1093 ( .A(G122), .ZN(n1324) );
endmodule


