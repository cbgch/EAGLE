//Key = 1010110101011100000011001000001011010000100100000010000000010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306;

XNOR2_X1 U719 ( .A(n997), .B(n998), .ZN(G9) );
XOR2_X1 U720 ( .A(KEYINPUT39), .B(G107), .Z(n998) );
NOR2_X1 U721 ( .A1(n999), .A2(n1000), .ZN(G75) );
XOR2_X1 U722 ( .A(n1001), .B(KEYINPUT40), .Z(n1000) );
NAND4_X1 U723 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n1001) );
NOR2_X1 U724 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
XOR2_X1 U725 ( .A(KEYINPUT55), .B(n1008), .Z(n1007) );
NOR3_X1 U726 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1008) );
INV_X1 U727 ( .A(n1012), .ZN(n1004) );
NAND4_X1 U728 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1003) );
NAND2_X1 U729 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND3_X1 U730 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NAND2_X1 U731 ( .A1(n1022), .A2(n1023), .ZN(n1002) );
NAND3_X1 U732 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
NAND2_X1 U733 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
INV_X1 U734 ( .A(KEYINPUT59), .ZN(n1028) );
NAND4_X1 U735 ( .A1(n1029), .A2(n1013), .A3(n1014), .A4(n1019), .ZN(n1027) );
NAND3_X1 U736 ( .A1(n1014), .A2(n1030), .A3(n1013), .ZN(n1025) );
NAND2_X1 U737 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U738 ( .A1(n1033), .A2(n1015), .ZN(n1032) );
XOR2_X1 U739 ( .A(n1034), .B(n1035), .Z(n1033) );
NAND2_X1 U740 ( .A1(n1019), .A2(n1036), .ZN(n1031) );
NAND2_X1 U741 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U742 ( .A1(KEYINPUT59), .A2(n1029), .ZN(n1038) );
OR2_X1 U743 ( .A1(n1010), .A2(n1039), .ZN(n1024) );
NAND3_X1 U744 ( .A1(n1019), .A2(n1015), .A3(n1014), .ZN(n1010) );
INV_X1 U745 ( .A(n1040), .ZN(n1014) );
NOR2_X1 U746 ( .A1(G952), .A2(n1012), .ZN(n999) );
NAND2_X1 U747 ( .A1(n1041), .A2(n1042), .ZN(n1012) );
NAND4_X1 U748 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
NOR4_X1 U749 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
XOR2_X1 U750 ( .A(n1051), .B(n1052), .Z(n1050) );
XOR2_X1 U751 ( .A(n1053), .B(n1054), .Z(n1049) );
NOR2_X1 U752 ( .A1(n1055), .A2(n1056), .ZN(n1045) );
XNOR2_X1 U753 ( .A(n1057), .B(n1058), .ZN(n1056) );
NAND2_X1 U754 ( .A1(KEYINPUT30), .A2(n1059), .ZN(n1057) );
XOR2_X1 U755 ( .A(n1060), .B(n1061), .Z(n1055) );
NOR2_X1 U756 ( .A1(n1062), .A2(KEYINPUT51), .ZN(n1061) );
XOR2_X1 U757 ( .A(n1063), .B(KEYINPUT58), .Z(n1060) );
XOR2_X1 U758 ( .A(n1064), .B(n1065), .Z(G72) );
NOR2_X1 U759 ( .A1(n1066), .A2(n1041), .ZN(n1065) );
AND2_X1 U760 ( .A1(G227), .A2(G900), .ZN(n1066) );
NOR3_X1 U761 ( .A1(KEYINPUT37), .A2(n1067), .A3(n1068), .ZN(n1064) );
NOR2_X1 U762 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XNOR2_X1 U763 ( .A(KEYINPUT48), .B(n1071), .ZN(n1070) );
NOR2_X1 U764 ( .A1(n1072), .A2(n1071), .ZN(n1067) );
NAND2_X1 U765 ( .A1(n1041), .A2(n1073), .ZN(n1071) );
INV_X1 U766 ( .A(n1069), .ZN(n1072) );
NOR2_X1 U767 ( .A1(n1074), .A2(n1075), .ZN(n1069) );
XNOR2_X1 U768 ( .A(n1076), .B(n1077), .ZN(n1074) );
XOR2_X1 U769 ( .A(n1078), .B(n1079), .Z(n1077) );
NAND2_X1 U770 ( .A1(n1080), .A2(KEYINPUT32), .ZN(n1078) );
XOR2_X1 U771 ( .A(n1081), .B(G143), .Z(n1080) );
XOR2_X1 U772 ( .A(G140), .B(G125), .Z(n1076) );
XOR2_X1 U773 ( .A(n1082), .B(n1083), .Z(G69) );
NOR3_X1 U774 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1083) );
NOR2_X1 U775 ( .A1(G898), .A2(n1087), .ZN(n1086) );
NOR2_X1 U776 ( .A1(n1088), .A2(n1089), .ZN(n1085) );
XOR2_X1 U777 ( .A(KEYINPUT61), .B(n1090), .Z(n1084) );
AND2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(n1090) );
XNOR2_X1 U779 ( .A(n1091), .B(n1092), .ZN(n1089) );
NAND2_X1 U780 ( .A1(KEYINPUT9), .A2(n1093), .ZN(n1091) );
XOR2_X1 U781 ( .A(n1094), .B(n1095), .Z(n1082) );
NOR2_X1 U782 ( .A1(KEYINPUT14), .A2(n1096), .ZN(n1095) );
NOR2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U784 ( .A(KEYINPUT27), .B(G953), .Z(n1098) );
NOR3_X1 U785 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1097) );
XOR2_X1 U786 ( .A(KEYINPUT3), .B(n1102), .Z(n1099) );
NAND2_X1 U787 ( .A1(G953), .A2(n1103), .ZN(n1094) );
NAND2_X1 U788 ( .A1(G224), .A2(n1104), .ZN(n1103) );
XOR2_X1 U789 ( .A(KEYINPUT38), .B(G898), .Z(n1104) );
NOR2_X1 U790 ( .A1(n1105), .A2(n1106), .ZN(G66) );
XOR2_X1 U791 ( .A(n1107), .B(n1108), .Z(n1106) );
XNOR2_X1 U792 ( .A(KEYINPUT28), .B(n1109), .ZN(n1108) );
NOR2_X1 U793 ( .A1(n1058), .A2(n1110), .ZN(n1107) );
NOR2_X1 U794 ( .A1(n1111), .A2(n1112), .ZN(G63) );
XNOR2_X1 U795 ( .A(n1113), .B(n1114), .ZN(n1112) );
XOR2_X1 U796 ( .A(KEYINPUT44), .B(n1115), .Z(n1114) );
NOR2_X1 U797 ( .A1(n1051), .A2(n1110), .ZN(n1115) );
INV_X1 U798 ( .A(G478), .ZN(n1051) );
NOR2_X1 U799 ( .A1(G952), .A2(n1116), .ZN(n1111) );
XOR2_X1 U800 ( .A(n1041), .B(KEYINPUT22), .Z(n1116) );
NOR2_X1 U801 ( .A1(n1105), .A2(n1117), .ZN(G60) );
XNOR2_X1 U802 ( .A(n1118), .B(n1119), .ZN(n1117) );
NOR2_X1 U803 ( .A1(n1120), .A2(n1110), .ZN(n1119) );
INV_X1 U804 ( .A(G475), .ZN(n1120) );
XNOR2_X1 U805 ( .A(G104), .B(n1121), .ZN(G6) );
NOR2_X1 U806 ( .A1(n1105), .A2(n1122), .ZN(G57) );
XOR2_X1 U807 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U808 ( .A(n1079), .B(n1125), .Z(n1124) );
XNOR2_X1 U809 ( .A(n1126), .B(n1127), .ZN(n1123) );
XOR2_X1 U810 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U811 ( .A1(n1130), .A2(n1110), .ZN(n1129) );
INV_X1 U812 ( .A(G472), .ZN(n1130) );
NOR2_X1 U813 ( .A1(KEYINPUT17), .A2(n1131), .ZN(n1128) );
XOR2_X1 U814 ( .A(n1132), .B(G101), .Z(n1131) );
NOR2_X1 U815 ( .A1(n1105), .A2(n1133), .ZN(G54) );
XOR2_X1 U816 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U817 ( .A(n1136), .B(n1137), .Z(n1135) );
NOR2_X1 U818 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR3_X1 U819 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
XOR2_X1 U820 ( .A(G101), .B(n1143), .Z(n1142) );
INV_X1 U821 ( .A(KEYINPUT41), .ZN(n1140) );
NOR2_X1 U822 ( .A1(KEYINPUT41), .A2(n1144), .ZN(n1138) );
XNOR2_X1 U823 ( .A(n1145), .B(n1143), .ZN(n1144) );
XNOR2_X1 U824 ( .A(n1081), .B(n1146), .ZN(n1143) );
XOR2_X1 U825 ( .A(G104), .B(n1147), .Z(n1146) );
XOR2_X1 U826 ( .A(n1148), .B(n1149), .Z(n1081) );
INV_X1 U827 ( .A(G146), .ZN(n1148) );
NOR2_X1 U828 ( .A1(n1053), .A2(n1110), .ZN(n1136) );
INV_X1 U829 ( .A(G469), .ZN(n1053) );
XOR2_X1 U830 ( .A(n1150), .B(n1151), .Z(n1134) );
NOR2_X1 U831 ( .A1(KEYINPUT23), .A2(n1152), .ZN(n1151) );
XOR2_X1 U832 ( .A(KEYINPUT54), .B(G110), .Z(n1152) );
XOR2_X1 U833 ( .A(n1153), .B(n1154), .Z(n1150) );
INV_X1 U834 ( .A(G140), .ZN(n1153) );
NOR2_X1 U835 ( .A1(n1105), .A2(n1155), .ZN(G51) );
XOR2_X1 U836 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U837 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U838 ( .A1(n1110), .A2(n1160), .ZN(n1158) );
NAND2_X1 U839 ( .A1(n1161), .A2(n1006), .ZN(n1110) );
OR4_X1 U840 ( .A1(n1101), .A2(n1073), .A3(n1100), .A4(n1102), .ZN(n1006) );
NAND4_X1 U841 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1100) );
NAND4_X1 U842 ( .A1(n1166), .A2(n1167), .A3(n1029), .A4(n1168), .ZN(n1163) );
NAND2_X1 U843 ( .A1(n1169), .A2(n1170), .ZN(n1162) );
XOR2_X1 U844 ( .A(n1171), .B(KEYINPUT20), .Z(n1169) );
NAND4_X1 U845 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1073) );
AND4_X1 U846 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1175) );
NAND2_X1 U847 ( .A1(n1180), .A2(n1181), .ZN(n1174) );
NAND4_X1 U848 ( .A1(n1166), .A2(n1167), .A3(n1182), .A4(n1183), .ZN(n1173) );
NAND2_X1 U849 ( .A1(n1184), .A2(n1185), .ZN(n1172) );
NAND2_X1 U850 ( .A1(n1186), .A2(n1037), .ZN(n1185) );
XOR2_X1 U851 ( .A(n1187), .B(KEYINPUT62), .Z(n1186) );
NAND3_X1 U852 ( .A1(n1188), .A2(n997), .A3(n1121), .ZN(n1101) );
NAND3_X1 U853 ( .A1(n1189), .A2(n1015), .A3(n1167), .ZN(n1121) );
NAND3_X1 U854 ( .A1(n1190), .A2(n1015), .A3(n1189), .ZN(n997) );
XOR2_X1 U855 ( .A(KEYINPUT45), .B(G902), .Z(n1161) );
NOR2_X1 U856 ( .A1(n1191), .A2(n1192), .ZN(n1156) );
NOR2_X1 U857 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XOR2_X1 U858 ( .A(KEYINPUT24), .B(n1195), .Z(n1194) );
NOR2_X1 U859 ( .A1(G125), .A2(n1195), .ZN(n1191) );
NOR2_X1 U860 ( .A1(n1041), .A2(G952), .ZN(n1105) );
XOR2_X1 U861 ( .A(G146), .B(n1196), .Z(G48) );
NOR2_X1 U862 ( .A1(n1171), .A2(n1197), .ZN(n1196) );
XOR2_X1 U863 ( .A(KEYINPUT2), .B(n1180), .Z(n1197) );
AND2_X1 U864 ( .A1(n1198), .A2(n1167), .ZN(n1180) );
XOR2_X1 U865 ( .A(n1199), .B(n1179), .Z(G45) );
NAND4_X1 U866 ( .A1(n1181), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1179) );
NOR2_X1 U867 ( .A1(n1187), .A2(n1203), .ZN(n1202) );
XOR2_X1 U868 ( .A(G140), .B(n1204), .Z(G42) );
NOR2_X1 U869 ( .A1(n1037), .A2(n1205), .ZN(n1204) );
XNOR2_X1 U870 ( .A(G137), .B(n1178), .ZN(G39) );
NAND3_X1 U871 ( .A1(n1022), .A2(n1013), .A3(n1198), .ZN(n1178) );
INV_X1 U872 ( .A(n1011), .ZN(n1022) );
XNOR2_X1 U873 ( .A(n1177), .B(n1206), .ZN(G36) );
NOR2_X1 U874 ( .A1(KEYINPUT34), .A2(n1207), .ZN(n1206) );
OR4_X1 U875 ( .A1(n1203), .A2(n1011), .A3(n1187), .A4(n1039), .ZN(n1177) );
XOR2_X1 U876 ( .A(G131), .B(n1208), .Z(G33) );
NOR2_X1 U877 ( .A1(n1187), .A2(n1205), .ZN(n1208) );
INV_X1 U878 ( .A(n1184), .ZN(n1205) );
NOR3_X1 U879 ( .A1(n1009), .A2(n1011), .A3(n1203), .ZN(n1184) );
NAND2_X1 U880 ( .A1(n1020), .A2(n1044), .ZN(n1011) );
XOR2_X1 U881 ( .A(n1209), .B(n1176), .Z(G30) );
NAND3_X1 U882 ( .A1(n1190), .A2(n1181), .A3(n1198), .ZN(n1176) );
NOR3_X1 U883 ( .A1(n1210), .A2(n1211), .A3(n1203), .ZN(n1198) );
NAND3_X1 U884 ( .A1(n1183), .A2(n1043), .A3(n1035), .ZN(n1203) );
XOR2_X1 U885 ( .A(G101), .B(n1102), .Z(G3) );
AND3_X1 U886 ( .A1(n1013), .A2(n1189), .A3(n1029), .ZN(n1102) );
XOR2_X1 U887 ( .A(n1193), .B(n1212), .Z(G27) );
NAND4_X1 U888 ( .A1(n1213), .A2(n1166), .A3(n1182), .A4(n1183), .ZN(n1212) );
NAND2_X1 U889 ( .A1(n1040), .A2(n1214), .ZN(n1183) );
NAND3_X1 U890 ( .A1(G902), .A2(n1215), .A3(n1075), .ZN(n1214) );
NOR2_X1 U891 ( .A1(n1087), .A2(G900), .ZN(n1075) );
XOR2_X1 U892 ( .A(n1009), .B(KEYINPUT21), .Z(n1213) );
XOR2_X1 U893 ( .A(n1164), .B(n1216), .Z(G24) );
XNOR2_X1 U894 ( .A(G122), .B(KEYINPUT47), .ZN(n1216) );
NAND3_X1 U895 ( .A1(n1166), .A2(n1015), .A3(n1217), .ZN(n1164) );
NOR3_X1 U896 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1217) );
NOR2_X1 U897 ( .A1(n1047), .A2(n1221), .ZN(n1015) );
XOR2_X1 U898 ( .A(G119), .B(n1222), .Z(G21) );
NOR2_X1 U899 ( .A1(n1223), .A2(n1171), .ZN(n1222) );
XNOR2_X1 U900 ( .A(n1170), .B(KEYINPUT56), .ZN(n1223) );
AND3_X1 U901 ( .A1(n1221), .A2(n1013), .A3(n1224), .ZN(n1170) );
NOR3_X1 U902 ( .A1(n1225), .A2(n1219), .A3(n1211), .ZN(n1224) );
XNOR2_X1 U903 ( .A(G116), .B(n1165), .ZN(G18) );
NAND4_X1 U904 ( .A1(n1166), .A2(n1029), .A3(n1190), .A4(n1168), .ZN(n1165) );
INV_X1 U905 ( .A(n1039), .ZN(n1190) );
NAND2_X1 U906 ( .A1(n1220), .A2(n1201), .ZN(n1039) );
INV_X1 U907 ( .A(n1187), .ZN(n1029) );
INV_X1 U908 ( .A(n1017), .ZN(n1166) );
NAND2_X1 U909 ( .A1(n1019), .A2(n1181), .ZN(n1017) );
XNOR2_X1 U910 ( .A(G113), .B(n1226), .ZN(G15) );
NAND3_X1 U911 ( .A1(n1227), .A2(n1167), .A3(n1228), .ZN(n1226) );
NOR3_X1 U912 ( .A1(n1187), .A2(n1219), .A3(n1225), .ZN(n1228) );
INV_X1 U913 ( .A(n1019), .ZN(n1225) );
NOR2_X1 U914 ( .A1(n1035), .A2(n1034), .ZN(n1019) );
INV_X1 U915 ( .A(n1043), .ZN(n1034) );
INV_X1 U916 ( .A(n1168), .ZN(n1219) );
NAND2_X1 U917 ( .A1(n1210), .A2(n1047), .ZN(n1187) );
INV_X1 U918 ( .A(n1211), .ZN(n1047) );
INV_X1 U919 ( .A(n1221), .ZN(n1210) );
INV_X1 U920 ( .A(n1009), .ZN(n1167) );
NAND2_X1 U921 ( .A1(n1218), .A2(n1200), .ZN(n1009) );
INV_X1 U922 ( .A(n1201), .ZN(n1218) );
XOR2_X1 U923 ( .A(n1171), .B(KEYINPUT33), .Z(n1227) );
INV_X1 U924 ( .A(n1181), .ZN(n1171) );
XNOR2_X1 U925 ( .A(G110), .B(n1188), .ZN(G12) );
NAND3_X1 U926 ( .A1(n1013), .A2(n1189), .A3(n1182), .ZN(n1188) );
INV_X1 U927 ( .A(n1037), .ZN(n1182) );
NAND2_X1 U928 ( .A1(n1221), .A2(n1211), .ZN(n1037) );
XOR2_X1 U929 ( .A(n1229), .B(G472), .Z(n1211) );
NAND2_X1 U930 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U931 ( .A(n1232), .B(n1233), .Z(n1230) );
XNOR2_X1 U932 ( .A(n1132), .B(n1234), .ZN(n1233) );
NOR2_X1 U933 ( .A1(KEYINPUT60), .A2(n1126), .ZN(n1234) );
XOR2_X1 U934 ( .A(n1235), .B(n1236), .Z(n1126) );
NOR2_X1 U935 ( .A1(G113), .A2(KEYINPUT26), .ZN(n1236) );
NAND3_X1 U936 ( .A1(n1237), .A2(n1041), .A3(G210), .ZN(n1132) );
XOR2_X1 U937 ( .A(n1145), .B(n1125), .Z(n1232) );
XNOR2_X1 U938 ( .A(n1238), .B(n1058), .ZN(n1221) );
NAND2_X1 U939 ( .A1(G217), .A2(n1239), .ZN(n1058) );
NAND2_X1 U940 ( .A1(KEYINPUT11), .A2(n1059), .ZN(n1238) );
NAND2_X1 U941 ( .A1(n1109), .A2(n1231), .ZN(n1059) );
NAND2_X1 U942 ( .A1(n1240), .A2(n1241), .ZN(n1109) );
NAND2_X1 U943 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U944 ( .A(n1244), .B(n1245), .Z(n1243) );
XOR2_X1 U945 ( .A(n1246), .B(KEYINPUT53), .Z(n1242) );
NAND2_X1 U946 ( .A1(n1247), .A2(n1248), .ZN(n1240) );
XNOR2_X1 U947 ( .A(n1245), .B(n1244), .ZN(n1248) );
NAND2_X1 U948 ( .A1(n1249), .A2(G221), .ZN(n1244) );
NOR2_X1 U949 ( .A1(KEYINPUT49), .A2(n1250), .ZN(n1245) );
XOR2_X1 U950 ( .A(n1246), .B(KEYINPUT50), .Z(n1247) );
XOR2_X1 U951 ( .A(n1251), .B(n1252), .Z(n1246) );
XNOR2_X1 U952 ( .A(n1253), .B(n1254), .ZN(n1251) );
NOR2_X1 U953 ( .A1(KEYINPUT6), .A2(n1193), .ZN(n1254) );
INV_X1 U954 ( .A(G125), .ZN(n1193) );
NOR2_X1 U955 ( .A1(KEYINPUT42), .A2(n1255), .ZN(n1253) );
XOR2_X1 U956 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U957 ( .A(G119), .B(G110), .Z(n1257) );
XOR2_X1 U958 ( .A(KEYINPUT5), .B(G128), .Z(n1256) );
AND4_X1 U959 ( .A1(n1035), .A2(n1181), .A3(n1168), .A4(n1043), .ZN(n1189) );
NAND2_X1 U960 ( .A1(G221), .A2(n1239), .ZN(n1043) );
NAND2_X1 U961 ( .A1(n1258), .A2(n1231), .ZN(n1239) );
NAND2_X1 U962 ( .A1(n1040), .A2(n1259), .ZN(n1168) );
OR4_X1 U963 ( .A1(n1087), .A2(n1231), .A3(n1260), .A4(G898), .ZN(n1259) );
INV_X1 U964 ( .A(n1215), .ZN(n1260) );
XNOR2_X1 U965 ( .A(n1041), .B(KEYINPUT43), .ZN(n1087) );
NAND3_X1 U966 ( .A1(n1215), .A2(n1041), .A3(G952), .ZN(n1040) );
NAND2_X1 U967 ( .A1(G237), .A2(n1258), .ZN(n1215) );
XOR2_X1 U968 ( .A(G234), .B(KEYINPUT19), .Z(n1258) );
NOR2_X1 U969 ( .A1(n1020), .A2(n1021), .ZN(n1181) );
INV_X1 U970 ( .A(n1044), .ZN(n1021) );
NAND2_X1 U971 ( .A1(G214), .A2(n1261), .ZN(n1044) );
XNOR2_X1 U972 ( .A(n1063), .B(n1262), .ZN(n1020) );
NOR2_X1 U973 ( .A1(n1062), .A2(KEYINPUT16), .ZN(n1262) );
INV_X1 U974 ( .A(n1160), .ZN(n1062) );
NAND2_X1 U975 ( .A1(G210), .A2(n1261), .ZN(n1160) );
NAND2_X1 U976 ( .A1(n1237), .A2(n1231), .ZN(n1261) );
NAND2_X1 U977 ( .A1(n1263), .A2(n1231), .ZN(n1063) );
XOR2_X1 U978 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U979 ( .A(KEYINPUT46), .B(G125), .Z(n1265) );
XNOR2_X1 U980 ( .A(n1159), .B(n1195), .ZN(n1264) );
XNOR2_X1 U981 ( .A(n1125), .B(n1266), .ZN(n1195) );
AND2_X1 U982 ( .A1(n1041), .A2(G224), .ZN(n1266) );
XNOR2_X1 U983 ( .A(n1149), .B(n1267), .ZN(n1125) );
NOR2_X1 U984 ( .A1(KEYINPUT36), .A2(n1268), .ZN(n1267) );
XOR2_X1 U985 ( .A(G146), .B(G143), .Z(n1268) );
XOR2_X1 U986 ( .A(n1269), .B(n1093), .Z(n1159) );
XOR2_X1 U987 ( .A(n1270), .B(n1235), .Z(n1093) );
XOR2_X1 U988 ( .A(G116), .B(G119), .Z(n1235) );
XNOR2_X1 U989 ( .A(KEYINPUT7), .B(n1271), .ZN(n1270) );
NOR2_X1 U990 ( .A1(G113), .A2(KEYINPUT25), .ZN(n1271) );
XOR2_X1 U991 ( .A(n1272), .B(n1088), .Z(n1269) );
XOR2_X1 U992 ( .A(G110), .B(n1273), .Z(n1088) );
NAND2_X1 U993 ( .A1(KEYINPUT0), .A2(n1092), .ZN(n1272) );
XNOR2_X1 U994 ( .A(n1274), .B(G101), .ZN(n1092) );
NAND2_X1 U995 ( .A1(KEYINPUT12), .A2(n1275), .ZN(n1274) );
XOR2_X1 U996 ( .A(G107), .B(G104), .Z(n1275) );
XOR2_X1 U997 ( .A(n1276), .B(G469), .Z(n1035) );
NAND2_X1 U998 ( .A1(KEYINPUT13), .A2(n1054), .ZN(n1276) );
NAND2_X1 U999 ( .A1(n1277), .A2(n1231), .ZN(n1054) );
XOR2_X1 U1000 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U1001 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U1002 ( .A(n1282), .B(n1149), .Z(n1281) );
XNOR2_X1 U1003 ( .A(n1209), .B(KEYINPUT31), .ZN(n1149) );
INV_X1 U1004 ( .A(G128), .ZN(n1209) );
INV_X1 U1005 ( .A(n1147), .ZN(n1282) );
XOR2_X1 U1006 ( .A(n1145), .B(n1283), .Z(n1278) );
XOR2_X1 U1007 ( .A(G110), .B(n1154), .Z(n1283) );
AND2_X1 U1008 ( .A1(G227), .A2(n1041), .ZN(n1154) );
XOR2_X1 U1009 ( .A(G101), .B(n1141), .Z(n1145) );
INV_X1 U1010 ( .A(n1079), .ZN(n1141) );
XOR2_X1 U1011 ( .A(n1284), .B(n1250), .Z(n1079) );
XOR2_X1 U1012 ( .A(G137), .B(KEYINPUT57), .Z(n1250) );
XOR2_X1 U1013 ( .A(n1207), .B(G131), .Z(n1284) );
NOR2_X1 U1014 ( .A1(n1200), .A2(n1201), .ZN(n1013) );
XOR2_X1 U1015 ( .A(n1052), .B(n1285), .Z(n1201) );
NOR2_X1 U1016 ( .A1(G478), .A2(KEYINPUT29), .ZN(n1285) );
NAND2_X1 U1017 ( .A1(n1113), .A2(n1231), .ZN(n1052) );
XNOR2_X1 U1018 ( .A(n1286), .B(n1287), .ZN(n1113) );
XOR2_X1 U1019 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U1020 ( .A(n1207), .B(G128), .Z(n1289) );
INV_X1 U1021 ( .A(G134), .ZN(n1207) );
NAND2_X1 U1022 ( .A1(G217), .A2(n1249), .ZN(n1288) );
AND2_X1 U1023 ( .A1(G234), .A2(n1041), .ZN(n1249) );
XOR2_X1 U1024 ( .A(n1290), .B(n1273), .Z(n1286) );
XOR2_X1 U1025 ( .A(n1291), .B(n1147), .Z(n1290) );
XOR2_X1 U1026 ( .A(G107), .B(G143), .Z(n1147) );
NAND2_X1 U1027 ( .A1(KEYINPUT4), .A2(G116), .ZN(n1291) );
INV_X1 U1028 ( .A(n1220), .ZN(n1200) );
XOR2_X1 U1029 ( .A(n1292), .B(n1048), .Z(n1220) );
XNOR2_X1 U1030 ( .A(n1293), .B(n1294), .ZN(n1048) );
XOR2_X1 U1031 ( .A(KEYINPUT52), .B(G475), .Z(n1294) );
NAND2_X1 U1032 ( .A1(n1118), .A2(n1231), .ZN(n1293) );
INV_X1 U1033 ( .A(G902), .ZN(n1231) );
XNOR2_X1 U1034 ( .A(n1295), .B(n1296), .ZN(n1118) );
XOR2_X1 U1035 ( .A(n1273), .B(n1297), .Z(n1296) );
INV_X1 U1036 ( .A(n1280), .ZN(n1297) );
XNOR2_X1 U1037 ( .A(G104), .B(n1252), .ZN(n1280) );
XOR2_X1 U1038 ( .A(G140), .B(G146), .Z(n1252) );
XOR2_X1 U1039 ( .A(G122), .B(KEYINPUT1), .Z(n1273) );
XOR2_X1 U1040 ( .A(n1298), .B(n1299), .Z(n1295) );
XOR2_X1 U1041 ( .A(G113), .B(n1300), .Z(n1299) );
NOR2_X1 U1042 ( .A1(KEYINPUT18), .A2(n1301), .ZN(n1300) );
XOR2_X1 U1043 ( .A(KEYINPUT63), .B(G125), .Z(n1301) );
NAND2_X1 U1044 ( .A1(n1302), .A2(n1303), .ZN(n1298) );
NAND2_X1 U1045 ( .A1(n1304), .A2(G131), .ZN(n1303) );
XOR2_X1 U1046 ( .A(n1305), .B(KEYINPUT15), .Z(n1302) );
OR2_X1 U1047 ( .A1(n1304), .A2(G131), .ZN(n1305) );
XNOR2_X1 U1048 ( .A(n1306), .B(n1199), .ZN(n1304) );
INV_X1 U1049 ( .A(G143), .ZN(n1199) );
NAND4_X1 U1050 ( .A1(KEYINPUT35), .A2(G214), .A3(n1237), .A4(n1041), .ZN(n1306) );
INV_X1 U1051 ( .A(G953), .ZN(n1041) );
INV_X1 U1052 ( .A(G237), .ZN(n1237) );
XNOR2_X1 U1053 ( .A(KEYINPUT8), .B(KEYINPUT10), .ZN(n1292) );
endmodule


