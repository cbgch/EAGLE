//Key = 1100101010001011011111111000001100010000110100101100100010010110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364;

XNOR2_X1 U757 ( .A(G107), .B(n1044), .ZN(G9) );
NOR2_X1 U758 ( .A1(n1045), .A2(n1046), .ZN(G75) );
NOR4_X1 U759 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
NOR2_X1 U760 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U761 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
XOR2_X1 U762 ( .A(KEYINPUT7), .B(n1055), .Z(n1054) );
AND3_X1 U763 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NOR2_X1 U764 ( .A1(n1059), .A2(n1060), .ZN(n1053) );
NOR2_X1 U765 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR3_X1 U766 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
NOR3_X1 U767 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1064) );
AND3_X1 U768 ( .A1(n1069), .A2(n1070), .A3(KEYINPUT58), .ZN(n1068) );
NOR2_X1 U769 ( .A1(n1071), .A2(n1069), .ZN(n1067) );
NOR2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U771 ( .A1(KEYINPUT58), .A2(n1074), .ZN(n1072) );
NOR2_X1 U772 ( .A1(n1075), .A2(n1076), .ZN(n1066) );
NOR4_X1 U773 ( .A1(n1077), .A2(n1078), .A3(n1076), .A4(n1069), .ZN(n1061) );
NOR2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR3_X1 U775 ( .A1(n1065), .A2(n1081), .A3(n1082), .ZN(n1077) );
NOR2_X1 U776 ( .A1(KEYINPUT17), .A2(n1063), .ZN(n1081) );
XOR2_X1 U777 ( .A(KEYINPUT14), .B(n1083), .Z(n1048) );
NAND3_X1 U778 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1047) );
NAND3_X1 U779 ( .A1(n1087), .A2(n1088), .A3(n1057), .ZN(n1086) );
NOR4_X1 U780 ( .A1(n1060), .A2(n1076), .A3(n1065), .A4(n1063), .ZN(n1057) );
NAND2_X1 U781 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND3_X1 U782 ( .A1(n1091), .A2(n1092), .A3(KEYINPUT17), .ZN(n1090) );
NOR3_X1 U783 ( .A1(n1093), .A2(G953), .A3(G952), .ZN(n1045) );
INV_X1 U784 ( .A(n1084), .ZN(n1093) );
NAND3_X1 U785 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1084) );
NOR3_X1 U786 ( .A1(n1097), .A2(n1092), .A3(n1056), .ZN(n1096) );
XOR2_X1 U787 ( .A(n1058), .B(KEYINPUT22), .Z(n1097) );
XOR2_X1 U788 ( .A(n1098), .B(KEYINPUT24), .Z(n1095) );
NAND4_X1 U789 ( .A1(n1099), .A2(n1080), .A3(n1100), .A4(n1079), .ZN(n1098) );
NOR2_X1 U790 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
AND2_X1 U791 ( .A1(n1103), .A2(G478), .ZN(n1102) );
XOR2_X1 U792 ( .A(n1091), .B(KEYINPUT27), .Z(n1094) );
XOR2_X1 U793 ( .A(n1104), .B(n1105), .Z(G72) );
XOR2_X1 U794 ( .A(n1106), .B(n1107), .Z(n1105) );
NAND2_X1 U795 ( .A1(G953), .A2(n1108), .ZN(n1107) );
NAND2_X1 U796 ( .A1(G900), .A2(G227), .ZN(n1108) );
NAND2_X1 U797 ( .A1(n1109), .A2(n1110), .ZN(n1106) );
NAND2_X1 U798 ( .A1(G953), .A2(n1111), .ZN(n1110) );
XOR2_X1 U799 ( .A(n1112), .B(n1113), .Z(n1109) );
XNOR2_X1 U800 ( .A(n1114), .B(n1115), .ZN(n1113) );
XOR2_X1 U801 ( .A(n1116), .B(KEYINPUT21), .Z(n1112) );
NAND3_X1 U802 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1116) );
NAND2_X1 U803 ( .A1(KEYINPUT30), .A2(n1120), .ZN(n1118) );
NAND2_X1 U804 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U805 ( .A1(n1123), .A2(n1124), .ZN(n1117) );
INV_X1 U806 ( .A(KEYINPUT30), .ZN(n1124) );
XNOR2_X1 U807 ( .A(n1125), .B(n1126), .ZN(n1123) );
NOR2_X1 U808 ( .A1(G134), .A2(n1127), .ZN(n1126) );
NOR2_X1 U809 ( .A1(n1083), .A2(G953), .ZN(n1104) );
XOR2_X1 U810 ( .A(n1128), .B(n1129), .Z(G69) );
XOR2_X1 U811 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U812 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XOR2_X1 U813 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U814 ( .A1(KEYINPUT56), .A2(n1136), .ZN(n1134) );
XOR2_X1 U815 ( .A(KEYINPUT18), .B(n1137), .Z(n1136) );
NOR2_X1 U816 ( .A1(n1138), .A2(n1085), .ZN(n1132) );
XNOR2_X1 U817 ( .A(G898), .B(KEYINPUT4), .ZN(n1138) );
NAND2_X1 U818 ( .A1(n1085), .A2(n1139), .ZN(n1130) );
NAND3_X1 U819 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
XNOR2_X1 U820 ( .A(KEYINPUT19), .B(n1044), .ZN(n1140) );
NAND2_X1 U821 ( .A1(G953), .A2(n1143), .ZN(n1128) );
NAND2_X1 U822 ( .A1(G898), .A2(G224), .ZN(n1143) );
NOR2_X1 U823 ( .A1(n1144), .A2(n1145), .ZN(G66) );
XOR2_X1 U824 ( .A(KEYINPUT2), .B(n1146), .Z(n1145) );
NOR2_X1 U825 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U826 ( .A(KEYINPUT36), .B(n1149), .Z(n1148) );
AND2_X1 U827 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NOR2_X1 U828 ( .A1(n1151), .A2(n1150), .ZN(n1147) );
NAND3_X1 U829 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1150) );
XNOR2_X1 U830 ( .A(G902), .B(KEYINPUT23), .ZN(n1154) );
XNOR2_X1 U831 ( .A(n1155), .B(KEYINPUT48), .ZN(n1151) );
NOR2_X1 U832 ( .A1(n1144), .A2(n1156), .ZN(G63) );
XNOR2_X1 U833 ( .A(n1157), .B(n1158), .ZN(n1156) );
NOR3_X1 U834 ( .A1(n1159), .A2(KEYINPUT54), .A3(n1160), .ZN(n1158) );
INV_X1 U835 ( .A(G478), .ZN(n1160) );
NOR2_X1 U836 ( .A1(n1144), .A2(n1161), .ZN(G60) );
XNOR2_X1 U837 ( .A(n1162), .B(n1163), .ZN(n1161) );
NOR2_X1 U838 ( .A1(n1164), .A2(n1159), .ZN(n1163) );
XOR2_X1 U839 ( .A(n1165), .B(n1166), .Z(G6) );
NAND2_X1 U840 ( .A1(KEYINPUT52), .A2(G104), .ZN(n1166) );
NOR2_X1 U841 ( .A1(n1144), .A2(n1167), .ZN(G57) );
XOR2_X1 U842 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U844 ( .A1(KEYINPUT55), .A2(n1172), .ZN(n1170) );
XOR2_X1 U845 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U846 ( .A(n1175), .B(n1176), .Z(n1173) );
NOR2_X1 U847 ( .A1(n1177), .A2(n1159), .ZN(n1176) );
NAND2_X1 U848 ( .A1(KEYINPUT49), .A2(n1178), .ZN(n1175) );
NAND2_X1 U849 ( .A1(KEYINPUT59), .A2(n1179), .ZN(n1168) );
NOR2_X1 U850 ( .A1(n1144), .A2(n1180), .ZN(G54) );
XOR2_X1 U851 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U852 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR3_X1 U853 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
NOR2_X1 U854 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
INV_X1 U855 ( .A(n1190), .ZN(n1189) );
NOR2_X1 U856 ( .A1(KEYINPUT51), .A2(n1191), .ZN(n1188) );
XNOR2_X1 U857 ( .A(KEYINPUT9), .B(n1192), .ZN(n1191) );
NOR3_X1 U858 ( .A1(n1190), .A2(KEYINPUT51), .A3(n1193), .ZN(n1186) );
XOR2_X1 U859 ( .A(n1194), .B(n1195), .Z(n1190) );
AND2_X1 U860 ( .A1(n1193), .A2(KEYINPUT51), .ZN(n1185) );
NOR2_X1 U861 ( .A1(n1196), .A2(n1159), .ZN(n1183) );
XOR2_X1 U862 ( .A(n1197), .B(n1198), .Z(n1181) );
NAND2_X1 U863 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND2_X1 U864 ( .A1(G140), .A2(n1201), .ZN(n1200) );
XOR2_X1 U865 ( .A(KEYINPUT20), .B(n1202), .Z(n1199) );
NOR2_X1 U866 ( .A1(G140), .A2(n1201), .ZN(n1202) );
XOR2_X1 U867 ( .A(KEYINPUT41), .B(G110), .Z(n1201) );
NOR3_X1 U868 ( .A1(n1203), .A2(n1144), .A3(n1204), .ZN(G51) );
NOR4_X1 U869 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1159), .ZN(n1204) );
NOR2_X1 U870 ( .A1(KEYINPUT25), .A2(n1208), .ZN(n1206) );
NOR2_X1 U871 ( .A1(n1209), .A2(n1210), .ZN(n1205) );
NOR2_X1 U872 ( .A1(KEYINPUT50), .A2(KEYINPUT25), .ZN(n1209) );
NOR2_X1 U873 ( .A1(n1085), .A2(G952), .ZN(n1144) );
NOR2_X1 U874 ( .A1(n1211), .A2(n1212), .ZN(n1203) );
NOR2_X1 U875 ( .A1(KEYINPUT50), .A2(n1210), .ZN(n1212) );
INV_X1 U876 ( .A(n1208), .ZN(n1210) );
XNOR2_X1 U877 ( .A(n1213), .B(n1214), .ZN(n1208) );
XOR2_X1 U878 ( .A(n1215), .B(n1216), .Z(n1213) );
NAND2_X1 U879 ( .A1(KEYINPUT12), .A2(n1217), .ZN(n1215) );
NOR2_X1 U880 ( .A1(n1207), .A2(n1159), .ZN(n1211) );
NAND2_X1 U881 ( .A1(G902), .A2(n1153), .ZN(n1159) );
NAND2_X1 U882 ( .A1(n1218), .A2(n1083), .ZN(n1153) );
AND4_X1 U883 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1083) );
AND4_X1 U884 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1222) );
NAND3_X1 U885 ( .A1(n1073), .A2(n1227), .A3(n1228), .ZN(n1221) );
NAND2_X1 U886 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
NAND2_X1 U887 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XNOR2_X1 U888 ( .A(n1233), .B(KEYINPUT11), .ZN(n1231) );
NAND2_X1 U889 ( .A1(n1234), .A2(n1079), .ZN(n1229) );
INV_X1 U890 ( .A(n1050), .ZN(n1218) );
NAND3_X1 U891 ( .A1(n1142), .A2(n1044), .A3(n1235), .ZN(n1050) );
XOR2_X1 U892 ( .A(n1141), .B(KEYINPUT34), .Z(n1235) );
NAND3_X1 U893 ( .A1(n1236), .A2(n1070), .A3(n1237), .ZN(n1044) );
NOR4_X1 U894 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1142) );
NAND3_X1 U895 ( .A1(n1242), .A2(n1243), .A3(n1165), .ZN(n1241) );
NAND3_X1 U896 ( .A1(n1236), .A2(n1237), .A3(n1073), .ZN(n1165) );
INV_X1 U897 ( .A(n1063), .ZN(n1236) );
OR3_X1 U898 ( .A1(n1244), .A2(n1245), .A3(n1082), .ZN(n1242) );
XOR2_X1 U899 ( .A(G146), .B(n1246), .Z(G48) );
NOR2_X1 U900 ( .A1(KEYINPUT60), .A2(n1219), .ZN(n1246) );
NAND4_X1 U901 ( .A1(n1234), .A2(n1073), .A3(n1247), .A4(n1065), .ZN(n1219) );
XOR2_X1 U902 ( .A(n1220), .B(n1248), .Z(G45) );
NAND2_X1 U903 ( .A1(KEYINPUT31), .A2(n1249), .ZN(n1248) );
XOR2_X1 U904 ( .A(KEYINPUT53), .B(G143), .Z(n1249) );
NAND3_X1 U905 ( .A1(n1250), .A2(n1251), .A3(n1232), .ZN(n1220) );
XNOR2_X1 U906 ( .A(G140), .B(n1252), .ZN(G42) );
NAND3_X1 U907 ( .A1(n1234), .A2(n1228), .A3(n1253), .ZN(n1252) );
NOR3_X1 U908 ( .A1(n1244), .A2(KEYINPUT26), .A3(n1065), .ZN(n1253) );
XOR2_X1 U909 ( .A(n1226), .B(n1254), .Z(G39) );
XNOR2_X1 U910 ( .A(KEYINPUT62), .B(n1127), .ZN(n1254) );
NAND4_X1 U911 ( .A1(n1234), .A2(n1228), .A3(n1255), .A4(n1065), .ZN(n1226) );
XNOR2_X1 U912 ( .A(G134), .B(n1225), .ZN(G36) );
NAND4_X1 U913 ( .A1(n1228), .A2(n1232), .A3(n1070), .A4(n1251), .ZN(n1225) );
XNOR2_X1 U914 ( .A(G131), .B(n1256), .ZN(G33) );
NAND3_X1 U915 ( .A1(n1228), .A2(n1232), .A3(n1257), .ZN(n1256) );
NOR3_X1 U916 ( .A1(n1244), .A2(KEYINPUT5), .A3(n1233), .ZN(n1257) );
INV_X1 U917 ( .A(n1073), .ZN(n1244) );
INV_X1 U918 ( .A(n1052), .ZN(n1228) );
NAND2_X1 U919 ( .A1(n1091), .A2(n1258), .ZN(n1052) );
NAND2_X1 U920 ( .A1(n1259), .A2(n1260), .ZN(G30) );
NAND2_X1 U921 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
INV_X1 U922 ( .A(G128), .ZN(n1262) );
NAND2_X1 U923 ( .A1(G128), .A2(n1263), .ZN(n1259) );
NAND2_X1 U924 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NAND2_X1 U925 ( .A1(KEYINPUT3), .A2(n1266), .ZN(n1265) );
INV_X1 U926 ( .A(n1223), .ZN(n1266) );
OR2_X1 U927 ( .A1(n1261), .A2(KEYINPUT3), .ZN(n1264) );
NOR2_X1 U928 ( .A1(KEYINPUT29), .A2(n1223), .ZN(n1261) );
NAND4_X1 U929 ( .A1(n1234), .A2(n1070), .A3(n1247), .A4(n1065), .ZN(n1223) );
INV_X1 U930 ( .A(n1074), .ZN(n1070) );
NOR3_X1 U931 ( .A1(n1080), .A2(n1233), .A3(n1075), .ZN(n1234) );
NAND2_X1 U932 ( .A1(n1267), .A2(n1268), .ZN(G3) );
NAND2_X1 U933 ( .A1(n1269), .A2(n1179), .ZN(n1268) );
XOR2_X1 U934 ( .A(n1270), .B(KEYINPUT42), .Z(n1267) );
OR2_X1 U935 ( .A1(n1269), .A2(n1179), .ZN(n1270) );
NAND2_X1 U936 ( .A1(n1271), .A2(n1272), .ZN(n1269) );
OR2_X1 U937 ( .A1(n1141), .A2(KEYINPUT57), .ZN(n1272) );
OR2_X1 U938 ( .A1(n1273), .A2(n1089), .ZN(n1141) );
NAND3_X1 U939 ( .A1(n1247), .A2(n1273), .A3(KEYINPUT57), .ZN(n1271) );
NAND3_X1 U940 ( .A1(n1255), .A2(n1274), .A3(n1232), .ZN(n1273) );
NOR3_X1 U941 ( .A1(n1075), .A2(n1079), .A3(n1082), .ZN(n1232) );
XNOR2_X1 U942 ( .A(G125), .B(n1224), .ZN(G27) );
NAND4_X1 U943 ( .A1(n1087), .A2(n1247), .A3(n1073), .A4(n1275), .ZN(n1224) );
NOR3_X1 U944 ( .A1(n1065), .A2(n1233), .A3(n1080), .ZN(n1275) );
INV_X1 U945 ( .A(n1251), .ZN(n1233) );
NAND2_X1 U946 ( .A1(n1060), .A2(n1276), .ZN(n1251) );
NAND4_X1 U947 ( .A1(n1277), .A2(G953), .A3(G902), .A4(n1111), .ZN(n1276) );
INV_X1 U948 ( .A(G900), .ZN(n1111) );
XOR2_X1 U949 ( .A(n1278), .B(KEYINPUT44), .Z(n1277) );
XNOR2_X1 U950 ( .A(G122), .B(n1243), .ZN(G24) );
NAND3_X1 U951 ( .A1(n1250), .A2(n1087), .A3(n1279), .ZN(n1243) );
NOR3_X1 U952 ( .A1(n1063), .A2(n1280), .A3(n1065), .ZN(n1279) );
XOR2_X1 U953 ( .A(n1082), .B(KEYINPUT45), .Z(n1063) );
NOR3_X1 U954 ( .A1(n1099), .A2(n1281), .A3(n1089), .ZN(n1250) );
XOR2_X1 U955 ( .A(G119), .B(n1240), .Z(G21) );
NOR3_X1 U956 ( .A1(n1076), .A2(n1080), .A3(n1245), .ZN(n1240) );
INV_X1 U957 ( .A(n1082), .ZN(n1080) );
XNOR2_X1 U958 ( .A(n1282), .B(n1238), .ZN(G18) );
NOR3_X1 U959 ( .A1(n1082), .A2(n1074), .A3(n1245), .ZN(n1238) );
NAND4_X1 U960 ( .A1(n1087), .A2(n1247), .A3(n1065), .A4(n1274), .ZN(n1245) );
NAND2_X1 U961 ( .A1(n1099), .A2(n1283), .ZN(n1074) );
XNOR2_X1 U962 ( .A(G113), .B(n1284), .ZN(G15) );
NAND4_X1 U963 ( .A1(n1073), .A2(n1087), .A3(n1285), .A4(n1286), .ZN(n1284) );
NOR3_X1 U964 ( .A1(n1082), .A2(n1280), .A3(n1079), .ZN(n1286) );
INV_X1 U965 ( .A(n1065), .ZN(n1079) );
XNOR2_X1 U966 ( .A(n1247), .B(KEYINPUT1), .ZN(n1285) );
INV_X1 U967 ( .A(n1069), .ZN(n1087) );
NAND2_X1 U968 ( .A1(n1058), .A2(n1287), .ZN(n1069) );
NOR2_X1 U969 ( .A1(n1283), .A2(n1099), .ZN(n1073) );
XOR2_X1 U970 ( .A(G110), .B(n1239), .Z(G12) );
AND3_X1 U971 ( .A1(n1237), .A2(n1082), .A3(n1255), .ZN(n1239) );
INV_X1 U972 ( .A(n1076), .ZN(n1255) );
NAND2_X1 U973 ( .A1(n1281), .A2(n1099), .ZN(n1076) );
XNOR2_X1 U974 ( .A(n1288), .B(n1164), .ZN(n1099) );
INV_X1 U975 ( .A(G475), .ZN(n1164) );
NAND2_X1 U976 ( .A1(n1289), .A2(n1162), .ZN(n1288) );
NAND2_X1 U977 ( .A1(n1290), .A2(n1291), .ZN(n1162) );
NAND2_X1 U978 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XOR2_X1 U979 ( .A(n1294), .B(KEYINPUT16), .Z(n1290) );
OR2_X1 U980 ( .A1(n1293), .A2(n1292), .ZN(n1294) );
XNOR2_X1 U981 ( .A(n1295), .B(n1296), .ZN(n1292) );
XOR2_X1 U982 ( .A(n1114), .B(n1297), .Z(n1296) );
XOR2_X1 U983 ( .A(n1298), .B(n1299), .Z(n1295) );
AND3_X1 U984 ( .A1(G214), .A2(n1085), .A3(n1300), .ZN(n1299) );
NAND2_X1 U985 ( .A1(KEYINPUT15), .A2(n1125), .ZN(n1298) );
XNOR2_X1 U986 ( .A(n1301), .B(n1302), .ZN(n1293) );
NOR2_X1 U987 ( .A1(KEYINPUT37), .A2(n1303), .ZN(n1302) );
XNOR2_X1 U988 ( .A(G113), .B(G122), .ZN(n1303) );
XNOR2_X1 U989 ( .A(G104), .B(KEYINPUT38), .ZN(n1301) );
INV_X1 U990 ( .A(n1283), .ZN(n1281) );
NAND3_X1 U991 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n1283) );
INV_X1 U992 ( .A(n1101), .ZN(n1306) );
NOR2_X1 U993 ( .A1(n1103), .A2(G478), .ZN(n1101) );
OR2_X1 U994 ( .A1(G478), .A2(KEYINPUT40), .ZN(n1305) );
NAND3_X1 U995 ( .A1(G478), .A2(n1103), .A3(KEYINPUT40), .ZN(n1304) );
NAND2_X1 U996 ( .A1(n1157), .A2(n1289), .ZN(n1103) );
XNOR2_X1 U997 ( .A(n1307), .B(n1308), .ZN(n1157) );
XOR2_X1 U998 ( .A(n1309), .B(n1310), .Z(n1308) );
NOR2_X1 U999 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NOR2_X1 U1000 ( .A1(KEYINPUT47), .A2(n1313), .ZN(n1312) );
INV_X1 U1001 ( .A(n1314), .ZN(n1313) );
NOR2_X1 U1002 ( .A1(KEYINPUT0), .A2(n1314), .ZN(n1311) );
NAND3_X1 U1003 ( .A1(G234), .A2(n1085), .A3(G217), .ZN(n1314) );
NOR2_X1 U1004 ( .A1(n1315), .A2(n1316), .ZN(n1309) );
XOR2_X1 U1005 ( .A(n1317), .B(KEYINPUT8), .Z(n1316) );
NAND2_X1 U1006 ( .A1(G122), .A2(n1282), .ZN(n1317) );
NOR2_X1 U1007 ( .A1(G122), .A2(n1282), .ZN(n1315) );
INV_X1 U1008 ( .A(G116), .ZN(n1282) );
XOR2_X1 U1009 ( .A(n1318), .B(G107), .Z(n1307) );
NAND2_X1 U1010 ( .A1(n1319), .A2(KEYINPUT46), .ZN(n1318) );
XNOR2_X1 U1011 ( .A(n1320), .B(n1321), .ZN(n1319) );
XNOR2_X1 U1012 ( .A(G143), .B(G134), .ZN(n1320) );
XNOR2_X1 U1013 ( .A(n1322), .B(n1152), .ZN(n1082) );
AND2_X1 U1014 ( .A1(G217), .A2(n1323), .ZN(n1152) );
NAND2_X1 U1015 ( .A1(n1155), .A2(n1289), .ZN(n1322) );
XOR2_X1 U1016 ( .A(n1324), .B(n1325), .Z(n1155) );
XOR2_X1 U1017 ( .A(n1326), .B(n1327), .Z(n1325) );
XNOR2_X1 U1018 ( .A(n1328), .B(n1329), .ZN(n1327) );
NOR2_X1 U1019 ( .A1(KEYINPUT63), .A2(G110), .ZN(n1329) );
NAND2_X1 U1020 ( .A1(KEYINPUT35), .A2(G119), .ZN(n1328) );
XNOR2_X1 U1021 ( .A(G146), .B(n1127), .ZN(n1326) );
XNOR2_X1 U1022 ( .A(n1330), .B(n1331), .ZN(n1324) );
XOR2_X1 U1023 ( .A(n1332), .B(n1114), .Z(n1331) );
XOR2_X1 U1024 ( .A(G125), .B(G140), .Z(n1114) );
AND3_X1 U1025 ( .A1(G221), .A2(n1085), .A3(G234), .ZN(n1332) );
NOR4_X1 U1026 ( .A1(n1089), .A2(n1075), .A3(n1065), .A4(n1280), .ZN(n1237) );
INV_X1 U1027 ( .A(n1274), .ZN(n1280) );
NAND2_X1 U1028 ( .A1(n1060), .A2(n1333), .ZN(n1274) );
NAND4_X1 U1029 ( .A1(G953), .A2(G902), .A3(n1278), .A4(n1334), .ZN(n1333) );
INV_X1 U1030 ( .A(G898), .ZN(n1334) );
NAND3_X1 U1031 ( .A1(n1278), .A2(n1085), .A3(G952), .ZN(n1060) );
NAND2_X1 U1032 ( .A1(G237), .A2(G234), .ZN(n1278) );
XOR2_X1 U1033 ( .A(n1335), .B(n1177), .Z(n1065) );
INV_X1 U1034 ( .A(G472), .ZN(n1177) );
NAND2_X1 U1035 ( .A1(n1336), .A2(n1289), .ZN(n1335) );
XOR2_X1 U1036 ( .A(n1337), .B(n1338), .Z(n1336) );
XNOR2_X1 U1037 ( .A(n1174), .B(n1178), .ZN(n1338) );
XOR2_X1 U1038 ( .A(n1192), .B(n1339), .Z(n1178) );
XNOR2_X1 U1039 ( .A(n1340), .B(G113), .ZN(n1174) );
NAND2_X1 U1040 ( .A1(KEYINPUT43), .A2(n1341), .ZN(n1340) );
XNOR2_X1 U1041 ( .A(n1179), .B(n1171), .ZN(n1337) );
AND3_X1 U1042 ( .A1(n1300), .A2(n1085), .A3(G210), .ZN(n1171) );
OR2_X1 U1043 ( .A1(n1058), .A2(n1056), .ZN(n1075) );
INV_X1 U1044 ( .A(n1287), .ZN(n1056) );
NAND2_X1 U1045 ( .A1(G221), .A2(n1323), .ZN(n1287) );
NAND2_X1 U1046 ( .A1(G234), .A2(n1342), .ZN(n1323) );
XNOR2_X1 U1047 ( .A(n1343), .B(n1196), .ZN(n1058) );
INV_X1 U1048 ( .A(G469), .ZN(n1196) );
NAND2_X1 U1049 ( .A1(n1289), .A2(n1344), .ZN(n1343) );
XOR2_X1 U1050 ( .A(n1345), .B(n1346), .Z(n1344) );
XOR2_X1 U1051 ( .A(n1195), .B(n1347), .Z(n1346) );
XNOR2_X1 U1052 ( .A(n1197), .B(n1348), .ZN(n1347) );
NAND2_X1 U1053 ( .A1(G227), .A2(n1085), .ZN(n1197) );
XOR2_X1 U1054 ( .A(n1115), .B(n1349), .Z(n1195) );
NOR2_X1 U1055 ( .A1(KEYINPUT32), .A2(n1179), .ZN(n1349) );
INV_X1 U1056 ( .A(G101), .ZN(n1179) );
XNOR2_X1 U1057 ( .A(n1297), .B(n1321), .ZN(n1115) );
XNOR2_X1 U1058 ( .A(n1193), .B(n1350), .ZN(n1345) );
XNOR2_X1 U1059 ( .A(G140), .B(KEYINPUT28), .ZN(n1350) );
INV_X1 U1060 ( .A(n1192), .ZN(n1193) );
NAND3_X1 U1061 ( .A1(n1122), .A2(n1121), .A3(n1119), .ZN(n1192) );
NAND3_X1 U1062 ( .A1(G134), .A2(n1127), .A3(G131), .ZN(n1119) );
NAND3_X1 U1063 ( .A1(n1351), .A2(n1127), .A3(n1125), .ZN(n1121) );
INV_X1 U1064 ( .A(G131), .ZN(n1125) );
INV_X1 U1065 ( .A(G137), .ZN(n1127) );
NAND2_X1 U1066 ( .A1(G137), .A2(n1352), .ZN(n1122) );
XNOR2_X1 U1067 ( .A(n1351), .B(G131), .ZN(n1352) );
INV_X1 U1068 ( .A(G134), .ZN(n1351) );
INV_X1 U1069 ( .A(n1247), .ZN(n1089) );
NOR2_X1 U1070 ( .A1(n1091), .A2(n1092), .ZN(n1247) );
INV_X1 U1071 ( .A(n1258), .ZN(n1092) );
NAND2_X1 U1072 ( .A1(G214), .A2(n1353), .ZN(n1258) );
XNOR2_X1 U1073 ( .A(n1354), .B(n1207), .ZN(n1091) );
NAND2_X1 U1074 ( .A1(G210), .A2(n1353), .ZN(n1207) );
NAND2_X1 U1075 ( .A1(n1300), .A2(n1342), .ZN(n1353) );
INV_X1 U1076 ( .A(G902), .ZN(n1342) );
INV_X1 U1077 ( .A(G237), .ZN(n1300) );
NAND2_X1 U1078 ( .A1(n1355), .A2(n1289), .ZN(n1354) );
XNOR2_X1 U1079 ( .A(G902), .B(KEYINPUT10), .ZN(n1289) );
XNOR2_X1 U1080 ( .A(n1217), .B(n1356), .ZN(n1355) );
XOR2_X1 U1081 ( .A(n1357), .B(n1216), .Z(n1356) );
AND2_X1 U1082 ( .A1(G224), .A2(n1085), .ZN(n1216) );
INV_X1 U1083 ( .A(G953), .ZN(n1085) );
NAND2_X1 U1084 ( .A1(KEYINPUT61), .A2(n1214), .ZN(n1357) );
XOR2_X1 U1085 ( .A(n1135), .B(n1137), .Z(n1214) );
XNOR2_X1 U1086 ( .A(n1358), .B(n1341), .ZN(n1137) );
XOR2_X1 U1087 ( .A(G119), .B(G116), .Z(n1341) );
INV_X1 U1088 ( .A(G113), .ZN(n1358) );
XNOR2_X1 U1089 ( .A(n1359), .B(n1360), .ZN(n1135) );
XOR2_X1 U1090 ( .A(KEYINPUT33), .B(G122), .Z(n1360) );
XNOR2_X1 U1091 ( .A(n1348), .B(G101), .ZN(n1359) );
XNOR2_X1 U1092 ( .A(G110), .B(n1361), .ZN(n1348) );
INV_X1 U1093 ( .A(n1194), .ZN(n1361) );
XOR2_X1 U1094 ( .A(G104), .B(G107), .Z(n1194) );
XOR2_X1 U1095 ( .A(G125), .B(n1339), .Z(n1217) );
XNOR2_X1 U1096 ( .A(n1362), .B(n1297), .ZN(n1339) );
XOR2_X1 U1097 ( .A(G143), .B(G146), .Z(n1297) );
NAND2_X1 U1098 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
NAND2_X1 U1099 ( .A1(KEYINPUT6), .A2(n1321), .ZN(n1364) );
INV_X1 U1100 ( .A(n1330), .ZN(n1321) );
NAND2_X1 U1101 ( .A1(KEYINPUT39), .A2(n1330), .ZN(n1363) );
XOR2_X1 U1102 ( .A(G128), .B(KEYINPUT13), .Z(n1330) );
endmodule


