//Key = 1001000101011100001100101110010111110011001110010110101101100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412;

XNOR2_X1 U765 ( .A(n1070), .B(n1071), .ZN(G9) );
NOR2_X1 U766 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U767 ( .A(n1074), .B(KEYINPUT45), .Z(n1072) );
NOR2_X1 U768 ( .A1(n1075), .A2(n1076), .ZN(G75) );
NOR3_X1 U769 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1076) );
NAND3_X1 U770 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1077) );
NAND2_X1 U771 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U772 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND3_X1 U773 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NAND2_X1 U774 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NAND2_X1 U775 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
OR2_X1 U776 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U777 ( .A1(n1096), .A2(n1097), .ZN(n1090) );
NAND2_X1 U778 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND3_X1 U779 ( .A1(G221), .A2(n1100), .A3(n1101), .ZN(n1099) );
NAND3_X1 U780 ( .A1(n1092), .A2(n1102), .A3(n1096), .ZN(n1085) );
NAND2_X1 U781 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND3_X1 U782 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1104) );
NAND2_X1 U783 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NAND3_X1 U784 ( .A1(n1110), .A2(n1073), .A3(n1111), .ZN(n1105) );
NAND2_X1 U785 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NAND2_X1 U786 ( .A1(n1089), .A2(n1114), .ZN(n1103) );
INV_X1 U787 ( .A(n1115), .ZN(n1083) );
NOR3_X1 U788 ( .A1(n1116), .A2(G953), .A3(G952), .ZN(n1075) );
INV_X1 U789 ( .A(n1080), .ZN(n1116) );
NAND4_X1 U790 ( .A1(n1117), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1080) );
NOR4_X1 U791 ( .A1(n1108), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1120) );
XNOR2_X1 U792 ( .A(G472), .B(n1124), .ZN(n1123) );
NAND2_X1 U793 ( .A1(KEYINPUT35), .A2(n1125), .ZN(n1124) );
NOR3_X1 U794 ( .A1(n1126), .A2(n1127), .A3(n1112), .ZN(n1119) );
NOR2_X1 U795 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NOR2_X1 U796 ( .A1(G902), .A2(n1130), .ZN(n1128) );
NAND2_X1 U797 ( .A1(n1131), .A2(n1132), .ZN(n1118) );
XOR2_X1 U798 ( .A(KEYINPUT22), .B(n1133), .Z(n1117) );
XOR2_X1 U799 ( .A(n1134), .B(n1135), .Z(G72) );
NOR2_X1 U800 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XOR2_X1 U801 ( .A(n1138), .B(KEYINPUT29), .Z(n1137) );
NAND3_X1 U802 ( .A1(n1078), .A2(n1081), .A3(n1139), .ZN(n1138) );
NOR3_X1 U803 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1136) );
NOR2_X1 U804 ( .A1(G953), .A2(n1142), .ZN(n1141) );
NOR2_X1 U805 ( .A1(G900), .A2(n1081), .ZN(n1140) );
XOR2_X1 U806 ( .A(n1143), .B(n1144), .Z(n1139) );
XNOR2_X1 U807 ( .A(G140), .B(n1145), .ZN(n1144) );
NAND2_X1 U808 ( .A1(n1146), .A2(KEYINPUT54), .ZN(n1145) );
XOR2_X1 U809 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U810 ( .A1(KEYINPUT21), .A2(n1149), .ZN(n1148) );
XNOR2_X1 U811 ( .A(n1150), .B(n1151), .ZN(n1147) );
NAND3_X1 U812 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1150) );
NAND2_X1 U813 ( .A1(G137), .A2(n1155), .ZN(n1154) );
NAND2_X1 U814 ( .A1(KEYINPUT56), .A2(n1156), .ZN(n1153) );
NAND2_X1 U815 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XNOR2_X1 U816 ( .A(KEYINPUT27), .B(n1155), .ZN(n1157) );
NAND2_X1 U817 ( .A1(n1159), .A2(n1160), .ZN(n1152) );
INV_X1 U818 ( .A(KEYINPUT56), .ZN(n1160) );
NAND2_X1 U819 ( .A1(n1161), .A2(n1162), .ZN(n1159) );
OR3_X1 U820 ( .A1(n1155), .A2(G137), .A3(KEYINPUT27), .ZN(n1162) );
NAND2_X1 U821 ( .A1(KEYINPUT27), .A2(n1155), .ZN(n1161) );
INV_X1 U822 ( .A(G134), .ZN(n1155) );
NAND2_X1 U823 ( .A1(KEYINPUT33), .A2(n1163), .ZN(n1143) );
NAND2_X1 U824 ( .A1(G953), .A2(n1164), .ZN(n1134) );
NAND2_X1 U825 ( .A1(G900), .A2(G227), .ZN(n1164) );
NAND3_X1 U826 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(G69) );
NAND2_X1 U827 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U828 ( .A1(KEYINPUT55), .A2(n1170), .ZN(n1169) );
XOR2_X1 U829 ( .A(KEYINPUT1), .B(n1171), .Z(n1170) );
NAND3_X1 U830 ( .A1(KEYINPUT55), .A2(n1172), .A3(n1171), .ZN(n1166) );
INV_X1 U831 ( .A(n1168), .ZN(n1172) );
XNOR2_X1 U832 ( .A(n1173), .B(n1174), .ZN(n1168) );
NOR2_X1 U833 ( .A1(n1175), .A2(G953), .ZN(n1174) );
NAND2_X1 U834 ( .A1(n1176), .A2(n1177), .ZN(n1173) );
NAND2_X1 U835 ( .A1(G953), .A2(n1178), .ZN(n1177) );
XOR2_X1 U836 ( .A(KEYINPUT47), .B(G898), .Z(n1178) );
XOR2_X1 U837 ( .A(n1179), .B(n1180), .Z(n1176) );
NOR2_X1 U838 ( .A1(KEYINPUT30), .A2(n1181), .ZN(n1180) );
OR2_X1 U839 ( .A1(n1171), .A2(KEYINPUT55), .ZN(n1165) );
AND2_X1 U840 ( .A1(G953), .A2(n1182), .ZN(n1171) );
NAND2_X1 U841 ( .A1(G898), .A2(G224), .ZN(n1182) );
NOR3_X1 U842 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(G66) );
NOR2_X1 U843 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
XOR2_X1 U844 ( .A(n1188), .B(KEYINPUT15), .Z(n1187) );
AND2_X1 U845 ( .A1(n1188), .A2(n1186), .ZN(n1184) );
NOR2_X1 U846 ( .A1(n1189), .A2(n1190), .ZN(n1186) );
NOR2_X1 U847 ( .A1(n1191), .A2(n1192), .ZN(G63) );
XNOR2_X1 U848 ( .A(n1183), .B(KEYINPUT19), .ZN(n1192) );
XNOR2_X1 U849 ( .A(n1193), .B(n1194), .ZN(n1191) );
NOR2_X1 U850 ( .A1(n1195), .A2(n1189), .ZN(n1194) );
INV_X1 U851 ( .A(G478), .ZN(n1195) );
NOR2_X1 U852 ( .A1(n1183), .A2(n1196), .ZN(G60) );
XNOR2_X1 U853 ( .A(n1197), .B(n1198), .ZN(n1196) );
NOR2_X1 U854 ( .A1(n1199), .A2(n1189), .ZN(n1198) );
XNOR2_X1 U855 ( .A(n1200), .B(n1201), .ZN(G6) );
XOR2_X1 U856 ( .A(KEYINPUT44), .B(G104), .Z(n1201) );
NOR2_X1 U857 ( .A1(n1183), .A2(n1202), .ZN(G57) );
XOR2_X1 U858 ( .A(n1203), .B(n1204), .Z(n1202) );
XNOR2_X1 U859 ( .A(G101), .B(n1205), .ZN(n1204) );
NAND2_X1 U860 ( .A1(n1206), .A2(n1207), .ZN(n1203) );
NAND2_X1 U861 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XNOR2_X1 U862 ( .A(KEYINPUT6), .B(n1210), .ZN(n1208) );
NAND2_X1 U863 ( .A1(n1211), .A2(n1212), .ZN(n1206) );
XOR2_X1 U864 ( .A(n1209), .B(n1213), .Z(n1212) );
XOR2_X1 U865 ( .A(KEYINPUT59), .B(KEYINPUT43), .Z(n1213) );
XNOR2_X1 U866 ( .A(n1214), .B(n1215), .ZN(n1209) );
XNOR2_X1 U867 ( .A(n1216), .B(n1217), .ZN(n1214) );
NOR2_X1 U868 ( .A1(n1218), .A2(n1189), .ZN(n1217) );
INV_X1 U869 ( .A(G472), .ZN(n1218) );
XOR2_X1 U870 ( .A(KEYINPUT6), .B(n1210), .Z(n1211) );
NOR2_X1 U871 ( .A1(n1183), .A2(n1219), .ZN(G54) );
XOR2_X1 U872 ( .A(n1220), .B(n1221), .Z(n1219) );
XNOR2_X1 U873 ( .A(n1222), .B(n1223), .ZN(n1221) );
XOR2_X1 U874 ( .A(KEYINPUT42), .B(n1224), .Z(n1223) );
NOR2_X1 U875 ( .A1(n1225), .A2(n1189), .ZN(n1224) );
XOR2_X1 U876 ( .A(n1226), .B(n1227), .Z(n1220) );
NOR2_X1 U877 ( .A1(n1183), .A2(n1228), .ZN(G51) );
XOR2_X1 U878 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U879 ( .A(n1231), .B(n1232), .Z(n1230) );
NAND2_X1 U880 ( .A1(n1233), .A2(KEYINPUT31), .ZN(n1231) );
XOR2_X1 U881 ( .A(n1234), .B(n1235), .Z(n1229) );
NOR2_X1 U882 ( .A1(n1132), .A2(n1189), .ZN(n1235) );
NAND2_X1 U883 ( .A1(G902), .A2(n1236), .ZN(n1189) );
NAND2_X1 U884 ( .A1(n1175), .A2(n1142), .ZN(n1236) );
INV_X1 U885 ( .A(n1078), .ZN(n1142) );
NAND4_X1 U886 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1078) );
NOR4_X1 U887 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1240) );
NOR2_X1 U888 ( .A1(KEYINPUT41), .A2(n1245), .ZN(n1244) );
NOR2_X1 U889 ( .A1(KEYINPUT37), .A2(n1246), .ZN(n1243) );
NOR3_X1 U890 ( .A1(n1109), .A2(n1247), .A3(n1248), .ZN(n1242) );
NOR2_X1 U891 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
AND4_X1 U892 ( .A1(n1251), .A2(n1095), .A3(n1114), .A4(KEYINPUT41), .ZN(n1250) );
NOR2_X1 U893 ( .A1(n1252), .A2(n1098), .ZN(n1247) );
INV_X1 U894 ( .A(n1249), .ZN(n1098) );
NOR3_X1 U895 ( .A1(n1253), .A2(n1251), .A3(n1254), .ZN(n1252) );
INV_X1 U896 ( .A(KEYINPUT37), .ZN(n1254) );
NAND3_X1 U897 ( .A1(n1107), .A2(n1108), .A3(n1094), .ZN(n1253) );
NOR3_X1 U898 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1239) );
INV_X1 U899 ( .A(n1079), .ZN(n1175) );
NAND2_X1 U900 ( .A1(n1258), .A2(n1259), .ZN(n1079) );
NOR4_X1 U901 ( .A1(n1260), .A2(n1200), .A3(n1261), .A4(n1262), .ZN(n1259) );
AND4_X1 U902 ( .A1(n1087), .A2(n1263), .A3(n1249), .A4(n1264), .ZN(n1200) );
NOR2_X1 U903 ( .A1(n1073), .A2(n1265), .ZN(n1264) );
INV_X1 U904 ( .A(n1266), .ZN(n1260) );
NOR4_X1 U905 ( .A1(n1267), .A2(n1268), .A3(n1269), .A4(n1270), .ZN(n1258) );
NOR2_X1 U906 ( .A1(n1074), .A2(n1073), .ZN(n1270) );
INV_X1 U907 ( .A(n1271), .ZN(n1073) );
NAND4_X1 U908 ( .A1(n1249), .A2(n1095), .A3(n1087), .A4(n1263), .ZN(n1074) );
NOR2_X1 U909 ( .A1(n1081), .A2(G952), .ZN(n1183) );
NAND3_X1 U910 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(G48) );
NAND2_X1 U911 ( .A1(G146), .A2(n1275), .ZN(n1274) );
NAND2_X1 U912 ( .A1(n1276), .A2(n1277), .ZN(n1273) );
INV_X1 U913 ( .A(KEYINPUT26), .ZN(n1277) );
NAND2_X1 U914 ( .A1(n1278), .A2(n1241), .ZN(n1276) );
INV_X1 U915 ( .A(n1275), .ZN(n1241) );
XNOR2_X1 U916 ( .A(KEYINPUT2), .B(G146), .ZN(n1278) );
NAND2_X1 U917 ( .A1(KEYINPUT26), .A2(n1279), .ZN(n1272) );
NAND2_X1 U918 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
OR3_X1 U919 ( .A1(n1275), .A2(G146), .A3(KEYINPUT2), .ZN(n1281) );
NAND3_X1 U920 ( .A1(n1094), .A2(n1271), .A3(n1282), .ZN(n1275) );
NAND2_X1 U921 ( .A1(KEYINPUT2), .A2(G146), .ZN(n1280) );
XNOR2_X1 U922 ( .A(G143), .B(n1237), .ZN(G45) );
NAND4_X1 U923 ( .A1(n1283), .A2(n1271), .A3(n1121), .A4(n1284), .ZN(n1237) );
XNOR2_X1 U924 ( .A(G140), .B(n1246), .ZN(G42) );
NAND3_X1 U925 ( .A1(n1089), .A2(n1249), .A3(n1285), .ZN(n1246) );
XNOR2_X1 U926 ( .A(n1158), .B(n1257), .ZN(G39) );
AND3_X1 U927 ( .A1(n1282), .A2(n1096), .A3(n1089), .ZN(n1257) );
XNOR2_X1 U928 ( .A(G134), .B(n1245), .ZN(G36) );
NAND3_X1 U929 ( .A1(n1089), .A2(n1095), .A3(n1283), .ZN(n1245) );
XNOR2_X1 U930 ( .A(G131), .B(n1238), .ZN(G33) );
NAND3_X1 U931 ( .A1(n1089), .A2(n1094), .A3(n1283), .ZN(n1238) );
AND3_X1 U932 ( .A1(n1249), .A2(n1251), .A3(n1114), .ZN(n1283) );
INV_X1 U933 ( .A(n1109), .ZN(n1089) );
NAND2_X1 U934 ( .A1(n1113), .A2(n1286), .ZN(n1109) );
XOR2_X1 U935 ( .A(n1256), .B(n1287), .Z(G30) );
NOR2_X1 U936 ( .A1(KEYINPUT40), .A2(n1288), .ZN(n1287) );
AND3_X1 U937 ( .A1(n1271), .A2(n1095), .A3(n1282), .ZN(n1256) );
AND4_X1 U938 ( .A1(n1249), .A2(n1289), .A3(n1108), .A4(n1251), .ZN(n1282) );
XNOR2_X1 U939 ( .A(n1290), .B(n1269), .ZN(G3) );
AND2_X1 U940 ( .A1(n1114), .A2(n1291), .ZN(n1269) );
NAND3_X1 U941 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(G27) );
NAND2_X1 U942 ( .A1(G125), .A2(n1295), .ZN(n1294) );
NAND2_X1 U943 ( .A1(KEYINPUT8), .A2(n1296), .ZN(n1293) );
NAND2_X1 U944 ( .A1(n1297), .A2(n1255), .ZN(n1296) );
INV_X1 U945 ( .A(n1295), .ZN(n1255) );
XNOR2_X1 U946 ( .A(KEYINPUT10), .B(G125), .ZN(n1297) );
NAND2_X1 U947 ( .A1(n1298), .A2(n1299), .ZN(n1292) );
INV_X1 U948 ( .A(KEYINPUT8), .ZN(n1299) );
NAND2_X1 U949 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
OR3_X1 U950 ( .A1(n1295), .A2(G125), .A3(KEYINPUT10), .ZN(n1301) );
NAND3_X1 U951 ( .A1(n1092), .A2(n1271), .A3(n1285), .ZN(n1295) );
AND4_X1 U952 ( .A1(n1107), .A2(n1094), .A3(n1108), .A4(n1251), .ZN(n1285) );
NAND2_X1 U953 ( .A1(n1115), .A2(n1302), .ZN(n1251) );
NAND4_X1 U954 ( .A1(G953), .A2(G902), .A3(n1303), .A4(n1304), .ZN(n1302) );
INV_X1 U955 ( .A(G900), .ZN(n1304) );
XNOR2_X1 U956 ( .A(KEYINPUT57), .B(n1305), .ZN(n1303) );
NAND2_X1 U957 ( .A1(KEYINPUT10), .A2(G125), .ZN(n1300) );
XNOR2_X1 U958 ( .A(G122), .B(n1266), .ZN(G24) );
NAND4_X1 U959 ( .A1(n1306), .A2(n1087), .A3(n1121), .A4(n1284), .ZN(n1266) );
AND2_X1 U960 ( .A1(n1111), .A2(n1107), .ZN(n1087) );
XNOR2_X1 U961 ( .A(G119), .B(n1307), .ZN(G21) );
NAND2_X1 U962 ( .A1(KEYINPUT12), .A2(n1268), .ZN(n1307) );
AND4_X1 U963 ( .A1(n1096), .A2(n1306), .A3(n1289), .A4(n1108), .ZN(n1268) );
XNOR2_X1 U964 ( .A(n1267), .B(n1308), .ZN(G18) );
NAND2_X1 U965 ( .A1(KEYINPUT50), .A2(G116), .ZN(n1308) );
AND3_X1 U966 ( .A1(n1306), .A2(n1095), .A3(n1114), .ZN(n1267) );
NOR2_X1 U967 ( .A1(n1121), .A2(n1309), .ZN(n1095) );
XOR2_X1 U968 ( .A(G113), .B(n1262), .Z(G15) );
AND3_X1 U969 ( .A1(n1094), .A2(n1306), .A3(n1114), .ZN(n1262) );
AND2_X1 U970 ( .A1(n1111), .A2(n1289), .ZN(n1114) );
XNOR2_X1 U971 ( .A(n1310), .B(KEYINPUT28), .ZN(n1289) );
AND3_X1 U972 ( .A1(n1271), .A2(n1263), .A3(n1092), .ZN(n1306) );
INV_X1 U973 ( .A(n1122), .ZN(n1092) );
NAND2_X1 U974 ( .A1(n1101), .A2(n1311), .ZN(n1122) );
NAND2_X1 U975 ( .A1(G221), .A2(n1100), .ZN(n1311) );
INV_X1 U976 ( .A(n1265), .ZN(n1094) );
NAND2_X1 U977 ( .A1(n1309), .A2(n1121), .ZN(n1265) );
XOR2_X1 U978 ( .A(G110), .B(n1261), .Z(G12) );
AND3_X1 U979 ( .A1(n1107), .A2(n1108), .A3(n1291), .ZN(n1261) );
AND4_X1 U980 ( .A1(n1096), .A2(n1271), .A3(n1249), .A4(n1263), .ZN(n1291) );
NAND2_X1 U981 ( .A1(n1115), .A2(n1312), .ZN(n1263) );
NAND4_X1 U982 ( .A1(G953), .A2(G902), .A3(n1305), .A4(n1313), .ZN(n1312) );
INV_X1 U983 ( .A(G898), .ZN(n1313) );
NAND3_X1 U984 ( .A1(n1305), .A2(n1081), .A3(G952), .ZN(n1115) );
NAND2_X1 U985 ( .A1(G237), .A2(G234), .ZN(n1305) );
NOR2_X1 U986 ( .A1(n1101), .A2(n1314), .ZN(n1249) );
AND2_X1 U987 ( .A1(G221), .A2(n1100), .ZN(n1314) );
XNOR2_X1 U988 ( .A(n1315), .B(n1225), .ZN(n1101) );
INV_X1 U989 ( .A(G469), .ZN(n1225) );
NAND2_X1 U990 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XOR2_X1 U991 ( .A(n1226), .B(n1318), .Z(n1316) );
XNOR2_X1 U992 ( .A(n1319), .B(n1320), .ZN(n1318) );
NOR2_X1 U993 ( .A1(KEYINPUT14), .A2(n1222), .ZN(n1320) );
NAND2_X1 U994 ( .A1(KEYINPUT38), .A2(n1321), .ZN(n1319) );
XOR2_X1 U995 ( .A(KEYINPUT63), .B(n1227), .Z(n1321) );
XNOR2_X1 U996 ( .A(n1322), .B(n1323), .ZN(n1227) );
XOR2_X1 U997 ( .A(G140), .B(G110), .Z(n1323) );
NAND2_X1 U998 ( .A1(G227), .A2(n1081), .ZN(n1322) );
XNOR2_X1 U999 ( .A(n1149), .B(n1324), .ZN(n1226) );
XNOR2_X1 U1000 ( .A(n1290), .B(n1325), .ZN(n1324) );
NOR2_X1 U1001 ( .A1(KEYINPUT16), .A2(n1326), .ZN(n1325) );
XNOR2_X1 U1002 ( .A(G104), .B(G107), .ZN(n1326) );
INV_X1 U1003 ( .A(G101), .ZN(n1290) );
XOR2_X1 U1004 ( .A(n1327), .B(n1328), .Z(n1149) );
XNOR2_X1 U1005 ( .A(G128), .B(KEYINPUT3), .ZN(n1327) );
NOR2_X1 U1006 ( .A1(n1112), .A2(n1113), .ZN(n1271) );
NOR2_X1 U1007 ( .A1(n1329), .A2(n1127), .ZN(n1113) );
NOR2_X1 U1008 ( .A1(n1132), .A2(n1131), .ZN(n1127) );
XNOR2_X1 U1009 ( .A(KEYINPUT24), .B(n1330), .ZN(n1329) );
NOR2_X1 U1010 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U1011 ( .A(KEYINPUT58), .B(n1131), .Z(n1332) );
AND2_X1 U1012 ( .A1(n1333), .A2(n1317), .ZN(n1131) );
XOR2_X1 U1013 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1014 ( .A(n1232), .B(n1234), .Z(n1335) );
AND2_X1 U1015 ( .A1(G224), .A2(n1081), .ZN(n1234) );
XNOR2_X1 U1016 ( .A(n1179), .B(n1181), .ZN(n1232) );
XNOR2_X1 U1017 ( .A(G110), .B(n1336), .ZN(n1181) );
XNOR2_X1 U1018 ( .A(KEYINPUT5), .B(n1337), .ZN(n1336) );
XOR2_X1 U1019 ( .A(n1338), .B(n1339), .Z(n1179) );
XOR2_X1 U1020 ( .A(n1340), .B(n1341), .Z(n1339) );
XNOR2_X1 U1021 ( .A(G104), .B(G101), .ZN(n1341) );
NAND2_X1 U1022 ( .A1(KEYINPUT61), .A2(n1070), .ZN(n1340) );
INV_X1 U1023 ( .A(G107), .ZN(n1070) );
XOR2_X1 U1024 ( .A(n1342), .B(n1343), .Z(n1338) );
NAND2_X1 U1025 ( .A1(KEYINPUT11), .A2(G113), .ZN(n1342) );
NAND2_X1 U1026 ( .A1(n1344), .A2(n1345), .ZN(n1334) );
NAND2_X1 U1027 ( .A1(KEYINPUT7), .A2(n1233), .ZN(n1345) );
XNOR2_X1 U1028 ( .A(G125), .B(n1215), .ZN(n1233) );
OR3_X1 U1029 ( .A1(n1163), .A2(n1215), .A3(KEYINPUT7), .ZN(n1344) );
INV_X1 U1030 ( .A(n1132), .ZN(n1331) );
NAND2_X1 U1031 ( .A1(G210), .A2(n1346), .ZN(n1132) );
INV_X1 U1032 ( .A(n1286), .ZN(n1112) );
NAND2_X1 U1033 ( .A1(G214), .A2(n1346), .ZN(n1286) );
NAND2_X1 U1034 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
NOR2_X1 U1035 ( .A1(n1284), .A2(n1121), .ZN(n1096) );
XOR2_X1 U1036 ( .A(n1349), .B(n1199), .Z(n1121) );
INV_X1 U1037 ( .A(G475), .ZN(n1199) );
NAND2_X1 U1038 ( .A1(n1197), .A2(n1317), .ZN(n1349) );
XNOR2_X1 U1039 ( .A(n1350), .B(n1351), .ZN(n1197) );
XOR2_X1 U1040 ( .A(n1352), .B(n1353), .Z(n1351) );
XNOR2_X1 U1041 ( .A(n1354), .B(n1355), .ZN(n1353) );
AND2_X1 U1042 ( .A1(G214), .A2(n1356), .ZN(n1355) );
XNOR2_X1 U1043 ( .A(G104), .B(G113), .ZN(n1352) );
XOR2_X1 U1044 ( .A(n1357), .B(n1358), .Z(n1350) );
XNOR2_X1 U1045 ( .A(G140), .B(n1151), .ZN(n1358) );
INV_X1 U1046 ( .A(G131), .ZN(n1151) );
XNOR2_X1 U1047 ( .A(G122), .B(G125), .ZN(n1357) );
INV_X1 U1048 ( .A(n1309), .ZN(n1284) );
NOR2_X1 U1049 ( .A1(n1359), .A2(n1133), .ZN(n1309) );
NOR3_X1 U1050 ( .A1(n1130), .A2(G902), .A3(n1360), .ZN(n1133) );
INV_X1 U1051 ( .A(n1193), .ZN(n1130) );
AND2_X1 U1052 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NAND2_X1 U1053 ( .A1(n1193), .A2(n1317), .ZN(n1361) );
XNOR2_X1 U1054 ( .A(n1362), .B(n1363), .ZN(n1193) );
NOR2_X1 U1055 ( .A1(KEYINPUT53), .A2(n1364), .ZN(n1363) );
XOR2_X1 U1056 ( .A(n1365), .B(n1366), .Z(n1364) );
XNOR2_X1 U1057 ( .A(G128), .B(n1367), .ZN(n1366) );
NAND2_X1 U1058 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
XOR2_X1 U1059 ( .A(KEYINPUT62), .B(KEYINPUT25), .Z(n1369) );
XNOR2_X1 U1060 ( .A(G107), .B(n1370), .ZN(n1368) );
XNOR2_X1 U1061 ( .A(n1337), .B(G116), .ZN(n1370) );
INV_X1 U1062 ( .A(G122), .ZN(n1337) );
XNOR2_X1 U1063 ( .A(n1371), .B(G134), .ZN(n1365) );
INV_X1 U1064 ( .A(G143), .ZN(n1371) );
NAND2_X1 U1065 ( .A1(G217), .A2(n1372), .ZN(n1362) );
INV_X1 U1066 ( .A(n1129), .ZN(n1360) );
XOR2_X1 U1067 ( .A(G478), .B(KEYINPUT32), .Z(n1129) );
INV_X1 U1068 ( .A(n1111), .ZN(n1108) );
XNOR2_X1 U1069 ( .A(n1373), .B(n1190), .ZN(n1111) );
NAND2_X1 U1070 ( .A1(G217), .A2(n1100), .ZN(n1190) );
NAND2_X1 U1071 ( .A1(G234), .A2(n1347), .ZN(n1100) );
XNOR2_X1 U1072 ( .A(n1317), .B(KEYINPUT9), .ZN(n1347) );
NAND2_X1 U1073 ( .A1(n1317), .A2(n1188), .ZN(n1373) );
NAND2_X1 U1074 ( .A1(n1374), .A2(n1375), .ZN(n1188) );
NAND2_X1 U1075 ( .A1(n1376), .A2(n1377), .ZN(n1375) );
XOR2_X1 U1076 ( .A(n1378), .B(KEYINPUT4), .Z(n1374) );
OR2_X1 U1077 ( .A1(n1377), .A2(n1376), .ZN(n1378) );
XNOR2_X1 U1078 ( .A(n1379), .B(n1380), .ZN(n1376) );
XNOR2_X1 U1079 ( .A(n1163), .B(n1381), .ZN(n1380) );
XNOR2_X1 U1080 ( .A(G146), .B(n1288), .ZN(n1381) );
INV_X1 U1081 ( .A(G128), .ZN(n1288) );
INV_X1 U1082 ( .A(G125), .ZN(n1163) );
XOR2_X1 U1083 ( .A(n1382), .B(n1383), .Z(n1379) );
XOR2_X1 U1084 ( .A(n1384), .B(G110), .Z(n1382) );
NAND2_X1 U1085 ( .A1(KEYINPUT18), .A2(G140), .ZN(n1384) );
XOR2_X1 U1086 ( .A(n1385), .B(n1158), .Z(n1377) );
NAND2_X1 U1087 ( .A1(n1372), .A2(G221), .ZN(n1385) );
AND2_X1 U1088 ( .A1(G234), .A2(n1081), .ZN(n1372) );
XOR2_X1 U1089 ( .A(n1310), .B(KEYINPUT36), .Z(n1107) );
XNOR2_X1 U1090 ( .A(n1125), .B(G472), .ZN(n1310) );
AND3_X1 U1091 ( .A1(n1386), .A2(n1387), .A3(n1317), .ZN(n1125) );
INV_X1 U1092 ( .A(G902), .ZN(n1317) );
NAND2_X1 U1093 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
NAND2_X1 U1094 ( .A1(n1390), .A2(n1391), .ZN(n1388) );
NAND2_X1 U1095 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
NAND2_X1 U1096 ( .A1(n1394), .A2(n1395), .ZN(n1390) );
INV_X1 U1097 ( .A(n1392), .ZN(n1395) );
XOR2_X1 U1098 ( .A(G101), .B(KEYINPUT60), .Z(n1392) );
NAND2_X1 U1099 ( .A1(n1205), .A2(n1396), .ZN(n1386) );
NAND2_X1 U1100 ( .A1(n1397), .A2(n1398), .ZN(n1396) );
NAND2_X1 U1101 ( .A1(n1399), .A2(n1393), .ZN(n1398) );
NAND2_X1 U1102 ( .A1(n1394), .A2(n1400), .ZN(n1397) );
INV_X1 U1103 ( .A(n1399), .ZN(n1400) );
XOR2_X1 U1104 ( .A(G101), .B(KEYINPUT39), .Z(n1399) );
XNOR2_X1 U1105 ( .A(n1393), .B(KEYINPUT48), .ZN(n1394) );
XOR2_X1 U1106 ( .A(n1401), .B(n1210), .Z(n1393) );
XOR2_X1 U1107 ( .A(G113), .B(n1402), .Z(n1210) );
NOR2_X1 U1108 ( .A1(KEYINPUT23), .A2(n1343), .ZN(n1402) );
XOR2_X1 U1109 ( .A(G116), .B(n1383), .Z(n1343) );
XOR2_X1 U1110 ( .A(G119), .B(KEYINPUT13), .Z(n1383) );
XNOR2_X1 U1111 ( .A(n1403), .B(n1222), .ZN(n1401) );
INV_X1 U1112 ( .A(n1216), .ZN(n1222) );
XNOR2_X1 U1113 ( .A(n1404), .B(n1405), .ZN(n1216) );
XOR2_X1 U1114 ( .A(KEYINPUT34), .B(n1406), .Z(n1405) );
XOR2_X1 U1115 ( .A(KEYINPUT49), .B(KEYINPUT46), .Z(n1406) );
XNOR2_X1 U1116 ( .A(G131), .B(n1407), .ZN(n1404) );
XNOR2_X1 U1117 ( .A(n1158), .B(G134), .ZN(n1407) );
INV_X1 U1118 ( .A(G137), .ZN(n1158) );
NAND2_X1 U1119 ( .A1(KEYINPUT52), .A2(n1408), .ZN(n1403) );
INV_X1 U1120 ( .A(n1215), .ZN(n1408) );
XOR2_X1 U1121 ( .A(G128), .B(n1409), .Z(n1215) );
NOR2_X1 U1122 ( .A1(KEYINPUT51), .A2(n1410), .ZN(n1409) );
XNOR2_X1 U1123 ( .A(n1411), .B(n1328), .ZN(n1410) );
INV_X1 U1124 ( .A(n1354), .ZN(n1328) );
XOR2_X1 U1125 ( .A(G143), .B(G146), .Z(n1354) );
XNOR2_X1 U1126 ( .A(KEYINPUT20), .B(KEYINPUT17), .ZN(n1411) );
INV_X1 U1127 ( .A(n1389), .ZN(n1205) );
NAND2_X1 U1128 ( .A1(n1356), .A2(G210), .ZN(n1389) );
AND2_X1 U1129 ( .A1(n1412), .A2(n1081), .ZN(n1356) );
INV_X1 U1130 ( .A(G953), .ZN(n1081) );
XNOR2_X1 U1131 ( .A(KEYINPUT0), .B(n1348), .ZN(n1412) );
INV_X1 U1132 ( .A(G237), .ZN(n1348) );
endmodule


