//Key = 1100110001011100111111100001101000100101010010110101101110101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378;

XNOR2_X1 U752 ( .A(G125), .B(G140), .ZN(n1034) );
NAND2_X1 U753 ( .A1(n1035), .A2(n1036), .ZN(G9) );
OR2_X1 U754 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
XOR2_X1 U755 ( .A(n1039), .B(KEYINPUT42), .Z(n1035) );
NAND2_X1 U756 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
NOR2_X1 U757 ( .A1(n1040), .A2(n1041), .ZN(G75) );
NOR4_X1 U758 ( .A1(G953), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1041) );
NOR2_X1 U759 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U760 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U761 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U762 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U763 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
INV_X1 U764 ( .A(n1055), .ZN(n1054) );
NOR3_X1 U765 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1053) );
NOR2_X1 U766 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR2_X1 U767 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR2_X1 U768 ( .A1(n1063), .A2(n1064), .ZN(n1057) );
XNOR2_X1 U769 ( .A(n1065), .B(KEYINPUT31), .ZN(n1063) );
NOR2_X1 U770 ( .A1(n1066), .A2(n1067), .ZN(n1056) );
NOR3_X1 U771 ( .A1(n1060), .A2(n1068), .A3(n1067), .ZN(n1051) );
NOR4_X1 U772 ( .A1(n1069), .A2(n1070), .A3(n1067), .A4(n1060), .ZN(n1047) );
NOR2_X1 U773 ( .A1(n1071), .A2(n1055), .ZN(n1070) );
NOR2_X1 U774 ( .A1(n1072), .A2(n1050), .ZN(n1071) );
NOR3_X1 U775 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1069) );
NOR2_X1 U776 ( .A1(n1076), .A2(n1077), .ZN(n1073) );
NOR3_X1 U777 ( .A1(n1042), .A2(G953), .A3(G952), .ZN(n1040) );
AND4_X1 U778 ( .A1(n1078), .A2(n1055), .A3(n1079), .A4(n1080), .ZN(n1042) );
NOR4_X1 U779 ( .A1(n1081), .A2(n1082), .A3(n1050), .A4(n1083), .ZN(n1080) );
AND2_X1 U780 ( .A1(n1084), .A2(KEYINPUT32), .ZN(n1081) );
XOR2_X1 U781 ( .A(n1085), .B(n1086), .Z(n1079) );
NOR2_X1 U782 ( .A1(KEYINPUT32), .A2(n1084), .ZN(n1086) );
XNOR2_X1 U783 ( .A(n1087), .B(KEYINPUT24), .ZN(n1078) );
XOR2_X1 U784 ( .A(n1088), .B(n1089), .Z(G72) );
NOR2_X1 U785 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U786 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NOR2_X1 U787 ( .A1(KEYINPUT59), .A2(n1094), .ZN(n1088) );
XOR2_X1 U788 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR3_X1 U789 ( .A1(n1097), .A2(KEYINPUT15), .A3(G953), .ZN(n1096) );
NOR2_X1 U790 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XNOR2_X1 U791 ( .A(n1100), .B(KEYINPUT52), .ZN(n1098) );
NAND4_X1 U792 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1095) );
NAND2_X1 U793 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
INV_X1 U794 ( .A(KEYINPUT55), .ZN(n1106) );
NAND2_X1 U795 ( .A1(n1034), .A2(n1107), .ZN(n1105) );
XNOR2_X1 U796 ( .A(KEYINPUT0), .B(n1108), .ZN(n1107) );
NAND2_X1 U797 ( .A1(KEYINPUT55), .A2(n1109), .ZN(n1103) );
NAND2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND3_X1 U799 ( .A1(KEYINPUT0), .A2(n1034), .A3(n1108), .ZN(n1111) );
OR2_X1 U800 ( .A1(n1108), .A2(KEYINPUT0), .ZN(n1110) );
OR2_X1 U801 ( .A1(n1108), .A2(n1034), .ZN(n1102) );
XOR2_X1 U802 ( .A(n1112), .B(n1113), .Z(n1108) );
XOR2_X1 U803 ( .A(G131), .B(n1114), .Z(n1113) );
XOR2_X1 U804 ( .A(KEYINPUT56), .B(G137), .Z(n1114) );
XOR2_X1 U805 ( .A(n1115), .B(n1116), .Z(n1112) );
NAND2_X1 U806 ( .A1(G953), .A2(n1093), .ZN(n1101) );
NAND2_X1 U807 ( .A1(n1117), .A2(n1118), .ZN(G69) );
NAND2_X1 U808 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U809 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U810 ( .A1(G953), .A2(n1123), .ZN(n1122) );
INV_X1 U811 ( .A(n1124), .ZN(n1121) );
NAND2_X1 U812 ( .A1(n1125), .A2(n1126), .ZN(n1117) );
NAND2_X1 U813 ( .A1(G953), .A2(n1127), .ZN(n1126) );
NAND2_X1 U814 ( .A1(G898), .A2(G224), .ZN(n1127) );
INV_X1 U815 ( .A(n1119), .ZN(n1125) );
XNOR2_X1 U816 ( .A(n1128), .B(n1129), .ZN(n1119) );
NOR2_X1 U817 ( .A1(n1124), .A2(n1130), .ZN(n1129) );
XNOR2_X1 U818 ( .A(n1131), .B(n1132), .ZN(n1130) );
XOR2_X1 U819 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U820 ( .A1(KEYINPUT22), .A2(n1135), .ZN(n1133) );
INV_X1 U821 ( .A(n1136), .ZN(n1135) );
NAND2_X1 U822 ( .A1(KEYINPUT21), .A2(n1137), .ZN(n1128) );
NAND2_X1 U823 ( .A1(n1138), .A2(n1091), .ZN(n1137) );
NOR2_X1 U824 ( .A1(n1139), .A2(n1140), .ZN(G66) );
XNOR2_X1 U825 ( .A(n1141), .B(n1142), .ZN(n1140) );
NOR2_X1 U826 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U827 ( .A(n1145), .B(KEYINPUT14), .Z(n1143) );
NOR2_X1 U828 ( .A1(n1139), .A2(n1146), .ZN(G63) );
XNOR2_X1 U829 ( .A(n1147), .B(n1148), .ZN(n1146) );
NOR2_X1 U830 ( .A1(n1084), .A2(n1144), .ZN(n1148) );
NOR2_X1 U831 ( .A1(n1139), .A2(n1149), .ZN(G60) );
XOR2_X1 U832 ( .A(n1150), .B(n1151), .Z(n1149) );
AND2_X1 U833 ( .A1(G475), .A2(n1152), .ZN(n1150) );
XNOR2_X1 U834 ( .A(n1153), .B(n1154), .ZN(G6) );
NOR2_X1 U835 ( .A1(n1155), .A2(n1156), .ZN(G57) );
XOR2_X1 U836 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U837 ( .A(G101), .B(n1159), .ZN(n1158) );
NAND3_X1 U838 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1157) );
NAND3_X1 U839 ( .A1(G472), .A2(n1163), .A3(n1152), .ZN(n1162) );
NAND2_X1 U840 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U841 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NAND3_X1 U842 ( .A1(n1168), .A2(n1169), .A3(n1164), .ZN(n1161) );
INV_X1 U843 ( .A(KEYINPUT7), .ZN(n1164) );
NAND3_X1 U844 ( .A1(G472), .A2(n1167), .A3(n1152), .ZN(n1168) );
INV_X1 U845 ( .A(KEYINPUT8), .ZN(n1167) );
NAND2_X1 U846 ( .A1(KEYINPUT7), .A2(n1166), .ZN(n1160) );
INV_X1 U847 ( .A(n1169), .ZN(n1166) );
NAND2_X1 U848 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NAND2_X1 U849 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XOR2_X1 U850 ( .A(KEYINPUT16), .B(n1174), .Z(n1173) );
XOR2_X1 U851 ( .A(KEYINPUT51), .B(n1175), .Z(n1172) );
XOR2_X1 U852 ( .A(n1176), .B(KEYINPUT50), .Z(n1170) );
NAND2_X1 U853 ( .A1(n1174), .A2(n1175), .ZN(n1176) );
NOR2_X1 U854 ( .A1(n1177), .A2(n1091), .ZN(n1155) );
XNOR2_X1 U855 ( .A(G952), .B(KEYINPUT39), .ZN(n1177) );
NOR2_X1 U856 ( .A1(n1139), .A2(n1178), .ZN(G54) );
XOR2_X1 U857 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U858 ( .A(n1181), .B(n1182), .Z(n1180) );
NAND3_X1 U859 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1181) );
NAND2_X1 U860 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NAND2_X1 U861 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XNOR2_X1 U862 ( .A(n1115), .B(n1190), .ZN(n1186) );
OR2_X1 U863 ( .A1(n1191), .A2(n1188), .ZN(n1184) );
NAND4_X1 U864 ( .A1(n1189), .A2(n1191), .A3(n1192), .A4(n1188), .ZN(n1183) );
XOR2_X1 U865 ( .A(n1193), .B(KEYINPUT34), .Z(n1188) );
XNOR2_X1 U866 ( .A(n1115), .B(n1131), .ZN(n1192) );
INV_X1 U867 ( .A(n1190), .ZN(n1131) );
INV_X1 U868 ( .A(KEYINPUT36), .ZN(n1191) );
INV_X1 U869 ( .A(KEYINPUT26), .ZN(n1189) );
XNOR2_X1 U870 ( .A(n1194), .B(n1195), .ZN(n1179) );
AND2_X1 U871 ( .A1(G469), .A2(n1152), .ZN(n1195) );
INV_X1 U872 ( .A(n1144), .ZN(n1152) );
NOR2_X1 U873 ( .A1(n1139), .A2(n1196), .ZN(G51) );
XOR2_X1 U874 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U875 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U876 ( .A1(n1201), .A2(n1144), .ZN(n1199) );
NAND2_X1 U877 ( .A1(n1202), .A2(n1044), .ZN(n1144) );
OR3_X1 U878 ( .A1(n1099), .A2(n1100), .A3(n1138), .ZN(n1044) );
NAND4_X1 U879 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1138) );
NOR4_X1 U880 ( .A1(n1207), .A2(n1208), .A3(n1154), .A4(n1038), .ZN(n1206) );
NOR3_X1 U881 ( .A1(n1067), .A2(n1066), .A3(n1209), .ZN(n1038) );
NOR3_X1 U882 ( .A1(n1209), .A2(n1067), .A3(n1064), .ZN(n1154) );
INV_X1 U883 ( .A(n1210), .ZN(n1064) );
INV_X1 U884 ( .A(n1065), .ZN(n1067) );
NOR2_X1 U885 ( .A1(n1211), .A2(n1212), .ZN(n1205) );
INV_X1 U886 ( .A(n1213), .ZN(n1212) );
NAND4_X1 U887 ( .A1(n1062), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1204) );
NAND2_X1 U888 ( .A1(KEYINPUT44), .A2(n1209), .ZN(n1216) );
NAND2_X1 U889 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
INV_X1 U890 ( .A(KEYINPUT44), .ZN(n1218) );
NAND2_X1 U891 ( .A1(n1219), .A2(n1068), .ZN(n1217) );
NAND3_X1 U892 ( .A1(n1220), .A2(n1061), .A3(n1210), .ZN(n1203) );
INV_X1 U893 ( .A(n1221), .ZN(n1100) );
NAND4_X1 U894 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1099) );
NOR3_X1 U895 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1225) );
NAND2_X1 U896 ( .A1(n1229), .A2(n1230), .ZN(n1224) );
NAND2_X1 U897 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND2_X1 U898 ( .A1(n1061), .A2(n1233), .ZN(n1232) );
NAND2_X1 U899 ( .A1(n1062), .A2(n1210), .ZN(n1231) );
XNOR2_X1 U900 ( .A(G902), .B(KEYINPUT28), .ZN(n1202) );
NAND2_X1 U901 ( .A1(n1234), .A2(n1235), .ZN(n1197) );
NAND2_X1 U902 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
INV_X1 U903 ( .A(n1238), .ZN(n1237) );
XOR2_X1 U904 ( .A(KEYINPUT58), .B(n1239), .Z(n1236) );
NAND2_X1 U905 ( .A1(n1238), .A2(n1240), .ZN(n1234) );
XNOR2_X1 U906 ( .A(n1239), .B(KEYINPUT18), .ZN(n1240) );
NOR2_X1 U907 ( .A1(n1091), .A2(G952), .ZN(n1139) );
XNOR2_X1 U908 ( .A(n1227), .B(n1241), .ZN(G48) );
NAND2_X1 U909 ( .A1(KEYINPUT11), .A2(G146), .ZN(n1241) );
AND2_X1 U910 ( .A1(n1242), .A2(n1210), .ZN(n1227) );
XNOR2_X1 U911 ( .A(G143), .B(n1221), .ZN(G45) );
NAND4_X1 U912 ( .A1(n1243), .A2(n1061), .A3(n1244), .A4(n1074), .ZN(n1221) );
NOR2_X1 U913 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
XNOR2_X1 U914 ( .A(G140), .B(n1247), .ZN(G42) );
NAND4_X1 U915 ( .A1(n1248), .A2(n1062), .A3(n1210), .A4(n1243), .ZN(n1247) );
XNOR2_X1 U916 ( .A(n1249), .B(KEYINPUT60), .ZN(n1248) );
XNOR2_X1 U917 ( .A(G137), .B(n1222), .ZN(G39) );
NAND2_X1 U918 ( .A1(n1229), .A2(n1250), .ZN(n1222) );
XNOR2_X1 U919 ( .A(G134), .B(n1251), .ZN(G36) );
NAND2_X1 U920 ( .A1(n1249), .A2(n1252), .ZN(n1251) );
XOR2_X1 U921 ( .A(KEYINPUT23), .B(n1253), .Z(n1252) );
NOR4_X1 U922 ( .A1(n1254), .A2(n1255), .A3(n1066), .A4(n1256), .ZN(n1253) );
INV_X1 U923 ( .A(n1233), .ZN(n1066) );
XNOR2_X1 U924 ( .A(n1257), .B(KEYINPUT38), .ZN(n1255) );
AND2_X1 U925 ( .A1(n1046), .A2(n1258), .ZN(n1254) );
XNOR2_X1 U926 ( .A(G131), .B(n1223), .ZN(G33) );
NAND3_X1 U927 ( .A1(n1210), .A2(n1061), .A3(n1229), .ZN(n1223) );
AND2_X1 U928 ( .A1(n1243), .A2(n1249), .ZN(n1229) );
INV_X1 U929 ( .A(n1050), .ZN(n1249) );
NAND2_X1 U930 ( .A1(n1259), .A2(n1077), .ZN(n1050) );
INV_X1 U931 ( .A(n1076), .ZN(n1259) );
XNOR2_X1 U932 ( .A(n1260), .B(n1226), .ZN(G30) );
AND2_X1 U933 ( .A1(n1242), .A2(n1233), .ZN(n1226) );
AND4_X1 U934 ( .A1(n1243), .A2(n1074), .A3(n1087), .A4(n1082), .ZN(n1242) );
AND2_X1 U935 ( .A1(n1257), .A2(n1261), .ZN(n1243) );
XNOR2_X1 U936 ( .A(n1262), .B(n1208), .ZN(G3) );
NOR3_X1 U937 ( .A1(n1256), .A2(n1209), .A3(n1060), .ZN(n1208) );
INV_X1 U938 ( .A(n1214), .ZN(n1060) );
XNOR2_X1 U939 ( .A(n1263), .B(n1228), .ZN(G27) );
AND3_X1 U940 ( .A1(n1062), .A2(n1261), .A3(n1264), .ZN(n1228) );
INV_X1 U941 ( .A(n1265), .ZN(n1264) );
NAND2_X1 U942 ( .A1(n1258), .A2(n1046), .ZN(n1261) );
NAND4_X1 U943 ( .A1(n1266), .A2(G902), .A3(n1267), .A4(n1093), .ZN(n1258) );
INV_X1 U944 ( .A(G900), .ZN(n1093) );
XNOR2_X1 U945 ( .A(G953), .B(KEYINPUT47), .ZN(n1266) );
XNOR2_X1 U946 ( .A(G122), .B(n1213), .ZN(G24) );
NAND4_X1 U947 ( .A1(n1220), .A2(n1065), .A3(n1268), .A4(n1269), .ZN(n1213) );
NOR2_X1 U948 ( .A1(n1082), .A2(n1087), .ZN(n1065) );
XOR2_X1 U949 ( .A(G119), .B(n1211), .Z(G21) );
AND2_X1 U950 ( .A1(n1250), .A2(n1220), .ZN(n1211) );
AND3_X1 U951 ( .A1(n1087), .A2(n1082), .A3(n1214), .ZN(n1250) );
XOR2_X1 U952 ( .A(G116), .B(n1207), .Z(G18) );
AND3_X1 U953 ( .A1(n1061), .A2(n1233), .A3(n1220), .ZN(n1207) );
AND2_X1 U954 ( .A1(n1055), .A2(n1219), .ZN(n1220) );
NOR2_X1 U955 ( .A1(n1083), .A2(n1245), .ZN(n1233) );
INV_X1 U956 ( .A(n1269), .ZN(n1245) );
XNOR2_X1 U957 ( .A(n1270), .B(n1271), .ZN(G15) );
NOR3_X1 U958 ( .A1(n1265), .A2(n1272), .A3(n1256), .ZN(n1271) );
INV_X1 U959 ( .A(n1061), .ZN(n1256) );
NOR2_X1 U960 ( .A1(n1082), .A2(n1273), .ZN(n1061) );
XOR2_X1 U961 ( .A(n1274), .B(KEYINPUT37), .Z(n1272) );
NAND3_X1 U962 ( .A1(n1055), .A2(n1074), .A3(n1210), .ZN(n1265) );
NOR2_X1 U963 ( .A1(n1269), .A2(n1246), .ZN(n1210) );
INV_X1 U964 ( .A(n1268), .ZN(n1246) );
XOR2_X1 U965 ( .A(n1083), .B(KEYINPUT63), .Z(n1268) );
NOR2_X1 U966 ( .A1(n1072), .A2(n1075), .ZN(n1055) );
INV_X1 U967 ( .A(n1275), .ZN(n1075) );
XNOR2_X1 U968 ( .A(G110), .B(n1276), .ZN(G12) );
NAND3_X1 U969 ( .A1(n1214), .A2(n1277), .A3(n1062), .ZN(n1276) );
AND2_X1 U970 ( .A1(n1273), .A2(n1082), .ZN(n1062) );
XOR2_X1 U971 ( .A(n1278), .B(n1145), .Z(n1082) );
NAND2_X1 U972 ( .A1(G217), .A2(n1279), .ZN(n1145) );
NAND2_X1 U973 ( .A1(n1141), .A2(n1280), .ZN(n1278) );
XNOR2_X1 U974 ( .A(n1281), .B(n1282), .ZN(n1141) );
XNOR2_X1 U975 ( .A(G137), .B(n1283), .ZN(n1282) );
NAND2_X1 U976 ( .A1(n1284), .A2(G221), .ZN(n1283) );
NAND2_X1 U977 ( .A1(n1285), .A2(KEYINPUT5), .ZN(n1281) );
XOR2_X1 U978 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U979 ( .A(G146), .B(n1194), .ZN(n1287) );
XNOR2_X1 U980 ( .A(n1288), .B(n1034), .ZN(n1286) );
NAND2_X1 U981 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
NAND2_X1 U982 ( .A1(G119), .A2(n1260), .ZN(n1290) );
XOR2_X1 U983 ( .A(KEYINPUT13), .B(n1291), .Z(n1289) );
NOR2_X1 U984 ( .A1(G119), .A2(n1260), .ZN(n1291) );
INV_X1 U985 ( .A(n1087), .ZN(n1273) );
XNOR2_X1 U986 ( .A(n1292), .B(G472), .ZN(n1087) );
NAND3_X1 U987 ( .A1(n1293), .A2(n1280), .A3(n1294), .ZN(n1292) );
NAND3_X1 U988 ( .A1(n1262), .A2(n1295), .A3(n1296), .ZN(n1294) );
XOR2_X1 U989 ( .A(n1297), .B(n1298), .Z(n1296) );
NOR2_X1 U990 ( .A1(n1299), .A2(n1159), .ZN(n1298) );
INV_X1 U991 ( .A(KEYINPUT4), .ZN(n1299) );
NAND2_X1 U992 ( .A1(n1300), .A2(n1301), .ZN(n1293) );
NAND2_X1 U993 ( .A1(n1262), .A2(n1295), .ZN(n1301) );
INV_X1 U994 ( .A(KEYINPUT62), .ZN(n1295) );
INV_X1 U995 ( .A(G101), .ZN(n1262) );
XOR2_X1 U996 ( .A(n1297), .B(n1302), .Z(n1300) );
AND2_X1 U997 ( .A1(n1159), .A2(KEYINPUT4), .ZN(n1302) );
NAND2_X1 U998 ( .A1(n1303), .A2(G210), .ZN(n1159) );
XNOR2_X1 U999 ( .A(n1175), .B(n1174), .ZN(n1297) );
XNOR2_X1 U1000 ( .A(n1304), .B(n1305), .ZN(n1174) );
NOR2_X1 U1001 ( .A1(G119), .A2(KEYINPUT57), .ZN(n1305) );
XNOR2_X1 U1002 ( .A(G113), .B(G116), .ZN(n1304) );
XOR2_X1 U1003 ( .A(n1193), .B(n1306), .Z(n1175) );
INV_X1 U1004 ( .A(n1209), .ZN(n1277) );
NAND2_X1 U1005 ( .A1(n1257), .A2(n1219), .ZN(n1209) );
AND2_X1 U1006 ( .A1(n1074), .A2(n1274), .ZN(n1219) );
NAND2_X1 U1007 ( .A1(n1046), .A2(n1307), .ZN(n1274) );
NAND3_X1 U1008 ( .A1(G902), .A2(n1267), .A3(n1124), .ZN(n1307) );
NOR2_X1 U1009 ( .A1(n1091), .A2(G898), .ZN(n1124) );
NAND3_X1 U1010 ( .A1(n1267), .A2(n1091), .A3(G952), .ZN(n1046) );
NAND2_X1 U1011 ( .A1(G237), .A2(G234), .ZN(n1267) );
AND2_X1 U1012 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NAND2_X1 U1013 ( .A1(G214), .A2(n1308), .ZN(n1077) );
XOR2_X1 U1014 ( .A(n1309), .B(n1201), .Z(n1076) );
NAND2_X1 U1015 ( .A1(G210), .A2(n1308), .ZN(n1201) );
NAND2_X1 U1016 ( .A1(n1310), .A2(n1280), .ZN(n1308) );
INV_X1 U1017 ( .A(G237), .ZN(n1310) );
NAND2_X1 U1018 ( .A1(n1311), .A2(n1280), .ZN(n1309) );
XOR2_X1 U1019 ( .A(n1200), .B(n1312), .Z(n1311) );
XNOR2_X1 U1020 ( .A(n1313), .B(n1238), .ZN(n1312) );
XOR2_X1 U1021 ( .A(G125), .B(n1306), .Z(n1238) );
XNOR2_X1 U1022 ( .A(n1260), .B(n1314), .ZN(n1306) );
NOR2_X1 U1023 ( .A1(KEYINPUT53), .A2(n1315), .ZN(n1314) );
XNOR2_X1 U1024 ( .A(G143), .B(G146), .ZN(n1315) );
NAND2_X1 U1025 ( .A1(KEYINPUT19), .A2(n1239), .ZN(n1313) );
NOR2_X1 U1026 ( .A1(n1123), .A2(G953), .ZN(n1239) );
INV_X1 U1027 ( .A(G224), .ZN(n1123) );
XNOR2_X1 U1028 ( .A(n1316), .B(n1317), .ZN(n1200) );
XNOR2_X1 U1029 ( .A(n1318), .B(KEYINPUT33), .ZN(n1317) );
NAND2_X1 U1030 ( .A1(KEYINPUT41), .A2(n1134), .ZN(n1318) );
XOR2_X1 U1031 ( .A(n1319), .B(n1320), .Z(n1134) );
XOR2_X1 U1032 ( .A(G119), .B(G116), .Z(n1320) );
NAND2_X1 U1033 ( .A1(KEYINPUT9), .A2(n1270), .ZN(n1319) );
INV_X1 U1034 ( .A(G113), .ZN(n1270) );
XNOR2_X1 U1035 ( .A(n1190), .B(n1136), .ZN(n1316) );
XNOR2_X1 U1036 ( .A(G110), .B(n1321), .ZN(n1136) );
INV_X1 U1037 ( .A(n1068), .ZN(n1257) );
NAND2_X1 U1038 ( .A1(n1072), .A2(n1275), .ZN(n1068) );
NAND2_X1 U1039 ( .A1(G221), .A2(n1279), .ZN(n1275) );
NAND2_X1 U1040 ( .A1(G234), .A2(n1280), .ZN(n1279) );
XNOR2_X1 U1041 ( .A(n1322), .B(G469), .ZN(n1072) );
NAND2_X1 U1042 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1043 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1044 ( .A(n1182), .B(n1327), .Z(n1326) );
XNOR2_X1 U1045 ( .A(n1190), .B(n1328), .ZN(n1327) );
NOR2_X1 U1046 ( .A1(KEYINPUT6), .A2(n1115), .ZN(n1328) );
NAND2_X1 U1047 ( .A1(n1329), .A2(n1330), .ZN(n1115) );
NAND2_X1 U1048 ( .A1(G128), .A2(n1331), .ZN(n1330) );
XOR2_X1 U1049 ( .A(KEYINPUT61), .B(n1332), .Z(n1329) );
NOR2_X1 U1050 ( .A1(G128), .A2(n1331), .ZN(n1332) );
XOR2_X1 U1051 ( .A(n1333), .B(G146), .Z(n1331) );
NAND2_X1 U1052 ( .A1(KEYINPUT12), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1053 ( .A(G101), .B(n1335), .Z(n1190) );
XNOR2_X1 U1054 ( .A(n1037), .B(G104), .ZN(n1335) );
XNOR2_X1 U1055 ( .A(G140), .B(n1336), .ZN(n1182) );
NOR2_X1 U1056 ( .A1(G953), .A2(n1092), .ZN(n1336) );
INV_X1 U1057 ( .A(G227), .ZN(n1092) );
XOR2_X1 U1058 ( .A(n1337), .B(n1338), .Z(n1325) );
XNOR2_X1 U1059 ( .A(KEYINPUT46), .B(n1339), .ZN(n1338) );
NOR2_X1 U1060 ( .A1(KEYINPUT45), .A2(n1193), .ZN(n1339) );
XNOR2_X1 U1061 ( .A(n1340), .B(n1341), .ZN(n1193) );
XOR2_X1 U1062 ( .A(n1342), .B(n1116), .Z(n1341) );
XOR2_X1 U1063 ( .A(G134), .B(KEYINPUT29), .Z(n1116) );
NOR2_X1 U1064 ( .A1(G137), .A2(KEYINPUT10), .ZN(n1342) );
XOR2_X1 U1065 ( .A(n1343), .B(G131), .Z(n1340) );
XNOR2_X1 U1066 ( .A(KEYINPUT43), .B(KEYINPUT3), .ZN(n1343) );
NAND2_X1 U1067 ( .A1(KEYINPUT49), .A2(n1194), .ZN(n1337) );
INV_X1 U1068 ( .A(G110), .ZN(n1194) );
XNOR2_X1 U1069 ( .A(KEYINPUT54), .B(n1280), .ZN(n1323) );
NOR2_X1 U1070 ( .A1(n1269), .A2(n1083), .ZN(n1214) );
XNOR2_X1 U1071 ( .A(n1344), .B(G475), .ZN(n1083) );
OR2_X1 U1072 ( .A1(n1151), .A2(G902), .ZN(n1344) );
XNOR2_X1 U1073 ( .A(n1345), .B(n1346), .ZN(n1151) );
XOR2_X1 U1074 ( .A(n1347), .B(n1348), .Z(n1346) );
XNOR2_X1 U1075 ( .A(n1321), .B(G113), .ZN(n1348) );
INV_X1 U1076 ( .A(G122), .ZN(n1321) );
XOR2_X1 U1077 ( .A(G146), .B(G131), .Z(n1347) );
XOR2_X1 U1078 ( .A(n1349), .B(n1350), .Z(n1345) );
XOR2_X1 U1079 ( .A(n1351), .B(n1352), .Z(n1350) );
NAND2_X1 U1080 ( .A1(KEYINPUT27), .A2(n1153), .ZN(n1352) );
INV_X1 U1081 ( .A(G104), .ZN(n1153) );
NAND2_X1 U1082 ( .A1(n1353), .A2(n1354), .ZN(n1351) );
OR2_X1 U1083 ( .A1(n1263), .A2(G140), .ZN(n1354) );
XOR2_X1 U1084 ( .A(n1355), .B(KEYINPUT40), .Z(n1353) );
NAND2_X1 U1085 ( .A1(G140), .A2(n1263), .ZN(n1355) );
INV_X1 U1086 ( .A(G125), .ZN(n1263) );
XOR2_X1 U1087 ( .A(n1356), .B(n1357), .Z(n1349) );
NOR2_X1 U1088 ( .A1(KEYINPUT35), .A2(G143), .ZN(n1357) );
NAND2_X1 U1089 ( .A1(n1303), .A2(G214), .ZN(n1356) );
NOR2_X1 U1090 ( .A1(G953), .A2(G237), .ZN(n1303) );
NAND3_X1 U1091 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1269) );
NAND2_X1 U1092 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
NAND2_X1 U1093 ( .A1(KEYINPUT17), .A2(n1363), .ZN(n1362) );
XNOR2_X1 U1094 ( .A(KEYINPUT20), .B(n1084), .ZN(n1363) );
NAND3_X1 U1095 ( .A1(KEYINPUT17), .A2(n1364), .A3(n1084), .ZN(n1359) );
INV_X1 U1096 ( .A(n1361), .ZN(n1364) );
XNOR2_X1 U1097 ( .A(n1085), .B(KEYINPUT1), .ZN(n1361) );
NAND2_X1 U1098 ( .A1(n1280), .A2(n1147), .ZN(n1085) );
NAND2_X1 U1099 ( .A1(n1365), .A2(n1366), .ZN(n1147) );
NAND2_X1 U1100 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
NAND2_X1 U1101 ( .A1(n1284), .A2(G217), .ZN(n1368) );
INV_X1 U1102 ( .A(n1369), .ZN(n1284) );
XOR2_X1 U1103 ( .A(KEYINPUT30), .B(n1370), .Z(n1365) );
NOR3_X1 U1104 ( .A1(n1367), .A2(n1371), .A3(n1369), .ZN(n1370) );
NAND2_X1 U1105 ( .A1(G234), .A2(n1091), .ZN(n1369) );
INV_X1 U1106 ( .A(G953), .ZN(n1091) );
INV_X1 U1107 ( .A(G217), .ZN(n1371) );
XNOR2_X1 U1108 ( .A(n1372), .B(n1373), .ZN(n1367) );
XOR2_X1 U1109 ( .A(n1374), .B(n1375), .Z(n1373) );
XNOR2_X1 U1110 ( .A(n1037), .B(n1376), .ZN(n1375) );
NOR2_X1 U1111 ( .A1(KEYINPUT48), .A2(n1377), .ZN(n1376) );
XNOR2_X1 U1112 ( .A(KEYINPUT2), .B(n1334), .ZN(n1377) );
INV_X1 U1113 ( .A(G143), .ZN(n1334) );
INV_X1 U1114 ( .A(G107), .ZN(n1037) );
NOR2_X1 U1115 ( .A1(G116), .A2(KEYINPUT25), .ZN(n1374) );
XNOR2_X1 U1116 ( .A(G122), .B(n1378), .ZN(n1372) );
XNOR2_X1 U1117 ( .A(G134), .B(n1260), .ZN(n1378) );
INV_X1 U1118 ( .A(G128), .ZN(n1260) );
INV_X1 U1119 ( .A(G902), .ZN(n1280) );
OR2_X1 U1120 ( .A1(n1084), .A2(KEYINPUT17), .ZN(n1358) );
INV_X1 U1121 ( .A(G478), .ZN(n1084) );
endmodule


