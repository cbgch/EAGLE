//Key = 0111000111101001010000100101100001001110111110011101010100110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270;

XNOR2_X1 U697 ( .A(G107), .B(n969), .ZN(G9) );
NOR2_X1 U698 ( .A1(n970), .A2(n971), .ZN(G75) );
NOR4_X1 U699 ( .A1(n972), .A2(n973), .A3(n974), .A4(n975), .ZN(n971) );
NAND4_X1 U700 ( .A1(n976), .A2(n977), .A3(n978), .A4(n979), .ZN(n972) );
NAND2_X1 U701 ( .A1(n980), .A2(n981), .ZN(n977) );
NAND2_X1 U702 ( .A1(n982), .A2(n983), .ZN(n981) );
NAND4_X1 U703 ( .A1(n984), .A2(n985), .A3(n986), .A4(n987), .ZN(n983) );
NAND3_X1 U704 ( .A1(n988), .A2(n989), .A3(n990), .ZN(n987) );
NAND2_X1 U705 ( .A1(n991), .A2(n992), .ZN(n990) );
OR2_X1 U706 ( .A1(n993), .A2(n994), .ZN(n992) );
NAND2_X1 U707 ( .A1(n995), .A2(n996), .ZN(n989) );
NAND3_X1 U708 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n996) );
NAND2_X1 U709 ( .A1(KEYINPUT44), .A2(n1000), .ZN(n999) );
OR3_X1 U710 ( .A1(n1001), .A2(n1002), .A3(KEYINPUT19), .ZN(n998) );
NAND2_X1 U711 ( .A1(KEYINPUT19), .A2(n991), .ZN(n997) );
NAND3_X1 U712 ( .A1(n1000), .A2(n1003), .A3(n1004), .ZN(n988) );
INV_X1 U713 ( .A(KEYINPUT44), .ZN(n1003) );
NAND3_X1 U714 ( .A1(n991), .A2(n1005), .A3(n995), .ZN(n982) );
NAND2_X1 U715 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NAND3_X1 U716 ( .A1(n1008), .A2(n1009), .A3(n986), .ZN(n1007) );
NAND2_X1 U717 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND3_X1 U718 ( .A1(n1012), .A2(n1013), .A3(n984), .ZN(n1008) );
NAND2_X1 U719 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NAND2_X1 U720 ( .A1(n1016), .A2(n985), .ZN(n1006) );
INV_X1 U721 ( .A(n1017), .ZN(n980) );
NOR3_X1 U722 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n970) );
XOR2_X1 U723 ( .A(n974), .B(KEYINPUT37), .Z(n1020) );
XNOR2_X1 U724 ( .A(KEYINPUT11), .B(n979), .ZN(n1018) );
NAND4_X1 U725 ( .A1(n1021), .A2(n1001), .A3(n1022), .A4(n1023), .ZN(n979) );
NOR4_X1 U726 ( .A1(n1024), .A2(n1025), .A3(n1011), .A4(n1026), .ZN(n1023) );
NOR3_X1 U727 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1025) );
AND2_X1 U728 ( .A1(n1030), .A2(KEYINPUT6), .ZN(n1028) );
INV_X1 U729 ( .A(n1031), .ZN(n1027) );
NOR2_X1 U730 ( .A1(n1032), .A2(n1031), .ZN(n1024) );
NAND2_X1 U731 ( .A1(KEYINPUT40), .A2(n1033), .ZN(n1031) );
INV_X1 U732 ( .A(n1030), .ZN(n1033) );
NOR2_X1 U733 ( .A1(KEYINPUT6), .A2(n1029), .ZN(n1032) );
NOR2_X1 U734 ( .A1(n1034), .A2(n1035), .ZN(n1022) );
XOR2_X1 U735 ( .A(n1036), .B(n1037), .Z(n1035) );
NOR2_X1 U736 ( .A1(KEYINPUT46), .A2(n1038), .ZN(n1037) );
XOR2_X1 U737 ( .A(n1039), .B(KEYINPUT36), .Z(n1038) );
XOR2_X1 U738 ( .A(n1040), .B(n1041), .Z(n1034) );
NOR2_X1 U739 ( .A1(G478), .A2(KEYINPUT45), .ZN(n1041) );
XNOR2_X1 U740 ( .A(n1042), .B(n1043), .ZN(n1021) );
NOR2_X1 U741 ( .A1(n1044), .A2(KEYINPUT24), .ZN(n1043) );
XOR2_X1 U742 ( .A(n1045), .B(n1046), .Z(G72) );
NOR2_X1 U743 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
AND2_X1 U744 ( .A1(G227), .A2(G900), .ZN(n1047) );
NOR2_X1 U745 ( .A1(KEYINPUT0), .A2(n1049), .ZN(n1045) );
XOR2_X1 U746 ( .A(n1050), .B(n1051), .Z(n1049) );
NOR2_X1 U747 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XOR2_X1 U748 ( .A(n1054), .B(n1055), .Z(n1053) );
XOR2_X1 U749 ( .A(n1056), .B(n1057), .Z(n1055) );
XOR2_X1 U750 ( .A(G131), .B(n1058), .Z(n1057) );
NAND2_X1 U751 ( .A1(KEYINPUT17), .A2(G134), .ZN(n1056) );
XOR2_X1 U752 ( .A(n1059), .B(n1060), .Z(n1054) );
NAND2_X1 U753 ( .A1(KEYINPUT12), .A2(n1061), .ZN(n1059) );
NOR2_X1 U754 ( .A1(G900), .A2(n1048), .ZN(n1052) );
NAND2_X1 U755 ( .A1(n1062), .A2(n1048), .ZN(n1050) );
NAND2_X1 U756 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
XOR2_X1 U757 ( .A(n978), .B(KEYINPUT35), .Z(n1063) );
XOR2_X1 U758 ( .A(n1065), .B(n1066), .Z(G69) );
NOR2_X1 U759 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U760 ( .A1(G953), .A2(n1069), .ZN(n1068) );
XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n975), .ZN(n1069) );
NOR2_X1 U762 ( .A1(n1070), .A2(n1048), .ZN(n1067) );
NOR2_X1 U763 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XNOR2_X1 U764 ( .A(G898), .B(KEYINPUT23), .ZN(n1071) );
NAND2_X1 U765 ( .A1(n1073), .A2(n1074), .ZN(n1065) );
NAND2_X1 U766 ( .A1(n1075), .A2(G953), .ZN(n1074) );
XNOR2_X1 U767 ( .A(n1076), .B(n1077), .ZN(n1073) );
XOR2_X1 U768 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(G66) );
XNOR2_X1 U770 ( .A(n1082), .B(n1083), .ZN(n1081) );
NOR2_X1 U771 ( .A1(n1030), .A2(n1084), .ZN(n1083) );
NOR2_X1 U772 ( .A1(n1080), .A2(n1085), .ZN(G63) );
XNOR2_X1 U773 ( .A(n1086), .B(n1087), .ZN(n1085) );
AND2_X1 U774 ( .A1(G478), .A2(n1088), .ZN(n1087) );
NOR2_X1 U775 ( .A1(n1080), .A2(n1089), .ZN(G60) );
NOR2_X1 U776 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U777 ( .A(KEYINPUT30), .B(n1092), .Z(n1091) );
NOR2_X1 U778 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
AND2_X1 U779 ( .A1(n1094), .A2(n1093), .ZN(n1090) );
XOR2_X1 U780 ( .A(n1095), .B(KEYINPUT13), .Z(n1093) );
NAND2_X1 U781 ( .A1(n1088), .A2(G475), .ZN(n1094) );
XNOR2_X1 U782 ( .A(G104), .B(n1096), .ZN(G6) );
NAND2_X1 U783 ( .A1(KEYINPUT15), .A2(n1097), .ZN(n1096) );
NOR2_X1 U784 ( .A1(n1080), .A2(n1098), .ZN(G57) );
XOR2_X1 U785 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U786 ( .A1(KEYINPUT32), .A2(n1101), .ZN(n1100) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(n1101) );
XNOR2_X1 U788 ( .A(n1104), .B(n1105), .ZN(n1103) );
XOR2_X1 U789 ( .A(n1106), .B(n1107), .Z(n1102) );
NOR2_X1 U790 ( .A1(n1039), .A2(n1084), .ZN(n1107) );
INV_X1 U791 ( .A(G472), .ZN(n1039) );
NAND2_X1 U792 ( .A1(KEYINPUT48), .A2(n1108), .ZN(n1106) );
NOR2_X1 U793 ( .A1(n1080), .A2(n1109), .ZN(G54) );
XOR2_X1 U794 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U795 ( .A(n1108), .B(n1112), .Z(n1111) );
XOR2_X1 U796 ( .A(n1113), .B(n1114), .Z(n1110) );
AND2_X1 U797 ( .A1(G469), .A2(n1088), .ZN(n1114) );
NAND2_X1 U798 ( .A1(KEYINPUT38), .A2(n1115), .ZN(n1113) );
NOR2_X1 U799 ( .A1(n1080), .A2(n1116), .ZN(G51) );
XOR2_X1 U800 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND3_X1 U801 ( .A1(G210), .A2(n1119), .A3(n1088), .ZN(n1118) );
INV_X1 U802 ( .A(n1084), .ZN(n1088) );
NAND2_X1 U803 ( .A1(n1120), .A2(n1121), .ZN(n1084) );
NAND3_X1 U804 ( .A1(n1122), .A2(n978), .A3(n1064), .ZN(n1121) );
INV_X1 U805 ( .A(n973), .ZN(n1064) );
NAND4_X1 U806 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n973) );
AND4_X1 U807 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1126) );
INV_X1 U808 ( .A(n975), .ZN(n1122) );
NAND4_X1 U809 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n975) );
AND4_X1 U810 ( .A1(n1135), .A2(n969), .A3(n1136), .A4(n1137), .ZN(n1134) );
NAND3_X1 U811 ( .A1(n984), .A2(n1138), .A3(n994), .ZN(n969) );
NOR2_X1 U812 ( .A1(n1097), .A2(n1139), .ZN(n1133) );
NOR4_X1 U813 ( .A1(n1013), .A2(n1140), .A3(n1141), .A4(n1004), .ZN(n1139) );
AND3_X1 U814 ( .A1(n984), .A2(n1138), .A3(n993), .ZN(n1097) );
XOR2_X1 U815 ( .A(n1142), .B(KEYINPUT22), .Z(n1120) );
NAND2_X1 U816 ( .A1(n1143), .A2(KEYINPUT62), .ZN(n1117) );
XNOR2_X1 U817 ( .A(n1144), .B(n1145), .ZN(n1143) );
XOR2_X1 U818 ( .A(n1146), .B(n1147), .Z(n1144) );
NOR2_X1 U819 ( .A1(n1048), .A2(G952), .ZN(n1080) );
XNOR2_X1 U820 ( .A(G146), .B(n978), .ZN(G48) );
NAND3_X1 U821 ( .A1(n1148), .A2(n1000), .A3(n993), .ZN(n978) );
NAND2_X1 U822 ( .A1(n1149), .A2(n1150), .ZN(G45) );
NAND2_X1 U823 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U824 ( .A(KEYINPUT59), .B(n1153), .Z(n1149) );
NOR2_X1 U825 ( .A1(n1151), .A2(n1152), .ZN(n1153) );
INV_X1 U826 ( .A(n1125), .ZN(n1151) );
NAND4_X1 U827 ( .A1(n1154), .A2(n1000), .A3(n1155), .A4(n1156), .ZN(n1125) );
XOR2_X1 U828 ( .A(n1157), .B(n1158), .Z(n1155) );
XNOR2_X1 U829 ( .A(G140), .B(n1123), .ZN(G42) );
NAND3_X1 U830 ( .A1(n1159), .A2(n1160), .A3(n991), .ZN(n1123) );
XOR2_X1 U831 ( .A(n1058), .B(n1124), .Z(G39) );
NAND3_X1 U832 ( .A1(n991), .A2(n1148), .A3(n995), .ZN(n1124) );
XNOR2_X1 U833 ( .A(G134), .B(n1130), .ZN(G36) );
NAND3_X1 U834 ( .A1(n1154), .A2(n994), .A3(n991), .ZN(n1130) );
XNOR2_X1 U835 ( .A(G131), .B(n1129), .ZN(G33) );
NAND3_X1 U836 ( .A1(n1154), .A2(n993), .A3(n991), .ZN(n1129) );
NOR2_X1 U837 ( .A1(n1002), .A2(n1161), .ZN(n991) );
INV_X1 U838 ( .A(n1001), .ZN(n1161) );
AND3_X1 U839 ( .A1(n1160), .A2(n1162), .A3(n1016), .ZN(n1154) );
XNOR2_X1 U840 ( .A(G128), .B(n1128), .ZN(G30) );
NAND3_X1 U841 ( .A1(n994), .A2(n1000), .A3(n1148), .ZN(n1128) );
AND4_X1 U842 ( .A1(n1160), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1148) );
NAND2_X1 U843 ( .A1(KEYINPUT29), .A2(n1141), .ZN(n1164) );
NAND2_X1 U844 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
INV_X1 U845 ( .A(KEYINPUT29), .ZN(n1166) );
NAND2_X1 U846 ( .A1(n1167), .A2(n1010), .ZN(n1165) );
XNOR2_X1 U847 ( .A(G101), .B(n1168), .ZN(G3) );
NAND4_X1 U848 ( .A1(n1169), .A2(n995), .A3(n1016), .A4(n1170), .ZN(n1168) );
INV_X1 U849 ( .A(n1140), .ZN(n1170) );
XOR2_X1 U850 ( .A(n1013), .B(KEYINPUT53), .Z(n1169) );
XOR2_X1 U851 ( .A(n1127), .B(n1171), .Z(G27) );
NAND2_X1 U852 ( .A1(KEYINPUT28), .A2(G125), .ZN(n1171) );
NAND3_X1 U853 ( .A1(n985), .A2(n1000), .A3(n1159), .ZN(n1127) );
AND4_X1 U854 ( .A1(n993), .A2(n986), .A3(n1010), .A4(n1162), .ZN(n1159) );
NAND2_X1 U855 ( .A1(n1017), .A2(n1172), .ZN(n1162) );
NAND4_X1 U856 ( .A1(G953), .A2(G902), .A3(n1173), .A4(n1174), .ZN(n1172) );
INV_X1 U857 ( .A(G900), .ZN(n1174) );
INV_X1 U858 ( .A(n1011), .ZN(n985) );
XNOR2_X1 U859 ( .A(n1175), .B(n1135), .ZN(G24) );
NAND4_X1 U860 ( .A1(n1176), .A2(n1177), .A3(n984), .A4(n986), .ZN(n1135) );
INV_X1 U861 ( .A(n1167), .ZN(n986) );
NOR2_X1 U862 ( .A1(n1178), .A2(n1179), .ZN(n1176) );
NOR2_X1 U863 ( .A1(n1180), .A2(n1157), .ZN(n1179) );
INV_X1 U864 ( .A(KEYINPUT8), .ZN(n1157) );
NOR2_X1 U865 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NOR2_X1 U866 ( .A1(KEYINPUT8), .A2(n994), .ZN(n1178) );
NAND2_X1 U867 ( .A1(KEYINPUT41), .A2(n1183), .ZN(n1175) );
INV_X1 U868 ( .A(G122), .ZN(n1183) );
XOR2_X1 U869 ( .A(n1184), .B(n1131), .Z(G21) );
NAND4_X1 U870 ( .A1(n1177), .A2(n995), .A3(n1167), .A4(n1185), .ZN(n1131) );
XOR2_X1 U871 ( .A(KEYINPUT29), .B(n1010), .Z(n1185) );
XOR2_X1 U872 ( .A(n1186), .B(n1132), .Z(G18) );
NAND3_X1 U873 ( .A1(n1016), .A2(n994), .A3(n1177), .ZN(n1132) );
NOR2_X1 U874 ( .A1(n1181), .A2(n1158), .ZN(n994) );
XOR2_X1 U875 ( .A(n1137), .B(n1187), .Z(G15) );
XOR2_X1 U876 ( .A(KEYINPUT10), .B(G113), .Z(n1187) );
NAND3_X1 U877 ( .A1(n1016), .A2(n993), .A3(n1177), .ZN(n1137) );
NOR2_X1 U878 ( .A1(n1011), .A2(n1140), .ZN(n1177) );
NAND2_X1 U879 ( .A1(n1015), .A2(n1188), .ZN(n1011) );
NOR2_X1 U880 ( .A1(n1182), .A2(n1156), .ZN(n993) );
INV_X1 U881 ( .A(n1181), .ZN(n1156) );
INV_X1 U882 ( .A(n1141), .ZN(n1016) );
NAND2_X1 U883 ( .A1(n1167), .A2(n984), .ZN(n1141) );
INV_X1 U884 ( .A(n1010), .ZN(n984) );
XNOR2_X1 U885 ( .A(G110), .B(n1136), .ZN(G12) );
NAND3_X1 U886 ( .A1(n1138), .A2(n1010), .A3(n995), .ZN(n1136) );
INV_X1 U887 ( .A(n1004), .ZN(n995) );
NAND2_X1 U888 ( .A1(n1181), .A2(n1182), .ZN(n1004) );
INV_X1 U889 ( .A(n1158), .ZN(n1182) );
XNOR2_X1 U890 ( .A(n1026), .B(KEYINPUT61), .ZN(n1158) );
XNOR2_X1 U891 ( .A(n1189), .B(G475), .ZN(n1026) );
NAND2_X1 U892 ( .A1(n1095), .A2(n1142), .ZN(n1189) );
XNOR2_X1 U893 ( .A(n1190), .B(n1191), .ZN(n1095) );
XOR2_X1 U894 ( .A(n1061), .B(n1192), .Z(n1191) );
XOR2_X1 U895 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U896 ( .A1(KEYINPUT56), .A2(n1195), .ZN(n1194) );
XOR2_X1 U897 ( .A(KEYINPUT5), .B(G146), .Z(n1195) );
NAND2_X1 U898 ( .A1(G214), .A2(n1196), .ZN(n1193) );
XNOR2_X1 U899 ( .A(G140), .B(G125), .ZN(n1061) );
XOR2_X1 U900 ( .A(n1197), .B(n1198), .Z(n1190) );
NOR2_X1 U901 ( .A1(KEYINPUT26), .A2(n1199), .ZN(n1198) );
XOR2_X1 U902 ( .A(n1200), .B(n1201), .Z(n1199) );
XNOR2_X1 U903 ( .A(G104), .B(n1202), .ZN(n1201) );
NOR2_X1 U904 ( .A1(G122), .A2(KEYINPUT20), .ZN(n1202) );
XOR2_X1 U905 ( .A(n1203), .B(KEYINPUT25), .Z(n1200) );
XOR2_X1 U906 ( .A(G131), .B(n1152), .Z(n1197) );
XOR2_X1 U907 ( .A(n1040), .B(G478), .Z(n1181) );
NAND2_X1 U908 ( .A1(n1086), .A2(n1142), .ZN(n1040) );
XNOR2_X1 U909 ( .A(n1204), .B(n1205), .ZN(n1086) );
XOR2_X1 U910 ( .A(G116), .B(n1206), .Z(n1205) );
XOR2_X1 U911 ( .A(G134), .B(G122), .Z(n1206) );
XOR2_X1 U912 ( .A(n1207), .B(n1208), .Z(n1204) );
XNOR2_X1 U913 ( .A(G107), .B(n1209), .ZN(n1208) );
NAND3_X1 U914 ( .A1(G217), .A2(n1048), .A3(G234), .ZN(n1209) );
NAND2_X1 U915 ( .A1(KEYINPUT47), .A2(n1210), .ZN(n1207) );
XOR2_X1 U916 ( .A(G143), .B(G128), .Z(n1210) );
XNOR2_X1 U917 ( .A(n1030), .B(n1211), .ZN(n1010) );
NOR2_X1 U918 ( .A1(KEYINPUT18), .A2(n1029), .ZN(n1211) );
NAND2_X1 U919 ( .A1(n1082), .A2(n1142), .ZN(n1029) );
XNOR2_X1 U920 ( .A(n1212), .B(n1213), .ZN(n1082) );
XOR2_X1 U921 ( .A(n1214), .B(n1215), .Z(n1213) );
XOR2_X1 U922 ( .A(G125), .B(G119), .Z(n1215) );
XOR2_X1 U923 ( .A(KEYINPUT5), .B(G137), .Z(n1214) );
XOR2_X1 U924 ( .A(n1216), .B(n1217), .Z(n1212) );
XOR2_X1 U925 ( .A(n1218), .B(n1219), .Z(n1216) );
NAND3_X1 U926 ( .A1(G234), .A2(n1048), .A3(G221), .ZN(n1218) );
NAND2_X1 U927 ( .A1(G217), .A2(n1220), .ZN(n1030) );
NOR3_X1 U928 ( .A1(n1013), .A2(n1167), .A3(n1140), .ZN(n1138) );
NAND2_X1 U929 ( .A1(n1000), .A2(n1221), .ZN(n1140) );
NAND2_X1 U930 ( .A1(n1017), .A2(n1222), .ZN(n1221) );
NAND4_X1 U931 ( .A1(n1075), .A2(G953), .A3(G902), .A4(n1173), .ZN(n1222) );
XNOR2_X1 U932 ( .A(G898), .B(KEYINPUT16), .ZN(n1075) );
NAND3_X1 U933 ( .A1(n976), .A2(n1173), .A3(n1223), .ZN(n1017) );
XOR2_X1 U934 ( .A(n974), .B(KEYINPUT51), .Z(n1223) );
INV_X1 U935 ( .A(G952), .ZN(n974) );
NAND2_X1 U936 ( .A1(G237), .A2(G234), .ZN(n1173) );
INV_X1 U937 ( .A(n1019), .ZN(n976) );
XOR2_X1 U938 ( .A(n1048), .B(KEYINPUT55), .Z(n1019) );
AND2_X1 U939 ( .A1(n1002), .A2(n1001), .ZN(n1000) );
NAND2_X1 U940 ( .A1(G214), .A2(n1119), .ZN(n1001) );
XNOR2_X1 U941 ( .A(n1042), .B(n1044), .ZN(n1002) );
AND2_X1 U942 ( .A1(n1224), .A2(n1119), .ZN(n1044) );
OR2_X1 U943 ( .A1(G902), .A2(G237), .ZN(n1119) );
XNOR2_X1 U944 ( .A(G210), .B(KEYINPUT9), .ZN(n1224) );
NAND2_X1 U945 ( .A1(n1225), .A2(n1142), .ZN(n1042) );
XOR2_X1 U946 ( .A(n1226), .B(n1227), .Z(n1225) );
INV_X1 U947 ( .A(n1146), .ZN(n1227) );
XOR2_X1 U948 ( .A(n1228), .B(n1078), .Z(n1146) );
XNOR2_X1 U949 ( .A(n1229), .B(G110), .ZN(n1078) );
NAND2_X1 U950 ( .A1(KEYINPUT3), .A2(G122), .ZN(n1229) );
XOR2_X1 U951 ( .A(n1230), .B(KEYINPUT4), .Z(n1228) );
NAND3_X1 U952 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1230) );
NAND2_X1 U953 ( .A1(KEYINPUT52), .A2(n1079), .ZN(n1233) );
NAND3_X1 U954 ( .A1(n1234), .A2(n1235), .A3(n1076), .ZN(n1232) );
INV_X1 U955 ( .A(KEYINPUT52), .ZN(n1235) );
OR2_X1 U956 ( .A1(n1076), .A2(n1234), .ZN(n1231) );
NOR2_X1 U957 ( .A1(KEYINPUT60), .A2(n1079), .ZN(n1234) );
XNOR2_X1 U958 ( .A(n1236), .B(n1237), .ZN(n1079) );
NAND2_X1 U959 ( .A1(KEYINPUT43), .A2(n1238), .ZN(n1236) );
XOR2_X1 U960 ( .A(n1239), .B(n1240), .Z(n1076) );
XOR2_X1 U961 ( .A(n1186), .B(n1241), .Z(n1240) );
NAND2_X1 U962 ( .A1(n1242), .A2(KEYINPUT2), .ZN(n1241) );
XOR2_X1 U963 ( .A(n1203), .B(KEYINPUT63), .Z(n1242) );
INV_X1 U964 ( .A(G113), .ZN(n1203) );
NAND2_X1 U965 ( .A1(KEYINPUT7), .A2(n1184), .ZN(n1239) );
XNOR2_X1 U966 ( .A(KEYINPUT1), .B(n1243), .ZN(n1226) );
NOR2_X1 U967 ( .A1(KEYINPUT31), .A2(n1244), .ZN(n1243) );
XNOR2_X1 U968 ( .A(n1147), .B(n1245), .ZN(n1244) );
NOR2_X1 U969 ( .A1(KEYINPUT39), .A2(n1145), .ZN(n1245) );
XNOR2_X1 U970 ( .A(G125), .B(n1105), .ZN(n1145) );
NOR2_X1 U971 ( .A1(n1072), .A2(G953), .ZN(n1147) );
INV_X1 U972 ( .A(G224), .ZN(n1072) );
XOR2_X1 U973 ( .A(n1246), .B(G472), .Z(n1167) );
NAND2_X1 U974 ( .A1(KEYINPUT42), .A2(n1036), .ZN(n1246) );
NAND2_X1 U975 ( .A1(n1247), .A2(n1142), .ZN(n1036) );
XOR2_X1 U976 ( .A(n1099), .B(n1248), .Z(n1247) );
XOR2_X1 U977 ( .A(n1249), .B(n1250), .Z(n1248) );
NAND2_X1 U978 ( .A1(KEYINPUT58), .A2(n1104), .ZN(n1250) );
XNOR2_X1 U979 ( .A(n1251), .B(n1252), .ZN(n1104) );
XOR2_X1 U980 ( .A(G113), .B(n1253), .Z(n1252) );
NOR2_X1 U981 ( .A1(KEYINPUT54), .A2(n1184), .ZN(n1253) );
INV_X1 U982 ( .A(G119), .ZN(n1184) );
XOR2_X1 U983 ( .A(n1186), .B(KEYINPUT14), .Z(n1251) );
INV_X1 U984 ( .A(G116), .ZN(n1186) );
NAND2_X1 U985 ( .A1(n1254), .A2(n1255), .ZN(n1249) );
OR2_X1 U986 ( .A1(n1108), .A2(n1105), .ZN(n1255) );
XOR2_X1 U987 ( .A(n1256), .B(KEYINPUT50), .Z(n1254) );
NAND2_X1 U988 ( .A1(n1108), .A2(n1105), .ZN(n1256) );
XOR2_X1 U989 ( .A(G128), .B(n1257), .Z(n1105) );
NOR2_X1 U990 ( .A1(KEYINPUT57), .A2(n1258), .ZN(n1257) );
XOR2_X1 U991 ( .A(G146), .B(G143), .Z(n1258) );
XOR2_X1 U992 ( .A(n1259), .B(n1238), .Z(n1099) );
NAND2_X1 U993 ( .A1(G210), .A2(n1196), .ZN(n1259) );
NOR2_X1 U994 ( .A1(G953), .A2(G237), .ZN(n1196) );
INV_X1 U995 ( .A(n1160), .ZN(n1013) );
NOR2_X1 U996 ( .A1(n1015), .A2(n1014), .ZN(n1160) );
INV_X1 U997 ( .A(n1188), .ZN(n1014) );
NAND2_X1 U998 ( .A1(G221), .A2(n1220), .ZN(n1188) );
NAND2_X1 U999 ( .A1(G234), .A2(n1142), .ZN(n1220) );
INV_X1 U1000 ( .A(G902), .ZN(n1142) );
XNOR2_X1 U1001 ( .A(G469), .B(n1260), .ZN(n1015) );
NOR2_X1 U1002 ( .A1(G902), .A2(n1261), .ZN(n1260) );
XNOR2_X1 U1003 ( .A(n1112), .B(n1262), .ZN(n1261) );
NOR2_X1 U1004 ( .A1(KEYINPUT34), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U1005 ( .A(n1108), .B(n1115), .ZN(n1263) );
XOR2_X1 U1006 ( .A(n1060), .B(n1264), .Z(n1115) );
XOR2_X1 U1007 ( .A(n1238), .B(n1237), .Z(n1264) );
XOR2_X1 U1008 ( .A(G104), .B(G107), .Z(n1237) );
XOR2_X1 U1009 ( .A(G101), .B(KEYINPUT49), .Z(n1238) );
XNOR2_X1 U1010 ( .A(n1152), .B(n1219), .ZN(n1060) );
XOR2_X1 U1011 ( .A(G128), .B(G146), .Z(n1219) );
INV_X1 U1012 ( .A(G143), .ZN(n1152) );
NAND2_X1 U1013 ( .A1(n1265), .A2(n1266), .ZN(n1108) );
NAND2_X1 U1014 ( .A1(n1267), .A2(G137), .ZN(n1266) );
NAND2_X1 U1015 ( .A1(n1268), .A2(n1058), .ZN(n1265) );
INV_X1 U1016 ( .A(G137), .ZN(n1058) );
XOR2_X1 U1017 ( .A(n1269), .B(n1267), .Z(n1268) );
XOR2_X1 U1018 ( .A(G131), .B(G134), .Z(n1267) );
XNOR2_X1 U1019 ( .A(KEYINPUT33), .B(KEYINPUT27), .ZN(n1269) );
XNOR2_X1 U1020 ( .A(n1270), .B(n1217), .ZN(n1112) );
XOR2_X1 U1021 ( .A(G110), .B(G140), .Z(n1217) );
NAND2_X1 U1022 ( .A1(G227), .A2(n1048), .ZN(n1270) );
INV_X1 U1023 ( .A(G953), .ZN(n1048) );
endmodule


