//Key = 1010001001000110011011001101001010101010110110110101100100101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374;

XNOR2_X1 U750 ( .A(G107), .B(n1044), .ZN(G9) );
NOR2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(G75) );
NOR4_X1 U752 ( .A1(G953), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1046) );
INV_X1 U753 ( .A(n1050), .ZN(n1049) );
NOR2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1048) );
NOR2_X1 U755 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR3_X1 U756 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NOR2_X1 U757 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U758 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR3_X1 U759 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1058) );
NOR3_X1 U760 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NOR2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U762 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U763 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
XOR2_X1 U764 ( .A(n1074), .B(KEYINPUT57), .Z(n1072) );
NOR2_X1 U765 ( .A1(n1075), .A2(n1076), .ZN(n1066) );
NOR2_X1 U766 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NOR2_X1 U767 ( .A1(n1079), .A2(n1080), .ZN(n1063) );
NOR4_X1 U768 ( .A1(n1065), .A2(n1081), .A3(n1062), .A4(n1061), .ZN(n1053) );
NOR2_X1 U769 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR3_X1 U770 ( .A1(n1047), .A2(G953), .A3(G952), .ZN(n1045) );
AND4_X1 U771 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1047) );
NOR4_X1 U772 ( .A1(n1065), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1087) );
XNOR2_X1 U773 ( .A(n1091), .B(n1092), .ZN(n1090) );
NOR2_X1 U774 ( .A1(KEYINPUT56), .A2(n1093), .ZN(n1092) );
XNOR2_X1 U775 ( .A(KEYINPUT39), .B(n1094), .ZN(n1093) );
XOR2_X1 U776 ( .A(n1095), .B(n1096), .Z(n1089) );
NOR2_X1 U777 ( .A1(KEYINPUT45), .A2(n1097), .ZN(n1096) );
INV_X1 U778 ( .A(n1073), .ZN(n1088) );
NOR2_X1 U779 ( .A1(n1098), .A2(n1099), .ZN(n1086) );
XNOR2_X1 U780 ( .A(G472), .B(n1100), .ZN(n1099) );
XOR2_X1 U781 ( .A(KEYINPUT4), .B(n1101), .Z(n1098) );
XOR2_X1 U782 ( .A(KEYINPUT40), .B(n1102), .Z(n1085) );
XOR2_X1 U783 ( .A(KEYINPUT25), .B(n1103), .Z(n1084) );
XOR2_X1 U784 ( .A(n1104), .B(n1105), .Z(G72) );
NOR2_X1 U785 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
AND3_X1 U786 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1107) );
NOR3_X1 U787 ( .A1(n1108), .A2(n1111), .A3(n1112), .ZN(n1106) );
XOR2_X1 U788 ( .A(n1113), .B(KEYINPUT18), .Z(n1112) );
NAND2_X1 U789 ( .A1(n1109), .A2(n1110), .ZN(n1113) );
NOR2_X1 U790 ( .A1(G900), .A2(n1109), .ZN(n1111) );
XNOR2_X1 U791 ( .A(n1114), .B(n1115), .ZN(n1108) );
XOR2_X1 U792 ( .A(G137), .B(G134), .Z(n1115) );
XOR2_X1 U793 ( .A(n1116), .B(G131), .Z(n1114) );
NAND3_X1 U794 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1116) );
NAND2_X1 U795 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND3_X1 U796 ( .A1(G125), .A2(n1122), .A3(G140), .ZN(n1118) );
NAND2_X1 U797 ( .A1(n1123), .A2(n1124), .ZN(n1117) );
XOR2_X1 U798 ( .A(G125), .B(n1122), .Z(n1123) );
NAND3_X1 U799 ( .A1(n1125), .A2(n1126), .A3(KEYINPUT32), .ZN(n1104) );
NAND2_X1 U800 ( .A1(G900), .A2(G227), .ZN(n1126) );
INV_X1 U801 ( .A(n1127), .ZN(n1125) );
XOR2_X1 U802 ( .A(n1128), .B(n1129), .Z(G69) );
NOR2_X1 U803 ( .A1(n1130), .A2(n1127), .ZN(n1129) );
XOR2_X1 U804 ( .A(n1109), .B(KEYINPUT26), .Z(n1127) );
AND2_X1 U805 ( .A1(G224), .A2(G898), .ZN(n1130) );
NAND2_X1 U806 ( .A1(n1131), .A2(n1132), .ZN(n1128) );
NAND2_X1 U807 ( .A1(n1133), .A2(n1109), .ZN(n1132) );
XOR2_X1 U808 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND3_X1 U809 ( .A1(G898), .A2(n1134), .A3(G953), .ZN(n1131) );
XNOR2_X1 U810 ( .A(n1136), .B(n1137), .ZN(n1134) );
XOR2_X1 U811 ( .A(n1138), .B(n1139), .Z(n1136) );
NOR2_X1 U812 ( .A1(n1140), .A2(n1141), .ZN(G66) );
XOR2_X1 U813 ( .A(KEYINPUT28), .B(n1142), .Z(n1141) );
NOR3_X1 U814 ( .A1(n1091), .A2(n1143), .A3(n1144), .ZN(n1140) );
AND3_X1 U815 ( .A1(n1145), .A2(G217), .A3(n1146), .ZN(n1144) );
NOR2_X1 U816 ( .A1(n1147), .A2(n1145), .ZN(n1143) );
NOR2_X1 U817 ( .A1(n1050), .A2(n1148), .ZN(n1147) );
NOR2_X1 U818 ( .A1(n1142), .A2(n1149), .ZN(G63) );
NOR3_X1 U819 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1149) );
NOR2_X1 U820 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U821 ( .A1(n1155), .A2(n1156), .ZN(n1153) );
XNOR2_X1 U822 ( .A(KEYINPUT49), .B(n1157), .ZN(n1156) );
NOR3_X1 U823 ( .A1(n1158), .A2(n1157), .A3(n1155), .ZN(n1151) );
AND2_X1 U824 ( .A1(n1155), .A2(n1157), .ZN(n1150) );
NAND2_X1 U825 ( .A1(n1146), .A2(G478), .ZN(n1157) );
INV_X1 U826 ( .A(KEYINPUT24), .ZN(n1155) );
NOR2_X1 U827 ( .A1(n1142), .A2(n1159), .ZN(G60) );
XOR2_X1 U828 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U829 ( .A(n1162), .B(KEYINPUT23), .Z(n1161) );
NAND2_X1 U830 ( .A1(n1146), .A2(G475), .ZN(n1162) );
XOR2_X1 U831 ( .A(n1163), .B(n1164), .Z(G6) );
NOR2_X1 U832 ( .A1(n1142), .A2(n1165), .ZN(G57) );
XOR2_X1 U833 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U834 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U835 ( .A(n1170), .B(n1171), .Z(n1168) );
NAND2_X1 U836 ( .A1(n1146), .A2(G472), .ZN(n1170) );
XOR2_X1 U837 ( .A(n1172), .B(n1173), .Z(n1166) );
NOR2_X1 U838 ( .A1(KEYINPUT22), .A2(n1174), .ZN(n1173) );
XOR2_X1 U839 ( .A(n1175), .B(KEYINPUT60), .Z(n1172) );
NOR2_X1 U840 ( .A1(n1142), .A2(n1176), .ZN(G54) );
XOR2_X1 U841 ( .A(n1177), .B(n1178), .Z(n1176) );
NOR3_X1 U842 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1178) );
INV_X1 U843 ( .A(G469), .ZN(n1180) );
XOR2_X1 U844 ( .A(KEYINPUT3), .B(n1050), .Z(n1179) );
NOR2_X1 U845 ( .A1(n1182), .A2(n1183), .ZN(n1177) );
XOR2_X1 U846 ( .A(n1184), .B(KEYINPUT27), .Z(n1183) );
NAND2_X1 U847 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NOR2_X1 U848 ( .A1(n1185), .A2(n1186), .ZN(n1182) );
XOR2_X1 U849 ( .A(n1187), .B(n1188), .Z(n1185) );
NAND2_X1 U850 ( .A1(KEYINPUT34), .A2(n1189), .ZN(n1187) );
NOR3_X1 U851 ( .A1(n1142), .A2(n1190), .A3(n1191), .ZN(G51) );
NOR2_X1 U852 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U853 ( .A(n1194), .B(n1195), .Z(n1193) );
AND2_X1 U854 ( .A1(n1196), .A2(KEYINPUT0), .ZN(n1195) );
NOR2_X1 U855 ( .A1(n1197), .A2(n1198), .ZN(n1190) );
XOR2_X1 U856 ( .A(n1194), .B(n1199), .Z(n1198) );
NOR2_X1 U857 ( .A1(n1200), .A2(n1196), .ZN(n1199) );
XNOR2_X1 U858 ( .A(n1201), .B(n1202), .ZN(n1196) );
NOR2_X1 U859 ( .A1(G125), .A2(KEYINPUT31), .ZN(n1202) );
INV_X1 U860 ( .A(KEYINPUT0), .ZN(n1200) );
XOR2_X1 U861 ( .A(n1203), .B(n1204), .Z(n1194) );
NAND2_X1 U862 ( .A1(n1146), .A2(n1205), .ZN(n1203) );
NOR2_X1 U863 ( .A1(n1181), .A2(n1050), .ZN(n1146) );
NOR2_X1 U864 ( .A1(n1135), .A2(n1110), .ZN(n1050) );
NAND4_X1 U865 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1110) );
AND4_X1 U866 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1209) );
OR2_X1 U867 ( .A1(n1214), .A2(KEYINPUT42), .ZN(n1208) );
NAND2_X1 U868 ( .A1(n1215), .A2(n1216), .ZN(n1207) );
NAND2_X1 U869 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NAND3_X1 U870 ( .A1(n1219), .A2(n1220), .A3(KEYINPUT42), .ZN(n1218) );
INV_X1 U871 ( .A(n1083), .ZN(n1220) );
NAND2_X1 U872 ( .A1(n1071), .A2(n1221), .ZN(n1206) );
NAND2_X1 U873 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
XOR2_X1 U874 ( .A(n1224), .B(KEYINPUT54), .Z(n1223) );
XOR2_X1 U875 ( .A(n1225), .B(KEYINPUT37), .Z(n1222) );
NAND4_X1 U876 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1135) );
AND4_X1 U877 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1044), .ZN(n1229) );
NAND3_X1 U878 ( .A1(n1077), .A2(n1233), .A3(n1234), .ZN(n1044) );
NOR3_X1 U879 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1228) );
AND4_X1 U880 ( .A1(KEYINPUT19), .A2(n1078), .A3(n1060), .A4(n1233), .ZN(n1237) );
NOR2_X1 U881 ( .A1(KEYINPUT19), .A2(n1164), .ZN(n1236) );
NAND3_X1 U882 ( .A1(n1234), .A2(n1233), .A3(n1078), .ZN(n1164) );
NOR4_X1 U883 ( .A1(n1238), .A2(n1055), .A3(n1057), .A4(n1239), .ZN(n1233) );
NOR2_X1 U884 ( .A1(n1240), .A2(n1238), .ZN(n1235) );
XOR2_X1 U885 ( .A(n1241), .B(KEYINPUT50), .Z(n1240) );
INV_X1 U886 ( .A(n1192), .ZN(n1197) );
NOR2_X1 U887 ( .A1(n1109), .A2(G952), .ZN(n1142) );
XOR2_X1 U888 ( .A(n1242), .B(n1212), .Z(G48) );
NAND3_X1 U889 ( .A1(n1078), .A2(n1071), .A3(n1243), .ZN(n1212) );
INV_X1 U890 ( .A(n1238), .ZN(n1071) );
XOR2_X1 U891 ( .A(G143), .B(n1244), .Z(G45) );
NOR2_X1 U892 ( .A1(n1238), .A2(n1225), .ZN(n1244) );
NAND4_X1 U893 ( .A1(n1245), .A2(n1082), .A3(n1102), .A4(n1101), .ZN(n1225) );
XOR2_X1 U894 ( .A(n1124), .B(n1214), .Z(G42) );
NAND3_X1 U895 ( .A1(n1215), .A2(n1083), .A3(n1219), .ZN(n1214) );
XOR2_X1 U896 ( .A(n1211), .B(n1246), .Z(G39) );
XOR2_X1 U897 ( .A(n1247), .B(KEYINPUT35), .Z(n1246) );
NAND2_X1 U898 ( .A1(n1243), .A2(n1079), .ZN(n1211) );
INV_X1 U899 ( .A(n1061), .ZN(n1079) );
NAND2_X1 U900 ( .A1(n1215), .A2(n1248), .ZN(n1061) );
XOR2_X1 U901 ( .A(n1249), .B(n1210), .Z(G36) );
NAND4_X1 U902 ( .A1(n1245), .A2(n1215), .A3(n1082), .A4(n1077), .ZN(n1210) );
INV_X1 U903 ( .A(n1076), .ZN(n1215) );
XOR2_X1 U904 ( .A(G131), .B(n1250), .Z(G33) );
NOR2_X1 U905 ( .A1(n1251), .A2(n1076), .ZN(n1250) );
NAND2_X1 U906 ( .A1(n1252), .A2(n1073), .ZN(n1076) );
INV_X1 U907 ( .A(n1074), .ZN(n1252) );
XOR2_X1 U908 ( .A(n1253), .B(KEYINPUT20), .Z(n1074) );
XOR2_X1 U909 ( .A(n1217), .B(KEYINPUT5), .Z(n1251) );
NAND2_X1 U910 ( .A1(n1219), .A2(n1082), .ZN(n1217) );
AND2_X1 U911 ( .A1(n1245), .A2(n1078), .ZN(n1219) );
XOR2_X1 U912 ( .A(G128), .B(n1254), .Z(G30) );
NOR2_X1 U913 ( .A1(n1238), .A2(n1224), .ZN(n1254) );
NAND2_X1 U914 ( .A1(n1243), .A2(n1077), .ZN(n1224) );
AND3_X1 U915 ( .A1(n1055), .A2(n1057), .A3(n1245), .ZN(n1243) );
AND2_X1 U916 ( .A1(n1234), .A2(n1255), .ZN(n1245) );
XNOR2_X1 U917 ( .A(G101), .B(n1232), .ZN(G3) );
NAND4_X1 U918 ( .A1(n1248), .A2(n1082), .A3(n1256), .A4(n1234), .ZN(n1232) );
NOR2_X1 U919 ( .A1(n1239), .A2(n1238), .ZN(n1256) );
INV_X1 U920 ( .A(n1257), .ZN(n1239) );
XOR2_X1 U921 ( .A(n1258), .B(n1213), .Z(G27) );
NAND4_X1 U922 ( .A1(n1083), .A2(n1078), .A3(n1259), .A4(n1255), .ZN(n1213) );
NAND2_X1 U923 ( .A1(n1052), .A2(n1260), .ZN(n1255) );
NAND4_X1 U924 ( .A1(G902), .A2(G953), .A3(n1261), .A4(n1262), .ZN(n1260) );
INV_X1 U925 ( .A(G900), .ZN(n1262) );
XNOR2_X1 U926 ( .A(G122), .B(n1231), .ZN(G24) );
NAND3_X1 U927 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1231) );
NOR3_X1 U928 ( .A1(n1057), .A2(n1266), .A3(n1267), .ZN(n1265) );
XNOR2_X1 U929 ( .A(G119), .B(n1226), .ZN(G21) );
NAND4_X1 U930 ( .A1(n1055), .A2(n1248), .A3(n1057), .A4(n1263), .ZN(n1226) );
NAND2_X1 U931 ( .A1(n1268), .A2(n1269), .ZN(G18) );
NAND2_X1 U932 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XOR2_X1 U933 ( .A(n1227), .B(KEYINPUT38), .Z(n1270) );
NAND2_X1 U934 ( .A1(n1272), .A2(G116), .ZN(n1268) );
XNOR2_X1 U935 ( .A(KEYINPUT13), .B(n1227), .ZN(n1272) );
NAND3_X1 U936 ( .A1(n1263), .A2(n1077), .A3(n1082), .ZN(n1227) );
NOR2_X1 U937 ( .A1(n1101), .A2(n1267), .ZN(n1077) );
INV_X1 U938 ( .A(n1266), .ZN(n1101) );
XOR2_X1 U939 ( .A(n1273), .B(n1230), .Z(G15) );
NAND3_X1 U940 ( .A1(n1078), .A2(n1263), .A3(n1082), .ZN(n1230) );
AND2_X1 U941 ( .A1(n1057), .A2(n1264), .ZN(n1082) );
AND2_X1 U942 ( .A1(n1259), .A2(n1257), .ZN(n1263) );
NOR3_X1 U943 ( .A1(n1062), .A2(n1065), .A3(n1238), .ZN(n1259) );
INV_X1 U944 ( .A(n1080), .ZN(n1065) );
NOR2_X1 U945 ( .A1(n1102), .A2(n1266), .ZN(n1078) );
INV_X1 U946 ( .A(n1267), .ZN(n1102) );
XOR2_X1 U947 ( .A(G110), .B(n1274), .Z(G12) );
NOR2_X1 U948 ( .A1(n1238), .A2(n1241), .ZN(n1274) );
NAND4_X1 U949 ( .A1(n1083), .A2(n1248), .A3(n1234), .A4(n1257), .ZN(n1241) );
NAND2_X1 U950 ( .A1(n1052), .A2(n1275), .ZN(n1257) );
NAND4_X1 U951 ( .A1(G902), .A2(G953), .A3(n1261), .A4(n1276), .ZN(n1275) );
INV_X1 U952 ( .A(G898), .ZN(n1276) );
NAND3_X1 U953 ( .A1(n1261), .A2(n1109), .A3(G952), .ZN(n1052) );
INV_X1 U954 ( .A(G953), .ZN(n1109) );
NAND2_X1 U955 ( .A1(G237), .A2(G234), .ZN(n1261) );
INV_X1 U956 ( .A(n1060), .ZN(n1234) );
NAND2_X1 U957 ( .A1(n1062), .A2(n1080), .ZN(n1060) );
NAND2_X1 U958 ( .A1(n1277), .A2(n1278), .ZN(n1080) );
NAND2_X1 U959 ( .A1(G234), .A2(n1181), .ZN(n1278) );
XOR2_X1 U960 ( .A(KEYINPUT1), .B(G221), .Z(n1277) );
XNOR2_X1 U961 ( .A(n1095), .B(n1097), .ZN(n1062) );
XNOR2_X1 U962 ( .A(G469), .B(KEYINPUT44), .ZN(n1097) );
NAND2_X1 U963 ( .A1(n1279), .A2(n1181), .ZN(n1095) );
XNOR2_X1 U964 ( .A(n1186), .B(n1280), .ZN(n1279) );
XOR2_X1 U965 ( .A(n1281), .B(n1188), .Z(n1280) );
XOR2_X1 U966 ( .A(G110), .B(G140), .Z(n1188) );
NOR2_X1 U967 ( .A1(KEYINPUT16), .A2(n1189), .ZN(n1281) );
NAND2_X1 U968 ( .A1(G227), .A2(n1282), .ZN(n1189) );
XNOR2_X1 U969 ( .A(n1169), .B(n1283), .ZN(n1186) );
XOR2_X1 U970 ( .A(n1284), .B(n1122), .Z(n1283) );
INV_X1 U971 ( .A(n1121), .ZN(n1122) );
XOR2_X1 U972 ( .A(n1285), .B(KEYINPUT51), .Z(n1121) );
NOR2_X1 U973 ( .A1(KEYINPUT10), .A2(n1286), .ZN(n1284) );
NOR2_X1 U974 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XOR2_X1 U975 ( .A(KEYINPUT29), .B(n1289), .Z(n1288) );
AND2_X1 U976 ( .A1(n1163), .A2(G107), .ZN(n1289) );
NOR2_X1 U977 ( .A1(G107), .A2(n1163), .ZN(n1287) );
XOR2_X1 U978 ( .A(n1290), .B(n1291), .Z(n1169) );
INV_X1 U979 ( .A(n1069), .ZN(n1248) );
NAND2_X1 U980 ( .A1(n1267), .A2(n1266), .ZN(n1069) );
XOR2_X1 U981 ( .A(n1292), .B(G475), .Z(n1266) );
NAND2_X1 U982 ( .A1(n1160), .A2(n1181), .ZN(n1292) );
XOR2_X1 U983 ( .A(n1293), .B(n1294), .Z(n1160) );
NOR3_X1 U984 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1294) );
NOR2_X1 U985 ( .A1(G113), .A2(n1298), .ZN(n1297) );
NOR2_X1 U986 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XNOR2_X1 U987 ( .A(G122), .B(KEYINPUT14), .ZN(n1299) );
NOR3_X1 U988 ( .A1(n1273), .A2(G122), .A3(n1300), .ZN(n1296) );
INV_X1 U989 ( .A(G113), .ZN(n1273) );
AND2_X1 U990 ( .A1(n1300), .A2(G122), .ZN(n1295) );
INV_X1 U991 ( .A(KEYINPUT9), .ZN(n1300) );
XOR2_X1 U992 ( .A(n1301), .B(G104), .Z(n1293) );
NAND2_X1 U993 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NAND2_X1 U994 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
XOR2_X1 U995 ( .A(KEYINPUT43), .B(n1306), .Z(n1302) );
NOR2_X1 U996 ( .A1(n1304), .A2(n1305), .ZN(n1306) );
XNOR2_X1 U997 ( .A(n1307), .B(n1308), .ZN(n1305) );
NOR2_X1 U998 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XNOR2_X1 U999 ( .A(n1120), .B(KEYINPUT52), .ZN(n1310) );
NOR2_X1 U1000 ( .A1(G140), .A2(n1258), .ZN(n1309) );
NAND2_X1 U1001 ( .A1(KEYINPUT61), .A2(n1242), .ZN(n1307) );
XNOR2_X1 U1002 ( .A(n1311), .B(n1312), .ZN(n1304) );
XOR2_X1 U1003 ( .A(G143), .B(G131), .Z(n1312) );
NAND3_X1 U1004 ( .A1(n1282), .A2(n1313), .A3(G214), .ZN(n1311) );
XOR2_X1 U1005 ( .A(n1314), .B(G478), .Z(n1267) );
NAND2_X1 U1006 ( .A1(n1315), .A2(n1181), .ZN(n1314) );
XOR2_X1 U1007 ( .A(KEYINPUT62), .B(n1158), .Z(n1315) );
INV_X1 U1008 ( .A(n1154), .ZN(n1158) );
XOR2_X1 U1009 ( .A(n1316), .B(n1317), .Z(n1154) );
XOR2_X1 U1010 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1011 ( .A(G107), .B(n1320), .Z(n1319) );
NOR2_X1 U1012 ( .A1(n1321), .A2(n1148), .ZN(n1320) );
INV_X1 U1013 ( .A(G217), .ZN(n1148) );
XOR2_X1 U1014 ( .A(n1271), .B(n1322), .Z(n1316) );
XOR2_X1 U1015 ( .A(G134), .B(G122), .Z(n1322) );
INV_X1 U1016 ( .A(G116), .ZN(n1271) );
NOR2_X1 U1017 ( .A1(n1264), .A2(n1057), .ZN(n1083) );
XNOR2_X1 U1018 ( .A(G472), .B(n1323), .ZN(n1057) );
NOR2_X1 U1019 ( .A1(KEYINPUT53), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1020 ( .A(n1100), .B(KEYINPUT47), .Z(n1324) );
NAND2_X1 U1021 ( .A1(n1325), .A2(n1181), .ZN(n1100) );
XOR2_X1 U1022 ( .A(n1326), .B(n1327), .Z(n1325) );
XOR2_X1 U1023 ( .A(n1328), .B(n1174), .Z(n1327) );
INV_X1 U1024 ( .A(n1201), .ZN(n1174) );
NOR2_X1 U1025 ( .A1(KEYINPUT48), .A2(n1329), .ZN(n1328) );
XNOR2_X1 U1026 ( .A(n1175), .B(n1291), .ZN(n1329) );
NAND3_X1 U1027 ( .A1(n1282), .A2(n1313), .A3(G210), .ZN(n1175) );
XOR2_X1 U1028 ( .A(n1290), .B(n1171), .Z(n1326) );
XOR2_X1 U1029 ( .A(G113), .B(n1330), .Z(n1171) );
NAND2_X1 U1030 ( .A1(n1331), .A2(n1332), .ZN(n1290) );
NAND2_X1 U1031 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
INV_X1 U1032 ( .A(G131), .ZN(n1334) );
XOR2_X1 U1033 ( .A(KEYINPUT36), .B(n1335), .Z(n1333) );
NAND2_X1 U1034 ( .A1(n1336), .A2(G131), .ZN(n1331) );
XOR2_X1 U1035 ( .A(KEYINPUT33), .B(n1335), .Z(n1336) );
XOR2_X1 U1036 ( .A(n1337), .B(n1247), .Z(n1335) );
INV_X1 U1037 ( .A(G137), .ZN(n1247) );
NAND2_X1 U1038 ( .A1(KEYINPUT58), .A2(n1249), .ZN(n1337) );
INV_X1 U1039 ( .A(G134), .ZN(n1249) );
INV_X1 U1040 ( .A(n1055), .ZN(n1264) );
XOR2_X1 U1041 ( .A(n1338), .B(n1091), .Z(n1055) );
NOR2_X1 U1042 ( .A1(n1145), .A2(G902), .ZN(n1091) );
XOR2_X1 U1043 ( .A(n1339), .B(n1340), .Z(n1145) );
XOR2_X1 U1044 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1045 ( .A(G110), .B(n1343), .Z(n1342) );
NOR2_X1 U1046 ( .A1(KEYINPUT15), .A2(n1344), .ZN(n1343) );
XOR2_X1 U1047 ( .A(n1345), .B(G146), .Z(n1344) );
NAND2_X1 U1048 ( .A1(KEYINPUT21), .A2(n1346), .ZN(n1345) );
NAND2_X1 U1049 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
NAND2_X1 U1050 ( .A1(G125), .A2(n1349), .ZN(n1348) );
NAND2_X1 U1051 ( .A1(KEYINPUT17), .A2(G140), .ZN(n1349) );
NAND2_X1 U1052 ( .A1(KEYINPUT17), .A2(n1120), .ZN(n1347) );
NOR2_X1 U1053 ( .A1(n1124), .A2(G125), .ZN(n1120) );
INV_X1 U1054 ( .A(G140), .ZN(n1124) );
NOR2_X1 U1055 ( .A1(n1350), .A2(n1321), .ZN(n1341) );
NAND2_X1 U1056 ( .A1(G234), .A2(n1282), .ZN(n1321) );
INV_X1 U1057 ( .A(G221), .ZN(n1350) );
XNOR2_X1 U1058 ( .A(G119), .B(n1351), .ZN(n1339) );
XOR2_X1 U1059 ( .A(G137), .B(G128), .Z(n1351) );
NAND2_X1 U1060 ( .A1(KEYINPUT2), .A2(n1094), .ZN(n1338) );
NAND2_X1 U1061 ( .A1(G217), .A2(n1352), .ZN(n1094) );
XOR2_X1 U1062 ( .A(KEYINPUT41), .B(n1353), .Z(n1352) );
AND2_X1 U1063 ( .A1(n1181), .A2(G234), .ZN(n1353) );
NAND2_X1 U1064 ( .A1(n1354), .A2(n1073), .ZN(n1238) );
NAND2_X1 U1065 ( .A1(G214), .A2(n1355), .ZN(n1073) );
INV_X1 U1066 ( .A(n1253), .ZN(n1354) );
XNOR2_X1 U1067 ( .A(n1103), .B(KEYINPUT63), .ZN(n1253) );
XNOR2_X1 U1068 ( .A(n1356), .B(n1205), .ZN(n1103) );
AND2_X1 U1069 ( .A1(G210), .A2(n1355), .ZN(n1205) );
NAND2_X1 U1070 ( .A1(n1313), .A2(n1181), .ZN(n1355) );
INV_X1 U1071 ( .A(G237), .ZN(n1313) );
NAND2_X1 U1072 ( .A1(n1357), .A2(n1181), .ZN(n1356) );
INV_X1 U1073 ( .A(G902), .ZN(n1181) );
XOR2_X1 U1074 ( .A(n1358), .B(n1359), .Z(n1357) );
XOR2_X1 U1075 ( .A(n1258), .B(n1192), .Z(n1359) );
NAND2_X1 U1076 ( .A1(G224), .A2(n1282), .ZN(n1192) );
XOR2_X1 U1077 ( .A(G953), .B(KEYINPUT46), .Z(n1282) );
INV_X1 U1078 ( .A(G125), .ZN(n1258) );
XOR2_X1 U1079 ( .A(n1204), .B(n1201), .Z(n1358) );
XOR2_X1 U1080 ( .A(n1285), .B(KEYINPUT8), .Z(n1201) );
XOR2_X1 U1081 ( .A(n1360), .B(n1318), .Z(n1285) );
XOR2_X1 U1082 ( .A(G128), .B(G143), .Z(n1318) );
XOR2_X1 U1083 ( .A(n1242), .B(KEYINPUT59), .Z(n1360) );
INV_X1 U1084 ( .A(G146), .ZN(n1242) );
XNOR2_X1 U1085 ( .A(n1361), .B(n1139), .ZN(n1204) );
XOR2_X1 U1086 ( .A(G110), .B(G122), .Z(n1139) );
NAND3_X1 U1087 ( .A1(n1362), .A2(n1363), .A3(n1364), .ZN(n1361) );
NAND2_X1 U1088 ( .A1(n1137), .A2(n1365), .ZN(n1364) );
INV_X1 U1089 ( .A(KEYINPUT55), .ZN(n1365) );
NAND3_X1 U1090 ( .A1(KEYINPUT55), .A2(n1366), .A3(n1138), .ZN(n1363) );
OR2_X1 U1091 ( .A1(n1138), .A2(n1366), .ZN(n1362) );
NOR2_X1 U1092 ( .A1(n1367), .A2(n1137), .ZN(n1366) );
XNOR2_X1 U1093 ( .A(n1368), .B(n1330), .ZN(n1137) );
XOR2_X1 U1094 ( .A(G119), .B(G116), .Z(n1330) );
NAND2_X1 U1095 ( .A1(KEYINPUT6), .A2(G113), .ZN(n1368) );
INV_X1 U1096 ( .A(KEYINPUT30), .ZN(n1367) );
NAND3_X1 U1097 ( .A1(n1369), .A2(n1370), .A3(n1371), .ZN(n1138) );
NAND2_X1 U1098 ( .A1(KEYINPUT7), .A2(n1372), .ZN(n1371) );
NAND3_X1 U1099 ( .A1(n1373), .A2(n1374), .A3(n1291), .ZN(n1370) );
INV_X1 U1100 ( .A(KEYINPUT7), .ZN(n1374) );
OR2_X1 U1101 ( .A1(n1291), .A2(n1373), .ZN(n1369) );
NOR2_X1 U1102 ( .A1(KEYINPUT12), .A2(n1372), .ZN(n1373) );
XOR2_X1 U1103 ( .A(n1163), .B(G107), .Z(n1372) );
INV_X1 U1104 ( .A(G104), .ZN(n1163) );
XNOR2_X1 U1105 ( .A(G101), .B(KEYINPUT11), .ZN(n1291) );
endmodule


