//Key = 1100000001000011001000011010111100101110000000110011011000100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308;

XOR2_X1 U733 ( .A(G107), .B(n1004), .Z(G9) );
NOR2_X1 U734 ( .A1(n1005), .A2(n1006), .ZN(G75) );
NOR3_X1 U735 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1006) );
NAND3_X1 U736 ( .A1(n1010), .A2(n1011), .A3(n1012), .ZN(n1007) );
NAND2_X1 U737 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U738 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND3_X1 U739 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1016) );
NAND3_X1 U740 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1018) );
NAND2_X1 U741 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U742 ( .A1(n1025), .A2(n1026), .ZN(n1020) );
NAND2_X1 U743 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U744 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND3_X1 U745 ( .A1(n1023), .A2(n1031), .A3(n1025), .ZN(n1015) );
NAND3_X1 U746 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NAND2_X1 U747 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
XNOR2_X1 U748 ( .A(KEYINPUT30), .B(n1017), .ZN(n1035) );
NAND2_X1 U749 ( .A1(n1019), .A2(n1037), .ZN(n1032) );
NAND2_X1 U750 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U751 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
INV_X1 U752 ( .A(n1042), .ZN(n1013) );
NOR3_X1 U753 ( .A1(n1043), .A2(G953), .A3(n1044), .ZN(n1005) );
INV_X1 U754 ( .A(n1010), .ZN(n1044) );
NAND4_X1 U755 ( .A1(n1023), .A2(n1019), .A3(n1045), .A4(n1046), .ZN(n1010) );
NOR3_X1 U756 ( .A1(n1047), .A2(n1040), .A3(n1048), .ZN(n1046) );
XOR2_X1 U757 ( .A(n1049), .B(n1050), .Z(n1048) );
NOR2_X1 U758 ( .A1(G478), .A2(KEYINPUT27), .ZN(n1050) );
XNOR2_X1 U759 ( .A(n1051), .B(KEYINPUT8), .ZN(n1045) );
XNOR2_X1 U760 ( .A(KEYINPUT43), .B(n1008), .ZN(n1043) );
INV_X1 U761 ( .A(G952), .ZN(n1008) );
XOR2_X1 U762 ( .A(n1052), .B(n1053), .Z(G72) );
NOR2_X1 U763 ( .A1(KEYINPUT39), .A2(n1054), .ZN(n1053) );
NOR2_X1 U764 ( .A1(n1055), .A2(n1011), .ZN(n1054) );
NOR2_X1 U765 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND3_X1 U766 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1052) );
NAND2_X1 U767 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
OR3_X1 U768 ( .A1(n1062), .A2(n1061), .A3(n1063), .ZN(n1059) );
OR2_X1 U769 ( .A1(KEYINPUT49), .A2(n1064), .ZN(n1061) );
NAND2_X1 U770 ( .A1(n1065), .A2(n1066), .ZN(n1062) );
NAND2_X1 U771 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XNOR2_X1 U772 ( .A(KEYINPUT63), .B(n1069), .ZN(n1068) );
XNOR2_X1 U773 ( .A(KEYINPUT47), .B(n1011), .ZN(n1065) );
NAND2_X1 U774 ( .A1(n1064), .A2(n1063), .ZN(n1058) );
INV_X1 U775 ( .A(KEYINPUT1), .ZN(n1063) );
NAND3_X1 U776 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1064) );
XOR2_X1 U777 ( .A(n1073), .B(KEYINPUT56), .Z(n1072) );
NAND2_X1 U778 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
OR2_X1 U779 ( .A1(n1075), .A2(n1074), .ZN(n1071) );
XOR2_X1 U780 ( .A(n1076), .B(n1077), .Z(n1074) );
XNOR2_X1 U781 ( .A(n1078), .B(G131), .ZN(n1077) );
XNOR2_X1 U782 ( .A(n1079), .B(n1080), .ZN(n1076) );
NOR2_X1 U783 ( .A1(KEYINPUT41), .A2(n1081), .ZN(n1080) );
NAND2_X1 U784 ( .A1(n1082), .A2(n1083), .ZN(n1075) );
NAND2_X1 U785 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XOR2_X1 U786 ( .A(KEYINPUT23), .B(n1086), .Z(n1082) );
NOR2_X1 U787 ( .A1(n1084), .A2(n1085), .ZN(n1086) );
NAND2_X1 U788 ( .A1(n1087), .A2(n1057), .ZN(n1070) );
XOR2_X1 U789 ( .A(n1088), .B(n1089), .Z(G69) );
XOR2_X1 U790 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U791 ( .A1(n1092), .A2(G953), .ZN(n1091) );
NOR2_X1 U792 ( .A1(n1093), .A2(n1094), .ZN(n1090) );
XNOR2_X1 U793 ( .A(n1095), .B(n1096), .ZN(n1094) );
NOR2_X1 U794 ( .A1(KEYINPUT48), .A2(n1097), .ZN(n1096) );
AND2_X1 U795 ( .A1(n1098), .A2(n1087), .ZN(n1093) );
NOR2_X1 U796 ( .A1(n1099), .A2(n1011), .ZN(n1088) );
AND2_X1 U797 ( .A1(G224), .A2(G898), .ZN(n1099) );
NOR2_X1 U798 ( .A1(n1100), .A2(n1101), .ZN(G66) );
XOR2_X1 U799 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND3_X1 U800 ( .A1(n1104), .A2(G217), .A3(KEYINPUT14), .ZN(n1102) );
NOR3_X1 U801 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(G63) );
AND2_X1 U802 ( .A1(KEYINPUT26), .A2(n1100), .ZN(n1107) );
NOR3_X1 U803 ( .A1(KEYINPUT26), .A2(G953), .A3(G952), .ZN(n1106) );
XOR2_X1 U804 ( .A(n1108), .B(n1109), .Z(n1105) );
NOR2_X1 U805 ( .A1(KEYINPUT2), .A2(n1110), .ZN(n1109) );
XOR2_X1 U806 ( .A(n1111), .B(n1112), .Z(n1110) );
NAND2_X1 U807 ( .A1(n1104), .A2(G478), .ZN(n1108) );
NOR2_X1 U808 ( .A1(n1100), .A2(n1113), .ZN(G60) );
NOR2_X1 U809 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U810 ( .A(n1116), .B(n1117), .Z(n1115) );
AND2_X1 U811 ( .A1(G475), .A2(n1104), .ZN(n1117) );
NOR2_X1 U812 ( .A1(KEYINPUT33), .A2(n1118), .ZN(n1116) );
AND2_X1 U813 ( .A1(n1118), .A2(KEYINPUT33), .ZN(n1114) );
XNOR2_X1 U814 ( .A(G104), .B(n1119), .ZN(G6) );
NOR2_X1 U815 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
AND2_X1 U816 ( .A1(KEYINPUT29), .A2(n1122), .ZN(n1121) );
NOR3_X1 U817 ( .A1(KEYINPUT29), .A2(n1123), .A3(n1124), .ZN(n1120) );
AND4_X1 U818 ( .A1(n1125), .A2(n1126), .A3(n1019), .A4(n1127), .ZN(n1123) );
NOR2_X1 U819 ( .A1(n1100), .A2(n1128), .ZN(G57) );
XOR2_X1 U820 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U821 ( .A(n1131), .B(n1132), .Z(n1130) );
AND2_X1 U822 ( .A1(G472), .A2(n1104), .ZN(n1131) );
XOR2_X1 U823 ( .A(n1133), .B(n1134), .Z(n1129) );
XOR2_X1 U824 ( .A(n1135), .B(n1136), .Z(n1134) );
NAND2_X1 U825 ( .A1(KEYINPUT62), .A2(G101), .ZN(n1136) );
NAND2_X1 U826 ( .A1(n1137), .A2(KEYINPUT0), .ZN(n1133) );
XOR2_X1 U827 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U828 ( .A1(KEYINPUT60), .A2(n1140), .ZN(n1139) );
NOR2_X1 U829 ( .A1(n1100), .A2(n1141), .ZN(G54) );
XOR2_X1 U830 ( .A(n1142), .B(n1143), .Z(n1141) );
AND2_X1 U831 ( .A1(G469), .A2(n1104), .ZN(n1143) );
INV_X1 U832 ( .A(n1144), .ZN(n1104) );
NAND2_X1 U833 ( .A1(n1145), .A2(n1146), .ZN(n1142) );
XOR2_X1 U834 ( .A(KEYINPUT31), .B(KEYINPUT19), .Z(n1146) );
XOR2_X1 U835 ( .A(n1147), .B(n1148), .Z(n1145) );
XNOR2_X1 U836 ( .A(n1149), .B(n1079), .ZN(n1148) );
NAND2_X1 U837 ( .A1(KEYINPUT28), .A2(n1150), .ZN(n1149) );
XOR2_X1 U838 ( .A(KEYINPUT12), .B(n1151), .Z(n1150) );
XOR2_X1 U839 ( .A(n1152), .B(n1153), .Z(n1147) );
NOR2_X1 U840 ( .A1(n1100), .A2(n1154), .ZN(G51) );
XOR2_X1 U841 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U842 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XOR2_X1 U843 ( .A(n1159), .B(KEYINPUT36), .Z(n1158) );
NAND2_X1 U844 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NOR2_X1 U845 ( .A1(n1161), .A2(n1160), .ZN(n1157) );
XNOR2_X1 U846 ( .A(n1162), .B(n1163), .ZN(n1160) );
NOR2_X1 U847 ( .A1(KEYINPUT11), .A2(n1164), .ZN(n1163) );
NOR2_X1 U848 ( .A1(n1165), .A2(n1144), .ZN(n1155) );
NAND2_X1 U849 ( .A1(G902), .A2(n1009), .ZN(n1144) );
NAND3_X1 U850 ( .A1(n1067), .A2(n1069), .A3(n1092), .ZN(n1009) );
AND2_X1 U851 ( .A1(n1166), .A2(n1167), .ZN(n1092) );
NOR4_X1 U852 ( .A1(n1168), .A2(n1004), .A3(n1122), .A4(n1169), .ZN(n1167) );
AND3_X1 U853 ( .A1(n1170), .A2(n1019), .A3(n1127), .ZN(n1122) );
AND3_X1 U854 ( .A1(n1019), .A2(n1024), .A3(n1170), .ZN(n1004) );
AND4_X1 U855 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1166) );
OR2_X1 U856 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
AND4_X1 U857 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1067) );
NOR3_X1 U858 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
INV_X1 U859 ( .A(n1184), .ZN(n1181) );
NAND2_X1 U860 ( .A1(n1185), .A2(n1186), .ZN(n1179) );
NAND2_X1 U861 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND3_X1 U862 ( .A1(n1036), .A2(n1189), .A3(n1190), .ZN(n1188) );
XNOR2_X1 U863 ( .A(KEYINPUT37), .B(n1191), .ZN(n1187) );
NAND3_X1 U864 ( .A1(n1192), .A2(n1017), .A3(n1025), .ZN(n1177) );
NOR2_X1 U865 ( .A1(n1011), .A2(G952), .ZN(n1100) );
XNOR2_X1 U866 ( .A(G146), .B(n1069), .ZN(G48) );
NAND3_X1 U867 ( .A1(n1192), .A2(n1185), .A3(n1127), .ZN(n1069) );
XNOR2_X1 U868 ( .A(G143), .B(n1178), .ZN(G45) );
NAND4_X1 U869 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1185), .ZN(n1178) );
NOR2_X1 U870 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND2_X1 U871 ( .A1(n1198), .A2(n1199), .ZN(G42) );
OR2_X1 U872 ( .A1(n1184), .A2(G140), .ZN(n1199) );
XOR2_X1 U873 ( .A(n1200), .B(KEYINPUT32), .Z(n1198) );
NAND2_X1 U874 ( .A1(G140), .A2(n1184), .ZN(n1200) );
NAND4_X1 U875 ( .A1(n1036), .A2(n1127), .A3(n1194), .A4(n1017), .ZN(n1184) );
XNOR2_X1 U876 ( .A(G137), .B(n1201), .ZN(G39) );
NAND3_X1 U877 ( .A1(n1025), .A2(n1192), .A3(n1202), .ZN(n1201) );
XNOR2_X1 U878 ( .A(KEYINPUT54), .B(n1017), .ZN(n1202) );
XOR2_X1 U879 ( .A(n1183), .B(n1203), .Z(G36) );
NOR2_X1 U880 ( .A1(KEYINPUT35), .A2(n1081), .ZN(n1203) );
AND3_X1 U881 ( .A1(n1194), .A2(n1024), .A3(n1204), .ZN(n1183) );
XNOR2_X1 U882 ( .A(G131), .B(n1205), .ZN(G33) );
NOR2_X1 U883 ( .A1(n1182), .A2(KEYINPUT55), .ZN(n1205) );
AND3_X1 U884 ( .A1(n1127), .A2(n1194), .A3(n1204), .ZN(n1182) );
INV_X1 U885 ( .A(n1033), .ZN(n1204) );
NAND2_X1 U886 ( .A1(n1193), .A2(n1017), .ZN(n1033) );
NAND2_X1 U887 ( .A1(n1206), .A2(n1207), .ZN(n1017) );
OR3_X1 U888 ( .A1(n1051), .A2(n1040), .A3(KEYINPUT44), .ZN(n1207) );
NAND2_X1 U889 ( .A1(KEYINPUT44), .A2(n1185), .ZN(n1206) );
XOR2_X1 U890 ( .A(n1208), .B(n1209), .Z(G30) );
NOR2_X1 U891 ( .A1(n1038), .A2(n1191), .ZN(n1209) );
NAND2_X1 U892 ( .A1(n1192), .A2(n1024), .ZN(n1191) );
AND3_X1 U893 ( .A1(n1210), .A2(n1211), .A3(n1194), .ZN(n1192) );
AND2_X1 U894 ( .A1(n1126), .A2(n1189), .ZN(n1194) );
INV_X1 U895 ( .A(n1185), .ZN(n1038) );
NOR2_X1 U896 ( .A1(KEYINPUT7), .A2(n1212), .ZN(n1208) );
XOR2_X1 U897 ( .A(n1173), .B(n1213), .Z(G3) );
NAND2_X1 U898 ( .A1(KEYINPUT24), .A2(G101), .ZN(n1213) );
NAND3_X1 U899 ( .A1(n1025), .A2(n1170), .A3(n1193), .ZN(n1173) );
XOR2_X1 U900 ( .A(n1214), .B(n1215), .Z(G27) );
XNOR2_X1 U901 ( .A(KEYINPUT59), .B(n1085), .ZN(n1215) );
INV_X1 U902 ( .A(G125), .ZN(n1085) );
NAND2_X1 U903 ( .A1(KEYINPUT46), .A2(n1216), .ZN(n1214) );
NAND4_X1 U904 ( .A1(n1190), .A2(n1185), .A3(n1217), .A4(n1189), .ZN(n1216) );
NAND2_X1 U905 ( .A1(n1042), .A2(n1218), .ZN(n1189) );
NAND4_X1 U906 ( .A1(n1087), .A2(G902), .A3(n1219), .A4(n1057), .ZN(n1218) );
INV_X1 U907 ( .A(G900), .ZN(n1057) );
XOR2_X1 U908 ( .A(KEYINPUT10), .B(n1036), .Z(n1217) );
XNOR2_X1 U909 ( .A(G122), .B(n1172), .ZN(G24) );
NAND4_X1 U910 ( .A1(n1220), .A2(n1019), .A3(n1221), .A4(n1047), .ZN(n1172) );
NOR2_X1 U911 ( .A1(n1211), .A2(n1210), .ZN(n1019) );
XNOR2_X1 U912 ( .A(G119), .B(n1171), .ZN(G21) );
NAND4_X1 U913 ( .A1(n1220), .A2(n1025), .A3(n1210), .A4(n1211), .ZN(n1171) );
XNOR2_X1 U914 ( .A(n1169), .B(n1222), .ZN(G18) );
NAND2_X1 U915 ( .A1(KEYINPUT9), .A2(G116), .ZN(n1222) );
AND3_X1 U916 ( .A1(n1220), .A2(n1024), .A3(n1193), .ZN(n1169) );
NOR2_X1 U917 ( .A1(n1047), .A2(n1197), .ZN(n1024) );
INV_X1 U918 ( .A(n1221), .ZN(n1197) );
AND3_X1 U919 ( .A1(n1185), .A2(n1125), .A3(n1023), .ZN(n1220) );
XOR2_X1 U920 ( .A(G113), .B(n1223), .Z(G15) );
NOR2_X1 U921 ( .A1(n1176), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U922 ( .A(KEYINPUT4), .B(n1125), .ZN(n1224) );
NAND3_X1 U923 ( .A1(n1193), .A2(n1225), .A3(n1190), .ZN(n1176) );
INV_X1 U924 ( .A(n1021), .ZN(n1190) );
NAND2_X1 U925 ( .A1(n1127), .A2(n1023), .ZN(n1021) );
NOR2_X1 U926 ( .A1(n1226), .A2(n1029), .ZN(n1023) );
NOR2_X1 U927 ( .A1(n1221), .A2(n1196), .ZN(n1127) );
INV_X1 U928 ( .A(n1047), .ZN(n1196) );
NOR2_X1 U929 ( .A1(n1211), .A2(n1227), .ZN(n1193) );
XOR2_X1 U930 ( .A(n1228), .B(n1229), .Z(G12) );
XNOR2_X1 U931 ( .A(G110), .B(KEYINPUT45), .ZN(n1229) );
NAND2_X1 U932 ( .A1(KEYINPUT53), .A2(n1168), .ZN(n1228) );
AND3_X1 U933 ( .A1(n1025), .A2(n1170), .A3(n1036), .ZN(n1168) );
AND2_X1 U934 ( .A1(n1227), .A2(n1211), .ZN(n1036) );
NAND3_X1 U935 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1211) );
OR2_X1 U936 ( .A1(n1233), .A2(n1103), .ZN(n1232) );
NAND3_X1 U937 ( .A1(n1103), .A2(n1233), .A3(n1234), .ZN(n1231) );
NAND2_X1 U938 ( .A1(G217), .A2(n1235), .ZN(n1233) );
XOR2_X1 U939 ( .A(n1236), .B(n1237), .Z(n1103) );
XOR2_X1 U940 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U941 ( .A(G119), .B(G110), .Z(n1239) );
XNOR2_X1 U942 ( .A(KEYINPUT17), .B(n1212), .ZN(n1238) );
INV_X1 U943 ( .A(G128), .ZN(n1212) );
XOR2_X1 U944 ( .A(n1240), .B(n1241), .Z(n1236) );
XNOR2_X1 U945 ( .A(n1242), .B(n1243), .ZN(n1241) );
NOR2_X1 U946 ( .A1(KEYINPUT16), .A2(G137), .ZN(n1243) );
NAND2_X1 U947 ( .A1(KEYINPUT50), .A2(n1244), .ZN(n1242) );
XNOR2_X1 U948 ( .A(n1245), .B(n1246), .ZN(n1244) );
INV_X1 U949 ( .A(n1247), .ZN(n1246) );
NOR2_X1 U950 ( .A1(KEYINPUT22), .A2(n1248), .ZN(n1245) );
NAND2_X1 U951 ( .A1(n1249), .A2(G221), .ZN(n1240) );
NAND2_X1 U952 ( .A1(G217), .A2(G902), .ZN(n1230) );
INV_X1 U953 ( .A(n1210), .ZN(n1227) );
XNOR2_X1 U954 ( .A(n1250), .B(G472), .ZN(n1210) );
NAND2_X1 U955 ( .A1(n1251), .A2(n1234), .ZN(n1250) );
XOR2_X1 U956 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U957 ( .A(n1138), .B(n1132), .Z(n1253) );
XNOR2_X1 U958 ( .A(n1254), .B(n1255), .ZN(n1132) );
NOR2_X1 U959 ( .A1(G116), .A2(KEYINPUT40), .ZN(n1255) );
XNOR2_X1 U960 ( .A(n1256), .B(n1257), .ZN(n1252) );
XOR2_X1 U961 ( .A(n1135), .B(G101), .Z(n1256) );
NAND2_X1 U962 ( .A1(n1258), .A2(G210), .ZN(n1135) );
NOR3_X1 U963 ( .A1(n1124), .A2(n1175), .A3(n1027), .ZN(n1170) );
INV_X1 U964 ( .A(n1126), .ZN(n1027) );
NOR2_X1 U965 ( .A1(n1030), .A2(n1029), .ZN(n1126) );
AND2_X1 U966 ( .A1(G221), .A2(n1259), .ZN(n1029) );
NAND2_X1 U967 ( .A1(G234), .A2(n1234), .ZN(n1259) );
INV_X1 U968 ( .A(n1226), .ZN(n1030) );
XNOR2_X1 U969 ( .A(n1260), .B(G469), .ZN(n1226) );
NAND2_X1 U970 ( .A1(n1261), .A2(n1234), .ZN(n1260) );
XOR2_X1 U971 ( .A(n1152), .B(n1262), .Z(n1261) );
XNOR2_X1 U972 ( .A(n1151), .B(n1263), .ZN(n1262) );
NOR2_X1 U973 ( .A1(KEYINPUT6), .A2(n1264), .ZN(n1263) );
XNOR2_X1 U974 ( .A(n1265), .B(n1266), .ZN(n1264) );
XNOR2_X1 U975 ( .A(n1267), .B(KEYINPUT21), .ZN(n1266) );
NAND2_X1 U976 ( .A1(KEYINPUT34), .A2(n1153), .ZN(n1267) );
XOR2_X1 U977 ( .A(G101), .B(n1268), .Z(n1153) );
INV_X1 U978 ( .A(n1079), .ZN(n1265) );
XOR2_X1 U979 ( .A(G110), .B(n1084), .Z(n1151) );
XOR2_X1 U980 ( .A(n1138), .B(n1269), .Z(n1152) );
NOR2_X1 U981 ( .A1(G953), .A2(n1056), .ZN(n1269) );
INV_X1 U982 ( .A(G227), .ZN(n1056) );
XOR2_X1 U983 ( .A(n1270), .B(G131), .Z(n1138) );
NAND2_X1 U984 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND2_X1 U985 ( .A1(G134), .A2(n1078), .ZN(n1272) );
XOR2_X1 U986 ( .A(KEYINPUT15), .B(n1273), .Z(n1271) );
NOR2_X1 U987 ( .A1(G134), .A2(n1078), .ZN(n1273) );
INV_X1 U988 ( .A(G137), .ZN(n1078) );
INV_X1 U989 ( .A(n1125), .ZN(n1175) );
NAND2_X1 U990 ( .A1(n1042), .A2(n1274), .ZN(n1125) );
NAND4_X1 U991 ( .A1(n1087), .A2(G902), .A3(n1219), .A4(n1098), .ZN(n1274) );
INV_X1 U992 ( .A(G898), .ZN(n1098) );
XNOR2_X1 U993 ( .A(G953), .B(KEYINPUT58), .ZN(n1087) );
NAND3_X1 U994 ( .A1(n1219), .A2(n1011), .A3(G952), .ZN(n1042) );
NAND2_X1 U995 ( .A1(G237), .A2(G234), .ZN(n1219) );
INV_X1 U996 ( .A(n1225), .ZN(n1124) );
XOR2_X1 U997 ( .A(n1185), .B(KEYINPUT52), .Z(n1225) );
NOR2_X1 U998 ( .A1(n1041), .A2(n1040), .ZN(n1185) );
AND2_X1 U999 ( .A1(G214), .A2(n1275), .ZN(n1040) );
INV_X1 U1000 ( .A(n1051), .ZN(n1041) );
XOR2_X1 U1001 ( .A(n1276), .B(n1165), .Z(n1051) );
NAND2_X1 U1002 ( .A1(G210), .A2(n1275), .ZN(n1165) );
NAND2_X1 U1003 ( .A1(n1277), .A2(n1234), .ZN(n1275) );
INV_X1 U1004 ( .A(G237), .ZN(n1277) );
NAND2_X1 U1005 ( .A1(n1278), .A2(n1234), .ZN(n1276) );
XNOR2_X1 U1006 ( .A(n1161), .B(n1279), .ZN(n1278) );
NOR2_X1 U1007 ( .A1(KEYINPUT3), .A2(n1280), .ZN(n1279) );
XOR2_X1 U1008 ( .A(n1281), .B(n1164), .Z(n1280) );
NAND2_X1 U1009 ( .A1(G224), .A2(n1011), .ZN(n1164) );
INV_X1 U1010 ( .A(G953), .ZN(n1011) );
NAND3_X1 U1011 ( .A1(n1282), .A2(n1283), .A3(KEYINPUT61), .ZN(n1281) );
OR2_X1 U1012 ( .A1(n1162), .A2(KEYINPUT20), .ZN(n1283) );
XOR2_X1 U1013 ( .A(n1284), .B(n1140), .Z(n1162) );
NAND3_X1 U1014 ( .A1(n1284), .A2(n1257), .A3(KEYINPUT20), .ZN(n1282) );
INV_X1 U1015 ( .A(n1140), .ZN(n1257) );
XOR2_X1 U1016 ( .A(n1079), .B(KEYINPUT5), .Z(n1140) );
XOR2_X1 U1017 ( .A(G128), .B(n1285), .Z(n1079) );
XNOR2_X1 U1018 ( .A(G125), .B(KEYINPUT18), .ZN(n1284) );
XNOR2_X1 U1019 ( .A(n1097), .B(n1286), .ZN(n1161) );
INV_X1 U1020 ( .A(n1095), .ZN(n1286) );
XNOR2_X1 U1021 ( .A(n1254), .B(n1287), .ZN(n1095) );
XOR2_X1 U1022 ( .A(G116), .B(n1288), .Z(n1287) );
NOR2_X1 U1023 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XOR2_X1 U1024 ( .A(n1291), .B(KEYINPUT51), .Z(n1290) );
NAND2_X1 U1025 ( .A1(G101), .A2(n1292), .ZN(n1291) );
NOR2_X1 U1026 ( .A1(G101), .A2(n1292), .ZN(n1289) );
XOR2_X1 U1027 ( .A(KEYINPUT42), .B(n1268), .Z(n1292) );
XOR2_X1 U1028 ( .A(G104), .B(G107), .Z(n1268) );
XNOR2_X1 U1029 ( .A(G113), .B(G119), .ZN(n1254) );
XNOR2_X1 U1030 ( .A(G110), .B(n1293), .ZN(n1097) );
INV_X1 U1031 ( .A(G122), .ZN(n1293) );
NOR2_X1 U1032 ( .A1(n1221), .A2(n1047), .ZN(n1025) );
XNOR2_X1 U1033 ( .A(n1294), .B(G475), .ZN(n1047) );
OR2_X1 U1034 ( .A1(n1118), .A2(G902), .ZN(n1294) );
XNOR2_X1 U1035 ( .A(n1295), .B(n1296), .ZN(n1118) );
XOR2_X1 U1036 ( .A(G104), .B(n1297), .Z(n1296) );
NOR2_X1 U1037 ( .A1(KEYINPUT13), .A2(n1298), .ZN(n1297) );
XOR2_X1 U1038 ( .A(n1299), .B(n1300), .Z(n1298) );
XNOR2_X1 U1039 ( .A(n1247), .B(n1285), .ZN(n1300) );
XNOR2_X1 U1040 ( .A(G143), .B(n1248), .ZN(n1285) );
INV_X1 U1041 ( .A(G146), .ZN(n1248) );
XOR2_X1 U1042 ( .A(G125), .B(n1084), .Z(n1247) );
XOR2_X1 U1043 ( .A(G140), .B(KEYINPUT57), .Z(n1084) );
XOR2_X1 U1044 ( .A(n1301), .B(G131), .Z(n1299) );
NAND2_X1 U1045 ( .A1(n1258), .A2(G214), .ZN(n1301) );
NOR2_X1 U1046 ( .A1(G953), .A2(G237), .ZN(n1258) );
XNOR2_X1 U1047 ( .A(G113), .B(G122), .ZN(n1295) );
XNOR2_X1 U1048 ( .A(n1049), .B(G478), .ZN(n1221) );
NAND2_X1 U1049 ( .A1(n1302), .A2(n1234), .ZN(n1049) );
INV_X1 U1050 ( .A(G902), .ZN(n1234) );
XNOR2_X1 U1051 ( .A(n1112), .B(n1111), .ZN(n1302) );
XOR2_X1 U1052 ( .A(n1303), .B(n1304), .Z(n1111) );
XOR2_X1 U1053 ( .A(G116), .B(G107), .Z(n1304) );
XOR2_X1 U1054 ( .A(n1305), .B(n1306), .Z(n1303) );
NOR2_X1 U1055 ( .A1(KEYINPUT25), .A2(G128), .ZN(n1306) );
NAND2_X1 U1056 ( .A1(n1249), .A2(G217), .ZN(n1305) );
NOR2_X1 U1057 ( .A1(n1235), .A2(G953), .ZN(n1249) );
INV_X1 U1058 ( .A(G234), .ZN(n1235) );
XNOR2_X1 U1059 ( .A(n1307), .B(n1308), .ZN(n1112) );
XNOR2_X1 U1060 ( .A(n1081), .B(G122), .ZN(n1308) );
INV_X1 U1061 ( .A(G134), .ZN(n1081) );
XNOR2_X1 U1062 ( .A(G143), .B(KEYINPUT38), .ZN(n1307) );
endmodule


