//Key = 0011110000100100101101010100110010011110110000000110001010101111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348;

XOR2_X1 U752 ( .A(G107), .B(n1035), .Z(G9) );
NOR2_X1 U753 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
XOR2_X1 U754 ( .A(KEYINPUT28), .B(n1038), .Z(n1037) );
NOR2_X1 U755 ( .A1(n1039), .A2(n1040), .ZN(G75) );
NOR4_X1 U756 ( .A1(n1041), .A2(n1042), .A3(G953), .A4(n1043), .ZN(n1040) );
NOR2_X1 U757 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U758 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR3_X1 U759 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
NOR2_X1 U760 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U761 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR2_X1 U762 ( .A1(n1055), .A2(n1056), .ZN(n1051) );
NOR2_X1 U763 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U764 ( .A1(n1059), .A2(n1054), .ZN(n1058) );
NOR2_X1 U765 ( .A1(n1060), .A2(n1061), .ZN(n1057) );
NOR2_X1 U766 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR4_X1 U767 ( .A1(n1064), .A2(n1061), .A3(n1054), .A4(n1056), .ZN(n1046) );
NOR2_X1 U768 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR2_X1 U769 ( .A1(n1067), .A2(n1050), .ZN(n1066) );
INV_X1 U770 ( .A(n1068), .ZN(n1050) );
NOR2_X1 U771 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR2_X1 U772 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR2_X1 U773 ( .A1(n1073), .A2(n1048), .ZN(n1065) );
NOR2_X1 U774 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND3_X1 U775 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1041) );
NOR3_X1 U776 ( .A1(n1043), .A2(G953), .A3(G952), .ZN(n1039) );
AND4_X1 U777 ( .A1(n1072), .A2(n1059), .A3(n1079), .A4(n1080), .ZN(n1043) );
NOR4_X1 U778 ( .A1(n1081), .A2(n1056), .A3(n1082), .A4(n1083), .ZN(n1080) );
XOR2_X1 U779 ( .A(n1084), .B(n1085), .Z(n1082) );
NOR2_X1 U780 ( .A1(n1086), .A2(KEYINPUT33), .ZN(n1085) );
NAND3_X1 U781 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1081) );
XNOR2_X1 U782 ( .A(G472), .B(n1090), .ZN(n1089) );
NOR2_X1 U783 ( .A1(KEYINPUT12), .A2(n1091), .ZN(n1090) );
OR2_X1 U784 ( .A1(G475), .A2(KEYINPUT29), .ZN(n1088) );
NAND3_X1 U785 ( .A1(G475), .A2(n1092), .A3(KEYINPUT29), .ZN(n1087) );
NOR3_X1 U786 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1079) );
XOR2_X1 U787 ( .A(n1096), .B(n1097), .Z(G72) );
XOR2_X1 U788 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U789 ( .A1(n1100), .A2(G953), .ZN(n1099) );
NOR2_X1 U790 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(n1098) );
XOR2_X1 U792 ( .A(n1105), .B(n1106), .Z(n1104) );
XOR2_X1 U793 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U794 ( .A(n1109), .B(KEYINPUT23), .Z(n1105) );
NAND2_X1 U795 ( .A1(KEYINPUT38), .A2(n1110), .ZN(n1109) );
XOR2_X1 U796 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U797 ( .A1(G137), .A2(KEYINPUT9), .ZN(n1111) );
NOR2_X1 U798 ( .A1(G900), .A2(n1113), .ZN(n1103) );
NOR2_X1 U799 ( .A1(n1114), .A2(n1115), .ZN(n1096) );
NOR2_X1 U800 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
XOR2_X1 U801 ( .A(n1118), .B(n1119), .Z(G69) );
XOR2_X1 U802 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U803 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XOR2_X1 U804 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U805 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U806 ( .A(n1128), .B(KEYINPUT52), .Z(n1124) );
NOR2_X1 U807 ( .A1(G898), .A2(n1113), .ZN(n1122) );
NAND2_X1 U808 ( .A1(n1115), .A2(n1129), .ZN(n1120) );
NAND2_X1 U809 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U810 ( .A1(G953), .A2(n1132), .ZN(n1118) );
NAND2_X1 U811 ( .A1(G898), .A2(G224), .ZN(n1132) );
NOR2_X1 U812 ( .A1(n1133), .A2(n1134), .ZN(G66) );
XOR2_X1 U813 ( .A(n1135), .B(n1136), .Z(n1134) );
NAND2_X1 U814 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
NOR2_X1 U815 ( .A1(n1133), .A2(n1139), .ZN(G63) );
XOR2_X1 U816 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR4_X1 U817 ( .A1(n1142), .A2(n1143), .A3(KEYINPUT48), .A4(n1144), .ZN(n1141) );
INV_X1 U818 ( .A(G478), .ZN(n1144) );
NOR2_X1 U819 ( .A1(n1145), .A2(n1146), .ZN(n1143) );
INV_X1 U820 ( .A(KEYINPUT59), .ZN(n1146) );
NOR2_X1 U821 ( .A1(G902), .A2(n1147), .ZN(n1145) );
NOR2_X1 U822 ( .A1(KEYINPUT59), .A2(n1137), .ZN(n1142) );
NOR2_X1 U823 ( .A1(n1148), .A2(n1149), .ZN(G60) );
XOR2_X1 U824 ( .A(KEYINPUT22), .B(n1133), .Z(n1149) );
XOR2_X1 U825 ( .A(n1150), .B(n1151), .Z(n1148) );
NAND2_X1 U826 ( .A1(n1137), .A2(G475), .ZN(n1150) );
XNOR2_X1 U827 ( .A(G104), .B(n1152), .ZN(G6) );
NOR2_X1 U828 ( .A1(n1133), .A2(n1153), .ZN(G57) );
XOR2_X1 U829 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U830 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U831 ( .A(n1158), .B(n1107), .Z(n1156) );
XOR2_X1 U832 ( .A(n1159), .B(n1160), .Z(n1154) );
XOR2_X1 U833 ( .A(KEYINPUT47), .B(n1161), .Z(n1160) );
AND2_X1 U834 ( .A1(G472), .A2(n1137), .ZN(n1161) );
NAND2_X1 U835 ( .A1(KEYINPUT19), .A2(n1162), .ZN(n1159) );
NOR2_X1 U836 ( .A1(n1133), .A2(n1163), .ZN(G54) );
XOR2_X1 U837 ( .A(n1164), .B(n1165), .Z(n1163) );
XNOR2_X1 U838 ( .A(n1166), .B(n1167), .ZN(n1165) );
XOR2_X1 U839 ( .A(n1168), .B(n1169), .Z(n1164) );
XOR2_X1 U840 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U841 ( .A1(KEYINPUT49), .A2(n1107), .ZN(n1171) );
NAND2_X1 U842 ( .A1(n1137), .A2(G469), .ZN(n1170) );
XOR2_X1 U843 ( .A(n1172), .B(KEYINPUT17), .Z(n1168) );
NOR2_X1 U844 ( .A1(n1133), .A2(n1173), .ZN(G51) );
XOR2_X1 U845 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U846 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U847 ( .A1(KEYINPUT13), .A2(n1178), .ZN(n1177) );
NAND2_X1 U848 ( .A1(n1137), .A2(n1086), .ZN(n1176) );
NOR2_X1 U849 ( .A1(n1179), .A2(n1147), .ZN(n1137) );
AND3_X1 U850 ( .A1(n1076), .A2(n1180), .A3(n1077), .ZN(n1147) );
INV_X1 U851 ( .A(n1102), .ZN(n1077) );
NAND3_X1 U852 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1102) );
NAND3_X1 U853 ( .A1(n1062), .A2(n1184), .A3(n1185), .ZN(n1183) );
NAND2_X1 U854 ( .A1(n1186), .A2(n1187), .ZN(n1184) );
NAND2_X1 U855 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XNOR2_X1 U856 ( .A(n1074), .B(KEYINPUT61), .ZN(n1188) );
NAND2_X1 U857 ( .A1(n1190), .A2(n1191), .ZN(n1186) );
XOR2_X1 U858 ( .A(n1192), .B(KEYINPUT7), .Z(n1191) );
XOR2_X1 U859 ( .A(KEYINPUT39), .B(n1070), .Z(n1190) );
XOR2_X1 U860 ( .A(KEYINPUT42), .B(n1078), .Z(n1180) );
AND2_X1 U861 ( .A1(n1193), .A2(n1130), .ZN(n1078) );
AND4_X1 U862 ( .A1(n1152), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1130) );
NOR4_X1 U863 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1196) );
OR2_X1 U864 ( .A1(n1036), .A2(n1053), .ZN(n1195) );
NAND3_X1 U865 ( .A1(n1062), .A2(n1068), .A3(n1201), .ZN(n1036) );
NAND4_X1 U866 ( .A1(n1063), .A2(n1038), .A3(n1201), .A4(n1068), .ZN(n1152) );
XOR2_X1 U867 ( .A(n1131), .B(KEYINPUT45), .Z(n1193) );
XOR2_X1 U868 ( .A(n1101), .B(KEYINPUT35), .Z(n1076) );
NAND4_X1 U869 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1101) );
NOR2_X1 U870 ( .A1(n1115), .A2(G952), .ZN(n1133) );
XNOR2_X1 U871 ( .A(G146), .B(n1203), .ZN(G48) );
OR2_X1 U872 ( .A1(n1206), .A2(n1207), .ZN(n1203) );
XOR2_X1 U873 ( .A(n1208), .B(n1209), .Z(G45) );
NAND2_X1 U874 ( .A1(KEYINPUT37), .A2(n1210), .ZN(n1209) );
INV_X1 U875 ( .A(n1202), .ZN(n1210) );
NAND4_X1 U876 ( .A1(n1211), .A2(n1070), .A3(n1212), .A4(n1213), .ZN(n1202) );
NAND2_X1 U877 ( .A1(n1214), .A2(n1215), .ZN(G42) );
NAND2_X1 U878 ( .A1(n1216), .A2(n1172), .ZN(n1215) );
NAND2_X1 U879 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NAND2_X1 U880 ( .A1(n1204), .A2(n1219), .ZN(n1218) );
INV_X1 U881 ( .A(KEYINPUT5), .ZN(n1219) );
NAND2_X1 U882 ( .A1(KEYINPUT5), .A2(n1220), .ZN(n1217) );
OR2_X1 U883 ( .A1(n1172), .A2(n1220), .ZN(n1214) );
NAND2_X1 U884 ( .A1(KEYINPUT63), .A2(n1204), .ZN(n1220) );
NAND4_X1 U885 ( .A1(n1189), .A2(n1185), .A3(n1063), .A4(n1075), .ZN(n1204) );
XOR2_X1 U886 ( .A(n1221), .B(n1205), .Z(G39) );
NAND4_X1 U887 ( .A1(n1189), .A2(n1185), .A3(n1222), .A4(n1192), .ZN(n1205) );
XOR2_X1 U888 ( .A(G134), .B(n1223), .Z(G36) );
NOR3_X1 U889 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1223) );
XOR2_X1 U890 ( .A(n1048), .B(KEYINPUT0), .Z(n1225) );
INV_X1 U891 ( .A(n1189), .ZN(n1048) );
XOR2_X1 U892 ( .A(n1227), .B(n1228), .Z(G33) );
NOR2_X1 U893 ( .A1(KEYINPUT51), .A2(n1182), .ZN(n1228) );
NAND3_X1 U894 ( .A1(n1189), .A2(n1063), .A3(n1211), .ZN(n1182) );
INV_X1 U895 ( .A(n1224), .ZN(n1211) );
NAND2_X1 U896 ( .A1(n1185), .A2(n1074), .ZN(n1224) );
NOR2_X1 U897 ( .A1(n1071), .A2(n1229), .ZN(n1189) );
INV_X1 U898 ( .A(n1072), .ZN(n1229) );
XNOR2_X1 U899 ( .A(G131), .B(KEYINPUT32), .ZN(n1227) );
XOR2_X1 U900 ( .A(G128), .B(n1230), .Z(G30) );
NOR2_X1 U901 ( .A1(n1226), .A2(n1206), .ZN(n1230) );
NAND3_X1 U902 ( .A1(n1070), .A2(n1192), .A3(n1185), .ZN(n1206) );
AND2_X1 U903 ( .A1(n1038), .A2(n1231), .ZN(n1185) );
XNOR2_X1 U904 ( .A(G101), .B(n1194), .ZN(G3) );
NAND4_X1 U905 ( .A1(n1074), .A2(n1222), .A3(n1038), .A4(n1201), .ZN(n1194) );
XNOR2_X1 U906 ( .A(n1181), .B(n1232), .ZN(G27) );
NOR2_X1 U907 ( .A1(KEYINPUT44), .A2(n1233), .ZN(n1232) );
NAND4_X1 U908 ( .A1(n1234), .A2(n1231), .A3(n1070), .A4(n1235), .ZN(n1181) );
NOR3_X1 U909 ( .A1(n1207), .A2(n1236), .A3(n1056), .ZN(n1235) );
NAND2_X1 U910 ( .A1(n1237), .A2(n1238), .ZN(n1231) );
NAND2_X1 U911 ( .A1(n1239), .A2(n1117), .ZN(n1237) );
INV_X1 U912 ( .A(G900), .ZN(n1117) );
XNOR2_X1 U913 ( .A(n1200), .B(n1240), .ZN(G24) );
NAND2_X1 U914 ( .A1(KEYINPUT4), .A2(G122), .ZN(n1240) );
AND4_X1 U915 ( .A1(n1241), .A2(n1068), .A3(n1212), .A4(n1213), .ZN(n1200) );
NOR2_X1 U916 ( .A1(n1242), .A2(n1083), .ZN(n1068) );
XOR2_X1 U917 ( .A(G119), .B(n1199), .Z(G21) );
AND3_X1 U918 ( .A1(n1222), .A2(n1192), .A3(n1241), .ZN(n1199) );
NAND2_X1 U919 ( .A1(n1243), .A2(n1244), .ZN(n1192) );
NAND3_X1 U920 ( .A1(n1083), .A2(n1242), .A3(n1245), .ZN(n1244) );
INV_X1 U921 ( .A(KEYINPUT8), .ZN(n1245) );
INV_X1 U922 ( .A(n1246), .ZN(n1242) );
NAND2_X1 U923 ( .A1(KEYINPUT8), .A2(n1074), .ZN(n1243) );
XNOR2_X1 U924 ( .A(G116), .B(n1131), .ZN(G18) );
NAND3_X1 U925 ( .A1(n1074), .A2(n1062), .A3(n1241), .ZN(n1131) );
INV_X1 U926 ( .A(n1226), .ZN(n1062) );
NAND2_X1 U927 ( .A1(n1247), .A2(n1212), .ZN(n1226) );
INV_X1 U928 ( .A(n1248), .ZN(n1212) );
XOR2_X1 U929 ( .A(n1198), .B(n1249), .Z(G15) );
NOR2_X1 U930 ( .A1(KEYINPUT53), .A2(n1250), .ZN(n1249) );
AND3_X1 U931 ( .A1(n1063), .A2(n1074), .A3(n1241), .ZN(n1198) );
AND3_X1 U932 ( .A1(n1201), .A2(n1234), .A3(n1251), .ZN(n1241) );
NOR2_X1 U933 ( .A1(n1083), .A2(n1246), .ZN(n1074) );
INV_X1 U934 ( .A(n1207), .ZN(n1063) );
NAND2_X1 U935 ( .A1(n1248), .A2(n1213), .ZN(n1207) );
INV_X1 U936 ( .A(n1247), .ZN(n1213) );
XOR2_X1 U937 ( .A(n1252), .B(G110), .Z(G12) );
NAND2_X1 U938 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NAND2_X1 U939 ( .A1(n1197), .A2(n1255), .ZN(n1254) );
INV_X1 U940 ( .A(KEYINPUT43), .ZN(n1255) );
AND2_X1 U941 ( .A1(n1256), .A2(n1038), .ZN(n1197) );
INV_X1 U942 ( .A(n1053), .ZN(n1038) );
NAND3_X1 U943 ( .A1(n1256), .A2(n1053), .A3(KEYINPUT43), .ZN(n1253) );
NAND2_X1 U944 ( .A1(n1234), .A2(n1056), .ZN(n1053) );
INV_X1 U945 ( .A(n1251), .ZN(n1056) );
XOR2_X1 U946 ( .A(n1257), .B(G469), .Z(n1251) );
NAND2_X1 U947 ( .A1(n1258), .A2(n1179), .ZN(n1257) );
XOR2_X1 U948 ( .A(n1259), .B(n1167), .Z(n1258) );
XOR2_X1 U949 ( .A(n1158), .B(n1260), .Z(n1167) );
XOR2_X1 U950 ( .A(n1261), .B(n1262), .Z(n1260) );
NOR2_X1 U951 ( .A1(G953), .A2(n1116), .ZN(n1262) );
INV_X1 U952 ( .A(G227), .ZN(n1116) );
XNOR2_X1 U953 ( .A(n1263), .B(n1264), .ZN(n1259) );
NOR2_X1 U954 ( .A1(G140), .A2(KEYINPUT27), .ZN(n1264) );
NOR2_X1 U955 ( .A1(KEYINPUT14), .A2(n1265), .ZN(n1263) );
XOR2_X1 U956 ( .A(n1166), .B(n1107), .Z(n1265) );
NAND2_X1 U957 ( .A1(n1266), .A2(n1267), .ZN(n1166) );
NAND2_X1 U958 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XOR2_X1 U959 ( .A(KEYINPUT58), .B(n1270), .Z(n1268) );
NAND2_X1 U960 ( .A1(n1270), .A2(G107), .ZN(n1266) );
INV_X1 U961 ( .A(n1061), .ZN(n1234) );
XOR2_X1 U962 ( .A(n1059), .B(KEYINPUT18), .Z(n1061) );
NAND2_X1 U963 ( .A1(G221), .A2(n1271), .ZN(n1059) );
AND3_X1 U964 ( .A1(n1075), .A2(n1201), .A3(n1222), .ZN(n1256) );
INV_X1 U965 ( .A(n1054), .ZN(n1222) );
NAND2_X1 U966 ( .A1(n1248), .A2(n1247), .ZN(n1054) );
NOR2_X1 U967 ( .A1(n1272), .A2(n1095), .ZN(n1247) );
NOR2_X1 U968 ( .A1(n1092), .A2(G475), .ZN(n1095) );
AND2_X1 U969 ( .A1(G475), .A2(n1092), .ZN(n1272) );
NAND2_X1 U970 ( .A1(n1151), .A2(n1179), .ZN(n1092) );
XOR2_X1 U971 ( .A(n1273), .B(n1274), .Z(n1151) );
XOR2_X1 U972 ( .A(n1275), .B(n1276), .Z(n1274) );
XOR2_X1 U973 ( .A(G131), .B(G104), .Z(n1276) );
XOR2_X1 U974 ( .A(G146), .B(G140), .Z(n1275) );
XOR2_X1 U975 ( .A(n1277), .B(n1278), .Z(n1273) );
XOR2_X1 U976 ( .A(n1279), .B(n1280), .Z(n1278) );
NAND2_X1 U977 ( .A1(KEYINPUT25), .A2(n1208), .ZN(n1280) );
NAND2_X1 U978 ( .A1(n1281), .A2(G214), .ZN(n1279) );
XNOR2_X1 U979 ( .A(n1282), .B(n1283), .ZN(n1277) );
NOR2_X1 U980 ( .A1(G125), .A2(KEYINPUT11), .ZN(n1283) );
NOR2_X1 U981 ( .A1(KEYINPUT57), .A2(n1284), .ZN(n1282) );
XOR2_X1 U982 ( .A(G122), .B(G113), .Z(n1284) );
NOR2_X1 U983 ( .A1(n1285), .A2(n1093), .ZN(n1248) );
NOR3_X1 U984 ( .A1(G478), .A2(G902), .A3(n1140), .ZN(n1093) );
XNOR2_X1 U985 ( .A(KEYINPUT21), .B(n1094), .ZN(n1285) );
AND2_X1 U986 ( .A1(G478), .A2(n1286), .ZN(n1094) );
NAND2_X1 U987 ( .A1(n1287), .A2(n1179), .ZN(n1286) );
INV_X1 U988 ( .A(n1140), .ZN(n1287) );
XOR2_X1 U989 ( .A(n1288), .B(n1289), .Z(n1140) );
NOR3_X1 U990 ( .A1(n1290), .A2(KEYINPUT55), .A3(n1291), .ZN(n1289) );
NOR2_X1 U991 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NOR2_X1 U992 ( .A1(n1294), .A2(n1295), .ZN(n1292) );
INV_X1 U993 ( .A(KEYINPUT56), .ZN(n1295) );
NOR2_X1 U994 ( .A1(KEYINPUT34), .A2(n1296), .ZN(n1294) );
NOR2_X1 U995 ( .A1(n1297), .A2(n1298), .ZN(n1290) );
INV_X1 U996 ( .A(n1296), .ZN(n1298) );
NAND2_X1 U997 ( .A1(n1299), .A2(n1300), .ZN(n1296) );
NAND2_X1 U998 ( .A1(G107), .A2(n1301), .ZN(n1300) );
XOR2_X1 U999 ( .A(n1302), .B(KEYINPUT46), .Z(n1299) );
OR2_X1 U1000 ( .A1(n1301), .A2(G107), .ZN(n1302) );
XOR2_X1 U1001 ( .A(G116), .B(G122), .Z(n1301) );
NOR2_X1 U1002 ( .A1(KEYINPUT34), .A2(n1303), .ZN(n1297) );
AND2_X1 U1003 ( .A1(KEYINPUT56), .A2(n1293), .ZN(n1303) );
XOR2_X1 U1004 ( .A(n1304), .B(n1305), .Z(n1293) );
XOR2_X1 U1005 ( .A(G143), .B(n1306), .Z(n1305) );
NOR2_X1 U1006 ( .A1(G128), .A2(KEYINPUT20), .ZN(n1306) );
NAND2_X1 U1007 ( .A1(KEYINPUT50), .A2(n1307), .ZN(n1304) );
INV_X1 U1008 ( .A(G134), .ZN(n1307) );
NAND3_X1 U1009 ( .A1(G234), .A2(n1308), .A3(G217), .ZN(n1288) );
XOR2_X1 U1010 ( .A(KEYINPUT60), .B(G953), .Z(n1308) );
AND2_X1 U1011 ( .A1(n1070), .A2(n1309), .ZN(n1201) );
NAND2_X1 U1012 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NAND2_X1 U1013 ( .A1(n1239), .A2(n1312), .ZN(n1311) );
INV_X1 U1014 ( .A(G898), .ZN(n1312) );
NOR3_X1 U1015 ( .A1(n1113), .A2(n1045), .A3(n1179), .ZN(n1239) );
AND2_X1 U1016 ( .A1(G234), .A2(G237), .ZN(n1045) );
XNOR2_X1 U1017 ( .A(n1115), .B(KEYINPUT54), .ZN(n1113) );
XOR2_X1 U1018 ( .A(n1238), .B(KEYINPUT1), .Z(n1310) );
NAND3_X1 U1019 ( .A1(n1313), .A2(n1115), .A3(n1314), .ZN(n1238) );
XNOR2_X1 U1020 ( .A(G952), .B(KEYINPUT62), .ZN(n1314) );
NAND2_X1 U1021 ( .A1(G237), .A2(G234), .ZN(n1313) );
AND2_X1 U1022 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U1023 ( .A1(G214), .A2(n1315), .ZN(n1072) );
XNOR2_X1 U1024 ( .A(n1084), .B(n1086), .ZN(n1071) );
AND2_X1 U1025 ( .A1(G210), .A2(n1315), .ZN(n1086) );
NAND2_X1 U1026 ( .A1(n1316), .A2(n1179), .ZN(n1315) );
INV_X1 U1027 ( .A(G237), .ZN(n1316) );
NAND2_X1 U1028 ( .A1(n1317), .A2(n1179), .ZN(n1084) );
XNOR2_X1 U1029 ( .A(n1174), .B(n1178), .ZN(n1317) );
AND2_X1 U1030 ( .A1(G224), .A2(n1115), .ZN(n1178) );
XNOR2_X1 U1031 ( .A(n1318), .B(n1319), .ZN(n1174) );
XOR2_X1 U1032 ( .A(n1107), .B(n1127), .Z(n1319) );
XNOR2_X1 U1033 ( .A(n1320), .B(G122), .ZN(n1127) );
NAND2_X1 U1034 ( .A1(KEYINPUT16), .A2(n1261), .ZN(n1320) );
INV_X1 U1035 ( .A(G110), .ZN(n1261) );
INV_X1 U1036 ( .A(n1321), .ZN(n1107) );
XOR2_X1 U1037 ( .A(n1322), .B(n1323), .Z(n1318) );
NOR2_X1 U1038 ( .A1(KEYINPUT6), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1039 ( .A(n1128), .B(n1325), .Z(n1324) );
NOR2_X1 U1040 ( .A1(KEYINPUT31), .A2(n1126), .ZN(n1325) );
XOR2_X1 U1041 ( .A(n1269), .B(n1270), .Z(n1126) );
XOR2_X1 U1042 ( .A(G101), .B(G104), .Z(n1270) );
INV_X1 U1043 ( .A(G107), .ZN(n1269) );
XOR2_X1 U1044 ( .A(n1326), .B(n1327), .Z(n1128) );
XOR2_X1 U1045 ( .A(G119), .B(G116), .Z(n1327) );
NAND2_X1 U1046 ( .A1(KEYINPUT2), .A2(n1328), .ZN(n1326) );
XOR2_X1 U1047 ( .A(n1233), .B(KEYINPUT30), .Z(n1322) );
INV_X1 U1048 ( .A(n1236), .ZN(n1075) );
NAND2_X1 U1049 ( .A1(n1246), .A2(n1329), .ZN(n1236) );
XOR2_X1 U1050 ( .A(KEYINPUT8), .B(n1083), .Z(n1329) );
XNOR2_X1 U1051 ( .A(n1330), .B(n1138), .ZN(n1083) );
AND2_X1 U1052 ( .A1(G217), .A2(n1271), .ZN(n1138) );
NAND2_X1 U1053 ( .A1(G234), .A2(n1179), .ZN(n1271) );
NAND2_X1 U1054 ( .A1(n1136), .A2(n1179), .ZN(n1330) );
XNOR2_X1 U1055 ( .A(n1331), .B(n1332), .ZN(n1136) );
XOR2_X1 U1056 ( .A(n1333), .B(n1334), .Z(n1332) );
XOR2_X1 U1057 ( .A(n1335), .B(G119), .Z(n1334) );
NAND3_X1 U1058 ( .A1(G234), .A2(n1115), .A3(G221), .ZN(n1335) );
INV_X1 U1059 ( .A(G953), .ZN(n1115) );
XOR2_X1 U1060 ( .A(n1221), .B(KEYINPUT3), .Z(n1333) );
XNOR2_X1 U1061 ( .A(n1108), .B(n1336), .ZN(n1331) );
XOR2_X1 U1062 ( .A(n1337), .B(n1338), .Z(n1336) );
NOR2_X1 U1063 ( .A1(G110), .A2(KEYINPUT15), .ZN(n1337) );
XOR2_X1 U1064 ( .A(n1233), .B(n1172), .Z(n1108) );
INV_X1 U1065 ( .A(G140), .ZN(n1172) );
INV_X1 U1066 ( .A(G125), .ZN(n1233) );
XOR2_X1 U1067 ( .A(n1091), .B(G472), .Z(n1246) );
NAND2_X1 U1068 ( .A1(n1339), .A2(n1179), .ZN(n1091) );
INV_X1 U1069 ( .A(G902), .ZN(n1179) );
XOR2_X1 U1070 ( .A(n1340), .B(n1341), .Z(n1339) );
XNOR2_X1 U1071 ( .A(n1342), .B(n1343), .ZN(n1341) );
NOR2_X1 U1072 ( .A1(KEYINPUT24), .A2(n1321), .ZN(n1343) );
XOR2_X1 U1073 ( .A(n1344), .B(n1338), .Z(n1321) );
XOR2_X1 U1074 ( .A(G128), .B(G146), .Z(n1338) );
XOR2_X1 U1075 ( .A(n1208), .B(KEYINPUT36), .Z(n1344) );
INV_X1 U1076 ( .A(G143), .ZN(n1208) );
NAND2_X1 U1077 ( .A1(KEYINPUT40), .A2(n1162), .ZN(n1342) );
XOR2_X1 U1078 ( .A(n1345), .B(G101), .Z(n1162) );
NAND2_X1 U1079 ( .A1(n1281), .A2(G210), .ZN(n1345) );
NOR2_X1 U1080 ( .A1(G953), .A2(G237), .ZN(n1281) );
XOR2_X1 U1081 ( .A(n1158), .B(n1157), .Z(n1340) );
XOR2_X1 U1082 ( .A(n1328), .B(n1346), .Z(n1157) );
XOR2_X1 U1083 ( .A(G116), .B(n1347), .Z(n1346) );
NOR2_X1 U1084 ( .A1(G119), .A2(KEYINPUT26), .ZN(n1347) );
XNOR2_X1 U1085 ( .A(n1250), .B(KEYINPUT10), .ZN(n1328) );
INV_X1 U1086 ( .A(G113), .ZN(n1250) );
XOR2_X1 U1087 ( .A(n1348), .B(n1112), .Z(n1158) );
XOR2_X1 U1088 ( .A(G131), .B(G134), .Z(n1112) );
NAND2_X1 U1089 ( .A1(KEYINPUT41), .A2(n1221), .ZN(n1348) );
INV_X1 U1090 ( .A(G137), .ZN(n1221) );
endmodule


