//Key = 0000100000001100111011010110101010000010111001101110111000111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322;

XNOR2_X1 U718 ( .A(G107), .B(n998), .ZN(G9) );
NOR2_X1 U719 ( .A1(n999), .A2(n1000), .ZN(G75) );
NOR4_X1 U720 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n1000) );
NAND4_X1 U721 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1001) );
NAND3_X1 U722 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1006) );
OR2_X1 U723 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NAND3_X1 U724 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1005) );
NAND2_X1 U725 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NAND3_X1 U726 ( .A1(n1019), .A2(n1020), .A3(n1009), .ZN(n1018) );
NAND3_X1 U727 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NAND4_X1 U728 ( .A1(KEYINPUT39), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1022) );
NAND3_X1 U729 ( .A1(n1027), .A2(n1028), .A3(KEYINPUT36), .ZN(n1021) );
NAND3_X1 U730 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1019) );
NAND2_X1 U731 ( .A1(n1028), .A2(n1032), .ZN(n1030) );
NAND2_X1 U732 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
OR2_X1 U733 ( .A1(n1035), .A2(KEYINPUT36), .ZN(n1034) );
NAND3_X1 U734 ( .A1(n1036), .A2(n1037), .A3(n1024), .ZN(n1029) );
NAND2_X1 U735 ( .A1(n1026), .A2(n1038), .ZN(n1037) );
NAND2_X1 U736 ( .A1(n1025), .A2(n1039), .ZN(n1038) );
INV_X1 U737 ( .A(KEYINPUT39), .ZN(n1039) );
XNOR2_X1 U738 ( .A(n1040), .B(KEYINPUT43), .ZN(n1025) );
NAND2_X1 U739 ( .A1(n1041), .A2(n1042), .ZN(n1036) );
NAND2_X1 U740 ( .A1(n1011), .A2(n1043), .ZN(n1017) );
NAND3_X1 U741 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
OR3_X1 U742 ( .A1(n1047), .A2(n1048), .A3(KEYINPUT57), .ZN(n1045) );
NAND2_X1 U743 ( .A1(KEYINPUT57), .A2(n1009), .ZN(n1044) );
AND3_X1 U744 ( .A1(n1024), .A2(n1028), .A3(n1031), .ZN(n1011) );
INV_X1 U745 ( .A(n1023), .ZN(n1031) );
NOR3_X1 U746 ( .A1(n1049), .A2(G953), .A3(G952), .ZN(n999) );
INV_X1 U747 ( .A(n1007), .ZN(n1049) );
NAND4_X1 U748 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1007) );
NOR4_X1 U749 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1053) );
XNOR2_X1 U750 ( .A(n1058), .B(n1059), .ZN(n1057) );
XOR2_X1 U751 ( .A(KEYINPUT22), .B(n1060), .Z(n1056) );
AND2_X1 U752 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
XOR2_X1 U753 ( .A(n1063), .B(n1064), .Z(n1055) );
XNOR2_X1 U754 ( .A(G472), .B(KEYINPUT21), .ZN(n1064) );
NAND2_X1 U755 ( .A1(KEYINPUT28), .A2(n1065), .ZN(n1063) );
NOR2_X1 U756 ( .A1(n1041), .A2(n1066), .ZN(n1052) );
NOR2_X1 U757 ( .A1(n1062), .A2(n1061), .ZN(n1066) );
XOR2_X1 U758 ( .A(KEYINPUT38), .B(n1067), .Z(n1051) );
XOR2_X1 U759 ( .A(n1068), .B(n1069), .Z(G72) );
NOR2_X1 U760 ( .A1(n1070), .A2(n1008), .ZN(n1069) );
NOR2_X1 U761 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XNOR2_X1 U762 ( .A(G227), .B(KEYINPUT51), .ZN(n1071) );
NAND2_X1 U763 ( .A1(n1073), .A2(n1074), .ZN(n1068) );
NAND2_X1 U764 ( .A1(n1075), .A2(n1008), .ZN(n1074) );
XOR2_X1 U765 ( .A(n1076), .B(n1077), .Z(n1075) );
NAND2_X1 U766 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
INV_X1 U767 ( .A(n1002), .ZN(n1078) );
NAND3_X1 U768 ( .A1(G900), .A2(n1077), .A3(G953), .ZN(n1073) );
XOR2_X1 U769 ( .A(n1080), .B(n1081), .Z(n1077) );
XNOR2_X1 U770 ( .A(n1082), .B(n1083), .ZN(n1081) );
NOR2_X1 U771 ( .A1(KEYINPUT35), .A2(n1084), .ZN(n1083) );
XOR2_X1 U772 ( .A(n1085), .B(n1086), .Z(n1084) );
XOR2_X1 U773 ( .A(n1087), .B(n1088), .Z(n1086) );
XNOR2_X1 U774 ( .A(G131), .B(KEYINPUT42), .ZN(n1085) );
NAND2_X1 U775 ( .A1(n1089), .A2(KEYINPUT60), .ZN(n1080) );
XNOR2_X1 U776 ( .A(G125), .B(KEYINPUT15), .ZN(n1089) );
XOR2_X1 U777 ( .A(n1090), .B(n1091), .Z(G69) );
XOR2_X1 U778 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND2_X1 U779 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
INV_X1 U780 ( .A(n1096), .ZN(n1095) );
NAND2_X1 U781 ( .A1(G953), .A2(n1097), .ZN(n1092) );
NAND2_X1 U782 ( .A1(n1098), .A2(G224), .ZN(n1097) );
XNOR2_X1 U783 ( .A(G898), .B(KEYINPUT49), .ZN(n1098) );
AND2_X1 U784 ( .A1(n1004), .A2(n1008), .ZN(n1090) );
NOR2_X1 U785 ( .A1(n1099), .A2(n1100), .ZN(G66) );
XNOR2_X1 U786 ( .A(n1101), .B(n1102), .ZN(n1100) );
NOR2_X1 U787 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(G63) );
XNOR2_X1 U789 ( .A(n1099), .B(KEYINPUT45), .ZN(n1106) );
XOR2_X1 U790 ( .A(n1107), .B(n1108), .Z(n1105) );
XNOR2_X1 U791 ( .A(KEYINPUT25), .B(n1109), .ZN(n1108) );
NAND3_X1 U792 ( .A1(n1110), .A2(G478), .A3(KEYINPUT48), .ZN(n1107) );
NOR2_X1 U793 ( .A1(n1099), .A2(n1111), .ZN(G60) );
XOR2_X1 U794 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U795 ( .A1(KEYINPUT1), .A2(n1114), .ZN(n1113) );
AND2_X1 U796 ( .A1(G475), .A2(n1110), .ZN(n1112) );
XNOR2_X1 U797 ( .A(G104), .B(n1115), .ZN(G6) );
NOR2_X1 U798 ( .A1(n1099), .A2(n1116), .ZN(G57) );
XOR2_X1 U799 ( .A(n1117), .B(KEYINPUT52), .Z(n1116) );
NAND2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U801 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U802 ( .A(KEYINPUT59), .B(n1122), .Z(n1118) );
NOR2_X1 U803 ( .A1(n1120), .A2(n1121), .ZN(n1122) );
XNOR2_X1 U804 ( .A(G101), .B(n1123), .ZN(n1121) );
XOR2_X1 U805 ( .A(n1124), .B(n1125), .Z(n1120) );
NOR2_X1 U806 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U807 ( .A(KEYINPUT11), .B(n1128), .Z(n1127) );
NOR2_X1 U808 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U809 ( .A1(n1131), .A2(n1132), .ZN(n1126) );
XOR2_X1 U810 ( .A(n1133), .B(n1134), .Z(n1124) );
NOR2_X1 U811 ( .A1(n1135), .A2(n1104), .ZN(n1134) );
NOR2_X1 U812 ( .A1(n1099), .A2(n1136), .ZN(G54) );
XOR2_X1 U813 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR3_X1 U815 ( .A1(n1141), .A2(KEYINPUT37), .A3(n1142), .ZN(n1140) );
NOR2_X1 U816 ( .A1(n1143), .A2(n1144), .ZN(n1139) );
NOR2_X1 U817 ( .A1(KEYINPUT37), .A2(n1142), .ZN(n1143) );
XOR2_X1 U818 ( .A(n1145), .B(n1146), .Z(n1137) );
AND2_X1 U819 ( .A1(G469), .A2(n1110), .ZN(n1146) );
INV_X1 U820 ( .A(n1104), .ZN(n1110) );
NAND2_X1 U821 ( .A1(KEYINPUT23), .A2(n1147), .ZN(n1145) );
NOR2_X1 U822 ( .A1(n1008), .A2(G952), .ZN(n1099) );
NOR2_X1 U823 ( .A1(n1148), .A2(n1149), .ZN(G51) );
XOR2_X1 U824 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U825 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U826 ( .A1(n1061), .A2(n1104), .ZN(n1153) );
NAND2_X1 U827 ( .A1(G902), .A2(n1154), .ZN(n1104) );
OR3_X1 U828 ( .A1(n1004), .A2(n1003), .A3(n1002), .ZN(n1154) );
NAND3_X1 U829 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1002) );
NAND2_X1 U830 ( .A1(n1027), .A2(n1158), .ZN(n1157) );
NAND2_X1 U831 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U832 ( .A(n1079), .B(KEYINPUT24), .ZN(n1003) );
AND4_X1 U833 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1079) );
AND2_X1 U834 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NAND2_X1 U835 ( .A1(n1167), .A2(n1168), .ZN(n1162) );
OR3_X1 U836 ( .A1(n1160), .A2(n1169), .A3(n1168), .ZN(n1161) );
INV_X1 U837 ( .A(KEYINPUT33), .ZN(n1168) );
NAND4_X1 U838 ( .A1(n1170), .A2(n998), .A3(n1171), .A4(n1172), .ZN(n1004) );
NOR4_X1 U839 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1172) );
NOR3_X1 U840 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1171) );
AND4_X1 U841 ( .A1(KEYINPUT55), .A2(n1027), .A3(n1046), .A4(n1180), .ZN(n1179) );
NOR2_X1 U842 ( .A1(KEYINPUT55), .A2(n1115), .ZN(n1178) );
NAND3_X1 U843 ( .A1(n1181), .A2(n1180), .A3(n1027), .ZN(n1115) );
NAND3_X1 U844 ( .A1(n1169), .A2(n1180), .A3(n1181), .ZN(n998) );
NOR2_X1 U845 ( .A1(KEYINPUT14), .A2(n1182), .ZN(n1152) );
XOR2_X1 U846 ( .A(KEYINPUT16), .B(n1183), .Z(n1182) );
NOR2_X1 U847 ( .A1(G952), .A2(n1184), .ZN(n1148) );
XNOR2_X1 U848 ( .A(KEYINPUT61), .B(n1008), .ZN(n1184) );
XNOR2_X1 U849 ( .A(n1185), .B(n1186), .ZN(G48) );
NOR2_X1 U850 ( .A1(n1035), .A2(n1160), .ZN(n1186) );
XNOR2_X1 U851 ( .A(G143), .B(n1155), .ZN(G45) );
NAND3_X1 U852 ( .A1(n1187), .A2(n1181), .A3(n1188), .ZN(n1155) );
AND3_X1 U853 ( .A1(n1012), .A2(n1189), .A3(n1067), .ZN(n1188) );
XNOR2_X1 U854 ( .A(G140), .B(n1190), .ZN(G42) );
NAND2_X1 U855 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
INV_X1 U856 ( .A(n1159), .ZN(n1192) );
NAND2_X1 U857 ( .A1(n1013), .A2(n1193), .ZN(n1159) );
XNOR2_X1 U858 ( .A(n1027), .B(KEYINPUT4), .ZN(n1191) );
XOR2_X1 U859 ( .A(n1156), .B(n1194), .Z(G39) );
NAND2_X1 U860 ( .A1(KEYINPUT32), .A2(G137), .ZN(n1194) );
NAND3_X1 U861 ( .A1(n1193), .A2(n1195), .A3(n1024), .ZN(n1156) );
XNOR2_X1 U862 ( .A(G134), .B(n1166), .ZN(G36) );
NAND3_X1 U863 ( .A1(n1169), .A2(n1012), .A3(n1193), .ZN(n1166) );
AND3_X1 U864 ( .A1(n1181), .A2(n1196), .A3(n1028), .ZN(n1193) );
XOR2_X1 U865 ( .A(n1197), .B(G131), .Z(G33) );
NAND2_X1 U866 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
OR2_X1 U867 ( .A1(n1163), .A2(KEYINPUT8), .ZN(n1199) );
NAND2_X1 U868 ( .A1(n1200), .A2(n1028), .ZN(n1163) );
INV_X1 U869 ( .A(n1201), .ZN(n1200) );
NAND3_X1 U870 ( .A1(n1028), .A2(n1201), .A3(KEYINPUT8), .ZN(n1198) );
NAND4_X1 U871 ( .A1(n1027), .A2(n1181), .A3(n1012), .A4(n1196), .ZN(n1201) );
NOR2_X1 U872 ( .A1(n1042), .A2(n1041), .ZN(n1028) );
INV_X1 U873 ( .A(n1040), .ZN(n1041) );
XOR2_X1 U874 ( .A(n1202), .B(n1167), .Z(G30) );
NOR2_X1 U875 ( .A1(n1160), .A2(n1033), .ZN(n1167) );
INV_X1 U876 ( .A(n1169), .ZN(n1033) );
NAND3_X1 U877 ( .A1(n1195), .A2(n1181), .A3(n1187), .ZN(n1160) );
NAND2_X1 U878 ( .A1(KEYINPUT46), .A2(n1203), .ZN(n1202) );
XNOR2_X1 U879 ( .A(n1204), .B(n1176), .ZN(G3) );
AND2_X1 U880 ( .A1(n1205), .A2(n1012), .ZN(n1176) );
XNOR2_X1 U881 ( .A(G125), .B(n1165), .ZN(G27) );
NAND4_X1 U882 ( .A1(n1027), .A2(n1013), .A3(n1187), .A4(n1009), .ZN(n1165) );
AND3_X1 U883 ( .A1(n1196), .A2(n1040), .A3(n1042), .ZN(n1187) );
NAND2_X1 U884 ( .A1(n1023), .A2(n1206), .ZN(n1196) );
NAND4_X1 U885 ( .A1(G953), .A2(G902), .A3(n1207), .A4(n1072), .ZN(n1206) );
INV_X1 U886 ( .A(G900), .ZN(n1072) );
NAND2_X1 U887 ( .A1(n1208), .A2(n1209), .ZN(G24) );
NAND2_X1 U888 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XNOR2_X1 U889 ( .A(n1177), .B(KEYINPUT12), .ZN(n1210) );
INV_X1 U890 ( .A(n1212), .ZN(n1177) );
NAND2_X1 U891 ( .A1(n1213), .A2(G122), .ZN(n1208) );
XNOR2_X1 U892 ( .A(KEYINPUT13), .B(n1212), .ZN(n1213) );
NAND4_X1 U893 ( .A1(n1009), .A2(n1180), .A3(n1067), .A4(n1189), .ZN(n1212) );
AND3_X1 U894 ( .A1(n1016), .A2(n1014), .A3(n1214), .ZN(n1180) );
NAND2_X1 U895 ( .A1(n1215), .A2(n1216), .ZN(G21) );
NAND2_X1 U896 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XOR2_X1 U897 ( .A(n1170), .B(KEYINPUT26), .Z(n1217) );
NAND2_X1 U898 ( .A1(n1219), .A2(G119), .ZN(n1215) );
XNOR2_X1 U899 ( .A(KEYINPUT53), .B(n1170), .ZN(n1219) );
NAND4_X1 U900 ( .A1(n1024), .A2(n1195), .A3(n1009), .A4(n1214), .ZN(n1170) );
XOR2_X1 U901 ( .A(G116), .B(n1175), .Z(G18) );
AND2_X1 U902 ( .A1(n1220), .A2(n1169), .ZN(n1175) );
NOR2_X1 U903 ( .A1(n1067), .A2(n1050), .ZN(n1169) );
XOR2_X1 U904 ( .A(G113), .B(n1174), .Z(G15) );
AND2_X1 U905 ( .A1(n1220), .A2(n1027), .ZN(n1174) );
INV_X1 U906 ( .A(n1035), .ZN(n1027) );
NAND2_X1 U907 ( .A1(n1050), .A2(n1067), .ZN(n1035) );
INV_X1 U908 ( .A(n1189), .ZN(n1050) );
AND3_X1 U909 ( .A1(n1214), .A2(n1012), .A3(n1009), .ZN(n1220) );
INV_X1 U910 ( .A(n1054), .ZN(n1009) );
NAND2_X1 U911 ( .A1(n1221), .A2(n1047), .ZN(n1054) );
NAND2_X1 U912 ( .A1(n1222), .A2(n1223), .ZN(n1012) );
OR3_X1 U913 ( .A1(n1016), .A2(n1224), .A3(KEYINPUT62), .ZN(n1223) );
NAND2_X1 U914 ( .A1(KEYINPUT62), .A2(n1195), .ZN(n1222) );
NOR2_X1 U915 ( .A1(n1014), .A2(n1016), .ZN(n1195) );
XOR2_X1 U916 ( .A(G110), .B(n1173), .Z(G12) );
AND2_X1 U917 ( .A1(n1205), .A2(n1013), .ZN(n1173) );
AND2_X1 U918 ( .A1(n1224), .A2(n1016), .ZN(n1013) );
XNOR2_X1 U919 ( .A(n1065), .B(n1135), .ZN(n1016) );
INV_X1 U920 ( .A(G472), .ZN(n1135) );
NAND2_X1 U921 ( .A1(n1225), .A2(n1226), .ZN(n1065) );
XOR2_X1 U922 ( .A(n1227), .B(n1228), .Z(n1225) );
XOR2_X1 U923 ( .A(n1229), .B(n1230), .Z(n1228) );
NAND2_X1 U924 ( .A1(KEYINPUT40), .A2(n1231), .ZN(n1230) );
INV_X1 U925 ( .A(n1123), .ZN(n1231) );
NAND3_X1 U926 ( .A1(G210), .A2(n1008), .A3(n1232), .ZN(n1123) );
XNOR2_X1 U927 ( .A(G237), .B(KEYINPUT10), .ZN(n1232) );
NAND2_X1 U928 ( .A1(n1233), .A2(n1234), .ZN(n1229) );
NAND2_X1 U929 ( .A1(n1131), .A2(n1235), .ZN(n1234) );
NAND2_X1 U930 ( .A1(n1129), .A2(n1236), .ZN(n1235) );
NAND2_X1 U931 ( .A1(KEYINPUT5), .A2(n1237), .ZN(n1236) );
INV_X1 U932 ( .A(n1130), .ZN(n1131) );
NAND3_X1 U933 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1233) );
INV_X1 U934 ( .A(KEYINPUT5), .ZN(n1240) );
NAND2_X1 U935 ( .A1(n1132), .A2(n1237), .ZN(n1239) );
NAND2_X1 U936 ( .A1(n1129), .A2(n1241), .ZN(n1238) );
NAND2_X1 U937 ( .A1(n1130), .A2(n1237), .ZN(n1241) );
INV_X1 U938 ( .A(KEYINPUT3), .ZN(n1237) );
INV_X1 U939 ( .A(n1132), .ZN(n1129) );
XNOR2_X1 U940 ( .A(n1242), .B(KEYINPUT18), .ZN(n1132) );
XNOR2_X1 U941 ( .A(G101), .B(n1133), .ZN(n1227) );
NAND2_X1 U942 ( .A1(n1243), .A2(n1244), .ZN(n1133) );
NAND2_X1 U943 ( .A1(G113), .A2(n1245), .ZN(n1244) );
XOR2_X1 U944 ( .A(n1246), .B(KEYINPUT19), .Z(n1243) );
OR2_X1 U945 ( .A1(n1245), .A2(G113), .ZN(n1246) );
XOR2_X1 U946 ( .A(G116), .B(n1247), .Z(n1245) );
XNOR2_X1 U947 ( .A(KEYINPUT27), .B(n1218), .ZN(n1247) );
INV_X1 U948 ( .A(n1014), .ZN(n1224) );
XNOR2_X1 U949 ( .A(n1058), .B(n1248), .ZN(n1014) );
NOR2_X1 U950 ( .A1(n1059), .A2(KEYINPUT47), .ZN(n1248) );
INV_X1 U951 ( .A(n1103), .ZN(n1059) );
NAND2_X1 U952 ( .A1(G217), .A2(n1249), .ZN(n1103) );
NAND2_X1 U953 ( .A1(n1101), .A2(n1226), .ZN(n1058) );
XNOR2_X1 U954 ( .A(n1250), .B(n1251), .ZN(n1101) );
XNOR2_X1 U955 ( .A(G128), .B(n1252), .ZN(n1251) );
XNOR2_X1 U956 ( .A(KEYINPUT20), .B(KEYINPUT17), .ZN(n1252) );
XNOR2_X1 U957 ( .A(n1253), .B(n1254), .ZN(n1250) );
XOR2_X1 U958 ( .A(n1255), .B(n1256), .Z(n1254) );
NAND2_X1 U959 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND4_X1 U960 ( .A1(G137), .A2(G221), .A3(G234), .A4(n1008), .ZN(n1258) );
XOR2_X1 U961 ( .A(n1259), .B(KEYINPUT0), .Z(n1257) );
NAND2_X1 U962 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND3_X1 U963 ( .A1(G234), .A2(n1008), .A3(G221), .ZN(n1261) );
NAND3_X1 U964 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1255) );
INV_X1 U965 ( .A(n1265), .ZN(n1264) );
OR2_X1 U966 ( .A1(n1266), .A2(n1185), .ZN(n1263) );
NAND3_X1 U967 ( .A1(n1266), .A2(n1267), .A3(n1185), .ZN(n1262) );
XOR2_X1 U968 ( .A(n1268), .B(KEYINPUT50), .Z(n1266) );
AND3_X1 U969 ( .A1(n1181), .A2(n1214), .A3(n1024), .ZN(n1205) );
NOR2_X1 U970 ( .A1(n1189), .A2(n1067), .ZN(n1024) );
XNOR2_X1 U971 ( .A(n1269), .B(G475), .ZN(n1067) );
NAND2_X1 U972 ( .A1(n1114), .A2(n1226), .ZN(n1269) );
XOR2_X1 U973 ( .A(n1270), .B(n1271), .Z(n1114) );
XNOR2_X1 U974 ( .A(n1211), .B(G113), .ZN(n1271) );
XOR2_X1 U975 ( .A(n1272), .B(n1273), .Z(n1270) );
NOR2_X1 U976 ( .A1(KEYINPUT44), .A2(n1274), .ZN(n1273) );
XOR2_X1 U977 ( .A(n1275), .B(n1276), .Z(n1274) );
NOR3_X1 U978 ( .A1(n1265), .A2(n1277), .A3(n1278), .ZN(n1276) );
NOR2_X1 U979 ( .A1(n1185), .A2(n1279), .ZN(n1278) );
INV_X1 U980 ( .A(n1268), .ZN(n1279) );
NOR3_X1 U981 ( .A1(G146), .A2(n1280), .A3(n1268), .ZN(n1277) );
NOR2_X1 U982 ( .A1(n1281), .A2(G140), .ZN(n1268) );
INV_X1 U983 ( .A(G125), .ZN(n1281) );
NOR2_X1 U984 ( .A1(n1185), .A2(n1267), .ZN(n1265) );
INV_X1 U985 ( .A(n1280), .ZN(n1267) );
NOR2_X1 U986 ( .A1(n1082), .A2(G125), .ZN(n1280) );
INV_X1 U987 ( .A(G140), .ZN(n1082) );
XNOR2_X1 U988 ( .A(G131), .B(n1282), .ZN(n1275) );
NOR2_X1 U989 ( .A1(KEYINPUT56), .A2(n1283), .ZN(n1282) );
XOR2_X1 U990 ( .A(G143), .B(n1284), .Z(n1283) );
AND3_X1 U991 ( .A1(G214), .A2(n1008), .A3(n1285), .ZN(n1284) );
XNOR2_X1 U992 ( .A(n1286), .B(G478), .ZN(n1189) );
NAND2_X1 U993 ( .A1(n1226), .A2(n1109), .ZN(n1286) );
NAND2_X1 U994 ( .A1(n1287), .A2(n1288), .ZN(n1109) );
NAND2_X1 U995 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XOR2_X1 U996 ( .A(n1291), .B(KEYINPUT9), .Z(n1287) );
OR2_X1 U997 ( .A1(n1290), .A2(n1289), .ZN(n1291) );
XNOR2_X1 U998 ( .A(n1292), .B(n1293), .ZN(n1289) );
XOR2_X1 U999 ( .A(KEYINPUT6), .B(G134), .Z(n1293) );
XNOR2_X1 U1000 ( .A(n1294), .B(n1295), .ZN(n1292) );
NAND3_X1 U1001 ( .A1(G234), .A2(n1008), .A3(G217), .ZN(n1290) );
AND3_X1 U1002 ( .A1(n1296), .A2(n1040), .A3(n1042), .ZN(n1214) );
INV_X1 U1003 ( .A(n1026), .ZN(n1042) );
XOR2_X1 U1004 ( .A(n1297), .B(n1061), .Z(n1026) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1298), .ZN(n1061) );
XNOR2_X1 U1006 ( .A(n1062), .B(KEYINPUT58), .ZN(n1297) );
AND2_X1 U1007 ( .A1(n1299), .A2(n1226), .ZN(n1062) );
XNOR2_X1 U1008 ( .A(n1150), .B(n1183), .ZN(n1299) );
XNOR2_X1 U1009 ( .A(n1242), .B(G125), .ZN(n1183) );
XNOR2_X1 U1010 ( .A(G146), .B(n1295), .ZN(n1242) );
XNOR2_X1 U1011 ( .A(n1203), .B(G143), .ZN(n1295) );
INV_X1 U1012 ( .A(G128), .ZN(n1203) );
XOR2_X1 U1013 ( .A(n1094), .B(n1300), .Z(n1150) );
AND2_X1 U1014 ( .A1(n1008), .A2(G224), .ZN(n1300) );
XNOR2_X1 U1015 ( .A(n1301), .B(n1302), .ZN(n1094) );
XNOR2_X1 U1016 ( .A(n1204), .B(n1303), .ZN(n1302) );
XOR2_X1 U1017 ( .A(KEYINPUT29), .B(G113), .Z(n1303) );
INV_X1 U1018 ( .A(G101), .ZN(n1204) );
XOR2_X1 U1019 ( .A(n1304), .B(n1294), .Z(n1301) );
XOR2_X1 U1020 ( .A(G107), .B(n1305), .Z(n1294) );
XNOR2_X1 U1021 ( .A(n1211), .B(G116), .ZN(n1305) );
INV_X1 U1022 ( .A(G122), .ZN(n1211) );
XOR2_X1 U1023 ( .A(n1306), .B(n1253), .Z(n1304) );
XNOR2_X1 U1024 ( .A(G110), .B(n1218), .ZN(n1253) );
INV_X1 U1025 ( .A(G119), .ZN(n1218) );
NAND2_X1 U1026 ( .A1(KEYINPUT54), .A2(n1272), .ZN(n1306) );
NAND2_X1 U1027 ( .A1(G214), .A2(n1298), .ZN(n1040) );
NAND2_X1 U1028 ( .A1(n1285), .A2(n1307), .ZN(n1298) );
INV_X1 U1029 ( .A(G237), .ZN(n1285) );
NAND2_X1 U1030 ( .A1(n1023), .A2(n1308), .ZN(n1296) );
NAND3_X1 U1031 ( .A1(G902), .A2(n1207), .A3(n1096), .ZN(n1308) );
NOR2_X1 U1032 ( .A1(n1008), .A2(G898), .ZN(n1096) );
NAND3_X1 U1033 ( .A1(n1207), .A2(n1008), .A3(G952), .ZN(n1023) );
NAND2_X1 U1034 ( .A1(G237), .A2(G234), .ZN(n1207) );
INV_X1 U1035 ( .A(n1046), .ZN(n1181) );
NAND2_X1 U1036 ( .A1(n1048), .A2(n1047), .ZN(n1046) );
NAND2_X1 U1037 ( .A1(G221), .A2(n1249), .ZN(n1047) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1307), .ZN(n1249) );
INV_X1 U1039 ( .A(n1221), .ZN(n1048) );
XOR2_X1 U1040 ( .A(n1309), .B(G469), .Z(n1221) );
NAND2_X1 U1041 ( .A1(n1310), .A2(n1226), .ZN(n1309) );
XNOR2_X1 U1042 ( .A(n1307), .B(KEYINPUT41), .ZN(n1226) );
INV_X1 U1043 ( .A(G902), .ZN(n1307) );
XOR2_X1 U1044 ( .A(n1142), .B(n1311), .Z(n1310) );
XNOR2_X1 U1045 ( .A(n1141), .B(n1312), .ZN(n1311) );
NOR2_X1 U1046 ( .A1(KEYINPUT7), .A2(n1147), .ZN(n1312) );
XNOR2_X1 U1047 ( .A(n1313), .B(n1314), .ZN(n1147) );
XNOR2_X1 U1048 ( .A(G101), .B(n1315), .ZN(n1314) );
NAND2_X1 U1049 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
NAND2_X1 U1050 ( .A1(G107), .A2(n1272), .ZN(n1317) );
XOR2_X1 U1051 ( .A(n1318), .B(KEYINPUT34), .Z(n1316) );
OR2_X1 U1052 ( .A1(n1272), .A2(G107), .ZN(n1318) );
XNOR2_X1 U1053 ( .A(G104), .B(KEYINPUT2), .ZN(n1272) );
XNOR2_X1 U1054 ( .A(n1130), .B(n1088), .ZN(n1313) );
XNOR2_X1 U1055 ( .A(n1319), .B(n1320), .ZN(n1088) );
XOR2_X1 U1056 ( .A(G143), .B(n1321), .Z(n1320) );
NOR2_X1 U1057 ( .A1(G128), .A2(KEYINPUT31), .ZN(n1321) );
NAND2_X1 U1058 ( .A1(KEYINPUT30), .A2(n1185), .ZN(n1319) );
INV_X1 U1059 ( .A(G146), .ZN(n1185) );
XNOR2_X1 U1060 ( .A(n1322), .B(n1087), .ZN(n1130) );
XNOR2_X1 U1061 ( .A(G134), .B(n1260), .ZN(n1087) );
INV_X1 U1062 ( .A(G137), .ZN(n1260) );
NAND2_X1 U1063 ( .A1(KEYINPUT63), .A2(G131), .ZN(n1322) );
INV_X1 U1064 ( .A(n1144), .ZN(n1141) );
NAND2_X1 U1065 ( .A1(G227), .A2(n1008), .ZN(n1144) );
INV_X1 U1066 ( .A(G953), .ZN(n1008) );
XNOR2_X1 U1067 ( .A(G110), .B(G140), .ZN(n1142) );
endmodule


