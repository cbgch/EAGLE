//Key = 1001000010100111111011100101011010011101100100000101101100010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343;

XNOR2_X1 U740 ( .A(G107), .B(n1025), .ZN(G9) );
NOR2_X1 U741 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR3_X1 U742 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
XOR2_X1 U743 ( .A(KEYINPUT4), .B(n1031), .Z(n1030) );
NOR3_X1 U744 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NAND3_X1 U745 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1032) );
NAND3_X1 U746 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1028) );
NAND2_X1 U747 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U748 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND3_X1 U749 ( .A1(n1036), .A2(n1045), .A3(n1046), .ZN(n1044) );
NAND2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND2_X1 U751 ( .A1(n1037), .A2(n1049), .ZN(n1048) );
NAND2_X1 U752 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U753 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
INV_X1 U754 ( .A(n1054), .ZN(n1050) );
NAND2_X1 U755 ( .A1(n1035), .A2(n1055), .ZN(n1047) );
NAND2_X1 U756 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U757 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND3_X1 U758 ( .A1(n1060), .A2(n1061), .A3(n1037), .ZN(n1043) );
NAND2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
OR2_X1 U760 ( .A1(n1064), .A2(KEYINPUT43), .ZN(n1062) );
NAND4_X1 U761 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1035), .ZN(n1060) );
NAND2_X1 U762 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U763 ( .A1(KEYINPUT43), .A2(n1070), .ZN(n1066) );
NAND2_X1 U764 ( .A1(n1071), .A2(n1036), .ZN(n1065) );
INV_X1 U765 ( .A(n1034), .ZN(n1041) );
NOR3_X1 U766 ( .A1(n1072), .A2(G953), .A3(G952), .ZN(n1026) );
INV_X1 U767 ( .A(n1038), .ZN(n1072) );
NAND4_X1 U768 ( .A1(n1037), .A2(n1035), .A3(n1073), .A4(n1074), .ZN(n1038) );
NOR3_X1 U769 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1074) );
XOR2_X1 U770 ( .A(n1078), .B(KEYINPUT54), .Z(n1076) );
XOR2_X1 U771 ( .A(n1079), .B(n1080), .Z(n1073) );
XOR2_X1 U772 ( .A(KEYINPUT21), .B(n1081), .Z(n1080) );
NAND2_X1 U773 ( .A1(KEYINPUT18), .A2(n1082), .ZN(n1079) );
XOR2_X1 U774 ( .A(n1083), .B(n1084), .Z(G72) );
XOR2_X1 U775 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U776 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XNOR2_X1 U777 ( .A(KEYINPUT57), .B(n1039), .ZN(n1088) );
INV_X1 U778 ( .A(n1089), .ZN(n1087) );
NAND2_X1 U779 ( .A1(n1090), .A2(n1091), .ZN(n1085) );
INV_X1 U780 ( .A(n1092), .ZN(n1091) );
XOR2_X1 U781 ( .A(n1093), .B(n1094), .Z(n1090) );
XOR2_X1 U782 ( .A(n1095), .B(n1096), .Z(n1094) );
XNOR2_X1 U783 ( .A(n1097), .B(n1098), .ZN(n1093) );
XNOR2_X1 U784 ( .A(n1099), .B(KEYINPUT62), .ZN(n1098) );
NAND2_X1 U785 ( .A1(KEYINPUT52), .A2(n1100), .ZN(n1099) );
XNOR2_X1 U786 ( .A(G134), .B(n1101), .ZN(n1100) );
NAND2_X1 U787 ( .A1(KEYINPUT32), .A2(G137), .ZN(n1101) );
NAND2_X1 U788 ( .A1(G953), .A2(n1102), .ZN(n1083) );
NAND2_X1 U789 ( .A1(G900), .A2(G227), .ZN(n1102) );
XOR2_X1 U790 ( .A(n1103), .B(n1104), .Z(G69) );
XOR2_X1 U791 ( .A(n1105), .B(n1106), .Z(n1104) );
NAND2_X1 U792 ( .A1(G953), .A2(n1107), .ZN(n1106) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1107) );
NAND2_X1 U794 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
NAND2_X1 U795 ( .A1(G953), .A2(n1110), .ZN(n1109) );
XOR2_X1 U796 ( .A(n1111), .B(n1112), .Z(n1108) );
NAND2_X1 U797 ( .A1(KEYINPUT10), .A2(n1113), .ZN(n1111) );
NOR2_X1 U798 ( .A1(n1114), .A2(G953), .ZN(n1103) );
NOR3_X1 U799 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
NOR2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XNOR2_X1 U801 ( .A(n1120), .B(n1121), .ZN(n1119) );
NOR2_X1 U802 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U803 ( .A1(n1118), .A2(n1124), .ZN(G63) );
NOR2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XOR2_X1 U805 ( .A(n1127), .B(KEYINPUT16), .Z(n1126) );
NAND2_X1 U806 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR2_X1 U807 ( .A1(n1128), .A2(n1129), .ZN(n1125) );
NAND3_X1 U808 ( .A1(G478), .A2(n1130), .A3(G902), .ZN(n1129) );
XNOR2_X1 U809 ( .A(KEYINPUT51), .B(n1029), .ZN(n1130) );
NOR2_X1 U810 ( .A1(n1118), .A2(n1131), .ZN(G60) );
XOR2_X1 U811 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U812 ( .A1(KEYINPUT8), .A2(n1134), .ZN(n1133) );
NAND3_X1 U813 ( .A1(G475), .A2(n1029), .A3(n1135), .ZN(n1132) );
XNOR2_X1 U814 ( .A(G902), .B(KEYINPUT40), .ZN(n1135) );
XOR2_X1 U815 ( .A(n1136), .B(n1137), .Z(G6) );
XNOR2_X1 U816 ( .A(G104), .B(KEYINPUT24), .ZN(n1137) );
NAND4_X1 U817 ( .A1(n1138), .A2(n1036), .A3(n1139), .A4(n1140), .ZN(n1136) );
OR2_X1 U818 ( .A1(n1141), .A2(KEYINPUT2), .ZN(n1140) );
NAND2_X1 U819 ( .A1(KEYINPUT2), .A2(n1142), .ZN(n1139) );
NAND2_X1 U820 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
INV_X1 U821 ( .A(n1145), .ZN(n1144) );
NOR2_X1 U822 ( .A1(n1118), .A2(n1146), .ZN(G57) );
XOR2_X1 U823 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U824 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U825 ( .A1(n1151), .A2(n1123), .ZN(n1150) );
XNOR2_X1 U826 ( .A(n1152), .B(n1153), .ZN(n1147) );
NOR2_X1 U827 ( .A1(KEYINPUT19), .A2(n1154), .ZN(n1153) );
NOR3_X1 U828 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(G54) );
AND2_X1 U829 ( .A1(KEYINPUT0), .A2(n1118), .ZN(n1157) );
NOR3_X1 U830 ( .A1(KEYINPUT0), .A2(G953), .A3(G952), .ZN(n1156) );
XNOR2_X1 U831 ( .A(n1158), .B(n1159), .ZN(n1155) );
XOR2_X1 U832 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U833 ( .A1(n1162), .A2(n1123), .ZN(n1161) );
NAND2_X1 U834 ( .A1(G902), .A2(n1029), .ZN(n1123) );
INV_X1 U835 ( .A(n1163), .ZN(n1029) );
NOR2_X1 U836 ( .A1(n1164), .A2(n1165), .ZN(n1160) );
NOR2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XNOR2_X1 U838 ( .A(n1168), .B(KEYINPUT27), .ZN(n1167) );
NOR2_X1 U839 ( .A1(n1118), .A2(n1169), .ZN(G51) );
XOR2_X1 U840 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND3_X1 U841 ( .A1(G902), .A2(G210), .A3(n1172), .ZN(n1171) );
XNOR2_X1 U842 ( .A(n1163), .B(KEYINPUT50), .ZN(n1172) );
NOR4_X1 U843 ( .A1(n1173), .A2(n1115), .A3(n1117), .A4(n1089), .ZN(n1163) );
NAND2_X1 U844 ( .A1(n1174), .A2(n1175), .ZN(n1089) );
AND4_X1 U845 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1175) );
AND4_X1 U846 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1174) );
NAND3_X1 U847 ( .A1(n1184), .A2(n1037), .A3(n1138), .ZN(n1183) );
NAND2_X1 U848 ( .A1(n1185), .A2(n1186), .ZN(n1117) );
NAND4_X1 U849 ( .A1(n1070), .A2(n1145), .A3(n1187), .A4(n1188), .ZN(n1186) );
XNOR2_X1 U850 ( .A(KEYINPUT1), .B(n1056), .ZN(n1187) );
INV_X1 U851 ( .A(n1189), .ZN(n1056) );
INV_X1 U852 ( .A(n1064), .ZN(n1070) );
NAND2_X1 U853 ( .A1(n1138), .A2(n1190), .ZN(n1185) );
NAND2_X1 U854 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NAND4_X1 U855 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1025), .ZN(n1115) );
NAND2_X1 U856 ( .A1(n1071), .A2(n1196), .ZN(n1025) );
INV_X1 U857 ( .A(n1192), .ZN(n1196) );
NAND2_X1 U858 ( .A1(n1141), .A2(n1036), .ZN(n1192) );
XOR2_X1 U859 ( .A(n1116), .B(KEYINPUT9), .Z(n1173) );
NAND2_X1 U860 ( .A1(n1197), .A2(n1198), .ZN(n1170) );
NAND2_X1 U861 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U862 ( .A(n1201), .B(KEYINPUT11), .Z(n1197) );
OR2_X1 U863 ( .A1(n1200), .A2(n1199), .ZN(n1201) );
NAND3_X1 U864 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1200) );
OR2_X1 U865 ( .A1(n1205), .A2(KEYINPUT31), .ZN(n1203) );
NAND2_X1 U866 ( .A1(KEYINPUT31), .A2(n1206), .ZN(n1202) );
NOR2_X1 U867 ( .A1(n1039), .A2(G952), .ZN(n1118) );
XNOR2_X1 U868 ( .A(G146), .B(n1182), .ZN(G48) );
NAND4_X1 U869 ( .A1(n1207), .A2(n1138), .A3(n1054), .A4(n1075), .ZN(n1182) );
XNOR2_X1 U870 ( .A(G143), .B(n1181), .ZN(G45) );
NAND4_X1 U871 ( .A1(n1208), .A2(n1184), .A3(n1209), .A4(n1189), .ZN(n1181) );
XNOR2_X1 U872 ( .A(G140), .B(n1180), .ZN(G42) );
NAND4_X1 U873 ( .A1(n1210), .A2(n1138), .A3(n1069), .A4(n1211), .ZN(n1180) );
XNOR2_X1 U874 ( .A(G137), .B(n1179), .ZN(G39) );
NAND3_X1 U875 ( .A1(n1068), .A2(n1075), .A3(n1210), .ZN(n1179) );
AND3_X1 U876 ( .A1(n1054), .A2(n1212), .A3(n1037), .ZN(n1210) );
XNOR2_X1 U877 ( .A(G134), .B(n1213), .ZN(G36) );
NAND2_X1 U878 ( .A1(KEYINPUT20), .A2(n1214), .ZN(n1213) );
INV_X1 U879 ( .A(n1178), .ZN(n1214) );
NAND3_X1 U880 ( .A1(n1037), .A2(n1071), .A3(n1184), .ZN(n1178) );
NAND2_X1 U881 ( .A1(n1215), .A2(n1216), .ZN(G33) );
NAND2_X1 U882 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
INV_X1 U883 ( .A(G131), .ZN(n1218) );
XOR2_X1 U884 ( .A(n1219), .B(KEYINPUT30), .Z(n1217) );
NAND2_X1 U885 ( .A1(G131), .A2(n1220), .ZN(n1215) );
XOR2_X1 U886 ( .A(n1219), .B(KEYINPUT56), .Z(n1220) );
NAND3_X1 U887 ( .A1(n1138), .A2(n1221), .A3(n1184), .ZN(n1219) );
AND3_X1 U888 ( .A1(n1054), .A2(n1212), .A3(n1222), .ZN(n1184) );
XOR2_X1 U889 ( .A(n1145), .B(KEYINPUT45), .Z(n1054) );
XOR2_X1 U890 ( .A(KEYINPUT60), .B(n1037), .Z(n1221) );
NOR2_X1 U891 ( .A1(n1223), .A2(n1058), .ZN(n1037) );
NAND2_X1 U892 ( .A1(n1224), .A2(n1225), .ZN(G30) );
NAND2_X1 U893 ( .A1(G128), .A2(n1177), .ZN(n1225) );
XOR2_X1 U894 ( .A(KEYINPUT22), .B(n1226), .Z(n1224) );
NOR2_X1 U895 ( .A1(G128), .A2(n1177), .ZN(n1226) );
NAND4_X1 U896 ( .A1(n1207), .A2(n1071), .A3(n1145), .A4(n1075), .ZN(n1177) );
XOR2_X1 U897 ( .A(G101), .B(n1227), .Z(G3) );
NOR2_X1 U898 ( .A1(n1228), .A2(n1064), .ZN(n1227) );
NAND2_X1 U899 ( .A1(n1046), .A2(n1222), .ZN(n1064) );
XOR2_X1 U900 ( .A(G125), .B(n1229), .Z(G27) );
NOR2_X1 U901 ( .A1(KEYINPUT46), .A2(n1176), .ZN(n1229) );
NAND4_X1 U902 ( .A1(n1207), .A2(n1138), .A3(n1069), .A4(n1035), .ZN(n1176) );
INV_X1 U903 ( .A(n1033), .ZN(n1138) );
AND3_X1 U904 ( .A1(n1189), .A2(n1212), .A3(n1211), .ZN(n1207) );
NAND2_X1 U905 ( .A1(n1034), .A2(n1230), .ZN(n1212) );
NAND3_X1 U906 ( .A1(G902), .A2(n1231), .A3(n1092), .ZN(n1230) );
NOR2_X1 U907 ( .A1(n1039), .A2(G900), .ZN(n1092) );
XNOR2_X1 U908 ( .A(G122), .B(n1194), .ZN(G24) );
NAND4_X1 U909 ( .A1(n1208), .A2(n1232), .A3(n1209), .A4(n1036), .ZN(n1194) );
NOR2_X1 U910 ( .A1(n1075), .A2(n1211), .ZN(n1036) );
XOR2_X1 U911 ( .A(G119), .B(n1116), .Z(G21) );
AND3_X1 U912 ( .A1(n1232), .A2(n1075), .A3(n1068), .ZN(n1116) );
XNOR2_X1 U913 ( .A(G116), .B(n1195), .ZN(G18) );
NAND2_X1 U914 ( .A1(n1233), .A2(n1071), .ZN(n1195) );
NOR2_X1 U915 ( .A1(n1234), .A2(n1235), .ZN(n1071) );
INV_X1 U916 ( .A(n1191), .ZN(n1233) );
NAND2_X1 U917 ( .A1(n1222), .A2(n1232), .ZN(n1191) );
INV_X1 U918 ( .A(n1236), .ZN(n1232) );
XNOR2_X1 U919 ( .A(n1237), .B(n1238), .ZN(G15) );
NOR3_X1 U920 ( .A1(n1239), .A2(n1236), .A3(n1033), .ZN(n1238) );
NAND2_X1 U921 ( .A1(n1208), .A2(n1234), .ZN(n1033) );
XOR2_X1 U922 ( .A(n1235), .B(KEYINPUT5), .Z(n1208) );
NAND2_X1 U923 ( .A1(n1035), .A2(n1143), .ZN(n1236) );
INV_X1 U924 ( .A(n1063), .ZN(n1035) );
NAND2_X1 U925 ( .A1(n1053), .A2(n1240), .ZN(n1063) );
XOR2_X1 U926 ( .A(KEYINPUT29), .B(n1222), .Z(n1239) );
NOR2_X1 U927 ( .A1(n1211), .A2(n1069), .ZN(n1222) );
XNOR2_X1 U928 ( .A(G110), .B(n1241), .ZN(G12) );
NAND2_X1 U929 ( .A1(KEYINPUT39), .A2(n1242), .ZN(n1241) );
INV_X1 U930 ( .A(n1193), .ZN(n1242) );
NAND3_X1 U931 ( .A1(n1069), .A2(n1141), .A3(n1068), .ZN(n1193) );
AND2_X1 U932 ( .A1(n1046), .A2(n1211), .ZN(n1068) );
XOR2_X1 U933 ( .A(n1078), .B(KEYINPUT3), .Z(n1211) );
XNOR2_X1 U934 ( .A(n1243), .B(n1122), .ZN(n1078) );
NAND2_X1 U935 ( .A1(G217), .A2(n1244), .ZN(n1122) );
NAND2_X1 U936 ( .A1(n1120), .A2(n1245), .ZN(n1243) );
XNOR2_X1 U937 ( .A(n1246), .B(n1247), .ZN(n1120) );
XOR2_X1 U938 ( .A(G137), .B(n1248), .Z(n1247) );
NOR2_X1 U939 ( .A1(KEYINPUT41), .A2(n1249), .ZN(n1248) );
XOR2_X1 U940 ( .A(n1250), .B(n1251), .Z(n1249) );
XOR2_X1 U941 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U942 ( .A(n1254), .B(n1255), .Z(n1250) );
XNOR2_X1 U943 ( .A(G146), .B(KEYINPUT13), .ZN(n1255) );
NAND2_X1 U944 ( .A1(n1256), .A2(n1257), .ZN(n1254) );
NAND2_X1 U945 ( .A1(G119), .A2(n1258), .ZN(n1257) );
XOR2_X1 U946 ( .A(KEYINPUT63), .B(n1259), .Z(n1256) );
NOR2_X1 U947 ( .A1(G119), .A2(n1258), .ZN(n1259) );
NAND4_X1 U948 ( .A1(KEYINPUT49), .A2(G221), .A3(G234), .A4(n1039), .ZN(n1246) );
NOR2_X1 U949 ( .A1(n1209), .A2(n1235), .ZN(n1046) );
XNOR2_X1 U950 ( .A(n1081), .B(n1082), .ZN(n1235) );
XOR2_X1 U951 ( .A(G475), .B(KEYINPUT25), .Z(n1082) );
NOR2_X1 U952 ( .A1(n1134), .A2(G902), .ZN(n1081) );
XNOR2_X1 U953 ( .A(n1260), .B(n1261), .ZN(n1134) );
XNOR2_X1 U954 ( .A(KEYINPUT38), .B(n1262), .ZN(n1261) );
XNOR2_X1 U955 ( .A(n1263), .B(n1264), .ZN(n1260) );
NOR2_X1 U956 ( .A1(KEYINPUT47), .A2(n1265), .ZN(n1264) );
XOR2_X1 U957 ( .A(n1266), .B(n1267), .Z(n1265) );
XNOR2_X1 U958 ( .A(n1268), .B(n1269), .ZN(n1267) );
NOR2_X1 U959 ( .A1(KEYINPUT33), .A2(n1270), .ZN(n1269) );
XOR2_X1 U960 ( .A(n1096), .B(G146), .Z(n1270) );
XNOR2_X1 U961 ( .A(G140), .B(n1252), .ZN(n1096) );
XNOR2_X1 U962 ( .A(n1271), .B(n1097), .ZN(n1266) );
INV_X1 U963 ( .A(n1272), .ZN(n1097) );
NAND2_X1 U964 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
XNOR2_X1 U965 ( .A(G214), .B(KEYINPUT35), .ZN(n1273) );
INV_X1 U966 ( .A(n1234), .ZN(n1209) );
XOR2_X1 U967 ( .A(n1077), .B(KEYINPUT36), .Z(n1234) );
XNOR2_X1 U968 ( .A(n1275), .B(G478), .ZN(n1077) );
NAND2_X1 U969 ( .A1(n1128), .A2(n1245), .ZN(n1275) );
XOR2_X1 U970 ( .A(n1276), .B(n1277), .Z(n1128) );
XOR2_X1 U971 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U972 ( .A(n1280), .B(n1281), .Z(n1279) );
AND3_X1 U973 ( .A1(n1282), .A2(G217), .A3(G234), .ZN(n1281) );
XNOR2_X1 U974 ( .A(KEYINPUT58), .B(G953), .ZN(n1282) );
NOR2_X1 U975 ( .A1(KEYINPUT53), .A2(n1283), .ZN(n1280) );
XNOR2_X1 U976 ( .A(G143), .B(G128), .ZN(n1283) );
NOR2_X1 U977 ( .A1(G107), .A2(KEYINPUT42), .ZN(n1278) );
XNOR2_X1 U978 ( .A(G116), .B(n1284), .ZN(n1276) );
XNOR2_X1 U979 ( .A(n1285), .B(G122), .ZN(n1284) );
INV_X1 U980 ( .A(n1228), .ZN(n1141) );
NAND2_X1 U981 ( .A1(n1145), .A2(n1143), .ZN(n1228) );
AND2_X1 U982 ( .A1(n1189), .A2(n1188), .ZN(n1143) );
NAND2_X1 U983 ( .A1(n1034), .A2(n1286), .ZN(n1188) );
NAND4_X1 U984 ( .A1(G902), .A2(G953), .A3(n1231), .A4(n1110), .ZN(n1286) );
INV_X1 U985 ( .A(G898), .ZN(n1110) );
NAND3_X1 U986 ( .A1(n1231), .A2(n1039), .A3(G952), .ZN(n1034) );
NAND2_X1 U987 ( .A1(G237), .A2(G234), .ZN(n1231) );
NOR2_X1 U988 ( .A1(n1059), .A2(n1058), .ZN(n1189) );
AND2_X1 U989 ( .A1(G214), .A2(n1287), .ZN(n1058) );
XOR2_X1 U990 ( .A(KEYINPUT37), .B(n1288), .Z(n1287) );
NOR2_X1 U991 ( .A1(G237), .A2(G902), .ZN(n1288) );
INV_X1 U992 ( .A(n1223), .ZN(n1059) );
NAND3_X1 U993 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1223) );
OR2_X1 U994 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND3_X1 U995 ( .A1(n1293), .A2(n1292), .A3(n1245), .ZN(n1290) );
NAND2_X1 U996 ( .A1(G237), .A2(G210), .ZN(n1292) );
XNOR2_X1 U997 ( .A(n1294), .B(n1199), .ZN(n1293) );
XNOR2_X1 U998 ( .A(n1112), .B(n1113), .ZN(n1199) );
XNOR2_X1 U999 ( .A(n1295), .B(G110), .ZN(n1113) );
NAND2_X1 U1000 ( .A1(KEYINPUT14), .A2(n1262), .ZN(n1295) );
INV_X1 U1001 ( .A(G122), .ZN(n1262) );
XOR2_X1 U1002 ( .A(n1296), .B(n1297), .Z(n1112) );
XOR2_X1 U1003 ( .A(G101), .B(n1298), .Z(n1297) );
XNOR2_X1 U1004 ( .A(KEYINPUT12), .B(n1299), .ZN(n1298) );
XOR2_X1 U1005 ( .A(n1300), .B(n1263), .Z(n1296) );
XNOR2_X1 U1006 ( .A(G104), .B(n1237), .ZN(n1263) );
NAND2_X1 U1007 ( .A1(n1204), .A2(n1205), .ZN(n1294) );
NAND3_X1 U1008 ( .A1(n1301), .A2(n1039), .A3(G224), .ZN(n1205) );
NAND2_X1 U1009 ( .A1(n1206), .A2(n1302), .ZN(n1204) );
NAND2_X1 U1010 ( .A1(G224), .A2(n1039), .ZN(n1302) );
INV_X1 U1011 ( .A(n1301), .ZN(n1206) );
XNOR2_X1 U1012 ( .A(n1252), .B(n1303), .ZN(n1301) );
XOR2_X1 U1013 ( .A(G125), .B(KEYINPUT61), .Z(n1252) );
NAND2_X1 U1014 ( .A1(G902), .A2(G210), .ZN(n1289) );
NOR2_X1 U1015 ( .A1(n1053), .A2(n1052), .ZN(n1145) );
INV_X1 U1016 ( .A(n1240), .ZN(n1052) );
NAND2_X1 U1017 ( .A1(n1304), .A2(n1244), .ZN(n1240) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1245), .ZN(n1244) );
XOR2_X1 U1019 ( .A(KEYINPUT28), .B(G221), .Z(n1304) );
XNOR2_X1 U1020 ( .A(n1305), .B(n1162), .ZN(n1053) );
INV_X1 U1021 ( .A(G469), .ZN(n1162) );
NAND4_X1 U1022 ( .A1(n1306), .A2(n1245), .A3(n1307), .A4(n1308), .ZN(n1305) );
NAND3_X1 U1023 ( .A1(n1168), .A2(n1309), .A3(n1158), .ZN(n1308) );
NAND2_X1 U1024 ( .A1(n1164), .A2(n1310), .ZN(n1307) );
INV_X1 U1025 ( .A(n1158), .ZN(n1310) );
NOR2_X1 U1026 ( .A1(n1309), .A2(n1311), .ZN(n1164) );
INV_X1 U1027 ( .A(n1166), .ZN(n1309) );
NAND2_X1 U1028 ( .A1(n1311), .A2(n1312), .ZN(n1306) );
XNOR2_X1 U1029 ( .A(n1166), .B(n1158), .ZN(n1312) );
XNOR2_X1 U1030 ( .A(n1313), .B(n1253), .ZN(n1158) );
XOR2_X1 U1031 ( .A(G110), .B(G140), .Z(n1253) );
NAND2_X1 U1032 ( .A1(G227), .A2(n1039), .ZN(n1313) );
INV_X1 U1033 ( .A(G953), .ZN(n1039) );
XOR2_X1 U1034 ( .A(G101), .B(n1314), .Z(n1166) );
NOR2_X1 U1035 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
AND3_X1 U1036 ( .A1(KEYINPUT7), .A2(n1299), .A3(G104), .ZN(n1316) );
NOR2_X1 U1037 ( .A1(KEYINPUT7), .A2(n1317), .ZN(n1315) );
XNOR2_X1 U1038 ( .A(n1299), .B(G104), .ZN(n1317) );
INV_X1 U1039 ( .A(G107), .ZN(n1299) );
INV_X1 U1040 ( .A(n1168), .ZN(n1311) );
XOR2_X1 U1041 ( .A(n1095), .B(n1318), .Z(n1168) );
INV_X1 U1042 ( .A(n1319), .ZN(n1318) );
XOR2_X1 U1043 ( .A(n1320), .B(KEYINPUT6), .Z(n1095) );
NAND3_X1 U1044 ( .A1(n1321), .A2(n1322), .A3(n1323), .ZN(n1320) );
NAND2_X1 U1045 ( .A1(G128), .A2(n1324), .ZN(n1323) );
NAND2_X1 U1046 ( .A1(n1325), .A2(n1326), .ZN(n1322) );
INV_X1 U1047 ( .A(KEYINPUT59), .ZN(n1326) );
NAND2_X1 U1048 ( .A1(n1327), .A2(n1258), .ZN(n1325) );
XNOR2_X1 U1049 ( .A(KEYINPUT26), .B(n1324), .ZN(n1327) );
NAND2_X1 U1050 ( .A1(KEYINPUT59), .A2(n1328), .ZN(n1321) );
NAND2_X1 U1051 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
OR3_X1 U1052 ( .A1(n1324), .A2(G128), .A3(KEYINPUT26), .ZN(n1330) );
NAND2_X1 U1053 ( .A1(KEYINPUT26), .A2(n1324), .ZN(n1329) );
INV_X1 U1054 ( .A(n1075), .ZN(n1069) );
XOR2_X1 U1055 ( .A(n1331), .B(n1151), .Z(n1075) );
INV_X1 U1056 ( .A(G472), .ZN(n1151) );
NAND2_X1 U1057 ( .A1(n1332), .A2(n1245), .ZN(n1331) );
INV_X1 U1058 ( .A(G902), .ZN(n1245) );
XOR2_X1 U1059 ( .A(n1333), .B(n1334), .Z(n1332) );
XOR2_X1 U1060 ( .A(n1149), .B(n1154), .Z(n1334) );
XOR2_X1 U1061 ( .A(n1335), .B(G101), .Z(n1154) );
NAND2_X1 U1062 ( .A1(G210), .A2(n1274), .ZN(n1335) );
NOR2_X1 U1063 ( .A1(G953), .A2(G237), .ZN(n1274) );
XNOR2_X1 U1064 ( .A(n1319), .B(n1303), .ZN(n1149) );
XNOR2_X1 U1065 ( .A(n1258), .B(n1336), .ZN(n1303) );
NOR2_X1 U1066 ( .A1(KEYINPUT23), .A2(n1324), .ZN(n1336) );
XNOR2_X1 U1067 ( .A(n1268), .B(G146), .ZN(n1324) );
INV_X1 U1068 ( .A(G143), .ZN(n1268) );
INV_X1 U1069 ( .A(G128), .ZN(n1258) );
XOR2_X1 U1070 ( .A(n1272), .B(n1337), .Z(n1319) );
XOR2_X1 U1071 ( .A(G137), .B(n1338), .Z(n1337) );
NOR2_X1 U1072 ( .A1(KEYINPUT34), .A2(n1285), .ZN(n1338) );
INV_X1 U1073 ( .A(G134), .ZN(n1285) );
XOR2_X1 U1074 ( .A(G131), .B(KEYINPUT48), .Z(n1272) );
XNOR2_X1 U1075 ( .A(n1339), .B(KEYINPUT55), .ZN(n1333) );
NAND2_X1 U1076 ( .A1(KEYINPUT15), .A2(n1152), .ZN(n1339) );
AND2_X1 U1077 ( .A1(n1340), .A2(n1341), .ZN(n1152) );
NAND2_X1 U1078 ( .A1(n1300), .A2(n1237), .ZN(n1341) );
XOR2_X1 U1079 ( .A(KEYINPUT17), .B(n1342), .Z(n1340) );
NOR2_X1 U1080 ( .A1(n1300), .A2(n1237), .ZN(n1342) );
INV_X1 U1081 ( .A(G113), .ZN(n1237) );
XNOR2_X1 U1082 ( .A(G116), .B(n1343), .ZN(n1300) );
XOR2_X1 U1083 ( .A(KEYINPUT44), .B(G119), .Z(n1343) );
endmodule


