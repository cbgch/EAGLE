//Key = 0100110101100101111111110110010101000011011010001111100110100101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325;

XNOR2_X1 U725 ( .A(G107), .B(n996), .ZN(G9) );
NOR2_X1 U726 ( .A1(n997), .A2(KEYINPUT36), .ZN(n996) );
INV_X1 U727 ( .A(n998), .ZN(n997) );
NOR2_X1 U728 ( .A1(n999), .A2(n1000), .ZN(G75) );
NOR3_X1 U729 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n1000) );
NOR2_X1 U730 ( .A1(n1004), .A2(n1005), .ZN(n1002) );
INV_X1 U731 ( .A(n1006), .ZN(n1005) );
NOR2_X1 U732 ( .A1(n1007), .A2(n1008), .ZN(n1004) );
XOR2_X1 U733 ( .A(n1009), .B(KEYINPUT16), .Z(n1008) );
NAND4_X1 U734 ( .A1(n1010), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1009) );
NOR3_X1 U735 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1007) );
NOR4_X1 U736 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
NOR4_X1 U737 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1020) );
INV_X1 U738 ( .A(KEYINPUT41), .ZN(n1023) );
NOR2_X1 U739 ( .A1(n1025), .A2(n1026), .ZN(n1018) );
INV_X1 U740 ( .A(n1011), .ZN(n1026) );
NOR2_X1 U741 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR2_X1 U742 ( .A1(n1029), .A2(n1030), .ZN(n1015) );
NOR4_X1 U743 ( .A1(KEYINPUT41), .A2(n1021), .A3(n1022), .A4(n1024), .ZN(n1030) );
NAND3_X1 U744 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1001) );
NAND4_X1 U745 ( .A1(n1010), .A2(n1011), .A3(n1013), .A4(n1034), .ZN(n1033) );
NAND2_X1 U746 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U747 ( .A1(n1029), .A2(n1037), .ZN(n1036) );
NAND2_X1 U748 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U749 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
XOR2_X1 U750 ( .A(KEYINPUT55), .B(n1042), .Z(n1041) );
NAND2_X1 U751 ( .A1(n1006), .A2(n1043), .ZN(n1035) );
INV_X1 U752 ( .A(n1014), .ZN(n1010) );
NOR3_X1 U753 ( .A1(n1044), .A2(G953), .A3(G952), .ZN(n999) );
INV_X1 U754 ( .A(n1031), .ZN(n1044) );
NAND4_X1 U755 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1031) );
NOR4_X1 U756 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
XOR2_X1 U757 ( .A(n1053), .B(n1054), .Z(n1052) );
XOR2_X1 U758 ( .A(n1055), .B(n1056), .Z(n1050) );
XOR2_X1 U759 ( .A(KEYINPUT61), .B(G475), .Z(n1056) );
XOR2_X1 U760 ( .A(n1057), .B(KEYINPUT44), .Z(n1049) );
NAND2_X1 U761 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR3_X1 U762 ( .A1(n1060), .A2(n1061), .A3(n1040), .ZN(n1047) );
NOR2_X1 U763 ( .A1(n1058), .A2(n1059), .ZN(n1060) );
XOR2_X1 U764 ( .A(G469), .B(KEYINPUT48), .Z(n1059) );
INV_X1 U765 ( .A(n1062), .ZN(n1058) );
XNOR2_X1 U766 ( .A(n1063), .B(n1064), .ZN(n1046) );
NOR2_X1 U767 ( .A1(n1065), .A2(KEYINPUT59), .ZN(n1064) );
XOR2_X1 U768 ( .A(n1066), .B(n1067), .Z(n1045) );
XNOR2_X1 U769 ( .A(n1068), .B(KEYINPUT22), .ZN(n1067) );
NAND3_X1 U770 ( .A1(n1069), .A2(n1070), .A3(KEYINPUT19), .ZN(n1068) );
XOR2_X1 U771 ( .A(n1071), .B(n1072), .Z(G72) );
NOR2_X1 U772 ( .A1(n1073), .A2(n1032), .ZN(n1072) );
AND2_X1 U773 ( .A1(G227), .A2(G900), .ZN(n1073) );
NAND2_X1 U774 ( .A1(n1074), .A2(n1075), .ZN(n1071) );
NAND2_X1 U775 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U776 ( .A(n1078), .B(KEYINPUT8), .Z(n1074) );
OR2_X1 U777 ( .A1(n1077), .A2(n1076), .ZN(n1078) );
AND2_X1 U778 ( .A1(n1079), .A2(n1080), .ZN(n1076) );
NAND2_X1 U779 ( .A1(G953), .A2(n1081), .ZN(n1080) );
XOR2_X1 U780 ( .A(n1082), .B(n1083), .Z(n1079) );
XOR2_X1 U781 ( .A(n1084), .B(n1085), .Z(n1083) );
NAND2_X1 U782 ( .A1(KEYINPUT10), .A2(n1086), .ZN(n1085) );
XOR2_X1 U783 ( .A(n1087), .B(n1088), .Z(n1082) );
NAND2_X1 U784 ( .A1(n1032), .A2(n1089), .ZN(n1077) );
NAND3_X1 U785 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
XOR2_X1 U786 ( .A(n1093), .B(KEYINPUT14), .Z(n1092) );
NAND2_X1 U787 ( .A1(n1094), .A2(n1095), .ZN(G69) );
NAND2_X1 U788 ( .A1(n1096), .A2(n1032), .ZN(n1095) );
XOR2_X1 U789 ( .A(n1097), .B(n1098), .Z(n1096) );
NAND2_X1 U790 ( .A1(n1099), .A2(G953), .ZN(n1094) );
XOR2_X1 U791 ( .A(n1097), .B(n1100), .Z(n1099) );
NOR2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U793 ( .A1(KEYINPUT35), .A2(n1103), .ZN(n1097) );
NOR2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XOR2_X1 U795 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U796 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U797 ( .A1(n1110), .A2(KEYINPUT5), .ZN(n1108) );
XNOR2_X1 U798 ( .A(n1111), .B(n1112), .ZN(n1110) );
XOR2_X1 U799 ( .A(G122), .B(G110), .Z(n1106) );
NOR2_X1 U800 ( .A1(G898), .A2(n1032), .ZN(n1104) );
NOR2_X1 U801 ( .A1(n1113), .A2(n1114), .ZN(G66) );
XOR2_X1 U802 ( .A(n1069), .B(n1115), .Z(n1114) );
XNOR2_X1 U803 ( .A(n1116), .B(KEYINPUT40), .ZN(n1115) );
NAND2_X1 U804 ( .A1(KEYINPUT20), .A2(n1117), .ZN(n1116) );
NAND2_X1 U805 ( .A1(n1118), .A2(n1066), .ZN(n1117) );
NOR2_X1 U806 ( .A1(n1113), .A2(n1119), .ZN(G63) );
XNOR2_X1 U807 ( .A(n1120), .B(n1121), .ZN(n1119) );
AND2_X1 U808 ( .A1(G478), .A2(n1118), .ZN(n1121) );
INV_X1 U809 ( .A(n1122), .ZN(n1118) );
NOR2_X1 U810 ( .A1(n1113), .A2(n1123), .ZN(G60) );
XNOR2_X1 U811 ( .A(n1124), .B(n1125), .ZN(n1123) );
NOR2_X1 U812 ( .A1(n1126), .A2(n1122), .ZN(n1125) );
XOR2_X1 U813 ( .A(G104), .B(n1127), .Z(G6) );
NOR2_X1 U814 ( .A1(n1128), .A2(n1038), .ZN(n1127) );
XOR2_X1 U815 ( .A(n1129), .B(KEYINPUT57), .Z(n1128) );
NOR2_X1 U816 ( .A1(n1113), .A2(n1130), .ZN(G57) );
XOR2_X1 U817 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U818 ( .A(n1133), .B(KEYINPUT53), .ZN(n1132) );
NAND2_X1 U819 ( .A1(KEYINPUT63), .A2(n1134), .ZN(n1133) );
XOR2_X1 U820 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U821 ( .A1(n1053), .A2(n1122), .ZN(n1136) );
INV_X1 U822 ( .A(G472), .ZN(n1053) );
NOR2_X1 U823 ( .A1(KEYINPUT6), .A2(n1137), .ZN(n1135) );
XOR2_X1 U824 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U825 ( .A(n1140), .B(n1141), .Z(n1138) );
NAND2_X1 U826 ( .A1(KEYINPUT49), .A2(n1142), .ZN(n1140) );
NOR2_X1 U827 ( .A1(n1113), .A2(n1143), .ZN(G54) );
XOR2_X1 U828 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U829 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U830 ( .A1(n1148), .A2(n1122), .ZN(n1147) );
NOR2_X1 U831 ( .A1(n1149), .A2(n1150), .ZN(n1146) );
XOR2_X1 U832 ( .A(n1151), .B(KEYINPUT52), .Z(n1150) );
NAND2_X1 U833 ( .A1(n1152), .A2(n1087), .ZN(n1151) );
NOR2_X1 U834 ( .A1(n1087), .A2(n1152), .ZN(n1149) );
XOR2_X1 U835 ( .A(n1153), .B(KEYINPUT12), .Z(n1152) );
XOR2_X1 U836 ( .A(n1154), .B(n1155), .Z(n1144) );
XOR2_X1 U837 ( .A(G140), .B(G110), .Z(n1155) );
NOR2_X1 U838 ( .A1(n1113), .A2(n1156), .ZN(G51) );
XOR2_X1 U839 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U840 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND2_X1 U841 ( .A1(n1161), .A2(KEYINPUT39), .ZN(n1160) );
XNOR2_X1 U842 ( .A(n1162), .B(n1163), .ZN(n1161) );
NAND2_X1 U843 ( .A1(n1164), .A2(n1165), .ZN(n1159) );
NAND2_X1 U844 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U845 ( .A(KEYINPUT13), .B(n1168), .Z(n1164) );
NOR2_X1 U846 ( .A1(n1167), .A2(n1166), .ZN(n1168) );
XOR2_X1 U847 ( .A(n1086), .B(n1141), .Z(n1166) );
NOR2_X1 U848 ( .A1(n1169), .A2(n1122), .ZN(n1157) );
NAND2_X1 U849 ( .A1(G902), .A2(n1003), .ZN(n1122) );
NAND4_X1 U850 ( .A1(n1098), .A2(n1090), .A3(n1170), .A4(n1093), .ZN(n1003) );
XNOR2_X1 U851 ( .A(KEYINPUT50), .B(n1091), .ZN(n1170) );
AND4_X1 U852 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1090) );
AND3_X1 U853 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1174) );
AND4_X1 U854 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1098) );
AND4_X1 U855 ( .A1(n998), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1181) );
NAND4_X1 U856 ( .A1(n1185), .A2(n1027), .A3(n1029), .A4(n1186), .ZN(n998) );
NAND2_X1 U857 ( .A1(n1187), .A2(n1019), .ZN(n1180) );
NAND2_X1 U858 ( .A1(n1188), .A2(n1189), .ZN(n1178) );
NAND2_X1 U859 ( .A1(n1190), .A2(n1129), .ZN(n1189) );
NAND4_X1 U860 ( .A1(n1185), .A2(n1029), .A3(n1028), .A4(n1191), .ZN(n1129) );
NOR2_X1 U861 ( .A1(n1032), .A2(G952), .ZN(n1113) );
XOR2_X1 U862 ( .A(n1192), .B(n1093), .Z(G48) );
NAND3_X1 U863 ( .A1(n1188), .A2(n1028), .A3(n1193), .ZN(n1093) );
XOR2_X1 U864 ( .A(G143), .B(n1194), .Z(G45) );
NOR2_X1 U865 ( .A1(KEYINPUT2), .A2(n1173), .ZN(n1194) );
NAND4_X1 U866 ( .A1(n1195), .A2(n1196), .A3(n1188), .A4(n1051), .ZN(n1173) );
XOR2_X1 U867 ( .A(n1084), .B(n1091), .Z(G42) );
NAND4_X1 U868 ( .A1(n1006), .A2(n1012), .A3(n1197), .A4(n1185), .ZN(n1091) );
NOR2_X1 U869 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U870 ( .A(n1200), .B(n1171), .Z(G39) );
NAND3_X1 U871 ( .A1(n1193), .A2(n1013), .A3(n1006), .ZN(n1171) );
XNOR2_X1 U872 ( .A(G134), .B(n1172), .ZN(G36) );
NAND3_X1 U873 ( .A1(n1006), .A2(n1027), .A3(n1196), .ZN(n1172) );
XNOR2_X1 U874 ( .A(G131), .B(n1175), .ZN(G33) );
NAND3_X1 U875 ( .A1(n1006), .A2(n1028), .A3(n1196), .ZN(n1175) );
AND3_X1 U876 ( .A1(n1185), .A2(n1201), .A3(n1043), .ZN(n1196) );
INV_X1 U877 ( .A(n1202), .ZN(n1185) );
NOR2_X1 U878 ( .A1(n1042), .A2(n1040), .ZN(n1006) );
INV_X1 U879 ( .A(n1203), .ZN(n1040) );
XOR2_X1 U880 ( .A(n1177), .B(n1204), .Z(G30) );
NAND2_X1 U881 ( .A1(KEYINPUT9), .A2(G128), .ZN(n1204) );
NAND3_X1 U882 ( .A1(n1027), .A2(n1188), .A3(n1193), .ZN(n1177) );
NOR4_X1 U883 ( .A1(n1202), .A2(n1205), .A3(n1206), .A4(n1198), .ZN(n1193) );
INV_X1 U884 ( .A(n1038), .ZN(n1188) );
XOR2_X1 U885 ( .A(G101), .B(n1207), .Z(G3) );
AND2_X1 U886 ( .A1(n1019), .A2(n1187), .ZN(n1207) );
XOR2_X1 U887 ( .A(n1176), .B(n1208), .Z(G27) );
NAND2_X1 U888 ( .A1(KEYINPUT38), .A2(G125), .ZN(n1208) );
NAND3_X1 U889 ( .A1(n1011), .A2(n1012), .A3(n1209), .ZN(n1176) );
NOR3_X1 U890 ( .A1(n1038), .A2(n1198), .A3(n1199), .ZN(n1209) );
INV_X1 U891 ( .A(n1028), .ZN(n1199) );
INV_X1 U892 ( .A(n1201), .ZN(n1198) );
NAND2_X1 U893 ( .A1(n1014), .A2(n1210), .ZN(n1201) );
NAND4_X1 U894 ( .A1(G953), .A2(G902), .A3(n1211), .A4(n1081), .ZN(n1210) );
INV_X1 U895 ( .A(G900), .ZN(n1081) );
XNOR2_X1 U896 ( .A(G122), .B(n1179), .ZN(G24) );
NAND3_X1 U897 ( .A1(n1195), .A2(n1011), .A3(n1212), .ZN(n1179) );
AND3_X1 U898 ( .A1(n1029), .A2(n1051), .A3(n1186), .ZN(n1212) );
INV_X1 U899 ( .A(n1017), .ZN(n1029) );
NAND2_X1 U900 ( .A1(n1213), .A2(n1206), .ZN(n1017) );
XOR2_X1 U901 ( .A(G119), .B(n1214), .Z(G21) );
NOR2_X1 U902 ( .A1(n1215), .A2(n1038), .ZN(n1214) );
XOR2_X1 U903 ( .A(n1190), .B(KEYINPUT32), .Z(n1215) );
NAND3_X1 U904 ( .A1(n1011), .A2(n1013), .A3(n1216), .ZN(n1190) );
NOR3_X1 U905 ( .A1(n1205), .A2(n1217), .A3(n1206), .ZN(n1216) );
XNOR2_X1 U906 ( .A(G116), .B(n1184), .ZN(G18) );
NAND3_X1 U907 ( .A1(n1011), .A2(n1027), .A3(n1187), .ZN(n1184) );
NOR2_X1 U908 ( .A1(n1195), .A2(n1218), .ZN(n1027) );
XOR2_X1 U909 ( .A(n1219), .B(n1183), .Z(G15) );
NAND3_X1 U910 ( .A1(n1011), .A2(n1028), .A3(n1187), .ZN(n1183) );
AND2_X1 U911 ( .A1(n1043), .A2(n1186), .ZN(n1187) );
AND2_X1 U912 ( .A1(n1213), .A2(n1220), .ZN(n1043) );
NAND2_X1 U913 ( .A1(n1221), .A2(n1222), .ZN(n1028) );
OR3_X1 U914 ( .A1(n1223), .A2(n1051), .A3(KEYINPUT62), .ZN(n1222) );
INV_X1 U915 ( .A(n1218), .ZN(n1051) );
NAND2_X1 U916 ( .A1(KEYINPUT62), .A2(n1013), .ZN(n1221) );
INV_X1 U917 ( .A(n1022), .ZN(n1013) );
NOR2_X1 U918 ( .A1(n1224), .A2(n1024), .ZN(n1011) );
XOR2_X1 U919 ( .A(n1061), .B(KEYINPUT28), .Z(n1224) );
INV_X1 U920 ( .A(n1021), .ZN(n1061) );
XOR2_X1 U921 ( .A(n1182), .B(n1225), .Z(G12) );
XOR2_X1 U922 ( .A(KEYINPUT4), .B(G110), .Z(n1225) );
NAND3_X1 U923 ( .A1(n1012), .A2(n1186), .A3(n1019), .ZN(n1182) );
NOR2_X1 U924 ( .A1(n1022), .A2(n1202), .ZN(n1019) );
NAND2_X1 U925 ( .A1(n1226), .A2(n1024), .ZN(n1202) );
XNOR2_X1 U926 ( .A(n1148), .B(n1227), .ZN(n1024) );
NOR2_X1 U927 ( .A1(KEYINPUT27), .A2(n1062), .ZN(n1227) );
NAND2_X1 U928 ( .A1(n1070), .A2(n1228), .ZN(n1062) );
XOR2_X1 U929 ( .A(n1229), .B(n1230), .Z(n1228) );
XNOR2_X1 U930 ( .A(n1231), .B(n1154), .ZN(n1230) );
NAND2_X1 U931 ( .A1(G227), .A2(n1032), .ZN(n1154) );
NAND2_X1 U932 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NAND4_X1 U933 ( .A1(KEYINPUT31), .A2(KEYINPUT15), .A3(n1234), .A4(n1084), .ZN(n1233) );
NAND2_X1 U934 ( .A1(n1235), .A2(n1236), .ZN(n1232) );
NAND2_X1 U935 ( .A1(n1237), .A2(n1084), .ZN(n1236) );
OR2_X1 U936 ( .A1(n1234), .A2(KEYINPUT15), .ZN(n1237) );
NAND2_X1 U937 ( .A1(KEYINPUT31), .A2(n1234), .ZN(n1235) );
INV_X1 U938 ( .A(G110), .ZN(n1234) );
NAND3_X1 U939 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1229) );
NAND2_X1 U940 ( .A1(KEYINPUT37), .A2(n1241), .ZN(n1240) );
NAND3_X1 U941 ( .A1(n1153), .A2(n1242), .A3(n1087), .ZN(n1239) );
NAND2_X1 U942 ( .A1(n1139), .A2(n1243), .ZN(n1238) );
NAND2_X1 U943 ( .A1(n1244), .A2(n1242), .ZN(n1243) );
INV_X1 U944 ( .A(KEYINPUT37), .ZN(n1242) );
XOR2_X1 U945 ( .A(KEYINPUT58), .B(n1241), .Z(n1244) );
INV_X1 U946 ( .A(n1153), .ZN(n1241) );
XOR2_X1 U947 ( .A(n1245), .B(n1246), .Z(n1153) );
XOR2_X1 U948 ( .A(n1247), .B(n1088), .Z(n1246) );
XOR2_X1 U949 ( .A(n1141), .B(KEYINPUT18), .Z(n1088) );
INV_X1 U950 ( .A(n1248), .ZN(n1141) );
XOR2_X1 U951 ( .A(n1249), .B(KEYINPUT25), .Z(n1245) );
INV_X1 U952 ( .A(n1087), .ZN(n1139) );
INV_X1 U953 ( .A(G469), .ZN(n1148) );
XOR2_X1 U954 ( .A(n1021), .B(KEYINPUT28), .Z(n1226) );
NAND2_X1 U955 ( .A1(G221), .A2(n1250), .ZN(n1021) );
NAND2_X1 U956 ( .A1(n1218), .A2(n1223), .ZN(n1022) );
INV_X1 U957 ( .A(n1195), .ZN(n1223) );
XNOR2_X1 U958 ( .A(n1251), .B(n1055), .ZN(n1195) );
NAND2_X1 U959 ( .A1(n1124), .A2(n1070), .ZN(n1055) );
XNOR2_X1 U960 ( .A(n1252), .B(n1253), .ZN(n1124) );
XOR2_X1 U961 ( .A(n1254), .B(n1255), .Z(n1253) );
NAND2_X1 U962 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND2_X1 U963 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
INV_X1 U964 ( .A(n1260), .ZN(n1259) );
NAND2_X1 U965 ( .A1(n1261), .A2(n1262), .ZN(n1258) );
NAND2_X1 U966 ( .A1(n1263), .A2(n1084), .ZN(n1262) );
NAND2_X1 U967 ( .A1(n1264), .A2(G140), .ZN(n1261) );
NAND2_X1 U968 ( .A1(n1260), .A2(n1265), .ZN(n1256) );
NAND2_X1 U969 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NAND2_X1 U970 ( .A1(G140), .A2(n1263), .ZN(n1267) );
XOR2_X1 U971 ( .A(n1192), .B(KEYINPUT45), .Z(n1263) );
NAND2_X1 U972 ( .A1(n1264), .A2(n1084), .ZN(n1266) );
INV_X1 U973 ( .A(G140), .ZN(n1084) );
XOR2_X1 U974 ( .A(G146), .B(KEYINPUT0), .Z(n1264) );
NOR2_X1 U975 ( .A1(KEYINPUT11), .A2(n1086), .ZN(n1260) );
NAND2_X1 U976 ( .A1(G214), .A2(n1268), .ZN(n1254) );
XOR2_X1 U977 ( .A(n1269), .B(n1270), .Z(n1252) );
XOR2_X1 U978 ( .A(G143), .B(G131), .Z(n1270) );
NAND2_X1 U979 ( .A1(n1271), .A2(KEYINPUT51), .ZN(n1269) );
XOR2_X1 U980 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U981 ( .A(G104), .B(n1274), .Z(n1273) );
NOR2_X1 U982 ( .A1(G122), .A2(KEYINPUT24), .ZN(n1274) );
XOR2_X1 U983 ( .A(n1275), .B(G113), .Z(n1272) );
XNOR2_X1 U984 ( .A(KEYINPUT7), .B(KEYINPUT21), .ZN(n1275) );
NAND2_X1 U985 ( .A1(KEYINPUT1), .A2(n1126), .ZN(n1251) );
INV_X1 U986 ( .A(G475), .ZN(n1126) );
XOR2_X1 U987 ( .A(n1276), .B(G478), .Z(n1218) );
NAND2_X1 U988 ( .A1(n1070), .A2(n1120), .ZN(n1276) );
XNOR2_X1 U989 ( .A(n1277), .B(n1278), .ZN(n1120) );
XOR2_X1 U990 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U991 ( .A(n1281), .B(n1282), .Z(n1277) );
XOR2_X1 U992 ( .A(G134), .B(G107), .Z(n1282) );
NAND2_X1 U993 ( .A1(G217), .A2(n1283), .ZN(n1281) );
NOR2_X1 U994 ( .A1(n1038), .A2(n1217), .ZN(n1186) );
INV_X1 U995 ( .A(n1191), .ZN(n1217) );
NAND2_X1 U996 ( .A1(n1284), .A2(n1014), .ZN(n1191) );
NAND3_X1 U997 ( .A1(n1211), .A2(n1032), .A3(G952), .ZN(n1014) );
XOR2_X1 U998 ( .A(n1285), .B(KEYINPUT60), .Z(n1284) );
NAND4_X1 U999 ( .A1(G953), .A2(G902), .A3(n1211), .A4(n1102), .ZN(n1285) );
INV_X1 U1000 ( .A(G898), .ZN(n1102) );
NAND2_X1 U1001 ( .A1(G237), .A2(G234), .ZN(n1211) );
NAND2_X1 U1002 ( .A1(n1042), .A2(n1203), .ZN(n1038) );
NAND2_X1 U1003 ( .A1(G214), .A2(n1286), .ZN(n1203) );
XNOR2_X1 U1004 ( .A(n1063), .B(n1065), .ZN(n1042) );
INV_X1 U1005 ( .A(n1169), .ZN(n1065) );
NAND2_X1 U1006 ( .A1(G210), .A2(n1286), .ZN(n1169) );
NAND2_X1 U1007 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XOR2_X1 U1008 ( .A(KEYINPUT26), .B(G237), .Z(n1287) );
NAND2_X1 U1009 ( .A1(n1070), .A2(n1289), .ZN(n1063) );
XOR2_X1 U1010 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U1011 ( .A(n1292), .B(n1163), .Z(n1291) );
XNOR2_X1 U1012 ( .A(n1109), .B(n1293), .ZN(n1163) );
XOR2_X1 U1013 ( .A(n1112), .B(n1280), .Z(n1293) );
XOR2_X1 U1014 ( .A(G116), .B(G122), .Z(n1280) );
XOR2_X1 U1015 ( .A(G113), .B(KEYINPUT30), .Z(n1112) );
XOR2_X1 U1016 ( .A(n1294), .B(KEYINPUT33), .Z(n1109) );
NAND3_X1 U1017 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1294) );
NAND2_X1 U1018 ( .A1(n1298), .A2(n1249), .ZN(n1297) );
NAND2_X1 U1019 ( .A1(KEYINPUT43), .A2(n1299), .ZN(n1296) );
NAND2_X1 U1020 ( .A1(n1300), .A2(n1247), .ZN(n1299) );
XOR2_X1 U1021 ( .A(KEYINPUT46), .B(G101), .Z(n1300) );
NAND2_X1 U1022 ( .A1(n1301), .A2(n1302), .ZN(n1295) );
INV_X1 U1023 ( .A(KEYINPUT43), .ZN(n1302) );
NAND2_X1 U1024 ( .A1(n1303), .A2(n1304), .ZN(n1301) );
NAND2_X1 U1025 ( .A1(KEYINPUT46), .A2(n1249), .ZN(n1304) );
OR3_X1 U1026 ( .A1(n1298), .A2(KEYINPUT46), .A3(n1249), .ZN(n1303) );
INV_X1 U1027 ( .A(n1247), .ZN(n1298) );
XOR2_X1 U1028 ( .A(G104), .B(G107), .Z(n1247) );
XOR2_X1 U1029 ( .A(n1305), .B(n1248), .Z(n1292) );
XOR2_X1 U1030 ( .A(n1306), .B(n1167), .Z(n1290) );
NOR2_X1 U1031 ( .A1(n1101), .A2(G953), .ZN(n1167) );
INV_X1 U1032 ( .A(G224), .ZN(n1101) );
XNOR2_X1 U1033 ( .A(KEYINPUT47), .B(KEYINPUT17), .ZN(n1306) );
NOR2_X1 U1034 ( .A1(n1220), .A2(n1205), .ZN(n1012) );
XOR2_X1 U1035 ( .A(n1213), .B(KEYINPUT3), .Z(n1205) );
XOR2_X1 U1036 ( .A(n1307), .B(n1066), .Z(n1213) );
AND2_X1 U1037 ( .A1(G217), .A2(n1250), .ZN(n1066) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1288), .ZN(n1250) );
NAND2_X1 U1039 ( .A1(n1069), .A2(n1070), .ZN(n1307) );
XOR2_X1 U1040 ( .A(n1308), .B(n1309), .Z(n1069) );
XOR2_X1 U1041 ( .A(G140), .B(n1310), .Z(n1309) );
XOR2_X1 U1042 ( .A(KEYINPUT56), .B(G146), .Z(n1310) );
XOR2_X1 U1043 ( .A(n1311), .B(n1305), .Z(n1308) );
XNOR2_X1 U1044 ( .A(n1086), .B(n1162), .ZN(n1305) );
XOR2_X1 U1045 ( .A(G119), .B(G110), .Z(n1162) );
INV_X1 U1046 ( .A(G125), .ZN(n1086) );
XNOR2_X1 U1047 ( .A(G128), .B(n1312), .ZN(n1311) );
NOR2_X1 U1048 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U1049 ( .A(n1315), .B(KEYINPUT42), .Z(n1314) );
NAND2_X1 U1050 ( .A1(n1200), .A2(n1316), .ZN(n1315) );
NAND2_X1 U1051 ( .A1(n1283), .A2(G221), .ZN(n1316) );
INV_X1 U1052 ( .A(G137), .ZN(n1200) );
AND3_X1 U1053 ( .A1(n1283), .A2(G137), .A3(G221), .ZN(n1313) );
AND2_X1 U1054 ( .A1(G234), .A2(n1032), .ZN(n1283) );
INV_X1 U1055 ( .A(G953), .ZN(n1032) );
INV_X1 U1056 ( .A(n1206), .ZN(n1220) );
XOR2_X1 U1057 ( .A(n1317), .B(G472), .Z(n1206) );
NAND2_X1 U1058 ( .A1(KEYINPUT23), .A2(n1318), .ZN(n1317) );
INV_X1 U1059 ( .A(n1054), .ZN(n1318) );
NAND2_X1 U1060 ( .A1(n1319), .A2(n1070), .ZN(n1054) );
XOR2_X1 U1061 ( .A(n1288), .B(KEYINPUT54), .Z(n1070) );
INV_X1 U1062 ( .A(G902), .ZN(n1288) );
XOR2_X1 U1063 ( .A(n1320), .B(n1321), .Z(n1319) );
XNOR2_X1 U1064 ( .A(n1322), .B(n1323), .ZN(n1321) );
NOR2_X1 U1065 ( .A1(KEYINPUT34), .A2(n1142), .ZN(n1323) );
XOR2_X1 U1066 ( .A(n1219), .B(n1111), .Z(n1142) );
XOR2_X1 U1067 ( .A(G116), .B(G119), .Z(n1111) );
INV_X1 U1068 ( .A(G113), .ZN(n1219) );
NAND2_X1 U1069 ( .A1(KEYINPUT29), .A2(n1248), .ZN(n1322) );
XOR2_X1 U1070 ( .A(n1192), .B(n1279), .Z(n1248) );
XOR2_X1 U1071 ( .A(G128), .B(G143), .Z(n1279) );
INV_X1 U1072 ( .A(G146), .ZN(n1192) );
XOR2_X1 U1073 ( .A(n1087), .B(n1131), .Z(n1320) );
XOR2_X1 U1074 ( .A(n1324), .B(n1249), .Z(n1131) );
INV_X1 U1075 ( .A(G101), .ZN(n1249) );
NAND2_X1 U1076 ( .A1(G210), .A2(n1268), .ZN(n1324) );
NOR2_X1 U1077 ( .A1(G953), .A2(G237), .ZN(n1268) );
XNOR2_X1 U1078 ( .A(G131), .B(n1325), .ZN(n1087) );
XOR2_X1 U1079 ( .A(G137), .B(G134), .Z(n1325) );
endmodule


