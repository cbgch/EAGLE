//Key = 0001110100101001010100001011000101010111101100001010011011011111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379;

NAND2_X1 U750 ( .A1(n1041), .A2(n1042), .ZN(G9) );
NAND2_X1 U751 ( .A1(G107), .A2(n1043), .ZN(n1042) );
XOR2_X1 U752 ( .A(KEYINPUT27), .B(n1044), .Z(n1041) );
NOR2_X1 U753 ( .A1(G107), .A2(n1043), .ZN(n1044) );
NOR2_X1 U754 ( .A1(n1045), .A2(n1046), .ZN(G75) );
NOR2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND4_X1 U756 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
NAND2_X1 U757 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
XOR2_X1 U758 ( .A(n1055), .B(KEYINPUT28), .Z(n1049) );
NAND3_X1 U759 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NAND4_X1 U760 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1047) );
NAND3_X1 U761 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1060) );
XNOR2_X1 U762 ( .A(n1053), .B(KEYINPUT38), .ZN(n1065) );
AND2_X1 U763 ( .A1(n1058), .A2(n1066), .ZN(n1053) );
AND3_X1 U764 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1058) );
NAND3_X1 U765 ( .A1(n1056), .A2(n1070), .A3(n1069), .ZN(n1059) );
INV_X1 U766 ( .A(n1071), .ZN(n1069) );
NAND2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NAND3_X1 U768 ( .A1(n1074), .A2(n1068), .A3(n1067), .ZN(n1073) );
NAND2_X1 U769 ( .A1(n1066), .A2(n1075), .ZN(n1072) );
NAND2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U771 ( .A1(n1068), .A2(n1078), .ZN(n1077) );
XNOR2_X1 U772 ( .A(n1079), .B(n1080), .ZN(n1078) );
NAND2_X1 U773 ( .A1(n1067), .A2(n1081), .ZN(n1076) );
NAND2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR3_X1 U775 ( .A1(n1084), .A2(G953), .A3(G952), .ZN(n1045) );
INV_X1 U776 ( .A(n1061), .ZN(n1084) );
NAND4_X1 U777 ( .A1(n1085), .A2(n1067), .A3(n1086), .A4(n1087), .ZN(n1061) );
NOR4_X1 U778 ( .A1(n1063), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1087) );
XOR2_X1 U779 ( .A(n1091), .B(KEYINPUT63), .Z(n1090) );
XOR2_X1 U780 ( .A(n1092), .B(n1093), .Z(n1089) );
NAND2_X1 U781 ( .A1(KEYINPUT19), .A2(n1094), .ZN(n1092) );
NOR2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(n1088) );
NOR2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1086) );
XNOR2_X1 U784 ( .A(KEYINPUT20), .B(n1099), .ZN(n1098) );
XNOR2_X1 U785 ( .A(n1100), .B(n1101), .ZN(n1097) );
XNOR2_X1 U786 ( .A(KEYINPUT32), .B(n1102), .ZN(n1101) );
XOR2_X1 U787 ( .A(n1103), .B(n1104), .Z(G72) );
XOR2_X1 U788 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U789 ( .A1(n1107), .A2(n1062), .ZN(n1106) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XOR2_X1 U791 ( .A(KEYINPUT57), .B(G227), .Z(n1109) );
NAND2_X1 U792 ( .A1(n1110), .A2(n1111), .ZN(n1105) );
NAND2_X1 U793 ( .A1(G953), .A2(n1108), .ZN(n1111) );
XOR2_X1 U794 ( .A(n1112), .B(n1113), .Z(n1110) );
XOR2_X1 U795 ( .A(n1114), .B(n1115), .Z(n1113) );
XNOR2_X1 U796 ( .A(G131), .B(KEYINPUT6), .ZN(n1115) );
NAND2_X1 U797 ( .A1(KEYINPUT50), .A2(n1116), .ZN(n1114) );
XNOR2_X1 U798 ( .A(n1117), .B(n1118), .ZN(n1112) );
NAND2_X1 U799 ( .A1(n1062), .A2(n1119), .ZN(n1103) );
NAND2_X1 U800 ( .A1(n1120), .A2(n1121), .ZN(G69) );
NAND2_X1 U801 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XOR2_X1 U802 ( .A(n1124), .B(KEYINPUT11), .Z(n1122) );
XOR2_X1 U803 ( .A(KEYINPUT40), .B(n1125), .Z(n1120) );
NOR2_X1 U804 ( .A1(n1123), .A2(n1124), .ZN(n1125) );
XOR2_X1 U805 ( .A(n1126), .B(n1127), .Z(n1124) );
NOR2_X1 U806 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR2_X1 U807 ( .A1(G898), .A2(n1062), .ZN(n1128) );
NAND2_X1 U808 ( .A1(n1130), .A2(n1062), .ZN(n1126) );
AND2_X1 U809 ( .A1(G953), .A2(n1131), .ZN(n1123) );
NAND2_X1 U810 ( .A1(G898), .A2(G224), .ZN(n1131) );
NOR3_X1 U811 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(G66) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NOR2_X1 U813 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
AND2_X1 U814 ( .A1(KEYINPUT16), .A2(n1139), .ZN(n1138) );
NOR3_X1 U815 ( .A1(KEYINPUT16), .A2(KEYINPUT51), .A3(n1139), .ZN(n1137) );
NOR2_X1 U816 ( .A1(n1140), .A2(n1141), .ZN(n1133) );
NOR2_X1 U817 ( .A1(KEYINPUT51), .A2(n1139), .ZN(n1140) );
AND2_X1 U818 ( .A1(n1142), .A2(n1143), .ZN(n1139) );
NOR2_X1 U819 ( .A1(n1132), .A2(n1144), .ZN(G63) );
NOR3_X1 U820 ( .A1(n1093), .A2(n1145), .A3(n1146), .ZN(n1144) );
AND3_X1 U821 ( .A1(n1147), .A2(G478), .A3(n1142), .ZN(n1146) );
NOR2_X1 U822 ( .A1(n1148), .A2(n1147), .ZN(n1145) );
NOR2_X1 U823 ( .A1(n1149), .A2(n1094), .ZN(n1148) );
NOR2_X1 U824 ( .A1(n1119), .A2(n1130), .ZN(n1149) );
NOR2_X1 U825 ( .A1(n1132), .A2(n1150), .ZN(G60) );
XOR2_X1 U826 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U827 ( .A(KEYINPUT15), .B(n1153), .Z(n1152) );
NOR2_X1 U828 ( .A1(n1096), .A2(n1154), .ZN(n1153) );
XOR2_X1 U829 ( .A(G104), .B(n1155), .Z(G6) );
NOR2_X1 U830 ( .A1(n1132), .A2(n1156), .ZN(G57) );
XOR2_X1 U831 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U832 ( .A(n1159), .B(n1160), .Z(n1158) );
XNOR2_X1 U833 ( .A(n1161), .B(n1162), .ZN(n1160) );
NOR2_X1 U834 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U835 ( .A(KEYINPUT8), .B(n1165), .Z(n1164) );
NOR2_X1 U836 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U837 ( .A(n1168), .B(KEYINPUT56), .Z(n1166) );
NOR3_X1 U838 ( .A1(n1154), .A2(KEYINPUT25), .A3(n1102), .ZN(n1159) );
INV_X1 U839 ( .A(G472), .ZN(n1102) );
XNOR2_X1 U840 ( .A(n1169), .B(n1170), .ZN(n1157) );
NAND2_X1 U841 ( .A1(KEYINPUT35), .A2(n1171), .ZN(n1169) );
NOR2_X1 U842 ( .A1(n1132), .A2(n1172), .ZN(G54) );
XOR2_X1 U843 ( .A(n1173), .B(n1174), .Z(n1172) );
XNOR2_X1 U844 ( .A(n1175), .B(n1176), .ZN(n1174) );
AND2_X1 U845 ( .A1(G469), .A2(n1142), .ZN(n1176) );
XOR2_X1 U846 ( .A(n1177), .B(n1178), .Z(n1173) );
NOR2_X1 U847 ( .A1(KEYINPUT13), .A2(n1179), .ZN(n1178) );
NOR2_X1 U848 ( .A1(n1180), .A2(n1181), .ZN(G51) );
XOR2_X1 U849 ( .A(n1182), .B(n1183), .Z(n1181) );
XNOR2_X1 U850 ( .A(n1184), .B(n1185), .ZN(n1183) );
XNOR2_X1 U851 ( .A(n1186), .B(n1167), .ZN(n1182) );
NAND3_X1 U852 ( .A1(n1142), .A2(n1187), .A3(KEYINPUT37), .ZN(n1186) );
INV_X1 U853 ( .A(n1154), .ZN(n1142) );
NAND2_X1 U854 ( .A1(G902), .A2(n1188), .ZN(n1154) );
NAND2_X1 U855 ( .A1(n1050), .A2(n1051), .ZN(n1188) );
INV_X1 U856 ( .A(n1119), .ZN(n1051) );
NAND2_X1 U857 ( .A1(n1189), .A2(n1190), .ZN(n1119) );
AND4_X1 U858 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1190) );
NOR4_X1 U859 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1189) );
NOR3_X1 U860 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1198) );
NOR2_X1 U861 ( .A1(n1056), .A2(n1202), .ZN(n1201) );
AND3_X1 U862 ( .A1(KEYINPUT47), .A2(n1057), .A3(n1203), .ZN(n1202) );
NOR2_X1 U863 ( .A1(n1204), .A2(n1205), .ZN(n1200) );
NOR2_X1 U864 ( .A1(n1206), .A2(n1207), .ZN(n1204) );
XNOR2_X1 U865 ( .A(n1208), .B(KEYINPUT52), .ZN(n1206) );
NOR2_X1 U866 ( .A1(KEYINPUT47), .A2(n1209), .ZN(n1195) );
INV_X1 U867 ( .A(n1130), .ZN(n1050) );
NAND4_X1 U868 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1130) );
NOR4_X1 U869 ( .A1(n1214), .A2(n1215), .A3(n1155), .A4(n1216), .ZN(n1213) );
NOR4_X1 U870 ( .A1(n1217), .A2(n1082), .A3(n1218), .A4(n1219), .ZN(n1216) );
NAND3_X1 U871 ( .A1(n1080), .A2(n1079), .A3(n1220), .ZN(n1217) );
XNOR2_X1 U872 ( .A(KEYINPUT10), .B(n1221), .ZN(n1220) );
AND3_X1 U873 ( .A1(n1222), .A2(n1068), .A3(n1057), .ZN(n1155) );
INV_X1 U874 ( .A(n1223), .ZN(n1214) );
AND2_X1 U875 ( .A1(n1043), .A2(n1224), .ZN(n1212) );
NAND3_X1 U876 ( .A1(n1074), .A2(n1068), .A3(n1222), .ZN(n1043) );
XNOR2_X1 U877 ( .A(n1132), .B(KEYINPUT61), .ZN(n1180) );
NOR2_X1 U878 ( .A1(n1062), .A2(G952), .ZN(n1132) );
XOR2_X1 U879 ( .A(G146), .B(n1197), .Z(G48) );
AND3_X1 U880 ( .A1(n1057), .A2(n1054), .A3(n1225), .ZN(n1197) );
NAND2_X1 U881 ( .A1(n1226), .A2(n1227), .ZN(G45) );
NAND2_X1 U882 ( .A1(n1196), .A2(n1228), .ZN(n1227) );
XOR2_X1 U883 ( .A(n1229), .B(KEYINPUT0), .Z(n1226) );
OR2_X1 U884 ( .A1(n1228), .A2(n1196), .ZN(n1229) );
NOR4_X1 U885 ( .A1(n1199), .A2(n1230), .A3(n1083), .A4(n1218), .ZN(n1196) );
INV_X1 U886 ( .A(n1054), .ZN(n1218) );
XOR2_X1 U887 ( .A(n1209), .B(n1231), .Z(G42) );
NOR2_X1 U888 ( .A1(G140), .A2(KEYINPUT30), .ZN(n1231) );
OR4_X1 U889 ( .A1(n1205), .A2(n1199), .A3(n1082), .A4(n1232), .ZN(n1209) );
XNOR2_X1 U890 ( .A(G137), .B(n1194), .ZN(G39) );
NAND3_X1 U891 ( .A1(n1225), .A2(n1066), .A3(n1056), .ZN(n1194) );
XNOR2_X1 U892 ( .A(G134), .B(n1233), .ZN(G36) );
NAND3_X1 U893 ( .A1(n1234), .A2(KEYINPUT33), .A3(n1235), .ZN(n1233) );
NOR3_X1 U894 ( .A1(n1199), .A2(n1207), .A3(n1083), .ZN(n1235) );
INV_X1 U895 ( .A(n1074), .ZN(n1207) );
XNOR2_X1 U896 ( .A(n1056), .B(KEYINPUT7), .ZN(n1234) );
INV_X1 U897 ( .A(n1205), .ZN(n1056) );
XNOR2_X1 U898 ( .A(G131), .B(n1193), .ZN(G33) );
OR4_X1 U899 ( .A1(n1205), .A2(n1199), .A3(n1083), .A4(n1232), .ZN(n1193) );
NAND2_X1 U900 ( .A1(n1064), .A2(n1236), .ZN(n1205) );
XNOR2_X1 U901 ( .A(G128), .B(n1192), .ZN(G30) );
NAND3_X1 U902 ( .A1(n1074), .A2(n1054), .A3(n1225), .ZN(n1192) );
NOR3_X1 U903 ( .A1(n1237), .A2(n1099), .A3(n1199), .ZN(n1225) );
NAND3_X1 U904 ( .A1(n1238), .A2(n1079), .A3(n1080), .ZN(n1199) );
NAND3_X1 U905 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(G3) );
OR2_X1 U906 ( .A1(n1161), .A2(n1215), .ZN(n1241) );
NAND2_X1 U907 ( .A1(n1242), .A2(n1243), .ZN(n1240) );
INV_X1 U908 ( .A(KEYINPUT43), .ZN(n1243) );
NAND2_X1 U909 ( .A1(n1215), .A2(n1244), .ZN(n1242) );
XNOR2_X1 U910 ( .A(KEYINPUT5), .B(n1161), .ZN(n1244) );
NAND2_X1 U911 ( .A1(KEYINPUT43), .A2(n1245), .ZN(n1239) );
NAND2_X1 U912 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
OR2_X1 U913 ( .A1(n1161), .A2(KEYINPUT5), .ZN(n1247) );
NAND3_X1 U914 ( .A1(n1215), .A2(n1161), .A3(KEYINPUT5), .ZN(n1246) );
NOR3_X1 U915 ( .A1(n1083), .A2(n1248), .A3(n1219), .ZN(n1215) );
INV_X1 U916 ( .A(n1208), .ZN(n1083) );
XNOR2_X1 U917 ( .A(G125), .B(n1191), .ZN(G27) );
NAND4_X1 U918 ( .A1(n1054), .A2(n1238), .A3(n1067), .A4(n1249), .ZN(n1191) );
NOR2_X1 U919 ( .A1(n1232), .A2(n1082), .ZN(n1249) );
INV_X1 U920 ( .A(n1203), .ZN(n1082) );
NAND2_X1 U921 ( .A1(n1071), .A2(n1250), .ZN(n1238) );
NAND2_X1 U922 ( .A1(n1251), .A2(n1108), .ZN(n1250) );
INV_X1 U923 ( .A(G900), .ZN(n1108) );
XNOR2_X1 U924 ( .A(G122), .B(n1252), .ZN(G24) );
NOR2_X1 U925 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NOR4_X1 U926 ( .A1(n1255), .A2(n1256), .A3(n1230), .A4(n1221), .ZN(n1254) );
NAND3_X1 U927 ( .A1(n1068), .A2(n1054), .A3(n1067), .ZN(n1256) );
INV_X1 U928 ( .A(KEYINPUT36), .ZN(n1255) );
NOR2_X1 U929 ( .A1(KEYINPUT36), .A2(n1223), .ZN(n1253) );
NAND3_X1 U930 ( .A1(n1257), .A2(n1068), .A3(n1258), .ZN(n1223) );
INV_X1 U931 ( .A(n1230), .ZN(n1258) );
NAND2_X1 U932 ( .A1(n1259), .A2(n1260), .ZN(n1230) );
NOR2_X1 U933 ( .A1(n1261), .A2(n1262), .ZN(n1068) );
XNOR2_X1 U934 ( .A(G119), .B(n1210), .ZN(G21) );
NAND4_X1 U935 ( .A1(n1066), .A2(n1257), .A3(n1262), .A4(n1261), .ZN(n1210) );
XNOR2_X1 U936 ( .A(G116), .B(n1263), .ZN(G18) );
NAND2_X1 U937 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NAND2_X1 U938 ( .A1(KEYINPUT1), .A2(n1266), .ZN(n1265) );
OR2_X1 U939 ( .A1(KEYINPUT41), .A2(n1266), .ZN(n1264) );
INV_X1 U940 ( .A(n1211), .ZN(n1266) );
NAND3_X1 U941 ( .A1(n1257), .A2(n1074), .A3(n1208), .ZN(n1211) );
NOR2_X1 U942 ( .A1(n1260), .A2(n1267), .ZN(n1074) );
XOR2_X1 U943 ( .A(n1224), .B(n1268), .Z(G15) );
XOR2_X1 U944 ( .A(KEYINPUT59), .B(G113), .Z(n1268) );
NAND3_X1 U945 ( .A1(n1057), .A2(n1257), .A3(n1208), .ZN(n1224) );
NOR2_X1 U946 ( .A1(n1237), .A2(n1261), .ZN(n1208) );
AND3_X1 U947 ( .A1(n1054), .A2(n1221), .A3(n1067), .ZN(n1257) );
AND2_X1 U948 ( .A1(n1269), .A2(n1079), .ZN(n1067) );
INV_X1 U949 ( .A(n1080), .ZN(n1269) );
INV_X1 U950 ( .A(n1232), .ZN(n1057) );
NAND2_X1 U951 ( .A1(n1267), .A2(n1260), .ZN(n1232) );
NAND2_X1 U952 ( .A1(n1270), .A2(n1271), .ZN(G12) );
NAND4_X1 U953 ( .A1(n1272), .A2(n1273), .A3(n1203), .A4(n1274), .ZN(n1271) );
NOR2_X1 U954 ( .A1(n1248), .A2(n1219), .ZN(n1274) );
INV_X1 U955 ( .A(n1066), .ZN(n1219) );
NAND2_X1 U956 ( .A1(G110), .A2(n1275), .ZN(n1273) );
OR2_X1 U957 ( .A1(G110), .A2(KEYINPUT53), .ZN(n1272) );
NAND3_X1 U958 ( .A1(n1276), .A2(n1275), .A3(G110), .ZN(n1270) );
INV_X1 U959 ( .A(KEYINPUT9), .ZN(n1275) );
NAND4_X1 U960 ( .A1(KEYINPUT53), .A2(n1203), .A3(n1066), .A4(n1222), .ZN(n1276) );
INV_X1 U961 ( .A(n1248), .ZN(n1222) );
NAND4_X1 U962 ( .A1(n1054), .A2(n1080), .A3(n1221), .A4(n1079), .ZN(n1248) );
NAND2_X1 U963 ( .A1(G221), .A2(n1277), .ZN(n1079) );
NAND2_X1 U964 ( .A1(n1278), .A2(n1071), .ZN(n1221) );
NAND3_X1 U965 ( .A1(n1279), .A2(n1062), .A3(G952), .ZN(n1071) );
XOR2_X1 U966 ( .A(n1280), .B(KEYINPUT58), .Z(n1278) );
NAND2_X1 U967 ( .A1(n1251), .A2(n1281), .ZN(n1280) );
INV_X1 U968 ( .A(G898), .ZN(n1281) );
AND3_X1 U969 ( .A1(n1282), .A2(n1279), .A3(G953), .ZN(n1251) );
NAND2_X1 U970 ( .A1(G237), .A2(G234), .ZN(n1279) );
XNOR2_X1 U971 ( .A(KEYINPUT2), .B(n1283), .ZN(n1282) );
XNOR2_X1 U972 ( .A(n1284), .B(G469), .ZN(n1080) );
NAND2_X1 U973 ( .A1(n1285), .A2(n1283), .ZN(n1284) );
XNOR2_X1 U974 ( .A(n1286), .B(n1287), .ZN(n1285) );
INV_X1 U975 ( .A(n1175), .ZN(n1287) );
XNOR2_X1 U976 ( .A(n1288), .B(n1289), .ZN(n1175) );
XOR2_X1 U977 ( .A(n1290), .B(n1118), .Z(n1289) );
XNOR2_X1 U978 ( .A(n1291), .B(KEYINPUT17), .ZN(n1118) );
NOR2_X1 U979 ( .A1(KEYINPUT49), .A2(n1161), .ZN(n1290) );
XOR2_X1 U980 ( .A(n1168), .B(n1292), .Z(n1288) );
NOR2_X1 U981 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
AND2_X1 U982 ( .A1(n1295), .A2(G104), .ZN(n1293) );
NAND2_X1 U983 ( .A1(KEYINPUT24), .A2(n1296), .ZN(n1286) );
XOR2_X1 U984 ( .A(n1179), .B(n1297), .Z(n1296) );
XNOR2_X1 U985 ( .A(KEYINPUT4), .B(n1177), .ZN(n1297) );
NAND2_X1 U986 ( .A1(G227), .A2(n1062), .ZN(n1177) );
NOR2_X1 U987 ( .A1(n1064), .A2(n1063), .ZN(n1054) );
INV_X1 U988 ( .A(n1236), .ZN(n1063) );
NAND2_X1 U989 ( .A1(G214), .A2(n1298), .ZN(n1236) );
XNOR2_X1 U990 ( .A(n1085), .B(KEYINPUT26), .ZN(n1064) );
XOR2_X1 U991 ( .A(n1299), .B(n1187), .Z(n1085) );
AND2_X1 U992 ( .A1(G210), .A2(n1298), .ZN(n1187) );
NAND2_X1 U993 ( .A1(n1300), .A2(n1283), .ZN(n1298) );
NAND2_X1 U994 ( .A1(n1301), .A2(n1283), .ZN(n1299) );
XOR2_X1 U995 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U996 ( .A(n1185), .B(n1304), .ZN(n1303) );
XOR2_X1 U997 ( .A(n1129), .B(n1305), .Z(n1185) );
AND2_X1 U998 ( .A1(n1062), .A2(G224), .ZN(n1305) );
XOR2_X1 U999 ( .A(n1306), .B(n1307), .Z(n1129) );
XNOR2_X1 U1000 ( .A(n1308), .B(n1309), .ZN(n1307) );
NAND2_X1 U1001 ( .A1(n1310), .A2(n1311), .ZN(n1308) );
NAND2_X1 U1002 ( .A1(G116), .A2(n1312), .ZN(n1311) );
XOR2_X1 U1003 ( .A(KEYINPUT54), .B(n1313), .Z(n1310) );
NOR2_X1 U1004 ( .A1(G116), .A2(n1314), .ZN(n1313) );
XNOR2_X1 U1005 ( .A(KEYINPUT62), .B(n1312), .ZN(n1314) );
XOR2_X1 U1006 ( .A(n1315), .B(G110), .Z(n1306) );
NAND2_X1 U1007 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
NAND2_X1 U1008 ( .A1(n1318), .A2(n1161), .ZN(n1317) );
XOR2_X1 U1009 ( .A(KEYINPUT48), .B(n1319), .Z(n1316) );
NOR2_X1 U1010 ( .A1(n1318), .A2(n1161), .ZN(n1319) );
NOR2_X1 U1011 ( .A1(n1320), .A2(n1294), .ZN(n1318) );
NOR2_X1 U1012 ( .A1(n1295), .A2(G104), .ZN(n1294) );
XNOR2_X1 U1013 ( .A(n1321), .B(KEYINPUT55), .ZN(n1320) );
NAND2_X1 U1014 ( .A1(n1322), .A2(n1295), .ZN(n1321) );
XNOR2_X1 U1015 ( .A(G104), .B(KEYINPUT42), .ZN(n1322) );
XNOR2_X1 U1016 ( .A(KEYINPUT22), .B(n1323), .ZN(n1302) );
NOR2_X1 U1017 ( .A1(KEYINPUT34), .A2(n1167), .ZN(n1323) );
NOR2_X1 U1018 ( .A1(n1259), .A2(n1260), .ZN(n1066) );
NAND2_X1 U1019 ( .A1(n1091), .A2(n1324), .ZN(n1260) );
NAND2_X1 U1020 ( .A1(G475), .A2(n1325), .ZN(n1324) );
NAND2_X1 U1021 ( .A1(n1095), .A2(n1096), .ZN(n1091) );
INV_X1 U1022 ( .A(G475), .ZN(n1096) );
INV_X1 U1023 ( .A(n1325), .ZN(n1095) );
NAND2_X1 U1024 ( .A1(n1151), .A2(n1283), .ZN(n1325) );
NAND2_X1 U1025 ( .A1(n1326), .A2(n1327), .ZN(n1151) );
NAND2_X1 U1026 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
XNOR2_X1 U1027 ( .A(n1330), .B(n1331), .ZN(n1328) );
XNOR2_X1 U1028 ( .A(KEYINPUT45), .B(KEYINPUT12), .ZN(n1331) );
NAND2_X1 U1029 ( .A1(n1330), .A2(n1332), .ZN(n1326) );
INV_X1 U1030 ( .A(n1329), .ZN(n1332) );
XNOR2_X1 U1031 ( .A(G104), .B(n1309), .ZN(n1329) );
XOR2_X1 U1032 ( .A(G113), .B(G122), .Z(n1309) );
XNOR2_X1 U1033 ( .A(n1333), .B(n1334), .ZN(n1330) );
XNOR2_X1 U1034 ( .A(n1228), .B(G131), .ZN(n1334) );
XOR2_X1 U1035 ( .A(n1335), .B(n1336), .Z(n1333) );
AND3_X1 U1036 ( .A1(G214), .A2(n1062), .A3(n1300), .ZN(n1336) );
NAND2_X1 U1037 ( .A1(n1337), .A2(KEYINPUT3), .ZN(n1335) );
XOR2_X1 U1038 ( .A(n1116), .B(G146), .Z(n1337) );
XNOR2_X1 U1039 ( .A(G140), .B(n1184), .ZN(n1116) );
INV_X1 U1040 ( .A(n1267), .ZN(n1259) );
XOR2_X1 U1041 ( .A(n1093), .B(n1094), .Z(n1267) );
INV_X1 U1042 ( .A(G478), .ZN(n1094) );
NOR2_X1 U1043 ( .A1(n1147), .A2(G902), .ZN(n1093) );
XNOR2_X1 U1044 ( .A(n1338), .B(n1339), .ZN(n1147) );
XNOR2_X1 U1045 ( .A(n1340), .B(n1341), .ZN(n1339) );
XOR2_X1 U1046 ( .A(n1342), .B(n1343), .Z(n1341) );
AND3_X1 U1047 ( .A1(G217), .A2(n1062), .A3(G234), .ZN(n1343) );
NAND2_X1 U1048 ( .A1(KEYINPUT31), .A2(G134), .ZN(n1342) );
XOR2_X1 U1049 ( .A(n1344), .B(n1345), .Z(n1338) );
XNOR2_X1 U1050 ( .A(G116), .B(n1295), .ZN(n1345) );
INV_X1 U1051 ( .A(G107), .ZN(n1295) );
XNOR2_X1 U1052 ( .A(G122), .B(KEYINPUT39), .ZN(n1344) );
NOR2_X1 U1053 ( .A1(n1262), .A2(n1099), .ZN(n1203) );
INV_X1 U1054 ( .A(n1261), .ZN(n1099) );
XNOR2_X1 U1055 ( .A(n1346), .B(n1143), .ZN(n1261) );
AND2_X1 U1056 ( .A1(G217), .A2(n1277), .ZN(n1143) );
NAND2_X1 U1057 ( .A1(G234), .A2(n1283), .ZN(n1277) );
NAND2_X1 U1058 ( .A1(n1136), .A2(n1283), .ZN(n1346) );
INV_X1 U1059 ( .A(n1141), .ZN(n1136) );
XNOR2_X1 U1060 ( .A(n1347), .B(n1348), .ZN(n1141) );
XNOR2_X1 U1061 ( .A(n1179), .B(n1349), .ZN(n1348) );
XNOR2_X1 U1062 ( .A(n1350), .B(n1304), .ZN(n1349) );
INV_X1 U1063 ( .A(n1184), .ZN(n1304) );
XOR2_X1 U1064 ( .A(G125), .B(KEYINPUT46), .Z(n1184) );
NAND2_X1 U1065 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
NAND2_X1 U1066 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
INV_X1 U1067 ( .A(G128), .ZN(n1354) );
XOR2_X1 U1068 ( .A(n1355), .B(KEYINPUT14), .Z(n1351) );
NAND2_X1 U1069 ( .A1(n1312), .A2(G128), .ZN(n1355) );
INV_X1 U1070 ( .A(n1353), .ZN(n1312) );
XOR2_X1 U1071 ( .A(G140), .B(G110), .Z(n1179) );
XOR2_X1 U1072 ( .A(n1356), .B(n1357), .Z(n1347) );
XOR2_X1 U1073 ( .A(G146), .B(G137), .Z(n1357) );
NAND3_X1 U1074 ( .A1(G234), .A2(n1062), .A3(G221), .ZN(n1356) );
INV_X1 U1075 ( .A(n1237), .ZN(n1262) );
XNOR2_X1 U1076 ( .A(n1100), .B(n1358), .ZN(n1237) );
NOR2_X1 U1077 ( .A1(G472), .A2(KEYINPUT18), .ZN(n1358) );
NAND2_X1 U1078 ( .A1(n1359), .A2(n1283), .ZN(n1100) );
INV_X1 U1079 ( .A(G902), .ZN(n1283) );
XOR2_X1 U1080 ( .A(n1360), .B(n1361), .Z(n1359) );
XNOR2_X1 U1081 ( .A(n1171), .B(n1362), .ZN(n1361) );
NAND3_X1 U1082 ( .A1(n1363), .A2(n1364), .A3(n1365), .ZN(n1362) );
NAND2_X1 U1083 ( .A1(n1163), .A2(n1170), .ZN(n1365) );
NOR2_X1 U1084 ( .A1(n1168), .A2(n1291), .ZN(n1163) );
OR3_X1 U1085 ( .A1(n1170), .A2(n1167), .A3(n1168), .ZN(n1364) );
NAND2_X1 U1086 ( .A1(n1366), .A2(n1168), .ZN(n1363) );
NAND3_X1 U1087 ( .A1(n1367), .A2(n1368), .A3(n1369), .ZN(n1168) );
NAND2_X1 U1088 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
NAND2_X1 U1089 ( .A1(KEYINPUT44), .A2(n1372), .ZN(n1368) );
NAND2_X1 U1090 ( .A1(n1373), .A2(n1117), .ZN(n1372) );
XNOR2_X1 U1091 ( .A(KEYINPUT29), .B(n1371), .ZN(n1373) );
NAND2_X1 U1092 ( .A1(n1374), .A2(n1375), .ZN(n1367) );
INV_X1 U1093 ( .A(KEYINPUT44), .ZN(n1375) );
NAND2_X1 U1094 ( .A1(n1376), .A2(n1377), .ZN(n1374) );
NAND2_X1 U1095 ( .A1(KEYINPUT29), .A2(n1371), .ZN(n1377) );
OR3_X1 U1096 ( .A1(n1370), .A2(KEYINPUT29), .A3(n1371), .ZN(n1376) );
INV_X1 U1097 ( .A(G131), .ZN(n1371) );
INV_X1 U1098 ( .A(n1117), .ZN(n1370) );
XOR2_X1 U1099 ( .A(G134), .B(G137), .Z(n1117) );
XNOR2_X1 U1100 ( .A(n1170), .B(n1291), .ZN(n1366) );
INV_X1 U1101 ( .A(n1167), .ZN(n1291) );
XOR2_X1 U1102 ( .A(G146), .B(n1340), .Z(n1167) );
XNOR2_X1 U1103 ( .A(G128), .B(n1228), .ZN(n1340) );
INV_X1 U1104 ( .A(G143), .ZN(n1228) );
XOR2_X1 U1105 ( .A(n1378), .B(n1379), .Z(n1170) );
XOR2_X1 U1106 ( .A(G116), .B(G113), .Z(n1379) );
NAND2_X1 U1107 ( .A1(KEYINPUT60), .A2(n1353), .ZN(n1378) );
XOR2_X1 U1108 ( .A(G119), .B(KEYINPUT23), .Z(n1353) );
AND3_X1 U1109 ( .A1(n1300), .A2(n1062), .A3(G210), .ZN(n1171) );
INV_X1 U1110 ( .A(G953), .ZN(n1062) );
INV_X1 U1111 ( .A(G237), .ZN(n1300) );
XNOR2_X1 U1112 ( .A(KEYINPUT21), .B(n1161), .ZN(n1360) );
INV_X1 U1113 ( .A(G101), .ZN(n1161) );
endmodule


