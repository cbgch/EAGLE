//Key = 1110010011100010011010110001100010100011100010000011000000001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368;

XOR2_X1 U761 ( .A(n1037), .B(n1038), .Z(G9) );
NOR2_X1 U762 ( .A1(n1039), .A2(n1040), .ZN(G75) );
NOR4_X1 U763 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1040) );
NOR3_X1 U764 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1043) );
NOR2_X1 U765 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U766 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U767 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U768 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U769 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U770 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U771 ( .A1(n1060), .A2(n1061), .ZN(n1052) );
NOR2_X1 U772 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
AND2_X1 U773 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR3_X1 U774 ( .A1(n1061), .A2(n1066), .A3(n1055), .ZN(n1048) );
NOR2_X1 U775 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND3_X1 U776 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1041) );
NAND3_X1 U777 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
NOR3_X1 U778 ( .A1(n1055), .A2(n1075), .A3(n1051), .ZN(n1074) );
NOR2_X1 U779 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U780 ( .A(KEYINPUT36), .B(n1078), .Z(n1077) );
INV_X1 U781 ( .A(n1045), .ZN(n1072) );
NOR3_X1 U782 ( .A1(n1079), .A2(G953), .A3(G952), .ZN(n1039) );
INV_X1 U783 ( .A(n1069), .ZN(n1079) );
NAND4_X1 U784 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1069) );
NOR3_X1 U785 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1083) );
NOR2_X1 U786 ( .A1(KEYINPUT32), .A2(n1087), .ZN(n1085) );
NAND3_X1 U787 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1084) );
XNOR2_X1 U788 ( .A(n1091), .B(G472), .ZN(n1090) );
NAND3_X1 U789 ( .A1(KEYINPUT32), .A2(n1087), .A3(G475), .ZN(n1089) );
NAND2_X1 U790 ( .A1(n1092), .A2(n1093), .ZN(n1088) );
NAND2_X1 U791 ( .A1(KEYINPUT32), .A2(n1094), .ZN(n1092) );
XOR2_X1 U792 ( .A(KEYINPUT8), .B(n1095), .Z(n1094) );
NOR3_X1 U793 ( .A1(n1096), .A2(n1065), .A3(n1097), .ZN(n1082) );
XNOR2_X1 U794 ( .A(n1098), .B(n1099), .ZN(n1096) );
NAND2_X1 U795 ( .A1(KEYINPUT23), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U796 ( .A(n1101), .B(n1102), .ZN(n1081) );
NOR2_X1 U797 ( .A1(G469), .A2(KEYINPUT35), .ZN(n1102) );
XNOR2_X1 U798 ( .A(n1103), .B(n1104), .ZN(n1080) );
XOR2_X1 U799 ( .A(KEYINPUT34), .B(n1105), .Z(n1104) );
XOR2_X1 U800 ( .A(n1106), .B(n1107), .Z(G72) );
NOR2_X1 U801 ( .A1(n1108), .A2(n1070), .ZN(n1107) );
NOR2_X1 U802 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U803 ( .A1(KEYINPUT48), .A2(n1111), .ZN(n1106) );
XOR2_X1 U804 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U805 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U806 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U807 ( .A(n1118), .B(n1119), .Z(n1117) );
XNOR2_X1 U808 ( .A(KEYINPUT51), .B(KEYINPUT19), .ZN(n1119) );
XNOR2_X1 U809 ( .A(n1120), .B(n1121), .ZN(n1116) );
XOR2_X1 U810 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U811 ( .A1(KEYINPUT52), .A2(n1124), .ZN(n1122) );
NOR2_X1 U812 ( .A1(G900), .A2(n1070), .ZN(n1114) );
NAND2_X1 U813 ( .A1(n1070), .A2(n1044), .ZN(n1112) );
NAND2_X1 U814 ( .A1(n1125), .A2(n1126), .ZN(G69) );
NAND2_X1 U815 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
INV_X1 U816 ( .A(n1129), .ZN(n1127) );
NAND2_X1 U817 ( .A1(n1129), .A2(n1130), .ZN(n1125) );
NAND2_X1 U818 ( .A1(n1131), .A2(n1128), .ZN(n1130) );
NAND2_X1 U819 ( .A1(G953), .A2(n1132), .ZN(n1128) );
INV_X1 U820 ( .A(G224), .ZN(n1132) );
XOR2_X1 U821 ( .A(n1133), .B(n1134), .Z(n1129) );
NOR2_X1 U822 ( .A1(G953), .A2(n1135), .ZN(n1134) );
XNOR2_X1 U823 ( .A(KEYINPUT46), .B(n1042), .ZN(n1135) );
NAND2_X1 U824 ( .A1(n1136), .A2(n1131), .ZN(n1133) );
INV_X1 U825 ( .A(n1137), .ZN(n1131) );
XOR2_X1 U826 ( .A(n1138), .B(n1139), .Z(n1136) );
NOR4_X1 U827 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(G66) );
NOR3_X1 U828 ( .A1(n1144), .A2(G953), .A3(G952), .ZN(n1143) );
AND2_X1 U829 ( .A1(n1144), .A2(n1145), .ZN(n1142) );
INV_X1 U830 ( .A(KEYINPUT7), .ZN(n1144) );
NOR2_X1 U831 ( .A1(n1146), .A2(n1147), .ZN(n1141) );
NOR2_X1 U832 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NOR3_X1 U833 ( .A1(n1150), .A2(KEYINPUT37), .A3(KEYINPUT24), .ZN(n1149) );
AND2_X1 U834 ( .A1(n1150), .A2(KEYINPUT37), .ZN(n1148) );
NOR2_X1 U835 ( .A1(n1151), .A2(n1152), .ZN(n1140) );
NOR2_X1 U836 ( .A1(KEYINPUT24), .A2(n1150), .ZN(n1151) );
OR2_X1 U837 ( .A1(n1153), .A2(n1103), .ZN(n1150) );
NOR2_X1 U838 ( .A1(n1145), .A2(n1154), .ZN(G63) );
XOR2_X1 U839 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND2_X1 U840 ( .A1(n1157), .A2(G478), .ZN(n1155) );
NOR2_X1 U841 ( .A1(n1145), .A2(n1158), .ZN(G60) );
NOR3_X1 U842 ( .A1(n1095), .A2(n1159), .A3(n1160), .ZN(n1158) );
AND3_X1 U843 ( .A1(n1161), .A2(G475), .A3(n1157), .ZN(n1160) );
NOR2_X1 U844 ( .A1(n1162), .A2(n1161), .ZN(n1159) );
NOR2_X1 U845 ( .A1(n1163), .A2(n1093), .ZN(n1162) );
NOR2_X1 U846 ( .A1(n1044), .A2(n1042), .ZN(n1163) );
XNOR2_X1 U847 ( .A(G104), .B(n1164), .ZN(G6) );
NOR2_X1 U848 ( .A1(n1145), .A2(n1165), .ZN(G57) );
XOR2_X1 U849 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U850 ( .A(n1168), .B(n1169), .Z(n1166) );
NOR2_X1 U851 ( .A1(KEYINPUT21), .A2(n1170), .ZN(n1169) );
NAND2_X1 U852 ( .A1(n1157), .A2(G472), .ZN(n1168) );
NOR2_X1 U853 ( .A1(n1171), .A2(n1172), .ZN(G54) );
XOR2_X1 U854 ( .A(n1173), .B(KEYINPUT2), .Z(n1172) );
NAND2_X1 U855 ( .A1(G953), .A2(n1174), .ZN(n1173) );
XOR2_X1 U856 ( .A(KEYINPUT0), .B(G952), .Z(n1174) );
XOR2_X1 U857 ( .A(n1175), .B(n1176), .Z(n1171) );
XNOR2_X1 U858 ( .A(n1177), .B(n1178), .ZN(n1176) );
XOR2_X1 U859 ( .A(n1179), .B(n1180), .Z(n1175) );
NOR2_X1 U860 ( .A1(KEYINPUT61), .A2(n1181), .ZN(n1180) );
NAND2_X1 U861 ( .A1(n1157), .A2(G469), .ZN(n1179) );
INV_X1 U862 ( .A(n1153), .ZN(n1157) );
NOR2_X1 U863 ( .A1(n1145), .A2(n1182), .ZN(G51) );
XOR2_X1 U864 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U865 ( .A(G125), .B(n1185), .Z(n1184) );
NOR2_X1 U866 ( .A1(n1186), .A2(KEYINPUT3), .ZN(n1185) );
NOR2_X1 U867 ( .A1(n1100), .A2(n1153), .ZN(n1186) );
NAND2_X1 U868 ( .A1(G902), .A2(n1187), .ZN(n1153) );
OR2_X1 U869 ( .A1(n1042), .A2(n1044), .ZN(n1187) );
NAND4_X1 U870 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1044) );
NOR4_X1 U871 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
NAND2_X1 U872 ( .A1(n1196), .A2(n1197), .ZN(n1190) );
INV_X1 U873 ( .A(KEYINPUT45), .ZN(n1197) );
NAND2_X1 U874 ( .A1(n1073), .A2(n1198), .ZN(n1189) );
NAND2_X1 U875 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND2_X1 U876 ( .A1(KEYINPUT45), .A2(n1201), .ZN(n1200) );
XNOR2_X1 U877 ( .A(n1202), .B(KEYINPUT31), .ZN(n1199) );
NAND2_X1 U878 ( .A1(n1057), .A2(n1203), .ZN(n1188) );
NAND2_X1 U879 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
XOR2_X1 U880 ( .A(n1206), .B(KEYINPUT33), .Z(n1204) );
NAND4_X1 U881 ( .A1(n1207), .A2(n1164), .A3(n1208), .A4(n1209), .ZN(n1042) );
AND4_X1 U882 ( .A1(n1038), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1209) );
NAND3_X1 U883 ( .A1(n1213), .A2(n1214), .A3(n1067), .ZN(n1038) );
NOR3_X1 U884 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1208) );
NOR3_X1 U885 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1217) );
NOR4_X1 U886 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1219) );
XOR2_X1 U887 ( .A(n1225), .B(n1055), .Z(n1224) );
INV_X1 U888 ( .A(KEYINPUT26), .ZN(n1218) );
NOR4_X1 U889 ( .A1(KEYINPUT26), .A2(n1223), .A3(n1226), .A4(n1227), .ZN(n1216) );
NOR2_X1 U890 ( .A1(KEYINPUT39), .A2(n1228), .ZN(n1227) );
NOR3_X1 U891 ( .A1(n1222), .A2(n1229), .A3(n1230), .ZN(n1228) );
NOR2_X1 U892 ( .A1(n1231), .A2(n1225), .ZN(n1226) );
INV_X1 U893 ( .A(KEYINPUT39), .ZN(n1225) );
AND2_X1 U894 ( .A1(n1067), .A2(n1231), .ZN(n1215) );
NAND3_X1 U895 ( .A1(n1213), .A2(n1214), .A3(n1068), .ZN(n1164) );
NAND2_X1 U896 ( .A1(n1232), .A2(n1229), .ZN(n1207) );
NOR2_X1 U897 ( .A1(n1070), .A2(G952), .ZN(n1145) );
XOR2_X1 U898 ( .A(G146), .B(n1195), .Z(G48) );
AND3_X1 U899 ( .A1(n1068), .A2(n1057), .A3(n1233), .ZN(n1195) );
XOR2_X1 U900 ( .A(G143), .B(n1234), .Z(G45) );
NOR3_X1 U901 ( .A1(n1205), .A2(KEYINPUT25), .A3(n1220), .ZN(n1234) );
NAND4_X1 U902 ( .A1(n1235), .A2(n1076), .A3(n1086), .A4(n1236), .ZN(n1205) );
XOR2_X1 U903 ( .A(G140), .B(n1194), .Z(G42) );
AND4_X1 U904 ( .A1(n1073), .A2(n1235), .A3(n1068), .A4(n1078), .ZN(n1194) );
XOR2_X1 U905 ( .A(n1237), .B(n1238), .Z(G39) );
XNOR2_X1 U906 ( .A(G137), .B(KEYINPUT55), .ZN(n1238) );
NAND2_X1 U907 ( .A1(n1202), .A2(n1073), .ZN(n1237) );
AND2_X1 U908 ( .A1(n1233), .A2(n1239), .ZN(n1202) );
XOR2_X1 U909 ( .A(G134), .B(n1193), .Z(G36) );
AND4_X1 U910 ( .A1(n1073), .A2(n1235), .A3(n1076), .A4(n1067), .ZN(n1193) );
NAND2_X1 U911 ( .A1(n1240), .A2(n1241), .ZN(G33) );
NAND2_X1 U912 ( .A1(n1242), .A2(n1118), .ZN(n1241) );
INV_X1 U913 ( .A(G131), .ZN(n1118) );
XOR2_X1 U914 ( .A(KEYINPUT57), .B(n1196), .Z(n1242) );
NAND2_X1 U915 ( .A1(n1243), .A2(G131), .ZN(n1240) );
XOR2_X1 U916 ( .A(KEYINPUT5), .B(n1196), .Z(n1243) );
NOR2_X1 U917 ( .A1(n1201), .A2(n1061), .ZN(n1196) );
INV_X1 U918 ( .A(n1073), .ZN(n1061) );
NOR2_X1 U919 ( .A1(n1058), .A2(n1097), .ZN(n1073) );
INV_X1 U920 ( .A(n1059), .ZN(n1097) );
NAND3_X1 U921 ( .A1(n1068), .A2(n1076), .A3(n1235), .ZN(n1201) );
XOR2_X1 U922 ( .A(G128), .B(n1192), .Z(G30) );
AND3_X1 U923 ( .A1(n1067), .A2(n1057), .A3(n1233), .ZN(n1192) );
AND3_X1 U924 ( .A1(n1244), .A2(n1245), .A3(n1235), .ZN(n1233) );
AND2_X1 U925 ( .A1(n1063), .A2(n1246), .ZN(n1235) );
INV_X1 U926 ( .A(n1220), .ZN(n1057) );
XOR2_X1 U927 ( .A(n1247), .B(n1212), .Z(G3) );
NAND3_X1 U928 ( .A1(n1239), .A2(n1214), .A3(n1076), .ZN(n1212) );
XOR2_X1 U929 ( .A(G125), .B(n1248), .Z(G27) );
NOR2_X1 U930 ( .A1(n1220), .A2(n1206), .ZN(n1248) );
NAND4_X1 U931 ( .A1(n1068), .A2(n1229), .A3(n1078), .A4(n1246), .ZN(n1206) );
NAND2_X1 U932 ( .A1(n1045), .A2(n1249), .ZN(n1246) );
NAND4_X1 U933 ( .A1(G902), .A2(G953), .A3(n1250), .A4(n1110), .ZN(n1249) );
INV_X1 U934 ( .A(G900), .ZN(n1110) );
INV_X1 U935 ( .A(n1055), .ZN(n1229) );
XOR2_X1 U936 ( .A(n1251), .B(n1252), .Z(G24) );
NAND2_X1 U937 ( .A1(n1253), .A2(n1232), .ZN(n1252) );
NOR4_X1 U938 ( .A1(n1047), .A2(n1230), .A3(n1254), .A4(n1255), .ZN(n1232) );
INV_X1 U939 ( .A(n1213), .ZN(n1047) );
NOR2_X1 U940 ( .A1(n1245), .A2(n1244), .ZN(n1213) );
XOR2_X1 U941 ( .A(n1055), .B(KEYINPUT28), .Z(n1253) );
NAND3_X1 U942 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(G21) );
OR2_X1 U943 ( .A1(n1211), .A2(G119), .ZN(n1258) );
NAND2_X1 U944 ( .A1(KEYINPUT41), .A2(n1259), .ZN(n1257) );
NAND2_X1 U945 ( .A1(G119), .A2(n1260), .ZN(n1259) );
XNOR2_X1 U946 ( .A(KEYINPUT60), .B(n1211), .ZN(n1260) );
NAND2_X1 U947 ( .A1(n1261), .A2(n1262), .ZN(n1256) );
INV_X1 U948 ( .A(KEYINPUT41), .ZN(n1262) );
NAND2_X1 U949 ( .A1(n1263), .A2(n1264), .ZN(n1261) );
OR2_X1 U950 ( .A1(n1211), .A2(KEYINPUT60), .ZN(n1264) );
NAND3_X1 U951 ( .A1(G119), .A2(n1211), .A3(KEYINPUT60), .ZN(n1263) );
NAND4_X1 U952 ( .A1(n1265), .A2(n1245), .A3(n1239), .A4(n1266), .ZN(n1211) );
NOR2_X1 U953 ( .A1(n1055), .A2(n1267), .ZN(n1266) );
XNOR2_X1 U954 ( .A(G116), .B(n1268), .ZN(G18) );
NAND3_X1 U955 ( .A1(n1231), .A2(n1067), .A3(KEYINPUT22), .ZN(n1268) );
NOR2_X1 U956 ( .A1(n1236), .A2(n1254), .ZN(n1067) );
NAND3_X1 U957 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(G15) );
NAND3_X1 U958 ( .A1(n1068), .A2(n1272), .A3(n1231), .ZN(n1271) );
NAND2_X1 U959 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U960 ( .A1(KEYINPUT50), .A2(n1275), .ZN(n1274) );
NAND2_X1 U961 ( .A1(KEYINPUT47), .A2(n1275), .ZN(n1270) );
NAND3_X1 U962 ( .A1(n1276), .A2(n1273), .A3(G113), .ZN(n1269) );
INV_X1 U963 ( .A(KEYINPUT47), .ZN(n1273) );
NAND3_X1 U964 ( .A1(n1231), .A2(n1068), .A3(KEYINPUT50), .ZN(n1276) );
INV_X1 U965 ( .A(n1223), .ZN(n1068) );
NAND2_X1 U966 ( .A1(n1277), .A2(n1236), .ZN(n1223) );
INV_X1 U967 ( .A(n1255), .ZN(n1236) );
NOR3_X1 U968 ( .A1(n1055), .A2(n1230), .A3(n1222), .ZN(n1231) );
INV_X1 U969 ( .A(n1076), .ZN(n1222) );
NOR2_X1 U970 ( .A1(n1267), .A2(n1245), .ZN(n1076) );
INV_X1 U971 ( .A(n1265), .ZN(n1230) );
NAND2_X1 U972 ( .A1(n1064), .A2(n1278), .ZN(n1055) );
XNOR2_X1 U973 ( .A(G110), .B(n1210), .ZN(G12) );
NAND3_X1 U974 ( .A1(n1078), .A2(n1214), .A3(n1239), .ZN(n1210) );
INV_X1 U975 ( .A(n1051), .ZN(n1239) );
NAND2_X1 U976 ( .A1(n1255), .A2(n1277), .ZN(n1051) );
XOR2_X1 U977 ( .A(n1086), .B(KEYINPUT20), .Z(n1277) );
INV_X1 U978 ( .A(n1254), .ZN(n1086) );
XOR2_X1 U979 ( .A(n1279), .B(G478), .Z(n1254) );
NAND2_X1 U980 ( .A1(n1156), .A2(n1280), .ZN(n1279) );
XNOR2_X1 U981 ( .A(n1281), .B(n1282), .ZN(n1156) );
XOR2_X1 U982 ( .A(n1283), .B(n1284), .Z(n1282) );
NAND2_X1 U983 ( .A1(G217), .A2(n1285), .ZN(n1284) );
NAND2_X1 U984 ( .A1(n1286), .A2(n1287), .ZN(n1283) );
NAND2_X1 U985 ( .A1(n1288), .A2(n1037), .ZN(n1287) );
XOR2_X1 U986 ( .A(n1289), .B(KEYINPUT53), .Z(n1286) );
OR2_X1 U987 ( .A1(n1037), .A2(n1288), .ZN(n1289) );
XNOR2_X1 U988 ( .A(n1251), .B(n1290), .ZN(n1288) );
NOR2_X1 U989 ( .A1(KEYINPUT63), .A2(n1291), .ZN(n1290) );
XNOR2_X1 U990 ( .A(G116), .B(KEYINPUT44), .ZN(n1291) );
XOR2_X1 U991 ( .A(n1292), .B(n1293), .Z(n1281) );
XOR2_X1 U992 ( .A(G143), .B(G134), .Z(n1293) );
XNOR2_X1 U993 ( .A(n1087), .B(n1093), .ZN(n1255) );
INV_X1 U994 ( .A(G475), .ZN(n1093) );
INV_X1 U995 ( .A(n1095), .ZN(n1087) );
NOR2_X1 U996 ( .A1(n1161), .A2(G902), .ZN(n1095) );
XNOR2_X1 U997 ( .A(n1294), .B(n1295), .ZN(n1161) );
XOR2_X1 U998 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U999 ( .A(G122), .B(G113), .Z(n1297) );
XOR2_X1 U1000 ( .A(G143), .B(G131), .Z(n1296) );
XOR2_X1 U1001 ( .A(n1298), .B(n1299), .Z(n1294) );
XNOR2_X1 U1002 ( .A(G104), .B(n1300), .ZN(n1299) );
NAND2_X1 U1003 ( .A1(G214), .A2(n1301), .ZN(n1300) );
NAND2_X1 U1004 ( .A1(KEYINPUT1), .A2(n1302), .ZN(n1298) );
AND2_X1 U1005 ( .A1(n1063), .A2(n1265), .ZN(n1214) );
NOR2_X1 U1006 ( .A1(n1220), .A2(n1221), .ZN(n1265) );
AND2_X1 U1007 ( .A1(n1045), .A2(n1303), .ZN(n1221) );
NAND3_X1 U1008 ( .A1(n1137), .A2(n1250), .A3(G902), .ZN(n1303) );
NOR2_X1 U1009 ( .A1(G898), .A2(n1070), .ZN(n1137) );
NAND3_X1 U1010 ( .A1(n1250), .A2(n1070), .A3(G952), .ZN(n1045) );
NAND2_X1 U1011 ( .A1(G237), .A2(G234), .ZN(n1250) );
NAND2_X1 U1012 ( .A1(n1058), .A2(n1059), .ZN(n1220) );
NAND2_X1 U1013 ( .A1(G214), .A2(n1304), .ZN(n1059) );
XOR2_X1 U1014 ( .A(n1099), .B(n1100), .Z(n1058) );
NAND2_X1 U1015 ( .A1(G210), .A2(n1304), .ZN(n1100) );
NAND2_X1 U1016 ( .A1(n1305), .A2(n1280), .ZN(n1304) );
INV_X1 U1017 ( .A(G237), .ZN(n1305) );
NAND2_X1 U1018 ( .A1(n1306), .A2(n1280), .ZN(n1099) );
XNOR2_X1 U1019 ( .A(n1183), .B(n1307), .ZN(n1306) );
NOR2_X1 U1020 ( .A1(G125), .A2(KEYINPUT42), .ZN(n1307) );
XNOR2_X1 U1021 ( .A(n1308), .B(n1309), .ZN(n1183) );
XOR2_X1 U1022 ( .A(n1138), .B(n1310), .Z(n1309) );
XNOR2_X1 U1023 ( .A(n1311), .B(n1312), .ZN(n1138) );
XOR2_X1 U1024 ( .A(n1313), .B(n1314), .Z(n1312) );
NOR2_X1 U1025 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
AND3_X1 U1026 ( .A1(KEYINPUT13), .A2(n1037), .A3(G104), .ZN(n1316) );
INV_X1 U1027 ( .A(G107), .ZN(n1037) );
NOR2_X1 U1028 ( .A1(KEYINPUT13), .A2(n1317), .ZN(n1315) );
NOR2_X1 U1029 ( .A1(G101), .A2(KEYINPUT58), .ZN(n1313) );
XOR2_X1 U1030 ( .A(G110), .B(n1251), .Z(n1311) );
INV_X1 U1031 ( .A(G122), .ZN(n1251) );
XOR2_X1 U1032 ( .A(n1318), .B(KEYINPUT16), .Z(n1308) );
NAND2_X1 U1033 ( .A1(G224), .A2(n1070), .ZN(n1318) );
NOR2_X1 U1034 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
INV_X1 U1035 ( .A(n1278), .ZN(n1065) );
NAND2_X1 U1036 ( .A1(G221), .A2(n1319), .ZN(n1278) );
XOR2_X1 U1037 ( .A(n1101), .B(G469), .Z(n1064) );
NAND2_X1 U1038 ( .A1(n1320), .A2(n1280), .ZN(n1101) );
XOR2_X1 U1039 ( .A(n1321), .B(n1322), .Z(n1320) );
NOR2_X1 U1040 ( .A1(KEYINPUT4), .A2(n1323), .ZN(n1322) );
XNOR2_X1 U1041 ( .A(n1177), .B(KEYINPUT10), .ZN(n1323) );
XNOR2_X1 U1042 ( .A(n1324), .B(n1325), .ZN(n1177) );
XOR2_X1 U1043 ( .A(G110), .B(n1326), .Z(n1325) );
NOR2_X1 U1044 ( .A1(G953), .A2(n1109), .ZN(n1326) );
INV_X1 U1045 ( .A(G227), .ZN(n1109) );
XNOR2_X1 U1046 ( .A(G140), .B(KEYINPUT14), .ZN(n1324) );
NOR2_X1 U1047 ( .A1(n1327), .A2(n1328), .ZN(n1321) );
XOR2_X1 U1048 ( .A(n1329), .B(KEYINPUT38), .Z(n1328) );
NAND2_X1 U1049 ( .A1(n1178), .A2(n1330), .ZN(n1329) );
NOR2_X1 U1050 ( .A1(n1178), .A2(n1330), .ZN(n1327) );
XNOR2_X1 U1051 ( .A(KEYINPUT12), .B(n1181), .ZN(n1330) );
XNOR2_X1 U1052 ( .A(n1124), .B(n1331), .ZN(n1181) );
XOR2_X1 U1053 ( .A(G101), .B(n1317), .Z(n1331) );
XOR2_X1 U1054 ( .A(G104), .B(G107), .Z(n1317) );
XNOR2_X1 U1055 ( .A(n1332), .B(KEYINPUT27), .ZN(n1124) );
NAND2_X1 U1056 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
NAND2_X1 U1057 ( .A1(G128), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1058 ( .A(KEYINPUT17), .B(n1336), .Z(n1333) );
NOR2_X1 U1059 ( .A1(G128), .A2(n1335), .ZN(n1336) );
NAND3_X1 U1060 ( .A1(n1337), .A2(n1338), .A3(n1339), .ZN(n1335) );
NAND2_X1 U1061 ( .A1(KEYINPUT15), .A2(n1340), .ZN(n1339) );
NAND3_X1 U1062 ( .A1(n1341), .A2(n1342), .A3(G146), .ZN(n1338) );
NAND2_X1 U1063 ( .A1(n1343), .A2(n1344), .ZN(n1337) );
NAND2_X1 U1064 ( .A1(n1345), .A2(n1342), .ZN(n1343) );
INV_X1 U1065 ( .A(KEYINPUT15), .ZN(n1342) );
XOR2_X1 U1066 ( .A(KEYINPUT29), .B(n1341), .Z(n1345) );
INV_X1 U1067 ( .A(n1340), .ZN(n1341) );
XNOR2_X1 U1068 ( .A(G143), .B(KEYINPUT40), .ZN(n1340) );
AND2_X1 U1069 ( .A1(n1267), .A2(n1245), .ZN(n1078) );
XOR2_X1 U1070 ( .A(n1105), .B(n1346), .Z(n1245) );
NOR2_X1 U1071 ( .A1(KEYINPUT59), .A2(n1103), .ZN(n1346) );
NAND2_X1 U1072 ( .A1(G217), .A2(n1319), .ZN(n1103) );
NAND2_X1 U1073 ( .A1(G234), .A2(n1280), .ZN(n1319) );
NOR2_X1 U1074 ( .A1(n1146), .A2(G902), .ZN(n1105) );
INV_X1 U1075 ( .A(n1152), .ZN(n1146) );
XOR2_X1 U1076 ( .A(n1347), .B(n1348), .Z(n1152) );
XOR2_X1 U1077 ( .A(G110), .B(n1349), .Z(n1348) );
NOR2_X1 U1078 ( .A1(KEYINPUT11), .A2(n1350), .ZN(n1349) );
XOR2_X1 U1079 ( .A(n1351), .B(n1352), .Z(n1350) );
NOR2_X1 U1080 ( .A1(KEYINPUT62), .A2(G137), .ZN(n1352) );
NAND2_X1 U1081 ( .A1(G221), .A2(n1285), .ZN(n1351) );
AND2_X1 U1082 ( .A1(G234), .A2(n1070), .ZN(n1285) );
INV_X1 U1083 ( .A(G953), .ZN(n1070) );
XNOR2_X1 U1084 ( .A(n1353), .B(n1354), .ZN(n1347) );
NOR2_X1 U1085 ( .A1(KEYINPUT56), .A2(n1355), .ZN(n1354) );
XNOR2_X1 U1086 ( .A(G119), .B(n1356), .ZN(n1355) );
NAND2_X1 U1087 ( .A1(KEYINPUT18), .A2(n1292), .ZN(n1356) );
INV_X1 U1088 ( .A(G128), .ZN(n1292) );
NOR2_X1 U1089 ( .A1(KEYINPUT49), .A2(n1357), .ZN(n1353) );
XOR2_X1 U1090 ( .A(n1302), .B(KEYINPUT6), .Z(n1357) );
XOR2_X1 U1091 ( .A(n1344), .B(n1120), .Z(n1302) );
XOR2_X1 U1092 ( .A(G140), .B(G125), .Z(n1120) );
INV_X1 U1093 ( .A(G146), .ZN(n1344) );
INV_X1 U1094 ( .A(n1244), .ZN(n1267) );
XNOR2_X1 U1095 ( .A(G472), .B(n1358), .ZN(n1244) );
NOR2_X1 U1096 ( .A1(n1091), .A2(KEYINPUT30), .ZN(n1358) );
AND2_X1 U1097 ( .A1(n1359), .A2(n1280), .ZN(n1091) );
INV_X1 U1098 ( .A(G902), .ZN(n1280) );
XNOR2_X1 U1099 ( .A(n1170), .B(n1360), .ZN(n1359) );
XOR2_X1 U1100 ( .A(KEYINPUT43), .B(n1167), .Z(n1360) );
XNOR2_X1 U1101 ( .A(n1178), .B(n1310), .ZN(n1167) );
XOR2_X1 U1102 ( .A(n1139), .B(n1361), .Z(n1310) );
XOR2_X1 U1103 ( .A(G128), .B(n1362), .Z(n1361) );
NOR2_X1 U1104 ( .A1(KEYINPUT54), .A2(n1363), .ZN(n1362) );
XOR2_X1 U1105 ( .A(G146), .B(G143), .Z(n1363) );
XNOR2_X1 U1106 ( .A(n1275), .B(n1364), .ZN(n1139) );
XOR2_X1 U1107 ( .A(G119), .B(G116), .Z(n1364) );
INV_X1 U1108 ( .A(G113), .ZN(n1275) );
XOR2_X1 U1109 ( .A(n1365), .B(n1123), .Z(n1178) );
XOR2_X1 U1110 ( .A(G134), .B(G137), .Z(n1123) );
NAND2_X1 U1111 ( .A1(KEYINPUT9), .A2(G131), .ZN(n1365) );
AND2_X1 U1112 ( .A1(n1366), .A2(n1367), .ZN(n1170) );
NAND2_X1 U1113 ( .A1(n1368), .A2(n1247), .ZN(n1367) );
INV_X1 U1114 ( .A(G101), .ZN(n1247) );
NAND2_X1 U1115 ( .A1(G210), .A2(n1301), .ZN(n1368) );
NAND3_X1 U1116 ( .A1(G210), .A2(n1301), .A3(G101), .ZN(n1366) );
NOR2_X1 U1117 ( .A1(G953), .A2(G237), .ZN(n1301) );
endmodule


