//Key = 0111010000000111011000001101000100101100101000111110100001010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397;

XNOR2_X1 U755 ( .A(G107), .B(n1070), .ZN(G9) );
NOR2_X1 U756 ( .A1(n1071), .A2(n1072), .ZN(G75) );
NOR4_X1 U757 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1072) );
NOR2_X1 U758 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U759 ( .A(n1079), .B(KEYINPUT30), .Z(n1077) );
NAND4_X1 U760 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1079) );
XNOR2_X1 U761 ( .A(KEYINPUT22), .B(n1084), .ZN(n1083) );
NOR3_X1 U762 ( .A1(n1085), .A2(n1086), .A3(n1084), .ZN(n1075) );
NAND3_X1 U763 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1085) );
NAND2_X1 U764 ( .A1(n1090), .A2(n1091), .ZN(n1087) );
NAND2_X1 U765 ( .A1(n1092), .A2(n1082), .ZN(n1091) );
XNOR2_X1 U766 ( .A(n1093), .B(n1094), .ZN(n1092) );
NAND2_X1 U767 ( .A1(KEYINPUT48), .A2(n1095), .ZN(n1093) );
NAND2_X1 U768 ( .A1(n1081), .A2(n1096), .ZN(n1090) );
NAND2_X1 U769 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND3_X1 U770 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1073) );
NAND4_X1 U771 ( .A1(n1082), .A2(n1089), .A3(n1081), .A4(n1102), .ZN(n1101) );
NOR3_X1 U772 ( .A1(n1084), .A2(n1103), .A3(n1104), .ZN(n1102) );
NOR3_X1 U773 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1104) );
NOR2_X1 U774 ( .A1(n1080), .A2(n1088), .ZN(n1103) );
AND3_X1 U775 ( .A1(n1099), .A2(n1100), .A3(n1108), .ZN(n1071) );
NAND4_X1 U776 ( .A1(n1109), .A2(n1088), .A3(n1110), .A4(n1111), .ZN(n1099) );
NOR4_X1 U777 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1111) );
XNOR2_X1 U778 ( .A(n1116), .B(n1117), .ZN(n1112) );
NAND2_X1 U779 ( .A1(KEYINPUT15), .A2(n1118), .ZN(n1116) );
NOR3_X1 U780 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1110) );
NAND2_X1 U781 ( .A1(G475), .A2(n1122), .ZN(n1109) );
XOR2_X1 U782 ( .A(n1123), .B(n1124), .Z(G72) );
XOR2_X1 U783 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U784 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U785 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U786 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U787 ( .A(n1133), .B(n1134), .ZN(n1131) );
XOR2_X1 U788 ( .A(n1135), .B(KEYINPUT43), .Z(n1129) );
XNOR2_X1 U789 ( .A(KEYINPUT61), .B(KEYINPUT55), .ZN(n1135) );
NOR2_X1 U790 ( .A1(G900), .A2(n1100), .ZN(n1127) );
NAND2_X1 U791 ( .A1(n1100), .A2(n1136), .ZN(n1125) );
NAND2_X1 U792 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U793 ( .A1(G953), .A2(n1139), .ZN(n1123) );
NAND2_X1 U794 ( .A1(G900), .A2(G227), .ZN(n1139) );
NAND2_X1 U795 ( .A1(n1140), .A2(n1141), .ZN(G69) );
NAND2_X1 U796 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U797 ( .A1(n1144), .A2(n1145), .ZN(n1140) );
NAND2_X1 U798 ( .A1(n1146), .A2(n1143), .ZN(n1145) );
NAND2_X1 U799 ( .A1(G953), .A2(n1147), .ZN(n1143) );
INV_X1 U800 ( .A(G224), .ZN(n1147) );
INV_X1 U801 ( .A(n1148), .ZN(n1146) );
INV_X1 U802 ( .A(n1142), .ZN(n1144) );
XNOR2_X1 U803 ( .A(n1149), .B(n1150), .ZN(n1142) );
NOR2_X1 U804 ( .A1(n1148), .A2(n1151), .ZN(n1150) );
XNOR2_X1 U805 ( .A(n1152), .B(n1153), .ZN(n1151) );
NOR2_X1 U806 ( .A1(KEYINPUT60), .A2(n1154), .ZN(n1153) );
XOR2_X1 U807 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U808 ( .A1(KEYINPUT44), .A2(n1157), .ZN(n1156) );
NAND2_X1 U809 ( .A1(n1100), .A2(n1158), .ZN(n1149) );
NAND2_X1 U810 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U811 ( .A(n1161), .B(KEYINPUT11), .Z(n1159) );
NOR2_X1 U812 ( .A1(n1162), .A2(n1163), .ZN(G66) );
XOR2_X1 U813 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U814 ( .A1(n1166), .A2(n1167), .ZN(n1164) );
NOR2_X1 U815 ( .A1(n1162), .A2(n1168), .ZN(G63) );
XNOR2_X1 U816 ( .A(n1169), .B(n1170), .ZN(n1168) );
NOR2_X1 U817 ( .A1(n1171), .A2(n1167), .ZN(n1170) );
INV_X1 U818 ( .A(G478), .ZN(n1171) );
NOR2_X1 U819 ( .A1(n1162), .A2(n1172), .ZN(G60) );
XNOR2_X1 U820 ( .A(n1173), .B(n1174), .ZN(n1172) );
NOR2_X1 U821 ( .A1(n1175), .A2(n1167), .ZN(n1174) );
INV_X1 U822 ( .A(G475), .ZN(n1175) );
XNOR2_X1 U823 ( .A(G104), .B(n1176), .ZN(G6) );
NOR2_X1 U824 ( .A1(n1162), .A2(n1177), .ZN(G57) );
XOR2_X1 U825 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U826 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U827 ( .A1(n1182), .A2(n1167), .ZN(n1180) );
INV_X1 U828 ( .A(G472), .ZN(n1182) );
XNOR2_X1 U829 ( .A(n1183), .B(n1184), .ZN(n1178) );
NOR2_X1 U830 ( .A1(n1162), .A2(n1185), .ZN(G54) );
XOR2_X1 U831 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U832 ( .A(n1188), .B(n1189), .Z(n1187) );
NOR2_X1 U833 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U834 ( .A1(n1133), .A2(n1192), .ZN(n1191) );
XOR2_X1 U835 ( .A(n1193), .B(KEYINPUT10), .Z(n1192) );
INV_X1 U836 ( .A(n1184), .ZN(n1133) );
NOR2_X1 U837 ( .A1(n1184), .A2(n1194), .ZN(n1190) );
XOR2_X1 U838 ( .A(n1193), .B(KEYINPUT31), .Z(n1194) );
XOR2_X1 U839 ( .A(n1195), .B(n1196), .Z(n1193) );
XNOR2_X1 U840 ( .A(G140), .B(G110), .ZN(n1195) );
NOR2_X1 U841 ( .A1(n1197), .A2(n1167), .ZN(n1188) );
XNOR2_X1 U842 ( .A(G469), .B(KEYINPUT21), .ZN(n1197) );
XNOR2_X1 U843 ( .A(n1198), .B(KEYINPUT12), .ZN(n1186) );
NOR2_X1 U844 ( .A1(n1162), .A2(n1199), .ZN(G51) );
XOR2_X1 U845 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U846 ( .A(n1202), .B(n1203), .Z(n1201) );
NOR2_X1 U847 ( .A1(n1117), .A2(n1167), .ZN(n1203) );
NAND2_X1 U848 ( .A1(G902), .A2(n1074), .ZN(n1167) );
NAND4_X1 U849 ( .A1(n1137), .A2(n1160), .A3(n1204), .A4(n1161), .ZN(n1074) );
NAND2_X1 U850 ( .A1(n1205), .A2(n1206), .ZN(n1161) );
XNOR2_X1 U851 ( .A(n1107), .B(KEYINPUT47), .ZN(n1205) );
XNOR2_X1 U852 ( .A(KEYINPUT1), .B(n1138), .ZN(n1204) );
AND4_X1 U853 ( .A1(n1207), .A2(n1208), .A3(n1176), .A4(n1209), .ZN(n1160) );
NOR4_X1 U854 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1209) );
INV_X1 U855 ( .A(n1070), .ZN(n1213) );
NAND4_X1 U856 ( .A1(n1214), .A2(n1106), .A3(n1082), .A4(n1215), .ZN(n1070) );
NOR4_X1 U857 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1086), .ZN(n1211) );
NOR2_X1 U858 ( .A1(KEYINPUT63), .A2(n1219), .ZN(n1217) );
NOR3_X1 U859 ( .A1(n1078), .A2(n1081), .A3(n1220), .ZN(n1219) );
AND2_X1 U860 ( .A1(n1221), .A2(KEYINPUT63), .ZN(n1216) );
NAND4_X1 U861 ( .A1(n1107), .A2(n1214), .A3(n1082), .A4(n1215), .ZN(n1176) );
AND4_X1 U862 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1137) );
NOR4_X1 U863 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1225) );
INV_X1 U864 ( .A(n1230), .ZN(n1229) );
INV_X1 U865 ( .A(n1231), .ZN(n1228) );
NAND3_X1 U866 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1224) );
XNOR2_X1 U867 ( .A(n1080), .B(KEYINPUT27), .ZN(n1234) );
NAND2_X1 U868 ( .A1(n1235), .A2(n1236), .ZN(n1222) );
XNOR2_X1 U869 ( .A(KEYINPUT20), .B(n1078), .ZN(n1236) );
NOR2_X1 U870 ( .A1(n1237), .A2(n1238), .ZN(n1202) );
XOR2_X1 U871 ( .A(n1239), .B(KEYINPUT13), .Z(n1238) );
NAND2_X1 U872 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NOR2_X1 U873 ( .A1(n1241), .A2(n1240), .ZN(n1237) );
XNOR2_X1 U874 ( .A(G125), .B(n1183), .ZN(n1240) );
AND2_X1 U875 ( .A1(n1242), .A2(n1108), .ZN(n1162) );
XNOR2_X1 U876 ( .A(G953), .B(KEYINPUT25), .ZN(n1242) );
XNOR2_X1 U877 ( .A(G146), .B(n1223), .ZN(G48) );
NAND2_X1 U878 ( .A1(n1243), .A2(n1107), .ZN(n1223) );
XNOR2_X1 U879 ( .A(G143), .B(n1231), .ZN(G45) );
NAND4_X1 U880 ( .A1(n1244), .A2(n1245), .A3(n1214), .A4(n1246), .ZN(n1231) );
XNOR2_X1 U881 ( .A(n1247), .B(n1227), .ZN(G42) );
AND3_X1 U882 ( .A1(n1107), .A2(n1233), .A3(n1248), .ZN(n1227) );
NAND2_X1 U883 ( .A1(n1249), .A2(n1250), .ZN(G39) );
NAND2_X1 U884 ( .A1(G137), .A2(n1251), .ZN(n1250) );
XOR2_X1 U885 ( .A(n1252), .B(KEYINPUT53), .Z(n1249) );
OR2_X1 U886 ( .A1(n1251), .A2(G137), .ZN(n1252) );
NAND3_X1 U887 ( .A1(n1232), .A2(n1233), .A3(n1080), .ZN(n1251) );
XOR2_X1 U888 ( .A(G134), .B(n1226), .Z(G36) );
AND3_X1 U889 ( .A1(n1233), .A2(n1106), .A3(n1245), .ZN(n1226) );
NAND2_X1 U890 ( .A1(n1253), .A2(n1254), .ZN(G33) );
NAND2_X1 U891 ( .A1(G131), .A2(n1230), .ZN(n1254) );
XOR2_X1 U892 ( .A(KEYINPUT57), .B(n1255), .Z(n1253) );
NOR2_X1 U893 ( .A1(G131), .A2(n1230), .ZN(n1255) );
NAND3_X1 U894 ( .A1(n1245), .A2(n1233), .A3(n1107), .ZN(n1230) );
AND3_X1 U895 ( .A1(n1089), .A2(n1256), .A3(n1257), .ZN(n1233) );
NOR3_X1 U896 ( .A1(n1258), .A2(n1259), .A3(n1105), .ZN(n1257) );
XNOR2_X1 U897 ( .A(n1260), .B(KEYINPUT18), .ZN(n1089) );
XNOR2_X1 U898 ( .A(G128), .B(n1138), .ZN(G30) );
NAND2_X1 U899 ( .A1(n1243), .A2(n1106), .ZN(n1138) );
AND3_X1 U900 ( .A1(n1214), .A2(n1246), .A3(n1232), .ZN(n1243) );
INV_X1 U901 ( .A(n1218), .ZN(n1232) );
XNOR2_X1 U902 ( .A(G101), .B(n1207), .ZN(G3) );
NAND4_X1 U903 ( .A1(n1080), .A2(n1245), .A3(n1214), .A4(n1215), .ZN(n1207) );
XOR2_X1 U904 ( .A(G125), .B(n1261), .Z(G27) );
AND2_X1 U905 ( .A1(n1262), .A2(n1235), .ZN(n1261) );
NOR4_X1 U906 ( .A1(n1097), .A2(n1263), .A3(n1114), .A4(n1258), .ZN(n1235) );
INV_X1 U907 ( .A(n1246), .ZN(n1258) );
NAND2_X1 U908 ( .A1(n1084), .A2(n1264), .ZN(n1246) );
NAND4_X1 U909 ( .A1(n1265), .A2(G953), .A3(n1266), .A4(n1267), .ZN(n1264) );
INV_X1 U910 ( .A(G900), .ZN(n1267) );
XNOR2_X1 U911 ( .A(G902), .B(KEYINPUT37), .ZN(n1265) );
NAND2_X1 U912 ( .A1(n1268), .A2(n1269), .ZN(G24) );
NAND2_X1 U913 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XOR2_X1 U914 ( .A(n1272), .B(KEYINPUT6), .Z(n1268) );
OR2_X1 U915 ( .A1(n1270), .A2(n1271), .ZN(n1272) );
NAND2_X1 U916 ( .A1(n1273), .A2(n1274), .ZN(n1270) );
NAND2_X1 U917 ( .A1(n1210), .A2(n1275), .ZN(n1274) );
INV_X1 U918 ( .A(KEYINPUT28), .ZN(n1275) );
AND3_X1 U919 ( .A1(n1244), .A2(n1082), .A3(n1276), .ZN(n1210) );
INV_X1 U920 ( .A(n1277), .ZN(n1244) );
NAND4_X1 U921 ( .A1(n1082), .A2(n1277), .A3(n1276), .A4(KEYINPUT28), .ZN(n1273) );
NAND2_X1 U922 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NOR2_X1 U923 ( .A1(n1280), .A2(n1281), .ZN(n1082) );
XOR2_X1 U924 ( .A(G119), .B(n1282), .Z(G21) );
NOR3_X1 U925 ( .A1(n1221), .A2(n1218), .A3(n1086), .ZN(n1282) );
INV_X1 U926 ( .A(n1080), .ZN(n1086) );
NAND2_X1 U927 ( .A1(n1281), .A2(n1280), .ZN(n1218) );
INV_X1 U928 ( .A(n1283), .ZN(n1280) );
XNOR2_X1 U929 ( .A(G116), .B(n1208), .ZN(G18) );
NAND2_X1 U930 ( .A1(n1206), .A2(n1106), .ZN(n1208) );
NOR2_X1 U931 ( .A1(n1284), .A2(n1285), .ZN(n1106) );
XNOR2_X1 U932 ( .A(G113), .B(n1286), .ZN(G15) );
NAND2_X1 U933 ( .A1(n1206), .A2(n1107), .ZN(n1286) );
INV_X1 U934 ( .A(n1263), .ZN(n1107) );
NAND2_X1 U935 ( .A1(n1287), .A2(n1285), .ZN(n1263) );
XOR2_X1 U936 ( .A(n1278), .B(KEYINPUT51), .Z(n1287) );
XOR2_X1 U937 ( .A(n1284), .B(KEYINPUT45), .Z(n1278) );
NOR2_X1 U938 ( .A1(n1221), .A2(n1098), .ZN(n1206) );
INV_X1 U939 ( .A(n1245), .ZN(n1098) );
NOR2_X1 U940 ( .A1(n1283), .A2(n1281), .ZN(n1245) );
INV_X1 U941 ( .A(n1276), .ZN(n1221) );
NOR3_X1 U942 ( .A1(n1078), .A2(n1220), .A3(n1114), .ZN(n1276) );
INV_X1 U943 ( .A(n1081), .ZN(n1114) );
NOR2_X1 U944 ( .A1(n1256), .A2(n1259), .ZN(n1081) );
NAND2_X1 U945 ( .A1(n1288), .A2(n1289), .ZN(G12) );
NAND2_X1 U946 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
XOR2_X1 U947 ( .A(n1292), .B(KEYINPUT0), .Z(n1288) );
OR2_X1 U948 ( .A1(n1290), .A2(n1291), .ZN(n1292) );
NAND2_X1 U949 ( .A1(n1293), .A2(n1294), .ZN(n1290) );
NAND2_X1 U950 ( .A1(n1212), .A2(n1295), .ZN(n1294) );
INV_X1 U951 ( .A(KEYINPUT41), .ZN(n1295) );
AND2_X1 U952 ( .A1(n1296), .A2(n1215), .ZN(n1212) );
NAND3_X1 U953 ( .A1(n1220), .A2(n1296), .A3(KEYINPUT41), .ZN(n1293) );
AND3_X1 U954 ( .A1(n1248), .A2(n1214), .A3(n1080), .ZN(n1296) );
NOR2_X1 U955 ( .A1(n1279), .A2(n1284), .ZN(n1080) );
NAND3_X1 U956 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1284) );
INV_X1 U957 ( .A(n1119), .ZN(n1299) );
NOR2_X1 U958 ( .A1(n1122), .A2(G475), .ZN(n1119) );
OR2_X1 U959 ( .A1(G475), .A2(KEYINPUT36), .ZN(n1298) );
NAND3_X1 U960 ( .A1(G475), .A2(n1122), .A3(KEYINPUT36), .ZN(n1297) );
NAND2_X1 U961 ( .A1(n1173), .A2(n1300), .ZN(n1122) );
XNOR2_X1 U962 ( .A(n1301), .B(n1302), .ZN(n1173) );
XNOR2_X1 U963 ( .A(n1303), .B(n1304), .ZN(n1302) );
XNOR2_X1 U964 ( .A(n1134), .B(n1305), .ZN(n1304) );
XOR2_X1 U965 ( .A(n1306), .B(n1307), .Z(n1301) );
XOR2_X1 U966 ( .A(n1308), .B(n1309), .Z(n1307) );
NAND2_X1 U967 ( .A1(KEYINPUT52), .A2(n1310), .ZN(n1309) );
INV_X1 U968 ( .A(G131), .ZN(n1310) );
NAND2_X1 U969 ( .A1(n1311), .A2(G214), .ZN(n1308) );
XNOR2_X1 U970 ( .A(G113), .B(n1312), .ZN(n1306) );
NOR2_X1 U971 ( .A1(KEYINPUT58), .A2(G122), .ZN(n1312) );
INV_X1 U972 ( .A(n1285), .ZN(n1279) );
NOR2_X1 U973 ( .A1(n1313), .A2(n1121), .ZN(n1285) );
NOR3_X1 U974 ( .A1(G478), .A2(G902), .A3(n1314), .ZN(n1121) );
INV_X1 U975 ( .A(n1169), .ZN(n1314) );
XNOR2_X1 U976 ( .A(KEYINPUT59), .B(n1120), .ZN(n1313) );
AND2_X1 U977 ( .A1(G478), .A2(n1315), .ZN(n1120) );
NAND2_X1 U978 ( .A1(n1169), .A2(n1300), .ZN(n1315) );
XNOR2_X1 U979 ( .A(n1316), .B(n1317), .ZN(n1169) );
XOR2_X1 U980 ( .A(n1318), .B(n1319), .Z(n1317) );
XNOR2_X1 U981 ( .A(n1271), .B(G116), .ZN(n1319) );
INV_X1 U982 ( .A(G122), .ZN(n1271) );
XNOR2_X1 U983 ( .A(n1320), .B(G134), .ZN(n1318) );
XOR2_X1 U984 ( .A(n1321), .B(n1322), .Z(n1316) );
XNOR2_X1 U985 ( .A(n1323), .B(n1324), .ZN(n1321) );
INV_X1 U986 ( .A(G107), .ZN(n1324) );
NAND2_X1 U987 ( .A1(G217), .A2(n1325), .ZN(n1323) );
NOR3_X1 U988 ( .A1(n1095), .A2(n1259), .A3(n1078), .ZN(n1214) );
INV_X1 U989 ( .A(n1262), .ZN(n1078) );
NOR2_X1 U990 ( .A1(n1260), .A2(n1105), .ZN(n1262) );
INV_X1 U991 ( .A(n1088), .ZN(n1105) );
NAND2_X1 U992 ( .A1(G214), .A2(n1326), .ZN(n1088) );
XNOR2_X1 U993 ( .A(n1327), .B(n1117), .ZN(n1260) );
NAND2_X1 U994 ( .A1(G210), .A2(n1326), .ZN(n1117) );
NAND2_X1 U995 ( .A1(n1328), .A2(n1300), .ZN(n1326) );
XOR2_X1 U996 ( .A(n1118), .B(KEYINPUT8), .Z(n1327) );
NAND2_X1 U997 ( .A1(n1329), .A2(n1300), .ZN(n1118) );
XOR2_X1 U998 ( .A(n1330), .B(n1331), .Z(n1329) );
XNOR2_X1 U999 ( .A(n1332), .B(n1333), .ZN(n1331) );
NAND2_X1 U1000 ( .A1(KEYINPUT42), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1001 ( .A(KEYINPUT17), .B(n1200), .Z(n1334) );
XNOR2_X1 U1002 ( .A(n1335), .B(n1152), .ZN(n1200) );
XNOR2_X1 U1003 ( .A(G122), .B(n1291), .ZN(n1152) );
XNOR2_X1 U1004 ( .A(n1336), .B(n1157), .ZN(n1335) );
XNOR2_X1 U1005 ( .A(n1337), .B(n1303), .ZN(n1157) );
NAND2_X1 U1006 ( .A1(KEYINPUT50), .A2(n1155), .ZN(n1336) );
XOR2_X1 U1007 ( .A(n1338), .B(n1339), .Z(n1155) );
XNOR2_X1 U1008 ( .A(KEYINPUT14), .B(n1340), .ZN(n1339) );
XNOR2_X1 U1009 ( .A(G113), .B(n1341), .ZN(n1338) );
NAND2_X1 U1010 ( .A1(KEYINPUT24), .A2(n1342), .ZN(n1332) );
INV_X1 U1011 ( .A(n1183), .ZN(n1342) );
XNOR2_X1 U1012 ( .A(G125), .B(n1241), .ZN(n1330) );
AND2_X1 U1013 ( .A1(G224), .A2(n1343), .ZN(n1241) );
INV_X1 U1014 ( .A(n1094), .ZN(n1259) );
NAND2_X1 U1015 ( .A1(G221), .A2(n1344), .ZN(n1094) );
INV_X1 U1016 ( .A(n1256), .ZN(n1095) );
XNOR2_X1 U1017 ( .A(n1345), .B(G469), .ZN(n1256) );
NAND2_X1 U1018 ( .A1(n1300), .A2(n1346), .ZN(n1345) );
NAND2_X1 U1019 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
NAND3_X1 U1020 ( .A1(n1349), .A2(n1350), .A3(n1351), .ZN(n1348) );
XOR2_X1 U1021 ( .A(n1352), .B(KEYINPUT7), .Z(n1347) );
NAND2_X1 U1022 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
NAND2_X1 U1023 ( .A1(n1349), .A2(n1350), .ZN(n1354) );
NAND2_X1 U1024 ( .A1(n1355), .A2(n1356), .ZN(n1350) );
XNOR2_X1 U1025 ( .A(G140), .B(n1357), .ZN(n1356) );
XNOR2_X1 U1026 ( .A(n1198), .B(KEYINPUT4), .ZN(n1355) );
NAND2_X1 U1027 ( .A1(n1198), .A2(n1358), .ZN(n1349) );
XNOR2_X1 U1028 ( .A(n1247), .B(n1357), .ZN(n1358) );
NOR2_X1 U1029 ( .A1(G110), .A2(KEYINPUT23), .ZN(n1357) );
AND2_X1 U1030 ( .A1(G227), .A2(n1343), .ZN(n1198) );
INV_X1 U1031 ( .A(n1351), .ZN(n1353) );
XOR2_X1 U1032 ( .A(n1184), .B(n1196), .Z(n1351) );
XOR2_X1 U1033 ( .A(n1132), .B(n1359), .Z(n1196) );
XOR2_X1 U1034 ( .A(n1360), .B(n1337), .Z(n1359) );
XNOR2_X1 U1035 ( .A(G101), .B(G107), .ZN(n1337) );
NAND2_X1 U1036 ( .A1(KEYINPUT2), .A2(n1303), .ZN(n1360) );
XNOR2_X1 U1037 ( .A(G104), .B(KEYINPUT39), .ZN(n1303) );
XOR2_X1 U1038 ( .A(n1322), .B(n1361), .Z(n1132) );
NOR2_X1 U1039 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
XOR2_X1 U1040 ( .A(KEYINPUT26), .B(n1364), .Z(n1363) );
NOR2_X1 U1041 ( .A1(G146), .A2(n1365), .ZN(n1364) );
XNOR2_X1 U1042 ( .A(KEYINPUT40), .B(n1320), .ZN(n1365) );
INV_X1 U1043 ( .A(G143), .ZN(n1320) );
NOR2_X1 U1044 ( .A1(G143), .A2(n1366), .ZN(n1362) );
XOR2_X1 U1045 ( .A(KEYINPUT34), .B(G146), .Z(n1366) );
INV_X1 U1046 ( .A(n1097), .ZN(n1248) );
NAND2_X1 U1047 ( .A1(n1281), .A2(n1283), .ZN(n1097) );
XNOR2_X1 U1048 ( .A(n1367), .B(n1115), .ZN(n1283) );
XNOR2_X1 U1049 ( .A(n1368), .B(G472), .ZN(n1115) );
NAND2_X1 U1050 ( .A1(n1369), .A2(n1300), .ZN(n1368) );
XNOR2_X1 U1051 ( .A(n1370), .B(n1181), .ZN(n1369) );
XNOR2_X1 U1052 ( .A(n1371), .B(n1372), .ZN(n1181) );
XOR2_X1 U1053 ( .A(n1373), .B(n1374), .Z(n1372) );
NAND2_X1 U1054 ( .A1(n1311), .A2(G210), .ZN(n1374) );
AND2_X1 U1055 ( .A1(n1343), .A2(n1328), .ZN(n1311) );
INV_X1 U1056 ( .A(G237), .ZN(n1328) );
NAND2_X1 U1057 ( .A1(n1375), .A2(n1376), .ZN(n1373) );
OR2_X1 U1058 ( .A1(n1341), .A2(n1340), .ZN(n1376) );
XOR2_X1 U1059 ( .A(n1377), .B(KEYINPUT32), .Z(n1375) );
NAND2_X1 U1060 ( .A1(n1341), .A2(n1340), .ZN(n1377) );
INV_X1 U1061 ( .A(G116), .ZN(n1340) );
XNOR2_X1 U1062 ( .A(G101), .B(n1378), .ZN(n1371) );
XNOR2_X1 U1063 ( .A(KEYINPUT46), .B(n1379), .ZN(n1378) );
INV_X1 U1064 ( .A(G113), .ZN(n1379) );
NAND2_X1 U1065 ( .A1(n1380), .A2(n1381), .ZN(n1370) );
NAND2_X1 U1066 ( .A1(n1382), .A2(n1183), .ZN(n1381) );
XOR2_X1 U1067 ( .A(KEYINPUT49), .B(n1383), .Z(n1380) );
NOR2_X1 U1068 ( .A1(n1382), .A2(n1183), .ZN(n1383) );
XOR2_X1 U1069 ( .A(n1305), .B(n1384), .Z(n1183) );
XOR2_X1 U1070 ( .A(KEYINPUT16), .B(n1322), .Z(n1384) );
XOR2_X1 U1071 ( .A(G143), .B(G146), .Z(n1305) );
XNOR2_X1 U1072 ( .A(n1184), .B(KEYINPUT62), .ZN(n1382) );
XOR2_X1 U1073 ( .A(G131), .B(n1385), .Z(n1184) );
XOR2_X1 U1074 ( .A(G137), .B(G134), .Z(n1385) );
XNOR2_X1 U1075 ( .A(KEYINPUT5), .B(KEYINPUT35), .ZN(n1367) );
XNOR2_X1 U1076 ( .A(n1113), .B(KEYINPUT3), .ZN(n1281) );
XOR2_X1 U1077 ( .A(n1386), .B(n1166), .Z(n1113) );
NAND2_X1 U1078 ( .A1(G217), .A2(n1344), .ZN(n1166) );
NAND2_X1 U1079 ( .A1(G234), .A2(n1300), .ZN(n1344) );
INV_X1 U1080 ( .A(G902), .ZN(n1300) );
OR2_X1 U1081 ( .A1(n1165), .A2(G902), .ZN(n1386) );
XNOR2_X1 U1082 ( .A(n1387), .B(n1388), .ZN(n1165) );
XOR2_X1 U1083 ( .A(n1389), .B(n1390), .Z(n1388) );
XNOR2_X1 U1084 ( .A(G137), .B(n1291), .ZN(n1390) );
INV_X1 U1085 ( .A(G110), .ZN(n1291) );
XOR2_X1 U1086 ( .A(KEYINPUT56), .B(G146), .Z(n1389) );
XOR2_X1 U1087 ( .A(n1391), .B(n1392), .Z(n1387) );
XOR2_X1 U1088 ( .A(n1393), .B(n1394), .Z(n1392) );
NOR2_X1 U1089 ( .A1(KEYINPUT38), .A2(n1134), .ZN(n1394) );
XOR2_X1 U1090 ( .A(G125), .B(n1247), .Z(n1134) );
INV_X1 U1091 ( .A(G140), .ZN(n1247) );
NOR2_X1 U1092 ( .A1(KEYINPUT19), .A2(n1341), .ZN(n1393) );
XOR2_X1 U1093 ( .A(G119), .B(KEYINPUT33), .Z(n1341) );
XOR2_X1 U1094 ( .A(n1395), .B(n1322), .Z(n1391) );
XOR2_X1 U1095 ( .A(G128), .B(KEYINPUT54), .Z(n1322) );
NAND2_X1 U1096 ( .A1(n1325), .A2(G221), .ZN(n1395) );
AND2_X1 U1097 ( .A1(G234), .A2(n1343), .ZN(n1325) );
XNOR2_X1 U1098 ( .A(G953), .B(KEYINPUT29), .ZN(n1343) );
INV_X1 U1099 ( .A(n1215), .ZN(n1220) );
NAND2_X1 U1100 ( .A1(n1084), .A2(n1396), .ZN(n1215) );
NAND3_X1 U1101 ( .A1(n1148), .A2(n1266), .A3(G902), .ZN(n1396) );
NOR2_X1 U1102 ( .A1(G898), .A2(n1100), .ZN(n1148) );
NAND3_X1 U1103 ( .A1(n1266), .A2(n1100), .A3(n1397), .ZN(n1084) );
XNOR2_X1 U1104 ( .A(KEYINPUT9), .B(n1108), .ZN(n1397) );
INV_X1 U1105 ( .A(G952), .ZN(n1108) );
INV_X1 U1106 ( .A(G953), .ZN(n1100) );
NAND2_X1 U1107 ( .A1(G237), .A2(G234), .ZN(n1266) );
endmodule


