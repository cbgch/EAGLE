//Key = 0111111001110001010000100110000110110000100011000101011101010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351;

XNOR2_X1 U743 ( .A(G107), .B(n1029), .ZN(G9) );
NOR2_X1 U744 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U745 ( .A1(G953), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1031) );
XOR2_X1 U746 ( .A(n1035), .B(KEYINPUT43), .Z(n1033) );
NAND2_X1 U747 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U748 ( .A1(n1038), .A2(n1039), .A3(KEYINPUT12), .ZN(n1037) );
NAND4_X1 U749 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NAND2_X1 U750 ( .A1(n1041), .A2(n1044), .ZN(n1036) );
NAND2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND3_X1 U752 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND2_X1 U753 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND2_X1 U754 ( .A1(n1038), .A2(n1052), .ZN(n1051) );
NAND2_X1 U755 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U756 ( .A1(n1043), .A2(n1055), .ZN(n1050) );
NAND2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U758 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND3_X1 U759 ( .A1(n1043), .A2(n1060), .A3(n1038), .ZN(n1045) );
NAND3_X1 U760 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NAND2_X1 U761 ( .A1(n1047), .A2(n1064), .ZN(n1063) );
NAND2_X1 U762 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
INV_X1 U764 ( .A(n1069), .ZN(n1065) );
NAND3_X1 U765 ( .A1(n1042), .A2(n1070), .A3(n1040), .ZN(n1062) );
XNOR2_X1 U766 ( .A(n1049), .B(KEYINPUT59), .ZN(n1040) );
INV_X1 U767 ( .A(KEYINPUT12), .ZN(n1070) );
NAND3_X1 U768 ( .A1(n1071), .A2(n1049), .A3(n1072), .ZN(n1061) );
INV_X1 U769 ( .A(n1073), .ZN(n1041) );
NOR3_X1 U770 ( .A1(n1032), .A2(G953), .A3(G952), .ZN(n1030) );
AND4_X1 U771 ( .A1(n1074), .A2(n1049), .A3(n1075), .A4(n1076), .ZN(n1032) );
NOR4_X1 U772 ( .A1(n1058), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1076) );
XNOR2_X1 U773 ( .A(n1080), .B(n1081), .ZN(n1075) );
XNOR2_X1 U774 ( .A(n1082), .B(n1083), .ZN(n1074) );
XOR2_X1 U775 ( .A(n1084), .B(n1085), .Z(G72) );
NOR2_X1 U776 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
AND2_X1 U777 ( .A1(G227), .A2(G900), .ZN(n1086) );
NOR2_X1 U778 ( .A1(KEYINPUT46), .A2(n1088), .ZN(n1084) );
XOR2_X1 U779 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U780 ( .A1(n1091), .A2(G953), .ZN(n1090) );
NOR2_X1 U781 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U782 ( .A1(n1094), .A2(n1095), .ZN(n1089) );
NAND2_X1 U783 ( .A1(G953), .A2(n1096), .ZN(n1095) );
XNOR2_X1 U784 ( .A(n1097), .B(n1098), .ZN(n1094) );
XOR2_X1 U785 ( .A(n1099), .B(n1100), .Z(n1098) );
NAND3_X1 U786 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1099) );
OR2_X1 U787 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND3_X1 U788 ( .A1(n1105), .A2(n1104), .A3(n1106), .ZN(n1102) );
INV_X1 U789 ( .A(G131), .ZN(n1106) );
NAND2_X1 U790 ( .A1(G131), .A2(n1107), .ZN(n1101) );
NAND2_X1 U791 ( .A1(n1108), .A2(n1104), .ZN(n1107) );
INV_X1 U792 ( .A(KEYINPUT24), .ZN(n1104) );
XNOR2_X1 U793 ( .A(n1105), .B(KEYINPUT54), .ZN(n1108) );
XNOR2_X1 U794 ( .A(n1109), .B(G134), .ZN(n1105) );
NAND2_X1 U795 ( .A1(KEYINPUT49), .A2(n1110), .ZN(n1109) );
XOR2_X1 U796 ( .A(n1111), .B(n1112), .Z(G69) );
XOR2_X1 U797 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1087), .ZN(n1114) );
NOR2_X1 U799 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(n1113) );
NAND2_X1 U801 ( .A1(G953), .A2(n1117), .ZN(n1119) );
XOR2_X1 U802 ( .A(n1120), .B(n1121), .Z(n1118) );
XNOR2_X1 U803 ( .A(n1122), .B(n1123), .ZN(n1121) );
NAND2_X1 U804 ( .A1(n1087), .A2(n1124), .ZN(n1111) );
NAND3_X1 U805 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1124) );
XOR2_X1 U806 ( .A(n1128), .B(KEYINPUT16), .Z(n1127) );
XOR2_X1 U807 ( .A(n1129), .B(KEYINPUT7), .Z(n1125) );
NOR2_X1 U808 ( .A1(n1130), .A2(n1131), .ZN(G66) );
NOR3_X1 U809 ( .A1(n1080), .A2(n1132), .A3(n1133), .ZN(n1131) );
NOR3_X1 U810 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1133) );
NOR2_X1 U811 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
AND2_X1 U812 ( .A1(n1034), .A2(n1081), .ZN(n1137) );
NOR2_X1 U813 ( .A1(n1130), .A2(n1139), .ZN(G63) );
XNOR2_X1 U814 ( .A(n1140), .B(n1141), .ZN(n1139) );
NOR2_X1 U815 ( .A1(n1142), .A2(n1136), .ZN(n1141) );
NOR2_X1 U816 ( .A1(n1130), .A2(n1143), .ZN(G60) );
XOR2_X1 U817 ( .A(n1144), .B(n1145), .Z(n1143) );
NOR2_X1 U818 ( .A1(n1146), .A2(n1136), .ZN(n1144) );
XOR2_X1 U819 ( .A(n1147), .B(n1148), .Z(G6) );
XOR2_X1 U820 ( .A(KEYINPUT4), .B(G104), .Z(n1148) );
NAND3_X1 U821 ( .A1(n1149), .A2(n1150), .A3(KEYINPUT9), .ZN(n1147) );
NOR2_X1 U822 ( .A1(n1130), .A2(n1151), .ZN(G57) );
XOR2_X1 U823 ( .A(n1152), .B(n1153), .Z(n1151) );
XNOR2_X1 U824 ( .A(n1154), .B(n1155), .ZN(n1153) );
XOR2_X1 U825 ( .A(n1156), .B(n1157), .Z(n1152) );
XOR2_X1 U826 ( .A(KEYINPUT25), .B(n1158), .Z(n1157) );
NOR2_X1 U827 ( .A1(n1159), .A2(n1136), .ZN(n1158) );
NOR2_X1 U828 ( .A1(KEYINPUT38), .A2(n1160), .ZN(n1156) );
NOR2_X1 U829 ( .A1(n1130), .A2(n1161), .ZN(G54) );
XOR2_X1 U830 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U831 ( .A1(n1164), .A2(n1136), .ZN(n1163) );
NOR2_X1 U832 ( .A1(KEYINPUT48), .A2(n1165), .ZN(n1162) );
XOR2_X1 U833 ( .A(n1166), .B(n1167), .Z(n1165) );
XNOR2_X1 U834 ( .A(n1168), .B(KEYINPUT39), .ZN(n1167) );
NOR2_X1 U835 ( .A1(n1130), .A2(n1169), .ZN(G51) );
XOR2_X1 U836 ( .A(n1170), .B(n1171), .Z(n1169) );
XNOR2_X1 U837 ( .A(n1172), .B(n1173), .ZN(n1171) );
NOR2_X1 U838 ( .A1(KEYINPUT27), .A2(n1174), .ZN(n1173) );
XOR2_X1 U839 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U840 ( .A(G125), .B(n1177), .ZN(n1175) );
NOR2_X1 U841 ( .A1(n1178), .A2(n1136), .ZN(n1170) );
NAND2_X1 U842 ( .A1(G902), .A2(n1034), .ZN(n1136) );
NAND4_X1 U843 ( .A1(n1128), .A2(n1129), .A3(n1126), .A4(n1179), .ZN(n1034) );
NOR2_X1 U844 ( .A1(n1093), .A2(n1180), .ZN(n1179) );
XOR2_X1 U845 ( .A(KEYINPUT14), .B(n1092), .Z(n1180) );
NAND4_X1 U846 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1093) );
AND4_X1 U847 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1184) );
AND4_X1 U848 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1126) );
AND3_X1 U849 ( .A1(n1193), .A2(n1029), .A3(n1194), .ZN(n1192) );
NAND3_X1 U850 ( .A1(n1195), .A2(n1196), .A3(n1047), .ZN(n1029) );
NAND2_X1 U851 ( .A1(n1150), .A2(n1197), .ZN(n1191) );
XOR2_X1 U852 ( .A(KEYINPUT36), .B(n1149), .Z(n1197) );
AND4_X1 U853 ( .A1(n1198), .A2(n1047), .A3(n1069), .A4(n1199), .ZN(n1149) );
NAND4_X1 U854 ( .A1(n1042), .A2(n1198), .A3(n1200), .A4(n1201), .ZN(n1189) );
OR2_X1 U855 ( .A1(n1202), .A2(KEYINPUT63), .ZN(n1201) );
NAND2_X1 U856 ( .A1(KEYINPUT63), .A2(n1203), .ZN(n1200) );
NAND3_X1 U857 ( .A1(n1199), .A2(n1056), .A3(n1049), .ZN(n1203) );
INV_X1 U858 ( .A(n1150), .ZN(n1056) );
NOR2_X1 U859 ( .A1(n1087), .A2(G952), .ZN(n1130) );
XOR2_X1 U860 ( .A(G146), .B(n1204), .Z(G48) );
NOR2_X1 U861 ( .A1(KEYINPUT56), .A2(n1183), .ZN(n1204) );
NAND3_X1 U862 ( .A1(n1198), .A2(n1150), .A3(n1205), .ZN(n1183) );
XNOR2_X1 U863 ( .A(G143), .B(n1181), .ZN(G45) );
NAND4_X1 U864 ( .A1(n1206), .A2(n1150), .A3(n1079), .A4(n1078), .ZN(n1181) );
XOR2_X1 U865 ( .A(G140), .B(n1092), .Z(G42) );
AND3_X1 U866 ( .A1(n1207), .A2(n1069), .A3(n1038), .ZN(n1092) );
XNOR2_X1 U867 ( .A(G137), .B(n1182), .ZN(G39) );
NAND3_X1 U868 ( .A1(n1205), .A2(n1043), .A3(n1038), .ZN(n1182) );
XNOR2_X1 U869 ( .A(G134), .B(n1188), .ZN(G36) );
NAND3_X1 U870 ( .A1(n1206), .A2(n1195), .A3(n1038), .ZN(n1188) );
NAND2_X1 U871 ( .A1(n1208), .A2(n1209), .ZN(G33) );
NAND2_X1 U872 ( .A1(G131), .A2(n1187), .ZN(n1209) );
XOR2_X1 U873 ( .A(n1210), .B(KEYINPUT19), .Z(n1208) );
OR2_X1 U874 ( .A1(n1187), .A2(G131), .ZN(n1210) );
NAND3_X1 U875 ( .A1(n1206), .A2(n1198), .A3(n1038), .ZN(n1187) );
AND2_X1 U876 ( .A1(n1211), .A2(n1059), .ZN(n1038) );
AND3_X1 U877 ( .A1(n1069), .A2(n1212), .A3(n1042), .ZN(n1206) );
XNOR2_X1 U878 ( .A(G128), .B(n1186), .ZN(G30) );
NAND3_X1 U879 ( .A1(n1195), .A2(n1150), .A3(n1205), .ZN(n1186) );
AND4_X1 U880 ( .A1(n1072), .A2(n1069), .A3(n1213), .A4(n1212), .ZN(n1205) );
XNOR2_X1 U881 ( .A(G101), .B(n1128), .ZN(G3) );
NAND3_X1 U882 ( .A1(n1196), .A2(n1043), .A3(n1042), .ZN(n1128) );
XNOR2_X1 U883 ( .A(G125), .B(n1185), .ZN(G27) );
NAND3_X1 U884 ( .A1(n1049), .A2(n1150), .A3(n1207), .ZN(n1185) );
AND4_X1 U885 ( .A1(n1072), .A2(n1198), .A3(n1071), .A4(n1212), .ZN(n1207) );
NAND2_X1 U886 ( .A1(n1073), .A2(n1214), .ZN(n1212) );
NAND4_X1 U887 ( .A1(G953), .A2(G902), .A3(n1215), .A4(n1096), .ZN(n1214) );
INV_X1 U888 ( .A(G900), .ZN(n1096) );
XNOR2_X1 U889 ( .A(G122), .B(n1129), .ZN(G24) );
NAND4_X1 U890 ( .A1(n1202), .A2(n1047), .A3(n1079), .A4(n1078), .ZN(n1129) );
NOR2_X1 U891 ( .A1(n1213), .A2(n1072), .ZN(n1047) );
XNOR2_X1 U892 ( .A(n1190), .B(n1216), .ZN(G21) );
NOR2_X1 U893 ( .A1(KEYINPUT52), .A2(n1217), .ZN(n1216) );
NAND4_X1 U894 ( .A1(n1202), .A2(n1072), .A3(n1043), .A4(n1213), .ZN(n1190) );
XNOR2_X1 U895 ( .A(G116), .B(n1193), .ZN(G18) );
NAND3_X1 U896 ( .A1(n1042), .A2(n1195), .A3(n1202), .ZN(n1193) );
INV_X1 U897 ( .A(n1054), .ZN(n1195) );
NAND2_X1 U898 ( .A1(n1218), .A2(n1078), .ZN(n1054) );
XNOR2_X1 U899 ( .A(KEYINPUT2), .B(n1219), .ZN(n1218) );
XOR2_X1 U900 ( .A(n1220), .B(n1221), .Z(G15) );
AND3_X1 U901 ( .A1(n1202), .A2(n1198), .A3(n1042), .ZN(n1221) );
NOR2_X1 U902 ( .A1(n1071), .A2(n1072), .ZN(n1042) );
AND3_X1 U903 ( .A1(n1150), .A2(n1199), .A3(n1049), .ZN(n1202) );
NOR2_X1 U904 ( .A1(n1222), .A2(n1067), .ZN(n1049) );
XNOR2_X1 U905 ( .A(G113), .B(KEYINPUT6), .ZN(n1220) );
XNOR2_X1 U906 ( .A(G110), .B(n1194), .ZN(G12) );
NAND4_X1 U907 ( .A1(n1072), .A2(n1196), .A3(n1071), .A4(n1043), .ZN(n1194) );
NAND2_X1 U908 ( .A1(n1223), .A2(n1224), .ZN(n1043) );
OR2_X1 U909 ( .A1(n1053), .A2(KEYINPUT2), .ZN(n1224) );
INV_X1 U910 ( .A(n1198), .ZN(n1053) );
NOR2_X1 U911 ( .A1(n1078), .A2(n1219), .ZN(n1198) );
NAND3_X1 U912 ( .A1(n1219), .A2(n1225), .A3(KEYINPUT2), .ZN(n1223) );
INV_X1 U913 ( .A(n1078), .ZN(n1225) );
XOR2_X1 U914 ( .A(n1226), .B(n1142), .Z(n1078) );
INV_X1 U915 ( .A(G478), .ZN(n1142) );
NAND2_X1 U916 ( .A1(n1227), .A2(n1140), .ZN(n1226) );
NAND2_X1 U917 ( .A1(n1228), .A2(n1229), .ZN(n1140) );
OR2_X1 U918 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U919 ( .A(n1232), .B(KEYINPUT8), .Z(n1228) );
NAND2_X1 U920 ( .A1(n1231), .A2(n1233), .ZN(n1232) );
XOR2_X1 U921 ( .A(KEYINPUT42), .B(n1230), .Z(n1233) );
XNOR2_X1 U922 ( .A(n1234), .B(n1235), .ZN(n1230) );
XOR2_X1 U923 ( .A(n1236), .B(n1237), .Z(n1235) );
XNOR2_X1 U924 ( .A(n1238), .B(G107), .ZN(n1237) );
XNOR2_X1 U925 ( .A(G122), .B(n1239), .ZN(n1234) );
XOR2_X1 U926 ( .A(KEYINPUT51), .B(G134), .Z(n1239) );
NOR2_X1 U927 ( .A1(n1240), .A2(n1241), .ZN(n1231) );
INV_X1 U928 ( .A(G217), .ZN(n1240) );
INV_X1 U929 ( .A(n1079), .ZN(n1219) );
XNOR2_X1 U930 ( .A(n1242), .B(n1243), .ZN(n1079) );
XNOR2_X1 U931 ( .A(KEYINPUT47), .B(n1146), .ZN(n1243) );
INV_X1 U932 ( .A(G475), .ZN(n1146) );
OR2_X1 U933 ( .A1(n1145), .A2(G902), .ZN(n1242) );
XNOR2_X1 U934 ( .A(n1244), .B(n1245), .ZN(n1145) );
XOR2_X1 U935 ( .A(n1246), .B(n1247), .Z(n1245) );
XNOR2_X1 U936 ( .A(n1248), .B(G104), .ZN(n1247) );
XNOR2_X1 U937 ( .A(n1249), .B(G131), .ZN(n1246) );
XOR2_X1 U938 ( .A(n1250), .B(n1251), .Z(n1244) );
XOR2_X1 U939 ( .A(n1252), .B(n1253), .Z(n1251) );
NAND2_X1 U940 ( .A1(G214), .A2(n1254), .ZN(n1253) );
NAND2_X1 U941 ( .A1(n1255), .A2(KEYINPUT5), .ZN(n1252) );
XNOR2_X1 U942 ( .A(G146), .B(n1256), .ZN(n1255) );
NOR2_X1 U943 ( .A1(KEYINPUT21), .A2(n1097), .ZN(n1256) );
NAND2_X1 U944 ( .A1(KEYINPUT44), .A2(G113), .ZN(n1250) );
INV_X1 U945 ( .A(n1213), .ZN(n1071) );
XOR2_X1 U946 ( .A(n1077), .B(KEYINPUT41), .Z(n1213) );
XOR2_X1 U947 ( .A(n1257), .B(n1159), .Z(n1077) );
INV_X1 U948 ( .A(G472), .ZN(n1159) );
NAND2_X1 U949 ( .A1(n1258), .A2(n1227), .ZN(n1257) );
XNOR2_X1 U950 ( .A(n1259), .B(n1260), .ZN(n1258) );
INV_X1 U951 ( .A(n1154), .ZN(n1260) );
XOR2_X1 U952 ( .A(n1261), .B(n1262), .Z(n1154) );
NAND2_X1 U953 ( .A1(G210), .A2(n1254), .ZN(n1261) );
NOR2_X1 U954 ( .A1(G953), .A2(G237), .ZN(n1254) );
NOR2_X1 U955 ( .A1(KEYINPUT58), .A2(n1263), .ZN(n1259) );
XNOR2_X1 U956 ( .A(n1160), .B(n1155), .ZN(n1263) );
XNOR2_X1 U957 ( .A(n1264), .B(n1176), .ZN(n1155) );
XNOR2_X1 U958 ( .A(n1265), .B(n1266), .ZN(n1160) );
NOR2_X1 U959 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NOR2_X1 U960 ( .A1(n1269), .A2(n1238), .ZN(n1268) );
INV_X1 U961 ( .A(G116), .ZN(n1238) );
XOR2_X1 U962 ( .A(KEYINPUT13), .B(G113), .Z(n1269) );
NOR2_X1 U963 ( .A1(G116), .A2(n1270), .ZN(n1267) );
XOR2_X1 U964 ( .A(KEYINPUT34), .B(G113), .Z(n1270) );
XNOR2_X1 U965 ( .A(G119), .B(KEYINPUT35), .ZN(n1265) );
AND3_X1 U966 ( .A1(n1069), .A2(n1199), .A3(n1150), .ZN(n1196) );
NOR2_X1 U967 ( .A1(n1059), .A2(n1058), .ZN(n1150) );
INV_X1 U968 ( .A(n1211), .ZN(n1058) );
NAND2_X1 U969 ( .A1(n1271), .A2(G214), .ZN(n1211) );
XOR2_X1 U970 ( .A(n1272), .B(KEYINPUT29), .Z(n1271) );
NAND2_X1 U971 ( .A1(n1273), .A2(n1274), .ZN(n1059) );
NAND2_X1 U972 ( .A1(n1275), .A2(n1178), .ZN(n1274) );
NAND2_X1 U973 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND2_X1 U974 ( .A1(KEYINPUT61), .A2(n1278), .ZN(n1277) );
NAND2_X1 U975 ( .A1(n1082), .A2(n1279), .ZN(n1273) );
NAND2_X1 U976 ( .A1(KEYINPUT61), .A2(n1280), .ZN(n1279) );
NAND2_X1 U977 ( .A1(n1083), .A2(n1276), .ZN(n1280) );
INV_X1 U978 ( .A(KEYINPUT18), .ZN(n1276) );
INV_X1 U979 ( .A(n1178), .ZN(n1083) );
NAND2_X1 U980 ( .A1(G210), .A2(n1272), .ZN(n1178) );
NAND2_X1 U981 ( .A1(n1281), .A2(n1282), .ZN(n1272) );
INV_X1 U982 ( .A(G237), .ZN(n1282) );
XNOR2_X1 U983 ( .A(G902), .B(KEYINPUT33), .ZN(n1281) );
INV_X1 U984 ( .A(n1278), .ZN(n1082) );
NAND2_X1 U985 ( .A1(n1283), .A2(n1227), .ZN(n1278) );
XOR2_X1 U986 ( .A(n1284), .B(n1172), .Z(n1283) );
NAND2_X1 U987 ( .A1(n1285), .A2(n1286), .ZN(n1172) );
NAND2_X1 U988 ( .A1(n1287), .A2(n1123), .ZN(n1286) );
XOR2_X1 U989 ( .A(KEYINPUT53), .B(n1288), .Z(n1285) );
NOR2_X1 U990 ( .A1(n1287), .A2(n1123), .ZN(n1288) );
XNOR2_X1 U991 ( .A(G110), .B(n1248), .ZN(n1123) );
INV_X1 U992 ( .A(G122), .ZN(n1248) );
XOR2_X1 U993 ( .A(n1289), .B(n1120), .Z(n1287) );
XNOR2_X1 U994 ( .A(n1290), .B(n1291), .ZN(n1120) );
XNOR2_X1 U995 ( .A(G104), .B(n1292), .ZN(n1291) );
NAND2_X1 U996 ( .A1(KEYINPUT17), .A2(n1262), .ZN(n1292) );
NAND2_X1 U997 ( .A1(KEYINPUT45), .A2(n1293), .ZN(n1290) );
XNOR2_X1 U998 ( .A(KEYINPUT10), .B(n1294), .ZN(n1289) );
NOR2_X1 U999 ( .A1(KEYINPUT0), .A2(n1122), .ZN(n1294) );
NAND3_X1 U1000 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1122) );
NAND2_X1 U1001 ( .A1(KEYINPUT62), .A2(n1298), .ZN(n1297) );
INV_X1 U1002 ( .A(n1299), .ZN(n1298) );
OR3_X1 U1003 ( .A1(n1300), .A2(KEYINPUT62), .A3(G113), .ZN(n1296) );
NAND2_X1 U1004 ( .A1(G113), .A2(n1300), .ZN(n1295) );
NAND2_X1 U1005 ( .A1(KEYINPUT57), .A2(n1299), .ZN(n1300) );
XNOR2_X1 U1006 ( .A(G116), .B(n1217), .ZN(n1299) );
NAND2_X1 U1007 ( .A1(n1301), .A2(n1302), .ZN(n1284) );
NAND2_X1 U1008 ( .A1(n1177), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1009 ( .A(KEYINPUT22), .B(n1304), .Z(n1301) );
NOR2_X1 U1010 ( .A1(n1177), .A2(n1303), .ZN(n1304) );
XOR2_X1 U1011 ( .A(n1305), .B(n1306), .Z(n1303) );
XOR2_X1 U1012 ( .A(n1176), .B(KEYINPUT28), .Z(n1306) );
XNOR2_X1 U1013 ( .A(n1307), .B(n1236), .ZN(n1176) );
XNOR2_X1 U1014 ( .A(G128), .B(n1249), .ZN(n1236) );
XNOR2_X1 U1015 ( .A(G146), .B(KEYINPUT50), .ZN(n1307) );
NOR2_X1 U1016 ( .A1(n1308), .A2(G125), .ZN(n1305) );
INV_X1 U1017 ( .A(KEYINPUT3), .ZN(n1308) );
NOR2_X1 U1018 ( .A1(n1116), .A2(G953), .ZN(n1177) );
INV_X1 U1019 ( .A(G224), .ZN(n1116) );
NAND2_X1 U1020 ( .A1(n1073), .A2(n1309), .ZN(n1199) );
NAND4_X1 U1021 ( .A1(n1310), .A2(G902), .A3(n1215), .A4(n1117), .ZN(n1309) );
INV_X1 U1022 ( .A(G898), .ZN(n1117) );
XNOR2_X1 U1023 ( .A(G953), .B(KEYINPUT15), .ZN(n1310) );
NAND3_X1 U1024 ( .A1(n1215), .A2(n1087), .A3(G952), .ZN(n1073) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1215) );
NOR2_X1 U1026 ( .A1(n1068), .A2(n1067), .ZN(n1069) );
AND2_X1 U1027 ( .A1(G221), .A2(n1311), .ZN(n1067) );
INV_X1 U1028 ( .A(n1222), .ZN(n1068) );
XOR2_X1 U1029 ( .A(n1312), .B(n1164), .Z(n1222) );
INV_X1 U1030 ( .A(G469), .ZN(n1164) );
NAND2_X1 U1031 ( .A1(n1313), .A2(n1227), .ZN(n1312) );
XOR2_X1 U1032 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1033 ( .A(n1166), .B(KEYINPUT26), .Z(n1315) );
XOR2_X1 U1034 ( .A(n1316), .B(n1317), .Z(n1166) );
XNOR2_X1 U1035 ( .A(G140), .B(n1318), .ZN(n1317) );
NAND2_X1 U1036 ( .A1(G227), .A2(n1087), .ZN(n1316) );
NAND2_X1 U1037 ( .A1(n1319), .A2(n1320), .ZN(n1314) );
NAND2_X1 U1038 ( .A1(n1168), .A2(n1321), .ZN(n1320) );
INV_X1 U1039 ( .A(KEYINPUT60), .ZN(n1321) );
XNOR2_X1 U1040 ( .A(n1322), .B(n1323), .ZN(n1168) );
INV_X1 U1041 ( .A(n1264), .ZN(n1323) );
NAND3_X1 U1042 ( .A1(n1322), .A2(n1264), .A3(KEYINPUT60), .ZN(n1319) );
XNOR2_X1 U1043 ( .A(n1324), .B(n1325), .ZN(n1264) );
XNOR2_X1 U1044 ( .A(KEYINPUT11), .B(n1110), .ZN(n1325) );
INV_X1 U1045 ( .A(G137), .ZN(n1110) );
XOR2_X1 U1046 ( .A(n1326), .B(G134), .Z(n1324) );
NAND2_X1 U1047 ( .A1(KEYINPUT55), .A2(G131), .ZN(n1326) );
XNOR2_X1 U1048 ( .A(n1100), .B(n1327), .ZN(n1322) );
NOR2_X1 U1049 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NOR2_X1 U1050 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
XNOR2_X1 U1051 ( .A(KEYINPUT30), .B(n1262), .ZN(n1331) );
INV_X1 U1052 ( .A(G101), .ZN(n1262) );
AND2_X1 U1053 ( .A1(n1330), .A2(G101), .ZN(n1328) );
XOR2_X1 U1054 ( .A(n1332), .B(n1293), .Z(n1330) );
INV_X1 U1055 ( .A(G107), .ZN(n1293) );
NAND2_X1 U1056 ( .A1(KEYINPUT40), .A2(G104), .ZN(n1332) );
XOR2_X1 U1057 ( .A(n1333), .B(G128), .Z(n1100) );
NAND2_X1 U1058 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NAND2_X1 U1059 ( .A1(G146), .A2(n1249), .ZN(n1335) );
XOR2_X1 U1060 ( .A(KEYINPUT32), .B(n1336), .Z(n1334) );
NOR2_X1 U1061 ( .A1(G146), .A2(n1249), .ZN(n1336) );
INV_X1 U1062 ( .A(G143), .ZN(n1249) );
AND3_X1 U1063 ( .A1(n1337), .A2(n1338), .A3(n1339), .ZN(n1072) );
NAND2_X1 U1064 ( .A1(KEYINPUT23), .A2(n1081), .ZN(n1339) );
OR4_X1 U1065 ( .A1(KEYINPUT23), .A2(KEYINPUT37), .A3(n1081), .A4(n1080), .ZN(n1338) );
NAND2_X1 U1066 ( .A1(n1080), .A2(n1340), .ZN(n1337) );
OR2_X1 U1067 ( .A1(n1081), .A2(KEYINPUT37), .ZN(n1340) );
INV_X1 U1068 ( .A(n1135), .ZN(n1081) );
NAND2_X1 U1069 ( .A1(G217), .A2(n1311), .ZN(n1135) );
NAND2_X1 U1070 ( .A1(G234), .A2(n1227), .ZN(n1311) );
INV_X1 U1071 ( .A(G902), .ZN(n1227) );
NOR2_X1 U1072 ( .A1(n1138), .A2(G902), .ZN(n1080) );
INV_X1 U1073 ( .A(n1134), .ZN(n1138) );
XNOR2_X1 U1074 ( .A(n1341), .B(n1342), .ZN(n1134) );
XNOR2_X1 U1075 ( .A(n1343), .B(n1344), .ZN(n1342) );
XOR2_X1 U1076 ( .A(n1345), .B(n1346), .Z(n1344) );
NOR2_X1 U1077 ( .A1(n1241), .A2(n1347), .ZN(n1346) );
INV_X1 U1078 ( .A(G221), .ZN(n1347) );
NAND2_X1 U1079 ( .A1(G234), .A2(n1087), .ZN(n1241) );
INV_X1 U1080 ( .A(G953), .ZN(n1087) );
NAND2_X1 U1081 ( .A1(n1348), .A2(KEYINPUT1), .ZN(n1345) );
XOR2_X1 U1082 ( .A(n1349), .B(n1350), .Z(n1348) );
XNOR2_X1 U1083 ( .A(G128), .B(n1217), .ZN(n1350) );
INV_X1 U1084 ( .A(G119), .ZN(n1217) );
NAND2_X1 U1085 ( .A1(KEYINPUT31), .A2(n1318), .ZN(n1349) );
INV_X1 U1086 ( .A(G110), .ZN(n1318) );
INV_X1 U1087 ( .A(n1097), .ZN(n1343) );
XNOR2_X1 U1088 ( .A(G140), .B(G125), .ZN(n1097) );
XNOR2_X1 U1089 ( .A(G137), .B(n1351), .ZN(n1341) );
XOR2_X1 U1090 ( .A(KEYINPUT20), .B(G146), .Z(n1351) );
endmodule


