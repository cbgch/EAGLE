//Key = 1101010100101100100011111101101101000101011100101111000101110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342;

XOR2_X1 U739 ( .A(n1031), .B(n1032), .Z(G9) );
NAND2_X1 U740 ( .A1(KEYINPUT27), .A2(n1033), .ZN(n1032) );
INV_X1 U741 ( .A(n1034), .ZN(n1033) );
NAND4_X1 U742 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(G75) );
INV_X1 U743 ( .A(n1039), .ZN(n1038) );
NAND4_X1 U744 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1037) );
NOR4_X1 U745 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
XOR2_X1 U746 ( .A(n1048), .B(KEYINPUT3), .Z(n1047) );
NAND2_X1 U747 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U748 ( .A1(n1049), .A2(n1050), .ZN(n1046) );
NOR2_X1 U749 ( .A1(n1051), .A2(n1052), .ZN(n1042) );
XOR2_X1 U750 ( .A(n1053), .B(KEYINPUT6), .Z(n1041) );
NAND2_X1 U751 ( .A1(G952), .A2(n1054), .ZN(n1036) );
NAND4_X1 U752 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NAND4_X1 U753 ( .A1(n1053), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1058) );
NAND3_X1 U754 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1060) );
INV_X1 U755 ( .A(n1065), .ZN(n1062) );
NAND2_X1 U756 ( .A1(n1066), .A2(n1067), .ZN(n1059) );
NAND2_X1 U757 ( .A1(n1068), .A2(n1065), .ZN(n1066) );
NAND2_X1 U758 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
NAND2_X1 U759 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U760 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND3_X1 U761 ( .A1(n1063), .A2(n1067), .A3(n1075), .ZN(n1074) );
INV_X1 U762 ( .A(KEYINPUT61), .ZN(n1067) );
NAND3_X1 U763 ( .A1(n1076), .A2(n1077), .A3(n1045), .ZN(n1073) );
XOR2_X1 U764 ( .A(KEYINPUT62), .B(n1075), .Z(n1077) );
XOR2_X1 U765 ( .A(n1040), .B(n1078), .Z(n1076) );
NAND2_X1 U766 ( .A1(n1079), .A2(n1080), .ZN(n1069) );
NAND3_X1 U767 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1080) );
NAND2_X1 U768 ( .A1(n1084), .A2(n1071), .ZN(n1083) );
NAND2_X1 U769 ( .A1(n1085), .A2(n1086), .ZN(n1082) );
XOR2_X1 U770 ( .A(KEYINPUT4), .B(n1071), .Z(n1086) );
NAND2_X1 U771 ( .A1(n1075), .A2(n1087), .ZN(n1081) );
NAND2_X1 U772 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U773 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
INV_X1 U774 ( .A(n1092), .ZN(n1088) );
NAND3_X1 U775 ( .A1(n1079), .A2(n1093), .A3(n1064), .ZN(n1057) );
AND3_X1 U776 ( .A1(n1068), .A2(n1071), .A3(n1075), .ZN(n1064) );
INV_X1 U777 ( .A(n1094), .ZN(n1068) );
NAND2_X1 U778 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NAND2_X1 U779 ( .A1(n1044), .A2(n1053), .ZN(n1096) );
NAND2_X1 U780 ( .A1(KEYINPUT19), .A2(n1097), .ZN(n1056) );
OR2_X1 U781 ( .A1(n1097), .A2(KEYINPUT19), .ZN(n1035) );
XOR2_X1 U782 ( .A(n1098), .B(n1099), .Z(G72) );
NOR2_X1 U783 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XOR2_X1 U784 ( .A(n1102), .B(KEYINPUT10), .Z(n1101) );
NAND3_X1 U785 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
NAND2_X1 U786 ( .A1(G953), .A2(n1106), .ZN(n1104) );
XOR2_X1 U787 ( .A(KEYINPUT40), .B(n1107), .Z(n1103) );
NOR3_X1 U788 ( .A1(n1105), .A2(G953), .A3(n1107), .ZN(n1100) );
XOR2_X1 U789 ( .A(n1108), .B(n1109), .Z(n1105) );
XOR2_X1 U790 ( .A(KEYINPUT38), .B(G125), .Z(n1109) );
XOR2_X1 U791 ( .A(n1110), .B(n1111), .Z(n1108) );
NOR2_X1 U792 ( .A1(KEYINPUT34), .A2(n1112), .ZN(n1111) );
INV_X1 U793 ( .A(n1113), .ZN(n1112) );
NAND2_X1 U794 ( .A1(G953), .A2(n1114), .ZN(n1098) );
NAND2_X1 U795 ( .A1(G900), .A2(G227), .ZN(n1114) );
XOR2_X1 U796 ( .A(n1115), .B(n1116), .Z(G69) );
XOR2_X1 U797 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U798 ( .A1(n1119), .A2(G953), .ZN(n1118) );
NOR3_X1 U799 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1117) );
NOR2_X1 U800 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
INV_X1 U801 ( .A(n1125), .ZN(n1124) );
NOR2_X1 U802 ( .A1(n1125), .A2(n1126), .ZN(n1121) );
NOR2_X1 U803 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U804 ( .A1(KEYINPUT41), .A2(n1129), .ZN(n1128) );
AND2_X1 U805 ( .A1(n1123), .A2(KEYINPUT41), .ZN(n1127) );
NAND2_X1 U806 ( .A1(KEYINPUT33), .A2(n1130), .ZN(n1123) );
INV_X1 U807 ( .A(n1129), .ZN(n1130) );
NOR2_X1 U808 ( .A1(G898), .A2(n1097), .ZN(n1120) );
NOR2_X1 U809 ( .A1(n1131), .A2(n1097), .ZN(n1115) );
AND2_X1 U810 ( .A1(G224), .A2(G898), .ZN(n1131) );
NOR2_X1 U811 ( .A1(n1039), .A2(n1132), .ZN(G66) );
XOR2_X1 U812 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR3_X1 U813 ( .A1(n1135), .A2(KEYINPUT2), .A3(n1136), .ZN(n1133) );
NOR2_X1 U814 ( .A1(n1039), .A2(n1137), .ZN(G63) );
NOR3_X1 U815 ( .A1(n1138), .A2(n1049), .A3(n1139), .ZN(n1137) );
NOR2_X1 U816 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR2_X1 U817 ( .A1(n1055), .A2(n1050), .ZN(n1140) );
INV_X1 U818 ( .A(G478), .ZN(n1050) );
XOR2_X1 U819 ( .A(KEYINPUT47), .B(n1142), .Z(n1138) );
AND3_X1 U820 ( .A1(n1143), .A2(G478), .A3(n1141), .ZN(n1142) );
NOR2_X1 U821 ( .A1(n1039), .A2(n1144), .ZN(G60) );
XNOR2_X1 U822 ( .A(n1145), .B(n1146), .ZN(n1144) );
AND2_X1 U823 ( .A1(G475), .A2(n1143), .ZN(n1146) );
XOR2_X1 U824 ( .A(n1147), .B(n1148), .Z(G6) );
NAND2_X1 U825 ( .A1(KEYINPUT16), .A2(G104), .ZN(n1148) );
NOR2_X1 U826 ( .A1(n1039), .A2(n1149), .ZN(G57) );
XOR2_X1 U827 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U828 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U829 ( .A(n1154), .B(n1155), .Z(n1153) );
AND2_X1 U830 ( .A1(G472), .A2(n1143), .ZN(n1155) );
NOR3_X1 U831 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1154) );
NOR2_X1 U832 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U833 ( .A1(n1161), .A2(n1162), .ZN(n1159) );
INV_X1 U834 ( .A(KEYINPUT30), .ZN(n1162) );
XOR2_X1 U835 ( .A(n1163), .B(KEYINPUT21), .Z(n1161) );
AND3_X1 U836 ( .A1(n1160), .A2(n1163), .A3(KEYINPUT30), .ZN(n1157) );
NOR2_X1 U837 ( .A1(KEYINPUT30), .A2(n1163), .ZN(n1156) );
NOR2_X1 U838 ( .A1(KEYINPUT26), .A2(n1164), .ZN(n1152) );
XOR2_X1 U839 ( .A(n1165), .B(n1166), .Z(n1150) );
XOR2_X1 U840 ( .A(KEYINPUT14), .B(G101), .Z(n1166) );
NOR2_X1 U841 ( .A1(n1039), .A2(n1167), .ZN(G54) );
XOR2_X1 U842 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U844 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
INV_X1 U845 ( .A(n1174), .ZN(n1173) );
XOR2_X1 U846 ( .A(n1175), .B(KEYINPUT45), .Z(n1172) );
XNOR2_X1 U847 ( .A(KEYINPUT58), .B(n1176), .ZN(n1168) );
NOR2_X1 U848 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR2_X1 U849 ( .A1(n1179), .A2(KEYINPUT18), .ZN(n1178) );
NOR2_X1 U850 ( .A1(n1180), .A2(n1135), .ZN(n1179) );
NOR3_X1 U851 ( .A1(n1135), .A2(KEYINPUT42), .A3(n1180), .ZN(n1177) );
INV_X1 U852 ( .A(n1143), .ZN(n1135) );
NOR2_X1 U853 ( .A1(n1039), .A2(n1181), .ZN(G51) );
XOR2_X1 U854 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U855 ( .A(G125), .B(n1184), .Z(n1183) );
NOR2_X1 U856 ( .A1(KEYINPUT29), .A2(n1185), .ZN(n1184) );
INV_X1 U857 ( .A(n1163), .ZN(n1185) );
XOR2_X1 U858 ( .A(n1186), .B(n1187), .Z(n1182) );
NAND3_X1 U859 ( .A1(n1143), .A2(G210), .A3(KEYINPUT1), .ZN(n1186) );
NOR2_X1 U860 ( .A1(n1188), .A2(n1055), .ZN(n1143) );
AND2_X1 U861 ( .A1(n1107), .A2(n1119), .ZN(n1055) );
AND4_X1 U862 ( .A1(n1147), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1119) );
AND4_X1 U863 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1034), .ZN(n1191) );
NAND3_X1 U864 ( .A1(n1195), .A2(n1071), .A3(n1085), .ZN(n1034) );
AND2_X1 U865 ( .A1(n1196), .A2(n1197), .ZN(n1190) );
NAND3_X1 U866 ( .A1(n1195), .A2(n1071), .A3(n1084), .ZN(n1147) );
AND4_X1 U867 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1107) );
NOR4_X1 U868 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
NOR2_X1 U869 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
XNOR2_X1 U870 ( .A(n1084), .B(KEYINPUT8), .ZN(n1206) );
INV_X1 U871 ( .A(n1208), .ZN(n1202) );
NOR2_X1 U872 ( .A1(n1209), .A2(n1210), .ZN(n1200) );
NOR2_X1 U873 ( .A1(n1097), .A2(G952), .ZN(n1039) );
XOR2_X1 U874 ( .A(G146), .B(n1204), .Z(G48) );
AND3_X1 U875 ( .A1(n1211), .A2(n1084), .A3(n1212), .ZN(n1204) );
XOR2_X1 U876 ( .A(n1199), .B(n1213), .Z(G45) );
XOR2_X1 U877 ( .A(KEYINPUT22), .B(G143), .Z(n1213) );
NAND4_X1 U878 ( .A1(n1211), .A2(n1092), .A3(n1214), .A4(n1052), .ZN(n1199) );
XOR2_X1 U879 ( .A(G140), .B(n1203), .Z(G42) );
AND2_X1 U880 ( .A1(n1215), .A2(n1216), .ZN(n1203) );
NAND2_X1 U881 ( .A1(n1217), .A2(n1218), .ZN(G39) );
NAND2_X1 U882 ( .A1(G137), .A2(n1208), .ZN(n1218) );
XOR2_X1 U883 ( .A(KEYINPUT20), .B(n1219), .Z(n1217) );
NOR2_X1 U884 ( .A1(G137), .A2(n1208), .ZN(n1219) );
NAND3_X1 U885 ( .A1(n1212), .A2(n1075), .A3(n1215), .ZN(n1208) );
XNOR2_X1 U886 ( .A(n1210), .B(n1220), .ZN(G36) );
NAND2_X1 U887 ( .A1(KEYINPUT50), .A2(G134), .ZN(n1220) );
AND2_X1 U888 ( .A1(n1221), .A2(n1085), .ZN(n1210) );
XNOR2_X1 U889 ( .A(G131), .B(n1222), .ZN(G33) );
NAND2_X1 U890 ( .A1(n1221), .A2(n1084), .ZN(n1222) );
INV_X1 U891 ( .A(n1207), .ZN(n1221) );
NAND2_X1 U892 ( .A1(n1215), .A2(n1092), .ZN(n1207) );
AND4_X1 U893 ( .A1(n1053), .A2(n1063), .A3(n1223), .A4(n1061), .ZN(n1215) );
XOR2_X1 U894 ( .A(G128), .B(n1209), .Z(G30) );
AND3_X1 U895 ( .A1(n1211), .A2(n1085), .A3(n1212), .ZN(n1209) );
AND3_X1 U896 ( .A1(n1224), .A2(n1223), .A3(n1063), .ZN(n1211) );
XOR2_X1 U897 ( .A(n1225), .B(n1194), .Z(G3) );
NAND3_X1 U898 ( .A1(n1075), .A2(n1195), .A3(n1092), .ZN(n1194) );
XOR2_X1 U899 ( .A(n1226), .B(n1198), .Z(G27) );
NAND4_X1 U900 ( .A1(n1216), .A2(n1224), .A3(n1079), .A4(n1223), .ZN(n1198) );
NAND2_X1 U901 ( .A1(n1094), .A2(n1227), .ZN(n1223) );
NAND4_X1 U902 ( .A1(G902), .A2(G953), .A3(n1228), .A4(n1106), .ZN(n1227) );
INV_X1 U903 ( .A(G900), .ZN(n1106) );
AND3_X1 U904 ( .A1(n1090), .A2(n1091), .A3(n1084), .ZN(n1216) );
XNOR2_X1 U905 ( .A(G122), .B(n1189), .ZN(G24) );
NAND4_X1 U906 ( .A1(n1229), .A2(n1071), .A3(n1214), .A4(n1052), .ZN(n1189) );
INV_X1 U907 ( .A(n1051), .ZN(n1071) );
NAND2_X1 U908 ( .A1(n1230), .A2(n1090), .ZN(n1051) );
XOR2_X1 U909 ( .A(n1231), .B(n1197), .Z(G21) );
NAND3_X1 U910 ( .A1(n1212), .A2(n1075), .A3(n1229), .ZN(n1197) );
NOR2_X1 U911 ( .A1(n1090), .A2(n1230), .ZN(n1212) );
XNOR2_X1 U912 ( .A(G116), .B(n1193), .ZN(G18) );
NAND3_X1 U913 ( .A1(n1092), .A2(n1085), .A3(n1229), .ZN(n1193) );
AND2_X1 U914 ( .A1(n1232), .A2(n1214), .ZN(n1085) );
XNOR2_X1 U915 ( .A(G113), .B(n1192), .ZN(G15) );
NAND3_X1 U916 ( .A1(n1092), .A2(n1084), .A3(n1229), .ZN(n1192) );
AND2_X1 U917 ( .A1(n1233), .A2(n1079), .ZN(n1229) );
NAND2_X1 U918 ( .A1(n1234), .A2(n1235), .ZN(n1079) );
NAND2_X1 U919 ( .A1(n1063), .A2(n1078), .ZN(n1235) );
INV_X1 U920 ( .A(KEYINPUT37), .ZN(n1078) );
NAND3_X1 U921 ( .A1(n1040), .A2(n1236), .A3(KEYINPUT37), .ZN(n1234) );
NOR2_X1 U922 ( .A1(n1214), .A2(n1232), .ZN(n1084) );
NOR2_X1 U923 ( .A1(n1091), .A2(n1090), .ZN(n1092) );
XOR2_X1 U924 ( .A(n1237), .B(G110), .Z(G12) );
NAND2_X1 U925 ( .A1(KEYINPUT39), .A2(n1196), .ZN(n1237) );
NAND4_X1 U926 ( .A1(n1075), .A2(n1195), .A3(n1090), .A4(n1091), .ZN(n1196) );
INV_X1 U927 ( .A(n1230), .ZN(n1091) );
XNOR2_X1 U928 ( .A(n1238), .B(n1136), .ZN(n1230) );
NAND2_X1 U929 ( .A1(G217), .A2(n1239), .ZN(n1136) );
OR2_X1 U930 ( .A1(n1134), .A2(G902), .ZN(n1238) );
XNOR2_X1 U931 ( .A(n1240), .B(n1241), .ZN(n1134) );
XOR2_X1 U932 ( .A(G110), .B(n1242), .Z(n1241) );
XOR2_X1 U933 ( .A(KEYINPUT57), .B(G119), .Z(n1242) );
XOR2_X1 U934 ( .A(n1243), .B(n1244), .Z(n1240) );
XNOR2_X1 U935 ( .A(n1245), .B(n1246), .ZN(n1243) );
NAND3_X1 U936 ( .A1(n1247), .A2(n1248), .A3(KEYINPUT55), .ZN(n1246) );
NAND2_X1 U937 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
NAND2_X1 U938 ( .A1(n1251), .A2(n1252), .ZN(n1249) );
INV_X1 U939 ( .A(n1253), .ZN(n1251) );
NAND2_X1 U940 ( .A1(G146), .A2(n1254), .ZN(n1247) );
XOR2_X1 U941 ( .A(G140), .B(n1226), .Z(n1254) );
NAND2_X1 U942 ( .A1(n1255), .A2(KEYINPUT49), .ZN(n1245) );
XNOR2_X1 U943 ( .A(G137), .B(n1256), .ZN(n1255) );
AND3_X1 U944 ( .A1(G221), .A2(n1097), .A3(G234), .ZN(n1256) );
XOR2_X1 U945 ( .A(n1257), .B(G472), .Z(n1090) );
NAND2_X1 U946 ( .A1(n1258), .A2(n1188), .ZN(n1257) );
XOR2_X1 U947 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U948 ( .A(KEYINPUT25), .B(G101), .Z(n1260) );
XNOR2_X1 U949 ( .A(n1261), .B(n1164), .ZN(n1259) );
OR3_X1 U950 ( .A1(G237), .A2(G953), .A3(n1262), .ZN(n1164) );
NAND2_X1 U951 ( .A1(KEYINPUT31), .A2(n1263), .ZN(n1261) );
XOR2_X1 U952 ( .A(n1163), .B(n1264), .Z(n1263) );
XOR2_X1 U953 ( .A(n1165), .B(n1265), .Z(n1264) );
NOR2_X1 U954 ( .A1(KEYINPUT54), .A2(n1160), .ZN(n1265) );
NAND2_X1 U955 ( .A1(n1266), .A2(n1267), .ZN(n1165) );
NAND2_X1 U956 ( .A1(G113), .A2(n1268), .ZN(n1267) );
XOR2_X1 U957 ( .A(n1269), .B(KEYINPUT44), .Z(n1266) );
OR2_X1 U958 ( .A1(n1268), .A2(G113), .ZN(n1269) );
XOR2_X1 U959 ( .A(G116), .B(G119), .Z(n1268) );
AND2_X1 U960 ( .A1(n1233), .A2(n1063), .ZN(n1195) );
NOR2_X1 U961 ( .A1(n1040), .A2(n1045), .ZN(n1063) );
INV_X1 U962 ( .A(n1236), .ZN(n1045) );
NAND2_X1 U963 ( .A1(G221), .A2(n1239), .ZN(n1236) );
NAND2_X1 U964 ( .A1(n1270), .A2(n1188), .ZN(n1239) );
XNOR2_X1 U965 ( .A(G234), .B(KEYINPUT28), .ZN(n1270) );
AND2_X1 U966 ( .A1(n1271), .A2(n1272), .ZN(n1040) );
NAND2_X1 U967 ( .A1(G469), .A2(n1273), .ZN(n1272) );
NAND2_X1 U968 ( .A1(n1274), .A2(n1188), .ZN(n1273) );
NAND3_X1 U969 ( .A1(n1274), .A2(n1188), .A3(n1180), .ZN(n1271) );
INV_X1 U970 ( .A(G469), .ZN(n1180) );
XNOR2_X1 U971 ( .A(n1275), .B(n1276), .ZN(n1274) );
XOR2_X1 U972 ( .A(KEYINPUT7), .B(KEYINPUT5), .Z(n1276) );
XNOR2_X1 U973 ( .A(n1171), .B(n1277), .ZN(n1275) );
NOR2_X1 U974 ( .A1(n1174), .A2(n1278), .ZN(n1277) );
XOR2_X1 U975 ( .A(n1175), .B(KEYINPUT63), .Z(n1278) );
NAND2_X1 U976 ( .A1(n1279), .A2(n1113), .ZN(n1175) );
NOR2_X1 U977 ( .A1(n1113), .A2(n1279), .ZN(n1174) );
XOR2_X1 U978 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U979 ( .A(G104), .B(G101), .Z(n1281) );
XOR2_X1 U980 ( .A(n1282), .B(G107), .Z(n1280) );
XNOR2_X1 U981 ( .A(KEYINPUT56), .B(KEYINPUT23), .ZN(n1282) );
XNOR2_X1 U982 ( .A(n1283), .B(n1284), .ZN(n1113) );
XOR2_X1 U983 ( .A(KEYINPUT46), .B(n1244), .Z(n1284) );
XNOR2_X1 U984 ( .A(n1110), .B(n1285), .ZN(n1171) );
XOR2_X1 U985 ( .A(G110), .B(n1286), .Z(n1285) );
AND2_X1 U986 ( .A1(n1097), .A2(G227), .ZN(n1286) );
XOR2_X1 U987 ( .A(n1160), .B(G140), .Z(n1110) );
XNOR2_X1 U988 ( .A(G131), .B(n1287), .ZN(n1160) );
XOR2_X1 U989 ( .A(G137), .B(G134), .Z(n1287) );
AND2_X1 U990 ( .A1(n1224), .A2(n1288), .ZN(n1233) );
NAND2_X1 U991 ( .A1(n1094), .A2(n1289), .ZN(n1288) );
NAND4_X1 U992 ( .A1(G902), .A2(G953), .A3(n1228), .A4(n1290), .ZN(n1289) );
INV_X1 U993 ( .A(G898), .ZN(n1290) );
NAND3_X1 U994 ( .A1(n1228), .A2(n1097), .A3(G952), .ZN(n1094) );
NAND2_X1 U995 ( .A1(G237), .A2(G234), .ZN(n1228) );
INV_X1 U996 ( .A(n1095), .ZN(n1224) );
NAND2_X1 U997 ( .A1(n1291), .A2(n1061), .ZN(n1095) );
INV_X1 U998 ( .A(n1044), .ZN(n1061) );
NOR2_X1 U999 ( .A1(n1292), .A2(n1293), .ZN(n1044) );
INV_X1 U1000 ( .A(n1053), .ZN(n1291) );
XOR2_X1 U1001 ( .A(n1294), .B(n1295), .Z(n1053) );
NOR2_X1 U1002 ( .A1(n1293), .A2(n1262), .ZN(n1295) );
INV_X1 U1003 ( .A(G210), .ZN(n1262) );
NOR2_X1 U1004 ( .A1(G902), .A2(G237), .ZN(n1293) );
NAND2_X1 U1005 ( .A1(n1296), .A2(n1188), .ZN(n1294) );
XNOR2_X1 U1006 ( .A(n1187), .B(n1297), .ZN(n1296) );
XOR2_X1 U1007 ( .A(n1226), .B(n1163), .Z(n1297) );
XOR2_X1 U1008 ( .A(n1298), .B(n1244), .Z(n1163) );
NAND2_X1 U1009 ( .A1(KEYINPUT48), .A2(n1283), .ZN(n1298) );
XOR2_X1 U1010 ( .A(G143), .B(G146), .Z(n1283) );
XNOR2_X1 U1011 ( .A(n1299), .B(n1125), .ZN(n1187) );
XOR2_X1 U1012 ( .A(G110), .B(G122), .Z(n1125) );
XOR2_X1 U1013 ( .A(n1300), .B(n1301), .Z(n1299) );
NOR2_X1 U1014 ( .A1(KEYINPUT60), .A2(n1129), .ZN(n1301) );
XOR2_X1 U1015 ( .A(n1302), .B(n1303), .Z(n1129) );
XOR2_X1 U1016 ( .A(n1304), .B(n1305), .Z(n1303) );
NOR2_X1 U1017 ( .A1(KEYINPUT9), .A2(n1031), .ZN(n1305) );
NOR2_X1 U1018 ( .A1(n1306), .A2(n1307), .ZN(n1304) );
XOR2_X1 U1019 ( .A(n1308), .B(KEYINPUT51), .Z(n1307) );
NAND3_X1 U1020 ( .A1(n1309), .A2(n1310), .A3(G113), .ZN(n1308) );
NAND2_X1 U1021 ( .A1(G119), .A2(n1311), .ZN(n1310) );
NAND2_X1 U1022 ( .A1(n1312), .A2(n1231), .ZN(n1309) );
INV_X1 U1023 ( .A(G119), .ZN(n1231) );
XNOR2_X1 U1024 ( .A(KEYINPUT36), .B(n1311), .ZN(n1312) );
NOR2_X1 U1025 ( .A1(G113), .A2(n1313), .ZN(n1306) );
XNOR2_X1 U1026 ( .A(n1314), .B(n1311), .ZN(n1313) );
XNOR2_X1 U1027 ( .A(G116), .B(KEYINPUT0), .ZN(n1311) );
NOR2_X1 U1028 ( .A1(G119), .A2(KEYINPUT36), .ZN(n1314) );
XOR2_X1 U1029 ( .A(n1225), .B(n1315), .Z(n1302) );
XOR2_X1 U1030 ( .A(KEYINPUT59), .B(G104), .Z(n1315) );
INV_X1 U1031 ( .A(G101), .ZN(n1225) );
NAND2_X1 U1032 ( .A1(n1316), .A2(G224), .ZN(n1300) );
XOR2_X1 U1033 ( .A(n1097), .B(KEYINPUT52), .Z(n1316) );
NOR2_X1 U1034 ( .A1(n1052), .A2(n1214), .ZN(n1075) );
XNOR2_X1 U1035 ( .A(n1049), .B(n1317), .ZN(n1214) );
XOR2_X1 U1036 ( .A(KEYINPUT12), .B(G478), .Z(n1317) );
NOR2_X1 U1037 ( .A1(n1141), .A2(G902), .ZN(n1049) );
XOR2_X1 U1038 ( .A(n1318), .B(n1319), .Z(n1141) );
XOR2_X1 U1039 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1040 ( .A(n1322), .B(n1323), .Z(n1321) );
NAND3_X1 U1041 ( .A1(n1324), .A2(n1097), .A3(G217), .ZN(n1323) );
INV_X1 U1042 ( .A(G953), .ZN(n1097) );
XOR2_X1 U1043 ( .A(KEYINPUT35), .B(G234), .Z(n1324) );
NAND2_X1 U1044 ( .A1(n1325), .A2(KEYINPUT13), .ZN(n1322) );
XNOR2_X1 U1045 ( .A(G116), .B(n1326), .ZN(n1325) );
NOR2_X1 U1046 ( .A1(G122), .A2(KEYINPUT53), .ZN(n1326) );
NOR2_X1 U1047 ( .A1(n1327), .A2(n1328), .ZN(n1320) );
NOR2_X1 U1048 ( .A1(KEYINPUT32), .A2(n1244), .ZN(n1328) );
INV_X1 U1049 ( .A(n1329), .ZN(n1244) );
NOR2_X1 U1050 ( .A1(KEYINPUT24), .A2(n1329), .ZN(n1327) );
XNOR2_X1 U1051 ( .A(G128), .B(KEYINPUT15), .ZN(n1329) );
XOR2_X1 U1052 ( .A(n1031), .B(n1330), .Z(n1318) );
XOR2_X1 U1053 ( .A(G143), .B(G134), .Z(n1330) );
INV_X1 U1054 ( .A(G107), .ZN(n1031) );
INV_X1 U1055 ( .A(n1232), .ZN(n1052) );
XOR2_X1 U1056 ( .A(n1331), .B(G475), .Z(n1232) );
NAND2_X1 U1057 ( .A1(n1145), .A2(n1188), .ZN(n1331) );
INV_X1 U1058 ( .A(G902), .ZN(n1188) );
XNOR2_X1 U1059 ( .A(n1332), .B(n1333), .ZN(n1145) );
XOR2_X1 U1060 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1061 ( .A(G104), .B(n1336), .Z(n1335) );
NOR2_X1 U1062 ( .A1(KEYINPUT11), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1063 ( .A(n1338), .B(n1339), .Z(n1337) );
XOR2_X1 U1064 ( .A(KEYINPUT17), .B(G143), .Z(n1339) );
NOR3_X1 U1065 ( .A1(n1292), .A2(G953), .A3(G237), .ZN(n1338) );
INV_X1 U1066 ( .A(G214), .ZN(n1292) );
NOR2_X1 U1067 ( .A1(n1253), .A2(n1340), .ZN(n1334) );
XOR2_X1 U1068 ( .A(n1252), .B(KEYINPUT43), .Z(n1340) );
NAND2_X1 U1069 ( .A1(G140), .A2(n1226), .ZN(n1252) );
NOR2_X1 U1070 ( .A1(n1226), .A2(G140), .ZN(n1253) );
INV_X1 U1071 ( .A(G125), .ZN(n1226) );
XOR2_X1 U1072 ( .A(n1341), .B(n1342), .Z(n1332) );
XOR2_X1 U1073 ( .A(G122), .B(G113), .Z(n1342) );
XOR2_X1 U1074 ( .A(G131), .B(n1250), .Z(n1341) );
INV_X1 U1075 ( .A(G146), .ZN(n1250) );
endmodule


