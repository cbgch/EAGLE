//Key = 1011011111000001001110010111000100000001001111000101001011010110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;

XNOR2_X1 U775 ( .A(G107), .B(n1069), .ZN(G9) );
NOR2_X1 U776 ( .A1(n1070), .A2(n1071), .ZN(G75) );
NOR3_X1 U777 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
NAND3_X1 U778 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1072) );
NAND2_X1 U779 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U780 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U781 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U782 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U783 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U784 ( .A1(n1088), .A2(n1089), .ZN(n1080) );
NAND2_X1 U785 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U786 ( .A1(n1082), .A2(n1092), .ZN(n1091) );
NAND2_X1 U787 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U788 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U789 ( .A1(n1086), .A2(n1097), .ZN(n1090) );
NAND3_X1 U790 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1097) );
NAND2_X1 U791 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND3_X1 U792 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1099) );
XNOR2_X1 U793 ( .A(n1101), .B(KEYINPUT31), .ZN(n1105) );
NAND2_X1 U794 ( .A1(n1106), .A2(n1107), .ZN(n1098) );
NAND2_X1 U795 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
INV_X1 U796 ( .A(n1110), .ZN(n1078) );
NOR3_X1 U797 ( .A1(n1111), .A2(G953), .A3(G952), .ZN(n1070) );
INV_X1 U798 ( .A(n1075), .ZN(n1111) );
NAND3_X1 U799 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1075) );
NOR3_X1 U800 ( .A1(n1115), .A2(n1095), .A3(n1103), .ZN(n1114) );
NOR3_X1 U801 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
AND2_X1 U802 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NOR3_X1 U803 ( .A1(n1120), .A2(KEYINPUT53), .A3(n1119), .ZN(n1117) );
NAND2_X1 U804 ( .A1(KEYINPUT54), .A2(n1121), .ZN(n1119) );
NOR2_X1 U805 ( .A1(n1121), .A2(n1122), .ZN(n1116) );
INV_X1 U806 ( .A(KEYINPUT53), .ZN(n1122) );
XOR2_X1 U807 ( .A(KEYINPUT58), .B(n1123), .Z(n1113) );
NOR3_X1 U808 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
XOR2_X1 U809 ( .A(n1127), .B(n1128), .Z(n1125) );
XNOR2_X1 U810 ( .A(KEYINPUT61), .B(n1129), .ZN(n1128) );
XNOR2_X1 U811 ( .A(n1130), .B(n1131), .ZN(n1112) );
NAND2_X1 U812 ( .A1(KEYINPUT42), .A2(G469), .ZN(n1130) );
XOR2_X1 U813 ( .A(n1132), .B(n1133), .Z(G72) );
NOR2_X1 U814 ( .A1(n1134), .A2(n1076), .ZN(n1133) );
NOR2_X1 U815 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U816 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
NAND3_X1 U817 ( .A1(n1073), .A2(n1076), .A3(n1139), .ZN(n1138) );
NAND2_X1 U818 ( .A1(n1140), .A2(n1141), .ZN(n1137) );
NAND2_X1 U819 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U820 ( .A1(n1144), .A2(n1076), .ZN(n1143) );
NAND2_X1 U821 ( .A1(n1145), .A2(G953), .ZN(n1142) );
XNOR2_X1 U822 ( .A(G900), .B(KEYINPUT9), .ZN(n1145) );
INV_X1 U823 ( .A(n1139), .ZN(n1140) );
NAND2_X1 U824 ( .A1(n1146), .A2(n1147), .ZN(n1139) );
XOR2_X1 U825 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U826 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U827 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U828 ( .A(KEYINPUT29), .B(n1154), .Z(n1153) );
AND2_X1 U829 ( .A1(n1155), .A2(G140), .ZN(n1154) );
NOR2_X1 U830 ( .A1(G140), .A2(n1155), .ZN(n1152) );
NOR2_X1 U831 ( .A1(KEYINPUT60), .A2(n1156), .ZN(n1150) );
XNOR2_X1 U832 ( .A(G131), .B(n1157), .ZN(n1156) );
NOR2_X1 U833 ( .A1(KEYINPUT63), .A2(n1158), .ZN(n1157) );
XOR2_X1 U834 ( .A(KEYINPUT40), .B(KEYINPUT26), .Z(n1146) );
NAND2_X1 U835 ( .A1(n1159), .A2(n1160), .ZN(G69) );
NAND2_X1 U836 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U837 ( .A1(G953), .A2(n1163), .ZN(n1162) );
NAND3_X1 U838 ( .A1(G953), .A2(n1164), .A3(n1165), .ZN(n1159) );
INV_X1 U839 ( .A(n1161), .ZN(n1165) );
XNOR2_X1 U840 ( .A(n1166), .B(n1167), .ZN(n1161) );
NOR3_X1 U841 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1167) );
NOR2_X1 U842 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XNOR2_X1 U843 ( .A(n1173), .B(KEYINPUT44), .ZN(n1172) );
INV_X1 U844 ( .A(n1174), .ZN(n1171) );
NOR2_X1 U845 ( .A1(n1174), .A2(n1175), .ZN(n1169) );
XNOR2_X1 U846 ( .A(n1173), .B(KEYINPUT11), .ZN(n1175) );
XOR2_X1 U847 ( .A(n1176), .B(n1177), .Z(n1174) );
NAND3_X1 U848 ( .A1(n1074), .A2(n1076), .A3(KEYINPUT56), .ZN(n1166) );
NAND2_X1 U849 ( .A1(G898), .A2(G224), .ZN(n1164) );
NOR2_X1 U850 ( .A1(n1178), .A2(n1179), .ZN(G66) );
XOR2_X1 U851 ( .A(n1180), .B(n1181), .Z(n1179) );
NAND3_X1 U852 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1180) );
XOR2_X1 U853 ( .A(n1185), .B(KEYINPUT47), .Z(n1184) );
NOR2_X1 U854 ( .A1(n1178), .A2(n1186), .ZN(G63) );
NOR2_X1 U855 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U856 ( .A(n1189), .B(n1190), .Z(n1188) );
AND2_X1 U857 ( .A1(G478), .A2(n1191), .ZN(n1190) );
AND2_X1 U858 ( .A1(n1192), .A2(KEYINPUT5), .ZN(n1189) );
NOR2_X1 U859 ( .A1(KEYINPUT5), .A2(n1192), .ZN(n1187) );
NOR2_X1 U860 ( .A1(n1178), .A2(n1193), .ZN(G60) );
XOR2_X1 U861 ( .A(n1194), .B(n1195), .Z(n1193) );
NAND3_X1 U862 ( .A1(n1191), .A2(G475), .A3(KEYINPUT20), .ZN(n1194) );
XOR2_X1 U863 ( .A(G104), .B(n1196), .Z(G6) );
NOR2_X1 U864 ( .A1(n1178), .A2(n1197), .ZN(G57) );
NOR2_X1 U865 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U866 ( .A(KEYINPUT21), .B(n1200), .Z(n1199) );
NOR2_X1 U867 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
XNOR2_X1 U868 ( .A(n1203), .B(n1204), .ZN(n1201) );
NOR2_X1 U869 ( .A1(n1205), .A2(n1206), .ZN(n1198) );
XNOR2_X1 U870 ( .A(n1207), .B(n1204), .ZN(n1206) );
XNOR2_X1 U871 ( .A(n1208), .B(n1209), .ZN(n1204) );
NOR2_X1 U872 ( .A1(KEYINPUT30), .A2(n1210), .ZN(n1209) );
NAND2_X1 U873 ( .A1(n1191), .A2(G472), .ZN(n1208) );
INV_X1 U874 ( .A(n1202), .ZN(n1205) );
XNOR2_X1 U875 ( .A(n1211), .B(n1212), .ZN(n1202) );
NOR2_X1 U876 ( .A1(KEYINPUT4), .A2(n1213), .ZN(n1212) );
XNOR2_X1 U877 ( .A(G101), .B(KEYINPUT23), .ZN(n1211) );
NOR2_X1 U878 ( .A1(n1214), .A2(n1215), .ZN(G54) );
XNOR2_X1 U879 ( .A(n1216), .B(n1217), .ZN(n1215) );
XOR2_X1 U880 ( .A(n1218), .B(n1219), .Z(n1217) );
AND2_X1 U881 ( .A1(G469), .A2(n1191), .ZN(n1219) );
INV_X1 U882 ( .A(n1220), .ZN(n1191) );
XOR2_X1 U883 ( .A(n1221), .B(KEYINPUT59), .Z(n1214) );
NAND2_X1 U884 ( .A1(n1222), .A2(G953), .ZN(n1221) );
XNOR2_X1 U885 ( .A(G952), .B(KEYINPUT16), .ZN(n1222) );
NOR2_X1 U886 ( .A1(n1178), .A2(n1223), .ZN(G51) );
XOR2_X1 U887 ( .A(n1224), .B(n1225), .Z(n1223) );
XOR2_X1 U888 ( .A(n1226), .B(n1227), .Z(n1225) );
NOR2_X1 U889 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
INV_X1 U890 ( .A(n1230), .ZN(n1228) );
NOR2_X1 U891 ( .A1(n1121), .A2(n1220), .ZN(n1226) );
NAND2_X1 U892 ( .A1(n1185), .A2(n1183), .ZN(n1220) );
NAND2_X1 U893 ( .A1(n1231), .A2(n1144), .ZN(n1183) );
INV_X1 U894 ( .A(n1073), .ZN(n1144) );
NAND4_X1 U895 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1073) );
AND4_X1 U896 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235) );
NOR2_X1 U897 ( .A1(n1240), .A2(n1241), .ZN(n1234) );
NOR2_X1 U898 ( .A1(KEYINPUT55), .A2(n1242), .ZN(n1241) );
NOR2_X1 U899 ( .A1(n1243), .A2(n1109), .ZN(n1240) );
NOR2_X1 U900 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
AND3_X1 U901 ( .A1(n1246), .A2(n1102), .A3(n1247), .ZN(n1245) );
NOR3_X1 U902 ( .A1(n1248), .A2(n1106), .A3(n1249), .ZN(n1244) );
INV_X1 U903 ( .A(KEYINPUT55), .ZN(n1248) );
NAND2_X1 U904 ( .A1(n1106), .A2(n1250), .ZN(n1232) );
XOR2_X1 U905 ( .A(KEYINPUT10), .B(n1251), .Z(n1250) );
NOR2_X1 U906 ( .A1(n1249), .A2(n1252), .ZN(n1251) );
XNOR2_X1 U907 ( .A(KEYINPUT2), .B(n1108), .ZN(n1252) );
INV_X1 U908 ( .A(n1253), .ZN(n1249) );
INV_X1 U909 ( .A(n1074), .ZN(n1231) );
NAND4_X1 U910 ( .A1(n1254), .A2(n1069), .A3(n1255), .A4(n1256), .ZN(n1074) );
NOR4_X1 U911 ( .A1(n1257), .A2(n1258), .A3(n1259), .A4(n1196), .ZN(n1256) );
AND3_X1 U912 ( .A1(n1088), .A2(n1260), .A3(n1261), .ZN(n1196) );
NOR2_X1 U913 ( .A1(n1262), .A2(n1263), .ZN(n1255) );
NOR3_X1 U914 ( .A1(n1084), .A2(n1264), .A3(n1109), .ZN(n1263) );
NAND3_X1 U915 ( .A1(n1260), .A2(n1265), .A3(n1088), .ZN(n1069) );
XNOR2_X1 U916 ( .A(G902), .B(KEYINPUT3), .ZN(n1185) );
NOR2_X1 U917 ( .A1(KEYINPUT38), .A2(n1266), .ZN(n1224) );
NOR2_X1 U918 ( .A1(n1076), .A2(G952), .ZN(n1178) );
XNOR2_X1 U919 ( .A(G146), .B(n1233), .ZN(G48) );
NAND4_X1 U920 ( .A1(n1246), .A2(n1247), .A3(n1261), .A4(n1102), .ZN(n1233) );
NAND2_X1 U921 ( .A1(n1267), .A2(n1268), .ZN(G45) );
NAND2_X1 U922 ( .A1(G143), .A2(n1238), .ZN(n1268) );
XOR2_X1 U923 ( .A(n1269), .B(KEYINPUT33), .Z(n1267) );
OR2_X1 U924 ( .A1(n1238), .A2(G143), .ZN(n1269) );
NAND4_X1 U925 ( .A1(n1270), .A2(n1253), .A3(n1102), .A4(n1271), .ZN(n1238) );
XNOR2_X1 U926 ( .A(G140), .B(n1237), .ZN(G42) );
NAND4_X1 U927 ( .A1(n1246), .A2(n1106), .A3(n1261), .A4(n1087), .ZN(n1237) );
XNOR2_X1 U928 ( .A(n1236), .B(n1272), .ZN(G39) );
NOR2_X1 U929 ( .A1(KEYINPUT41), .A2(n1273), .ZN(n1272) );
INV_X1 U930 ( .A(G137), .ZN(n1273) );
NAND3_X1 U931 ( .A1(n1082), .A2(n1247), .A3(n1246), .ZN(n1236) );
INV_X1 U932 ( .A(n1274), .ZN(n1246) );
AND2_X1 U933 ( .A1(n1106), .A2(n1101), .ZN(n1082) );
XNOR2_X1 U934 ( .A(n1242), .B(n1275), .ZN(G36) );
NOR2_X1 U935 ( .A1(KEYINPUT12), .A2(n1276), .ZN(n1275) );
NAND2_X1 U936 ( .A1(n1277), .A2(n1265), .ZN(n1242) );
XNOR2_X1 U937 ( .A(G131), .B(n1278), .ZN(G33) );
NAND2_X1 U938 ( .A1(n1277), .A2(n1261), .ZN(n1278) );
AND2_X1 U939 ( .A1(n1253), .A2(n1106), .ZN(n1277) );
NOR2_X1 U940 ( .A1(n1279), .A2(n1103), .ZN(n1106) );
NOR3_X1 U941 ( .A1(n1126), .A2(n1280), .A3(n1274), .ZN(n1253) );
NAND2_X1 U942 ( .A1(n1281), .A2(n1282), .ZN(n1274) );
XNOR2_X1 U943 ( .A(G128), .B(n1283), .ZN(G30) );
NAND4_X1 U944 ( .A1(n1284), .A2(n1282), .A3(n1102), .A4(n1285), .ZN(n1283) );
NOR2_X1 U945 ( .A1(n1109), .A2(n1286), .ZN(n1285) );
XNOR2_X1 U946 ( .A(KEYINPUT28), .B(n1093), .ZN(n1284) );
INV_X1 U947 ( .A(n1281), .ZN(n1093) );
XNOR2_X1 U948 ( .A(n1287), .B(n1259), .ZN(G3) );
NOR4_X1 U949 ( .A1(n1280), .A2(n1124), .A3(n1126), .A4(n1288), .ZN(n1259) );
XNOR2_X1 U950 ( .A(G125), .B(n1239), .ZN(G27) );
NAND3_X1 U951 ( .A1(n1261), .A2(n1086), .A3(n1289), .ZN(n1239) );
AND3_X1 U952 ( .A1(n1102), .A2(n1282), .A3(n1087), .ZN(n1289) );
NAND2_X1 U953 ( .A1(n1290), .A2(n1110), .ZN(n1282) );
NAND4_X1 U954 ( .A1(G953), .A2(G902), .A3(n1291), .A4(n1136), .ZN(n1290) );
INV_X1 U955 ( .A(G900), .ZN(n1136) );
INV_X1 U956 ( .A(n1108), .ZN(n1261) );
XOR2_X1 U957 ( .A(n1262), .B(n1292), .Z(G24) );
NOR2_X1 U958 ( .A1(KEYINPUT37), .A2(n1293), .ZN(n1292) );
AND4_X1 U959 ( .A1(n1294), .A2(n1271), .A3(n1088), .A4(n1295), .ZN(n1262) );
AND2_X1 U960 ( .A1(n1086), .A2(n1270), .ZN(n1295) );
XNOR2_X1 U961 ( .A(n1296), .B(KEYINPUT62), .ZN(n1270) );
XOR2_X1 U962 ( .A(n1254), .B(n1297), .Z(G21) );
NAND2_X1 U963 ( .A1(KEYINPUT18), .A2(G119), .ZN(n1297) );
NAND4_X1 U964 ( .A1(n1247), .A2(n1086), .A3(n1101), .A4(n1294), .ZN(n1254) );
INV_X1 U965 ( .A(n1298), .ZN(n1086) );
INV_X1 U966 ( .A(n1286), .ZN(n1247) );
NAND2_X1 U967 ( .A1(n1299), .A2(n1300), .ZN(n1286) );
XNOR2_X1 U968 ( .A(KEYINPUT27), .B(n1126), .ZN(n1299) );
XNOR2_X1 U969 ( .A(G116), .B(n1301), .ZN(G18) );
NAND4_X1 U970 ( .A1(n1302), .A2(n1265), .A3(n1303), .A4(n1304), .ZN(n1301) );
XOR2_X1 U971 ( .A(KEYINPUT22), .B(n1102), .Z(n1303) );
INV_X1 U972 ( .A(n1109), .ZN(n1265) );
NAND2_X1 U973 ( .A1(n1305), .A2(n1271), .ZN(n1109) );
XNOR2_X1 U974 ( .A(n1306), .B(KEYINPUT1), .ZN(n1271) );
XNOR2_X1 U975 ( .A(n1296), .B(KEYINPUT13), .ZN(n1305) );
XOR2_X1 U976 ( .A(G113), .B(n1258), .Z(G15) );
NOR3_X1 U977 ( .A1(n1084), .A2(n1264), .A3(n1108), .ZN(n1258) );
NAND2_X1 U978 ( .A1(n1306), .A2(n1296), .ZN(n1108) );
INV_X1 U979 ( .A(n1302), .ZN(n1084) );
NOR3_X1 U980 ( .A1(n1126), .A2(n1280), .A3(n1298), .ZN(n1302) );
NAND2_X1 U981 ( .A1(n1096), .A2(n1307), .ZN(n1298) );
XOR2_X1 U982 ( .A(G110), .B(n1257), .Z(G12) );
AND3_X1 U983 ( .A1(n1260), .A2(n1087), .A3(n1101), .ZN(n1257) );
INV_X1 U984 ( .A(n1124), .ZN(n1101) );
NAND2_X1 U985 ( .A1(n1308), .A2(n1306), .ZN(n1124) );
XOR2_X1 U986 ( .A(n1309), .B(G478), .Z(n1306) );
NAND2_X1 U987 ( .A1(n1192), .A2(n1310), .ZN(n1309) );
XOR2_X1 U988 ( .A(n1311), .B(n1312), .Z(n1192) );
NOR2_X1 U989 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U990 ( .A(n1315), .B(KEYINPUT25), .Z(n1314) );
NAND2_X1 U991 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
NOR2_X1 U992 ( .A1(n1317), .A2(n1316), .ZN(n1313) );
XOR2_X1 U993 ( .A(n1318), .B(n1319), .Z(n1316) );
AND2_X1 U994 ( .A1(KEYINPUT15), .A2(n1276), .ZN(n1318) );
XOR2_X1 U995 ( .A(G107), .B(n1320), .Z(n1317) );
XNOR2_X1 U996 ( .A(n1293), .B(G116), .ZN(n1320) );
NAND2_X1 U997 ( .A1(n1321), .A2(G217), .ZN(n1311) );
INV_X1 U998 ( .A(n1296), .ZN(n1308) );
XNOR2_X1 U999 ( .A(n1322), .B(G475), .ZN(n1296) );
NAND2_X1 U1000 ( .A1(n1195), .A2(n1310), .ZN(n1322) );
XOR2_X1 U1001 ( .A(n1323), .B(n1324), .Z(n1195) );
XOR2_X1 U1002 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1003 ( .A(n1327), .B(n1328), .Z(n1326) );
AND3_X1 U1004 ( .A1(G214), .A2(n1076), .A3(n1329), .ZN(n1328) );
NAND2_X1 U1005 ( .A1(n1330), .A2(KEYINPUT49), .ZN(n1327) );
XNOR2_X1 U1006 ( .A(G113), .B(n1331), .ZN(n1330) );
NOR2_X1 U1007 ( .A1(G122), .A2(KEYINPUT46), .ZN(n1331) );
NAND2_X1 U1008 ( .A1(n1332), .A2(KEYINPUT39), .ZN(n1325) );
XOR2_X1 U1009 ( .A(n1333), .B(n1334), .Z(n1332) );
XNOR2_X1 U1010 ( .A(n1335), .B(G125), .ZN(n1334) );
NAND2_X1 U1011 ( .A1(KEYINPUT6), .A2(G140), .ZN(n1333) );
XNOR2_X1 U1012 ( .A(G104), .B(n1336), .ZN(n1323) );
XOR2_X1 U1013 ( .A(G143), .B(G131), .Z(n1336) );
NAND2_X1 U1014 ( .A1(n1337), .A2(n1338), .ZN(n1087) );
NAND2_X1 U1015 ( .A1(n1088), .A2(n1339), .ZN(n1338) );
INV_X1 U1016 ( .A(KEYINPUT27), .ZN(n1339) );
NOR2_X1 U1017 ( .A1(n1126), .A2(n1300), .ZN(n1088) );
INV_X1 U1018 ( .A(n1280), .ZN(n1300) );
NAND3_X1 U1019 ( .A1(n1280), .A2(n1126), .A3(KEYINPUT27), .ZN(n1337) );
XNOR2_X1 U1020 ( .A(n1340), .B(n1182), .ZN(n1126) );
AND2_X1 U1021 ( .A1(G217), .A2(n1341), .ZN(n1182) );
NAND2_X1 U1022 ( .A1(n1181), .A2(n1310), .ZN(n1340) );
XOR2_X1 U1023 ( .A(n1342), .B(n1343), .Z(n1181) );
XOR2_X1 U1024 ( .A(n1344), .B(n1345), .Z(n1343) );
XNOR2_X1 U1025 ( .A(n1346), .B(n1347), .ZN(n1345) );
NOR2_X1 U1026 ( .A1(G128), .A2(KEYINPUT48), .ZN(n1347) );
NAND2_X1 U1027 ( .A1(KEYINPUT45), .A2(G125), .ZN(n1346) );
XOR2_X1 U1028 ( .A(n1348), .B(n1349), .Z(n1342) );
XNOR2_X1 U1029 ( .A(n1335), .B(G137), .ZN(n1349) );
INV_X1 U1030 ( .A(G146), .ZN(n1335) );
XOR2_X1 U1031 ( .A(n1350), .B(G119), .Z(n1348) );
NAND2_X1 U1032 ( .A1(G221), .A2(n1321), .ZN(n1350) );
AND2_X1 U1033 ( .A1(G234), .A2(n1076), .ZN(n1321) );
XOR2_X1 U1034 ( .A(n1351), .B(n1127), .Z(n1280) );
NAND2_X1 U1035 ( .A1(n1352), .A2(n1310), .ZN(n1127) );
XOR2_X1 U1036 ( .A(n1353), .B(n1354), .Z(n1352) );
XNOR2_X1 U1037 ( .A(n1287), .B(n1213), .ZN(n1354) );
NAND3_X1 U1038 ( .A1(n1329), .A2(n1076), .A3(G210), .ZN(n1213) );
INV_X1 U1039 ( .A(G101), .ZN(n1287) );
NAND2_X1 U1040 ( .A1(KEYINPUT8), .A2(n1355), .ZN(n1353) );
XNOR2_X1 U1041 ( .A(n1210), .B(n1207), .ZN(n1355) );
INV_X1 U1042 ( .A(n1203), .ZN(n1207) );
XNOR2_X1 U1043 ( .A(n1356), .B(n1357), .ZN(n1203) );
XNOR2_X1 U1044 ( .A(G113), .B(KEYINPUT35), .ZN(n1356) );
XNOR2_X1 U1045 ( .A(n1358), .B(n1359), .ZN(n1210) );
NAND2_X1 U1046 ( .A1(KEYINPUT0), .A2(n1129), .ZN(n1351) );
INV_X1 U1047 ( .A(G472), .ZN(n1129) );
INV_X1 U1048 ( .A(n1288), .ZN(n1260) );
NAND2_X1 U1049 ( .A1(n1281), .A2(n1294), .ZN(n1288) );
INV_X1 U1050 ( .A(n1264), .ZN(n1294) );
NAND2_X1 U1051 ( .A1(n1102), .A2(n1304), .ZN(n1264) );
NAND2_X1 U1052 ( .A1(n1110), .A2(n1360), .ZN(n1304) );
NAND3_X1 U1053 ( .A1(n1168), .A2(G902), .A3(n1361), .ZN(n1360) );
XOR2_X1 U1054 ( .A(n1291), .B(KEYINPUT24), .Z(n1361) );
NOR2_X1 U1055 ( .A1(n1076), .A2(G898), .ZN(n1168) );
NAND3_X1 U1056 ( .A1(n1291), .A2(n1076), .A3(G952), .ZN(n1110) );
NAND2_X1 U1057 ( .A1(G237), .A2(G234), .ZN(n1291) );
NOR2_X1 U1058 ( .A1(n1104), .A2(n1103), .ZN(n1102) );
AND2_X1 U1059 ( .A1(G214), .A2(n1362), .ZN(n1103) );
INV_X1 U1060 ( .A(n1279), .ZN(n1104) );
NAND3_X1 U1061 ( .A1(n1363), .A2(n1364), .A3(n1365), .ZN(n1279) );
NAND2_X1 U1062 ( .A1(n1120), .A2(n1366), .ZN(n1365) );
OR3_X1 U1063 ( .A1(n1366), .A2(n1120), .A3(n1121), .ZN(n1364) );
INV_X1 U1064 ( .A(KEYINPUT43), .ZN(n1366) );
NAND2_X1 U1065 ( .A1(n1367), .A2(n1121), .ZN(n1363) );
NAND2_X1 U1066 ( .A1(G210), .A2(n1362), .ZN(n1121) );
NAND2_X1 U1067 ( .A1(n1329), .A2(n1368), .ZN(n1362) );
INV_X1 U1068 ( .A(G237), .ZN(n1329) );
NAND2_X1 U1069 ( .A1(n1369), .A2(KEYINPUT43), .ZN(n1367) );
XNOR2_X1 U1070 ( .A(n1120), .B(KEYINPUT32), .ZN(n1369) );
AND2_X1 U1071 ( .A1(n1370), .A2(n1310), .ZN(n1120) );
XNOR2_X1 U1072 ( .A(n1371), .B(n1266), .ZN(n1370) );
AND2_X1 U1073 ( .A1(n1372), .A2(n1373), .ZN(n1266) );
NAND2_X1 U1074 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
NAND2_X1 U1075 ( .A1(n1376), .A2(n1176), .ZN(n1372) );
INV_X1 U1076 ( .A(n1375), .ZN(n1176) );
NAND2_X1 U1077 ( .A1(n1377), .A2(n1378), .ZN(n1375) );
OR2_X1 U1078 ( .A1(n1357), .A2(G113), .ZN(n1378) );
XOR2_X1 U1079 ( .A(n1379), .B(KEYINPUT50), .Z(n1377) );
NAND2_X1 U1080 ( .A1(G113), .A2(n1357), .ZN(n1379) );
XOR2_X1 U1081 ( .A(G116), .B(G119), .Z(n1357) );
XOR2_X1 U1082 ( .A(KEYINPUT57), .B(n1374), .Z(n1376) );
XOR2_X1 U1083 ( .A(n1177), .B(n1173), .Z(n1374) );
XNOR2_X1 U1084 ( .A(G110), .B(n1293), .ZN(n1173) );
INV_X1 U1085 ( .A(G122), .ZN(n1293) );
NAND3_X1 U1086 ( .A1(n1380), .A2(n1381), .A3(n1230), .ZN(n1371) );
NAND2_X1 U1087 ( .A1(n1382), .A2(n1383), .ZN(n1230) );
NAND2_X1 U1088 ( .A1(n1229), .A2(n1384), .ZN(n1381) );
INV_X1 U1089 ( .A(KEYINPUT36), .ZN(n1384) );
NOR2_X1 U1090 ( .A1(n1383), .A2(n1382), .ZN(n1229) );
XNOR2_X1 U1091 ( .A(n1385), .B(n1155), .ZN(n1383) );
INV_X1 U1092 ( .A(G125), .ZN(n1155) );
NAND2_X1 U1093 ( .A1(KEYINPUT36), .A2(n1382), .ZN(n1380) );
NOR2_X1 U1094 ( .A1(n1163), .A2(G953), .ZN(n1382) );
INV_X1 U1095 ( .A(G224), .ZN(n1163) );
NOR2_X1 U1096 ( .A1(n1096), .A2(n1095), .ZN(n1281) );
INV_X1 U1097 ( .A(n1307), .ZN(n1095) );
NAND2_X1 U1098 ( .A1(G221), .A2(n1341), .ZN(n1307) );
NAND2_X1 U1099 ( .A1(G234), .A2(n1368), .ZN(n1341) );
XNOR2_X1 U1100 ( .A(n1131), .B(n1386), .ZN(n1096) );
NOR2_X1 U1101 ( .A1(G469), .A2(KEYINPUT14), .ZN(n1386) );
NAND2_X1 U1102 ( .A1(n1387), .A2(n1310), .ZN(n1131) );
XNOR2_X1 U1103 ( .A(n1368), .B(KEYINPUT7), .ZN(n1310) );
INV_X1 U1104 ( .A(G902), .ZN(n1368) );
XOR2_X1 U1105 ( .A(n1388), .B(n1389), .Z(n1387) );
NOR2_X1 U1106 ( .A1(KEYINPUT17), .A2(n1216), .ZN(n1389) );
AND2_X1 U1107 ( .A1(n1390), .A2(n1391), .ZN(n1216) );
NAND2_X1 U1108 ( .A1(n1344), .A2(n1392), .ZN(n1391) );
NAND2_X1 U1109 ( .A1(G227), .A2(n1076), .ZN(n1392) );
INV_X1 U1110 ( .A(G953), .ZN(n1076) );
OR3_X1 U1111 ( .A1(n1135), .A2(G953), .A3(n1344), .ZN(n1390) );
XOR2_X1 U1112 ( .A(G110), .B(G140), .Z(n1344) );
INV_X1 U1113 ( .A(G227), .ZN(n1135) );
NAND2_X1 U1114 ( .A1(n1393), .A2(n1394), .ZN(n1388) );
OR2_X1 U1115 ( .A1(n1218), .A2(KEYINPUT52), .ZN(n1394) );
XNOR2_X1 U1116 ( .A(n1395), .B(n1358), .ZN(n1218) );
NAND3_X1 U1117 ( .A1(n1395), .A2(n1358), .A3(KEYINPUT52), .ZN(n1393) );
XNOR2_X1 U1118 ( .A(G131), .B(n1158), .ZN(n1358) );
XNOR2_X1 U1119 ( .A(n1276), .B(G137), .ZN(n1158) );
INV_X1 U1120 ( .A(G134), .ZN(n1276) );
XOR2_X1 U1121 ( .A(n1396), .B(n1148), .Z(n1395) );
XNOR2_X1 U1122 ( .A(n1385), .B(n1397), .ZN(n1148) );
XOR2_X1 U1123 ( .A(KEYINPUT51), .B(KEYINPUT34), .Z(n1397) );
INV_X1 U1124 ( .A(n1359), .ZN(n1385) );
XOR2_X1 U1125 ( .A(G146), .B(n1319), .Z(n1359) );
XOR2_X1 U1126 ( .A(G128), .B(G143), .Z(n1319) );
XNOR2_X1 U1127 ( .A(n1177), .B(KEYINPUT19), .ZN(n1396) );
XOR2_X1 U1128 ( .A(G101), .B(n1398), .Z(n1177) );
XOR2_X1 U1129 ( .A(G107), .B(G104), .Z(n1398) );
endmodule


