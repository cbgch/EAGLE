//Key = 0011101110110010111000110001111001110000100110011001010000010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374;

XOR2_X1 U750 ( .A(G107), .B(n1040), .Z(G9) );
NOR2_X1 U751 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR3_X1 U752 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
INV_X1 U753 ( .A(n1046), .ZN(n1045) );
INV_X1 U754 ( .A(G952), .ZN(n1044) );
NAND3_X1 U755 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1043) );
NAND2_X1 U756 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U757 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND3_X1 U758 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NAND2_X1 U759 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
OR3_X1 U760 ( .A1(n1059), .A2(KEYINPUT2), .A3(n1060), .ZN(n1057) );
NAND3_X1 U761 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1054) );
NAND2_X1 U762 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND2_X1 U763 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1061) );
NAND2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U766 ( .A1(KEYINPUT2), .A2(n1072), .ZN(n1071) );
NAND3_X1 U767 ( .A1(n1064), .A2(n1073), .A3(n1068), .ZN(n1052) );
NAND3_X1 U768 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
NAND2_X1 U769 ( .A1(n1056), .A2(n1077), .ZN(n1076) );
NAND3_X1 U770 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1075) );
XNOR2_X1 U771 ( .A(KEYINPUT41), .B(n1081), .ZN(n1079) );
NAND2_X1 U772 ( .A1(n1063), .A2(n1082), .ZN(n1074) );
NAND2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U774 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
INV_X1 U775 ( .A(n1087), .ZN(n1050) );
NOR3_X1 U776 ( .A1(n1088), .A2(G953), .A3(n1089), .ZN(n1041) );
INV_X1 U777 ( .A(n1047), .ZN(n1089) );
NAND4_X1 U778 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1047) );
NOR4_X1 U779 ( .A1(n1094), .A2(n1095), .A3(n1058), .A4(n1096), .ZN(n1093) );
XNOR2_X1 U780 ( .A(n1097), .B(KEYINPUT11), .ZN(n1094) );
NOR3_X1 U781 ( .A1(n1085), .A2(n1098), .A3(n1099), .ZN(n1092) );
INV_X1 U782 ( .A(n1100), .ZN(n1099) );
NAND2_X1 U783 ( .A1(n1101), .A2(n1102), .ZN(n1091) );
NAND2_X1 U784 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NAND2_X1 U785 ( .A1(KEYINPUT38), .A2(KEYINPUT14), .ZN(n1104) );
NAND3_X1 U786 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1090) );
INV_X1 U787 ( .A(KEYINPUT38), .ZN(n1107) );
NAND2_X1 U788 ( .A1(KEYINPUT14), .A2(n1108), .ZN(n1106) );
NAND2_X1 U789 ( .A1(n1103), .A2(G475), .ZN(n1108) );
NAND2_X1 U790 ( .A1(n1103), .A2(n1109), .ZN(n1105) );
INV_X1 U791 ( .A(KEYINPUT14), .ZN(n1109) );
XNOR2_X1 U792 ( .A(n1110), .B(KEYINPUT1), .ZN(n1103) );
XNOR2_X1 U793 ( .A(G952), .B(KEYINPUT27), .ZN(n1088) );
XOR2_X1 U794 ( .A(n1111), .B(n1112), .Z(G72) );
XOR2_X1 U795 ( .A(n1113), .B(n1114), .Z(n1112) );
NAND2_X1 U796 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XNOR2_X1 U797 ( .A(n1117), .B(n1118), .ZN(n1115) );
NAND2_X1 U798 ( .A1(G953), .A2(n1119), .ZN(n1113) );
NAND2_X1 U799 ( .A1(G900), .A2(n1120), .ZN(n1119) );
XOR2_X1 U800 ( .A(KEYINPUT50), .B(G227), .Z(n1120) );
NOR2_X1 U801 ( .A1(G953), .A2(n1121), .ZN(n1111) );
NOR2_X1 U802 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XNOR2_X1 U803 ( .A(n1124), .B(KEYINPUT7), .ZN(n1122) );
NAND2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(G69) );
NAND2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U806 ( .A(KEYINPUT62), .B(n1129), .Z(n1125) );
NOR2_X1 U807 ( .A1(n1127), .A2(n1130), .ZN(n1129) );
NOR2_X1 U808 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
INV_X1 U809 ( .A(n1128), .ZN(n1132) );
NAND3_X1 U810 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1128) );
NAND2_X1 U811 ( .A1(n1136), .A2(n1048), .ZN(n1134) );
NAND2_X1 U812 ( .A1(n1137), .A2(G953), .ZN(n1133) );
XNOR2_X1 U813 ( .A(G898), .B(KEYINPUT60), .ZN(n1137) );
NOR2_X1 U814 ( .A1(n1138), .A2(n1135), .ZN(n1131) );
XNOR2_X1 U815 ( .A(n1139), .B(n1140), .ZN(n1135) );
XOR2_X1 U816 ( .A(G110), .B(n1141), .Z(n1140) );
NOR2_X1 U817 ( .A1(KEYINPUT24), .A2(n1142), .ZN(n1141) );
XNOR2_X1 U818 ( .A(G119), .B(n1143), .ZN(n1142) );
INV_X1 U819 ( .A(n1136), .ZN(n1138) );
AND2_X1 U820 ( .A1(G953), .A2(n1144), .ZN(n1127) );
NAND2_X1 U821 ( .A1(G898), .A2(G224), .ZN(n1144) );
NOR2_X1 U822 ( .A1(n1145), .A2(n1146), .ZN(G66) );
XOR2_X1 U823 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U824 ( .A(n1149), .B(n1150), .Z(n1148) );
NAND3_X1 U825 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1149) );
OR2_X1 U826 ( .A1(n1154), .A2(KEYINPUT46), .ZN(n1152) );
NAND2_X1 U827 ( .A1(KEYINPUT46), .A2(n1155), .ZN(n1151) );
NAND2_X1 U828 ( .A1(n1046), .A2(G902), .ZN(n1155) );
XOR2_X1 U829 ( .A(KEYINPUT53), .B(KEYINPUT23), .Z(n1147) );
NOR2_X1 U830 ( .A1(n1145), .A2(n1156), .ZN(G63) );
XOR2_X1 U831 ( .A(n1157), .B(n1158), .Z(n1156) );
AND2_X1 U832 ( .A1(G478), .A2(n1154), .ZN(n1157) );
NOR2_X1 U833 ( .A1(n1145), .A2(n1159), .ZN(G60) );
NOR3_X1 U834 ( .A1(n1110), .A2(n1160), .A3(n1161), .ZN(n1159) );
AND3_X1 U835 ( .A1(n1162), .A2(G475), .A3(n1154), .ZN(n1161) );
NOR2_X1 U836 ( .A1(n1163), .A2(n1162), .ZN(n1160) );
NOR2_X1 U837 ( .A1(n1046), .A2(n1102), .ZN(n1163) );
XNOR2_X1 U838 ( .A(G104), .B(n1164), .ZN(G6) );
NOR2_X1 U839 ( .A1(n1145), .A2(n1165), .ZN(G57) );
XOR2_X1 U840 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U841 ( .A1(KEYINPUT19), .A2(n1168), .ZN(n1167) );
XOR2_X1 U842 ( .A(n1169), .B(n1170), .Z(n1166) );
NOR3_X1 U843 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1170) );
NOR2_X1 U844 ( .A1(KEYINPUT56), .A2(n1174), .ZN(n1173) );
NOR2_X1 U845 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
AND2_X1 U846 ( .A1(n1177), .A2(KEYINPUT39), .ZN(n1176) );
NOR3_X1 U847 ( .A1(KEYINPUT39), .A2(n1178), .A3(n1177), .ZN(n1175) );
NOR2_X1 U848 ( .A1(n1179), .A2(n1180), .ZN(n1172) );
INV_X1 U849 ( .A(KEYINPUT56), .ZN(n1180) );
NOR2_X1 U850 ( .A1(n1178), .A2(n1181), .ZN(n1179) );
XOR2_X1 U851 ( .A(KEYINPUT39), .B(n1177), .Z(n1181) );
AND2_X1 U852 ( .A1(n1178), .A2(n1177), .ZN(n1171) );
NAND2_X1 U853 ( .A1(n1154), .A2(G472), .ZN(n1169) );
NOR2_X1 U854 ( .A1(n1145), .A2(n1182), .ZN(G54) );
XOR2_X1 U855 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U856 ( .A(n1185), .B(n1186), .Z(n1184) );
XNOR2_X1 U857 ( .A(n1187), .B(n1188), .ZN(n1186) );
NOR2_X1 U858 ( .A1(KEYINPUT49), .A2(G110), .ZN(n1185) );
XOR2_X1 U859 ( .A(n1189), .B(n1190), .Z(n1183) );
NOR2_X1 U860 ( .A1(KEYINPUT25), .A2(n1191), .ZN(n1190) );
NAND2_X1 U861 ( .A1(n1154), .A2(G469), .ZN(n1189) );
NOR2_X1 U862 ( .A1(n1145), .A2(n1192), .ZN(G51) );
XNOR2_X1 U863 ( .A(n1193), .B(n1194), .ZN(n1192) );
XOR2_X1 U864 ( .A(n1195), .B(n1196), .Z(n1194) );
NOR2_X1 U865 ( .A1(n1197), .A2(n1198), .ZN(n1195) );
INV_X1 U866 ( .A(n1154), .ZN(n1198) );
NOR2_X1 U867 ( .A1(n1199), .A2(n1046), .ZN(n1154) );
NOR3_X1 U868 ( .A1(n1123), .A2(n1124), .A3(n1136), .ZN(n1046) );
NAND4_X1 U869 ( .A1(n1164), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1136) );
NOR4_X1 U870 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1040), .ZN(n1202) );
AND4_X1 U871 ( .A1(n1077), .A2(n1206), .A3(n1064), .A4(n1207), .ZN(n1040) );
NAND2_X1 U872 ( .A1(n1208), .A2(n1209), .ZN(n1201) );
NAND2_X1 U873 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND2_X1 U874 ( .A1(n1212), .A2(n1063), .ZN(n1211) );
NAND2_X1 U875 ( .A1(n1068), .A2(n1077), .ZN(n1210) );
INV_X1 U876 ( .A(n1213), .ZN(n1208) );
NAND4_X1 U877 ( .A1(n1212), .A2(n1077), .A3(n1206), .A4(n1064), .ZN(n1164) );
AND4_X1 U878 ( .A1(n1214), .A2(n1215), .A3(n1072), .A4(n1216), .ZN(n1124) );
NOR2_X1 U879 ( .A1(n1067), .A2(n1081), .ZN(n1216) );
NAND2_X1 U880 ( .A1(KEYINPUT6), .A2(n1217), .ZN(n1215) );
NAND2_X1 U881 ( .A1(n1218), .A2(n1219), .ZN(n1214) );
INV_X1 U882 ( .A(KEYINPUT6), .ZN(n1219) );
NAND2_X1 U883 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
NAND4_X1 U884 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1123) );
AND2_X1 U885 ( .A1(n1226), .A2(n1227), .ZN(n1224) );
NAND2_X1 U886 ( .A1(n1228), .A2(n1229), .ZN(n1222) );
NAND2_X1 U887 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND2_X1 U888 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
XNOR2_X1 U889 ( .A(n1234), .B(KEYINPUT43), .ZN(n1232) );
NAND2_X1 U890 ( .A1(n1056), .A2(n1235), .ZN(n1230) );
NAND2_X1 U891 ( .A1(n1236), .A2(n1059), .ZN(n1235) );
XNOR2_X1 U892 ( .A(KEYINPUT34), .B(n1070), .ZN(n1236) );
NOR2_X1 U893 ( .A1(n1048), .A2(G952), .ZN(n1145) );
XOR2_X1 U894 ( .A(G146), .B(n1237), .Z(G48) );
NOR3_X1 U895 ( .A1(n1238), .A2(n1083), .A3(n1239), .ZN(n1237) );
XNOR2_X1 U896 ( .A(G143), .B(n1223), .ZN(G45) );
NAND3_X1 U897 ( .A1(n1240), .A2(n1072), .A3(n1241), .ZN(n1223) );
NOR3_X1 U898 ( .A1(n1083), .A2(n1242), .A3(n1243), .ZN(n1241) );
XNOR2_X1 U899 ( .A(G140), .B(n1244), .ZN(G42) );
NAND2_X1 U900 ( .A1(n1056), .A2(n1245), .ZN(n1244) );
XOR2_X1 U901 ( .A(KEYINPUT54), .B(n1246), .Z(n1245) );
NOR2_X1 U902 ( .A1(n1070), .A2(n1238), .ZN(n1246) );
INV_X1 U903 ( .A(n1228), .ZN(n1238) );
INV_X1 U904 ( .A(n1247), .ZN(n1070) );
XNOR2_X1 U905 ( .A(G137), .B(n1225), .ZN(G39) );
NAND4_X1 U906 ( .A1(n1240), .A2(n1234), .A3(n1068), .A4(n1056), .ZN(n1225) );
INV_X1 U907 ( .A(n1217), .ZN(n1240) );
XOR2_X1 U908 ( .A(n1248), .B(n1249), .Z(G36) );
XOR2_X1 U909 ( .A(KEYINPUT16), .B(G134), .Z(n1249) );
NOR2_X1 U910 ( .A1(KEYINPUT37), .A2(n1250), .ZN(n1248) );
NOR4_X1 U911 ( .A1(n1067), .A2(n1081), .A3(n1059), .A4(n1217), .ZN(n1250) );
XNOR2_X1 U912 ( .A(G131), .B(n1251), .ZN(G33) );
NAND3_X1 U913 ( .A1(n1056), .A2(n1252), .A3(n1228), .ZN(n1251) );
NOR2_X1 U914 ( .A1(n1217), .A2(n1066), .ZN(n1228) );
XNOR2_X1 U915 ( .A(KEYINPUT15), .B(n1059), .ZN(n1252) );
INV_X1 U916 ( .A(n1081), .ZN(n1056) );
NAND2_X1 U917 ( .A1(n1253), .A2(n1254), .ZN(n1081) );
XNOR2_X1 U918 ( .A(n1095), .B(KEYINPUT5), .ZN(n1253) );
NAND2_X1 U919 ( .A1(n1255), .A2(n1256), .ZN(G30) );
NAND2_X1 U920 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND2_X1 U921 ( .A1(n1259), .A2(G128), .ZN(n1255) );
NAND2_X1 U922 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND2_X1 U923 ( .A1(KEYINPUT31), .A2(n1262), .ZN(n1261) );
OR2_X1 U924 ( .A1(n1257), .A2(KEYINPUT31), .ZN(n1260) );
NOR2_X1 U925 ( .A1(KEYINPUT12), .A2(n1226), .ZN(n1257) );
INV_X1 U926 ( .A(n1262), .ZN(n1226) );
NOR4_X1 U927 ( .A1(n1217), .A2(n1239), .A3(n1067), .A4(n1083), .ZN(n1262) );
INV_X1 U928 ( .A(n1233), .ZN(n1083) );
NAND2_X1 U929 ( .A1(n1077), .A2(n1220), .ZN(n1217) );
XNOR2_X1 U930 ( .A(n1263), .B(n1264), .ZN(G3) );
NOR4_X1 U931 ( .A1(KEYINPUT57), .A2(n1060), .A3(n1213), .A4(n1265), .ZN(n1264) );
XNOR2_X1 U932 ( .A(KEYINPUT35), .B(n1221), .ZN(n1265) );
INV_X1 U933 ( .A(n1077), .ZN(n1221) );
INV_X1 U934 ( .A(n1068), .ZN(n1060) );
XNOR2_X1 U935 ( .A(G125), .B(n1227), .ZN(G27) );
NAND3_X1 U936 ( .A1(n1212), .A2(n1247), .A3(n1266), .ZN(n1227) );
AND3_X1 U937 ( .A1(n1063), .A2(n1220), .A3(n1233), .ZN(n1266) );
NAND2_X1 U938 ( .A1(n1087), .A2(n1267), .ZN(n1220) );
NAND3_X1 U939 ( .A1(G902), .A2(n1268), .A3(n1269), .ZN(n1267) );
INV_X1 U940 ( .A(n1116), .ZN(n1269) );
NAND2_X1 U941 ( .A1(G953), .A2(n1270), .ZN(n1116) );
XOR2_X1 U942 ( .A(KEYINPUT47), .B(G900), .Z(n1270) );
XNOR2_X1 U943 ( .A(G122), .B(n1200), .ZN(G24) );
NAND4_X1 U944 ( .A1(n1063), .A2(n1206), .A3(n1271), .A4(n1064), .ZN(n1200) );
NOR2_X1 U945 ( .A1(n1272), .A2(n1097), .ZN(n1064) );
NOR2_X1 U946 ( .A1(n1242), .A2(n1243), .ZN(n1271) );
XOR2_X1 U947 ( .A(G119), .B(n1205), .Z(G21) );
AND4_X1 U948 ( .A1(n1234), .A2(n1068), .A3(n1063), .A4(n1206), .ZN(n1205) );
INV_X1 U949 ( .A(n1058), .ZN(n1063) );
INV_X1 U950 ( .A(n1239), .ZN(n1234) );
NAND2_X1 U951 ( .A1(n1097), .A2(n1272), .ZN(n1239) );
XNOR2_X1 U952 ( .A(G116), .B(n1273), .ZN(G18) );
NAND2_X1 U953 ( .A1(KEYINPUT29), .A2(n1204), .ZN(n1273) );
NOR3_X1 U954 ( .A1(n1058), .A2(n1067), .A3(n1213), .ZN(n1204) );
INV_X1 U955 ( .A(n1207), .ZN(n1067) );
NOR2_X1 U956 ( .A1(n1274), .A2(n1243), .ZN(n1207) );
INV_X1 U957 ( .A(n1096), .ZN(n1243) );
XNOR2_X1 U958 ( .A(n1275), .B(n1276), .ZN(G15) );
NOR4_X1 U959 ( .A1(KEYINPUT0), .A2(n1058), .A3(n1213), .A4(n1066), .ZN(n1276) );
INV_X1 U960 ( .A(n1212), .ZN(n1066) );
NOR2_X1 U961 ( .A1(n1096), .A2(n1242), .ZN(n1212) );
NAND2_X1 U962 ( .A1(n1072), .A2(n1206), .ZN(n1213) );
INV_X1 U963 ( .A(n1059), .ZN(n1072) );
NAND2_X1 U964 ( .A1(n1277), .A2(n1097), .ZN(n1059) );
NAND2_X1 U965 ( .A1(n1078), .A2(n1278), .ZN(n1058) );
XNOR2_X1 U966 ( .A(G110), .B(n1279), .ZN(G12) );
NAND2_X1 U967 ( .A1(KEYINPUT59), .A2(n1203), .ZN(n1279) );
AND4_X1 U968 ( .A1(n1068), .A2(n1247), .A3(n1077), .A4(n1206), .ZN(n1203) );
AND2_X1 U969 ( .A1(n1233), .A2(n1280), .ZN(n1206) );
NAND2_X1 U970 ( .A1(n1087), .A2(n1281), .ZN(n1280) );
NAND4_X1 U971 ( .A1(G953), .A2(G902), .A3(n1268), .A4(n1282), .ZN(n1281) );
INV_X1 U972 ( .A(G898), .ZN(n1282) );
NAND3_X1 U973 ( .A1(n1268), .A2(n1048), .A3(G952), .ZN(n1087) );
NAND2_X1 U974 ( .A1(G237), .A2(G234), .ZN(n1268) );
NOR2_X1 U975 ( .A1(n1086), .A2(n1085), .ZN(n1233) );
INV_X1 U976 ( .A(n1254), .ZN(n1085) );
NAND2_X1 U977 ( .A1(G214), .A2(n1283), .ZN(n1254) );
INV_X1 U978 ( .A(n1095), .ZN(n1086) );
XOR2_X1 U979 ( .A(n1284), .B(n1197), .Z(n1095) );
NAND2_X1 U980 ( .A1(G210), .A2(n1283), .ZN(n1197) );
NAND2_X1 U981 ( .A1(n1285), .A2(n1199), .ZN(n1283) );
XOR2_X1 U982 ( .A(KEYINPUT44), .B(G237), .Z(n1285) );
NAND2_X1 U983 ( .A1(n1286), .A2(n1199), .ZN(n1284) );
XNOR2_X1 U984 ( .A(n1196), .B(n1287), .ZN(n1286) );
NOR2_X1 U985 ( .A1(KEYINPUT13), .A2(n1193), .ZN(n1287) );
XOR2_X1 U986 ( .A(n1288), .B(n1289), .Z(n1193) );
XNOR2_X1 U987 ( .A(G125), .B(n1290), .ZN(n1289) );
XOR2_X1 U988 ( .A(n1291), .B(n1292), .Z(n1288) );
NAND2_X1 U989 ( .A1(G224), .A2(n1048), .ZN(n1291) );
XNOR2_X1 U990 ( .A(n1143), .B(n1293), .ZN(n1196) );
XNOR2_X1 U991 ( .A(n1294), .B(n1139), .ZN(n1293) );
XOR2_X1 U992 ( .A(n1295), .B(n1296), .Z(n1139) );
NOR2_X1 U993 ( .A1(KEYINPUT52), .A2(n1297), .ZN(n1296) );
XNOR2_X1 U994 ( .A(G104), .B(n1298), .ZN(n1297) );
XOR2_X1 U995 ( .A(KEYINPUT26), .B(G107), .Z(n1298) );
XNOR2_X1 U996 ( .A(G101), .B(G122), .ZN(n1295) );
XOR2_X1 U997 ( .A(n1299), .B(n1300), .Z(n1143) );
XNOR2_X1 U998 ( .A(n1301), .B(G113), .ZN(n1300) );
XNOR2_X1 U999 ( .A(KEYINPUT8), .B(KEYINPUT63), .ZN(n1299) );
NOR2_X1 U1000 ( .A1(n1078), .A2(n1080), .ZN(n1077) );
INV_X1 U1001 ( .A(n1278), .ZN(n1080) );
NAND2_X1 U1002 ( .A1(G221), .A2(n1302), .ZN(n1278) );
XOR2_X1 U1003 ( .A(n1303), .B(G469), .Z(n1078) );
NAND3_X1 U1004 ( .A1(n1304), .A2(n1305), .A3(n1199), .ZN(n1303) );
NAND3_X1 U1005 ( .A1(n1306), .A2(n1191), .A3(n1307), .ZN(n1305) );
INV_X1 U1006 ( .A(KEYINPUT18), .ZN(n1307) );
NAND2_X1 U1007 ( .A1(n1308), .A2(KEYINPUT18), .ZN(n1304) );
XNOR2_X1 U1008 ( .A(n1309), .B(n1191), .ZN(n1308) );
XOR2_X1 U1009 ( .A(n1118), .B(n1310), .Z(n1191) );
NOR2_X1 U1010 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U1011 ( .A(KEYINPUT45), .B(n1313), .Z(n1312) );
NOR2_X1 U1012 ( .A1(n1314), .A2(n1263), .ZN(n1313) );
AND2_X1 U1013 ( .A1(n1263), .A2(n1314), .ZN(n1311) );
NAND3_X1 U1014 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n1314) );
NAND2_X1 U1015 ( .A1(KEYINPUT58), .A2(G104), .ZN(n1317) );
OR3_X1 U1016 ( .A1(n1318), .A2(KEYINPUT58), .A3(G107), .ZN(n1316) );
NAND2_X1 U1017 ( .A1(G107), .A2(n1318), .ZN(n1315) );
NAND2_X1 U1018 ( .A1(KEYINPUT17), .A2(n1319), .ZN(n1318) );
INV_X1 U1019 ( .A(G101), .ZN(n1263) );
XNOR2_X1 U1020 ( .A(n1320), .B(n1258), .ZN(n1118) );
NOR2_X1 U1021 ( .A1(KEYINPUT36), .A2(n1306), .ZN(n1309) );
XOR2_X1 U1022 ( .A(n1321), .B(n1322), .Z(n1306) );
XOR2_X1 U1023 ( .A(KEYINPUT30), .B(G110), .Z(n1322) );
XOR2_X1 U1024 ( .A(n1323), .B(n1188), .Z(n1321) );
AND2_X1 U1025 ( .A1(G227), .A2(n1048), .ZN(n1188) );
NAND2_X1 U1026 ( .A1(KEYINPUT33), .A2(n1187), .ZN(n1323) );
NOR2_X1 U1027 ( .A1(n1097), .A2(n1277), .ZN(n1247) );
INV_X1 U1028 ( .A(n1272), .ZN(n1277) );
NAND2_X1 U1029 ( .A1(n1324), .A2(n1100), .ZN(n1272) );
NAND3_X1 U1030 ( .A1(n1325), .A2(n1199), .A3(n1150), .ZN(n1100) );
XOR2_X1 U1031 ( .A(KEYINPUT48), .B(n1098), .Z(n1324) );
AND2_X1 U1032 ( .A1(n1153), .A2(n1326), .ZN(n1098) );
NAND2_X1 U1033 ( .A1(n1150), .A2(n1199), .ZN(n1326) );
XOR2_X1 U1034 ( .A(n1327), .B(n1328), .Z(n1150) );
XOR2_X1 U1035 ( .A(n1294), .B(n1117), .Z(n1328) );
XNOR2_X1 U1036 ( .A(G125), .B(n1187), .ZN(n1117) );
XOR2_X1 U1037 ( .A(G110), .B(G119), .Z(n1294) );
XOR2_X1 U1038 ( .A(n1329), .B(n1330), .Z(n1327) );
NOR2_X1 U1039 ( .A1(G128), .A2(KEYINPUT55), .ZN(n1330) );
XOR2_X1 U1040 ( .A(n1331), .B(G146), .Z(n1329) );
NAND3_X1 U1041 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1331) );
NAND2_X1 U1042 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
OR3_X1 U1043 ( .A1(n1336), .A2(n1335), .A3(n1337), .ZN(n1333) );
INV_X1 U1044 ( .A(KEYINPUT3), .ZN(n1336) );
NAND2_X1 U1045 ( .A1(n1338), .A2(n1337), .ZN(n1332) );
INV_X1 U1046 ( .A(G137), .ZN(n1337) );
NAND2_X1 U1047 ( .A1(KEYINPUT3), .A2(n1339), .ZN(n1338) );
XNOR2_X1 U1048 ( .A(KEYINPUT9), .B(n1335), .ZN(n1339) );
NAND2_X1 U1049 ( .A1(n1340), .A2(G221), .ZN(n1335) );
INV_X1 U1050 ( .A(n1325), .ZN(n1153) );
NAND2_X1 U1051 ( .A1(G217), .A2(n1302), .ZN(n1325) );
NAND2_X1 U1052 ( .A1(G234), .A2(n1199), .ZN(n1302) );
XNOR2_X1 U1053 ( .A(n1341), .B(G472), .ZN(n1097) );
NAND2_X1 U1054 ( .A1(n1342), .A2(n1199), .ZN(n1341) );
INV_X1 U1055 ( .A(G902), .ZN(n1199) );
XNOR2_X1 U1056 ( .A(n1168), .B(n1343), .ZN(n1342) );
XOR2_X1 U1057 ( .A(n1178), .B(n1177), .Z(n1343) );
XNOR2_X1 U1058 ( .A(n1275), .B(n1344), .ZN(n1177) );
NOR2_X1 U1059 ( .A1(KEYINPUT32), .A2(n1345), .ZN(n1344) );
XNOR2_X1 U1060 ( .A(G116), .B(G119), .ZN(n1345) );
XOR2_X1 U1061 ( .A(n1320), .B(n1290), .Z(n1178) );
NAND2_X1 U1062 ( .A1(KEYINPUT22), .A2(n1258), .ZN(n1290) );
INV_X1 U1063 ( .A(G128), .ZN(n1258) );
XOR2_X1 U1064 ( .A(n1346), .B(n1347), .Z(n1320) );
XNOR2_X1 U1065 ( .A(n1348), .B(n1292), .ZN(n1347) );
XOR2_X1 U1066 ( .A(G143), .B(G146), .Z(n1292) );
INV_X1 U1067 ( .A(n1349), .ZN(n1348) );
XNOR2_X1 U1068 ( .A(G134), .B(G137), .ZN(n1346) );
XOR2_X1 U1069 ( .A(n1350), .B(G101), .Z(n1168) );
NAND2_X1 U1070 ( .A1(n1351), .A2(G210), .ZN(n1350) );
NOR2_X1 U1071 ( .A1(n1096), .A2(n1274), .ZN(n1068) );
INV_X1 U1072 ( .A(n1242), .ZN(n1274) );
XOR2_X1 U1073 ( .A(n1110), .B(n1102), .Z(n1242) );
INV_X1 U1074 ( .A(G475), .ZN(n1102) );
NOR2_X1 U1075 ( .A1(n1162), .A2(G902), .ZN(n1110) );
XOR2_X1 U1076 ( .A(n1352), .B(n1353), .Z(n1162) );
XNOR2_X1 U1077 ( .A(n1319), .B(n1354), .ZN(n1353) );
XNOR2_X1 U1078 ( .A(KEYINPUT42), .B(n1187), .ZN(n1354) );
INV_X1 U1079 ( .A(G140), .ZN(n1187) );
INV_X1 U1080 ( .A(G104), .ZN(n1319) );
XOR2_X1 U1081 ( .A(n1355), .B(n1356), .Z(n1352) );
NOR2_X1 U1082 ( .A1(KEYINPUT21), .A2(n1357), .ZN(n1356) );
XNOR2_X1 U1083 ( .A(G143), .B(n1358), .ZN(n1357) );
NAND2_X1 U1084 ( .A1(n1351), .A2(G214), .ZN(n1358) );
NOR2_X1 U1085 ( .A1(G953), .A2(G237), .ZN(n1351) );
XOR2_X1 U1086 ( .A(n1359), .B(n1360), .Z(n1355) );
XOR2_X1 U1087 ( .A(n1361), .B(n1362), .Z(n1360) );
XOR2_X1 U1088 ( .A(G146), .B(G122), .Z(n1362) );
XOR2_X1 U1089 ( .A(KEYINPUT40), .B(KEYINPUT10), .Z(n1361) );
XNOR2_X1 U1090 ( .A(n1349), .B(n1363), .ZN(n1359) );
XNOR2_X1 U1091 ( .A(n1364), .B(n1365), .ZN(n1363) );
NOR2_X1 U1092 ( .A1(G125), .A2(KEYINPUT20), .ZN(n1365) );
NAND2_X1 U1093 ( .A1(KEYINPUT4), .A2(n1275), .ZN(n1364) );
INV_X1 U1094 ( .A(G113), .ZN(n1275) );
XOR2_X1 U1095 ( .A(G131), .B(KEYINPUT61), .Z(n1349) );
XNOR2_X1 U1096 ( .A(n1366), .B(G478), .ZN(n1096) );
OR2_X1 U1097 ( .A1(n1158), .A2(G902), .ZN(n1366) );
XNOR2_X1 U1098 ( .A(n1367), .B(n1368), .ZN(n1158) );
XOR2_X1 U1099 ( .A(n1369), .B(n1370), .Z(n1368) );
XNOR2_X1 U1100 ( .A(n1371), .B(n1372), .ZN(n1370) );
NAND2_X1 U1101 ( .A1(KEYINPUT51), .A2(n1301), .ZN(n1372) );
INV_X1 U1102 ( .A(G116), .ZN(n1301) );
NAND2_X1 U1103 ( .A1(KEYINPUT28), .A2(G128), .ZN(n1371) );
NAND2_X1 U1104 ( .A1(n1340), .A2(G217), .ZN(n1369) );
AND2_X1 U1105 ( .A1(G234), .A2(n1048), .ZN(n1340) );
INV_X1 U1106 ( .A(G953), .ZN(n1048) );
XOR2_X1 U1107 ( .A(n1373), .B(n1374), .Z(n1367) );
XOR2_X1 U1108 ( .A(G122), .B(G107), .Z(n1374) );
XNOR2_X1 U1109 ( .A(G134), .B(G143), .ZN(n1373) );
endmodule


