//Key = 0110001000011011001100001100010001110101001101011100010011010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326;

XNOR2_X1 U728 ( .A(G107), .B(n1002), .ZN(G9) );
NAND3_X1 U729 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1002) );
NOR2_X1 U730 ( .A1(n1006), .A2(n1007), .ZN(G75) );
NOR4_X1 U731 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1007) );
NAND3_X1 U732 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1008) );
NAND2_X1 U733 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U734 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND4_X1 U735 ( .A1(n1019), .A2(n1020), .A3(n1004), .A4(n1021), .ZN(n1018) );
XOR2_X1 U736 ( .A(KEYINPUT34), .B(n1022), .Z(n1017) );
NOR3_X1 U737 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NAND3_X1 U738 ( .A1(n1026), .A2(n1004), .A3(n1020), .ZN(n1023) );
NAND4_X1 U739 ( .A1(n1019), .A2(n1027), .A3(n1028), .A4(n1025), .ZN(n1012) );
NAND2_X1 U740 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND3_X1 U741 ( .A1(n1004), .A2(n1031), .A3(n1015), .ZN(n1030) );
NAND2_X1 U742 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U743 ( .A1(n1020), .A2(n1034), .ZN(n1029) );
NAND2_X1 U744 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U745 ( .A1(n1015), .A2(n1037), .ZN(n1036) );
OR2_X1 U746 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U747 ( .A1(n1004), .A2(n1040), .ZN(n1035) );
NAND2_X1 U748 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U749 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
INV_X1 U750 ( .A(n1024), .ZN(n1019) );
NOR3_X1 U751 ( .A1(n1011), .A2(G952), .A3(n1045), .ZN(n1006) );
INV_X1 U752 ( .A(n1013), .ZN(n1045) );
NAND4_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1013) );
NOR4_X1 U754 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1049) );
XNOR2_X1 U755 ( .A(n1054), .B(n1055), .ZN(n1053) );
NAND2_X1 U756 ( .A1(KEYINPUT59), .A2(n1056), .ZN(n1054) );
INV_X1 U757 ( .A(n1057), .ZN(n1050) );
NOR2_X1 U758 ( .A1(n1058), .A2(n1059), .ZN(n1048) );
XOR2_X1 U759 ( .A(n1060), .B(n1061), .Z(n1059) );
XOR2_X1 U760 ( .A(KEYINPUT47), .B(n1062), .Z(n1061) );
NOR2_X1 U761 ( .A1(KEYINPUT46), .A2(G478), .ZN(n1060) );
XNOR2_X1 U762 ( .A(KEYINPUT37), .B(n1026), .ZN(n1047) );
NAND2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(G72) );
NAND2_X1 U764 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1063) );
INV_X1 U766 ( .A(n1065), .ZN(n1068) );
NOR2_X1 U767 ( .A1(KEYINPUT5), .A2(n1069), .ZN(n1065) );
XOR2_X1 U768 ( .A(n1070), .B(n1071), .Z(n1069) );
NOR2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XNOR2_X1 U770 ( .A(n1074), .B(n1075), .ZN(n1073) );
NOR2_X1 U771 ( .A1(KEYINPUT51), .A2(n1076), .ZN(n1075) );
XNOR2_X1 U772 ( .A(n1077), .B(n1078), .ZN(n1076) );
XOR2_X1 U773 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND2_X1 U774 ( .A1(n1081), .A2(n1082), .ZN(n1070) );
NAND2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XNOR2_X1 U776 ( .A(KEYINPUT33), .B(n1085), .ZN(n1084) );
NAND2_X1 U777 ( .A1(n1086), .A2(n1066), .ZN(n1067) );
NAND2_X1 U778 ( .A1(G953), .A2(n1087), .ZN(n1066) );
INV_X1 U779 ( .A(G227), .ZN(n1087) );
INV_X1 U780 ( .A(n1072), .ZN(n1086) );
XOR2_X1 U781 ( .A(n1088), .B(n1089), .Z(G69) );
NOR2_X1 U782 ( .A1(n1090), .A2(n1081), .ZN(n1089) );
NOR2_X1 U783 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U784 ( .A1(n1093), .A2(n1094), .ZN(n1088) );
NAND2_X1 U785 ( .A1(n1095), .A2(n1081), .ZN(n1094) );
XNOR2_X1 U786 ( .A(n1010), .B(n1096), .ZN(n1095) );
OR3_X1 U787 ( .A1(n1092), .A2(n1096), .A3(n1081), .ZN(n1093) );
XNOR2_X1 U788 ( .A(n1097), .B(n1098), .ZN(n1096) );
XOR2_X1 U789 ( .A(n1099), .B(KEYINPUT19), .Z(n1097) );
NAND2_X1 U790 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U791 ( .A1(n1102), .A2(n1103), .ZN(G66) );
XOR2_X1 U792 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U793 ( .A1(KEYINPUT24), .A2(n1106), .ZN(n1105) );
NAND2_X1 U794 ( .A1(n1107), .A2(n1108), .ZN(n1104) );
XOR2_X1 U795 ( .A(n1109), .B(KEYINPUT45), .Z(n1107) );
NAND2_X1 U796 ( .A1(KEYINPUT56), .A2(G217), .ZN(n1109) );
NOR2_X1 U797 ( .A1(n1102), .A2(n1110), .ZN(G63) );
NOR3_X1 U798 ( .A1(n1062), .A2(n1111), .A3(n1112), .ZN(n1110) );
AND3_X1 U799 ( .A1(n1113), .A2(G478), .A3(n1108), .ZN(n1112) );
NOR2_X1 U800 ( .A1(n1114), .A2(n1113), .ZN(n1111) );
NOR2_X1 U801 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U802 ( .A1(n1102), .A2(n1117), .ZN(G60) );
XOR2_X1 U803 ( .A(n1118), .B(n1119), .Z(n1117) );
AND2_X1 U804 ( .A1(G475), .A2(n1108), .ZN(n1118) );
XOR2_X1 U805 ( .A(n1120), .B(n1121), .Z(G6) );
XNOR2_X1 U806 ( .A(G104), .B(KEYINPUT21), .ZN(n1121) );
NOR2_X1 U807 ( .A1(n1102), .A2(n1122), .ZN(G57) );
XOR2_X1 U808 ( .A(n1123), .B(n1124), .Z(n1122) );
XNOR2_X1 U809 ( .A(n1125), .B(n1126), .ZN(n1124) );
XNOR2_X1 U810 ( .A(n1127), .B(n1128), .ZN(n1126) );
NOR2_X1 U811 ( .A1(n1056), .A2(n1129), .ZN(n1128) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1123) );
XNOR2_X1 U813 ( .A(G137), .B(n1132), .ZN(n1131) );
NOR2_X1 U814 ( .A1(KEYINPUT41), .A2(n1133), .ZN(n1132) );
XNOR2_X1 U815 ( .A(G101), .B(n1134), .ZN(n1133) );
NAND2_X1 U816 ( .A1(KEYINPUT11), .A2(n1135), .ZN(n1130) );
XOR2_X1 U817 ( .A(KEYINPUT35), .B(n1136), .Z(n1135) );
NOR2_X1 U818 ( .A1(n1102), .A2(n1137), .ZN(G54) );
XOR2_X1 U819 ( .A(n1138), .B(n1139), .Z(n1137) );
XNOR2_X1 U820 ( .A(G140), .B(n1140), .ZN(n1139) );
NAND2_X1 U821 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XOR2_X1 U822 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U823 ( .A(KEYINPUT58), .B(KEYINPUT38), .ZN(n1141) );
XOR2_X1 U824 ( .A(n1145), .B(n1146), .Z(n1138) );
AND2_X1 U825 ( .A1(G469), .A2(n1108), .ZN(n1146) );
NOR2_X1 U826 ( .A1(n1102), .A2(n1147), .ZN(G51) );
XNOR2_X1 U827 ( .A(n1148), .B(n1149), .ZN(n1147) );
XOR2_X1 U828 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR3_X1 U829 ( .A1(n1129), .A2(KEYINPUT8), .A3(n1152), .ZN(n1151) );
INV_X1 U830 ( .A(n1108), .ZN(n1129) );
NOR2_X1 U831 ( .A1(n1153), .A2(n1115), .ZN(n1108) );
NOR2_X1 U832 ( .A1(n1009), .A2(n1154), .ZN(n1115) );
XOR2_X1 U833 ( .A(KEYINPUT31), .B(n1010), .Z(n1154) );
NAND4_X1 U834 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1010) );
AND4_X1 U835 ( .A1(n1159), .A2(n1160), .A3(n1120), .A4(n1161), .ZN(n1158) );
NAND3_X1 U836 ( .A1(n1003), .A2(n1004), .A3(n1162), .ZN(n1120) );
NOR3_X1 U837 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1157) );
NOR2_X1 U838 ( .A1(n1041), .A2(n1166), .ZN(n1165) );
NOR4_X1 U839 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1164) );
NOR2_X1 U840 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR3_X1 U841 ( .A1(n1033), .A2(n1173), .A3(n1174), .ZN(n1172) );
AND3_X1 U842 ( .A1(KEYINPUT28), .A2(n1020), .A3(n1039), .ZN(n1171) );
NOR2_X1 U843 ( .A1(KEYINPUT28), .A2(n1175), .ZN(n1163) );
OR4_X1 U844 ( .A1(n1033), .A2(n1174), .A3(n1173), .A4(KEYINPUT23), .ZN(n1155) );
NOR2_X1 U845 ( .A1(n1003), .A2(KEYINPUT23), .ZN(n1173) );
INV_X1 U846 ( .A(n1004), .ZN(n1174) );
INV_X1 U847 ( .A(n1005), .ZN(n1033) );
NAND2_X1 U848 ( .A1(n1083), .A2(n1085), .ZN(n1009) );
AND4_X1 U849 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1083) );
AND4_X1 U850 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1179) );
NAND4_X1 U851 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1162), .ZN(n1178) );
XNOR2_X1 U852 ( .A(n1187), .B(KEYINPUT26), .ZN(n1184) );
NOR2_X1 U853 ( .A1(n1188), .A2(n1189), .ZN(n1150) );
XNOR2_X1 U854 ( .A(KEYINPUT9), .B(n1190), .ZN(n1189) );
NOR2_X1 U855 ( .A1(n1081), .A2(G952), .ZN(n1102) );
XNOR2_X1 U856 ( .A(G146), .B(n1176), .ZN(G48) );
NAND4_X1 U857 ( .A1(n1162), .A2(n1191), .A3(n1021), .A4(n1192), .ZN(n1176) );
XNOR2_X1 U858 ( .A(G143), .B(n1085), .ZN(G45) );
NAND2_X1 U859 ( .A1(n1193), .A2(n1194), .ZN(n1085) );
XNOR2_X1 U860 ( .A(G140), .B(n1195), .ZN(G42) );
NAND3_X1 U861 ( .A1(n1039), .A2(n1162), .A3(n1196), .ZN(n1195) );
NOR3_X1 U862 ( .A1(n1197), .A2(n1187), .A3(n1198), .ZN(n1196) );
XNOR2_X1 U863 ( .A(n1015), .B(KEYINPUT4), .ZN(n1197) );
XNOR2_X1 U864 ( .A(n1177), .B(n1199), .ZN(G39) );
NOR2_X1 U865 ( .A1(KEYINPUT44), .A2(n1200), .ZN(n1199) );
INV_X1 U866 ( .A(G137), .ZN(n1200) );
NAND4_X1 U867 ( .A1(n1020), .A2(n1185), .A3(n1192), .A4(n1201), .ZN(n1177) );
NOR3_X1 U868 ( .A1(n1198), .A2(n1202), .A3(n1058), .ZN(n1185) );
INV_X1 U869 ( .A(n1021), .ZN(n1198) );
XNOR2_X1 U870 ( .A(G134), .B(n1183), .ZN(G36) );
NAND3_X1 U871 ( .A1(n1015), .A2(n1005), .A3(n1193), .ZN(n1183) );
XNOR2_X1 U872 ( .A(G131), .B(n1182), .ZN(G33) );
NAND3_X1 U873 ( .A1(n1193), .A2(n1015), .A3(n1162), .ZN(n1182) );
INV_X1 U874 ( .A(n1058), .ZN(n1015) );
NAND2_X1 U875 ( .A1(n1044), .A2(n1203), .ZN(n1058) );
AND3_X1 U876 ( .A1(n1021), .A2(n1201), .A3(n1038), .ZN(n1193) );
XOR2_X1 U877 ( .A(n1204), .B(KEYINPUT52), .Z(n1021) );
XOR2_X1 U878 ( .A(n1181), .B(n1205), .Z(G30) );
XNOR2_X1 U879 ( .A(KEYINPUT57), .B(n1206), .ZN(n1205) );
NAND4_X1 U880 ( .A1(n1191), .A2(n1005), .A3(n1204), .A4(n1192), .ZN(n1181) );
XNOR2_X1 U881 ( .A(G101), .B(n1156), .ZN(G3) );
NAND3_X1 U882 ( .A1(n1038), .A2(n1003), .A3(n1020), .ZN(n1156) );
XNOR2_X1 U883 ( .A(G125), .B(n1180), .ZN(G27) );
NAND3_X1 U884 ( .A1(n1162), .A2(n1191), .A3(n1207), .ZN(n1180) );
AND3_X1 U885 ( .A1(n1186), .A2(n1025), .A3(n1027), .ZN(n1207) );
NOR3_X1 U886 ( .A1(n1202), .A2(n1187), .A3(n1041), .ZN(n1191) );
INV_X1 U887 ( .A(n1201), .ZN(n1187) );
NAND2_X1 U888 ( .A1(n1208), .A2(n1024), .ZN(n1201) );
NAND3_X1 U889 ( .A1(G902), .A2(n1209), .A3(n1072), .ZN(n1208) );
NOR2_X1 U890 ( .A1(G900), .A2(n1081), .ZN(n1072) );
XNOR2_X1 U891 ( .A(G122), .B(n1161), .ZN(G24) );
NAND3_X1 U892 ( .A1(n1194), .A2(n1004), .A3(n1210), .ZN(n1161) );
NOR2_X1 U893 ( .A1(n1211), .A2(n1192), .ZN(n1004) );
AND3_X1 U894 ( .A1(n1212), .A2(n1213), .A3(n1167), .ZN(n1194) );
NAND2_X1 U895 ( .A1(n1214), .A2(n1215), .ZN(G21) );
NAND2_X1 U896 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U897 ( .A1(G119), .A2(n1218), .ZN(n1214) );
NAND2_X1 U898 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NAND2_X1 U899 ( .A1(KEYINPUT32), .A2(n1221), .ZN(n1220) );
OR2_X1 U900 ( .A1(n1216), .A2(KEYINPUT32), .ZN(n1219) );
AND2_X1 U901 ( .A1(KEYINPUT29), .A2(n1221), .ZN(n1216) );
INV_X1 U902 ( .A(n1160), .ZN(n1221) );
NAND3_X1 U903 ( .A1(n1210), .A2(n1020), .A3(n1222), .ZN(n1160) );
NOR3_X1 U904 ( .A1(n1041), .A2(n1202), .A3(n1186), .ZN(n1222) );
XNOR2_X1 U905 ( .A(G116), .B(n1223), .ZN(G18) );
NAND2_X1 U906 ( .A1(n1167), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U907 ( .A(KEYINPUT0), .B(n1166), .ZN(n1224) );
NAND3_X1 U908 ( .A1(n1038), .A2(n1005), .A3(n1210), .ZN(n1166) );
NOR2_X1 U909 ( .A1(n1212), .A2(n1225), .ZN(n1005) );
XOR2_X1 U910 ( .A(n1159), .B(n1226), .Z(G15) );
XNOR2_X1 U911 ( .A(KEYINPUT2), .B(n1227), .ZN(n1226) );
NAND4_X1 U912 ( .A1(n1210), .A2(n1162), .A3(n1038), .A4(n1167), .ZN(n1159) );
NOR2_X1 U913 ( .A1(n1211), .A2(n1186), .ZN(n1038) );
INV_X1 U914 ( .A(n1192), .ZN(n1186) );
INV_X1 U915 ( .A(n1032), .ZN(n1162) );
NAND2_X1 U916 ( .A1(n1225), .A2(n1212), .ZN(n1032) );
AND3_X1 U917 ( .A1(n1025), .A2(n1228), .A3(n1027), .ZN(n1210) );
XOR2_X1 U918 ( .A(n1229), .B(KEYINPUT25), .Z(n1027) );
XOR2_X1 U919 ( .A(n1175), .B(n1230), .Z(G12) );
XNOR2_X1 U920 ( .A(G110), .B(KEYINPUT17), .ZN(n1230) );
NAND3_X1 U921 ( .A1(n1020), .A2(n1003), .A3(n1039), .ZN(n1175) );
NOR2_X1 U922 ( .A1(n1192), .A2(n1202), .ZN(n1039) );
INV_X1 U923 ( .A(n1211), .ZN(n1202) );
NAND3_X1 U924 ( .A1(n1231), .A2(n1232), .A3(n1057), .ZN(n1211) );
NAND2_X1 U925 ( .A1(n1233), .A2(n1234), .ZN(n1057) );
NAND2_X1 U926 ( .A1(KEYINPUT3), .A2(n1234), .ZN(n1232) );
NAND2_X1 U927 ( .A1(n1052), .A2(n1235), .ZN(n1231) );
INV_X1 U928 ( .A(KEYINPUT3), .ZN(n1235) );
NOR2_X1 U929 ( .A1(n1234), .A2(n1233), .ZN(n1052) );
NOR2_X1 U930 ( .A1(n1106), .A2(G902), .ZN(n1233) );
XOR2_X1 U931 ( .A(n1236), .B(n1237), .Z(n1106) );
XOR2_X1 U932 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U933 ( .A(n1240), .B(n1080), .Z(n1239) );
AND3_X1 U934 ( .A1(G221), .A2(n1081), .A3(G234), .ZN(n1240) );
XOR2_X1 U935 ( .A(n1241), .B(n1242), .Z(n1236) );
NOR2_X1 U936 ( .A1(KEYINPUT20), .A2(n1243), .ZN(n1242) );
XNOR2_X1 U937 ( .A(G119), .B(KEYINPUT42), .ZN(n1241) );
NAND2_X1 U938 ( .A1(G217), .A2(n1244), .ZN(n1234) );
XOR2_X1 U939 ( .A(n1055), .B(n1056), .Z(n1192) );
INV_X1 U940 ( .A(G472), .ZN(n1056) );
NAND2_X1 U941 ( .A1(n1245), .A2(n1153), .ZN(n1055) );
XOR2_X1 U942 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U943 ( .A(n1248), .B(n1249), .Z(n1247) );
XNOR2_X1 U944 ( .A(n1250), .B(n1251), .ZN(n1248) );
INV_X1 U945 ( .A(n1127), .ZN(n1251) );
XNOR2_X1 U946 ( .A(n1252), .B(n1253), .ZN(n1127) );
XNOR2_X1 U947 ( .A(KEYINPUT50), .B(n1217), .ZN(n1253) );
XNOR2_X1 U948 ( .A(n1254), .B(n1227), .ZN(n1252) );
NAND2_X1 U949 ( .A1(KEYINPUT43), .A2(n1255), .ZN(n1254) );
INV_X1 U950 ( .A(G116), .ZN(n1255) );
NAND2_X1 U951 ( .A1(n1256), .A2(n1257), .ZN(n1250) );
OR2_X1 U952 ( .A1(n1134), .A2(n1258), .ZN(n1257) );
XOR2_X1 U953 ( .A(n1259), .B(KEYINPUT22), .Z(n1256) );
NAND2_X1 U954 ( .A1(n1258), .A2(n1134), .ZN(n1259) );
NAND3_X1 U955 ( .A1(n1260), .A2(n1081), .A3(G210), .ZN(n1134) );
XOR2_X1 U956 ( .A(G101), .B(KEYINPUT15), .Z(n1258) );
XOR2_X1 U957 ( .A(n1261), .B(n1262), .Z(n1246) );
XOR2_X1 U958 ( .A(KEYINPUT62), .B(KEYINPUT35), .Z(n1262) );
NOR3_X1 U959 ( .A1(n1168), .A2(n1169), .A3(n1041), .ZN(n1003) );
INV_X1 U960 ( .A(n1167), .ZN(n1041) );
NOR2_X1 U961 ( .A1(n1044), .A2(n1043), .ZN(n1167) );
INV_X1 U962 ( .A(n1203), .ZN(n1043) );
NAND2_X1 U963 ( .A1(G214), .A2(n1263), .ZN(n1203) );
XOR2_X1 U964 ( .A(KEYINPUT18), .B(n1264), .Z(n1263) );
NOR2_X1 U965 ( .A1(G237), .A2(G902), .ZN(n1264) );
XNOR2_X1 U966 ( .A(n1265), .B(n1152), .ZN(n1044) );
NAND2_X1 U967 ( .A1(G210), .A2(n1266), .ZN(n1152) );
NAND2_X1 U968 ( .A1(n1260), .A2(n1153), .ZN(n1266) );
NAND2_X1 U969 ( .A1(n1267), .A2(n1268), .ZN(n1265) );
XNOR2_X1 U970 ( .A(KEYINPUT53), .B(n1153), .ZN(n1268) );
XNOR2_X1 U971 ( .A(n1269), .B(n1270), .ZN(n1267) );
INV_X1 U972 ( .A(n1148), .ZN(n1270) );
XNOR2_X1 U973 ( .A(n1271), .B(n1098), .ZN(n1148) );
XNOR2_X1 U974 ( .A(n1272), .B(n1238), .ZN(n1098) );
NAND2_X1 U975 ( .A1(n1273), .A2(n1101), .ZN(n1271) );
NAND2_X1 U976 ( .A1(n1274), .A2(n1275), .ZN(n1101) );
XNOR2_X1 U977 ( .A(n1227), .B(n1276), .ZN(n1275) );
INV_X1 U978 ( .A(G113), .ZN(n1227) );
XNOR2_X1 U979 ( .A(n1277), .B(n1278), .ZN(n1274) );
INV_X1 U980 ( .A(G101), .ZN(n1277) );
XOR2_X1 U981 ( .A(n1100), .B(KEYINPUT55), .Z(n1273) );
NAND2_X1 U982 ( .A1(n1279), .A2(n1280), .ZN(n1100) );
XNOR2_X1 U983 ( .A(G113), .B(n1276), .ZN(n1280) );
NOR2_X1 U984 ( .A1(KEYINPUT13), .A2(n1281), .ZN(n1276) );
XNOR2_X1 U985 ( .A(G116), .B(n1282), .ZN(n1281) );
XNOR2_X1 U986 ( .A(KEYINPUT61), .B(n1217), .ZN(n1282) );
INV_X1 U987 ( .A(G119), .ZN(n1217) );
XNOR2_X1 U988 ( .A(G101), .B(n1278), .ZN(n1279) );
XOR2_X1 U989 ( .A(n1283), .B(KEYINPUT6), .Z(n1269) );
NAND2_X1 U990 ( .A1(n1190), .A2(n1284), .ZN(n1283) );
INV_X1 U991 ( .A(n1188), .ZN(n1284) );
NOR3_X1 U992 ( .A1(n1285), .A2(G953), .A3(n1091), .ZN(n1188) );
INV_X1 U993 ( .A(G224), .ZN(n1091) );
NAND2_X1 U994 ( .A1(n1285), .A2(n1286), .ZN(n1190) );
NAND2_X1 U995 ( .A1(G224), .A2(n1081), .ZN(n1286) );
XOR2_X1 U996 ( .A(G125), .B(n1136), .Z(n1285) );
XNOR2_X1 U997 ( .A(n1261), .B(G128), .ZN(n1136) );
NAND3_X1 U998 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n1261) );
NAND2_X1 U999 ( .A1(KEYINPUT40), .A2(G143), .ZN(n1289) );
OR3_X1 U1000 ( .A1(n1290), .A2(KEYINPUT40), .A3(G146), .ZN(n1288) );
NAND2_X1 U1001 ( .A1(G146), .A2(n1290), .ZN(n1287) );
NAND2_X1 U1002 ( .A1(KEYINPUT14), .A2(n1291), .ZN(n1290) );
INV_X1 U1003 ( .A(n1228), .ZN(n1169) );
NAND2_X1 U1004 ( .A1(n1024), .A2(n1292), .ZN(n1228) );
NAND4_X1 U1005 ( .A1(G953), .A2(G902), .A3(n1209), .A4(n1092), .ZN(n1292) );
INV_X1 U1006 ( .A(G898), .ZN(n1092) );
NAND3_X1 U1007 ( .A1(n1293), .A2(n1209), .A3(G952), .ZN(n1024) );
NAND2_X1 U1008 ( .A1(G237), .A2(G234), .ZN(n1209) );
INV_X1 U1009 ( .A(n1011), .ZN(n1293) );
XOR2_X1 U1010 ( .A(G953), .B(KEYINPUT36), .Z(n1011) );
INV_X1 U1011 ( .A(n1204), .ZN(n1168) );
NOR2_X1 U1012 ( .A1(n1026), .A2(n1051), .ZN(n1204) );
INV_X1 U1013 ( .A(n1025), .ZN(n1051) );
NAND2_X1 U1014 ( .A1(G221), .A2(n1244), .ZN(n1025) );
NAND2_X1 U1015 ( .A1(G234), .A2(n1153), .ZN(n1244) );
INV_X1 U1016 ( .A(n1229), .ZN(n1026) );
XNOR2_X1 U1017 ( .A(n1294), .B(G469), .ZN(n1229) );
NAND2_X1 U1018 ( .A1(n1295), .A2(n1153), .ZN(n1294) );
INV_X1 U1019 ( .A(G902), .ZN(n1153) );
XOR2_X1 U1020 ( .A(n1296), .B(n1297), .Z(n1295) );
XNOR2_X1 U1021 ( .A(n1298), .B(KEYINPUT16), .ZN(n1297) );
NAND2_X1 U1022 ( .A1(KEYINPUT63), .A2(n1299), .ZN(n1298) );
XOR2_X1 U1023 ( .A(n1300), .B(n1145), .Z(n1299) );
XOR2_X1 U1024 ( .A(n1301), .B(n1238), .Z(n1145) );
XOR2_X1 U1025 ( .A(G110), .B(KEYINPUT1), .Z(n1238) );
NAND2_X1 U1026 ( .A1(G227), .A2(n1081), .ZN(n1301) );
NAND2_X1 U1027 ( .A1(KEYINPUT12), .A2(n1302), .ZN(n1300) );
XOR2_X1 U1028 ( .A(n1143), .B(n1303), .Z(n1296) );
NOR2_X1 U1029 ( .A1(KEYINPUT10), .A2(n1144), .ZN(n1303) );
XNOR2_X1 U1030 ( .A(n1304), .B(G101), .ZN(n1144) );
NAND2_X1 U1031 ( .A1(KEYINPUT49), .A2(n1278), .ZN(n1304) );
XOR2_X1 U1032 ( .A(G107), .B(G104), .Z(n1278) );
XNOR2_X1 U1033 ( .A(n1249), .B(n1077), .ZN(n1143) );
XOR2_X1 U1034 ( .A(G143), .B(n1305), .Z(n1077) );
XOR2_X1 U1035 ( .A(KEYINPUT60), .B(G146), .Z(n1305) );
XNOR2_X1 U1036 ( .A(n1080), .B(n1306), .ZN(n1249) );
INV_X1 U1037 ( .A(n1125), .ZN(n1306) );
XNOR2_X1 U1038 ( .A(n1079), .B(KEYINPUT30), .ZN(n1125) );
XNOR2_X1 U1039 ( .A(G131), .B(G134), .ZN(n1079) );
XNOR2_X1 U1040 ( .A(G137), .B(n1206), .ZN(n1080) );
INV_X1 U1041 ( .A(G128), .ZN(n1206) );
NOR2_X1 U1042 ( .A1(n1213), .A2(n1212), .ZN(n1020) );
XNOR2_X1 U1043 ( .A(n1046), .B(KEYINPUT7), .ZN(n1212) );
XOR2_X1 U1044 ( .A(n1307), .B(G475), .Z(n1046) );
OR2_X1 U1045 ( .A1(n1119), .A2(G902), .ZN(n1307) );
XNOR2_X1 U1046 ( .A(n1308), .B(n1309), .ZN(n1119) );
XNOR2_X1 U1047 ( .A(n1310), .B(n1311), .ZN(n1309) );
NOR2_X1 U1048 ( .A1(KEYINPUT27), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U1049 ( .A(n1291), .B(n1313), .ZN(n1312) );
AND3_X1 U1050 ( .A1(G214), .A2(n1081), .A3(n1260), .ZN(n1313) );
INV_X1 U1051 ( .A(G237), .ZN(n1260) );
INV_X1 U1052 ( .A(G131), .ZN(n1310) );
XNOR2_X1 U1053 ( .A(n1314), .B(n1243), .ZN(n1308) );
XNOR2_X1 U1054 ( .A(G146), .B(n1074), .ZN(n1243) );
XNOR2_X1 U1055 ( .A(G125), .B(n1302), .ZN(n1074) );
INV_X1 U1056 ( .A(G140), .ZN(n1302) );
NAND2_X1 U1057 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
OR2_X1 U1058 ( .A1(n1317), .A2(G104), .ZN(n1316) );
XOR2_X1 U1059 ( .A(n1318), .B(KEYINPUT54), .Z(n1315) );
NAND2_X1 U1060 ( .A1(G104), .A2(n1317), .ZN(n1318) );
XNOR2_X1 U1061 ( .A(G113), .B(n1272), .ZN(n1317) );
INV_X1 U1062 ( .A(n1225), .ZN(n1213) );
XOR2_X1 U1063 ( .A(n1062), .B(n1116), .Z(n1225) );
INV_X1 U1064 ( .A(G478), .ZN(n1116) );
NOR2_X1 U1065 ( .A1(n1113), .A2(G902), .ZN(n1062) );
XOR2_X1 U1066 ( .A(n1319), .B(n1320), .Z(n1113) );
XOR2_X1 U1067 ( .A(n1321), .B(n1322), .Z(n1320) );
XNOR2_X1 U1068 ( .A(n1272), .B(G116), .ZN(n1322) );
INV_X1 U1069 ( .A(G122), .ZN(n1272) );
XNOR2_X1 U1070 ( .A(n1291), .B(G134), .ZN(n1321) );
INV_X1 U1071 ( .A(G143), .ZN(n1291) );
XOR2_X1 U1072 ( .A(n1323), .B(n1324), .Z(n1319) );
XOR2_X1 U1073 ( .A(G107), .B(n1325), .Z(n1324) );
AND3_X1 U1074 ( .A1(G234), .A2(n1081), .A3(G217), .ZN(n1325) );
INV_X1 U1075 ( .A(G953), .ZN(n1081) );
NAND2_X1 U1076 ( .A1(n1326), .A2(KEYINPUT48), .ZN(n1323) );
XNOR2_X1 U1077 ( .A(G128), .B(KEYINPUT39), .ZN(n1326) );
endmodule


