//Key = 0111000001010101001101101111010001000011011000101010011001101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360;

XNOR2_X1 U749 ( .A(G107), .B(n1039), .ZN(G9) );
NOR2_X1 U750 ( .A1(n1040), .A2(n1041), .ZN(G75) );
NOR4_X1 U751 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1041) );
NAND4_X1 U752 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1042) );
NAND2_X1 U753 ( .A1(n1050), .A2(n1051), .ZN(n1047) );
NAND2_X1 U754 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND4_X1 U755 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1053) );
NAND2_X1 U756 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U757 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
OR2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U759 ( .A1(n1064), .A2(n1065), .ZN(n1058) );
NAND2_X1 U760 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND3_X1 U762 ( .A1(n1064), .A2(n1070), .A3(n1060), .ZN(n1052) );
NAND2_X1 U763 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U764 ( .A1(n1073), .A2(n1074), .A3(n1056), .ZN(n1072) );
NAND2_X1 U765 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND3_X1 U766 ( .A1(n1077), .A2(n1078), .A3(n1054), .ZN(n1073) );
INV_X1 U767 ( .A(n1079), .ZN(n1078) );
NAND2_X1 U768 ( .A1(n1080), .A2(n1081), .ZN(n1077) );
NAND2_X1 U769 ( .A1(n1055), .A2(n1082), .ZN(n1071) );
INV_X1 U770 ( .A(n1083), .ZN(n1050) );
NOR3_X1 U771 ( .A1(n1084), .A2(G953), .A3(n1085), .ZN(n1040) );
INV_X1 U772 ( .A(n1048), .ZN(n1085) );
NAND4_X1 U773 ( .A1(n1054), .A2(n1060), .A3(n1086), .A4(n1087), .ZN(n1048) );
NOR4_X1 U774 ( .A1(n1080), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1087) );
XNOR2_X1 U775 ( .A(n1091), .B(n1092), .ZN(n1090) );
XNOR2_X1 U776 ( .A(KEYINPUT33), .B(KEYINPUT0), .ZN(n1091) );
XNOR2_X1 U777 ( .A(n1093), .B(n1094), .ZN(n1089) );
NAND2_X1 U778 ( .A1(KEYINPUT57), .A2(n1095), .ZN(n1093) );
NOR2_X1 U779 ( .A1(n1096), .A2(n1097), .ZN(n1088) );
NOR2_X1 U780 ( .A1(n1098), .A2(G472), .ZN(n1097) );
NOR2_X1 U781 ( .A1(KEYINPUT59), .A2(n1099), .ZN(n1098) );
NOR2_X1 U782 ( .A1(n1100), .A2(KEYINPUT16), .ZN(n1099) );
NOR2_X1 U783 ( .A1(n1101), .A2(n1102), .ZN(n1096) );
NOR2_X1 U784 ( .A1(n1103), .A2(KEYINPUT16), .ZN(n1101) );
NOR2_X1 U785 ( .A1(KEYINPUT59), .A2(n1104), .ZN(n1103) );
XOR2_X1 U786 ( .A(n1105), .B(KEYINPUT15), .Z(n1086) );
NAND2_X1 U787 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U788 ( .A(n1108), .B(KEYINPUT56), .Z(n1106) );
XNOR2_X1 U789 ( .A(KEYINPUT31), .B(n1044), .ZN(n1084) );
INV_X1 U790 ( .A(G952), .ZN(n1044) );
XOR2_X1 U791 ( .A(n1109), .B(n1110), .Z(G72) );
XOR2_X1 U792 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U793 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U794 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U795 ( .A(n1117), .B(n1118), .Z(n1116) );
XNOR2_X1 U796 ( .A(G140), .B(n1119), .ZN(n1115) );
NOR2_X1 U797 ( .A1(G125), .A2(KEYINPUT36), .ZN(n1119) );
XOR2_X1 U798 ( .A(KEYINPUT20), .B(n1120), .Z(n1113) );
NAND3_X1 U799 ( .A1(n1121), .A2(n1122), .A3(KEYINPUT60), .ZN(n1111) );
OR2_X1 U800 ( .A1(n1043), .A2(n1123), .ZN(n1122) );
XNOR2_X1 U801 ( .A(KEYINPUT13), .B(n1049), .ZN(n1121) );
NAND2_X1 U802 ( .A1(G953), .A2(n1124), .ZN(n1109) );
NAND2_X1 U803 ( .A1(G900), .A2(G227), .ZN(n1124) );
NAND2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(G69) );
NAND2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U806 ( .A1(n1129), .A2(n1130), .ZN(n1125) );
NAND2_X1 U807 ( .A1(n1131), .A2(n1128), .ZN(n1130) );
NAND2_X1 U808 ( .A1(G953), .A2(n1132), .ZN(n1128) );
INV_X1 U809 ( .A(G224), .ZN(n1132) );
INV_X1 U810 ( .A(n1133), .ZN(n1131) );
INV_X1 U811 ( .A(n1127), .ZN(n1129) );
XNOR2_X1 U812 ( .A(n1134), .B(n1135), .ZN(n1127) );
NOR2_X1 U813 ( .A1(n1133), .A2(n1136), .ZN(n1135) );
XOR2_X1 U814 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U815 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U816 ( .A1(KEYINPUT30), .A2(n1141), .ZN(n1139) );
XOR2_X1 U817 ( .A(n1142), .B(KEYINPUT42), .Z(n1137) );
NAND2_X1 U818 ( .A1(n1143), .A2(n1049), .ZN(n1134) );
XOR2_X1 U819 ( .A(n1045), .B(KEYINPUT47), .Z(n1143) );
NOR2_X1 U820 ( .A1(n1144), .A2(n1145), .ZN(G66) );
XNOR2_X1 U821 ( .A(n1146), .B(n1147), .ZN(n1145) );
NOR2_X1 U822 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NOR2_X1 U823 ( .A1(n1144), .A2(n1150), .ZN(G63) );
NOR2_X1 U824 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U825 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U826 ( .A1(KEYINPUT35), .A2(n1155), .ZN(n1154) );
NOR2_X1 U827 ( .A1(n1156), .A2(n1149), .ZN(n1153) );
AND2_X1 U828 ( .A1(n1155), .A2(KEYINPUT35), .ZN(n1151) );
INV_X1 U829 ( .A(n1157), .ZN(n1155) );
NOR2_X1 U830 ( .A1(n1144), .A2(n1158), .ZN(G60) );
XOR2_X1 U831 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR3_X1 U832 ( .A1(n1149), .A2(KEYINPUT51), .A3(n1161), .ZN(n1159) );
XNOR2_X1 U833 ( .A(G104), .B(n1162), .ZN(G6) );
NOR2_X1 U834 ( .A1(n1144), .A2(n1163), .ZN(G57) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(n1163) );
XNOR2_X1 U836 ( .A(n1166), .B(n1167), .ZN(n1165) );
NAND2_X1 U837 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U838 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
INV_X1 U839 ( .A(KEYINPUT45), .ZN(n1171) );
XOR2_X1 U840 ( .A(n1118), .B(n1172), .Z(n1170) );
NAND3_X1 U841 ( .A1(n1172), .A2(n1118), .A3(KEYINPUT45), .ZN(n1168) );
XOR2_X1 U842 ( .A(n1173), .B(n1174), .Z(n1164) );
NOR2_X1 U843 ( .A1(n1104), .A2(n1149), .ZN(n1174) );
NAND2_X1 U844 ( .A1(n1175), .A2(KEYINPUT25), .ZN(n1173) );
XNOR2_X1 U845 ( .A(G101), .B(n1176), .ZN(n1175) );
NOR2_X1 U846 ( .A1(KEYINPUT12), .A2(n1177), .ZN(n1176) );
NOR2_X1 U847 ( .A1(n1144), .A2(n1178), .ZN(G54) );
XNOR2_X1 U848 ( .A(n1179), .B(n1180), .ZN(n1178) );
XNOR2_X1 U849 ( .A(n1181), .B(n1182), .ZN(n1180) );
NOR3_X1 U850 ( .A1(n1095), .A2(KEYINPUT8), .A3(n1149), .ZN(n1182) );
INV_X1 U851 ( .A(G469), .ZN(n1095) );
NAND2_X1 U852 ( .A1(KEYINPUT48), .A2(n1117), .ZN(n1181) );
NOR2_X1 U853 ( .A1(n1144), .A2(n1183), .ZN(G51) );
XOR2_X1 U854 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U855 ( .A1(n1186), .A2(n1149), .ZN(n1185) );
NAND2_X1 U856 ( .A1(G902), .A2(n1187), .ZN(n1149) );
NAND3_X1 U857 ( .A1(n1188), .A2(n1046), .A3(n1189), .ZN(n1187) );
XOR2_X1 U858 ( .A(n1045), .B(KEYINPUT58), .Z(n1189) );
NAND4_X1 U859 ( .A1(n1190), .A2(n1162), .A3(n1191), .A4(n1192), .ZN(n1045) );
NOR4_X1 U860 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
INV_X1 U861 ( .A(n1039), .ZN(n1196) );
NAND4_X1 U862 ( .A1(n1197), .A2(n1198), .A3(n1054), .A4(n1062), .ZN(n1039) );
NAND2_X1 U863 ( .A1(n1197), .A2(n1199), .ZN(n1191) );
NAND2_X1 U864 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XNOR2_X1 U865 ( .A(n1202), .B(KEYINPUT43), .ZN(n1200) );
NAND4_X1 U866 ( .A1(n1063), .A2(n1197), .A3(n1054), .A4(n1198), .ZN(n1162) );
NAND3_X1 U867 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1190) );
INV_X1 U868 ( .A(n1206), .ZN(n1205) );
OR2_X1 U869 ( .A1(n1207), .A2(KEYINPUT14), .ZN(n1204) );
NAND2_X1 U870 ( .A1(KEYINPUT14), .A2(n1208), .ZN(n1203) );
NAND3_X1 U871 ( .A1(n1209), .A2(n1066), .A3(n1055), .ZN(n1208) );
XNOR2_X1 U872 ( .A(n1123), .B(KEYINPUT4), .ZN(n1046) );
NAND4_X1 U873 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1123) );
OR2_X1 U874 ( .A1(n1214), .A2(n1215), .ZN(n1211) );
NAND2_X1 U875 ( .A1(n1216), .A2(n1197), .ZN(n1210) );
INV_X1 U876 ( .A(n1043), .ZN(n1188) );
NAND4_X1 U877 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1043) );
OR2_X1 U878 ( .A1(n1221), .A2(n1066), .ZN(n1217) );
INV_X1 U879 ( .A(n1197), .ZN(n1066) );
INV_X1 U880 ( .A(G210), .ZN(n1186) );
NOR2_X1 U881 ( .A1(n1222), .A2(n1223), .ZN(n1184) );
XOR2_X1 U882 ( .A(n1224), .B(KEYINPUT39), .Z(n1223) );
NAND2_X1 U883 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
NOR2_X1 U884 ( .A1(n1225), .A2(n1226), .ZN(n1222) );
XOR2_X1 U885 ( .A(n1227), .B(n1172), .Z(n1225) );
XNOR2_X1 U886 ( .A(n1228), .B(n1229), .ZN(n1227) );
NAND2_X1 U887 ( .A1(KEYINPUT21), .A2(n1230), .ZN(n1228) );
INV_X1 U888 ( .A(G125), .ZN(n1230) );
AND2_X1 U889 ( .A1(n1231), .A2(G953), .ZN(n1144) );
XNOR2_X1 U890 ( .A(G952), .B(KEYINPUT44), .ZN(n1231) );
XNOR2_X1 U891 ( .A(G146), .B(n1218), .ZN(G48) );
NAND3_X1 U892 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1218) );
XOR2_X1 U893 ( .A(n1235), .B(n1236), .Z(G45) );
NAND2_X1 U894 ( .A1(KEYINPUT38), .A2(G143), .ZN(n1236) );
NAND2_X1 U895 ( .A1(n1237), .A2(n1197), .ZN(n1235) );
XOR2_X1 U896 ( .A(n1221), .B(KEYINPUT3), .Z(n1237) );
NAND4_X1 U897 ( .A1(n1082), .A2(n1232), .A3(n1238), .A4(n1239), .ZN(n1221) );
XNOR2_X1 U898 ( .A(G140), .B(n1219), .ZN(G42) );
NAND3_X1 U899 ( .A1(n1056), .A2(n1240), .A3(n1063), .ZN(n1219) );
XNOR2_X1 U900 ( .A(G137), .B(n1220), .ZN(G39) );
NAND3_X1 U901 ( .A1(n1064), .A2(n1233), .A3(n1240), .ZN(n1220) );
AND3_X1 U902 ( .A1(n1060), .A2(n1075), .A3(n1232), .ZN(n1240) );
XOR2_X1 U903 ( .A(G134), .B(n1241), .Z(G36) );
NOR2_X1 U904 ( .A1(n1242), .A2(n1215), .ZN(n1241) );
XOR2_X1 U905 ( .A(n1214), .B(KEYINPUT5), .Z(n1242) );
NAND3_X1 U906 ( .A1(n1232), .A2(n1062), .A3(n1082), .ZN(n1214) );
XNOR2_X1 U907 ( .A(G131), .B(n1212), .ZN(G33) );
NAND4_X1 U908 ( .A1(n1082), .A2(n1063), .A3(n1232), .A4(n1060), .ZN(n1212) );
INV_X1 U909 ( .A(n1215), .ZN(n1060) );
NAND2_X1 U910 ( .A1(n1069), .A2(n1243), .ZN(n1215) );
XOR2_X1 U911 ( .A(n1244), .B(n1245), .Z(G30) );
NAND2_X1 U912 ( .A1(KEYINPUT22), .A2(G128), .ZN(n1245) );
NAND2_X1 U913 ( .A1(n1197), .A2(n1246), .ZN(n1244) );
XOR2_X1 U914 ( .A(KEYINPUT7), .B(n1216), .Z(n1246) );
AND4_X1 U915 ( .A1(n1232), .A2(n1062), .A3(n1075), .A4(n1233), .ZN(n1216) );
AND2_X1 U916 ( .A1(n1079), .A2(n1247), .ZN(n1232) );
XOR2_X1 U917 ( .A(n1248), .B(n1249), .Z(G3) );
XOR2_X1 U918 ( .A(KEYINPUT11), .B(G101), .Z(n1249) );
NAND3_X1 U919 ( .A1(n1202), .A2(n1197), .A3(KEYINPUT19), .ZN(n1248) );
AND4_X1 U920 ( .A1(n1082), .A2(n1064), .A3(n1079), .A4(n1209), .ZN(n1202) );
XOR2_X1 U921 ( .A(n1213), .B(n1250), .Z(G27) );
NAND2_X1 U922 ( .A1(KEYINPUT54), .A2(G125), .ZN(n1250) );
NAND4_X1 U923 ( .A1(n1055), .A2(n1234), .A3(n1056), .A4(n1247), .ZN(n1213) );
NAND2_X1 U924 ( .A1(n1083), .A2(n1251), .ZN(n1247) );
NAND3_X1 U925 ( .A1(n1120), .A2(n1252), .A3(n1253), .ZN(n1251) );
XNOR2_X1 U926 ( .A(G902), .B(KEYINPUT27), .ZN(n1253) );
NOR2_X1 U927 ( .A1(n1049), .A2(G900), .ZN(n1120) );
AND3_X1 U928 ( .A1(n1197), .A2(n1075), .A3(n1063), .ZN(n1234) );
XOR2_X1 U929 ( .A(G122), .B(n1195), .Z(G24) );
AND3_X1 U930 ( .A1(n1054), .A2(n1207), .A3(n1254), .ZN(n1195) );
NOR3_X1 U931 ( .A1(n1233), .A2(n1255), .A3(n1092), .ZN(n1254) );
INV_X1 U932 ( .A(n1238), .ZN(n1092) );
INV_X1 U933 ( .A(n1075), .ZN(n1054) );
XOR2_X1 U934 ( .A(G119), .B(n1256), .Z(G21) );
NOR3_X1 U935 ( .A1(n1206), .A2(KEYINPUT55), .A3(n1257), .ZN(n1256) );
NAND3_X1 U936 ( .A1(n1075), .A2(n1233), .A3(n1064), .ZN(n1206) );
XOR2_X1 U937 ( .A(G116), .B(n1194), .Z(G18) );
AND3_X1 U938 ( .A1(n1082), .A2(n1062), .A3(n1207), .ZN(n1194) );
NAND2_X1 U939 ( .A1(n1258), .A2(n1259), .ZN(n1062) );
NAND2_X1 U940 ( .A1(n1064), .A2(n1260), .ZN(n1259) );
INV_X1 U941 ( .A(KEYINPUT63), .ZN(n1260) );
NAND3_X1 U942 ( .A1(n1255), .A2(n1238), .A3(KEYINPUT63), .ZN(n1258) );
XOR2_X1 U943 ( .A(G113), .B(n1193), .Z(G15) );
AND3_X1 U944 ( .A1(n1082), .A2(n1063), .A3(n1207), .ZN(n1193) );
INV_X1 U945 ( .A(n1257), .ZN(n1207) );
NAND3_X1 U946 ( .A1(n1197), .A2(n1209), .A3(n1055), .ZN(n1257) );
INV_X1 U947 ( .A(n1076), .ZN(n1055) );
NAND2_X1 U948 ( .A1(n1081), .A2(n1261), .ZN(n1076) );
NOR2_X1 U949 ( .A1(n1238), .A2(n1255), .ZN(n1063) );
INV_X1 U950 ( .A(n1239), .ZN(n1255) );
NOR2_X1 U951 ( .A1(n1075), .A2(n1056), .ZN(n1082) );
XNOR2_X1 U952 ( .A(G110), .B(n1262), .ZN(G12) );
NAND2_X1 U953 ( .A1(n1263), .A2(n1197), .ZN(n1262) );
NOR2_X1 U954 ( .A1(n1069), .A2(n1068), .ZN(n1197) );
INV_X1 U955 ( .A(n1243), .ZN(n1068) );
NAND2_X1 U956 ( .A1(G214), .A2(n1264), .ZN(n1243) );
XOR2_X1 U957 ( .A(n1265), .B(n1266), .Z(n1069) );
AND2_X1 U958 ( .A1(n1264), .A2(G210), .ZN(n1266) );
NAND2_X1 U959 ( .A1(n1267), .A2(n1268), .ZN(n1264) );
XNOR2_X1 U960 ( .A(G237), .B(KEYINPUT37), .ZN(n1267) );
NAND2_X1 U961 ( .A1(n1269), .A2(n1268), .ZN(n1265) );
XOR2_X1 U962 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U963 ( .A(n1272), .B(n1226), .Z(n1271) );
XNOR2_X1 U964 ( .A(n1273), .B(n1274), .ZN(n1226) );
XNOR2_X1 U965 ( .A(n1141), .B(n1140), .ZN(n1274) );
XNOR2_X1 U966 ( .A(n1275), .B(G122), .ZN(n1140) );
NAND2_X1 U967 ( .A1(n1276), .A2(n1277), .ZN(n1141) );
NAND2_X1 U968 ( .A1(G101), .A2(n1278), .ZN(n1277) );
XOR2_X1 U969 ( .A(n1279), .B(KEYINPUT62), .Z(n1276) );
OR2_X1 U970 ( .A1(n1278), .A2(G101), .ZN(n1279) );
XNOR2_X1 U971 ( .A(G104), .B(n1280), .ZN(n1278) );
XOR2_X1 U972 ( .A(n1142), .B(KEYINPUT9), .Z(n1273) );
NAND2_X1 U973 ( .A1(n1281), .A2(n1282), .ZN(n1142) );
NAND2_X1 U974 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NAND2_X1 U975 ( .A1(G113), .A2(n1285), .ZN(n1284) );
OR2_X1 U976 ( .A1(KEYINPUT32), .A2(KEYINPUT53), .ZN(n1285) );
NAND3_X1 U977 ( .A1(n1286), .A2(n1287), .A3(KEYINPUT53), .ZN(n1281) );
OR2_X1 U978 ( .A1(G113), .A2(KEYINPUT32), .ZN(n1287) );
NAND2_X1 U979 ( .A1(G113), .A2(n1288), .ZN(n1286) );
OR2_X1 U980 ( .A1(n1283), .A2(KEYINPUT32), .ZN(n1288) );
NAND2_X1 U981 ( .A1(n1289), .A2(n1290), .ZN(n1272) );
OR2_X1 U982 ( .A1(KEYINPUT23), .A2(n1229), .ZN(n1290) );
NAND2_X1 U983 ( .A1(KEYINPUT17), .A2(n1229), .ZN(n1289) );
NAND2_X1 U984 ( .A1(G224), .A2(n1049), .ZN(n1229) );
XNOR2_X1 U985 ( .A(G125), .B(n1172), .ZN(n1270) );
XOR2_X1 U986 ( .A(n1201), .B(KEYINPUT2), .Z(n1263) );
NAND3_X1 U987 ( .A1(n1064), .A2(n1075), .A3(n1198), .ZN(n1201) );
AND3_X1 U988 ( .A1(n1056), .A2(n1209), .A3(n1079), .ZN(n1198) );
NOR2_X1 U989 ( .A1(n1081), .A2(n1080), .ZN(n1079) );
INV_X1 U990 ( .A(n1261), .ZN(n1080) );
NAND2_X1 U991 ( .A1(G221), .A2(n1291), .ZN(n1261) );
XNOR2_X1 U992 ( .A(n1094), .B(n1292), .ZN(n1081) );
NOR2_X1 U993 ( .A1(G469), .A2(KEYINPUT28), .ZN(n1292) );
NAND3_X1 U994 ( .A1(n1293), .A2(n1294), .A3(n1268), .ZN(n1094) );
NAND3_X1 U995 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1294) );
INV_X1 U996 ( .A(KEYINPUT41), .ZN(n1297) );
XNOR2_X1 U997 ( .A(n1298), .B(n1299), .ZN(n1295) );
NAND2_X1 U998 ( .A1(n1300), .A2(KEYINPUT41), .ZN(n1293) );
XNOR2_X1 U999 ( .A(n1301), .B(n1179), .ZN(n1300) );
XNOR2_X1 U1000 ( .A(n1296), .B(n1299), .ZN(n1179) );
XOR2_X1 U1001 ( .A(n1302), .B(n1303), .Z(n1299) );
XNOR2_X1 U1002 ( .A(n1304), .B(n1305), .ZN(n1303) );
NOR2_X1 U1003 ( .A1(G107), .A2(KEYINPUT10), .ZN(n1305) );
XNOR2_X1 U1004 ( .A(n1306), .B(n1307), .ZN(n1296) );
XNOR2_X1 U1005 ( .A(G140), .B(n1275), .ZN(n1307) );
NAND2_X1 U1006 ( .A1(G227), .A2(n1049), .ZN(n1306) );
INV_X1 U1007 ( .A(n1298), .ZN(n1301) );
XOR2_X1 U1008 ( .A(n1117), .B(KEYINPUT24), .Z(n1298) );
XOR2_X1 U1009 ( .A(G128), .B(n1308), .Z(n1117) );
NOR2_X1 U1010 ( .A1(KEYINPUT34), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1011 ( .A(n1310), .B(n1311), .Z(n1309) );
NOR2_X1 U1012 ( .A1(KEYINPUT40), .A2(n1312), .ZN(n1311) );
XOR2_X1 U1013 ( .A(KEYINPUT61), .B(G143), .Z(n1312) );
XNOR2_X1 U1014 ( .A(G146), .B(KEYINPUT1), .ZN(n1310) );
NAND2_X1 U1015 ( .A1(n1083), .A2(n1313), .ZN(n1209) );
NAND3_X1 U1016 ( .A1(n1133), .A2(n1252), .A3(G902), .ZN(n1313) );
NOR2_X1 U1017 ( .A1(G898), .A2(n1049), .ZN(n1133) );
NAND3_X1 U1018 ( .A1(n1252), .A2(n1049), .A3(G952), .ZN(n1083) );
NAND2_X1 U1019 ( .A1(G234), .A2(G237), .ZN(n1252) );
INV_X1 U1020 ( .A(n1233), .ZN(n1056) );
XNOR2_X1 U1021 ( .A(n1100), .B(n1104), .ZN(n1233) );
INV_X1 U1022 ( .A(G472), .ZN(n1104) );
INV_X1 U1023 ( .A(n1102), .ZN(n1100) );
NAND2_X1 U1024 ( .A1(n1314), .A2(n1268), .ZN(n1102) );
XOR2_X1 U1025 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1026 ( .A(n1166), .B(n1172), .Z(n1316) );
XNOR2_X1 U1027 ( .A(n1317), .B(n1318), .ZN(n1172) );
XNOR2_X1 U1028 ( .A(KEYINPUT61), .B(G146), .ZN(n1317) );
XNOR2_X1 U1029 ( .A(G113), .B(n1283), .ZN(n1166) );
XNOR2_X1 U1030 ( .A(G116), .B(G119), .ZN(n1283) );
XNOR2_X1 U1031 ( .A(n1302), .B(n1177), .ZN(n1315) );
NAND2_X1 U1032 ( .A1(n1319), .A2(G210), .ZN(n1177) );
XOR2_X1 U1033 ( .A(G101), .B(n1118), .Z(n1302) );
XOR2_X1 U1034 ( .A(n1320), .B(n1321), .Z(n1118) );
XNOR2_X1 U1035 ( .A(KEYINPUT29), .B(n1322), .ZN(n1321) );
XNOR2_X1 U1036 ( .A(G131), .B(G134), .ZN(n1320) );
XOR2_X1 U1037 ( .A(n1323), .B(n1148), .Z(n1075) );
NAND2_X1 U1038 ( .A1(G217), .A2(n1291), .ZN(n1148) );
NAND2_X1 U1039 ( .A1(G234), .A2(n1268), .ZN(n1291) );
NAND2_X1 U1040 ( .A1(n1146), .A2(n1268), .ZN(n1323) );
XNOR2_X1 U1041 ( .A(n1324), .B(n1325), .ZN(n1146) );
XOR2_X1 U1042 ( .A(n1326), .B(n1327), .Z(n1325) );
NAND2_X1 U1043 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NAND2_X1 U1044 ( .A1(n1330), .A2(n1322), .ZN(n1329) );
XOR2_X1 U1045 ( .A(KEYINPUT50), .B(n1331), .Z(n1328) );
NOR2_X1 U1046 ( .A1(n1322), .A2(n1330), .ZN(n1331) );
NAND3_X1 U1047 ( .A1(G234), .A2(n1049), .A3(G221), .ZN(n1330) );
INV_X1 U1048 ( .A(G137), .ZN(n1322) );
NAND2_X1 U1049 ( .A1(n1332), .A2(n1333), .ZN(n1326) );
OR2_X1 U1050 ( .A1(n1334), .A2(n1275), .ZN(n1333) );
XOR2_X1 U1051 ( .A(n1335), .B(KEYINPUT6), .Z(n1332) );
NAND2_X1 U1052 ( .A1(n1334), .A2(n1275), .ZN(n1335) );
INV_X1 U1053 ( .A(G110), .ZN(n1275) );
XNOR2_X1 U1054 ( .A(n1336), .B(G119), .ZN(n1334) );
NAND2_X1 U1055 ( .A1(KEYINPUT18), .A2(n1337), .ZN(n1336) );
NOR2_X1 U1056 ( .A1(n1238), .A2(n1239), .ZN(n1064) );
NAND2_X1 U1057 ( .A1(n1108), .A2(n1107), .ZN(n1239) );
NAND2_X1 U1058 ( .A1(G475), .A2(n1338), .ZN(n1107) );
INV_X1 U1059 ( .A(n1339), .ZN(n1338) );
NAND2_X1 U1060 ( .A1(n1339), .A2(n1161), .ZN(n1108) );
INV_X1 U1061 ( .A(G475), .ZN(n1161) );
NOR2_X1 U1062 ( .A1(n1160), .A2(G902), .ZN(n1339) );
XNOR2_X1 U1063 ( .A(n1340), .B(n1341), .ZN(n1160) );
XNOR2_X1 U1064 ( .A(n1304), .B(n1342), .ZN(n1341) );
NOR2_X1 U1065 ( .A1(KEYINPUT52), .A2(n1343), .ZN(n1342) );
XNOR2_X1 U1066 ( .A(G122), .B(G113), .ZN(n1343) );
INV_X1 U1067 ( .A(G104), .ZN(n1304) );
NAND2_X1 U1068 ( .A1(KEYINPUT26), .A2(n1344), .ZN(n1340) );
XOR2_X1 U1069 ( .A(n1345), .B(n1346), .Z(n1344) );
XOR2_X1 U1070 ( .A(n1324), .B(n1347), .Z(n1346) );
AND2_X1 U1071 ( .A1(G214), .A2(n1319), .ZN(n1347) );
NOR2_X1 U1072 ( .A1(G953), .A2(G237), .ZN(n1319) );
XNOR2_X1 U1073 ( .A(G125), .B(n1348), .ZN(n1324) );
XNOR2_X1 U1074 ( .A(n1349), .B(G140), .ZN(n1348) );
INV_X1 U1075 ( .A(G146), .ZN(n1349) );
XNOR2_X1 U1076 ( .A(G131), .B(n1350), .ZN(n1345) );
XOR2_X1 U1077 ( .A(KEYINPUT46), .B(G143), .Z(n1350) );
XOR2_X1 U1078 ( .A(n1351), .B(n1156), .Z(n1238) );
INV_X1 U1079 ( .A(G478), .ZN(n1156) );
NAND2_X1 U1080 ( .A1(n1157), .A2(n1268), .ZN(n1351) );
INV_X1 U1081 ( .A(G902), .ZN(n1268) );
NAND2_X1 U1082 ( .A1(n1352), .A2(n1353), .ZN(n1157) );
NAND2_X1 U1083 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NAND3_X1 U1084 ( .A1(G234), .A2(n1049), .A3(G217), .ZN(n1355) );
NAND4_X1 U1085 ( .A1(G234), .A2(n1049), .A3(G217), .A4(n1356), .ZN(n1352) );
INV_X1 U1086 ( .A(n1354), .ZN(n1356) );
XNOR2_X1 U1087 ( .A(n1357), .B(n1358), .ZN(n1354) );
XOR2_X1 U1088 ( .A(n1318), .B(n1359), .Z(n1358) );
XNOR2_X1 U1089 ( .A(G116), .B(n1280), .ZN(n1359) );
INV_X1 U1090 ( .A(G107), .ZN(n1280) );
XNOR2_X1 U1091 ( .A(n1337), .B(G143), .ZN(n1318) );
INV_X1 U1092 ( .A(G128), .ZN(n1337) );
XNOR2_X1 U1093 ( .A(G122), .B(n1360), .ZN(n1357) );
XOR2_X1 U1094 ( .A(KEYINPUT49), .B(G134), .Z(n1360) );
INV_X1 U1095 ( .A(G953), .ZN(n1049) );
endmodule


