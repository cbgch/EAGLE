//Key = 1110011000001010000100111010110110101111101101000101001110110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279;

XNOR2_X1 U709 ( .A(G107), .B(n981), .ZN(G9) );
NOR2_X1 U710 ( .A1(n982), .A2(n983), .ZN(G75) );
NOR3_X1 U711 ( .A1(n984), .A2(n985), .A3(n986), .ZN(n983) );
INV_X1 U712 ( .A(n987), .ZN(n986) );
XOR2_X1 U713 ( .A(n988), .B(KEYINPUT28), .Z(n985) );
NAND3_X1 U714 ( .A1(n989), .A2(n990), .A3(n991), .ZN(n988) );
NAND2_X1 U715 ( .A1(n992), .A2(n993), .ZN(n990) );
NAND3_X1 U716 ( .A1(n994), .A2(n995), .A3(n996), .ZN(n993) );
NAND2_X1 U717 ( .A1(n997), .A2(n998), .ZN(n992) );
NAND3_X1 U718 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n998) );
NAND2_X1 U719 ( .A1(n996), .A2(n1002), .ZN(n1001) );
NAND3_X1 U720 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1000) );
XNOR2_X1 U721 ( .A(KEYINPUT11), .B(n1006), .ZN(n1004) );
NAND3_X1 U722 ( .A1(n995), .A2(n1007), .A3(n1008), .ZN(n999) );
NAND3_X1 U723 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n984) );
NAND2_X1 U724 ( .A1(n991), .A2(n1012), .ZN(n1011) );
NAND2_X1 U725 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND3_X1 U726 ( .A1(n1015), .A2(n1016), .A3(n996), .ZN(n1014) );
NOR2_X1 U727 ( .A1(n1017), .A2(n1005), .ZN(n996) );
NAND3_X1 U728 ( .A1(n1008), .A2(n1018), .A3(n997), .ZN(n1013) );
NAND2_X1 U729 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND3_X1 U730 ( .A1(n1021), .A2(n1015), .A3(n1022), .ZN(n1020) );
NAND3_X1 U731 ( .A1(n1023), .A2(n1024), .A3(n1003), .ZN(n1019) );
NAND2_X1 U732 ( .A1(n989), .A2(n1025), .ZN(n1024) );
NAND2_X1 U733 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U734 ( .A1(n1028), .A2(n1006), .ZN(n1023) );
AND3_X1 U735 ( .A1(n1009), .A2(n1010), .A3(n1029), .ZN(n982) );
NAND4_X1 U736 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1009) );
NOR4_X1 U737 ( .A1(n1034), .A2(n1035), .A3(n1017), .A4(n1006), .ZN(n1033) );
XOR2_X1 U738 ( .A(n1036), .B(KEYINPUT39), .Z(n1035) );
NAND2_X1 U739 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U740 ( .A1(n1037), .A2(n1038), .ZN(n1034) );
XNOR2_X1 U741 ( .A(n1039), .B(n1040), .ZN(n1032) );
XNOR2_X1 U742 ( .A(n1041), .B(n1042), .ZN(n1031) );
XOR2_X1 U743 ( .A(n1043), .B(n1044), .Z(n1030) );
XOR2_X1 U744 ( .A(KEYINPUT18), .B(G472), .Z(n1044) );
XOR2_X1 U745 ( .A(n1045), .B(n1046), .Z(G72) );
XOR2_X1 U746 ( .A(n1047), .B(n1048), .Z(n1046) );
NOR2_X1 U747 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U748 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
XOR2_X1 U749 ( .A(KEYINPUT2), .B(G227), .Z(n1052) );
NAND2_X1 U750 ( .A1(n1053), .A2(n1054), .ZN(n1047) );
NAND2_X1 U751 ( .A1(n1055), .A2(n1051), .ZN(n1054) );
XNOR2_X1 U752 ( .A(KEYINPUT41), .B(n1010), .ZN(n1055) );
XOR2_X1 U753 ( .A(n1056), .B(n1057), .Z(n1053) );
XOR2_X1 U754 ( .A(n1058), .B(n1059), .Z(n1057) );
XOR2_X1 U755 ( .A(n1060), .B(n1061), .Z(n1059) );
XOR2_X1 U756 ( .A(n1062), .B(n1063), .Z(n1056) );
NOR2_X1 U757 ( .A1(KEYINPUT35), .A2(n1064), .ZN(n1063) );
XNOR2_X1 U758 ( .A(KEYINPUT61), .B(KEYINPUT10), .ZN(n1062) );
NAND2_X1 U759 ( .A1(n1010), .A2(n1065), .ZN(n1045) );
XOR2_X1 U760 ( .A(n1066), .B(n1067), .Z(G69) );
XOR2_X1 U761 ( .A(n1068), .B(n1069), .Z(n1067) );
NOR2_X1 U762 ( .A1(n1070), .A2(n1050), .ZN(n1069) );
XNOR2_X1 U763 ( .A(n1010), .B(KEYINPUT38), .ZN(n1050) );
AND2_X1 U764 ( .A1(G224), .A2(G898), .ZN(n1070) );
NAND2_X1 U765 ( .A1(n1071), .A2(n1072), .ZN(n1068) );
NAND2_X1 U766 ( .A1(G953), .A2(n1073), .ZN(n1072) );
XOR2_X1 U767 ( .A(n1074), .B(n1075), .Z(n1071) );
XNOR2_X1 U768 ( .A(n1076), .B(n1077), .ZN(n1075) );
XOR2_X1 U769 ( .A(n1078), .B(n1079), .Z(n1074) );
XNOR2_X1 U770 ( .A(KEYINPUT8), .B(KEYINPUT6), .ZN(n1079) );
NAND2_X1 U771 ( .A1(KEYINPUT29), .A2(n1080), .ZN(n1078) );
NAND2_X1 U772 ( .A1(n1010), .A2(n1081), .ZN(n1066) );
NOR2_X1 U773 ( .A1(n1082), .A2(n1083), .ZN(G66) );
XOR2_X1 U774 ( .A(n1084), .B(n1085), .Z(n1083) );
NAND2_X1 U775 ( .A1(n1086), .A2(n1040), .ZN(n1084) );
NOR2_X1 U776 ( .A1(n1082), .A2(n1087), .ZN(G63) );
NOR3_X1 U777 ( .A1(n1088), .A2(n1037), .A3(n1089), .ZN(n1087) );
NOR4_X1 U778 ( .A1(n1090), .A2(n1091), .A3(n1038), .A4(n1092), .ZN(n1089) );
NOR2_X1 U779 ( .A1(n1093), .A2(n1094), .ZN(n1088) );
NOR2_X1 U780 ( .A1(n1090), .A2(n1091), .ZN(n1094) );
NOR2_X1 U781 ( .A1(n987), .A2(n1038), .ZN(n1093) );
NOR2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(G60) );
XOR2_X1 U783 ( .A(n1097), .B(n1098), .Z(n1096) );
NAND2_X1 U784 ( .A1(n1086), .A2(G475), .ZN(n1097) );
NOR2_X1 U785 ( .A1(n1099), .A2(n1100), .ZN(n1095) );
XNOR2_X1 U786 ( .A(KEYINPUT60), .B(n1029), .ZN(n1100) );
XNOR2_X1 U787 ( .A(KEYINPUT50), .B(G953), .ZN(n1099) );
XNOR2_X1 U788 ( .A(n1101), .B(n1102), .ZN(G6) );
NOR2_X1 U789 ( .A1(KEYINPUT46), .A2(n1103), .ZN(n1102) );
NOR2_X1 U790 ( .A1(n1082), .A2(n1104), .ZN(G57) );
XOR2_X1 U791 ( .A(n1105), .B(n1106), .Z(n1104) );
XNOR2_X1 U792 ( .A(n1107), .B(n1108), .ZN(n1106) );
XOR2_X1 U793 ( .A(n1109), .B(n1110), .Z(n1105) );
NOR2_X1 U794 ( .A1(KEYINPUT57), .A2(n1111), .ZN(n1110) );
XOR2_X1 U795 ( .A(n1112), .B(n1113), .Z(n1111) );
XNOR2_X1 U796 ( .A(G101), .B(KEYINPUT4), .ZN(n1113) );
NAND2_X1 U797 ( .A1(n1086), .A2(G472), .ZN(n1109) );
NOR2_X1 U798 ( .A1(n1082), .A2(n1114), .ZN(G54) );
XOR2_X1 U799 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U800 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U801 ( .A1(KEYINPUT43), .A2(n1119), .ZN(n1118) );
NAND2_X1 U802 ( .A1(n1086), .A2(G469), .ZN(n1117) );
NOR2_X1 U803 ( .A1(n1082), .A2(n1120), .ZN(G51) );
XOR2_X1 U804 ( .A(n1121), .B(n1122), .Z(n1120) );
XNOR2_X1 U805 ( .A(n1123), .B(n1124), .ZN(n1122) );
XNOR2_X1 U806 ( .A(G125), .B(KEYINPUT27), .ZN(n1124) );
XNOR2_X1 U807 ( .A(n1125), .B(n1126), .ZN(n1121) );
XNOR2_X1 U808 ( .A(n1127), .B(n1064), .ZN(n1126) );
NAND3_X1 U809 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1127) );
NAND2_X1 U810 ( .A1(KEYINPUT23), .A2(n1092), .ZN(n1129) );
INV_X1 U811 ( .A(n1086), .ZN(n1092) );
NOR2_X1 U812 ( .A1(n1131), .A2(n987), .ZN(n1086) );
NAND2_X1 U813 ( .A1(n1132), .A2(n1133), .ZN(n1128) );
INV_X1 U814 ( .A(KEYINPUT23), .ZN(n1133) );
NAND2_X1 U815 ( .A1(n987), .A2(G902), .ZN(n1132) );
NOR2_X1 U816 ( .A1(n1081), .A2(n1065), .ZN(n987) );
NAND4_X1 U817 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1065) );
NOR4_X1 U818 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1137) );
INV_X1 U819 ( .A(n1142), .ZN(n1140) );
NOR2_X1 U820 ( .A1(n1143), .A2(n1144), .ZN(n1136) );
NAND3_X1 U821 ( .A1(n1016), .A2(n1007), .A3(n1145), .ZN(n1134) );
NAND4_X1 U822 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1081) );
AND4_X1 U823 ( .A1(n1150), .A2(n1101), .A3(n981), .A4(n1151), .ZN(n1149) );
NAND3_X1 U824 ( .A1(n1016), .A2(n1152), .A3(n1002), .ZN(n981) );
NAND3_X1 U825 ( .A1(n1002), .A2(n1152), .A3(n994), .ZN(n1101) );
NAND2_X1 U826 ( .A1(n1153), .A2(n1016), .ZN(n1148) );
NAND2_X1 U827 ( .A1(n1154), .A2(n1155), .ZN(n1146) );
NAND2_X1 U828 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND3_X1 U829 ( .A1(n995), .A2(n1158), .A3(KEYINPUT15), .ZN(n1157) );
NAND3_X1 U830 ( .A1(n1159), .A2(n1160), .A3(n1028), .ZN(n1156) );
OR2_X1 U831 ( .A1(n1005), .A2(n1002), .ZN(n1160) );
NAND2_X1 U832 ( .A1(n1161), .A2(n1005), .ZN(n1159) );
OR2_X1 U833 ( .A1(n1006), .A2(KEYINPUT15), .ZN(n1161) );
AND2_X1 U834 ( .A1(n1162), .A2(n1029), .ZN(n1082) );
INV_X1 U835 ( .A(G952), .ZN(n1029) );
XNOR2_X1 U836 ( .A(KEYINPUT50), .B(n1010), .ZN(n1162) );
XNOR2_X1 U837 ( .A(n1163), .B(n1139), .ZN(G48) );
AND3_X1 U838 ( .A1(n994), .A2(n1007), .A3(n1145), .ZN(n1139) );
XNOR2_X1 U839 ( .A(G143), .B(n1135), .ZN(G45) );
NAND4_X1 U840 ( .A1(n1164), .A2(n1165), .A3(n1007), .A4(n1166), .ZN(n1135) );
XOR2_X1 U841 ( .A(G140), .B(n1144), .Z(G42) );
AND3_X1 U842 ( .A1(n1003), .A2(n1002), .A3(n1167), .ZN(n1144) );
XOR2_X1 U843 ( .A(G137), .B(n1138), .Z(G39) );
AND3_X1 U844 ( .A1(n997), .A2(n1003), .A3(n1145), .ZN(n1138) );
INV_X1 U845 ( .A(n1168), .ZN(n1145) );
XOR2_X1 U846 ( .A(G134), .B(n1143), .Z(G36) );
AND3_X1 U847 ( .A1(n1003), .A2(n1016), .A3(n1165), .ZN(n1143) );
INV_X1 U848 ( .A(n1169), .ZN(n1016) );
XOR2_X1 U849 ( .A(G131), .B(n1141), .Z(G33) );
AND3_X1 U850 ( .A1(n994), .A2(n1003), .A3(n1165), .ZN(n1141) );
AND4_X1 U851 ( .A1(n1002), .A2(n989), .A3(n1170), .A4(n1005), .ZN(n1165) );
INV_X1 U852 ( .A(n1017), .ZN(n1003) );
NAND2_X1 U853 ( .A1(n1021), .A2(n1171), .ZN(n1017) );
XOR2_X1 U854 ( .A(G128), .B(n1172), .Z(G30) );
NOR3_X1 U855 ( .A1(n1168), .A2(n1173), .A3(n1169), .ZN(n1172) );
XNOR2_X1 U856 ( .A(n1007), .B(KEYINPUT3), .ZN(n1173) );
NAND3_X1 U857 ( .A1(n1002), .A2(n1170), .A3(n1174), .ZN(n1168) );
XNOR2_X1 U858 ( .A(n1175), .B(n1176), .ZN(G3) );
NOR2_X1 U859 ( .A1(n1177), .A2(n1151), .ZN(n1176) );
NAND4_X1 U860 ( .A1(n1154), .A2(n1002), .A3(n989), .A4(n1005), .ZN(n1151) );
XNOR2_X1 U861 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n1177) );
XNOR2_X1 U862 ( .A(n1178), .B(n1179), .ZN(G27) );
NOR2_X1 U863 ( .A1(KEYINPUT48), .A2(n1142), .ZN(n1179) );
NAND3_X1 U864 ( .A1(n995), .A2(n1007), .A3(n1167), .ZN(n1142) );
AND4_X1 U865 ( .A1(n1028), .A2(n994), .A3(n1008), .A4(n1170), .ZN(n1167) );
NAND2_X1 U866 ( .A1(n1180), .A2(n1181), .ZN(n1170) );
NAND4_X1 U867 ( .A1(n1182), .A2(G902), .A3(G953), .A4(n1051), .ZN(n1181) );
INV_X1 U868 ( .A(G900), .ZN(n1051) );
XOR2_X1 U869 ( .A(n1183), .B(KEYINPUT25), .Z(n1182) );
XNOR2_X1 U870 ( .A(G122), .B(n1150), .ZN(G24) );
NAND4_X1 U871 ( .A1(n1164), .A2(n995), .A3(n1152), .A4(n1166), .ZN(n1150) );
AND3_X1 U872 ( .A1(n1008), .A2(n989), .A3(n1184), .ZN(n1152) );
INV_X1 U873 ( .A(n1006), .ZN(n995) );
XOR2_X1 U874 ( .A(G119), .B(n1185), .Z(G21) );
NOR4_X1 U875 ( .A1(KEYINPUT9), .A2(n1006), .A3(n1186), .A4(n1158), .ZN(n1185) );
INV_X1 U876 ( .A(n1174), .ZN(n1158) );
NOR2_X1 U877 ( .A1(n989), .A2(n1008), .ZN(n1174) );
XNOR2_X1 U878 ( .A(n1187), .B(n1188), .ZN(G18) );
NOR3_X1 U879 ( .A1(n1189), .A2(n1169), .A3(n1190), .ZN(n1188) );
NAND2_X1 U880 ( .A1(n1191), .A2(n1166), .ZN(n1169) );
XOR2_X1 U881 ( .A(KEYINPUT37), .B(KEYINPUT32), .Z(n1189) );
XNOR2_X1 U882 ( .A(n1147), .B(n1192), .ZN(G15) );
NOR2_X1 U883 ( .A1(KEYINPUT33), .A2(n1193), .ZN(n1192) );
NAND2_X1 U884 ( .A1(n1153), .A2(n994), .ZN(n1147) );
NOR2_X1 U885 ( .A1(n1166), .A2(n1191), .ZN(n994) );
INV_X1 U886 ( .A(n1190), .ZN(n1153) );
NAND3_X1 U887 ( .A1(n1184), .A2(n1005), .A3(n1015), .ZN(n1190) );
NOR2_X1 U888 ( .A1(n1006), .A2(n1028), .ZN(n1015) );
NAND2_X1 U889 ( .A1(n1027), .A2(n1194), .ZN(n1006) );
XNOR2_X1 U890 ( .A(G110), .B(n1195), .ZN(G12) );
NAND4_X1 U891 ( .A1(n1028), .A2(n1154), .A3(n1008), .A4(n1196), .ZN(n1195) );
XOR2_X1 U892 ( .A(KEYINPUT44), .B(n1002), .Z(n1196) );
NOR2_X1 U893 ( .A1(n1027), .A2(n1026), .ZN(n1002) );
INV_X1 U894 ( .A(n1194), .ZN(n1026) );
NAND2_X1 U895 ( .A1(G221), .A2(n1197), .ZN(n1194) );
XOR2_X1 U896 ( .A(n1198), .B(G469), .Z(n1027) );
NAND2_X1 U897 ( .A1(n1199), .A2(n1131), .ZN(n1198) );
XOR2_X1 U898 ( .A(n1200), .B(n1201), .Z(n1199) );
XNOR2_X1 U899 ( .A(n1115), .B(G110), .ZN(n1201) );
XNOR2_X1 U900 ( .A(n1202), .B(n1203), .ZN(n1115) );
XOR2_X1 U901 ( .A(n1204), .B(n1108), .Z(n1203) );
XNOR2_X1 U902 ( .A(n1064), .B(n1205), .ZN(n1108) );
XNOR2_X1 U903 ( .A(n1060), .B(n1206), .ZN(n1202) );
XNOR2_X1 U904 ( .A(n1175), .B(n1207), .ZN(n1206) );
AND2_X1 U905 ( .A1(n1010), .A2(G227), .ZN(n1207) );
INV_X1 U906 ( .A(G101), .ZN(n1175) );
XNOR2_X1 U907 ( .A(KEYINPUT7), .B(KEYINPUT52), .ZN(n1200) );
INV_X1 U908 ( .A(n1005), .ZN(n1008) );
NAND2_X1 U909 ( .A1(n1208), .A2(n1209), .ZN(n1005) );
NAND2_X1 U910 ( .A1(G472), .A2(n1043), .ZN(n1209) );
XOR2_X1 U911 ( .A(KEYINPUT54), .B(n1210), .Z(n1208) );
NOR2_X1 U912 ( .A1(G472), .A2(n1043), .ZN(n1210) );
NAND2_X1 U913 ( .A1(n1211), .A2(n1131), .ZN(n1043) );
XOR2_X1 U914 ( .A(n1212), .B(n1213), .Z(n1211) );
XNOR2_X1 U915 ( .A(n1214), .B(n1215), .ZN(n1213) );
INV_X1 U916 ( .A(n1107), .ZN(n1215) );
XNOR2_X1 U917 ( .A(n1080), .B(KEYINPUT0), .ZN(n1107) );
NAND2_X1 U918 ( .A1(n1216), .A2(KEYINPUT63), .ZN(n1214) );
XOR2_X1 U919 ( .A(n1217), .B(n1218), .Z(n1216) );
NOR2_X1 U920 ( .A1(KEYINPUT53), .A2(n1112), .ZN(n1218) );
NAND2_X1 U921 ( .A1(G210), .A2(n1219), .ZN(n1112) );
XNOR2_X1 U922 ( .A(G101), .B(KEYINPUT34), .ZN(n1217) );
XOR2_X1 U923 ( .A(n1220), .B(KEYINPUT59), .Z(n1212) );
NAND2_X1 U924 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NAND2_X1 U925 ( .A1(n1205), .A2(n1064), .ZN(n1222) );
XOR2_X1 U926 ( .A(KEYINPUT62), .B(n1223), .Z(n1221) );
NOR2_X1 U927 ( .A1(n1205), .A2(n1064), .ZN(n1223) );
XOR2_X1 U928 ( .A(n1058), .B(n1224), .Z(n1205) );
NOR2_X1 U929 ( .A1(G137), .A2(KEYINPUT30), .ZN(n1224) );
XNOR2_X1 U930 ( .A(G131), .B(G134), .ZN(n1058) );
INV_X1 U931 ( .A(n1186), .ZN(n1154) );
NAND2_X1 U932 ( .A1(n997), .A2(n1184), .ZN(n1186) );
AND2_X1 U933 ( .A1(n1007), .A2(n1225), .ZN(n1184) );
NAND2_X1 U934 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
NAND4_X1 U935 ( .A1(G902), .A2(G953), .A3(n1183), .A4(n1073), .ZN(n1227) );
INV_X1 U936 ( .A(G898), .ZN(n1073) );
XNOR2_X1 U937 ( .A(n991), .B(KEYINPUT47), .ZN(n1226) );
INV_X1 U938 ( .A(n1180), .ZN(n991) );
NAND3_X1 U939 ( .A1(n1183), .A2(n1010), .A3(G952), .ZN(n1180) );
NAND2_X1 U940 ( .A1(G237), .A2(G234), .ZN(n1183) );
NOR2_X1 U941 ( .A1(n1021), .A2(n1022), .ZN(n1007) );
INV_X1 U942 ( .A(n1171), .ZN(n1022) );
NAND2_X1 U943 ( .A1(G214), .A2(n1228), .ZN(n1171) );
XOR2_X1 U944 ( .A(n1229), .B(n1130), .Z(n1021) );
AND2_X1 U945 ( .A1(G210), .A2(n1228), .ZN(n1130) );
NAND2_X1 U946 ( .A1(n1230), .A2(n1131), .ZN(n1228) );
INV_X1 U947 ( .A(G237), .ZN(n1230) );
NAND2_X1 U948 ( .A1(n1231), .A2(n1131), .ZN(n1229) );
XOR2_X1 U949 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U950 ( .A(n1234), .B(n1235), .Z(n1233) );
NAND2_X1 U951 ( .A1(KEYINPUT49), .A2(n1123), .ZN(n1235) );
AND2_X1 U952 ( .A1(G224), .A2(n1236), .ZN(n1123) );
XNOR2_X1 U953 ( .A(KEYINPUT12), .B(n1010), .ZN(n1236) );
NAND2_X1 U954 ( .A1(n1237), .A2(n1238), .ZN(n1234) );
NAND2_X1 U955 ( .A1(n1064), .A2(n1178), .ZN(n1238) );
XOR2_X1 U956 ( .A(KEYINPUT26), .B(n1239), .Z(n1237) );
NOR2_X1 U957 ( .A1(n1064), .A2(n1178), .ZN(n1239) );
INV_X1 U958 ( .A(G125), .ZN(n1178) );
XOR2_X1 U959 ( .A(G146), .B(n1240), .Z(n1064) );
NAND2_X1 U960 ( .A1(KEYINPUT56), .A2(n1125), .ZN(n1232) );
XOR2_X1 U961 ( .A(n1241), .B(n1242), .Z(n1125) );
INV_X1 U962 ( .A(n1076), .ZN(n1242) );
XNOR2_X1 U963 ( .A(n1243), .B(n1204), .ZN(n1076) );
XNOR2_X1 U964 ( .A(n1103), .B(G107), .ZN(n1204) );
NAND2_X1 U965 ( .A1(KEYINPUT45), .A2(G101), .ZN(n1243) );
XNOR2_X1 U966 ( .A(n1244), .B(n1080), .ZN(n1241) );
XNOR2_X1 U967 ( .A(G113), .B(n1245), .ZN(n1080) );
XNOR2_X1 U968 ( .A(G119), .B(n1187), .ZN(n1245) );
NAND2_X1 U969 ( .A1(KEYINPUT5), .A2(n1077), .ZN(n1244) );
XOR2_X1 U970 ( .A(n1246), .B(n1247), .Z(n1077) );
NAND2_X1 U971 ( .A1(KEYINPUT42), .A2(n1119), .ZN(n1246) );
NOR2_X1 U972 ( .A1(n1166), .A2(n1164), .ZN(n997) );
INV_X1 U973 ( .A(n1191), .ZN(n1164) );
XOR2_X1 U974 ( .A(n1248), .B(n1041), .Z(n1191) );
NAND2_X1 U975 ( .A1(n1098), .A2(n1131), .ZN(n1041) );
XNOR2_X1 U976 ( .A(n1249), .B(n1250), .ZN(n1098) );
XNOR2_X1 U977 ( .A(n1247), .B(n1251), .ZN(n1250) );
XOR2_X1 U978 ( .A(n1252), .B(n1253), .Z(n1251) );
NOR2_X1 U979 ( .A1(G131), .A2(KEYINPUT21), .ZN(n1253) );
NAND2_X1 U980 ( .A1(G214), .A2(n1219), .ZN(n1252) );
NOR2_X1 U981 ( .A1(G953), .A2(G237), .ZN(n1219) );
XOR2_X1 U982 ( .A(n1254), .B(n1255), .Z(n1249) );
XNOR2_X1 U983 ( .A(G143), .B(n1193), .ZN(n1255) );
INV_X1 U984 ( .A(G113), .ZN(n1193) );
XNOR2_X1 U985 ( .A(n1256), .B(n1103), .ZN(n1254) );
INV_X1 U986 ( .A(G104), .ZN(n1103) );
NAND2_X1 U987 ( .A1(n1257), .A2(KEYINPUT51), .ZN(n1256) );
XNOR2_X1 U988 ( .A(n1258), .B(n1163), .ZN(n1257) );
NAND2_X1 U989 ( .A1(n1259), .A2(KEYINPUT14), .ZN(n1258) );
XNOR2_X1 U990 ( .A(G125), .B(n1060), .ZN(n1259) );
NAND2_X1 U991 ( .A1(KEYINPUT40), .A2(n1042), .ZN(n1248) );
INV_X1 U992 ( .A(G475), .ZN(n1042) );
XOR2_X1 U993 ( .A(n1037), .B(n1260), .Z(n1166) );
XNOR2_X1 U994 ( .A(KEYINPUT13), .B(n1038), .ZN(n1260) );
INV_X1 U995 ( .A(G478), .ZN(n1038) );
AND2_X1 U996 ( .A1(n1261), .A2(n1131), .ZN(n1037) );
OR2_X1 U997 ( .A1(n1090), .A2(n1091), .ZN(n1261) );
NOR2_X1 U998 ( .A1(n1262), .A2(n1263), .ZN(n1091) );
AND2_X1 U999 ( .A1(n1263), .A2(n1262), .ZN(n1090) );
NAND3_X1 U1000 ( .A1(G234), .A2(n1264), .A3(G217), .ZN(n1262) );
XNOR2_X1 U1001 ( .A(KEYINPUT36), .B(n1010), .ZN(n1264) );
XNOR2_X1 U1002 ( .A(n1265), .B(n1266), .ZN(n1263) );
XOR2_X1 U1003 ( .A(G107), .B(n1267), .Z(n1266) );
XOR2_X1 U1004 ( .A(KEYINPUT31), .B(G134), .Z(n1267) );
XOR2_X1 U1005 ( .A(n1268), .B(n1247), .Z(n1265) );
XOR2_X1 U1006 ( .A(G122), .B(KEYINPUT16), .Z(n1247) );
XOR2_X1 U1007 ( .A(n1269), .B(n1240), .Z(n1268) );
XOR2_X1 U1008 ( .A(G128), .B(G143), .Z(n1240) );
NAND2_X1 U1009 ( .A1(KEYINPUT58), .A2(n1187), .ZN(n1269) );
INV_X1 U1010 ( .A(G116), .ZN(n1187) );
INV_X1 U1011 ( .A(n989), .ZN(n1028) );
XOR2_X1 U1012 ( .A(n1040), .B(n1270), .Z(n989) );
NOR2_X1 U1013 ( .A1(n1039), .A2(KEYINPUT20), .ZN(n1270) );
AND2_X1 U1014 ( .A1(n1271), .A2(n1131), .ZN(n1039) );
XNOR2_X1 U1015 ( .A(n1085), .B(KEYINPUT24), .ZN(n1271) );
XNOR2_X1 U1016 ( .A(n1272), .B(n1273), .ZN(n1085) );
XOR2_X1 U1017 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U1018 ( .A(G128), .B(G119), .Z(n1275) );
XNOR2_X1 U1019 ( .A(KEYINPUT55), .B(n1163), .ZN(n1274) );
INV_X1 U1020 ( .A(G146), .ZN(n1163) );
XOR2_X1 U1021 ( .A(n1276), .B(n1277), .Z(n1272) );
XOR2_X1 U1022 ( .A(n1278), .B(n1061), .Z(n1277) );
XOR2_X1 U1023 ( .A(G137), .B(G125), .Z(n1061) );
AND3_X1 U1024 ( .A1(G221), .A2(n1010), .A3(G234), .ZN(n1278) );
INV_X1 U1025 ( .A(G953), .ZN(n1010) );
XNOR2_X1 U1026 ( .A(n1279), .B(n1119), .ZN(n1276) );
INV_X1 U1027 ( .A(G110), .ZN(n1119) );
NAND2_X1 U1028 ( .A1(KEYINPUT22), .A2(n1060), .ZN(n1279) );
XOR2_X1 U1029 ( .A(G140), .B(KEYINPUT1), .Z(n1060) );
AND2_X1 U1030 ( .A1(G217), .A2(n1197), .ZN(n1040) );
NAND2_X1 U1031 ( .A1(G234), .A2(n1131), .ZN(n1197) );
INV_X1 U1032 ( .A(G902), .ZN(n1131) );
endmodule


