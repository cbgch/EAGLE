//Key = 0100101111010101110001100010011001010011110001010100110100111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382;

XOR2_X1 U747 ( .A(n1037), .B(n1038), .Z(G9) );
NAND2_X1 U748 ( .A1(KEYINPUT58), .A2(G107), .ZN(n1038) );
NAND2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
XOR2_X1 U750 ( .A(KEYINPUT3), .B(n1041), .Z(n1040) );
NOR2_X1 U751 ( .A1(n1042), .A2(n1043), .ZN(G75) );
NOR3_X1 U752 ( .A1(n1044), .A2(G953), .A3(n1045), .ZN(n1043) );
XNOR2_X1 U753 ( .A(KEYINPUT54), .B(n1046), .ZN(n1044) );
NOR4_X1 U754 ( .A1(n1047), .A2(n1048), .A3(n1045), .A4(n1046), .ZN(n1042) );
INV_X1 U755 ( .A(G952), .ZN(n1046) );
AND4_X1 U756 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1045) );
NOR4_X1 U757 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
XNOR2_X1 U758 ( .A(G475), .B(n1057), .ZN(n1056) );
XOR2_X1 U759 ( .A(n1058), .B(n1059), .Z(n1053) );
NOR2_X1 U760 ( .A1(KEYINPUT37), .A2(n1060), .ZN(n1059) );
XOR2_X1 U761 ( .A(KEYINPUT51), .B(G469), .Z(n1060) );
AND2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(n1051) );
XNOR2_X1 U763 ( .A(G472), .B(n1063), .ZN(n1049) );
NAND2_X1 U764 ( .A1(n1064), .A2(KEYINPUT29), .ZN(n1063) );
XOR2_X1 U765 ( .A(n1065), .B(KEYINPUT20), .Z(n1064) );
NAND4_X1 U766 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1047) );
NAND2_X1 U767 ( .A1(n1070), .A2(n1039), .ZN(n1068) );
NAND3_X1 U768 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1067) );
XNOR2_X1 U769 ( .A(n1070), .B(KEYINPUT61), .ZN(n1073) );
AND3_X1 U770 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1070) );
NAND2_X1 U771 ( .A1(n1077), .A2(n1078), .ZN(n1066) );
NAND2_X1 U772 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U773 ( .A1(n1081), .A2(n1075), .ZN(n1080) );
NAND2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U775 ( .A1(n1074), .A2(n1084), .ZN(n1083) );
NAND2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U778 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U780 ( .A1(n1093), .A2(n1094), .ZN(n1085) );
OR2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U782 ( .A1(n1076), .A2(n1097), .ZN(n1082) );
NAND2_X1 U783 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U784 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
INV_X1 U785 ( .A(KEYINPUT44), .ZN(n1101) );
NAND2_X1 U786 ( .A1(KEYINPUT44), .A2(n1102), .ZN(n1079) );
NAND3_X1 U787 ( .A1(n1076), .A2(n1075), .A3(n1100), .ZN(n1102) );
XOR2_X1 U788 ( .A(n1103), .B(n1104), .Z(G72) );
NAND2_X1 U789 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U790 ( .A1(n1107), .A2(n1069), .ZN(n1106) );
XOR2_X1 U791 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND3_X1 U792 ( .A1(G900), .A2(n1109), .A3(G953), .ZN(n1105) );
XNOR2_X1 U793 ( .A(n1110), .B(n1111), .ZN(n1109) );
NAND3_X1 U794 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1110) );
NAND2_X1 U795 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
OR3_X1 U796 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1113) );
INV_X1 U797 ( .A(KEYINPUT41), .ZN(n1116) );
NAND2_X1 U798 ( .A1(n1118), .A2(n1117), .ZN(n1112) );
NAND2_X1 U799 ( .A1(KEYINPUT45), .A2(n1119), .ZN(n1117) );
NAND2_X1 U800 ( .A1(KEYINPUT55), .A2(n1120), .ZN(n1103) );
NAND2_X1 U801 ( .A1(G953), .A2(n1121), .ZN(n1120) );
NAND2_X1 U802 ( .A1(G900), .A2(G227), .ZN(n1121) );
NAND2_X1 U803 ( .A1(n1122), .A2(n1123), .ZN(G69) );
NAND2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND3_X1 U805 ( .A1(G953), .A2(n1126), .A3(n1127), .ZN(n1125) );
XNOR2_X1 U806 ( .A(G224), .B(KEYINPUT57), .ZN(n1127) );
NAND4_X1 U807 ( .A1(n1128), .A2(n1126), .A3(G953), .A4(n1129), .ZN(n1122) );
INV_X1 U808 ( .A(n1124), .ZN(n1129) );
XNOR2_X1 U809 ( .A(n1130), .B(n1131), .ZN(n1124) );
NOR2_X1 U810 ( .A1(n1132), .A2(G953), .ZN(n1131) );
NOR2_X1 U811 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XNOR2_X1 U812 ( .A(n1135), .B(KEYINPUT21), .ZN(n1133) );
NAND3_X1 U813 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1130) );
XOR2_X1 U814 ( .A(n1139), .B(KEYINPUT14), .Z(n1138) );
NAND2_X1 U815 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
INV_X1 U816 ( .A(n1142), .ZN(n1141) );
XNOR2_X1 U817 ( .A(n1143), .B(n1144), .ZN(n1140) );
INV_X1 U818 ( .A(n1145), .ZN(n1137) );
NAND2_X1 U819 ( .A1(n1146), .A2(n1142), .ZN(n1136) );
XNOR2_X1 U820 ( .A(n1143), .B(n1147), .ZN(n1146) );
INV_X1 U821 ( .A(KEYINPUT36), .ZN(n1126) );
NAND2_X1 U822 ( .A1(G898), .A2(n1148), .ZN(n1128) );
XNOR2_X1 U823 ( .A(KEYINPUT57), .B(n1149), .ZN(n1148) );
NOR2_X1 U824 ( .A1(n1150), .A2(n1151), .ZN(G66) );
XOR2_X1 U825 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U826 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NOR2_X1 U827 ( .A1(n1150), .A2(n1156), .ZN(G63) );
XOR2_X1 U828 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U829 ( .A1(n1154), .A2(G478), .ZN(n1158) );
NAND2_X1 U830 ( .A1(n1159), .A2(KEYINPUT7), .ZN(n1157) );
XOR2_X1 U831 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U832 ( .A1(n1150), .A2(n1162), .ZN(G60) );
XOR2_X1 U833 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U834 ( .A1(n1165), .A2(KEYINPUT12), .ZN(n1163) );
AND2_X1 U835 ( .A1(G475), .A2(n1154), .ZN(n1165) );
XNOR2_X1 U836 ( .A(G104), .B(n1166), .ZN(G6) );
NOR2_X1 U837 ( .A1(n1150), .A2(n1167), .ZN(G57) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U839 ( .A(n1170), .B(n1171), .Z(n1168) );
AND3_X1 U840 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1171) );
OR2_X1 U841 ( .A1(n1147), .A2(n1175), .ZN(n1172) );
XOR2_X1 U842 ( .A(n1176), .B(KEYINPUT16), .Z(n1175) );
NAND2_X1 U843 ( .A1(n1154), .A2(G472), .ZN(n1170) );
NOR2_X1 U844 ( .A1(n1150), .A2(n1177), .ZN(G54) );
XOR2_X1 U845 ( .A(n1178), .B(n1179), .Z(n1177) );
NAND2_X1 U846 ( .A1(n1154), .A2(G469), .ZN(n1179) );
NAND2_X1 U847 ( .A1(n1180), .A2(n1181), .ZN(n1178) );
NAND2_X1 U848 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
XOR2_X1 U849 ( .A(KEYINPUT47), .B(n1184), .Z(n1180) );
NOR2_X1 U850 ( .A1(n1182), .A2(n1183), .ZN(n1184) );
XNOR2_X1 U851 ( .A(n1185), .B(KEYINPUT33), .ZN(n1183) );
AND2_X1 U852 ( .A1(n1186), .A2(n1187), .ZN(n1182) );
NAND3_X1 U853 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
INV_X1 U854 ( .A(n1191), .ZN(n1190) );
NAND2_X1 U855 ( .A1(n1192), .A2(n1193), .ZN(n1189) );
NAND2_X1 U856 ( .A1(G140), .A2(n1194), .ZN(n1192) );
NAND2_X1 U857 ( .A1(KEYINPUT1), .A2(n1195), .ZN(n1188) );
XOR2_X1 U858 ( .A(n1196), .B(KEYINPUT18), .Z(n1186) );
NAND3_X1 U859 ( .A1(n1197), .A2(n1198), .A3(n1191), .ZN(n1196) );
OR2_X1 U860 ( .A1(n1193), .A2(n1195), .ZN(n1198) );
NAND3_X1 U861 ( .A1(G140), .A2(n1194), .A3(n1193), .ZN(n1197) );
INV_X1 U862 ( .A(KEYINPUT1), .ZN(n1193) );
NOR2_X1 U863 ( .A1(n1150), .A2(n1199), .ZN(G51) );
XOR2_X1 U864 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U865 ( .A(n1202), .B(n1203), .Z(n1201) );
NAND2_X1 U866 ( .A1(n1154), .A2(n1204), .ZN(n1203) );
AND2_X1 U867 ( .A1(G902), .A2(n1048), .ZN(n1154) );
OR3_X1 U868 ( .A1(n1134), .A2(n1135), .A3(n1108), .ZN(n1048) );
NAND4_X1 U869 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1108) );
NOR3_X1 U870 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1208) );
INV_X1 U871 ( .A(n1212), .ZN(n1210) );
NAND2_X1 U872 ( .A1(n1077), .A2(n1213), .ZN(n1207) );
NAND2_X1 U873 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND2_X1 U874 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U875 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NAND2_X1 U876 ( .A1(n1220), .A2(n1095), .ZN(n1219) );
XNOR2_X1 U877 ( .A(n1221), .B(KEYINPUT30), .ZN(n1220) );
NAND2_X1 U878 ( .A1(n1096), .A2(n1100), .ZN(n1218) );
XOR2_X1 U879 ( .A(n1222), .B(KEYINPUT0), .Z(n1214) );
NAND3_X1 U880 ( .A1(n1100), .A2(n1223), .A3(n1224), .ZN(n1205) );
INV_X1 U881 ( .A(n1225), .ZN(n1135) );
NAND4_X1 U882 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1134) );
AND4_X1 U883 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1166), .ZN(n1229) );
NAND4_X1 U884 ( .A1(n1233), .A2(n1100), .A3(n1234), .A4(n1087), .ZN(n1166) );
NAND2_X1 U885 ( .A1(n1039), .A2(n1041), .ZN(n1228) );
AND4_X1 U886 ( .A1(n1234), .A2(n1221), .A3(n1087), .A4(n1235), .ZN(n1041) );
NAND3_X1 U887 ( .A1(n1236), .A2(n1234), .A3(n1096), .ZN(n1227) );
NAND2_X1 U888 ( .A1(n1237), .A2(n1233), .ZN(n1226) );
INV_X1 U889 ( .A(n1238), .ZN(n1237) );
NAND2_X1 U890 ( .A1(KEYINPUT63), .A2(n1239), .ZN(n1202) );
XNOR2_X1 U891 ( .A(n1240), .B(n1241), .ZN(n1200) );
NOR2_X1 U892 ( .A1(n1069), .A2(G952), .ZN(n1150) );
XNOR2_X1 U893 ( .A(G146), .B(n1242), .ZN(G48) );
NAND4_X1 U894 ( .A1(KEYINPUT9), .A2(n1224), .A3(n1100), .A4(n1223), .ZN(n1242) );
NAND2_X1 U895 ( .A1(n1243), .A2(n1244), .ZN(G45) );
OR2_X1 U896 ( .A1(n1206), .A2(G143), .ZN(n1244) );
XOR2_X1 U897 ( .A(n1245), .B(KEYINPUT25), .Z(n1243) );
NAND2_X1 U898 ( .A1(G143), .A2(n1206), .ZN(n1245) );
NAND4_X1 U899 ( .A1(n1246), .A2(n1224), .A3(n1095), .A4(n1054), .ZN(n1206) );
NAND3_X1 U900 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(G42) );
NAND2_X1 U901 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
INV_X1 U902 ( .A(KEYINPUT40), .ZN(n1251) );
NAND2_X1 U903 ( .A1(G140), .A2(n1252), .ZN(n1250) );
NAND3_X1 U904 ( .A1(KEYINPUT40), .A2(n1253), .A3(G140), .ZN(n1248) );
NAND2_X1 U905 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND3_X1 U906 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1247) );
XOR2_X1 U907 ( .A(KEYINPUT38), .B(KEYINPUT34), .Z(n1255) );
INV_X1 U908 ( .A(n1252), .ZN(n1254) );
NAND4_X1 U909 ( .A1(n1257), .A2(n1216), .A3(n1096), .A4(n1100), .ZN(n1252) );
XNOR2_X1 U910 ( .A(n1077), .B(KEYINPUT53), .ZN(n1257) );
XOR2_X1 U911 ( .A(G137), .B(n1209), .Z(G39) );
AND4_X1 U912 ( .A1(n1216), .A2(n1077), .A3(n1223), .A4(n1074), .ZN(n1209) );
XNOR2_X1 U913 ( .A(G134), .B(n1258), .ZN(G36) );
NAND4_X1 U914 ( .A1(n1216), .A2(n1077), .A3(n1221), .A4(n1095), .ZN(n1258) );
INV_X1 U915 ( .A(n1055), .ZN(n1077) );
XNOR2_X1 U916 ( .A(n1259), .B(n1260), .ZN(G33) );
NOR2_X1 U917 ( .A1(n1055), .A2(n1222), .ZN(n1260) );
NAND3_X1 U918 ( .A1(n1100), .A2(n1095), .A3(n1216), .ZN(n1222) );
NAND2_X1 U919 ( .A1(n1071), .A2(n1261), .ZN(n1055) );
XNOR2_X1 U920 ( .A(n1262), .B(n1211), .ZN(G30) );
AND3_X1 U921 ( .A1(n1223), .A2(n1221), .A3(n1224), .ZN(n1211) );
AND2_X1 U922 ( .A1(n1216), .A2(n1039), .ZN(n1224) );
NOR2_X1 U923 ( .A1(n1089), .A2(n1263), .ZN(n1216) );
INV_X1 U924 ( .A(n1234), .ZN(n1089) );
XNOR2_X1 U925 ( .A(G101), .B(n1232), .ZN(G3) );
NAND3_X1 U926 ( .A1(n1234), .A2(n1095), .A3(n1236), .ZN(n1232) );
NAND2_X1 U927 ( .A1(n1264), .A2(n1265), .ZN(G27) );
OR2_X1 U928 ( .A1(n1212), .A2(G125), .ZN(n1265) );
XOR2_X1 U929 ( .A(n1266), .B(KEYINPUT2), .Z(n1264) );
NAND2_X1 U930 ( .A1(G125), .A2(n1212), .ZN(n1266) );
NAND4_X1 U931 ( .A1(n1096), .A2(n1100), .A3(n1267), .A4(n1093), .ZN(n1212) );
NOR2_X1 U932 ( .A1(n1263), .A2(n1268), .ZN(n1267) );
AND2_X1 U933 ( .A1(n1269), .A2(n1270), .ZN(n1263) );
NAND4_X1 U934 ( .A1(G902), .A2(G953), .A3(n1075), .A4(n1271), .ZN(n1270) );
INV_X1 U935 ( .A(G900), .ZN(n1271) );
XNOR2_X1 U936 ( .A(KEYINPUT52), .B(n1272), .ZN(n1269) );
XOR2_X1 U937 ( .A(G122), .B(n1273), .Z(G24) );
NOR3_X1 U938 ( .A1(n1238), .A2(n1274), .A3(n1268), .ZN(n1273) );
INV_X1 U939 ( .A(n1039), .ZN(n1268) );
XOR2_X1 U940 ( .A(n1235), .B(KEYINPUT8), .Z(n1274) );
NAND3_X1 U941 ( .A1(n1246), .A2(n1054), .A3(n1076), .ZN(n1238) );
AND2_X1 U942 ( .A1(n1093), .A2(n1087), .ZN(n1076) );
AND2_X1 U943 ( .A1(n1275), .A2(n1276), .ZN(n1087) );
XNOR2_X1 U944 ( .A(KEYINPUT23), .B(n1277), .ZN(n1276) );
XOR2_X1 U945 ( .A(G119), .B(n1278), .Z(G21) );
NOR3_X1 U946 ( .A1(KEYINPUT43), .A2(n1279), .A3(n1280), .ZN(n1278) );
NOR2_X1 U947 ( .A1(KEYINPUT6), .A2(n1281), .ZN(n1280) );
NOR3_X1 U948 ( .A1(n1282), .A2(n1093), .A3(n1283), .ZN(n1281) );
INV_X1 U949 ( .A(n1223), .ZN(n1283) );
AND2_X1 U950 ( .A1(n1225), .A2(KEYINPUT6), .ZN(n1279) );
NAND3_X1 U951 ( .A1(n1223), .A2(n1093), .A3(n1236), .ZN(n1225) );
XNOR2_X1 U952 ( .A(G116), .B(n1231), .ZN(G18) );
NAND2_X1 U953 ( .A1(n1284), .A2(n1221), .ZN(n1231) );
INV_X1 U954 ( .A(n1098), .ZN(n1221) );
NAND2_X1 U955 ( .A1(n1285), .A2(n1054), .ZN(n1098) );
XNOR2_X1 U956 ( .A(KEYINPUT27), .B(n1246), .ZN(n1285) );
XOR2_X1 U957 ( .A(n1230), .B(n1286), .Z(G15) );
XNOR2_X1 U958 ( .A(KEYINPUT39), .B(n1287), .ZN(n1286) );
NAND2_X1 U959 ( .A1(n1284), .A2(n1100), .ZN(n1230) );
NOR2_X1 U960 ( .A1(n1054), .A2(n1288), .ZN(n1100) );
AND3_X1 U961 ( .A1(n1093), .A2(n1095), .A3(n1233), .ZN(n1284) );
NAND2_X1 U962 ( .A1(n1289), .A2(n1290), .ZN(n1095) );
OR3_X1 U963 ( .A1(n1277), .A2(n1275), .A3(KEYINPUT23), .ZN(n1290) );
NAND2_X1 U964 ( .A1(KEYINPUT23), .A2(n1223), .ZN(n1289) );
NOR2_X1 U965 ( .A1(n1275), .A2(n1291), .ZN(n1223) );
INV_X1 U966 ( .A(n1292), .ZN(n1275) );
NOR2_X1 U967 ( .A1(n1293), .A2(n1091), .ZN(n1093) );
XOR2_X1 U968 ( .A(n1294), .B(n1295), .Z(G12) );
XNOR2_X1 U969 ( .A(G110), .B(KEYINPUT48), .ZN(n1295) );
NAND4_X1 U970 ( .A1(KEYINPUT11), .A2(n1096), .A3(n1236), .A4(n1234), .ZN(n1294) );
NOR2_X1 U971 ( .A1(n1092), .A2(n1091), .ZN(n1234) );
INV_X1 U972 ( .A(n1050), .ZN(n1091) );
NAND2_X1 U973 ( .A1(G221), .A2(n1296), .ZN(n1050) );
INV_X1 U974 ( .A(n1293), .ZN(n1092) );
XNOR2_X1 U975 ( .A(n1058), .B(G469), .ZN(n1293) );
NAND3_X1 U976 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1058) );
NAND2_X1 U977 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
INV_X1 U978 ( .A(KEYINPUT19), .ZN(n1301) );
XNOR2_X1 U979 ( .A(n1302), .B(n1185), .ZN(n1300) );
NAND2_X1 U980 ( .A1(KEYINPUT19), .A2(n1303), .ZN(n1297) );
NAND2_X1 U981 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND3_X1 U982 ( .A1(KEYINPUT50), .A2(n1306), .A3(n1185), .ZN(n1305) );
INV_X1 U983 ( .A(n1307), .ZN(n1185) );
NAND2_X1 U984 ( .A1(n1302), .A2(n1307), .ZN(n1304) );
XOR2_X1 U985 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U986 ( .A(n1176), .B(n1310), .Z(n1308) );
NOR2_X1 U987 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U988 ( .A(n1313), .B(KEYINPUT60), .Z(n1312) );
NAND2_X1 U989 ( .A1(G107), .A2(n1314), .ZN(n1313) );
XNOR2_X1 U990 ( .A(n1119), .B(n1315), .ZN(n1176) );
NOR2_X1 U991 ( .A1(n1316), .A2(KEYINPUT50), .ZN(n1302) );
INV_X1 U992 ( .A(n1306), .ZN(n1316) );
XNOR2_X1 U993 ( .A(n1195), .B(n1317), .ZN(n1306) );
XNOR2_X1 U994 ( .A(KEYINPUT22), .B(n1191), .ZN(n1317) );
NAND2_X1 U995 ( .A1(G227), .A2(n1069), .ZN(n1191) );
XNOR2_X1 U996 ( .A(G110), .B(n1256), .ZN(n1195) );
INV_X1 U997 ( .A(n1282), .ZN(n1236) );
NAND2_X1 U998 ( .A1(n1233), .A2(n1074), .ZN(n1282) );
NOR2_X1 U999 ( .A1(n1054), .A2(n1246), .ZN(n1074) );
INV_X1 U1000 ( .A(n1288), .ZN(n1246) );
XNOR2_X1 U1001 ( .A(n1057), .B(n1318), .ZN(n1288) );
NOR2_X1 U1002 ( .A1(G475), .A2(KEYINPUT28), .ZN(n1318) );
NAND2_X1 U1003 ( .A1(n1164), .A2(n1299), .ZN(n1057) );
XNOR2_X1 U1004 ( .A(n1319), .B(n1320), .ZN(n1164) );
XOR2_X1 U1005 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1006 ( .A(n1323), .B(n1324), .Z(n1322) );
NOR2_X1 U1007 ( .A1(KEYINPUT62), .A2(n1325), .ZN(n1324) );
XOR2_X1 U1008 ( .A(G146), .B(n1111), .Z(n1325) );
NAND2_X1 U1009 ( .A1(n1326), .A2(G214), .ZN(n1323) );
NAND2_X1 U1010 ( .A1(KEYINPUT15), .A2(n1287), .ZN(n1321) );
INV_X1 U1011 ( .A(G113), .ZN(n1287) );
XOR2_X1 U1012 ( .A(n1327), .B(n1328), .Z(n1319) );
XNOR2_X1 U1013 ( .A(G122), .B(n1314), .ZN(n1328) );
XNOR2_X1 U1014 ( .A(G131), .B(G143), .ZN(n1327) );
XNOR2_X1 U1015 ( .A(n1329), .B(G478), .ZN(n1054) );
NAND2_X1 U1016 ( .A1(n1330), .A2(n1299), .ZN(n1329) );
XNOR2_X1 U1017 ( .A(n1160), .B(n1161), .ZN(n1330) );
XOR2_X1 U1018 ( .A(G107), .B(n1331), .Z(n1161) );
XOR2_X1 U1019 ( .A(G122), .B(G116), .Z(n1331) );
XOR2_X1 U1020 ( .A(n1332), .B(n1333), .Z(n1160) );
AND2_X1 U1021 ( .A1(n1334), .A2(G217), .ZN(n1333) );
NAND2_X1 U1022 ( .A1(n1335), .A2(KEYINPUT59), .ZN(n1332) );
XOR2_X1 U1023 ( .A(n1336), .B(n1337), .Z(n1335) );
XNOR2_X1 U1024 ( .A(G128), .B(G143), .ZN(n1336) );
AND2_X1 U1025 ( .A1(n1039), .A2(n1235), .ZN(n1233) );
NAND2_X1 U1026 ( .A1(n1272), .A2(n1338), .ZN(n1235) );
NAND3_X1 U1027 ( .A1(n1145), .A2(n1075), .A3(G902), .ZN(n1338) );
NOR2_X1 U1028 ( .A1(n1069), .A2(G898), .ZN(n1145) );
NAND3_X1 U1029 ( .A1(G952), .A2(n1075), .A3(n1339), .ZN(n1272) );
XNOR2_X1 U1030 ( .A(G953), .B(KEYINPUT5), .ZN(n1339) );
NAND2_X1 U1031 ( .A1(G237), .A2(n1340), .ZN(n1075) );
XOR2_X1 U1032 ( .A(KEYINPUT42), .B(G234), .Z(n1340) );
NOR2_X1 U1033 ( .A1(n1071), .A2(n1072), .ZN(n1039) );
INV_X1 U1034 ( .A(n1261), .ZN(n1072) );
NAND2_X1 U1035 ( .A1(G214), .A2(n1341), .ZN(n1261) );
XOR2_X1 U1036 ( .A(n1342), .B(n1204), .Z(n1071) );
AND2_X1 U1037 ( .A1(G210), .A2(n1341), .ZN(n1204) );
NAND2_X1 U1038 ( .A1(n1343), .A2(n1299), .ZN(n1341) );
INV_X1 U1039 ( .A(G237), .ZN(n1343) );
NAND2_X1 U1040 ( .A1(n1344), .A2(n1299), .ZN(n1342) );
XNOR2_X1 U1041 ( .A(n1345), .B(n1346), .ZN(n1344) );
XOR2_X1 U1042 ( .A(n1239), .B(n1241), .Z(n1346) );
XNOR2_X1 U1043 ( .A(G125), .B(n1347), .ZN(n1241) );
NOR2_X1 U1044 ( .A1(n1149), .A2(G953), .ZN(n1239) );
INV_X1 U1045 ( .A(G224), .ZN(n1149) );
INV_X1 U1046 ( .A(n1240), .ZN(n1345) );
XOR2_X1 U1047 ( .A(n1348), .B(n1142), .Z(n1240) );
XOR2_X1 U1048 ( .A(G122), .B(n1194), .Z(n1142) );
NAND2_X1 U1049 ( .A1(n1349), .A2(KEYINPUT4), .ZN(n1348) );
XOR2_X1 U1050 ( .A(n1143), .B(n1350), .Z(n1349) );
NOR2_X1 U1051 ( .A1(KEYINPUT10), .A2(n1144), .ZN(n1350) );
NAND3_X1 U1052 ( .A1(n1351), .A2(n1352), .A3(n1353), .ZN(n1143) );
NAND2_X1 U1053 ( .A1(n1311), .A2(n1354), .ZN(n1353) );
NOR2_X1 U1054 ( .A1(n1314), .A2(G107), .ZN(n1311) );
OR3_X1 U1055 ( .A1(n1354), .A2(G104), .A3(G107), .ZN(n1352) );
NAND2_X1 U1056 ( .A1(n1355), .A2(G107), .ZN(n1351) );
XNOR2_X1 U1057 ( .A(n1314), .B(n1354), .ZN(n1355) );
NOR2_X1 U1058 ( .A1(KEYINPUT24), .A2(n1309), .ZN(n1354) );
XNOR2_X1 U1059 ( .A(G101), .B(KEYINPUT13), .ZN(n1309) );
INV_X1 U1060 ( .A(G104), .ZN(n1314) );
NOR2_X1 U1061 ( .A1(n1292), .A2(n1291), .ZN(n1096) );
INV_X1 U1062 ( .A(n1277), .ZN(n1291) );
NAND2_X1 U1063 ( .A1(n1356), .A2(n1062), .ZN(n1277) );
NAND3_X1 U1064 ( .A1(n1357), .A2(n1299), .A3(n1153), .ZN(n1062) );
XOR2_X1 U1065 ( .A(n1061), .B(KEYINPUT56), .Z(n1356) );
NAND2_X1 U1066 ( .A1(n1155), .A2(n1358), .ZN(n1061) );
NAND2_X1 U1067 ( .A1(n1153), .A2(n1299), .ZN(n1358) );
XNOR2_X1 U1068 ( .A(n1359), .B(n1360), .ZN(n1153) );
XNOR2_X1 U1069 ( .A(n1361), .B(n1362), .ZN(n1360) );
NAND2_X1 U1070 ( .A1(n1334), .A2(G221), .ZN(n1361) );
AND2_X1 U1071 ( .A1(G234), .A2(n1069), .ZN(n1334) );
INV_X1 U1072 ( .A(G953), .ZN(n1069) );
XNOR2_X1 U1073 ( .A(KEYINPUT49), .B(n1363), .ZN(n1359) );
NOR2_X1 U1074 ( .A1(KEYINPUT32), .A2(n1364), .ZN(n1363) );
XOR2_X1 U1075 ( .A(n1365), .B(n1366), .Z(n1364) );
XNOR2_X1 U1076 ( .A(n1194), .B(n1367), .ZN(n1366) );
XOR2_X1 U1077 ( .A(KEYINPUT35), .B(G119), .Z(n1367) );
INV_X1 U1078 ( .A(G110), .ZN(n1194) );
XOR2_X1 U1079 ( .A(n1368), .B(n1369), .Z(n1365) );
NAND2_X1 U1080 ( .A1(KEYINPUT17), .A2(n1111), .ZN(n1368) );
XNOR2_X1 U1081 ( .A(G125), .B(n1256), .ZN(n1111) );
INV_X1 U1082 ( .A(G140), .ZN(n1256) );
INV_X1 U1083 ( .A(n1357), .ZN(n1155) );
NAND2_X1 U1084 ( .A1(G217), .A2(n1296), .ZN(n1357) );
NAND2_X1 U1085 ( .A1(G234), .A2(n1299), .ZN(n1296) );
XNOR2_X1 U1086 ( .A(n1065), .B(G472), .ZN(n1292) );
NAND2_X1 U1087 ( .A1(n1370), .A2(n1299), .ZN(n1065) );
INV_X1 U1088 ( .A(G902), .ZN(n1299) );
XNOR2_X1 U1089 ( .A(n1371), .B(n1169), .ZN(n1370) );
XNOR2_X1 U1090 ( .A(n1372), .B(G101), .ZN(n1169) );
NAND2_X1 U1091 ( .A1(n1326), .A2(G210), .ZN(n1372) );
NOR2_X1 U1092 ( .A1(G953), .A2(G237), .ZN(n1326) );
NAND3_X1 U1093 ( .A1(n1373), .A2(n1374), .A3(n1173), .ZN(n1371) );
NAND3_X1 U1094 ( .A1(n1147), .A2(n1347), .A3(n1118), .ZN(n1173) );
NAND2_X1 U1095 ( .A1(n1375), .A2(n1376), .ZN(n1374) );
INV_X1 U1096 ( .A(KEYINPUT31), .ZN(n1376) );
NAND2_X1 U1097 ( .A1(n1174), .A2(n1377), .ZN(n1375) );
NAND2_X1 U1098 ( .A1(n1378), .A2(n1144), .ZN(n1377) );
XNOR2_X1 U1099 ( .A(n1347), .B(n1315), .ZN(n1378) );
NAND2_X1 U1100 ( .A1(n1379), .A2(n1147), .ZN(n1174) );
INV_X1 U1101 ( .A(n1144), .ZN(n1147) );
NAND2_X1 U1102 ( .A1(KEYINPUT31), .A2(n1380), .ZN(n1373) );
XNOR2_X1 U1103 ( .A(n1379), .B(n1144), .ZN(n1380) );
XOR2_X1 U1104 ( .A(G113), .B(n1381), .Z(n1144) );
XOR2_X1 U1105 ( .A(G119), .B(G116), .Z(n1381) );
NOR2_X1 U1106 ( .A1(n1118), .A2(n1347), .ZN(n1379) );
XOR2_X1 U1107 ( .A(KEYINPUT16), .B(n1115), .Z(n1347) );
INV_X1 U1108 ( .A(n1119), .ZN(n1115) );
XOR2_X1 U1109 ( .A(G143), .B(n1369), .Z(n1119) );
XNOR2_X1 U1110 ( .A(n1262), .B(G146), .ZN(n1369) );
INV_X1 U1111 ( .A(G128), .ZN(n1262) );
INV_X1 U1112 ( .A(n1315), .ZN(n1118) );
XOR2_X1 U1113 ( .A(n1337), .B(n1382), .Z(n1315) );
XNOR2_X1 U1114 ( .A(n1259), .B(n1362), .ZN(n1382) );
XOR2_X1 U1115 ( .A(G137), .B(KEYINPUT46), .Z(n1362) );
INV_X1 U1116 ( .A(G131), .ZN(n1259) );
XOR2_X1 U1117 ( .A(G134), .B(KEYINPUT26), .Z(n1337) );
endmodule


