//Key = 0111010011111111110001111000011100000001001111100101010100101111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312;

NAND2_X1 U717 ( .A1(n997), .A2(n998), .ZN(G9) );
NAND2_X1 U718 ( .A1(n999), .A2(n1000), .ZN(n998) );
XOR2_X1 U719 ( .A(KEYINPUT14), .B(G107), .Z(n1000) );
XOR2_X1 U720 ( .A(n1001), .B(KEYINPUT63), .Z(n999) );
NAND2_X1 U721 ( .A1(n1002), .A2(G107), .ZN(n997) );
XOR2_X1 U722 ( .A(n1001), .B(KEYINPUT50), .Z(n1002) );
NOR2_X1 U723 ( .A1(n1003), .A2(n1004), .ZN(G75) );
NOR4_X1 U724 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1004) );
NOR2_X1 U725 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U726 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR3_X1 U727 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NOR2_X1 U728 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR2_X1 U729 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NOR2_X1 U730 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR2_X1 U731 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U732 ( .A1(n1024), .A2(n1025), .ZN(n1016) );
NOR2_X1 U733 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR3_X1 U734 ( .A1(n1019), .A2(n1028), .A3(n1025), .ZN(n1011) );
NOR3_X1 U735 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NOR2_X1 U736 ( .A1(n1032), .A2(n1013), .ZN(n1031) );
NOR2_X1 U737 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR2_X1 U738 ( .A1(KEYINPUT37), .A2(n1035), .ZN(n1033) );
NOR3_X1 U739 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1030) );
XNOR2_X1 U740 ( .A(KEYINPUT17), .B(n1015), .ZN(n1036) );
NOR2_X1 U741 ( .A1(n1039), .A2(n1015), .ZN(n1029) );
INV_X1 U742 ( .A(n1040), .ZN(n1015) );
NAND4_X1 U743 ( .A1(n1041), .A2(n1042), .A3(n1001), .A4(n1043), .ZN(n1005) );
NAND3_X1 U744 ( .A1(n1044), .A2(n1045), .A3(KEYINPUT37), .ZN(n1041) );
OR4_X1 U745 ( .A1(n1010), .A2(n1035), .A3(n1013), .A4(n1019), .ZN(n1045) );
NOR3_X1 U746 ( .A1(n1046), .A2(G953), .A3(G952), .ZN(n1003) );
INV_X1 U747 ( .A(n1042), .ZN(n1046) );
NAND4_X1 U748 ( .A1(n1047), .A2(n1044), .A3(n1048), .A4(n1049), .ZN(n1042) );
NOR4_X1 U749 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1049) );
XNOR2_X1 U750 ( .A(n1054), .B(KEYINPUT42), .ZN(n1053) );
XNOR2_X1 U751 ( .A(n1055), .B(n1056), .ZN(n1052) );
NAND2_X1 U752 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
XNOR2_X1 U753 ( .A(KEYINPUT9), .B(KEYINPUT30), .ZN(n1057) );
NOR3_X1 U754 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1048) );
NOR3_X1 U755 ( .A1(n1062), .A2(KEYINPUT32), .A3(n1063), .ZN(n1061) );
AND2_X1 U756 ( .A1(n1062), .A2(KEYINPUT32), .ZN(n1060) );
XNOR2_X1 U757 ( .A(KEYINPUT47), .B(n1064), .ZN(n1059) );
XOR2_X1 U758 ( .A(n1065), .B(n1066), .Z(G72) );
XOR2_X1 U759 ( .A(n1067), .B(n1068), .Z(n1066) );
NOR2_X1 U760 ( .A1(n1069), .A2(G953), .ZN(n1068) );
NOR2_X1 U761 ( .A1(n1070), .A2(n1071), .ZN(n1067) );
XOR2_X1 U762 ( .A(n1072), .B(n1073), .Z(n1071) );
XNOR2_X1 U763 ( .A(n1074), .B(n1075), .ZN(n1073) );
XOR2_X1 U764 ( .A(n1076), .B(n1077), .Z(n1075) );
XOR2_X1 U765 ( .A(n1078), .B(n1079), .Z(n1072) );
XNOR2_X1 U766 ( .A(KEYINPUT62), .B(n1080), .ZN(n1079) );
NAND2_X1 U767 ( .A1(KEYINPUT5), .A2(G140), .ZN(n1078) );
AND2_X1 U768 ( .A1(n1081), .A2(n1082), .ZN(n1070) );
NOR2_X1 U769 ( .A1(n1083), .A2(n1043), .ZN(n1065) );
AND2_X1 U770 ( .A1(G227), .A2(G900), .ZN(n1083) );
XOR2_X1 U771 ( .A(n1084), .B(n1085), .Z(G69) );
NAND2_X1 U772 ( .A1(G953), .A2(n1086), .ZN(n1085) );
NAND2_X1 U773 ( .A1(G898), .A2(G224), .ZN(n1086) );
NAND3_X1 U774 ( .A1(n1087), .A2(n1088), .A3(KEYINPUT55), .ZN(n1084) );
OR2_X1 U775 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U776 ( .A1(n1089), .A2(n1091), .ZN(n1087) );
NAND2_X1 U777 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U778 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
INV_X1 U779 ( .A(KEYINPUT23), .ZN(n1095) );
NAND2_X1 U780 ( .A1(KEYINPUT23), .A2(n1090), .ZN(n1092) );
NOR2_X1 U781 ( .A1(KEYINPUT25), .A2(n1094), .ZN(n1090) );
NAND2_X1 U782 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NAND2_X1 U783 ( .A1(n1082), .A2(n1098), .ZN(n1097) );
XOR2_X1 U784 ( .A(n1099), .B(n1100), .Z(n1096) );
AND2_X1 U785 ( .A1(n1043), .A2(n1101), .ZN(n1089) );
NAND2_X1 U786 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U787 ( .A(n1001), .B(KEYINPUT6), .Z(n1102) );
NOR2_X1 U788 ( .A1(n1104), .A2(n1105), .ZN(G66) );
XNOR2_X1 U789 ( .A(n1106), .B(n1107), .ZN(n1105) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U791 ( .A1(n1104), .A2(n1110), .ZN(G63) );
XNOR2_X1 U792 ( .A(n1111), .B(n1112), .ZN(n1110) );
NOR2_X1 U793 ( .A1(n1113), .A2(n1109), .ZN(n1112) );
NOR2_X1 U794 ( .A1(n1104), .A2(n1114), .ZN(G60) );
XOR2_X1 U795 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U796 ( .A1(n1062), .A2(n1109), .ZN(n1115) );
XNOR2_X1 U797 ( .A(G104), .B(n1117), .ZN(G6) );
NOR2_X1 U798 ( .A1(n1118), .A2(n1119), .ZN(G57) );
XOR2_X1 U799 ( .A(n1120), .B(n1121), .Z(n1119) );
XOR2_X1 U800 ( .A(n1122), .B(n1123), .Z(n1120) );
NOR2_X1 U801 ( .A1(n1124), .A2(n1109), .ZN(n1123) );
NAND3_X1 U802 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1122) );
NAND2_X1 U803 ( .A1(KEYINPUT36), .A2(n1128), .ZN(n1127) );
NAND3_X1 U804 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1126) );
NAND2_X1 U805 ( .A1(n1132), .A2(n1133), .ZN(n1125) );
NAND2_X1 U806 ( .A1(n1134), .A2(n1130), .ZN(n1133) );
INV_X1 U807 ( .A(KEYINPUT36), .ZN(n1130) );
XNOR2_X1 U808 ( .A(KEYINPUT3), .B(n1129), .ZN(n1134) );
NOR2_X1 U809 ( .A1(n1043), .A2(n1135), .ZN(n1118) );
XOR2_X1 U810 ( .A(KEYINPUT0), .B(G952), .Z(n1135) );
NOR2_X1 U811 ( .A1(n1104), .A2(n1136), .ZN(G54) );
XOR2_X1 U812 ( .A(n1137), .B(n1138), .Z(n1136) );
XNOR2_X1 U813 ( .A(n1139), .B(n1140), .ZN(n1138) );
XNOR2_X1 U814 ( .A(n1141), .B(G110), .ZN(n1140) );
XNOR2_X1 U815 ( .A(n1142), .B(n1143), .ZN(n1137) );
XNOR2_X1 U816 ( .A(n1144), .B(n1145), .ZN(n1143) );
NOR2_X1 U817 ( .A1(n1056), .A2(n1109), .ZN(n1144) );
NOR2_X1 U818 ( .A1(n1104), .A2(n1146), .ZN(G51) );
XOR2_X1 U819 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U820 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U821 ( .A1(n1151), .A2(n1109), .ZN(n1149) );
NAND2_X1 U822 ( .A1(n1152), .A2(n1153), .ZN(n1109) );
NAND3_X1 U823 ( .A1(n1069), .A2(n1001), .A3(n1103), .ZN(n1153) );
INV_X1 U824 ( .A(n1006), .ZN(n1103) );
NAND4_X1 U825 ( .A1(n1154), .A2(n1155), .A3(n1117), .A4(n1156), .ZN(n1006) );
AND4_X1 U826 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1156) );
NAND3_X1 U827 ( .A1(n1161), .A2(n1040), .A3(n1027), .ZN(n1117) );
NAND3_X1 U828 ( .A1(n1026), .A2(n1040), .A3(n1161), .ZN(n1001) );
INV_X1 U829 ( .A(n1008), .ZN(n1069) );
NAND4_X1 U830 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1008) );
NOR4_X1 U831 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
NOR2_X1 U832 ( .A1(n1170), .A2(n1171), .ZN(n1164) );
NOR4_X1 U833 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1171) );
NOR2_X1 U834 ( .A1(n1176), .A2(n1177), .ZN(n1173) );
NOR2_X1 U835 ( .A1(n1039), .A2(n1025), .ZN(n1176) );
NOR2_X1 U836 ( .A1(n1027), .A2(n1178), .ZN(n1172) );
NOR3_X1 U837 ( .A1(n1179), .A2(KEYINPUT60), .A3(n1013), .ZN(n1178) );
INV_X1 U838 ( .A(n1180), .ZN(n1013) );
NAND3_X1 U839 ( .A1(n1181), .A2(n1044), .A3(n1182), .ZN(n1163) );
NAND2_X1 U840 ( .A1(KEYINPUT60), .A2(n1183), .ZN(n1162) );
INV_X1 U841 ( .A(n1184), .ZN(n1183) );
XNOR2_X1 U842 ( .A(KEYINPUT40), .B(n1185), .ZN(n1152) );
XOR2_X1 U843 ( .A(n1186), .B(n1187), .Z(n1147) );
NOR2_X1 U844 ( .A1(KEYINPUT56), .A2(n1188), .ZN(n1186) );
XNOR2_X1 U845 ( .A(n1189), .B(n1080), .ZN(n1188) );
NOR2_X1 U846 ( .A1(n1043), .A2(G952), .ZN(n1104) );
XNOR2_X1 U847 ( .A(n1166), .B(n1190), .ZN(G48) );
NAND2_X1 U848 ( .A1(KEYINPUT2), .A2(G146), .ZN(n1190) );
NOR3_X1 U849 ( .A1(n1179), .A2(n1177), .A3(n1191), .ZN(n1166) );
XOR2_X1 U850 ( .A(G143), .B(n1170), .Z(G45) );
AND2_X1 U851 ( .A1(n1192), .A2(n1193), .ZN(n1170) );
XNOR2_X1 U852 ( .A(G140), .B(n1194), .ZN(G42) );
NAND4_X1 U853 ( .A1(KEYINPUT31), .A2(n1195), .A3(n1044), .A4(n1196), .ZN(n1194) );
XOR2_X1 U854 ( .A(n1197), .B(n1198), .Z(G39) );
NOR2_X1 U855 ( .A1(KEYINPUT33), .A2(n1199), .ZN(n1198) );
NOR3_X1 U856 ( .A1(n1200), .A2(n1019), .A3(n1191), .ZN(n1197) );
INV_X1 U857 ( .A(n1182), .ZN(n1191) );
XNOR2_X1 U858 ( .A(KEYINPUT44), .B(n1025), .ZN(n1200) );
XOR2_X1 U859 ( .A(n1201), .B(n1169), .Z(G36) );
AND3_X1 U860 ( .A1(n1044), .A2(n1026), .A3(n1192), .ZN(n1169) );
XNOR2_X1 U861 ( .A(G134), .B(KEYINPUT61), .ZN(n1201) );
XOR2_X1 U862 ( .A(G131), .B(n1168), .Z(G33) );
AND3_X1 U863 ( .A1(n1027), .A2(n1044), .A3(n1192), .ZN(n1168) );
NOR3_X1 U864 ( .A1(n1039), .A2(n1174), .A3(n1035), .ZN(n1192) );
INV_X1 U865 ( .A(n1202), .ZN(n1035) );
INV_X1 U866 ( .A(n1025), .ZN(n1044) );
NAND2_X1 U867 ( .A1(n1203), .A2(n1023), .ZN(n1025) );
INV_X1 U868 ( .A(n1022), .ZN(n1203) );
XOR2_X1 U869 ( .A(G128), .B(n1167), .Z(G30) );
AND3_X1 U870 ( .A1(n1021), .A2(n1026), .A3(n1182), .ZN(n1167) );
NOR4_X1 U871 ( .A1(n1039), .A2(n1064), .A3(n1204), .A4(n1174), .ZN(n1182) );
XNOR2_X1 U872 ( .A(G101), .B(n1205), .ZN(G3) );
NAND2_X1 U873 ( .A1(KEYINPUT39), .A2(n1206), .ZN(n1205) );
INV_X1 U874 ( .A(n1154), .ZN(n1206) );
NAND3_X1 U875 ( .A1(n1181), .A2(n1161), .A3(n1202), .ZN(n1154) );
XNOR2_X1 U876 ( .A(G125), .B(n1184), .ZN(G27) );
NAND3_X1 U877 ( .A1(n1021), .A2(n1180), .A3(n1195), .ZN(n1184) );
NOR3_X1 U878 ( .A1(n1175), .A2(n1174), .A3(n1177), .ZN(n1195) );
AND2_X1 U879 ( .A1(n1010), .A2(n1207), .ZN(n1174) );
NAND4_X1 U880 ( .A1(n1082), .A2(G902), .A3(n1208), .A4(n1081), .ZN(n1207) );
INV_X1 U881 ( .A(G900), .ZN(n1081) );
INV_X1 U882 ( .A(n1034), .ZN(n1175) );
XNOR2_X1 U883 ( .A(G122), .B(n1155), .ZN(G24) );
NAND3_X1 U884 ( .A1(n1209), .A2(n1040), .A3(n1193), .ZN(n1155) );
AND3_X1 U885 ( .A1(n1210), .A2(n1211), .A3(n1021), .ZN(n1193) );
NOR2_X1 U886 ( .A1(n1054), .A2(n1212), .ZN(n1040) );
XNOR2_X1 U887 ( .A(n1160), .B(n1213), .ZN(G21) );
NOR2_X1 U888 ( .A1(KEYINPUT19), .A2(n1214), .ZN(n1213) );
NAND3_X1 U889 ( .A1(n1021), .A2(n1209), .A3(n1215), .ZN(n1160) );
NOR3_X1 U890 ( .A1(n1019), .A2(n1204), .A3(n1064), .ZN(n1215) );
XNOR2_X1 U891 ( .A(G116), .B(n1159), .ZN(G18) );
NAND4_X1 U892 ( .A1(n1021), .A2(n1202), .A3(n1209), .A4(n1026), .ZN(n1159) );
AND2_X1 U893 ( .A1(n1216), .A2(n1210), .ZN(n1026) );
XOR2_X1 U894 ( .A(n1047), .B(KEYINPUT12), .Z(n1210) );
INV_X1 U895 ( .A(n1179), .ZN(n1021) );
XOR2_X1 U896 ( .A(n1217), .B(KEYINPUT8), .Z(n1179) );
XOR2_X1 U897 ( .A(n1158), .B(n1218), .Z(G15) );
NOR2_X1 U898 ( .A1(G113), .A2(KEYINPUT41), .ZN(n1218) );
NAND4_X1 U899 ( .A1(n1202), .A2(n1027), .A3(n1209), .A4(n1217), .ZN(n1158) );
AND2_X1 U900 ( .A1(n1180), .A2(n1219), .ZN(n1209) );
NOR2_X1 U901 ( .A1(n1037), .A2(n1051), .ZN(n1180) );
INV_X1 U902 ( .A(n1038), .ZN(n1051) );
INV_X1 U903 ( .A(n1177), .ZN(n1027) );
NAND2_X1 U904 ( .A1(n1047), .A2(n1211), .ZN(n1177) );
XOR2_X1 U905 ( .A(n1216), .B(KEYINPUT16), .Z(n1211) );
NOR2_X1 U906 ( .A1(n1212), .A2(n1204), .ZN(n1202) );
INV_X1 U907 ( .A(n1054), .ZN(n1204) );
XNOR2_X1 U908 ( .A(G110), .B(n1157), .ZN(G12) );
NAND3_X1 U909 ( .A1(n1034), .A2(n1161), .A3(n1181), .ZN(n1157) );
INV_X1 U910 ( .A(n1019), .ZN(n1181) );
NAND2_X1 U911 ( .A1(n1216), .A2(n1047), .ZN(n1019) );
XNOR2_X1 U912 ( .A(n1220), .B(n1113), .ZN(n1047) );
INV_X1 U913 ( .A(G478), .ZN(n1113) );
NAND2_X1 U914 ( .A1(n1111), .A2(n1185), .ZN(n1220) );
XNOR2_X1 U915 ( .A(n1221), .B(n1222), .ZN(n1111) );
XOR2_X1 U916 ( .A(n1223), .B(n1224), .Z(n1222) );
XNOR2_X1 U917 ( .A(n1225), .B(n1226), .ZN(n1224) );
NOR2_X1 U918 ( .A1(G128), .A2(KEYINPUT27), .ZN(n1226) );
NAND2_X1 U919 ( .A1(KEYINPUT45), .A2(n1227), .ZN(n1225) );
INV_X1 U920 ( .A(G134), .ZN(n1227) );
XOR2_X1 U921 ( .A(n1228), .B(n1229), .Z(n1221) );
XOR2_X1 U922 ( .A(G143), .B(G122), .Z(n1229) );
NAND2_X1 U923 ( .A1(G217), .A2(n1230), .ZN(n1228) );
NOR2_X1 U924 ( .A1(n1050), .A2(n1231), .ZN(n1216) );
NOR2_X1 U925 ( .A1(n1062), .A2(n1063), .ZN(n1231) );
AND2_X1 U926 ( .A1(n1063), .A2(n1062), .ZN(n1050) );
INV_X1 U927 ( .A(G475), .ZN(n1062) );
NOR2_X1 U928 ( .A1(n1116), .A2(G902), .ZN(n1063) );
XNOR2_X1 U929 ( .A(n1232), .B(n1233), .ZN(n1116) );
XOR2_X1 U930 ( .A(n1234), .B(n1235), .Z(n1233) );
XNOR2_X1 U931 ( .A(G122), .B(n1236), .ZN(n1235) );
NOR2_X1 U932 ( .A1(n1237), .A2(n1238), .ZN(n1234) );
XOR2_X1 U933 ( .A(n1239), .B(KEYINPUT29), .Z(n1238) );
NAND2_X1 U934 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
XOR2_X1 U935 ( .A(KEYINPUT1), .B(n1242), .Z(n1240) );
NOR2_X1 U936 ( .A1(n1243), .A2(n1241), .ZN(n1237) );
XNOR2_X1 U937 ( .A(n1242), .B(KEYINPUT4), .ZN(n1243) );
XNOR2_X1 U938 ( .A(G125), .B(n1141), .ZN(n1242) );
XNOR2_X1 U939 ( .A(n1244), .B(n1245), .ZN(n1232) );
NAND2_X1 U940 ( .A1(KEYINPUT21), .A2(n1246), .ZN(n1245) );
NAND2_X1 U941 ( .A1(n1247), .A2(KEYINPUT15), .ZN(n1244) );
XNOR2_X1 U942 ( .A(n1076), .B(n1248), .ZN(n1247) );
XOR2_X1 U943 ( .A(G143), .B(n1249), .Z(n1248) );
AND3_X1 U944 ( .A1(n1250), .A2(n1043), .A3(G214), .ZN(n1249) );
AND3_X1 U945 ( .A1(n1196), .A2(n1219), .A3(n1217), .ZN(n1161) );
AND2_X1 U946 ( .A1(n1022), .A2(n1023), .ZN(n1217) );
NAND2_X1 U947 ( .A1(G214), .A2(n1251), .ZN(n1023) );
XOR2_X1 U948 ( .A(n1252), .B(n1151), .Z(n1022) );
NAND2_X1 U949 ( .A1(G210), .A2(n1251), .ZN(n1151) );
NAND2_X1 U950 ( .A1(n1253), .A2(n1185), .ZN(n1251) );
NAND2_X1 U951 ( .A1(n1254), .A2(n1185), .ZN(n1252) );
XNOR2_X1 U952 ( .A(n1150), .B(n1255), .ZN(n1254) );
XNOR2_X1 U953 ( .A(KEYINPUT51), .B(n1256), .ZN(n1255) );
NOR3_X1 U954 ( .A1(KEYINPUT54), .A2(n1257), .A3(n1258), .ZN(n1256) );
NOR2_X1 U955 ( .A1(n1259), .A2(n1080), .ZN(n1258) );
XOR2_X1 U956 ( .A(KEYINPUT58), .B(n1260), .Z(n1259) );
NOR2_X1 U957 ( .A1(G125), .A2(n1260), .ZN(n1257) );
XNOR2_X1 U958 ( .A(n1189), .B(n1187), .ZN(n1260) );
AND2_X1 U959 ( .A1(G224), .A2(n1043), .ZN(n1187) );
XNOR2_X1 U960 ( .A(n1099), .B(n1261), .ZN(n1150) );
NOR2_X1 U961 ( .A1(KEYINPUT52), .A2(n1100), .ZN(n1261) );
XNOR2_X1 U962 ( .A(n1262), .B(G122), .ZN(n1100) );
XOR2_X1 U963 ( .A(n1263), .B(n1264), .Z(n1099) );
XOR2_X1 U964 ( .A(n1223), .B(n1265), .Z(n1264) );
XOR2_X1 U965 ( .A(G116), .B(G107), .Z(n1223) );
XNOR2_X1 U966 ( .A(G113), .B(n1266), .ZN(n1263) );
NAND2_X1 U967 ( .A1(n1010), .A2(n1267), .ZN(n1219) );
NAND4_X1 U968 ( .A1(n1082), .A2(G902), .A3(n1208), .A4(n1098), .ZN(n1267) );
INV_X1 U969 ( .A(G898), .ZN(n1098) );
XNOR2_X1 U970 ( .A(G953), .B(KEYINPUT49), .ZN(n1082) );
NAND3_X1 U971 ( .A1(n1208), .A2(n1043), .A3(G952), .ZN(n1010) );
NAND2_X1 U972 ( .A1(G237), .A2(G234), .ZN(n1208) );
INV_X1 U973 ( .A(n1039), .ZN(n1196) );
NAND2_X1 U974 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
NAND2_X1 U975 ( .A1(n1268), .A2(n1269), .ZN(n1037) );
OR2_X1 U976 ( .A1(n1058), .A2(G469), .ZN(n1269) );
XOR2_X1 U977 ( .A(n1270), .B(KEYINPUT34), .Z(n1268) );
NAND2_X1 U978 ( .A1(n1271), .A2(n1058), .ZN(n1270) );
NAND2_X1 U979 ( .A1(n1272), .A2(n1185), .ZN(n1058) );
XOR2_X1 U980 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U981 ( .A(n1275), .B(n1276), .ZN(n1274) );
INV_X1 U982 ( .A(n1142), .ZN(n1276) );
XOR2_X1 U983 ( .A(n1277), .B(n1278), .Z(n1142) );
INV_X1 U984 ( .A(n1074), .ZN(n1278) );
XNOR2_X1 U985 ( .A(n1279), .B(n1280), .ZN(n1074) );
NOR2_X1 U986 ( .A1(G128), .A2(KEYINPUT26), .ZN(n1280) );
NOR2_X1 U987 ( .A1(KEYINPUT20), .A2(n1141), .ZN(n1275) );
XOR2_X1 U988 ( .A(n1281), .B(n1282), .Z(n1273) );
XNOR2_X1 U989 ( .A(n1262), .B(n1283), .ZN(n1282) );
NOR2_X1 U990 ( .A1(KEYINPUT48), .A2(n1145), .ZN(n1283) );
XNOR2_X1 U991 ( .A(G107), .B(n1265), .ZN(n1145) );
XNOR2_X1 U992 ( .A(G101), .B(n1246), .ZN(n1265) );
INV_X1 U993 ( .A(G104), .ZN(n1246) );
INV_X1 U994 ( .A(G110), .ZN(n1262) );
NOR2_X1 U995 ( .A1(KEYINPUT7), .A2(n1139), .ZN(n1281) );
NAND2_X1 U996 ( .A1(G227), .A2(n1043), .ZN(n1139) );
XNOR2_X1 U997 ( .A(KEYINPUT59), .B(n1056), .ZN(n1271) );
INV_X1 U998 ( .A(G469), .ZN(n1056) );
NAND2_X1 U999 ( .A1(G221), .A2(n1284), .ZN(n1038) );
NOR2_X1 U1000 ( .A1(n1054), .A2(n1064), .ZN(n1034) );
INV_X1 U1001 ( .A(n1212), .ZN(n1064) );
XOR2_X1 U1002 ( .A(n1285), .B(n1108), .Z(n1212) );
NAND2_X1 U1003 ( .A1(G217), .A2(n1284), .ZN(n1108) );
NAND2_X1 U1004 ( .A1(G234), .A2(n1185), .ZN(n1284) );
NAND2_X1 U1005 ( .A1(n1106), .A2(n1185), .ZN(n1285) );
XNOR2_X1 U1006 ( .A(n1286), .B(n1287), .ZN(n1106) );
XOR2_X1 U1007 ( .A(n1288), .B(n1289), .Z(n1287) );
XNOR2_X1 U1008 ( .A(n1080), .B(G119), .ZN(n1289) );
INV_X1 U1009 ( .A(G125), .ZN(n1080) );
XNOR2_X1 U1010 ( .A(n1199), .B(G128), .ZN(n1288) );
XOR2_X1 U1011 ( .A(n1290), .B(n1291), .Z(n1286) );
XNOR2_X1 U1012 ( .A(G110), .B(n1292), .ZN(n1291) );
NAND2_X1 U1013 ( .A1(n1230), .A2(G221), .ZN(n1292) );
AND2_X1 U1014 ( .A1(G234), .A2(n1043), .ZN(n1230) );
XOR2_X1 U1015 ( .A(n1293), .B(n1241), .Z(n1290) );
NAND2_X1 U1016 ( .A1(KEYINPUT10), .A2(n1141), .ZN(n1293) );
INV_X1 U1017 ( .A(G140), .ZN(n1141) );
XOR2_X1 U1018 ( .A(n1294), .B(n1124), .Z(n1054) );
INV_X1 U1019 ( .A(G472), .ZN(n1124) );
NAND2_X1 U1020 ( .A1(n1295), .A2(n1185), .ZN(n1294) );
INV_X1 U1021 ( .A(G902), .ZN(n1185) );
XNOR2_X1 U1022 ( .A(n1296), .B(n1121), .ZN(n1295) );
XNOR2_X1 U1023 ( .A(n1297), .B(G101), .ZN(n1121) );
NAND3_X1 U1024 ( .A1(G210), .A2(n1043), .A3(n1250), .ZN(n1297) );
XOR2_X1 U1025 ( .A(n1253), .B(KEYINPUT38), .Z(n1250) );
INV_X1 U1026 ( .A(G237), .ZN(n1253) );
INV_X1 U1027 ( .A(G953), .ZN(n1043) );
NAND2_X1 U1028 ( .A1(KEYINPUT46), .A2(n1298), .ZN(n1296) );
XNOR2_X1 U1029 ( .A(n1128), .B(n1131), .ZN(n1298) );
INV_X1 U1030 ( .A(n1132), .ZN(n1131) );
XOR2_X1 U1031 ( .A(n1189), .B(n1277), .Z(n1132) );
NAND2_X1 U1032 ( .A1(n1299), .A2(n1300), .ZN(n1277) );
NAND2_X1 U1033 ( .A1(n1301), .A2(n1076), .ZN(n1300) );
XOR2_X1 U1034 ( .A(n1302), .B(KEYINPUT57), .Z(n1299) );
OR2_X1 U1035 ( .A1(n1076), .A2(n1301), .ZN(n1302) );
XOR2_X1 U1036 ( .A(n1077), .B(KEYINPUT11), .Z(n1301) );
XNOR2_X1 U1037 ( .A(G134), .B(n1199), .ZN(n1077) );
INV_X1 U1038 ( .A(G137), .ZN(n1199) );
XOR2_X1 U1039 ( .A(G131), .B(KEYINPUT13), .Z(n1076) );
NAND2_X1 U1040 ( .A1(n1303), .A2(n1304), .ZN(n1189) );
NAND2_X1 U1041 ( .A1(n1305), .A2(G128), .ZN(n1304) );
XOR2_X1 U1042 ( .A(KEYINPUT22), .B(n1306), .Z(n1303) );
NOR2_X1 U1043 ( .A1(G128), .A2(n1305), .ZN(n1306) );
XOR2_X1 U1044 ( .A(n1279), .B(KEYINPUT28), .Z(n1305) );
XNOR2_X1 U1045 ( .A(G143), .B(n1241), .ZN(n1279) );
XOR2_X1 U1046 ( .A(G146), .B(KEYINPUT43), .Z(n1241) );
INV_X1 U1047 ( .A(n1129), .ZN(n1128) );
NAND2_X1 U1048 ( .A1(n1307), .A2(n1308), .ZN(n1129) );
NAND2_X1 U1049 ( .A1(n1309), .A2(n1236), .ZN(n1308) );
XOR2_X1 U1050 ( .A(KEYINPUT24), .B(n1310), .Z(n1309) );
XOR2_X1 U1051 ( .A(KEYINPUT53), .B(n1311), .Z(n1307) );
NOR2_X1 U1052 ( .A1(n1312), .A2(n1236), .ZN(n1311) );
INV_X1 U1053 ( .A(G113), .ZN(n1236) );
XNOR2_X1 U1054 ( .A(n1310), .B(KEYINPUT35), .ZN(n1312) );
XOR2_X1 U1055 ( .A(G116), .B(n1266), .Z(n1310) );
XNOR2_X1 U1056 ( .A(n1214), .B(KEYINPUT18), .ZN(n1266) );
INV_X1 U1057 ( .A(G119), .ZN(n1214) );
endmodule


