//Key = 1001000010110100011011000011011111111101111110011000000111111111
module c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, 
        G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, 
        G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, 
        G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, 
        G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, 
        G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, 
        G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, 
        G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, 
        G136, G137, G138, G139, G140, G141, G142, G452, G483, G543, G559, G567, 
        G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, 
        G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, 
        G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, 
        G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, G350, G335, 
        G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, 
        G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, 
        G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, 
        G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, 
        G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, 
        G308, G225, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, 
        KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, 
        KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, 
        KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, 
        KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, 
        KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, 
        KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, 
        KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, 
        KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, 
        KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, 
        KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63 );
  
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G452, G483, G543,
         G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956,
         G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067,
         G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427,
         G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678,
         KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
         KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
         KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
         KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
         KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
         KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
         KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
         KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
         KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
         KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
         KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
         KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
         KEYINPUT62, KEYINPUT63;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;

  wire   n1548, n1555, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036;

  INV_X1 U1125 ( .A(G452), .ZN(n1548) );
  INV_X1 U1126 ( .A(n1548), .ZN(G335) );
  INV_X1 U1127 ( .A(n1548), .ZN(G350) );
  INV_X1 U1128 ( .A(n1548), .ZN(G409) );
  INV_X1 U1129 ( .A(n1548), .ZN(G391) );
  BUF_X1 U1130 ( .A(G1083), .Z(G369) );
  BUF_X1 U1131 ( .A(G1083), .Z(G367) );
  INV_X1 U1132 ( .A(G2066), .ZN(n1555) );
  INV_X1 U1133 ( .A(n1555), .ZN(G337) );
  INV_X1 U1134 ( .A(n1555), .ZN(G411) );
  INV_X1 U1135 ( .A(n1555), .ZN(G384) );
  BUF_X1 U1136 ( .A(G321), .Z(G284) );
  BUF_X1 U1137 ( .A(G323), .Z(G282) );
  BUF_X1 U1138 ( .A(G331), .Z(G295) );
  BUF_X1 U1139 ( .A(G297), .Z(G280) );
  NAND2_X1 U1140 ( .A1(n1563), .A2(n1564), .ZN(G331) );
  NAND2_X1 U1141 ( .A1(n1565), .A2(n1566), .ZN(n1564) );
  NAND2_X1 U1142 ( .A1(G868), .A2(n1567), .ZN(n1563) );
  XOR2_X1 U1143 ( .A(n1568), .B(n1569), .Z(n1567) );
  XOR2_X1 U1144 ( .A(n1570), .B(n1571), .Z(n1569) );
  NAND2_X1 U1145 ( .A1(n1572), .A2(n1573), .ZN(n1570) );
  NAND2_X1 U1146 ( .A1(n1574), .A2(n1575), .ZN(n1573) );
  NAND2_X1 U1147 ( .A1(n1576), .A2(KEYINPUT32), .ZN(n1574) );
  NAND2_X1 U1148 ( .A1(n1576), .A2(n1577), .ZN(n1572) );
  XNOR2_X1 U1149 ( .A(KEYINPUT59), .B(n1578), .ZN(n1576) );
  XOR2_X1 U1150 ( .A(n1579), .B(n1580), .Z(n1568) );
  XOR2_X1 U1151 ( .A(G303), .B(n1581), .Z(n1580) );
  NAND2_X1 U1152 ( .A1(n1582), .A2(n1583), .ZN(G323) );
  NAND2_X1 U1153 ( .A1(n1584), .A2(n1566), .ZN(n1583) );
  NAND2_X1 U1154 ( .A1(G868), .A2(n1575), .ZN(n1582) );
  NAND2_X1 U1155 ( .A1(n1585), .A2(n1586), .ZN(G321) );
  NAND2_X1 U1156 ( .A1(n1587), .A2(n1566), .ZN(n1586) );
  NAND2_X1 U1157 ( .A1(G868), .A2(G301), .ZN(n1585) );
  INV_X1 U1158 ( .A(G150), .ZN(G311) );
  INV_X1 U1159 ( .A(G225), .ZN(G308) );
  NAND2_X1 U1160 ( .A1(n1588), .A2(n1589), .ZN(G297) );
  NAND2_X1 U1161 ( .A1(G868), .A2(n1590), .ZN(n1589) );
  NAND2_X1 U1162 ( .A1(n1591), .A2(n1566), .ZN(n1588) );
  INV_X1 U1163 ( .A(G868), .ZN(n1566) );
  XOR2_X1 U1164 ( .A(KEYINPUT18), .B(n1592), .Z(n1591) );
  XOR2_X1 U1165 ( .A(n1590), .B(KEYINPUT9), .Z(G286) );
  INV_X1 U1166 ( .A(G325), .ZN(G261) );
  NOR2_X1 U1167 ( .A1(n1593), .A2(n1594), .ZN(G325) );
  NAND3_X1 U1168 ( .A1(G2), .A2(G15), .A3(G661), .ZN(G259) );
  INV_X1 U1169 ( .A(G108), .ZN(G238) );
  INV_X1 U1170 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1171 ( .A(G120), .B(KEYINPUT25), .ZN(G236) );
  INV_X1 U1172 ( .A(G69), .ZN(G235) );
  NAND2_X1 U1173 ( .A1(G567), .A2(n1595), .ZN(G234) );
  INV_X1 U1174 ( .A(n1596), .ZN(G231) );
  NAND4_X1 U1175 ( .A1(n1596), .A2(n1597), .A3(G319), .A4(n1598), .ZN(G225) );
  NOR4_X1 U1176 ( .A1(G401), .A2(G397), .A3(G395), .A4(G227), .ZN(n1598) );
  XNOR2_X1 U1177 ( .A(n1599), .B(n1600), .ZN(G227) );
  NOR2_X1 U1178 ( .A1(KEYINPUT19), .A2(n1601), .ZN(n1600) );
  INV_X1 U1179 ( .A(G2100), .ZN(n1601) );
  XOR2_X1 U1180 ( .A(n1602), .B(G2096), .Z(n1599) );
  NAND2_X1 U1181 ( .A1(n1603), .A2(n1604), .ZN(n1602) );
  NAND3_X1 U1182 ( .A1(n1605), .A2(n1606), .A3(n1607), .ZN(n1604) );
  NAND2_X1 U1183 ( .A1(n1608), .A2(KEYINPUT62), .ZN(n1607) );
  NAND2_X1 U1184 ( .A1(n1609), .A2(n1610), .ZN(n1606) );
  NAND2_X1 U1185 ( .A1(KEYINPUT27), .A2(n1611), .ZN(n1610) );
  NAND2_X1 U1186 ( .A1(n1612), .A2(n1611), .ZN(n1605) );
  NAND4_X1 U1187 ( .A1(n1608), .A2(n1613), .A3(n1614), .A4(n1615), .ZN(n1603) );
  NAND2_X1 U1188 ( .A1(n1616), .A2(KEYINPUT27), .ZN(n1615) );
  OR2_X1 U1189 ( .A1(n1616), .A2(KEYINPUT62), .ZN(n1614) );
  AND2_X1 U1190 ( .A1(n1609), .A2(n1611), .ZN(n1616) );
  OR2_X1 U1191 ( .A1(n1611), .A2(n1609), .ZN(n1613) );
  INV_X1 U1192 ( .A(n1612), .ZN(n1609) );
  XOR2_X1 U1193 ( .A(n1617), .B(G2678), .Z(n1612) );
  XOR2_X1 U1194 ( .A(n1618), .B(n1619), .Z(n1611) );
  XNOR2_X1 U1195 ( .A(G2072), .B(G2078), .ZN(n1608) );
  AND2_X1 U1196 ( .A1(n1620), .A2(n1621), .ZN(G395) );
  XOR2_X1 U1197 ( .A(n1622), .B(n1623), .Z(n1620) );
  XOR2_X1 U1198 ( .A(n1624), .B(n1625), .Z(n1623) );
  NOR2_X1 U1199 ( .A1(n1626), .A2(n1627), .ZN(n1625) );
  XOR2_X1 U1200 ( .A(KEYINPUT52), .B(n1628), .Z(n1627) );
  NOR2_X1 U1201 ( .A1(G160), .A2(n1629), .ZN(n1628) );
  NOR2_X1 U1202 ( .A1(G162), .A2(n1630), .ZN(n1626) );
  NAND2_X1 U1203 ( .A1(n1631), .A2(n1632), .ZN(n1624) );
  NAND2_X1 U1204 ( .A1(n1633), .A2(n1634), .ZN(n1632) );
  NAND2_X1 U1205 ( .A1(KEYINPUT56), .A2(n1635), .ZN(n1634) );
  INV_X1 U1206 ( .A(n1636), .ZN(n1633) );
  NAND2_X1 U1207 ( .A1(n1635), .A2(n1636), .ZN(n1631) );
  NAND2_X1 U1208 ( .A1(n1637), .A2(n1638), .ZN(n1636) );
  NAND2_X1 U1209 ( .A1(n1639), .A2(n1640), .ZN(n1638) );
  XOR2_X1 U1210 ( .A(KEYINPUT40), .B(n1641), .Z(n1637) );
  NOR2_X1 U1211 ( .A1(n1639), .A2(n1640), .ZN(n1641) );
  XOR2_X1 U1212 ( .A(n1642), .B(n1643), .Z(n1635) );
  NAND4_X1 U1213 ( .A1(n1644), .A2(n1645), .A3(n1646), .A4(n1647), .ZN(n1643) );
  NAND3_X1 U1214 ( .A1(n1648), .A2(n1649), .A3(G142), .ZN(n1647) );
  OR2_X1 U1215 ( .A1(n1650), .A2(KEYINPUT0), .ZN(n1649) );
  NAND2_X1 U1216 ( .A1(KEYINPUT0), .A2(n1651), .ZN(n1648) );
  NAND2_X1 U1217 ( .A1(G106), .A2(n1652), .ZN(n1646) );
  NAND2_X1 U1218 ( .A1(G118), .A2(n1653), .ZN(n1645) );
  NAND2_X1 U1219 ( .A1(G130), .A2(n1650), .ZN(n1644) );
  XOR2_X1 U1220 ( .A(n1654), .B(n1655), .Z(n1622) );
  XNOR2_X1 U1221 ( .A(G164), .B(n1656), .ZN(n1655) );
  AND3_X1 U1222 ( .A1(n1657), .A2(n1658), .A3(n1621), .ZN(G397) );
  INV_X1 U1223 ( .A(G37), .ZN(n1621) );
  NAND2_X1 U1224 ( .A1(n1659), .A2(n1660), .ZN(n1658) );
  NAND2_X1 U1225 ( .A1(n1661), .A2(n1662), .ZN(n1660) );
  NAND3_X1 U1226 ( .A1(n1661), .A2(n1662), .A3(n1663), .ZN(n1657) );
  INV_X1 U1227 ( .A(n1659), .ZN(n1663) );
  XOR2_X1 U1228 ( .A(n1664), .B(n1665), .Z(n1659) );
  XOR2_X1 U1229 ( .A(G168), .B(n1571), .Z(n1665) );
  XOR2_X1 U1230 ( .A(n1666), .B(n1667), .Z(n1571) );
  XOR2_X1 U1231 ( .A(G301), .B(n1578), .Z(n1664) );
  XOR2_X1 U1232 ( .A(n1668), .B(n1592), .Z(n1578) );
  NAND2_X1 U1233 ( .A1(n1579), .A2(n1669), .ZN(n1662) );
  INV_X1 U1234 ( .A(n1670), .ZN(n1579) );
  XNOR2_X1 U1235 ( .A(KEYINPUT16), .B(n1671), .ZN(n1661) );
  AND2_X1 U1236 ( .A1(n1672), .A2(n1670), .ZN(n1671) );
  XNOR2_X1 U1237 ( .A(G290), .B(n1673), .ZN(n1670) );
  XNOR2_X1 U1238 ( .A(n1669), .B(n1674), .ZN(n1672) );
  XOR2_X1 U1239 ( .A(KEYINPUT28), .B(KEYINPUT14), .Z(n1674) );
  XNOR2_X1 U1240 ( .A(n1675), .B(n1581), .ZN(n1669) );
  XNOR2_X1 U1241 ( .A(n1676), .B(KEYINPUT37), .ZN(n1581) );
  NAND2_X1 U1242 ( .A1(KEYINPUT36), .A2(G166), .ZN(n1675) );
  AND2_X1 U1243 ( .A1(n1677), .A2(G14), .ZN(G401) );
  XOR2_X1 U1244 ( .A(n1678), .B(n1679), .Z(n1677) );
  XOR2_X1 U1245 ( .A(n1680), .B(n1681), .Z(n1679) );
  XNOR2_X1 U1246 ( .A(G2427), .B(n1682), .ZN(n1681) );
  NOR2_X1 U1247 ( .A1(KEYINPUT53), .A2(n1683), .ZN(n1682) );
  XOR2_X1 U1248 ( .A(n1684), .B(n1685), .Z(n1683) );
  XOR2_X1 U1249 ( .A(G1348), .B(G1341), .Z(n1685) );
  XNOR2_X1 U1250 ( .A(G2454), .B(G2451), .ZN(n1684) );
  NAND3_X1 U1251 ( .A1(n1686), .A2(n1687), .A3(n1688), .ZN(n1680) );
  OR2_X1 U1252 ( .A1(n1689), .A2(G2446), .ZN(n1688) );
  NAND3_X1 U1253 ( .A1(G2446), .A2(n1689), .A3(KEYINPUT41), .ZN(n1687) );
  NOR2_X1 U1254 ( .A1(KEYINPUT22), .A2(n1690), .ZN(n1689) );
  INV_X1 U1255 ( .A(G2443), .ZN(n1690) );
  OR2_X1 U1256 ( .A1(G2443), .A2(KEYINPUT41), .ZN(n1686) );
  XOR2_X1 U1257 ( .A(n1691), .B(G2430), .Z(n1678) );
  XNOR2_X1 U1258 ( .A(G2438), .B(G2435), .ZN(n1691) );
  INV_X1 U1259 ( .A(G229), .ZN(n1597) );
  XOR2_X1 U1260 ( .A(n1692), .B(n1693), .Z(G229) );
  XOR2_X1 U1261 ( .A(G1971), .B(G1966), .Z(n1693) );
  XOR2_X1 U1262 ( .A(n1694), .B(n1695), .Z(n1692) );
  XOR2_X1 U1263 ( .A(n1696), .B(n1697), .Z(n1695) );
  XNOR2_X1 U1264 ( .A(n1698), .B(n1699), .ZN(n1697) );
  NAND2_X1 U1265 ( .A1(KEYINPUT44), .A2(G1981), .ZN(n1699) );
  NAND2_X1 U1266 ( .A1(KEYINPUT10), .A2(G2474), .ZN(n1698) );
  XOR2_X1 U1267 ( .A(n1700), .B(G1956), .Z(n1696) );
  XOR2_X1 U1268 ( .A(n1701), .B(n1702), .Z(n1694) );
  XOR2_X1 U1269 ( .A(G1996), .B(G1991), .Z(n1702) );
  XOR2_X1 U1270 ( .A(G1986), .B(n1703), .Z(n1701) );
  XOR2_X1 U1271 ( .A(G329), .B(n1704), .Z(n1596) );
  NOR2_X1 U1272 ( .A1(n1705), .A2(n1706), .ZN(n1704) );
  NOR2_X1 U1273 ( .A1(n1707), .A2(G2067), .ZN(n1706) );
  NOR2_X1 U1274 ( .A1(n1708), .A2(n1709), .ZN(n1707) );
  AND2_X1 U1275 ( .A1(n1710), .A2(n1711), .ZN(n1708) );
  AND2_X1 U1276 ( .A1(n1710), .A2(n1709), .ZN(n1705) );
  NAND2_X1 U1277 ( .A1(n1712), .A2(n1713), .ZN(n1709) );
  NAND3_X1 U1278 ( .A1(n1639), .A2(n1714), .A3(n1711), .ZN(n1713) );
  NAND2_X1 U1279 ( .A1(n1715), .A2(n1716), .ZN(n1712) );
  NAND2_X1 U1280 ( .A1(n1711), .A2(n1717), .ZN(n1716) );
  NAND2_X1 U1281 ( .A1(n1718), .A2(n1719), .ZN(n1717) );
  NAND2_X1 U1282 ( .A1(n1720), .A2(n1721), .ZN(n1719) );
  NAND2_X1 U1283 ( .A1(KEYINPUT58), .A2(n1714), .ZN(n1720) );
  XOR2_X1 U1284 ( .A(G1996), .B(KEYINPUT42), .Z(n1714) );
  NAND2_X1 U1285 ( .A1(G1991), .A2(n1642), .ZN(n1718) );
  NAND2_X1 U1286 ( .A1(n1722), .A2(n1723), .ZN(n1715) );
  NAND3_X1 U1287 ( .A1(n1724), .A2(n1725), .A3(n1726), .ZN(n1723) );
  OR2_X1 U1288 ( .A1(n1727), .A2(n1728), .ZN(n1726) );
  NAND3_X1 U1289 ( .A1(n1711), .A2(G290), .A3(n1729), .ZN(n1725) );
  NAND2_X1 U1290 ( .A1(n1730), .A2(n1731), .ZN(n1724) );
  NAND2_X1 U1291 ( .A1(n1732), .A2(n1733), .ZN(n1731) );
  NAND2_X1 U1292 ( .A1(n1728), .A2(n1734), .ZN(n1733) );
  NAND2_X1 U1293 ( .A1(n1735), .A2(n1736), .ZN(n1734) );
  NAND2_X1 U1294 ( .A1(n1737), .A2(G288), .ZN(n1736) );
  NAND2_X1 U1295 ( .A1(n1738), .A2(n1727), .ZN(n1737) );
  XOR2_X1 U1296 ( .A(KEYINPUT5), .B(n1739), .Z(n1738) );
  OR2_X1 U1297 ( .A1(n1727), .A2(n1739), .ZN(n1732) );
  XNOR2_X1 U1298 ( .A(n1703), .B(KEYINPUT61), .ZN(n1739) );
  NAND2_X1 U1299 ( .A1(n1740), .A2(n1741), .ZN(n1727) );
  NAND2_X1 U1300 ( .A1(n1742), .A2(n1743), .ZN(n1741) );
  NAND2_X1 U1301 ( .A1(n1744), .A2(n1745), .ZN(n1743) );
  NAND2_X1 U1302 ( .A1(KEYINPUT33), .A2(n1746), .ZN(n1745) );
  INV_X1 U1303 ( .A(n1747), .ZN(n1744) );
  NAND2_X1 U1304 ( .A1(n1748), .A2(n1749), .ZN(n1742) );
  NAND3_X1 U1305 ( .A1(n1750), .A2(n1751), .A3(n1752), .ZN(n1748) );
  NAND2_X1 U1306 ( .A1(n1753), .A2(n1754), .ZN(n1752) );
  NAND3_X1 U1307 ( .A1(n1755), .A2(n1756), .A3(n1757), .ZN(n1754) );
  OR2_X1 U1308 ( .A1(n1758), .A2(KEYINPUT30), .ZN(n1756) );
  NAND3_X1 U1309 ( .A1(n1759), .A2(n1758), .A3(KEYINPUT30), .ZN(n1755) );
  NAND2_X1 U1310 ( .A1(n1760), .A2(n1761), .ZN(n1751) );
  XOR2_X1 U1311 ( .A(n1762), .B(KEYINPUT43), .Z(n1760) );
  NAND2_X1 U1312 ( .A1(G301), .A2(n1763), .ZN(n1750) );
  NAND2_X1 U1313 ( .A1(n1758), .A2(n1757), .ZN(n1763) );
  XNOR2_X1 U1314 ( .A(n1753), .B(KEYINPUT50), .ZN(n1758) );
  NAND2_X1 U1315 ( .A1(n1747), .A2(n1746), .ZN(n1740) );
  NAND3_X1 U1316 ( .A1(n1764), .A2(G303), .A3(G8), .ZN(n1747) );
  OR2_X1 U1317 ( .A1(KEYINPUT63), .A2(n1765), .ZN(n1764) );
  NAND2_X1 U1318 ( .A1(n1711), .A2(n1766), .ZN(n1722) );
  NAND2_X1 U1319 ( .A1(n1767), .A2(n1768), .ZN(n1766) );
  NAND2_X1 U1320 ( .A1(n1769), .A2(n1770), .ZN(n1767) );
  NAND2_X1 U1321 ( .A1(n1771), .A2(n1772), .ZN(G329) );
  NAND3_X1 U1322 ( .A1(n1710), .A2(n1617), .A3(n1773), .ZN(n1772) );
  NAND4_X1 U1323 ( .A1(n1774), .A2(n1775), .A3(n1776), .A4(n1777), .ZN(n1771) );
  NAND4_X1 U1324 ( .A1(n1778), .A2(n1779), .A3(n1773), .A4(n1780), .ZN(n1777) );
  INV_X1 U1325 ( .A(KEYINPUT39), .ZN(n1780) );
  NAND2_X1 U1326 ( .A1(n1781), .A2(n1782), .ZN(n1778) );
  NAND2_X1 U1327 ( .A1(n1639), .A2(n1783), .ZN(n1782) );
  INV_X1 U1328 ( .A(n1721), .ZN(n1639) );
  NAND3_X1 U1329 ( .A1(n1784), .A2(n1785), .A3(KEYINPUT39), .ZN(n1776) );
  NAND2_X1 U1330 ( .A1(n1781), .A2(n1783), .ZN(n1785) );
  INV_X1 U1331 ( .A(KEYINPUT54), .ZN(n1783) );
  NAND2_X1 U1332 ( .A1(n1773), .A2(n1779), .ZN(n1784) );
  NAND3_X1 U1333 ( .A1(n1786), .A2(n1721), .A3(n1711), .ZN(n1775) );
  NAND3_X1 U1334 ( .A1(n1781), .A2(n1779), .A3(KEYINPUT8), .ZN(n1786) );
  NAND3_X1 U1335 ( .A1(n1787), .A2(n1788), .A3(n1789), .ZN(n1781) );
  NAND2_X1 U1336 ( .A1(n1790), .A2(n1791), .ZN(n1789) );
  NAND2_X1 U1337 ( .A1(n1792), .A2(n1793), .ZN(n1791) );
  NAND3_X1 U1338 ( .A1(n1769), .A2(n1794), .A3(n1773), .ZN(n1793) );
  NAND2_X1 U1339 ( .A1(n1795), .A2(n1796), .ZN(n1792) );
  NAND2_X1 U1340 ( .A1(n1797), .A2(n1798), .ZN(n1796) );
  NAND2_X1 U1341 ( .A1(n1773), .A2(n1769), .ZN(n1798) );
  INV_X1 U1342 ( .A(n1794), .ZN(n1797) );
  NAND2_X1 U1343 ( .A1(n1799), .A2(n1800), .ZN(n1794) );
  NAND2_X1 U1344 ( .A1(n1728), .A2(n1801), .ZN(n1800) );
  NAND2_X1 U1345 ( .A1(n1730), .A2(n1802), .ZN(n1801) );
  NAND3_X1 U1346 ( .A1(n1676), .A2(n1703), .A3(n1735), .ZN(n1802) );
  INV_X1 U1347 ( .A(G288), .ZN(n1676) );
  NAND2_X1 U1348 ( .A1(n1803), .A2(n1673), .ZN(n1730) );
  NAND3_X1 U1349 ( .A1(n1804), .A2(n1805), .A3(n1806), .ZN(n1799) );
  OR2_X1 U1350 ( .A1(n1746), .A2(n1807), .ZN(n1806) );
  NAND3_X1 U1351 ( .A1(n1808), .A2(G303), .A3(G8), .ZN(n1805) );
  NAND2_X1 U1352 ( .A1(n1746), .A2(n1807), .ZN(n1808) );
  NAND3_X1 U1353 ( .A1(n1809), .A2(n1810), .A3(n1749), .ZN(n1807) );
  NAND2_X1 U1354 ( .A1(n1811), .A2(n1762), .ZN(n1749) );
  NAND3_X1 U1355 ( .A1(n1812), .A2(n1757), .A3(n1813), .ZN(n1810) );
  XOR2_X1 U1356 ( .A(n1814), .B(KEYINPUT1), .Z(n1813) );
  NAND2_X1 U1357 ( .A1(n1815), .A2(n1816), .ZN(n1757) );
  NAND3_X1 U1358 ( .A1(n1817), .A2(n1818), .A3(n1819), .ZN(n1816) );
  NAND2_X1 U1359 ( .A1(n1820), .A2(n1821), .ZN(n1818) );
  NAND3_X1 U1360 ( .A1(n1822), .A2(n1823), .A3(n1824), .ZN(n1820) );
  NAND2_X1 U1361 ( .A1(G1956), .A2(G299), .ZN(n1824) );
  NAND2_X1 U1362 ( .A1(G1348), .A2(n1825), .ZN(n1823) );
  NAND2_X1 U1363 ( .A1(n1826), .A2(n1827), .ZN(n1825) );
  INV_X1 U1364 ( .A(G1341), .ZN(n1827) );
  NAND2_X1 U1365 ( .A1(G1341), .A2(n1587), .ZN(n1822) );
  NAND2_X1 U1366 ( .A1(n1765), .A2(n1828), .ZN(n1817) );
  NAND3_X1 U1367 ( .A1(n1829), .A2(n1830), .A3(n1831), .ZN(n1828) );
  NAND2_X1 U1368 ( .A1(G2072), .A2(G299), .ZN(n1831) );
  NAND2_X1 U1369 ( .A1(G2067), .A2(n1832), .ZN(n1830) );
  NAND2_X1 U1370 ( .A1(n1826), .A2(n1779), .ZN(n1832) );
  INV_X1 U1371 ( .A(G1996), .ZN(n1779) );
  NAND2_X1 U1372 ( .A1(G1996), .A2(n1587), .ZN(n1829) );
  NAND3_X1 U1373 ( .A1(n1833), .A2(n1834), .A3(n1592), .ZN(n1815) );
  NAND2_X1 U1374 ( .A1(G1956), .A2(n1821), .ZN(n1834) );
  NAND2_X1 U1375 ( .A1(n1765), .A2(G2072), .ZN(n1833) );
  XOR2_X1 U1376 ( .A(n1835), .B(G301), .Z(n1812) );
  NAND2_X1 U1377 ( .A1(KEYINPUT48), .A2(n1836), .ZN(n1835) );
  NAND3_X1 U1378 ( .A1(n1759), .A2(n1814), .A3(n1837), .ZN(n1809) );
  XOR2_X1 U1379 ( .A(KEYINPUT55), .B(n1753), .Z(n1837) );
  INV_X1 U1380 ( .A(n1836), .ZN(n1753) );
  NAND2_X1 U1381 ( .A1(n1838), .A2(n1839), .ZN(n1836) );
  OR2_X1 U1382 ( .A1(n1821), .A2(G2078), .ZN(n1839) );
  NAND2_X1 U1383 ( .A1(n1821), .A2(n1700), .ZN(n1838) );
  NAND2_X1 U1384 ( .A1(n1840), .A2(n1841), .ZN(n1814) );
  OR2_X1 U1385 ( .A1(KEYINPUT24), .A2(n1761), .ZN(n1841) );
  INV_X1 U1386 ( .A(n1811), .ZN(n1761) );
  NAND2_X1 U1387 ( .A1(G8), .A2(n1590), .ZN(n1811) );
  INV_X1 U1388 ( .A(n1762), .ZN(n1840) );
  NAND2_X1 U1389 ( .A1(n1842), .A2(n1843), .ZN(n1762) );
  NAND3_X1 U1390 ( .A1(G8), .A2(n1618), .A3(n1765), .ZN(n1843) );
  INV_X1 U1391 ( .A(G2084), .ZN(n1618) );
  OR2_X1 U1392 ( .A1(n1844), .A2(G1966), .ZN(n1842) );
  INV_X1 U1393 ( .A(G301), .ZN(n1759) );
  XNOR2_X1 U1394 ( .A(G171), .B(KEYINPUT45), .ZN(G301) );
  NAND2_X1 U1395 ( .A1(n1845), .A2(n1846), .ZN(n1746) );
  NAND3_X1 U1396 ( .A1(G8), .A2(n1619), .A3(n1765), .ZN(n1846) );
  INV_X1 U1397 ( .A(G2090), .ZN(n1619) );
  NAND2_X1 U1398 ( .A1(n1728), .A2(n1847), .ZN(n1845) );
  NAND2_X1 U1399 ( .A1(n1728), .A2(n1848), .ZN(n1804) );
  NAND2_X1 U1400 ( .A1(n1735), .A2(n1849), .ZN(n1848) );
  NAND2_X1 U1401 ( .A1(G1976), .A2(G288), .ZN(n1849) );
  OR2_X1 U1402 ( .A1(n1803), .A2(n1673), .ZN(n1735) );
  INV_X1 U1403 ( .A(n1844), .ZN(n1728) );
  NAND2_X1 U1404 ( .A1(G8), .A2(n1821), .ZN(n1844) );
  XOR2_X1 U1405 ( .A(KEYINPUT60), .B(n1850), .Z(n1795) );
  NOR3_X1 U1406 ( .A1(n1851), .A2(n1770), .A3(n1765), .ZN(n1850) );
  INV_X1 U1407 ( .A(n1821), .ZN(n1765) );
  NAND3_X1 U1408 ( .A1(G40), .A2(G160), .A3(n1852), .ZN(n1821) );
  INV_X1 U1409 ( .A(G290), .ZN(n1770) );
  XOR2_X1 U1410 ( .A(KEYINPUT13), .B(n1711), .Z(n1851) );
  XOR2_X1 U1411 ( .A(n1853), .B(n1854), .Z(n1790) );
  NOR3_X1 U1412 ( .A1(n1855), .A2(KEYINPUT49), .A3(n1856), .ZN(n1854) );
  XOR2_X1 U1413 ( .A(n1857), .B(KEYINPUT7), .Z(n1853) );
  NAND2_X1 U1414 ( .A1(n1858), .A2(n1859), .ZN(n1788) );
  NAND2_X1 U1415 ( .A1(n1860), .A2(n1773), .ZN(n1858) );
  OR3_X1 U1416 ( .A1(n1857), .A2(n1642), .A3(n1859), .ZN(n1787) );
  INV_X1 U1417 ( .A(KEYINPUT34), .ZN(n1859) );
  NAND2_X1 U1418 ( .A1(n1773), .A2(n1861), .ZN(n1857) );
  XOR2_X1 U1419 ( .A(n1862), .B(n1863), .Z(n1774) );
  XNOR2_X1 U1420 ( .A(KEYINPUT6), .B(n1710), .ZN(n1863) );
  NAND2_X1 U1421 ( .A1(n1864), .A2(n1711), .ZN(n1710) );
  XOR2_X1 U1422 ( .A(n1640), .B(KEYINPUT51), .Z(n1864) );
  NAND2_X1 U1423 ( .A1(n1773), .A2(n1617), .ZN(n1862) );
  AND2_X1 U1424 ( .A1(KEYINPUT8), .A2(n1711), .ZN(n1773) );
  INV_X1 U1425 ( .A(n1855), .ZN(n1711) );
  NAND3_X1 U1426 ( .A1(G160), .A2(n1865), .A3(G40), .ZN(n1855) );
  INV_X1 U1427 ( .A(n1852), .ZN(n1865) );
  NOR2_X1 U1428 ( .A1(G164), .A2(G1384), .ZN(n1852) );
  INV_X1 U1429 ( .A(G96), .ZN(G221) );
  INV_X1 U1430 ( .A(G82), .ZN(G220) );
  INV_X1 U1431 ( .A(G132), .ZN(G219) );
  INV_X1 U1432 ( .A(G44), .ZN(G218) );
  NAND2_X1 U1433 ( .A1(G2106), .A2(n1595), .ZN(G217) );
  INV_X1 U1434 ( .A(G223), .ZN(n1595) );
  NAND2_X1 U1435 ( .A1(G7), .A2(n1866), .ZN(G223) );
  XOR2_X1 U1436 ( .A(KEYINPUT23), .B(G661), .Z(n1866) );
  NAND2_X1 U1437 ( .A1(n1867), .A2(n1868), .ZN(G188) );
  NAND2_X1 U1438 ( .A1(G3), .A2(G1), .ZN(n1868) );
  NAND2_X1 U1439 ( .A1(G36), .A2(n1867), .ZN(G176) );
  AND3_X1 U1440 ( .A1(G661), .A2(G319), .A3(G483), .ZN(n1867) );
  AND2_X1 U1441 ( .A1(n1869), .A2(n1870), .ZN(G319) );
  NAND2_X1 U1442 ( .A1(G2106), .A2(n1593), .ZN(n1870) );
  NAND4_X1 U1443 ( .A1(G44), .A2(G132), .A3(G82), .A4(G96), .ZN(n1593) );
  NAND2_X1 U1444 ( .A1(G567), .A2(n1594), .ZN(n1869) );
  NAND4_X1 U1445 ( .A1(G120), .A2(G69), .A3(G57), .A4(G108), .ZN(n1594) );
  AND2_X1 U1446 ( .A1(G94), .A2(G452), .ZN(G173) );
  INV_X1 U1447 ( .A(n1590), .ZN(G168) );
  INV_X1 U1448 ( .A(G303), .ZN(G166) );
  INV_X1 U1449 ( .A(n1629), .ZN(G162) );
  INV_X1 U1450 ( .A(n1630), .ZN(G160) );
  NAND4_X1 U1451 ( .A1(G2090), .A2(G2084), .A3(G2078), .A4(G2072), .ZN(G158) );
  NAND2_X1 U1452 ( .A1(n1871), .A2(n1872), .ZN(G156) );
  XOR2_X1 U1453 ( .A(KEYINPUT57), .B(G2100), .Z(n1872) );
  XOR2_X1 U1454 ( .A(n1656), .B(G2096), .Z(n1871) );
  NAND2_X1 U1455 ( .A1(G860), .A2(n1666), .ZN(G153) );
  INV_X1 U1456 ( .A(n1584), .ZN(n1666) );
  NAND4_X1 U1457 ( .A1(n1873), .A2(G11), .A3(n1874), .A4(n1875), .ZN(G150) );
  NOR3_X1 U1458 ( .A1(n1876), .A2(n1877), .A3(n1878), .ZN(n1875) );
  NOR2_X1 U1459 ( .A1(n1879), .A2(n1880), .ZN(n1878) );
  NOR4_X1 U1460 ( .A1(n1881), .A2(n1882), .A3(n1883), .A4(n1884), .ZN(n1879) );
  XOR2_X1 U1461 ( .A(n1703), .B(G288), .Z(n1884) );
  NAND4_X1 U1462 ( .A1(n1885), .A2(n1886), .A3(n1887), .A4(n1888), .ZN(G288) );
  NAND2_X1 U1463 ( .A1(G49), .A2(n1889), .ZN(n1887) );
  NAND2_X1 U1464 ( .A1(G87), .A2(n1890), .ZN(n1886) );
  NAND2_X1 U1465 ( .A1(G74), .A2(G651), .ZN(n1885) );
  XOR2_X1 U1466 ( .A(n1847), .B(G303), .Z(n1883) );
  NAND4_X1 U1467 ( .A1(n1891), .A2(n1892), .A3(n1893), .A4(n1894), .ZN(G303) );
  NAND2_X1 U1468 ( .A1(G88), .A2(n1895), .ZN(n1894) );
  NAND2_X1 U1469 ( .A1(G75), .A2(n1896), .ZN(n1893) );
  NAND2_X1 U1470 ( .A1(G50), .A2(n1889), .ZN(n1892) );
  NAND2_X1 U1471 ( .A1(G62), .A2(n1897), .ZN(n1891) );
  INV_X1 U1472 ( .A(G1971), .ZN(n1847) );
  XOR2_X1 U1473 ( .A(G1956), .B(n1592), .Z(n1882) );
  INV_X1 U1474 ( .A(G299), .ZN(n1592) );
  NAND4_X1 U1475 ( .A1(n1898), .A2(n1899), .A3(n1900), .A4(n1901), .ZN(G299) );
  NAND2_X1 U1476 ( .A1(G91), .A2(n1895), .ZN(n1901) );
  NAND2_X1 U1477 ( .A1(G78), .A2(n1896), .ZN(n1900) );
  NAND2_X1 U1478 ( .A1(G53), .A2(n1889), .ZN(n1899) );
  NAND2_X1 U1479 ( .A1(G65), .A2(n1897), .ZN(n1898) );
  NAND4_X1 U1480 ( .A1(n1902), .A2(n1903), .A3(n1904), .A4(n1905), .ZN(n1881) );
  XNOR2_X1 U1481 ( .A(G171), .B(n1906), .ZN(n1905) );
  AND4_X1 U1482 ( .A1(n1907), .A2(n1908), .A3(n1909), .A4(n1910), .ZN(G171) );
  NAND2_X1 U1483 ( .A1(G90), .A2(n1895), .ZN(n1910) );
  NAND2_X1 U1484 ( .A1(G77), .A2(n1896), .ZN(n1909) );
  NAND2_X1 U1485 ( .A1(G52), .A2(n1889), .ZN(n1908) );
  NAND2_X1 U1486 ( .A1(G64), .A2(n1897), .ZN(n1907) );
  XOR2_X1 U1487 ( .A(G290), .B(n1729), .Z(n1904) );
  NAND4_X1 U1488 ( .A1(n1911), .A2(n1912), .A3(n1913), .A4(n1914), .ZN(G290) );
  NAND2_X1 U1489 ( .A1(n1889), .A2(n1915), .ZN(n1914) );
  XOR2_X1 U1490 ( .A(KEYINPUT4), .B(G47), .Z(n1915) );
  NAND2_X1 U1491 ( .A1(G85), .A2(n1895), .ZN(n1913) );
  NAND2_X1 U1492 ( .A1(G72), .A2(n1896), .ZN(n1912) );
  NAND2_X1 U1493 ( .A1(G60), .A2(n1897), .ZN(n1911) );
  XOR2_X1 U1494 ( .A(n1590), .B(G1966), .Z(n1903) );
  NAND4_X1 U1495 ( .A1(n1916), .A2(n1917), .A3(n1918), .A4(n1919), .ZN(n1590) );
  NAND2_X1 U1496 ( .A1(G89), .A2(n1895), .ZN(n1919) );
  NAND2_X1 U1497 ( .A1(G76), .A2(n1896), .ZN(n1918) );
  NAND2_X1 U1498 ( .A1(G51), .A2(n1889), .ZN(n1917) );
  NAND2_X1 U1499 ( .A1(G63), .A2(n1897), .ZN(n1916) );
  XOR2_X1 U1500 ( .A(n1584), .B(G1341), .Z(n1902) );
  NOR2_X1 U1501 ( .A1(G16), .A2(n1920), .ZN(n1877) );
  NOR4_X1 U1502 ( .A1(n1921), .A2(n1922), .A3(n1923), .A4(n1924), .ZN(n1920) );
  XOR2_X1 U1503 ( .A(G24), .B(n1769), .Z(n1924) );
  INV_X1 U1504 ( .A(n1729), .ZN(n1769) );
  XNOR2_X1 U1505 ( .A(G1986), .B(KEYINPUT29), .ZN(n1729) );
  XOR2_X1 U1506 ( .A(n1703), .B(G23), .Z(n1923) );
  INV_X1 U1507 ( .A(G1976), .ZN(n1703) );
  XNOR2_X1 U1508 ( .A(G5), .B(n1906), .ZN(n1922) );
  NAND2_X1 U1509 ( .A1(KEYINPUT3), .A2(n1700), .ZN(n1906) );
  INV_X1 U1510 ( .A(G1961), .ZN(n1700) );
  NAND4_X1 U1511 ( .A1(n1925), .A2(n1926), .A3(n1927), .A4(n1928), .ZN(n1921) );
  XOR2_X1 U1512 ( .A(G19), .B(G1341), .Z(n1928) );
  XOR2_X1 U1513 ( .A(G20), .B(G1956), .Z(n1927) );
  XOR2_X1 U1514 ( .A(G21), .B(G1966), .Z(n1926) );
  XOR2_X1 U1515 ( .A(G22), .B(G1971), .Z(n1925) );
  NAND4_X1 U1516 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .ZN(n1876) );
  NAND2_X1 U1517 ( .A1(G29), .A2(n1933), .ZN(n1932) );
  NAND4_X1 U1518 ( .A1(n1934), .A2(n1935), .A3(n1936), .A4(n1656), .ZN(n1933) );
  NAND4_X1 U1519 ( .A1(n1937), .A2(n1938), .A3(n1939), .A4(n1940), .ZN(n1656) );
  NAND2_X1 U1520 ( .A1(G135), .A2(n1941), .ZN(n1940) );
  NAND2_X1 U1521 ( .A1(G99), .A2(n1652), .ZN(n1939) );
  NAND2_X1 U1522 ( .A1(G111), .A2(n1653), .ZN(n1938) );
  NAND2_X1 U1523 ( .A1(G123), .A2(n1650), .ZN(n1937) );
  XOR2_X1 U1524 ( .A(n1630), .B(G2084), .Z(n1936) );
  NAND4_X1 U1525 ( .A1(n1942), .A2(n1943), .A3(n1944), .A4(n1945), .ZN(n1630) );
  NAND3_X1 U1526 ( .A1(n1946), .A2(n1947), .A3(G101), .ZN(n1945) );
  OR2_X1 U1527 ( .A1(n1941), .A2(KEYINPUT47), .ZN(n1947) );
  NAND2_X1 U1528 ( .A1(KEYINPUT47), .A2(n1948), .ZN(n1946) );
  NAND2_X1 U1529 ( .A1(G137), .A2(n1941), .ZN(n1944) );
  NAND2_X1 U1530 ( .A1(G113), .A2(n1653), .ZN(n1943) );
  NAND2_X1 U1531 ( .A1(G125), .A2(n1650), .ZN(n1942) );
  XOR2_X1 U1532 ( .A(n1629), .B(G2090), .Z(n1935) );
  NAND4_X1 U1533 ( .A1(n1949), .A2(n1950), .A3(n1951), .A4(n1952), .ZN(n1629) );
  NAND2_X1 U1534 ( .A1(G136), .A2(n1941), .ZN(n1952) );
  NAND2_X1 U1535 ( .A1(G100), .A2(n1652), .ZN(n1951) );
  NAND2_X1 U1536 ( .A1(G112), .A2(n1653), .ZN(n1950) );
  NAND2_X1 U1537 ( .A1(G124), .A2(n1650), .ZN(n1949) );
  XNOR2_X1 U1538 ( .A(G164), .B(G2078), .ZN(n1934) );
  AND4_X1 U1539 ( .A1(n1953), .A2(n1954), .A3(n1955), .A4(n1956), .ZN(G164) );
  NAND3_X1 U1540 ( .A1(n1957), .A2(n1958), .A3(G114), .ZN(n1956) );
  OR2_X1 U1541 ( .A1(n1653), .A2(KEYINPUT2), .ZN(n1958) );
  NAND2_X1 U1542 ( .A1(KEYINPUT2), .A2(n1948), .ZN(n1957) );
  NAND2_X1 U1543 ( .A1(G138), .A2(n1941), .ZN(n1955) );
  NAND2_X1 U1544 ( .A1(G102), .A2(n1652), .ZN(n1954) );
  NAND2_X1 U1545 ( .A1(G126), .A2(n1650), .ZN(n1953) );
  NAND2_X1 U1546 ( .A1(n1959), .A2(n1960), .ZN(n1931) );
  NAND4_X1 U1547 ( .A1(G28), .A2(n1961), .A3(n1962), .A4(n1963), .ZN(n1959) );
  XOR2_X1 U1548 ( .A(G27), .B(G2078), .Z(n1963) );
  XOR2_X1 U1549 ( .A(G34), .B(G2084), .Z(n1962) );
  XOR2_X1 U1550 ( .A(G35), .B(G2090), .Z(n1961) );
  NAND2_X1 U1551 ( .A1(n1964), .A2(n1965), .ZN(n1930) );
  NAND4_X1 U1552 ( .A1(n1966), .A2(n1967), .A3(n1968), .A4(n1969), .ZN(n1965) );
  XOR2_X1 U1553 ( .A(G25), .B(G1991), .Z(n1969) );
  XOR2_X1 U1554 ( .A(G32), .B(G1996), .Z(n1968) );
  XOR2_X1 U1555 ( .A(G33), .B(G2072), .Z(n1967) );
  XOR2_X1 U1556 ( .A(n1970), .B(G26), .Z(n1966) );
  INV_X1 U1557 ( .A(n1971), .ZN(n1964) );
  NAND2_X1 U1558 ( .A1(n1971), .A2(n1972), .ZN(n1929) );
  NAND4_X1 U1559 ( .A1(n1973), .A2(n1974), .A3(n1975), .A4(n1976), .ZN(n1972) );
  XOR2_X1 U1560 ( .A(n1970), .B(n1640), .Z(n1976) );
  NAND4_X1 U1561 ( .A1(n1977), .A2(n1978), .A3(n1979), .A4(n1980), .ZN(n1640) );
  NAND2_X1 U1562 ( .A1(G140), .A2(n1941), .ZN(n1980) );
  NAND2_X1 U1563 ( .A1(G104), .A2(n1652), .ZN(n1979) );
  NAND2_X1 U1564 ( .A1(G116), .A2(n1653), .ZN(n1978) );
  NAND2_X1 U1565 ( .A1(G128), .A2(n1650), .ZN(n1977) );
  NAND2_X1 U1566 ( .A1(KEYINPUT17), .A2(n1617), .ZN(n1970) );
  INV_X1 U1567 ( .A(G2067), .ZN(n1617) );
  NOR2_X1 U1568 ( .A1(n1860), .A2(n1981), .ZN(n1975) );
  NOR2_X1 U1569 ( .A1(n1856), .A2(n1861), .ZN(n1981) );
  INV_X1 U1570 ( .A(n1768), .ZN(n1860) );
  NAND2_X1 U1571 ( .A1(n1856), .A2(n1861), .ZN(n1768) );
  INV_X1 U1572 ( .A(G1991), .ZN(n1861) );
  INV_X1 U1573 ( .A(n1642), .ZN(n1856) );
  NAND4_X1 U1574 ( .A1(n1982), .A2(n1983), .A3(n1984), .A4(n1985), .ZN(n1642) );
  NAND2_X1 U1575 ( .A1(G131), .A2(n1941), .ZN(n1985) );
  NAND2_X1 U1576 ( .A1(G95), .A2(n1652), .ZN(n1984) );
  NAND2_X1 U1577 ( .A1(G107), .A2(n1653), .ZN(n1983) );
  NAND2_X1 U1578 ( .A1(G119), .A2(n1650), .ZN(n1982) );
  XOR2_X1 U1579 ( .A(n1654), .B(G2072), .Z(n1974) );
  NAND4_X1 U1580 ( .A1(n1986), .A2(n1987), .A3(n1988), .A4(n1989), .ZN(n1654) );
  NAND2_X1 U1581 ( .A1(G139), .A2(n1941), .ZN(n1989) );
  NAND2_X1 U1582 ( .A1(G103), .A2(n1652), .ZN(n1988) );
  NAND2_X1 U1583 ( .A1(G115), .A2(n1653), .ZN(n1987) );
  NAND2_X1 U1584 ( .A1(G127), .A2(n1650), .ZN(n1986) );
  XOR2_X1 U1585 ( .A(n1721), .B(G1996), .Z(n1973) );
  NAND4_X1 U1586 ( .A1(n1990), .A2(n1991), .A3(n1992), .A4(n1993), .ZN(n1721) );
  NAND2_X1 U1587 ( .A1(G141), .A2(n1941), .ZN(n1993) );
  INV_X1 U1588 ( .A(n1651), .ZN(n1941) );
  NAND2_X1 U1589 ( .A1(n1994), .A2(n1995), .ZN(n1651) );
  NAND2_X1 U1590 ( .A1(G105), .A2(n1652), .ZN(n1992) );
  INV_X1 U1591 ( .A(n1948), .ZN(n1652) );
  NAND2_X1 U1592 ( .A1(G2104), .A2(n1995), .ZN(n1948) );
  NAND2_X1 U1593 ( .A1(G117), .A2(n1653), .ZN(n1991) );
  NOR2_X1 U1594 ( .A1(n1995), .A2(n1994), .ZN(n1653) );
  INV_X1 U1595 ( .A(G2104), .ZN(n1994) );
  NAND2_X1 U1596 ( .A1(G129), .A2(n1650), .ZN(n1990) );
  NOR2_X1 U1597 ( .A1(n1995), .A2(G2104), .ZN(n1650) );
  INV_X1 U1598 ( .A(G2105), .ZN(n1995) );
  XOR2_X1 U1599 ( .A(n1960), .B(KEYINPUT21), .Z(n1971) );
  INV_X1 U1600 ( .A(G29), .ZN(n1960) );
  XNOR2_X1 U1601 ( .A(n1996), .B(n1803), .ZN(n1874) );
  XNOR2_X1 U1602 ( .A(G1981), .B(KEYINPUT12), .ZN(n1803) );
  NAND2_X1 U1603 ( .A1(n1997), .A2(n1998), .ZN(n1996) );
  NAND2_X1 U1604 ( .A1(G6), .A2(n1880), .ZN(n1998) );
  XOR2_X1 U1605 ( .A(KEYINPUT31), .B(n1999), .Z(n1997) );
  NOR2_X1 U1606 ( .A1(n1673), .A2(n1880), .ZN(n1999) );
  INV_X1 U1607 ( .A(G305), .ZN(n1673) );
  NAND4_X1 U1608 ( .A1(n2000), .A2(n2001), .A3(n2002), .A4(n2003), .ZN(G305) );
  NAND2_X1 U1609 ( .A1(G86), .A2(n1895), .ZN(n2003) );
  NAND2_X1 U1610 ( .A1(G73), .A2(n1896), .ZN(n2002) );
  NAND2_X1 U1611 ( .A1(G48), .A2(n1889), .ZN(n2001) );
  NAND2_X1 U1612 ( .A1(G61), .A2(n1897), .ZN(n2000) );
  XOR2_X1 U1613 ( .A(n2004), .B(G1348), .Z(n1873) );
  NAND2_X1 U1614 ( .A1(n2005), .A2(n2006), .ZN(n2004) );
  NAND2_X1 U1615 ( .A1(G4), .A2(n1880), .ZN(n2006) );
  INV_X1 U1616 ( .A(G16), .ZN(n1880) );
  XOR2_X1 U1617 ( .A(n2007), .B(KEYINPUT38), .Z(n2005) );
  NAND2_X1 U1618 ( .A1(G16), .A2(n1587), .ZN(n2007) );
  NAND2_X1 U1619 ( .A1(n1668), .A2(n2008), .ZN(G148) );
  NAND2_X1 U1620 ( .A1(n1575), .A2(n2009), .ZN(n2008) );
  NAND2_X1 U1621 ( .A1(n2010), .A2(n2011), .ZN(G145) );
  NAND2_X1 U1622 ( .A1(G860), .A2(n2012), .ZN(n2011) );
  NAND2_X1 U1623 ( .A1(n1667), .A2(n2013), .ZN(n2012) );
  NAND2_X1 U1624 ( .A1(n2014), .A2(n2015), .ZN(n2013) );
  INV_X1 U1625 ( .A(KEYINPUT11), .ZN(n2015) );
  NAND3_X1 U1626 ( .A1(n2016), .A2(n2017), .A3(KEYINPUT11), .ZN(n2010) );
  NAND2_X1 U1627 ( .A1(n2014), .A2(n2018), .ZN(n2017) );
  NAND2_X1 U1628 ( .A1(n1667), .A2(n2009), .ZN(n2018) );
  INV_X1 U1629 ( .A(G860), .ZN(n2009) );
  INV_X1 U1630 ( .A(n1565), .ZN(n1667) );
  OR2_X1 U1631 ( .A1(n2014), .A2(n1565), .ZN(n2016) );
  NAND4_X1 U1632 ( .A1(n2019), .A2(n2020), .A3(n2021), .A4(n2022), .ZN(n1565) );
  NAND2_X1 U1633 ( .A1(G93), .A2(n1895), .ZN(n2022) );
  NAND2_X1 U1634 ( .A1(G80), .A2(n1896), .ZN(n2021) );
  NAND2_X1 U1635 ( .A1(G55), .A2(n1889), .ZN(n2020) );
  NAND2_X1 U1636 ( .A1(G67), .A2(n1897), .ZN(n2019) );
  XNOR2_X1 U1637 ( .A(n2023), .B(n2024), .ZN(n2014) );
  NOR3_X1 U1638 ( .A1(n1826), .A2(n2025), .A3(n2026), .ZN(n2024) );
  NOR2_X1 U1639 ( .A1(n2027), .A2(n1819), .ZN(n2026) );
  NAND2_X1 U1640 ( .A1(n1587), .A2(n1584), .ZN(n1819) );
  AND2_X1 U1641 ( .A1(n1668), .A2(n2027), .ZN(n2025) );
  XNOR2_X1 U1642 ( .A(KEYINPUT46), .B(KEYINPUT20), .ZN(n2027) );
  NOR2_X1 U1643 ( .A1(n1587), .A2(n1584), .ZN(n1826) );
  NAND4_X1 U1644 ( .A1(n2028), .A2(n2029), .A3(n2030), .A4(n2031), .ZN(n1584) );
  NAND2_X1 U1645 ( .A1(G81), .A2(n1895), .ZN(n2031) );
  NAND2_X1 U1646 ( .A1(G68), .A2(n1896), .ZN(n2030) );
  NAND2_X1 U1647 ( .A1(G43), .A2(n1889), .ZN(n2029) );
  NAND2_X1 U1648 ( .A1(G56), .A2(n1897), .ZN(n2028) );
  NAND2_X1 U1649 ( .A1(KEYINPUT26), .A2(n1577), .ZN(n2023) );
  INV_X1 U1650 ( .A(n1575), .ZN(n1577) );
  NAND2_X1 U1651 ( .A1(n2032), .A2(n1668), .ZN(n1575) );
  INV_X1 U1652 ( .A(n1587), .ZN(n1668) );
  NAND4_X1 U1653 ( .A1(n2033), .A2(n2034), .A3(n2035), .A4(n2036), .ZN(n1587) );
  NAND2_X1 U1654 ( .A1(G92), .A2(n1895), .ZN(n2036) );
  NOR2_X1 U1655 ( .A1(G543), .A2(G651), .ZN(n1895) );
  NAND2_X1 U1656 ( .A1(G79), .A2(n1896), .ZN(n2035) );
  AND2_X1 U1657 ( .A1(G651), .A2(G543), .ZN(n1896) );
  NAND2_X1 U1658 ( .A1(G54), .A2(n1889), .ZN(n2034) );
  NOR2_X1 U1659 ( .A1(n1890), .A2(G651), .ZN(n1889) );
  NAND2_X1 U1660 ( .A1(G66), .A2(n1897), .ZN(n2033) );
  INV_X1 U1661 ( .A(n1888), .ZN(n1897) );
  NAND2_X1 U1662 ( .A1(G651), .A2(n1890), .ZN(n1888) );
  INV_X1 U1663 ( .A(G543), .ZN(n1890) );
  XNOR2_X1 U1664 ( .A(KEYINPUT15), .B(G559), .ZN(n2032) );
endmodule

