//Key = 0010000101010100111100101001000011111001010011100111001000101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291;

NAND2_X1 U711 ( .A1(n980), .A2(n981), .ZN(G9) );
NAND2_X1 U712 ( .A1(G107), .A2(n982), .ZN(n981) );
XOR2_X1 U713 ( .A(n983), .B(KEYINPUT14), .Z(n980) );
OR2_X1 U714 ( .A1(n982), .A2(G107), .ZN(n983) );
NOR2_X1 U715 ( .A1(n984), .A2(n985), .ZN(G75) );
NOR4_X1 U716 ( .A1(n986), .A2(n987), .A3(n988), .A4(n989), .ZN(n985) );
XOR2_X1 U717 ( .A(n990), .B(KEYINPUT51), .Z(n989) );
NAND3_X1 U718 ( .A1(n991), .A2(n992), .A3(n993), .ZN(n990) );
NOR2_X1 U719 ( .A1(n994), .A2(n995), .ZN(n988) );
INV_X1 U720 ( .A(n996), .ZN(n994) );
NAND4_X1 U721 ( .A1(n997), .A2(n998), .A3(n999), .A4(n1000), .ZN(n986) );
NAND3_X1 U722 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n998) );
XOR2_X1 U723 ( .A(n995), .B(KEYINPUT60), .Z(n1003) );
NAND3_X1 U724 ( .A1(n1004), .A2(n1005), .A3(n991), .ZN(n995) );
INV_X1 U725 ( .A(n1006), .ZN(n1004) );
NAND2_X1 U726 ( .A1(n993), .A2(n1007), .ZN(n997) );
NAND2_X1 U727 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND2_X1 U728 ( .A1(n991), .A2(n1010), .ZN(n1009) );
AND2_X1 U729 ( .A1(n1011), .A2(n1012), .ZN(n991) );
NAND2_X1 U730 ( .A1(n1005), .A2(n1013), .ZN(n1008) );
NAND2_X1 U731 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND2_X1 U732 ( .A1(n1016), .A2(n1012), .ZN(n1015) );
XNOR2_X1 U733 ( .A(n1017), .B(n1018), .ZN(n1016) );
NOR2_X1 U734 ( .A1(KEYINPUT26), .A2(n1019), .ZN(n1018) );
NAND2_X1 U735 ( .A1(n1011), .A2(n1020), .ZN(n1014) );
NAND2_X1 U736 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U737 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR3_X1 U738 ( .A1(n1025), .A2(n1001), .A3(n1006), .ZN(n993) );
NOR3_X1 U739 ( .A1(n1026), .A2(G953), .A3(G952), .ZN(n984) );
INV_X1 U740 ( .A(n999), .ZN(n1026) );
NAND4_X1 U741 ( .A1(n1027), .A2(n1011), .A3(n1028), .A4(n1029), .ZN(n999) );
NOR4_X1 U742 ( .A1(n1001), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1029) );
AND2_X1 U743 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U744 ( .A1(n1035), .A2(n1036), .ZN(n1028) );
XNOR2_X1 U745 ( .A(n1037), .B(KEYINPUT4), .ZN(n1027) );
XOR2_X1 U746 ( .A(n1038), .B(n1039), .Z(G72) );
NOR3_X1 U747 ( .A1(n1000), .A2(KEYINPUT31), .A3(n1040), .ZN(n1039) );
NOR2_X1 U748 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U749 ( .A1(n1043), .A2(n1044), .ZN(n1038) );
NAND2_X1 U750 ( .A1(n1045), .A2(n1000), .ZN(n1044) );
XOR2_X1 U751 ( .A(n1046), .B(n1047), .Z(n1045) );
NAND2_X1 U752 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NAND3_X1 U753 ( .A1(n1047), .A2(G900), .A3(G953), .ZN(n1043) );
NOR2_X1 U754 ( .A1(KEYINPUT29), .A2(n1050), .ZN(n1047) );
XOR2_X1 U755 ( .A(KEYINPUT33), .B(n1051), .Z(n1050) );
NOR2_X1 U756 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XOR2_X1 U757 ( .A(n1054), .B(KEYINPUT63), .Z(n1053) );
NAND3_X1 U758 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
OR2_X1 U759 ( .A1(n1058), .A2(G125), .ZN(n1055) );
NOR2_X1 U760 ( .A1(n1059), .A2(n1060), .ZN(n1052) );
XNOR2_X1 U761 ( .A(KEYINPUT58), .B(n1057), .ZN(n1060) );
XOR2_X1 U762 ( .A(n1061), .B(n1062), .Z(n1057) );
XNOR2_X1 U763 ( .A(n1063), .B(n1064), .ZN(n1061) );
NAND2_X1 U764 ( .A1(KEYINPUT36), .A2(n1065), .ZN(n1063) );
NOR2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1059) );
NOR2_X1 U766 ( .A1(G125), .A2(n1058), .ZN(n1067) );
XNOR2_X1 U767 ( .A(n1068), .B(G140), .ZN(n1058) );
XNOR2_X1 U768 ( .A(KEYINPUT9), .B(KEYINPUT27), .ZN(n1068) );
XOR2_X1 U769 ( .A(n1069), .B(n1070), .Z(G69) );
NOR2_X1 U770 ( .A1(G953), .A2(n1071), .ZN(n1070) );
XOR2_X1 U771 ( .A(KEYINPUT48), .B(n1072), .Z(n1071) );
NAND2_X1 U772 ( .A1(n1073), .A2(n1074), .ZN(n1069) );
NAND2_X1 U773 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U774 ( .A1(G953), .A2(n1077), .ZN(n1076) );
NAND2_X1 U775 ( .A1(G953), .A2(n1078), .ZN(n1073) );
NAND2_X1 U776 ( .A1(G898), .A2(n1079), .ZN(n1078) );
OR2_X1 U777 ( .A1(n1075), .A2(G224), .ZN(n1079) );
XNOR2_X1 U778 ( .A(n1080), .B(n1081), .ZN(n1075) );
XNOR2_X1 U779 ( .A(KEYINPUT40), .B(n1082), .ZN(n1080) );
NOR2_X1 U780 ( .A1(KEYINPUT25), .A2(n1083), .ZN(n1082) );
XOR2_X1 U781 ( .A(n1084), .B(n1085), .Z(n1083) );
NOR2_X1 U782 ( .A1(KEYINPUT59), .A2(n1086), .ZN(n1084) );
NOR2_X1 U783 ( .A1(n1087), .A2(n1088), .ZN(G66) );
XOR2_X1 U784 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U785 ( .A1(n1091), .A2(KEYINPUT57), .ZN(n1089) );
NOR2_X1 U786 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR2_X1 U787 ( .A1(n1087), .A2(n1094), .ZN(G63) );
XNOR2_X1 U788 ( .A(n1095), .B(n1096), .ZN(n1094) );
NOR2_X1 U789 ( .A1(n1097), .A2(n1093), .ZN(n1096) );
NOR2_X1 U790 ( .A1(n1087), .A2(n1098), .ZN(G60) );
NOR2_X1 U791 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U792 ( .A(KEYINPUT8), .B(n1101), .Z(n1100) );
NOR2_X1 U793 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U794 ( .A(KEYINPUT42), .B(n1104), .Z(n1103) );
AND2_X1 U795 ( .A1(n1102), .A2(n1104), .ZN(n1099) );
NOR2_X1 U796 ( .A1(n1093), .A2(n1105), .ZN(n1104) );
INV_X1 U797 ( .A(G475), .ZN(n1105) );
XOR2_X1 U798 ( .A(n1106), .B(n1107), .Z(G6) );
NOR2_X1 U799 ( .A1(KEYINPUT53), .A2(n1108), .ZN(n1107) );
NOR2_X1 U800 ( .A1(n1087), .A2(n1109), .ZN(G57) );
XOR2_X1 U801 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U802 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U803 ( .A(n1114), .B(n1115), .Z(n1110) );
NOR2_X1 U804 ( .A1(n1116), .A2(n1093), .ZN(n1115) );
XOR2_X1 U805 ( .A(n1117), .B(KEYINPUT17), .Z(n1114) );
NOR2_X1 U806 ( .A1(n1087), .A2(n1118), .ZN(G54) );
XOR2_X1 U807 ( .A(n1119), .B(n1120), .Z(n1118) );
NOR2_X1 U808 ( .A1(n1121), .A2(n1093), .ZN(n1120) );
NOR2_X1 U809 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
XOR2_X1 U810 ( .A(KEYINPUT15), .B(n1124), .Z(n1123) );
NOR2_X1 U811 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
AND2_X1 U812 ( .A1(n1126), .A2(n1125), .ZN(n1122) );
XNOR2_X1 U813 ( .A(n1127), .B(n1128), .ZN(n1125) );
XOR2_X1 U814 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U815 ( .A1(n1131), .A2(KEYINPUT10), .ZN(n1129) );
XNOR2_X1 U816 ( .A(KEYINPUT61), .B(KEYINPUT56), .ZN(n1127) );
XNOR2_X1 U817 ( .A(n1132), .B(n1133), .ZN(n1126) );
NAND2_X1 U818 ( .A1(KEYINPUT35), .A2(n1062), .ZN(n1132) );
NOR2_X1 U819 ( .A1(n1087), .A2(n1134), .ZN(G51) );
XOR2_X1 U820 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U821 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U822 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
INV_X1 U823 ( .A(n1141), .ZN(n1140) );
XOR2_X1 U824 ( .A(KEYINPUT32), .B(n1142), .Z(n1139) );
NOR2_X1 U825 ( .A1(n1141), .A2(n1143), .ZN(n1137) );
XOR2_X1 U826 ( .A(KEYINPUT20), .B(n1142), .Z(n1143) );
XNOR2_X1 U827 ( .A(n1144), .B(n1145), .ZN(n1135) );
NOR2_X1 U828 ( .A1(n1146), .A2(n1093), .ZN(n1145) );
NAND2_X1 U829 ( .A1(G902), .A2(n987), .ZN(n1093) );
NAND3_X1 U830 ( .A1(n1072), .A2(n1048), .A3(n1147), .ZN(n987) );
XOR2_X1 U831 ( .A(n1049), .B(KEYINPUT55), .Z(n1147) );
NAND2_X1 U832 ( .A1(n1148), .A2(n996), .ZN(n1049) );
XNOR2_X1 U833 ( .A(n1149), .B(KEYINPUT34), .ZN(n1148) );
AND4_X1 U834 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1048) );
AND4_X1 U835 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1153) );
NAND2_X1 U836 ( .A1(n1158), .A2(n992), .ZN(n1152) );
AND4_X1 U837 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1072) );
AND4_X1 U838 ( .A1(n982), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1162) );
NAND3_X1 U839 ( .A1(n1010), .A2(n1012), .A3(n1166), .ZN(n982) );
NOR2_X1 U840 ( .A1(n1167), .A2(n1106), .ZN(n1161) );
AND3_X1 U841 ( .A1(n1166), .A2(n1012), .A3(n992), .ZN(n1106) );
NOR3_X1 U842 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1167) );
INV_X1 U843 ( .A(n1010), .ZN(n1169) );
XNOR2_X1 U844 ( .A(KEYINPUT49), .B(n1021), .ZN(n1168) );
NAND3_X1 U845 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1160) );
INV_X1 U846 ( .A(n1174), .ZN(n1173) );
NAND2_X1 U847 ( .A1(KEYINPUT50), .A2(n1170), .ZN(n1172) );
NAND2_X1 U848 ( .A1(n1175), .A2(n1176), .ZN(n1171) );
INV_X1 U849 ( .A(KEYINPUT50), .ZN(n1176) );
NAND2_X1 U850 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
INV_X1 U851 ( .A(n1011), .ZN(n1178) );
NOR2_X1 U852 ( .A1(n1000), .A2(G952), .ZN(n1087) );
XOR2_X1 U853 ( .A(G146), .B(n1179), .Z(G48) );
NOR2_X1 U854 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U855 ( .A(KEYINPUT16), .B(n992), .Z(n1181) );
XNOR2_X1 U856 ( .A(G143), .B(n1150), .ZN(G45) );
NAND4_X1 U857 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n996), .ZN(n1150) );
NOR2_X1 U858 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XNOR2_X1 U859 ( .A(G140), .B(n1151), .ZN(G42) );
NAND4_X1 U860 ( .A1(n1187), .A2(n992), .A3(n1024), .A4(n1023), .ZN(n1151) );
XNOR2_X1 U861 ( .A(G137), .B(n1157), .ZN(G39) );
NAND3_X1 U862 ( .A1(n1188), .A2(n1036), .A3(n1187), .ZN(n1157) );
XOR2_X1 U863 ( .A(n1156), .B(n1189), .Z(G36) );
NAND2_X1 U864 ( .A1(KEYINPUT2), .A2(G134), .ZN(n1189) );
NAND3_X1 U865 ( .A1(n1183), .A2(n1010), .A3(n1187), .ZN(n1156) );
XNOR2_X1 U866 ( .A(G131), .B(n1155), .ZN(G33) );
NAND3_X1 U867 ( .A1(n992), .A2(n1183), .A3(n1187), .ZN(n1155) );
AND3_X1 U868 ( .A1(n1182), .A2(n1190), .A3(n1002), .ZN(n1187) );
XOR2_X1 U869 ( .A(n1154), .B(n1191), .Z(G30) );
NAND2_X1 U870 ( .A1(KEYINPUT18), .A2(G128), .ZN(n1191) );
NAND2_X1 U871 ( .A1(n1158), .A2(n1010), .ZN(n1154) );
INV_X1 U872 ( .A(n1180), .ZN(n1158) );
NAND4_X1 U873 ( .A1(n1023), .A2(n1182), .A3(n996), .A4(n1036), .ZN(n1180) );
AND3_X1 U874 ( .A1(n1192), .A2(n1193), .A3(n1019), .ZN(n1182) );
XNOR2_X1 U875 ( .A(G101), .B(n1165), .ZN(G3) );
NAND3_X1 U876 ( .A1(n1005), .A2(n1166), .A3(n1183), .ZN(n1165) );
XNOR2_X1 U877 ( .A(G125), .B(n1194), .ZN(G27) );
NAND3_X1 U878 ( .A1(n1149), .A2(n996), .A3(KEYINPUT22), .ZN(n1194) );
AND4_X1 U879 ( .A1(n1024), .A2(n1192), .A3(n1011), .A4(n1195), .ZN(n1149) );
AND2_X1 U880 ( .A1(n992), .A2(n1023), .ZN(n1195) );
NAND2_X1 U881 ( .A1(n1006), .A2(n1196), .ZN(n1192) );
NAND4_X1 U882 ( .A1(G953), .A2(G902), .A3(n1197), .A4(n1042), .ZN(n1196) );
INV_X1 U883 ( .A(G900), .ZN(n1042) );
XNOR2_X1 U884 ( .A(n1198), .B(n1199), .ZN(G24) );
NOR2_X1 U885 ( .A1(n1170), .A2(n1174), .ZN(n1199) );
NAND3_X1 U886 ( .A1(n1037), .A2(n1200), .A3(n1012), .ZN(n1174) );
NOR2_X1 U887 ( .A1(n1036), .A2(n1023), .ZN(n1012) );
XNOR2_X1 U888 ( .A(G119), .B(n1164), .ZN(G21) );
OR3_X1 U889 ( .A1(n1201), .A2(n1024), .A3(n1170), .ZN(n1164) );
XNOR2_X1 U890 ( .A(G116), .B(n1202), .ZN(G18) );
NAND2_X1 U891 ( .A1(n1203), .A2(n1010), .ZN(n1202) );
NOR2_X1 U892 ( .A1(n1037), .A2(n1185), .ZN(n1010) );
INV_X1 U893 ( .A(n1200), .ZN(n1185) );
XNOR2_X1 U894 ( .A(n1204), .B(n1205), .ZN(G15) );
NOR2_X1 U895 ( .A1(KEYINPUT3), .A2(n1159), .ZN(n1205) );
NAND2_X1 U896 ( .A1(n1203), .A2(n992), .ZN(n1159) );
NOR2_X1 U897 ( .A1(n1200), .A2(n1186), .ZN(n992) );
NOR2_X1 U898 ( .A1(n1021), .A2(n1170), .ZN(n1203) );
NAND2_X1 U899 ( .A1(n1011), .A2(n1177), .ZN(n1170) );
NOR2_X1 U900 ( .A1(n1019), .A2(n1017), .ZN(n1011) );
INV_X1 U901 ( .A(n1193), .ZN(n1017) );
INV_X1 U902 ( .A(n1183), .ZN(n1021) );
NOR2_X1 U903 ( .A1(n1023), .A2(n1024), .ZN(n1183) );
XOR2_X1 U904 ( .A(n1163), .B(n1206), .Z(G12) );
XNOR2_X1 U905 ( .A(G110), .B(KEYINPUT0), .ZN(n1206) );
NAND3_X1 U906 ( .A1(n1024), .A2(n1166), .A3(n1188), .ZN(n1163) );
INV_X1 U907 ( .A(n1201), .ZN(n1188) );
NAND2_X1 U908 ( .A1(n1005), .A2(n1023), .ZN(n1201) );
XNOR2_X1 U909 ( .A(n1035), .B(KEYINPUT45), .ZN(n1023) );
XOR2_X1 U910 ( .A(n1207), .B(n1092), .Z(n1035) );
NAND2_X1 U911 ( .A1(G217), .A2(n1208), .ZN(n1092) );
NAND2_X1 U912 ( .A1(n1090), .A2(n1209), .ZN(n1207) );
XNOR2_X1 U913 ( .A(n1210), .B(n1211), .ZN(n1090) );
XOR2_X1 U914 ( .A(n1212), .B(n1213), .Z(n1211) );
XNOR2_X1 U915 ( .A(n1214), .B(G110), .ZN(n1213) );
INV_X1 U916 ( .A(G119), .ZN(n1214) );
XOR2_X1 U917 ( .A(G146), .B(G137), .Z(n1212) );
XOR2_X1 U918 ( .A(n1215), .B(n1216), .Z(n1210) );
XOR2_X1 U919 ( .A(n1217), .B(n1218), .Z(n1216) );
NOR2_X1 U920 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
INV_X1 U921 ( .A(G221), .ZN(n1219) );
NOR2_X1 U922 ( .A1(KEYINPUT21), .A2(n1221), .ZN(n1217) );
NOR4_X1 U923 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1221) );
AND2_X1 U924 ( .A1(KEYINPUT41), .A2(n1066), .ZN(n1225) );
NOR2_X1 U925 ( .A1(KEYINPUT41), .A2(G140), .ZN(n1224) );
AND2_X1 U926 ( .A1(KEYINPUT7), .A2(n1226), .ZN(n1223) );
NOR2_X1 U927 ( .A1(KEYINPUT7), .A2(n1227), .ZN(n1222) );
INV_X1 U928 ( .A(G125), .ZN(n1227) );
NAND2_X1 U929 ( .A1(KEYINPUT13), .A2(n1228), .ZN(n1215) );
NOR2_X1 U930 ( .A1(n1200), .A2(n1037), .ZN(n1005) );
INV_X1 U931 ( .A(n1186), .ZN(n1037) );
XOR2_X1 U932 ( .A(n1229), .B(G475), .Z(n1186) );
OR2_X1 U933 ( .A1(n1102), .A2(G902), .ZN(n1229) );
XOR2_X1 U934 ( .A(n1230), .B(n1231), .Z(n1102) );
XOR2_X1 U935 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U936 ( .A(n1234), .B(n1235), .Z(n1233) );
NOR3_X1 U937 ( .A1(n1226), .A2(KEYINPUT6), .A3(n1066), .ZN(n1235) );
INV_X1 U938 ( .A(n1056), .ZN(n1066) );
NAND2_X1 U939 ( .A1(G140), .A2(G125), .ZN(n1056) );
NOR2_X1 U940 ( .A1(G140), .A2(G125), .ZN(n1226) );
NAND2_X1 U941 ( .A1(n1236), .A2(G214), .ZN(n1234) );
XNOR2_X1 U942 ( .A(G104), .B(G113), .ZN(n1232) );
XOR2_X1 U943 ( .A(n1237), .B(n1238), .Z(n1230) );
XNOR2_X1 U944 ( .A(n1064), .B(G122), .ZN(n1238) );
INV_X1 U945 ( .A(G131), .ZN(n1064) );
XNOR2_X1 U946 ( .A(G143), .B(G146), .ZN(n1237) );
XOR2_X1 U947 ( .A(n1032), .B(KEYINPUT1), .Z(n1200) );
XOR2_X1 U948 ( .A(n1239), .B(n1097), .Z(n1032) );
INV_X1 U949 ( .A(G478), .ZN(n1097) );
NAND2_X1 U950 ( .A1(n1095), .A2(n1209), .ZN(n1239) );
XNOR2_X1 U951 ( .A(n1240), .B(n1241), .ZN(n1095) );
NOR2_X1 U952 ( .A1(n1220), .A2(n1242), .ZN(n1241) );
INV_X1 U953 ( .A(G217), .ZN(n1242) );
NAND2_X1 U954 ( .A1(G234), .A2(n1000), .ZN(n1220) );
NAND2_X1 U955 ( .A1(KEYINPUT39), .A2(n1243), .ZN(n1240) );
NAND2_X1 U956 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
NAND2_X1 U957 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XNOR2_X1 U958 ( .A(n1248), .B(n1249), .ZN(n1247) );
XNOR2_X1 U959 ( .A(G134), .B(n1250), .ZN(n1246) );
XOR2_X1 U960 ( .A(n1251), .B(KEYINPUT62), .Z(n1244) );
NAND2_X1 U961 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
XOR2_X1 U962 ( .A(G134), .B(n1250), .Z(n1253) );
XOR2_X1 U963 ( .A(n1248), .B(n1249), .Z(n1252) );
XNOR2_X1 U964 ( .A(G116), .B(n1198), .ZN(n1249) );
NAND2_X1 U965 ( .A1(KEYINPUT11), .A2(G107), .ZN(n1248) );
AND3_X1 U966 ( .A1(n1019), .A2(n1193), .A3(n1177), .ZN(n1166) );
AND2_X1 U967 ( .A1(n996), .A2(n1254), .ZN(n1177) );
NAND2_X1 U968 ( .A1(n1255), .A2(n1006), .ZN(n1254) );
NAND3_X1 U969 ( .A1(n1197), .A2(n1000), .A3(G952), .ZN(n1006) );
INV_X1 U970 ( .A(G953), .ZN(n1000) );
NAND4_X1 U971 ( .A1(G953), .A2(G902), .A3(n1197), .A4(n1256), .ZN(n1255) );
INV_X1 U972 ( .A(G898), .ZN(n1256) );
NAND2_X1 U973 ( .A1(G237), .A2(n1257), .ZN(n1197) );
XOR2_X1 U974 ( .A(KEYINPUT5), .B(G234), .Z(n1257) );
NOR2_X1 U975 ( .A1(n1001), .A2(n1002), .ZN(n996) );
INV_X1 U976 ( .A(n1025), .ZN(n1002) );
NAND3_X1 U977 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1025) );
INV_X1 U978 ( .A(n1030), .ZN(n1260) );
NOR2_X1 U979 ( .A1(n1033), .A2(n1034), .ZN(n1030) );
NAND3_X1 U980 ( .A1(KEYINPUT54), .A2(n1034), .A3(n1033), .ZN(n1259) );
INV_X1 U981 ( .A(n1146), .ZN(n1034) );
NAND2_X1 U982 ( .A1(G210), .A2(n1261), .ZN(n1146) );
OR2_X1 U983 ( .A1(n1033), .A2(KEYINPUT54), .ZN(n1258) );
NAND2_X1 U984 ( .A1(n1262), .A2(n1209), .ZN(n1033) );
XOR2_X1 U985 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U986 ( .A(n1142), .B(n1265), .ZN(n1264) );
XNOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT38), .ZN(n1265) );
NOR2_X1 U988 ( .A1(n1077), .A2(G953), .ZN(n1142) );
INV_X1 U989 ( .A(G224), .ZN(n1077) );
XNOR2_X1 U990 ( .A(n1141), .B(n1144), .ZN(n1263) );
XNOR2_X1 U991 ( .A(n1086), .B(n1266), .ZN(n1144) );
XOR2_X1 U992 ( .A(n1085), .B(n1081), .Z(n1266) );
XOR2_X1 U993 ( .A(G110), .B(n1267), .Z(n1081) );
NOR2_X1 U994 ( .A1(KEYINPUT30), .A2(n1198), .ZN(n1267) );
INV_X1 U995 ( .A(G122), .ZN(n1198) );
XNOR2_X1 U996 ( .A(n1268), .B(n1269), .ZN(n1085) );
NOR2_X1 U997 ( .A1(G101), .A2(KEYINPUT28), .ZN(n1269) );
XNOR2_X1 U998 ( .A(G107), .B(n1270), .ZN(n1268) );
NOR2_X1 U999 ( .A1(G104), .A2(KEYINPUT23), .ZN(n1270) );
XOR2_X1 U1000 ( .A(n1271), .B(n1272), .Z(n1086) );
NOR2_X1 U1001 ( .A1(KEYINPUT52), .A2(n1273), .ZN(n1272) );
XNOR2_X1 U1002 ( .A(G113), .B(KEYINPUT37), .ZN(n1271) );
XOR2_X1 U1003 ( .A(G125), .B(n1062), .Z(n1141) );
INV_X1 U1004 ( .A(n1190), .ZN(n1001) );
NAND2_X1 U1005 ( .A1(G214), .A2(n1261), .ZN(n1190) );
NAND2_X1 U1006 ( .A1(n1274), .A2(n1209), .ZN(n1261) );
INV_X1 U1007 ( .A(G237), .ZN(n1274) );
NAND2_X1 U1008 ( .A1(G221), .A2(n1208), .ZN(n1193) );
NAND2_X1 U1009 ( .A1(G234), .A2(n1209), .ZN(n1208) );
XOR2_X1 U1010 ( .A(n1275), .B(n1121), .Z(n1019) );
INV_X1 U1011 ( .A(G469), .ZN(n1121) );
NAND2_X1 U1012 ( .A1(n1276), .A2(n1209), .ZN(n1275) );
XOR2_X1 U1013 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U1014 ( .A(n1062), .B(n1279), .Z(n1278) );
XOR2_X1 U1015 ( .A(KEYINPUT44), .B(n1131), .Z(n1279) );
NOR2_X1 U1016 ( .A1(n1041), .A2(G953), .ZN(n1131) );
INV_X1 U1017 ( .A(G227), .ZN(n1041) );
XNOR2_X1 U1018 ( .A(n1133), .B(n1130), .ZN(n1277) );
XOR2_X1 U1019 ( .A(G110), .B(G140), .Z(n1130) );
XOR2_X1 U1020 ( .A(n1113), .B(n1280), .Z(n1133) );
XNOR2_X1 U1021 ( .A(G107), .B(n1108), .ZN(n1280) );
INV_X1 U1022 ( .A(G104), .ZN(n1108) );
XOR2_X1 U1023 ( .A(G101), .B(n1281), .Z(n1113) );
INV_X1 U1024 ( .A(n1036), .ZN(n1024) );
XOR2_X1 U1025 ( .A(n1282), .B(n1116), .Z(n1036) );
INV_X1 U1026 ( .A(G472), .ZN(n1116) );
NAND2_X1 U1027 ( .A1(n1283), .A2(n1209), .ZN(n1282) );
INV_X1 U1028 ( .A(G902), .ZN(n1209) );
XOR2_X1 U1029 ( .A(n1284), .B(n1285), .Z(n1283) );
XOR2_X1 U1030 ( .A(n1117), .B(G101), .Z(n1285) );
NAND2_X1 U1031 ( .A1(n1236), .A2(G210), .ZN(n1117) );
NOR2_X1 U1032 ( .A1(G953), .A2(G237), .ZN(n1236) );
NAND2_X1 U1033 ( .A1(KEYINPUT24), .A2(n1286), .ZN(n1284) );
XOR2_X1 U1034 ( .A(n1287), .B(n1112), .Z(n1286) );
XOR2_X1 U1035 ( .A(n1288), .B(n1289), .Z(n1112) );
XNOR2_X1 U1036 ( .A(KEYINPUT43), .B(n1204), .ZN(n1289) );
INV_X1 U1037 ( .A(G113), .ZN(n1204) );
XOR2_X1 U1038 ( .A(n1273), .B(n1062), .Z(n1288) );
XNOR2_X1 U1039 ( .A(n1290), .B(n1250), .ZN(n1062) );
XNOR2_X1 U1040 ( .A(n1228), .B(G143), .ZN(n1250) );
INV_X1 U1041 ( .A(G128), .ZN(n1228) );
XNOR2_X1 U1042 ( .A(G146), .B(KEYINPUT12), .ZN(n1290) );
XNOR2_X1 U1043 ( .A(G116), .B(G119), .ZN(n1273) );
NAND2_X1 U1044 ( .A1(KEYINPUT19), .A2(n1281), .ZN(n1287) );
XNOR2_X1 U1045 ( .A(n1291), .B(n1065), .ZN(n1281) );
XOR2_X1 U1046 ( .A(G137), .B(G134), .Z(n1065) );
XNOR2_X1 U1047 ( .A(G131), .B(KEYINPUT47), .ZN(n1291) );
endmodule


