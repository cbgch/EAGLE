//Key = 0000100011011001001001111101001001101111100001100100001100110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298;

XOR2_X1 U705 ( .A(n982), .B(n983), .Z(G9) );
NOR2_X1 U706 ( .A1(KEYINPUT19), .A2(n984), .ZN(n983) );
INV_X1 U707 ( .A(G107), .ZN(n984) );
NOR2_X1 U708 ( .A1(n985), .A2(n986), .ZN(G75) );
NOR4_X1 U709 ( .A1(n987), .A2(n988), .A3(G953), .A4(n989), .ZN(n986) );
NOR3_X1 U710 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n988) );
NOR2_X1 U711 ( .A1(n993), .A2(n994), .ZN(n991) );
NOR2_X1 U712 ( .A1(n995), .A2(n996), .ZN(n994) );
NOR3_X1 U713 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n995) );
NOR3_X1 U714 ( .A1(n1000), .A2(KEYINPUT61), .A3(n1001), .ZN(n999) );
NOR2_X1 U715 ( .A1(n1002), .A2(n1003), .ZN(n998) );
INV_X1 U716 ( .A(n1000), .ZN(n1003) );
NOR2_X1 U717 ( .A1(n1004), .A2(n1005), .ZN(n1002) );
NOR2_X1 U718 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
AND2_X1 U719 ( .A1(n1008), .A2(KEYINPUT61), .ZN(n1004) );
NOR2_X1 U720 ( .A1(n1009), .A2(n1010), .ZN(n993) );
NAND2_X1 U721 ( .A1(n1011), .A2(n1012), .ZN(n987) );
NAND2_X1 U722 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND3_X1 U723 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NAND2_X1 U724 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
INV_X1 U725 ( .A(KEYINPUT40), .ZN(n1019) );
NAND4_X1 U726 ( .A1(n1020), .A2(n1021), .A3(n1000), .A4(n1022), .ZN(n1018) );
NAND4_X1 U727 ( .A1(n1020), .A2(n1023), .A3(n1022), .A4(n1024), .ZN(n1016) );
NAND2_X1 U728 ( .A1(n1000), .A2(n1025), .ZN(n1015) );
NAND2_X1 U729 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND4_X1 U730 ( .A1(n1028), .A2(n1029), .A3(n1024), .A4(n1030), .ZN(n1027) );
XNOR2_X1 U731 ( .A(KEYINPUT48), .B(n990), .ZN(n1030) );
NAND2_X1 U732 ( .A1(n1020), .A2(n1031), .ZN(n1026) );
NAND2_X1 U733 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND3_X1 U734 ( .A1(n1021), .A2(n1022), .A3(KEYINPUT40), .ZN(n1033) );
NAND2_X1 U735 ( .A1(n1024), .A2(n1034), .ZN(n1032) );
INV_X1 U736 ( .A(n990), .ZN(n1020) );
NAND2_X1 U737 ( .A1(KEYINPUT18), .A2(n1035), .ZN(n990) );
NOR3_X1 U738 ( .A1(n989), .A2(G953), .A3(G952), .ZN(n985) );
AND3_X1 U739 ( .A1(n1036), .A2(n1000), .A3(n1037), .ZN(n989) );
NOR3_X1 U740 ( .A1(n992), .A2(n1038), .A3(n996), .ZN(n1037) );
XNOR2_X1 U741 ( .A(n1039), .B(n1040), .ZN(n1036) );
NAND2_X1 U742 ( .A1(KEYINPUT36), .A2(n1041), .ZN(n1039) );
XOR2_X1 U743 ( .A(n1042), .B(n1043), .Z(G72) );
NOR2_X1 U744 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
AND2_X1 U745 ( .A1(G227), .A2(G900), .ZN(n1044) );
NOR2_X1 U746 ( .A1(KEYINPUT43), .A2(n1046), .ZN(n1042) );
XOR2_X1 U747 ( .A(n1047), .B(n1048), .Z(n1046) );
NOR2_X1 U748 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
XOR2_X1 U749 ( .A(n1051), .B(n1052), .Z(n1050) );
XNOR2_X1 U750 ( .A(n1053), .B(n1054), .ZN(n1051) );
NOR2_X1 U751 ( .A1(G900), .A2(n1045), .ZN(n1049) );
NAND2_X1 U752 ( .A1(n1045), .A2(n1055), .ZN(n1047) );
NAND2_X1 U753 ( .A1(n1056), .A2(n1057), .ZN(G69) );
NAND2_X1 U754 ( .A1(G953), .A2(n1058), .ZN(n1057) );
XOR2_X1 U755 ( .A(n1059), .B(n1060), .Z(n1056) );
NAND2_X1 U756 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U757 ( .A1(G953), .A2(n1063), .ZN(n1062) );
INV_X1 U758 ( .A(n1064), .ZN(n1061) );
NAND2_X1 U759 ( .A1(n1065), .A2(KEYINPUT30), .ZN(n1059) );
XOR2_X1 U760 ( .A(n1066), .B(n1067), .Z(n1065) );
XOR2_X1 U761 ( .A(G101), .B(n1068), .Z(n1067) );
NOR2_X1 U762 ( .A1(KEYINPUT1), .A2(n1069), .ZN(n1068) );
XOR2_X1 U763 ( .A(n1070), .B(n1071), .Z(n1066) );
NOR2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(G66) );
XOR2_X1 U765 ( .A(n1074), .B(n1075), .Z(n1073) );
NAND2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U767 ( .A1(n1072), .A2(n1078), .ZN(G63) );
XOR2_X1 U768 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND2_X1 U769 ( .A1(n1076), .A2(G478), .ZN(n1080) );
NOR2_X1 U770 ( .A1(n1072), .A2(n1081), .ZN(G60) );
NOR2_X1 U771 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XOR2_X1 U772 ( .A(KEYINPUT35), .B(n1084), .Z(n1083) );
NOR2_X1 U773 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
AND2_X1 U774 ( .A1(n1086), .A2(n1085), .ZN(n1082) );
NAND2_X1 U775 ( .A1(n1076), .A2(n1087), .ZN(n1085) );
XOR2_X1 U776 ( .A(KEYINPUT53), .B(G475), .Z(n1087) );
XOR2_X1 U777 ( .A(G104), .B(n1088), .Z(G6) );
NOR2_X1 U778 ( .A1(n1089), .A2(n1090), .ZN(G57) );
XOR2_X1 U779 ( .A(n1091), .B(n1092), .Z(n1090) );
XNOR2_X1 U780 ( .A(n1093), .B(n1094), .ZN(n1092) );
XOR2_X1 U781 ( .A(n1095), .B(n1096), .Z(n1091) );
XOR2_X1 U782 ( .A(n1097), .B(KEYINPUT49), .Z(n1096) );
NAND2_X1 U783 ( .A1(n1076), .A2(G472), .ZN(n1097) );
NAND2_X1 U784 ( .A1(KEYINPUT63), .A2(n1053), .ZN(n1095) );
NOR2_X1 U785 ( .A1(n1098), .A2(n1099), .ZN(n1089) );
XOR2_X1 U786 ( .A(KEYINPUT47), .B(G952), .Z(n1099) );
XOR2_X1 U787 ( .A(KEYINPUT54), .B(n1100), .Z(n1098) );
NOR2_X1 U788 ( .A1(n1072), .A2(n1101), .ZN(G54) );
XOR2_X1 U789 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U790 ( .A(KEYINPUT32), .B(n1104), .Z(n1103) );
NOR2_X1 U791 ( .A1(KEYINPUT52), .A2(n1105), .ZN(n1104) );
XNOR2_X1 U792 ( .A(KEYINPUT38), .B(n1106), .ZN(n1105) );
XOR2_X1 U793 ( .A(n1107), .B(n1108), .Z(n1102) );
NAND2_X1 U794 ( .A1(n1076), .A2(G469), .ZN(n1107) );
NOR2_X1 U795 ( .A1(n1072), .A2(n1109), .ZN(G51) );
XOR2_X1 U796 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U797 ( .A1(n1076), .A2(n1041), .ZN(n1111) );
NOR2_X1 U798 ( .A1(n1112), .A2(n1011), .ZN(n1076) );
NOR2_X1 U799 ( .A1(n1055), .A2(n1064), .ZN(n1011) );
NAND4_X1 U800 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1064) );
NOR4_X1 U801 ( .A1(n1117), .A2(n1118), .A3(n1088), .A4(n982), .ZN(n1116) );
AND3_X1 U802 ( .A1(n1119), .A2(n1024), .A3(n1120), .ZN(n982) );
AND3_X1 U803 ( .A1(n1120), .A2(n1024), .A3(n1023), .ZN(n1088) );
NOR2_X1 U804 ( .A1(n1121), .A2(n1122), .ZN(n1115) );
NOR2_X1 U805 ( .A1(n1001), .A2(n1123), .ZN(n1122) );
NAND4_X1 U806 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1055) );
AND3_X1 U807 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1127) );
NAND4_X1 U808 ( .A1(n1021), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1126) );
NAND2_X1 U809 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
INV_X1 U810 ( .A(n1034), .ZN(n1135) );
OR2_X1 U811 ( .A1(n1136), .A2(KEYINPUT9), .ZN(n1134) );
NAND4_X1 U812 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1034), .ZN(n1132) );
NAND2_X1 U813 ( .A1(KEYINPUT9), .A2(n997), .ZN(n1139) );
INV_X1 U814 ( .A(n1136), .ZN(n997) );
NAND3_X1 U815 ( .A1(n1008), .A2(n1140), .A3(n1141), .ZN(n1138) );
NAND2_X1 U816 ( .A1(n1142), .A2(n1023), .ZN(n1137) );
XNOR2_X1 U817 ( .A(n1013), .B(KEYINPUT58), .ZN(n1142) );
NAND2_X1 U818 ( .A1(n1143), .A2(n1144), .ZN(n1110) );
OR2_X1 U819 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U820 ( .A(n1147), .B(KEYINPUT3), .Z(n1143) );
NAND2_X1 U821 ( .A1(n1145), .A2(n1146), .ZN(n1147) );
XOR2_X1 U822 ( .A(n1148), .B(n1149), .Z(n1145) );
NOR2_X1 U823 ( .A1(KEYINPUT26), .A2(n1150), .ZN(n1149) );
XNOR2_X1 U824 ( .A(KEYINPUT10), .B(n1151), .ZN(n1150) );
AND2_X1 U825 ( .A1(n1152), .A2(n1100), .ZN(n1072) );
XNOR2_X1 U826 ( .A(n1045), .B(KEYINPUT29), .ZN(n1100) );
XNOR2_X1 U827 ( .A(KEYINPUT47), .B(G952), .ZN(n1152) );
NAND3_X1 U828 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(G48) );
OR2_X1 U829 ( .A1(n1124), .A2(G146), .ZN(n1155) );
NAND2_X1 U830 ( .A1(n1156), .A2(n1157), .ZN(n1154) );
INV_X1 U831 ( .A(KEYINPUT8), .ZN(n1157) );
NAND2_X1 U832 ( .A1(G146), .A2(n1158), .ZN(n1156) );
XNOR2_X1 U833 ( .A(KEYINPUT39), .B(n1124), .ZN(n1158) );
NAND2_X1 U834 ( .A1(KEYINPUT8), .A2(n1159), .ZN(n1153) );
NAND2_X1 U835 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND3_X1 U836 ( .A1(KEYINPUT39), .A2(G146), .A3(n1124), .ZN(n1161) );
OR2_X1 U837 ( .A1(n1124), .A2(KEYINPUT39), .ZN(n1160) );
NAND3_X1 U838 ( .A1(n1162), .A2(n1023), .A3(n1163), .ZN(n1124) );
XNOR2_X1 U839 ( .A(G143), .B(n1164), .ZN(G45) );
NAND3_X1 U840 ( .A1(n1165), .A2(KEYINPUT22), .A3(n1166), .ZN(n1164) );
NOR3_X1 U841 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1166) );
XNOR2_X1 U842 ( .A(n1008), .B(KEYINPUT46), .ZN(n1165) );
XNOR2_X1 U843 ( .A(G140), .B(n1125), .ZN(G42) );
NAND3_X1 U844 ( .A1(n1170), .A2(n1034), .A3(n1013), .ZN(n1125) );
XOR2_X1 U845 ( .A(n1128), .B(n1171), .Z(G39) );
XOR2_X1 U846 ( .A(KEYINPUT62), .B(G137), .Z(n1171) );
NAND3_X1 U847 ( .A1(n1162), .A2(n1172), .A3(n1173), .ZN(n1128) );
INV_X1 U848 ( .A(n1010), .ZN(n1173) );
NAND3_X1 U849 ( .A1(n1174), .A2(n1000), .A3(n1013), .ZN(n1010) );
XNOR2_X1 U850 ( .A(n1175), .B(n1176), .ZN(G36) );
NOR2_X1 U851 ( .A1(n1136), .A2(n1167), .ZN(n1176) );
NAND2_X1 U852 ( .A1(n1013), .A2(n1119), .ZN(n1136) );
XNOR2_X1 U853 ( .A(G131), .B(n1177), .ZN(G33) );
NAND3_X1 U854 ( .A1(n1013), .A2(n1023), .A3(n1178), .ZN(n1177) );
INV_X1 U855 ( .A(n1167), .ZN(n1178) );
NAND2_X1 U856 ( .A1(n1021), .A2(n1162), .ZN(n1167) );
NOR2_X1 U857 ( .A1(n1006), .A2(n1038), .ZN(n1013) );
INV_X1 U858 ( .A(n1007), .ZN(n1038) );
XNOR2_X1 U859 ( .A(G128), .B(n1130), .ZN(G30) );
NAND3_X1 U860 ( .A1(n1162), .A2(n1119), .A3(n1163), .ZN(n1130) );
AND2_X1 U861 ( .A1(n1034), .A2(n1131), .ZN(n1162) );
XNOR2_X1 U862 ( .A(n1118), .B(n1179), .ZN(G3) );
NAND2_X1 U863 ( .A1(KEYINPUT33), .A2(G101), .ZN(n1179) );
AND3_X1 U864 ( .A1(n1000), .A2(n1120), .A3(n1021), .ZN(n1118) );
XNOR2_X1 U865 ( .A(G125), .B(n1180), .ZN(G27) );
NAND2_X1 U866 ( .A1(KEYINPUT23), .A2(n1181), .ZN(n1180) );
INV_X1 U867 ( .A(n1129), .ZN(n1181) );
NAND3_X1 U868 ( .A1(n1022), .A2(n1008), .A3(n1170), .ZN(n1129) );
AND4_X1 U869 ( .A1(n1174), .A2(n1023), .A3(n1182), .A4(n1131), .ZN(n1170) );
NAND2_X1 U870 ( .A1(n1183), .A2(n1184), .ZN(n1131) );
NAND2_X1 U871 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
INV_X1 U872 ( .A(G900), .ZN(n1186) );
XNOR2_X1 U873 ( .A(n1121), .B(n1187), .ZN(G24) );
XNOR2_X1 U874 ( .A(G122), .B(KEYINPUT31), .ZN(n1187) );
AND4_X1 U875 ( .A1(n1008), .A2(n1140), .A3(n1024), .A4(n1188), .ZN(n1121) );
NOR2_X1 U876 ( .A1(n1189), .A2(n1169), .ZN(n1188) );
INV_X1 U877 ( .A(n996), .ZN(n1024) );
NAND2_X1 U878 ( .A1(n1182), .A2(n1190), .ZN(n996) );
NAND3_X1 U879 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(G21) );
NAND2_X1 U880 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NAND2_X1 U881 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
XNOR2_X1 U882 ( .A(KEYINPUT44), .B(n1198), .ZN(n1196) );
INV_X1 U883 ( .A(n1113), .ZN(n1194) );
NAND3_X1 U884 ( .A1(G119), .A2(n1113), .A3(n1197), .ZN(n1192) );
INV_X1 U885 ( .A(KEYINPUT42), .ZN(n1197) );
NAND3_X1 U886 ( .A1(n1163), .A2(n1000), .A3(n1199), .ZN(n1113) );
AND3_X1 U887 ( .A1(n1008), .A2(n1172), .A3(n1174), .ZN(n1163) );
NAND2_X1 U888 ( .A1(KEYINPUT42), .A2(n1198), .ZN(n1191) );
NAND2_X1 U889 ( .A1(n1200), .A2(n1201), .ZN(G18) );
NAND2_X1 U890 ( .A1(n1117), .A2(n1202), .ZN(n1201) );
XOR2_X1 U891 ( .A(KEYINPUT4), .B(n1203), .Z(n1200) );
NOR2_X1 U892 ( .A1(n1117), .A2(n1202), .ZN(n1203) );
INV_X1 U893 ( .A(G116), .ZN(n1202) );
AND4_X1 U894 ( .A1(n1199), .A2(n1021), .A3(n1119), .A4(n1008), .ZN(n1117) );
NOR2_X1 U895 ( .A1(n1141), .A2(n1168), .ZN(n1119) );
INV_X1 U896 ( .A(n1140), .ZN(n1168) );
XOR2_X1 U897 ( .A(G113), .B(n1204), .Z(G15) );
NOR3_X1 U898 ( .A1(n1205), .A2(KEYINPUT16), .A3(n1001), .ZN(n1204) );
XNOR2_X1 U899 ( .A(KEYINPUT27), .B(n1123), .ZN(n1205) );
NAND3_X1 U900 ( .A1(n1021), .A2(n1023), .A3(n1199), .ZN(n1123) );
INV_X1 U901 ( .A(n1189), .ZN(n1199) );
NAND2_X1 U902 ( .A1(n1022), .A2(n1206), .ZN(n1189) );
INV_X1 U903 ( .A(n992), .ZN(n1022) );
NAND2_X1 U904 ( .A1(n1028), .A2(n1207), .ZN(n992) );
NOR2_X1 U905 ( .A1(n1169), .A2(n1140), .ZN(n1023) );
AND2_X1 U906 ( .A1(n1190), .A2(n1172), .ZN(n1021) );
XNOR2_X1 U907 ( .A(n1182), .B(KEYINPUT5), .ZN(n1172) );
XNOR2_X1 U908 ( .A(n1208), .B(n1209), .ZN(G12) );
NOR2_X1 U909 ( .A1(KEYINPUT60), .A2(n1114), .ZN(n1209) );
NAND4_X1 U910 ( .A1(n1174), .A2(n1000), .A3(n1182), .A4(n1120), .ZN(n1114) );
AND3_X1 U911 ( .A1(n1008), .A2(n1206), .A3(n1034), .ZN(n1120) );
NOR2_X1 U912 ( .A1(n1028), .A2(n1029), .ZN(n1034) );
INV_X1 U913 ( .A(n1207), .ZN(n1029) );
NAND2_X1 U914 ( .A1(G221), .A2(n1210), .ZN(n1207) );
XOR2_X1 U915 ( .A(n1211), .B(G469), .Z(n1028) );
NAND2_X1 U916 ( .A1(n1212), .A2(n1112), .ZN(n1211) );
XNOR2_X1 U917 ( .A(n1108), .B(n1213), .ZN(n1212) );
NOR2_X1 U918 ( .A1(KEYINPUT50), .A2(n1214), .ZN(n1213) );
XNOR2_X1 U919 ( .A(n1053), .B(KEYINPUT38), .ZN(n1214) );
XNOR2_X1 U920 ( .A(n1215), .B(n1216), .ZN(n1108) );
XOR2_X1 U921 ( .A(G104), .B(n1217), .Z(n1216) );
XNOR2_X1 U922 ( .A(n1208), .B(G107), .ZN(n1217) );
XNOR2_X1 U923 ( .A(n1052), .B(n1218), .ZN(n1215) );
XOR2_X1 U924 ( .A(n1219), .B(n1220), .Z(n1218) );
NOR2_X1 U925 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
XNOR2_X1 U926 ( .A(G227), .B(KEYINPUT28), .ZN(n1221) );
NOR2_X1 U927 ( .A1(G101), .A2(n1223), .ZN(n1219) );
XNOR2_X1 U928 ( .A(KEYINPUT57), .B(KEYINPUT55), .ZN(n1223) );
XNOR2_X1 U929 ( .A(n1224), .B(n1225), .ZN(n1052) );
NAND2_X1 U930 ( .A1(KEYINPUT21), .A2(n1226), .ZN(n1224) );
NAND2_X1 U931 ( .A1(n1183), .A2(n1227), .ZN(n1206) );
NAND2_X1 U932 ( .A1(n1185), .A2(n1058), .ZN(n1227) );
INV_X1 U933 ( .A(G898), .ZN(n1058) );
AND3_X1 U934 ( .A1(G953), .A2(n1035), .A3(G902), .ZN(n1185) );
NAND3_X1 U935 ( .A1(n1035), .A2(n1045), .A3(G952), .ZN(n1183) );
INV_X1 U936 ( .A(G953), .ZN(n1045) );
NAND2_X1 U937 ( .A1(G237), .A2(G234), .ZN(n1035) );
INV_X1 U938 ( .A(n1001), .ZN(n1008) );
NAND2_X1 U939 ( .A1(n1006), .A2(n1007), .ZN(n1001) );
NAND2_X1 U940 ( .A1(G214), .A2(n1228), .ZN(n1007) );
XNOR2_X1 U941 ( .A(n1040), .B(n1041), .ZN(n1006) );
AND2_X1 U942 ( .A1(G210), .A2(n1228), .ZN(n1041) );
OR2_X1 U943 ( .A1(G902), .A2(G237), .ZN(n1228) );
NAND2_X1 U944 ( .A1(n1229), .A2(n1112), .ZN(n1040) );
XNOR2_X1 U945 ( .A(n1230), .B(n1231), .ZN(n1229) );
INV_X1 U946 ( .A(n1148), .ZN(n1231) );
XOR2_X1 U947 ( .A(n1054), .B(n1232), .Z(n1148) );
NOR2_X1 U948 ( .A1(n1222), .A2(n1063), .ZN(n1232) );
INV_X1 U949 ( .A(G224), .ZN(n1063) );
XNOR2_X1 U950 ( .A(n1146), .B(n1151), .ZN(n1230) );
NAND2_X1 U951 ( .A1(n1233), .A2(n1234), .ZN(n1146) );
NAND2_X1 U952 ( .A1(n1235), .A2(n1071), .ZN(n1234) );
XOR2_X1 U953 ( .A(n1236), .B(KEYINPUT20), .Z(n1233) );
OR2_X1 U954 ( .A1(n1071), .A2(n1235), .ZN(n1236) );
XNOR2_X1 U955 ( .A(n1237), .B(n1070), .ZN(n1235) );
XNOR2_X1 U956 ( .A(G107), .B(n1238), .ZN(n1070) );
NOR2_X1 U957 ( .A1(G104), .A2(KEYINPUT56), .ZN(n1238) );
XOR2_X1 U958 ( .A(n1239), .B(KEYINPUT41), .Z(n1237) );
XOR2_X1 U959 ( .A(G122), .B(n1240), .Z(n1071) );
NOR2_X1 U960 ( .A1(G110), .A2(KEYINPUT2), .ZN(n1240) );
INV_X1 U961 ( .A(n1009), .ZN(n1182) );
XNOR2_X1 U962 ( .A(n1241), .B(G472), .ZN(n1009) );
NAND2_X1 U963 ( .A1(n1242), .A2(n1112), .ZN(n1241) );
XOR2_X1 U964 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U965 ( .A(n1245), .B(n1093), .Z(n1244) );
XOR2_X1 U966 ( .A(n1239), .B(n1246), .Z(n1093) );
AND2_X1 U967 ( .A1(G210), .A2(n1247), .ZN(n1246) );
XOR2_X1 U968 ( .A(n1069), .B(G101), .Z(n1239) );
XNOR2_X1 U969 ( .A(G113), .B(n1248), .ZN(n1069) );
XNOR2_X1 U970 ( .A(n1198), .B(G116), .ZN(n1248) );
NAND3_X1 U971 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1245) );
NAND2_X1 U972 ( .A1(n1094), .A2(n1053), .ZN(n1251) );
NAND2_X1 U973 ( .A1(KEYINPUT13), .A2(n1252), .ZN(n1250) );
NAND2_X1 U974 ( .A1(n1106), .A2(n1253), .ZN(n1252) );
XNOR2_X1 U975 ( .A(KEYINPUT34), .B(n1151), .ZN(n1253) );
NAND2_X1 U976 ( .A1(n1254), .A2(n1255), .ZN(n1249) );
INV_X1 U977 ( .A(KEYINPUT13), .ZN(n1255) );
NAND2_X1 U978 ( .A1(n1256), .A2(n1257), .ZN(n1254) );
NAND3_X1 U979 ( .A1(KEYINPUT34), .A2(n1106), .A3(n1151), .ZN(n1257) );
INV_X1 U980 ( .A(n1053), .ZN(n1106) );
XOR2_X1 U981 ( .A(G131), .B(n1258), .Z(n1053) );
XNOR2_X1 U982 ( .A(G137), .B(n1175), .ZN(n1258) );
OR2_X1 U983 ( .A1(n1151), .A2(KEYINPUT34), .ZN(n1256) );
INV_X1 U984 ( .A(n1094), .ZN(n1151) );
XOR2_X1 U985 ( .A(G143), .B(n1259), .Z(n1094) );
XOR2_X1 U986 ( .A(KEYINPUT37), .B(KEYINPUT24), .Z(n1243) );
NOR2_X1 U987 ( .A1(n1140), .A2(n1141), .ZN(n1000) );
INV_X1 U988 ( .A(n1169), .ZN(n1141) );
XNOR2_X1 U989 ( .A(n1260), .B(n1261), .ZN(n1169) );
XOR2_X1 U990 ( .A(KEYINPUT11), .B(G475), .Z(n1261) );
NAND2_X1 U991 ( .A1(n1112), .A2(n1086), .ZN(n1260) );
NAND2_X1 U992 ( .A1(n1262), .A2(n1263), .ZN(n1086) );
NAND2_X1 U993 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
XOR2_X1 U994 ( .A(n1266), .B(KEYINPUT7), .Z(n1262) );
OR2_X1 U995 ( .A1(n1265), .A2(n1264), .ZN(n1266) );
XNOR2_X1 U996 ( .A(n1267), .B(n1268), .ZN(n1264) );
XOR2_X1 U997 ( .A(G122), .B(G113), .Z(n1268) );
NAND2_X1 U998 ( .A1(KEYINPUT12), .A2(n1269), .ZN(n1267) );
XOR2_X1 U999 ( .A(KEYINPUT59), .B(G104), .Z(n1269) );
XNOR2_X1 U1000 ( .A(n1270), .B(n1271), .ZN(n1265) );
XOR2_X1 U1001 ( .A(G140), .B(n1272), .Z(n1271) );
XNOR2_X1 U1002 ( .A(G146), .B(n1226), .ZN(n1272) );
XNOR2_X1 U1003 ( .A(n1273), .B(n1274), .ZN(n1270) );
XOR2_X1 U1004 ( .A(n1275), .B(G131), .Z(n1273) );
NAND2_X1 U1005 ( .A1(n1247), .A2(G214), .ZN(n1275) );
NOR2_X1 U1006 ( .A1(n1222), .A2(G237), .ZN(n1247) );
XNOR2_X1 U1007 ( .A(n1276), .B(G478), .ZN(n1140) );
NAND2_X1 U1008 ( .A1(n1112), .A2(n1079), .ZN(n1276) );
NAND2_X1 U1009 ( .A1(n1277), .A2(n1278), .ZN(n1079) );
NAND2_X1 U1010 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND2_X1 U1011 ( .A1(G217), .A2(n1281), .ZN(n1280) );
XOR2_X1 U1012 ( .A(n1282), .B(n1283), .Z(n1279) );
XOR2_X1 U1013 ( .A(n1284), .B(KEYINPUT14), .Z(n1277) );
NAND3_X1 U1014 ( .A1(G217), .A2(n1281), .A3(n1285), .ZN(n1284) );
XNOR2_X1 U1015 ( .A(n1282), .B(n1283), .ZN(n1285) );
XNOR2_X1 U1016 ( .A(n1286), .B(n1287), .ZN(n1283) );
NOR2_X1 U1017 ( .A1(KEYINPUT6), .A2(n1175), .ZN(n1287) );
INV_X1 U1018 ( .A(G134), .ZN(n1175) );
XNOR2_X1 U1019 ( .A(G107), .B(G116), .ZN(n1286) );
XOR2_X1 U1020 ( .A(G122), .B(n1288), .Z(n1282) );
XNOR2_X1 U1021 ( .A(n1226), .B(G128), .ZN(n1288) );
INV_X1 U1022 ( .A(G143), .ZN(n1226) );
XOR2_X1 U1023 ( .A(n1190), .B(KEYINPUT45), .Z(n1174) );
XOR2_X1 U1024 ( .A(n1289), .B(n1077), .Z(n1190) );
AND2_X1 U1025 ( .A1(G217), .A2(n1210), .ZN(n1077) );
NAND2_X1 U1026 ( .A1(n1290), .A2(n1112), .ZN(n1210) );
XNOR2_X1 U1027 ( .A(G234), .B(KEYINPUT15), .ZN(n1290) );
NAND2_X1 U1028 ( .A1(n1075), .A2(n1112), .ZN(n1289) );
INV_X1 U1029 ( .A(G902), .ZN(n1112) );
XOR2_X1 U1030 ( .A(n1291), .B(n1292), .Z(n1075) );
XOR2_X1 U1031 ( .A(n1225), .B(n1293), .Z(n1292) );
XNOR2_X1 U1032 ( .A(n1294), .B(n1274), .ZN(n1293) );
INV_X1 U1033 ( .A(n1054), .ZN(n1274) );
XOR2_X1 U1034 ( .A(G125), .B(KEYINPUT0), .Z(n1054) );
NOR2_X1 U1035 ( .A1(KEYINPUT17), .A2(n1208), .ZN(n1294) );
XOR2_X1 U1036 ( .A(G140), .B(n1259), .Z(n1225) );
XOR2_X1 U1037 ( .A(G128), .B(G146), .Z(n1259) );
XOR2_X1 U1038 ( .A(n1295), .B(n1296), .Z(n1291) );
XOR2_X1 U1039 ( .A(KEYINPUT25), .B(G137), .Z(n1296) );
XNOR2_X1 U1040 ( .A(n1297), .B(n1198), .ZN(n1295) );
INV_X1 U1041 ( .A(G119), .ZN(n1198) );
NAND2_X1 U1042 ( .A1(n1281), .A2(G221), .ZN(n1297) );
NOR2_X1 U1043 ( .A1(n1222), .A2(n1298), .ZN(n1281) );
INV_X1 U1044 ( .A(G234), .ZN(n1298) );
XOR2_X1 U1045 ( .A(G953), .B(KEYINPUT51), .Z(n1222) );
INV_X1 U1046 ( .A(G110), .ZN(n1208) );
endmodule


