//Key = 0101110001011101110101100011001000001101110011111110100000101101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373;

XNOR2_X1 U764 ( .A(G107), .B(n1041), .ZN(G9) );
NOR2_X1 U765 ( .A1(n1042), .A2(n1043), .ZN(G75) );
NOR4_X1 U766 ( .A1(G953), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1043) );
NOR2_X1 U767 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U768 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U769 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
INV_X1 U770 ( .A(n1053), .ZN(n1052) );
NOR2_X1 U771 ( .A1(n1054), .A2(n1055), .ZN(n1051) );
NOR2_X1 U772 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U773 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U774 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U775 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U776 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U777 ( .A1(n1066), .A2(n1067), .ZN(n1058) );
NOR2_X1 U778 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR3_X1 U779 ( .A1(n1067), .A2(n1070), .A3(n1061), .ZN(n1054) );
NOR2_X1 U780 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U781 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR4_X1 U782 ( .A1(n1075), .A2(n1061), .A3(n1057), .A4(n1067), .ZN(n1049) );
INV_X1 U783 ( .A(n1076), .ZN(n1067) );
INV_X1 U784 ( .A(n1077), .ZN(n1061) );
NOR2_X1 U785 ( .A1(n1078), .A2(n1079), .ZN(n1075) );
NOR3_X1 U786 ( .A1(n1044), .A2(G953), .A3(G952), .ZN(n1042) );
AND4_X1 U787 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1044) );
NOR4_X1 U788 ( .A1(n1084), .A2(n1085), .A3(n1057), .A4(n1086), .ZN(n1083) );
XNOR2_X1 U789 ( .A(n1087), .B(KEYINPUT63), .ZN(n1085) );
XNOR2_X1 U790 ( .A(n1088), .B(G478), .ZN(n1082) );
XOR2_X1 U791 ( .A(n1089), .B(n1090), .Z(G72) );
NOR2_X1 U792 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U793 ( .A(n1093), .B(n1094), .Z(n1092) );
XNOR2_X1 U794 ( .A(n1095), .B(n1096), .ZN(n1094) );
XNOR2_X1 U795 ( .A(G134), .B(G137), .ZN(n1093) );
NAND2_X1 U796 ( .A1(n1097), .A2(n1098), .ZN(n1089) );
NAND2_X1 U797 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND3_X1 U798 ( .A1(KEYINPUT30), .A2(n1101), .A3(G953), .ZN(n1097) );
NAND2_X1 U799 ( .A1(G900), .A2(G227), .ZN(n1101) );
NAND2_X1 U800 ( .A1(n1102), .A2(n1103), .ZN(G69) );
NAND2_X1 U801 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U802 ( .A1(G953), .A2(n1106), .ZN(n1105) );
NAND3_X1 U803 ( .A1(G953), .A2(n1107), .A3(n1108), .ZN(n1102) );
INV_X1 U804 ( .A(n1104), .ZN(n1108) );
NAND2_X1 U805 ( .A1(n1109), .A2(n1110), .ZN(n1104) );
NAND3_X1 U806 ( .A1(n1111), .A2(KEYINPUT36), .A3(n1112), .ZN(n1110) );
NAND2_X1 U807 ( .A1(n1113), .A2(n1114), .ZN(n1109) );
NAND2_X1 U808 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U809 ( .A1(KEYINPUT50), .A2(n1117), .ZN(n1116) );
INV_X1 U810 ( .A(n1111), .ZN(n1117) );
NAND2_X1 U811 ( .A1(n1111), .A2(n1118), .ZN(n1115) );
NAND2_X1 U812 ( .A1(KEYINPUT50), .A2(KEYINPUT36), .ZN(n1118) );
NOR2_X1 U813 ( .A1(n1119), .A2(n1120), .ZN(n1111) );
XOR2_X1 U814 ( .A(n1121), .B(n1122), .Z(n1119) );
XOR2_X1 U815 ( .A(KEYINPUT31), .B(KEYINPUT1), .Z(n1122) );
INV_X1 U816 ( .A(n1112), .ZN(n1113) );
NAND2_X1 U817 ( .A1(n1100), .A2(n1123), .ZN(n1112) );
NAND2_X1 U818 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U819 ( .A(n1126), .B(KEYINPUT33), .Z(n1124) );
NAND2_X1 U820 ( .A1(G898), .A2(G224), .ZN(n1107) );
NOR2_X1 U821 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XOR2_X1 U822 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U823 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
XNOR2_X1 U824 ( .A(n1133), .B(KEYINPUT27), .ZN(n1127) );
NOR2_X1 U825 ( .A1(n1133), .A2(n1134), .ZN(G63) );
NOR3_X1 U826 ( .A1(n1088), .A2(n1135), .A3(n1136), .ZN(n1134) );
AND3_X1 U827 ( .A1(n1137), .A2(G478), .A3(n1131), .ZN(n1136) );
NOR2_X1 U828 ( .A1(n1138), .A2(n1137), .ZN(n1135) );
NOR2_X1 U829 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR2_X1 U830 ( .A1(n1133), .A2(n1141), .ZN(G60) );
XOR2_X1 U831 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND2_X1 U832 ( .A1(n1131), .A2(G475), .ZN(n1142) );
XNOR2_X1 U833 ( .A(G104), .B(n1144), .ZN(G6) );
NOR2_X1 U834 ( .A1(n1133), .A2(n1145), .ZN(G57) );
XOR2_X1 U835 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U836 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U837 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
OR2_X1 U838 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U839 ( .A(n1154), .B(KEYINPUT62), .Z(n1150) );
NAND2_X1 U840 ( .A1(n1153), .A2(n1152), .ZN(n1154) );
XOR2_X1 U841 ( .A(n1155), .B(n1156), .Z(n1146) );
NOR2_X1 U842 ( .A1(KEYINPUT6), .A2(n1157), .ZN(n1156) );
XNOR2_X1 U843 ( .A(n1158), .B(n1159), .ZN(n1157) );
NOR2_X1 U844 ( .A1(KEYINPUT56), .A2(n1160), .ZN(n1159) );
INV_X1 U845 ( .A(n1161), .ZN(n1160) );
NAND2_X1 U846 ( .A1(n1131), .A2(G472), .ZN(n1155) );
NOR2_X1 U847 ( .A1(n1133), .A2(n1162), .ZN(G54) );
NOR2_X1 U848 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U849 ( .A(KEYINPUT8), .B(n1165), .Z(n1164) );
NOR2_X1 U850 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
AND2_X1 U851 ( .A1(n1167), .A2(n1166), .ZN(n1163) );
XNOR2_X1 U852 ( .A(n1168), .B(n1169), .ZN(n1166) );
XNOR2_X1 U853 ( .A(n1170), .B(n1171), .ZN(n1169) );
XNOR2_X1 U854 ( .A(KEYINPUT47), .B(n1172), .ZN(n1168) );
NOR2_X1 U855 ( .A1(KEYINPUT2), .A2(n1173), .ZN(n1172) );
NAND2_X1 U856 ( .A1(n1131), .A2(G469), .ZN(n1167) );
NOR2_X1 U857 ( .A1(n1133), .A2(n1174), .ZN(G51) );
XOR2_X1 U858 ( .A(n1121), .B(n1175), .Z(n1174) );
XOR2_X1 U859 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U860 ( .A1(KEYINPUT10), .A2(n1178), .ZN(n1177) );
XNOR2_X1 U861 ( .A(n1161), .B(n1179), .ZN(n1178) );
XOR2_X1 U862 ( .A(G125), .B(n1180), .Z(n1179) );
NAND2_X1 U863 ( .A1(n1131), .A2(n1181), .ZN(n1176) );
NOR2_X1 U864 ( .A1(n1182), .A2(n1139), .ZN(n1131) );
INV_X1 U865 ( .A(n1046), .ZN(n1139) );
NAND3_X1 U866 ( .A1(n1183), .A2(n1126), .A3(n1125), .ZN(n1046) );
AND4_X1 U867 ( .A1(n1184), .A2(n1185), .A3(n1144), .A4(n1186), .ZN(n1125) );
AND4_X1 U868 ( .A1(n1041), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1186) );
NAND3_X1 U869 ( .A1(n1190), .A2(n1077), .A3(n1078), .ZN(n1041) );
NAND3_X1 U870 ( .A1(n1190), .A2(n1077), .A3(n1079), .ZN(n1144) );
NAND2_X1 U871 ( .A1(n1063), .A2(n1191), .ZN(n1126) );
XNOR2_X1 U872 ( .A(KEYINPUT29), .B(n1192), .ZN(n1191) );
INV_X1 U873 ( .A(n1099), .ZN(n1183) );
NAND2_X1 U874 ( .A1(n1193), .A2(n1194), .ZN(n1099) );
NOR4_X1 U875 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1194) );
NOR4_X1 U876 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1193) );
NOR2_X1 U877 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
INV_X1 U878 ( .A(n1205), .ZN(n1199) );
NOR2_X1 U879 ( .A1(n1100), .A2(G952), .ZN(n1133) );
XNOR2_X1 U880 ( .A(G146), .B(n1206), .ZN(G48) );
NAND2_X1 U881 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U882 ( .A1(KEYINPUT22), .A2(n1209), .ZN(n1208) );
NAND2_X1 U883 ( .A1(KEYINPUT24), .A2(n1201), .ZN(n1207) );
INV_X1 U884 ( .A(n1209), .ZN(n1201) );
NAND3_X1 U885 ( .A1(n1079), .A2(n1063), .A3(n1210), .ZN(n1209) );
XOR2_X1 U886 ( .A(G143), .B(n1200), .Z(G45) );
AND4_X1 U887 ( .A1(n1211), .A2(n1069), .A3(n1212), .A4(n1063), .ZN(n1200) );
NOR2_X1 U888 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND2_X1 U889 ( .A1(n1215), .A2(n1216), .ZN(G42) );
NAND2_X1 U890 ( .A1(G140), .A2(n1205), .ZN(n1216) );
XOR2_X1 U891 ( .A(n1217), .B(KEYINPUT59), .Z(n1215) );
OR2_X1 U892 ( .A1(n1205), .A2(G140), .ZN(n1217) );
NAND4_X1 U893 ( .A1(n1076), .A2(n1211), .A3(n1079), .A4(n1068), .ZN(n1205) );
XOR2_X1 U894 ( .A(G137), .B(n1198), .Z(G39) );
AND3_X1 U895 ( .A1(n1210), .A2(n1053), .A3(n1076), .ZN(n1198) );
XOR2_X1 U896 ( .A(n1218), .B(n1197), .Z(G36) );
AND2_X1 U897 ( .A1(n1219), .A2(n1078), .ZN(n1197) );
XNOR2_X1 U898 ( .A(G134), .B(KEYINPUT58), .ZN(n1218) );
XNOR2_X1 U899 ( .A(G131), .B(n1220), .ZN(G33) );
NAND2_X1 U900 ( .A1(KEYINPUT5), .A2(n1196), .ZN(n1220) );
AND2_X1 U901 ( .A1(n1219), .A2(n1079), .ZN(n1196) );
AND3_X1 U902 ( .A1(n1211), .A2(n1069), .A3(n1076), .ZN(n1219) );
NOR2_X1 U903 ( .A1(n1064), .A2(n1084), .ZN(n1076) );
INV_X1 U904 ( .A(n1065), .ZN(n1084) );
XNOR2_X1 U905 ( .A(n1195), .B(n1221), .ZN(G30) );
NAND2_X1 U906 ( .A1(n1222), .A2(G128), .ZN(n1221) );
XNOR2_X1 U907 ( .A(KEYINPUT40), .B(KEYINPUT16), .ZN(n1222) );
AND3_X1 U908 ( .A1(n1078), .A2(n1063), .A3(n1210), .ZN(n1195) );
AND3_X1 U909 ( .A1(n1223), .A2(n1224), .A3(n1211), .ZN(n1210) );
AND2_X1 U910 ( .A1(n1072), .A2(n1225), .ZN(n1211) );
XNOR2_X1 U911 ( .A(n1153), .B(n1226), .ZN(G3) );
NOR2_X1 U912 ( .A1(n1227), .A2(n1192), .ZN(n1226) );
NAND4_X1 U913 ( .A1(n1053), .A2(n1069), .A3(n1072), .A4(n1228), .ZN(n1192) );
XOR2_X1 U914 ( .A(G125), .B(n1229), .Z(G27) );
NOR2_X1 U915 ( .A1(n1230), .A2(n1204), .ZN(n1229) );
NAND4_X1 U916 ( .A1(n1079), .A2(n1068), .A3(n1063), .A4(n1231), .ZN(n1204) );
XNOR2_X1 U917 ( .A(n1203), .B(KEYINPUT37), .ZN(n1230) );
INV_X1 U918 ( .A(n1225), .ZN(n1203) );
NAND2_X1 U919 ( .A1(n1048), .A2(n1232), .ZN(n1225) );
NAND3_X1 U920 ( .A1(G902), .A2(n1233), .A3(n1091), .ZN(n1232) );
NOR2_X1 U921 ( .A1(n1100), .A2(G900), .ZN(n1091) );
XNOR2_X1 U922 ( .A(G122), .B(n1184), .ZN(G24) );
NAND4_X1 U923 ( .A1(n1234), .A2(n1235), .A3(n1077), .A4(n1087), .ZN(n1184) );
NAND2_X1 U924 ( .A1(n1236), .A2(n1237), .ZN(n1077) );
NAND2_X1 U925 ( .A1(n1069), .A2(n1238), .ZN(n1237) );
INV_X1 U926 ( .A(KEYINPUT41), .ZN(n1238) );
NAND3_X1 U927 ( .A1(n1080), .A2(n1239), .A3(KEYINPUT41), .ZN(n1236) );
NAND2_X1 U928 ( .A1(n1240), .A2(n1241), .ZN(G21) );
NAND2_X1 U929 ( .A1(n1242), .A2(n1185), .ZN(n1241) );
NAND2_X1 U930 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
NAND2_X1 U931 ( .A1(KEYINPUT54), .A2(n1245), .ZN(n1244) );
NAND3_X1 U932 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1240) );
INV_X1 U933 ( .A(KEYINPUT54), .ZN(n1248) );
NAND2_X1 U934 ( .A1(G119), .A2(n1245), .ZN(n1247) );
INV_X1 U935 ( .A(KEYINPUT53), .ZN(n1245) );
NAND2_X1 U936 ( .A1(n1249), .A2(n1243), .ZN(n1246) );
OR2_X1 U937 ( .A1(n1185), .A2(KEYINPUT53), .ZN(n1249) );
NAND4_X1 U938 ( .A1(n1235), .A2(n1053), .A3(n1223), .A4(n1224), .ZN(n1185) );
NAND3_X1 U939 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(G18) );
NAND2_X1 U940 ( .A1(KEYINPUT43), .A2(n1189), .ZN(n1252) );
OR3_X1 U941 ( .A1(n1189), .A2(KEYINPUT43), .A3(G116), .ZN(n1251) );
NAND2_X1 U942 ( .A1(G116), .A2(n1253), .ZN(n1250) );
NAND2_X1 U943 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
INV_X1 U944 ( .A(KEYINPUT43), .ZN(n1255) );
XOR2_X1 U945 ( .A(n1189), .B(KEYINPUT9), .Z(n1254) );
NAND3_X1 U946 ( .A1(n1078), .A2(n1069), .A3(n1235), .ZN(n1189) );
NOR2_X1 U947 ( .A1(n1087), .A2(n1214), .ZN(n1078) );
NAND2_X1 U948 ( .A1(n1256), .A2(n1257), .ZN(G15) );
NAND3_X1 U949 ( .A1(KEYINPUT44), .A2(n1188), .A3(n1258), .ZN(n1257) );
INV_X1 U950 ( .A(n1259), .ZN(n1258) );
NAND2_X1 U951 ( .A1(n1259), .A2(n1260), .ZN(n1256) );
NAND2_X1 U952 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
OR2_X1 U953 ( .A1(n1188), .A2(KEYINPUT7), .ZN(n1262) );
NAND2_X1 U954 ( .A1(n1263), .A2(n1188), .ZN(n1261) );
NAND3_X1 U955 ( .A1(n1079), .A2(n1069), .A3(n1235), .ZN(n1188) );
AND3_X1 U956 ( .A1(n1231), .A2(n1228), .A3(n1063), .ZN(n1235) );
NOR2_X1 U957 ( .A1(n1223), .A2(n1080), .ZN(n1069) );
INV_X1 U958 ( .A(n1224), .ZN(n1080) );
NOR2_X1 U959 ( .A1(n1234), .A2(n1213), .ZN(n1079) );
INV_X1 U960 ( .A(n1087), .ZN(n1213) );
NAND2_X1 U961 ( .A1(KEYINPUT44), .A2(n1264), .ZN(n1263) );
INV_X1 U962 ( .A(KEYINPUT7), .ZN(n1264) );
XOR2_X1 U963 ( .A(G113), .B(KEYINPUT12), .Z(n1259) );
XNOR2_X1 U964 ( .A(G110), .B(n1187), .ZN(G12) );
NAND3_X1 U965 ( .A1(n1068), .A2(n1190), .A3(n1053), .ZN(n1187) );
NOR2_X1 U966 ( .A1(n1087), .A2(n1234), .ZN(n1053) );
INV_X1 U967 ( .A(n1214), .ZN(n1234) );
NAND2_X1 U968 ( .A1(n1265), .A2(n1266), .ZN(n1214) );
NAND2_X1 U969 ( .A1(n1267), .A2(n1140), .ZN(n1266) );
INV_X1 U970 ( .A(G478), .ZN(n1140) );
XOR2_X1 U971 ( .A(KEYINPUT11), .B(n1088), .Z(n1267) );
NAND2_X1 U972 ( .A1(n1268), .A2(G478), .ZN(n1265) );
XOR2_X1 U973 ( .A(KEYINPUT32), .B(n1088), .Z(n1268) );
NOR2_X1 U974 ( .A1(n1137), .A2(G902), .ZN(n1088) );
XNOR2_X1 U975 ( .A(n1269), .B(n1270), .ZN(n1137) );
XOR2_X1 U976 ( .A(n1271), .B(n1272), .Z(n1270) );
NAND2_X1 U977 ( .A1(G217), .A2(n1273), .ZN(n1272) );
NAND2_X1 U978 ( .A1(KEYINPUT46), .A2(n1274), .ZN(n1271) );
NAND2_X1 U979 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NAND2_X1 U980 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
XNOR2_X1 U981 ( .A(G134), .B(KEYINPUT19), .ZN(n1277) );
XOR2_X1 U982 ( .A(KEYINPUT52), .B(n1279), .Z(n1275) );
NOR2_X1 U983 ( .A1(G134), .A2(n1278), .ZN(n1279) );
NOR2_X1 U984 ( .A1(n1280), .A2(n1281), .ZN(n1278) );
AND2_X1 U985 ( .A1(n1282), .A2(G143), .ZN(n1281) );
XNOR2_X1 U986 ( .A(G128), .B(KEYINPUT17), .ZN(n1282) );
XNOR2_X1 U987 ( .A(G107), .B(n1283), .ZN(n1269) );
XOR2_X1 U988 ( .A(G122), .B(G116), .Z(n1283) );
XNOR2_X1 U989 ( .A(n1284), .B(G475), .ZN(n1087) );
NAND2_X1 U990 ( .A1(n1143), .A2(n1182), .ZN(n1284) );
XOR2_X1 U991 ( .A(n1285), .B(n1286), .Z(n1143) );
XOR2_X1 U992 ( .A(n1287), .B(n1288), .Z(n1286) );
XNOR2_X1 U993 ( .A(G113), .B(G143), .ZN(n1288) );
NAND2_X1 U994 ( .A1(G214), .A2(n1289), .ZN(n1287) );
XOR2_X1 U995 ( .A(n1096), .B(n1290), .Z(n1285) );
XOR2_X1 U996 ( .A(n1291), .B(n1292), .Z(n1290) );
NOR2_X1 U997 ( .A1(KEYINPUT38), .A2(n1293), .ZN(n1291) );
XOR2_X1 U998 ( .A(n1294), .B(n1295), .Z(n1096) );
AND3_X1 U999 ( .A1(n1072), .A2(n1228), .A3(n1063), .ZN(n1190) );
INV_X1 U1000 ( .A(n1227), .ZN(n1063) );
NAND2_X1 U1001 ( .A1(n1064), .A2(n1065), .ZN(n1227) );
NAND2_X1 U1002 ( .A1(G214), .A2(n1296), .ZN(n1065) );
XNOR2_X1 U1003 ( .A(n1086), .B(KEYINPUT39), .ZN(n1064) );
XNOR2_X1 U1004 ( .A(n1297), .B(n1181), .ZN(n1086) );
AND2_X1 U1005 ( .A1(G210), .A2(n1296), .ZN(n1181) );
NAND2_X1 U1006 ( .A1(n1298), .A2(n1182), .ZN(n1296) );
XOR2_X1 U1007 ( .A(KEYINPUT15), .B(G237), .Z(n1298) );
NAND2_X1 U1008 ( .A1(n1299), .A2(n1300), .ZN(n1297) );
XNOR2_X1 U1009 ( .A(KEYINPUT60), .B(n1182), .ZN(n1300) );
XOR2_X1 U1010 ( .A(n1121), .B(n1301), .Z(n1299) );
XNOR2_X1 U1011 ( .A(n1180), .B(n1302), .ZN(n1301) );
NAND3_X1 U1012 ( .A1(KEYINPUT26), .A2(n1303), .A3(n1304), .ZN(n1302) );
XOR2_X1 U1013 ( .A(n1305), .B(KEYINPUT23), .Z(n1304) );
OR2_X1 U1014 ( .A1(n1161), .A2(G125), .ZN(n1305) );
NAND2_X1 U1015 ( .A1(G125), .A2(n1161), .ZN(n1303) );
NOR2_X1 U1016 ( .A1(n1106), .A2(G953), .ZN(n1180) );
INV_X1 U1017 ( .A(G224), .ZN(n1106) );
XOR2_X1 U1018 ( .A(n1306), .B(n1307), .Z(n1121) );
XOR2_X1 U1019 ( .A(n1308), .B(n1292), .Z(n1307) );
XNOR2_X1 U1020 ( .A(n1309), .B(G122), .ZN(n1292) );
XNOR2_X1 U1021 ( .A(n1149), .B(n1310), .ZN(n1306) );
NAND2_X1 U1022 ( .A1(n1311), .A2(n1312), .ZN(n1228) );
NAND3_X1 U1023 ( .A1(n1120), .A2(n1313), .A3(G902), .ZN(n1312) );
XNOR2_X1 U1024 ( .A(KEYINPUT13), .B(n1233), .ZN(n1313) );
NOR2_X1 U1025 ( .A1(n1100), .A2(G898), .ZN(n1120) );
XNOR2_X1 U1026 ( .A(KEYINPUT49), .B(n1048), .ZN(n1311) );
NAND3_X1 U1027 ( .A1(n1233), .A2(n1100), .A3(G952), .ZN(n1048) );
NAND2_X1 U1028 ( .A1(G237), .A2(G234), .ZN(n1233) );
NAND2_X1 U1029 ( .A1(n1314), .A2(n1315), .ZN(n1072) );
NAND3_X1 U1030 ( .A1(n1073), .A2(n1074), .A3(n1316), .ZN(n1315) );
INV_X1 U1031 ( .A(KEYINPUT28), .ZN(n1316) );
NAND2_X1 U1032 ( .A1(KEYINPUT28), .A2(n1231), .ZN(n1314) );
INV_X1 U1033 ( .A(n1057), .ZN(n1231) );
NAND2_X1 U1034 ( .A1(n1317), .A2(n1074), .ZN(n1057) );
NAND2_X1 U1035 ( .A1(G221), .A2(n1318), .ZN(n1074) );
INV_X1 U1036 ( .A(n1073), .ZN(n1317) );
XNOR2_X1 U1037 ( .A(n1319), .B(G469), .ZN(n1073) );
NAND2_X1 U1038 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
XNOR2_X1 U1039 ( .A(KEYINPUT45), .B(n1182), .ZN(n1321) );
XOR2_X1 U1040 ( .A(n1322), .B(n1170), .Z(n1320) );
XNOR2_X1 U1041 ( .A(n1323), .B(n1324), .ZN(n1170) );
XNOR2_X1 U1042 ( .A(n1325), .B(n1326), .ZN(n1324) );
AND2_X1 U1043 ( .A1(n1100), .A2(G227), .ZN(n1325) );
XNOR2_X1 U1044 ( .A(G110), .B(n1327), .ZN(n1323) );
XOR2_X1 U1045 ( .A(KEYINPUT25), .B(G140), .Z(n1327) );
NAND3_X1 U1046 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1322) );
NAND2_X1 U1047 ( .A1(n1171), .A2(n1173), .ZN(n1330) );
INV_X1 U1048 ( .A(n1331), .ZN(n1173) );
INV_X1 U1049 ( .A(n1095), .ZN(n1171) );
NAND2_X1 U1050 ( .A1(KEYINPUT20), .A2(n1332), .ZN(n1329) );
NAND2_X1 U1051 ( .A1(n1333), .A2(n1331), .ZN(n1332) );
XNOR2_X1 U1052 ( .A(n1095), .B(KEYINPUT4), .ZN(n1333) );
NAND2_X1 U1053 ( .A1(n1334), .A2(n1335), .ZN(n1328) );
INV_X1 U1054 ( .A(KEYINPUT20), .ZN(n1335) );
NAND2_X1 U1055 ( .A1(n1336), .A2(n1337), .ZN(n1334) );
OR2_X1 U1056 ( .A1(n1095), .A2(KEYINPUT4), .ZN(n1337) );
NAND3_X1 U1057 ( .A1(n1331), .A2(n1095), .A3(KEYINPUT4), .ZN(n1336) );
XOR2_X1 U1058 ( .A(n1338), .B(n1293), .Z(n1095) );
NAND2_X1 U1059 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
NAND2_X1 U1060 ( .A1(G143), .A2(n1341), .ZN(n1340) );
NAND2_X1 U1061 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NAND2_X1 U1062 ( .A1(n1280), .A2(n1342), .ZN(n1339) );
INV_X1 U1063 ( .A(KEYINPUT35), .ZN(n1342) );
XNOR2_X1 U1064 ( .A(n1344), .B(n1308), .ZN(n1331) );
XNOR2_X1 U1065 ( .A(G107), .B(n1153), .ZN(n1308) );
NAND2_X1 U1066 ( .A1(KEYINPUT48), .A2(n1309), .ZN(n1344) );
INV_X1 U1067 ( .A(G104), .ZN(n1309) );
NOR2_X1 U1068 ( .A1(n1224), .A2(n1239), .ZN(n1068) );
INV_X1 U1069 ( .A(n1223), .ZN(n1239) );
XNOR2_X1 U1070 ( .A(n1081), .B(n1345), .ZN(n1223) );
XOR2_X1 U1071 ( .A(KEYINPUT55), .B(KEYINPUT51), .Z(n1345) );
XOR2_X1 U1072 ( .A(n1346), .B(n1132), .Z(n1081) );
AND2_X1 U1073 ( .A1(G217), .A2(n1318), .ZN(n1132) );
NAND2_X1 U1074 ( .A1(G234), .A2(n1182), .ZN(n1318) );
NAND2_X1 U1075 ( .A1(n1130), .A2(n1182), .ZN(n1346) );
XOR2_X1 U1076 ( .A(n1347), .B(n1348), .Z(n1130) );
XOR2_X1 U1077 ( .A(n1349), .B(n1350), .Z(n1348) );
NAND2_X1 U1078 ( .A1(n1351), .A2(KEYINPUT61), .ZN(n1350) );
XNOR2_X1 U1079 ( .A(n1352), .B(n1353), .ZN(n1351) );
XOR2_X1 U1080 ( .A(KEYINPUT42), .B(n1295), .Z(n1353) );
XOR2_X1 U1081 ( .A(G125), .B(G140), .Z(n1295) );
NAND2_X1 U1082 ( .A1(G221), .A2(n1273), .ZN(n1349) );
AND2_X1 U1083 ( .A1(G234), .A2(n1100), .ZN(n1273) );
INV_X1 U1084 ( .A(G953), .ZN(n1100) );
XOR2_X1 U1085 ( .A(n1354), .B(n1355), .Z(n1347) );
XNOR2_X1 U1086 ( .A(G137), .B(n1310), .ZN(n1355) );
INV_X1 U1087 ( .A(G110), .ZN(n1310) );
NAND2_X1 U1088 ( .A1(n1356), .A2(n1357), .ZN(n1354) );
NAND2_X1 U1089 ( .A1(G119), .A2(n1343), .ZN(n1357) );
INV_X1 U1090 ( .A(G128), .ZN(n1343) );
XOR2_X1 U1091 ( .A(n1358), .B(KEYINPUT34), .Z(n1356) );
NAND2_X1 U1092 ( .A1(G128), .A2(n1243), .ZN(n1358) );
XNOR2_X1 U1093 ( .A(n1359), .B(G472), .ZN(n1224) );
NAND2_X1 U1094 ( .A1(n1360), .A2(n1182), .ZN(n1359) );
INV_X1 U1095 ( .A(G902), .ZN(n1182) );
XOR2_X1 U1096 ( .A(n1361), .B(n1362), .Z(n1360) );
XOR2_X1 U1097 ( .A(n1363), .B(n1149), .Z(n1362) );
XNOR2_X1 U1098 ( .A(G113), .B(n1364), .ZN(n1149) );
XNOR2_X1 U1099 ( .A(n1243), .B(G116), .ZN(n1364) );
INV_X1 U1100 ( .A(G119), .ZN(n1243) );
NAND2_X1 U1101 ( .A1(KEYINPUT21), .A2(n1152), .ZN(n1363) );
NAND2_X1 U1102 ( .A1(G210), .A2(n1289), .ZN(n1152) );
NOR2_X1 U1103 ( .A1(G953), .A2(G237), .ZN(n1289) );
XNOR2_X1 U1104 ( .A(n1153), .B(n1365), .ZN(n1361) );
NOR2_X1 U1105 ( .A1(KEYINPUT0), .A2(n1366), .ZN(n1365) );
XNOR2_X1 U1106 ( .A(n1161), .B(n1326), .ZN(n1366) );
INV_X1 U1107 ( .A(n1158), .ZN(n1326) );
XNOR2_X1 U1108 ( .A(n1294), .B(n1367), .ZN(n1158) );
XOR2_X1 U1109 ( .A(G134), .B(n1368), .Z(n1367) );
NOR2_X1 U1110 ( .A1(G137), .A2(KEYINPUT18), .ZN(n1368) );
XNOR2_X1 U1111 ( .A(G131), .B(KEYINPUT14), .ZN(n1294) );
XOR2_X1 U1112 ( .A(n1369), .B(n1293), .Z(n1161) );
INV_X1 U1113 ( .A(n1352), .ZN(n1293) );
XOR2_X1 U1114 ( .A(G146), .B(KEYINPUT3), .Z(n1352) );
NAND2_X1 U1115 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
NAND2_X1 U1116 ( .A1(G128), .A2(n1372), .ZN(n1371) );
OR2_X1 U1117 ( .A1(KEYINPUT57), .A2(G143), .ZN(n1372) );
NAND2_X1 U1118 ( .A1(n1280), .A2(n1373), .ZN(n1370) );
INV_X1 U1119 ( .A(KEYINPUT57), .ZN(n1373) );
NOR2_X1 U1120 ( .A1(G128), .A2(G143), .ZN(n1280) );
INV_X1 U1121 ( .A(G101), .ZN(n1153) );
endmodule


