//Key = 1111010011111001100011101100110110011010100000111001111111100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346;

XNOR2_X1 U729 ( .A(G107), .B(n1019), .ZN(G9) );
NOR2_X1 U730 ( .A1(n1020), .A2(n1021), .ZN(G75) );
NOR4_X1 U731 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1021) );
NAND3_X1 U732 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1022) );
XNOR2_X1 U733 ( .A(KEYINPUT13), .B(n1029), .ZN(n1028) );
NAND2_X1 U734 ( .A1(n1030), .A2(n1031), .ZN(n1026) );
NAND2_X1 U735 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND3_X1 U736 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NAND2_X1 U737 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NAND2_X1 U738 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
OR2_X1 U739 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U740 ( .A1(n1043), .A2(n1044), .ZN(n1037) );
NAND2_X1 U741 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U742 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U743 ( .A1(n1039), .A2(n1049), .A3(n1043), .ZN(n1032) );
NAND2_X1 U744 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U745 ( .A1(n1034), .A2(n1052), .ZN(n1051) );
NAND2_X1 U746 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U747 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
INV_X1 U748 ( .A(n1057), .ZN(n1053) );
NAND2_X1 U749 ( .A1(n1036), .A2(n1058), .ZN(n1050) );
NAND2_X1 U750 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U751 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR3_X1 U752 ( .A1(n1025), .A2(G952), .A3(n1063), .ZN(n1020) );
INV_X1 U753 ( .A(n1027), .ZN(n1063) );
NAND4_X1 U754 ( .A1(n1064), .A2(n1039), .A3(n1065), .A4(n1066), .ZN(n1027) );
NOR4_X1 U755 ( .A1(n1067), .A2(n1061), .A3(n1068), .A4(n1069), .ZN(n1066) );
XOR2_X1 U756 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND2_X1 U757 ( .A1(KEYINPUT10), .A2(n1072), .ZN(n1070) );
NOR2_X1 U758 ( .A1(n1073), .A2(n1074), .ZN(n1068) );
XOR2_X1 U759 ( .A(n1075), .B(KEYINPUT29), .Z(n1073) );
NOR2_X1 U760 ( .A1(n1076), .A2(n1077), .ZN(n1065) );
XNOR2_X1 U761 ( .A(G478), .B(n1078), .ZN(n1077) );
XOR2_X1 U762 ( .A(n1079), .B(n1080), .Z(n1076) );
XNOR2_X1 U763 ( .A(G472), .B(n1081), .ZN(n1064) );
NOR2_X1 U764 ( .A1(KEYINPUT50), .A2(n1082), .ZN(n1081) );
XOR2_X1 U765 ( .A(n1083), .B(n1084), .Z(G72) );
XOR2_X1 U766 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U767 ( .A1(G953), .A2(n1087), .ZN(n1086) );
NAND2_X1 U768 ( .A1(G900), .A2(G227), .ZN(n1087) );
NAND2_X1 U769 ( .A1(n1088), .A2(n1089), .ZN(n1085) );
NAND2_X1 U770 ( .A1(G953), .A2(n1090), .ZN(n1089) );
XOR2_X1 U771 ( .A(n1091), .B(n1092), .Z(n1088) );
XNOR2_X1 U772 ( .A(n1093), .B(n1094), .ZN(n1092) );
NAND2_X1 U773 ( .A1(KEYINPUT25), .A2(n1095), .ZN(n1093) );
XOR2_X1 U774 ( .A(n1096), .B(n1097), .Z(n1091) );
XNOR2_X1 U775 ( .A(n1098), .B(G131), .ZN(n1097) );
NAND3_X1 U776 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1096) );
NAND2_X1 U777 ( .A1(KEYINPUT7), .A2(G134), .ZN(n1101) );
NAND3_X1 U778 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1100) );
INV_X1 U779 ( .A(KEYINPUT7), .ZN(n1103) );
OR2_X1 U780 ( .A1(n1104), .A2(n1102), .ZN(n1099) );
NOR2_X1 U781 ( .A1(G134), .A2(KEYINPUT43), .ZN(n1102) );
XNOR2_X1 U782 ( .A(n1105), .B(KEYINPUT48), .ZN(n1104) );
AND2_X1 U783 ( .A1(n1029), .A2(n1106), .ZN(n1083) );
XOR2_X1 U784 ( .A(n1107), .B(n1108), .Z(G69) );
XOR2_X1 U785 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U786 ( .A1(G953), .A2(n1111), .ZN(n1110) );
NOR2_X1 U787 ( .A1(n1112), .A2(n1024), .ZN(n1111) );
XOR2_X1 U788 ( .A(n1023), .B(KEYINPUT49), .Z(n1112) );
NAND2_X1 U789 ( .A1(n1113), .A2(n1114), .ZN(n1109) );
NAND2_X1 U790 ( .A1(G953), .A2(n1115), .ZN(n1114) );
XNOR2_X1 U791 ( .A(n1116), .B(n1117), .ZN(n1113) );
NAND2_X1 U792 ( .A1(G953), .A2(n1118), .ZN(n1107) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1118) );
NOR3_X1 U794 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(G66) );
AND2_X1 U795 ( .A1(KEYINPUT22), .A2(n1122), .ZN(n1121) );
NOR3_X1 U796 ( .A1(KEYINPUT22), .A2(G953), .A3(G952), .ZN(n1120) );
XOR2_X1 U797 ( .A(n1123), .B(n1124), .Z(n1119) );
XNOR2_X1 U798 ( .A(KEYINPUT27), .B(n1125), .ZN(n1124) );
NOR3_X1 U799 ( .A1(n1126), .A2(KEYINPUT44), .A3(n1127), .ZN(n1123) );
INV_X1 U800 ( .A(G217), .ZN(n1127) );
NOR2_X1 U801 ( .A1(n1122), .A2(n1128), .ZN(G63) );
XNOR2_X1 U802 ( .A(n1129), .B(n1130), .ZN(n1128) );
NAND2_X1 U803 ( .A1(n1131), .A2(G478), .ZN(n1129) );
NOR2_X1 U804 ( .A1(n1122), .A2(n1132), .ZN(G60) );
XOR2_X1 U805 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U806 ( .A1(n1131), .A2(G475), .ZN(n1133) );
XNOR2_X1 U807 ( .A(G104), .B(n1135), .ZN(G6) );
NOR2_X1 U808 ( .A1(n1122), .A2(n1136), .ZN(G57) );
XOR2_X1 U809 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U810 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U811 ( .A1(KEYINPUT36), .A2(n1141), .ZN(n1140) );
NAND2_X1 U812 ( .A1(n1131), .A2(G472), .ZN(n1139) );
XNOR2_X1 U813 ( .A(n1142), .B(n1143), .ZN(n1137) );
NAND2_X1 U814 ( .A1(n1144), .A2(n1145), .ZN(n1142) );
XOR2_X1 U815 ( .A(KEYINPUT57), .B(KEYINPUT30), .Z(n1145) );
XNOR2_X1 U816 ( .A(n1146), .B(n1147), .ZN(n1144) );
NOR2_X1 U817 ( .A1(n1122), .A2(n1148), .ZN(G54) );
XOR2_X1 U818 ( .A(n1149), .B(n1150), .Z(n1148) );
NAND2_X1 U819 ( .A1(n1131), .A2(G469), .ZN(n1150) );
NAND2_X1 U820 ( .A1(n1151), .A2(KEYINPUT9), .ZN(n1149) );
XOR2_X1 U821 ( .A(n1152), .B(n1153), .Z(n1151) );
XNOR2_X1 U822 ( .A(n1154), .B(n1155), .ZN(n1153) );
NAND2_X1 U823 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
OR2_X1 U824 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U825 ( .A(n1160), .B(KEYINPUT6), .Z(n1156) );
NAND2_X1 U826 ( .A1(n1158), .A2(n1159), .ZN(n1160) );
XNOR2_X1 U827 ( .A(G110), .B(n1161), .ZN(n1152) );
XNOR2_X1 U828 ( .A(KEYINPUT63), .B(n1098), .ZN(n1161) );
NOR2_X1 U829 ( .A1(n1122), .A2(n1162), .ZN(G51) );
XOR2_X1 U830 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U831 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND2_X1 U832 ( .A1(n1131), .A2(n1079), .ZN(n1166) );
INV_X1 U833 ( .A(n1126), .ZN(n1131) );
NAND2_X1 U834 ( .A1(G902), .A2(n1167), .ZN(n1126) );
OR3_X1 U835 ( .A1(n1024), .A2(n1029), .A3(n1023), .ZN(n1167) );
NAND4_X1 U836 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1023) );
NAND4_X1 U837 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1029) );
NOR4_X1 U838 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1175) );
NOR2_X1 U839 ( .A1(n1180), .A2(n1181), .ZN(n1174) );
NAND3_X1 U840 ( .A1(n1041), .A2(n1182), .A3(n1183), .ZN(n1172) );
NAND4_X1 U841 ( .A1(n1184), .A2(n1135), .A3(n1185), .A4(n1019), .ZN(n1024) );
NAND3_X1 U842 ( .A1(n1036), .A2(n1186), .A3(n1042), .ZN(n1019) );
NAND3_X1 U843 ( .A1(n1036), .A2(n1186), .A3(n1041), .ZN(n1135) );
NAND2_X1 U844 ( .A1(n1187), .A2(n1188), .ZN(n1184) );
XOR2_X1 U845 ( .A(KEYINPUT14), .B(n1189), .Z(n1188) );
NAND2_X1 U846 ( .A1(n1190), .A2(n1191), .ZN(n1165) );
NAND2_X1 U847 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U848 ( .A(n1194), .B(KEYINPUT39), .Z(n1190) );
NAND2_X1 U849 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XOR2_X1 U850 ( .A(KEYINPUT56), .B(n1193), .Z(n1195) );
NOR2_X1 U851 ( .A1(n1106), .A2(G952), .ZN(n1122) );
XNOR2_X1 U852 ( .A(G146), .B(n1197), .ZN(G48) );
NAND4_X1 U853 ( .A1(KEYINPUT40), .A2(n1183), .A3(n1041), .A4(n1182), .ZN(n1197) );
XNOR2_X1 U854 ( .A(G143), .B(n1173), .ZN(G45) );
NAND4_X1 U855 ( .A1(n1198), .A2(n1199), .A3(n1182), .A4(n1200), .ZN(n1173) );
XOR2_X1 U856 ( .A(n1181), .B(n1201), .Z(G42) );
XNOR2_X1 U857 ( .A(KEYINPUT34), .B(n1098), .ZN(n1201) );
AND3_X1 U858 ( .A1(n1202), .A2(n1034), .A3(n1203), .ZN(n1181) );
XOR2_X1 U859 ( .A(G137), .B(n1180), .Z(G39) );
AND3_X1 U860 ( .A1(n1043), .A2(n1034), .A3(n1183), .ZN(n1180) );
XNOR2_X1 U861 ( .A(n1204), .B(n1177), .ZN(G36) );
AND3_X1 U862 ( .A1(n1042), .A2(n1034), .A3(n1199), .ZN(n1177) );
XNOR2_X1 U863 ( .A(n1205), .B(n1176), .ZN(G33) );
AND3_X1 U864 ( .A1(n1041), .A2(n1034), .A3(n1199), .ZN(n1176) );
AND3_X1 U865 ( .A1(n1202), .A2(n1206), .A3(n1057), .ZN(n1199) );
NAND2_X1 U866 ( .A1(n1207), .A2(n1208), .ZN(n1034) );
OR2_X1 U867 ( .A1(n1209), .A2(KEYINPUT0), .ZN(n1208) );
NAND3_X1 U868 ( .A1(n1062), .A2(n1210), .A3(KEYINPUT0), .ZN(n1207) );
XOR2_X1 U869 ( .A(n1211), .B(n1179), .Z(G30) );
AND3_X1 U870 ( .A1(n1042), .A2(n1182), .A3(n1183), .ZN(n1179) );
AND4_X1 U871 ( .A1(n1202), .A2(n1212), .A3(n1056), .A4(n1206), .ZN(n1183) );
NAND2_X1 U872 ( .A1(KEYINPUT12), .A2(n1213), .ZN(n1211) );
XNOR2_X1 U873 ( .A(G101), .B(n1185), .ZN(G3) );
NAND3_X1 U874 ( .A1(n1057), .A2(n1186), .A3(n1043), .ZN(n1185) );
NOR3_X1 U875 ( .A1(n1045), .A2(n1214), .A3(n1209), .ZN(n1186) );
INV_X1 U876 ( .A(n1202), .ZN(n1045) );
XNOR2_X1 U877 ( .A(n1095), .B(n1178), .ZN(G27) );
AND3_X1 U878 ( .A1(n1039), .A2(n1182), .A3(n1203), .ZN(n1178) );
AND4_X1 U879 ( .A1(n1055), .A2(n1041), .A3(n1056), .A4(n1206), .ZN(n1203) );
NAND2_X1 U880 ( .A1(n1215), .A2(n1216), .ZN(n1206) );
NAND2_X1 U881 ( .A1(n1217), .A2(n1090), .ZN(n1216) );
INV_X1 U882 ( .A(G900), .ZN(n1090) );
INV_X1 U883 ( .A(n1218), .ZN(n1039) );
INV_X1 U884 ( .A(G125), .ZN(n1095) );
XOR2_X1 U885 ( .A(n1168), .B(n1219), .Z(G24) );
XNOR2_X1 U886 ( .A(KEYINPUT46), .B(n1220), .ZN(n1219) );
NAND4_X1 U887 ( .A1(n1221), .A2(n1036), .A3(n1198), .A4(n1200), .ZN(n1168) );
NOR2_X1 U888 ( .A1(n1056), .A2(n1212), .ZN(n1036) );
XNOR2_X1 U889 ( .A(G119), .B(n1169), .ZN(G21) );
NAND4_X1 U890 ( .A1(n1043), .A2(n1221), .A3(n1212), .A4(n1056), .ZN(n1169) );
XNOR2_X1 U891 ( .A(G116), .B(n1170), .ZN(G18) );
NAND3_X1 U892 ( .A1(n1057), .A2(n1042), .A3(n1221), .ZN(n1170) );
NOR3_X1 U893 ( .A1(n1059), .A2(n1214), .A3(n1218), .ZN(n1221) );
INV_X1 U894 ( .A(n1182), .ZN(n1059) );
XOR2_X1 U895 ( .A(n1187), .B(KEYINPUT45), .Z(n1182) );
AND2_X1 U896 ( .A1(n1222), .A2(n1198), .ZN(n1042) );
XOR2_X1 U897 ( .A(n1171), .B(n1223), .Z(G15) );
XNOR2_X1 U898 ( .A(KEYINPUT8), .B(n1224), .ZN(n1223) );
NAND3_X1 U899 ( .A1(n1057), .A2(n1041), .A3(n1225), .ZN(n1171) );
NOR3_X1 U900 ( .A1(n1218), .A2(n1214), .A3(n1209), .ZN(n1225) );
INV_X1 U901 ( .A(n1187), .ZN(n1209) );
INV_X1 U902 ( .A(n1226), .ZN(n1214) );
NAND2_X1 U903 ( .A1(n1048), .A2(n1227), .ZN(n1218) );
NOR2_X1 U904 ( .A1(n1198), .A2(n1222), .ZN(n1041) );
NOR2_X1 U905 ( .A1(n1056), .A2(n1055), .ZN(n1057) );
XNOR2_X1 U906 ( .A(G110), .B(n1228), .ZN(G12) );
NAND2_X1 U907 ( .A1(n1189), .A2(n1187), .ZN(n1228) );
NOR2_X1 U908 ( .A1(n1062), .A2(n1061), .ZN(n1187) );
INV_X1 U909 ( .A(n1210), .ZN(n1061) );
NAND2_X1 U910 ( .A1(G214), .A2(n1229), .ZN(n1210) );
XOR2_X1 U911 ( .A(n1079), .B(n1230), .Z(n1062) );
NOR2_X1 U912 ( .A1(n1080), .A2(KEYINPUT37), .ZN(n1230) );
AND3_X1 U913 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1080) );
NAND2_X1 U914 ( .A1(n1234), .A2(n1192), .ZN(n1232) );
INV_X1 U915 ( .A(n1196), .ZN(n1192) );
NAND2_X1 U916 ( .A1(n1235), .A2(n1196), .ZN(n1231) );
XNOR2_X1 U917 ( .A(G125), .B(n1094), .ZN(n1196) );
XNOR2_X1 U918 ( .A(n1234), .B(KEYINPUT23), .ZN(n1235) );
XOR2_X1 U919 ( .A(n1163), .B(n1236), .Z(n1234) );
XOR2_X1 U920 ( .A(KEYINPUT28), .B(n1193), .Z(n1236) );
AND2_X1 U921 ( .A1(G224), .A2(n1106), .ZN(n1193) );
XOR2_X1 U922 ( .A(n1237), .B(n1238), .Z(n1163) );
INV_X1 U923 ( .A(n1116), .ZN(n1238) );
XNOR2_X1 U924 ( .A(n1239), .B(n1240), .ZN(n1116) );
XNOR2_X1 U925 ( .A(n1241), .B(G101), .ZN(n1240) );
INV_X1 U926 ( .A(G110), .ZN(n1241) );
XOR2_X1 U927 ( .A(n1242), .B(n1243), .Z(n1239) );
NAND2_X1 U928 ( .A1(KEYINPUT38), .A2(n1220), .ZN(n1242) );
NAND2_X1 U929 ( .A1(KEYINPUT52), .A2(n1117), .ZN(n1237) );
XNOR2_X1 U930 ( .A(n1244), .B(n1245), .ZN(n1117) );
XNOR2_X1 U931 ( .A(n1246), .B(G113), .ZN(n1245) );
NAND2_X1 U932 ( .A1(KEYINPUT5), .A2(n1247), .ZN(n1244) );
AND2_X1 U933 ( .A1(G210), .A2(n1229), .ZN(n1079) );
NAND2_X1 U934 ( .A1(n1248), .A2(n1233), .ZN(n1229) );
INV_X1 U935 ( .A(G237), .ZN(n1248) );
AND4_X1 U936 ( .A1(n1043), .A2(n1202), .A3(n1249), .A4(n1055), .ZN(n1189) );
INV_X1 U937 ( .A(n1212), .ZN(n1055) );
XNOR2_X1 U938 ( .A(G472), .B(n1082), .ZN(n1212) );
NAND2_X1 U939 ( .A1(n1250), .A2(n1233), .ZN(n1082) );
XOR2_X1 U940 ( .A(KEYINPUT3), .B(n1251), .Z(n1250) );
NOR3_X1 U941 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1251) );
NOR2_X1 U942 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
INV_X1 U943 ( .A(n1257), .ZN(n1256) );
NOR2_X1 U944 ( .A1(n1258), .A2(n1259), .ZN(n1255) );
XOR2_X1 U945 ( .A(KEYINPUT59), .B(n1260), .Z(n1259) );
NOR3_X1 U946 ( .A1(n1257), .A2(n1260), .A3(n1258), .ZN(n1253) );
XOR2_X1 U947 ( .A(n1143), .B(n1141), .Z(n1257) );
NAND2_X1 U948 ( .A1(n1261), .A2(n1262), .ZN(n1143) );
XNOR2_X1 U949 ( .A(G210), .B(KEYINPUT2), .ZN(n1261) );
AND2_X1 U950 ( .A1(n1258), .A2(n1260), .ZN(n1252) );
XNOR2_X1 U951 ( .A(n1263), .B(n1147), .ZN(n1260) );
XNOR2_X1 U952 ( .A(n1264), .B(n1159), .ZN(n1147) );
NAND2_X1 U953 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NAND2_X1 U954 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
XNOR2_X1 U955 ( .A(n1269), .B(n1246), .ZN(n1268) );
XNOR2_X1 U956 ( .A(G113), .B(KEYINPUT11), .ZN(n1267) );
XOR2_X1 U957 ( .A(n1270), .B(KEYINPUT41), .Z(n1265) );
NAND2_X1 U958 ( .A1(n1271), .A2(n1224), .ZN(n1270) );
INV_X1 U959 ( .A(G113), .ZN(n1224) );
XNOR2_X1 U960 ( .A(G119), .B(n1269), .ZN(n1271) );
NAND2_X1 U961 ( .A1(KEYINPUT35), .A2(n1247), .ZN(n1269) );
XNOR2_X1 U962 ( .A(KEYINPUT17), .B(n1272), .ZN(n1263) );
NOR2_X1 U963 ( .A1(KEYINPUT18), .A2(n1146), .ZN(n1272) );
INV_X1 U964 ( .A(KEYINPUT58), .ZN(n1258) );
AND2_X1 U965 ( .A1(n1226), .A2(n1056), .ZN(n1249) );
XNOR2_X1 U966 ( .A(n1273), .B(n1071), .ZN(n1056) );
AND2_X1 U967 ( .A1(G217), .A2(n1274), .ZN(n1071) );
NAND2_X1 U968 ( .A1(KEYINPUT21), .A2(n1275), .ZN(n1273) );
INV_X1 U969 ( .A(n1072), .ZN(n1275) );
NAND2_X1 U970 ( .A1(n1233), .A2(n1125), .ZN(n1072) );
NAND2_X1 U971 ( .A1(n1276), .A2(n1277), .ZN(n1125) );
NAND2_X1 U972 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
XOR2_X1 U973 ( .A(KEYINPUT47), .B(n1280), .Z(n1276) );
NOR2_X1 U974 ( .A1(n1278), .A2(n1279), .ZN(n1280) );
XNOR2_X1 U975 ( .A(n1281), .B(n1282), .ZN(n1279) );
XOR2_X1 U976 ( .A(n1283), .B(n1284), .Z(n1282) );
XNOR2_X1 U977 ( .A(G110), .B(G125), .ZN(n1284) );
NAND2_X1 U978 ( .A1(KEYINPUT53), .A2(n1098), .ZN(n1283) );
XOR2_X1 U979 ( .A(n1285), .B(n1286), .Z(n1281) );
NAND2_X1 U980 ( .A1(KEYINPUT31), .A2(n1246), .ZN(n1285) );
INV_X1 U981 ( .A(G119), .ZN(n1246) );
XNOR2_X1 U982 ( .A(n1287), .B(n1105), .ZN(n1278) );
NAND2_X1 U983 ( .A1(G221), .A2(n1288), .ZN(n1287) );
NAND2_X1 U984 ( .A1(n1215), .A2(n1289), .ZN(n1226) );
NAND2_X1 U985 ( .A1(n1217), .A2(n1115), .ZN(n1289) );
INV_X1 U986 ( .A(G898), .ZN(n1115) );
NOR3_X1 U987 ( .A1(n1233), .A2(n1290), .A3(n1106), .ZN(n1217) );
INV_X1 U988 ( .A(n1030), .ZN(n1215) );
NOR3_X1 U989 ( .A1(n1025), .A2(n1290), .A3(n1291), .ZN(n1030) );
INV_X1 U990 ( .A(G952), .ZN(n1291) );
AND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1290) );
XOR2_X1 U992 ( .A(G953), .B(KEYINPUT26), .Z(n1025) );
NOR2_X1 U993 ( .A1(n1048), .A2(n1047), .ZN(n1202) );
INV_X1 U994 ( .A(n1227), .ZN(n1047) );
NAND2_X1 U995 ( .A1(G221), .A2(n1274), .ZN(n1227) );
NAND2_X1 U996 ( .A1(G234), .A2(n1233), .ZN(n1274) );
XOR2_X1 U997 ( .A(n1292), .B(G469), .Z(n1048) );
NAND2_X1 U998 ( .A1(n1293), .A2(n1233), .ZN(n1292) );
XOR2_X1 U999 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U1000 ( .A(n1159), .B(n1158), .Z(n1295) );
XOR2_X1 U1001 ( .A(n1296), .B(n1094), .Z(n1158) );
INV_X1 U1002 ( .A(n1146), .ZN(n1094) );
XOR2_X1 U1003 ( .A(G143), .B(n1286), .Z(n1146) );
XNOR2_X1 U1004 ( .A(n1213), .B(G146), .ZN(n1286) );
NAND3_X1 U1005 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1296) );
NAND2_X1 U1006 ( .A1(KEYINPUT19), .A2(G101), .ZN(n1299) );
OR3_X1 U1007 ( .A1(G101), .A2(KEYINPUT19), .A3(n1243), .ZN(n1298) );
NAND2_X1 U1008 ( .A1(n1243), .A2(n1300), .ZN(n1297) );
NAND2_X1 U1009 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
INV_X1 U1010 ( .A(KEYINPUT19), .ZN(n1302) );
XNOR2_X1 U1011 ( .A(KEYINPUT20), .B(n1141), .ZN(n1301) );
INV_X1 U1012 ( .A(G101), .ZN(n1141) );
XOR2_X1 U1013 ( .A(G104), .B(G107), .Z(n1243) );
XOR2_X1 U1014 ( .A(n1303), .B(n1205), .Z(n1159) );
NAND2_X1 U1015 ( .A1(n1304), .A2(KEYINPUT32), .ZN(n1303) );
XNOR2_X1 U1016 ( .A(G134), .B(n1105), .ZN(n1304) );
XOR2_X1 U1017 ( .A(G137), .B(KEYINPUT15), .Z(n1105) );
XOR2_X1 U1018 ( .A(n1305), .B(n1306), .Z(n1294) );
NOR3_X1 U1019 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1306) );
NOR2_X1 U1020 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
INV_X1 U1021 ( .A(KEYINPUT51), .ZN(n1311) );
NOR2_X1 U1022 ( .A1(n1312), .A2(n1313), .ZN(n1310) );
NOR3_X1 U1023 ( .A1(n1098), .A2(KEYINPUT60), .A3(n1314), .ZN(n1313) );
AND2_X1 U1024 ( .A1(n1098), .A2(KEYINPUT60), .ZN(n1312) );
NOR2_X1 U1025 ( .A1(KEYINPUT51), .A2(n1315), .ZN(n1308) );
NOR2_X1 U1026 ( .A1(n1314), .A2(n1316), .ZN(n1315) );
XNOR2_X1 U1027 ( .A(KEYINPUT60), .B(G140), .ZN(n1316) );
AND2_X1 U1028 ( .A1(n1098), .A2(n1314), .ZN(n1307) );
XNOR2_X1 U1029 ( .A(G110), .B(KEYINPUT24), .ZN(n1314) );
NAND2_X1 U1030 ( .A1(KEYINPUT62), .A2(n1154), .ZN(n1305) );
AND2_X1 U1031 ( .A1(G227), .A2(n1106), .ZN(n1154) );
NOR2_X1 U1032 ( .A1(n1200), .A2(n1198), .ZN(n1043) );
XNOR2_X1 U1033 ( .A(n1317), .B(n1078), .ZN(n1198) );
NAND2_X1 U1034 ( .A1(n1318), .A2(n1233), .ZN(n1078) );
XNOR2_X1 U1035 ( .A(KEYINPUT55), .B(n1319), .ZN(n1318) );
INV_X1 U1036 ( .A(n1130), .ZN(n1319) );
XNOR2_X1 U1037 ( .A(n1320), .B(n1321), .ZN(n1130) );
XOR2_X1 U1038 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1039 ( .A(n1247), .B(G107), .ZN(n1323) );
INV_X1 U1040 ( .A(G116), .ZN(n1247) );
XNOR2_X1 U1041 ( .A(n1213), .B(G122), .ZN(n1322) );
INV_X1 U1042 ( .A(G128), .ZN(n1213) );
XOR2_X1 U1043 ( .A(n1324), .B(n1325), .Z(n1320) );
XNOR2_X1 U1044 ( .A(n1326), .B(n1327), .ZN(n1325) );
NOR2_X1 U1045 ( .A1(KEYINPUT33), .A2(n1204), .ZN(n1327) );
INV_X1 U1046 ( .A(G134), .ZN(n1204) );
NAND2_X1 U1047 ( .A1(KEYINPUT54), .A2(n1328), .ZN(n1326) );
NAND2_X1 U1048 ( .A1(G217), .A2(n1288), .ZN(n1324) );
AND2_X1 U1049 ( .A1(G234), .A2(n1106), .ZN(n1288) );
INV_X1 U1050 ( .A(G953), .ZN(n1106) );
NAND2_X1 U1051 ( .A1(KEYINPUT16), .A2(n1329), .ZN(n1317) );
INV_X1 U1052 ( .A(G478), .ZN(n1329) );
INV_X1 U1053 ( .A(n1222), .ZN(n1200) );
NOR2_X1 U1054 ( .A1(n1330), .A2(n1067), .ZN(n1222) );
NOR2_X1 U1055 ( .A1(n1075), .A2(G475), .ZN(n1067) );
AND2_X1 U1056 ( .A1(n1331), .A2(n1075), .ZN(n1330) );
NAND2_X1 U1057 ( .A1(n1134), .A2(n1233), .ZN(n1075) );
INV_X1 U1058 ( .A(G902), .ZN(n1233) );
XOR2_X1 U1059 ( .A(n1332), .B(n1333), .Z(n1134) );
NOR2_X1 U1060 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
XOR2_X1 U1061 ( .A(n1336), .B(KEYINPUT1), .Z(n1335) );
NAND2_X1 U1062 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
NOR2_X1 U1063 ( .A1(n1337), .A2(n1338), .ZN(n1334) );
XNOR2_X1 U1064 ( .A(G125), .B(n1339), .ZN(n1338) );
XNOR2_X1 U1065 ( .A(G146), .B(n1098), .ZN(n1339) );
INV_X1 U1066 ( .A(G140), .ZN(n1098) );
AND2_X1 U1067 ( .A1(n1340), .A2(n1341), .ZN(n1337) );
NAND2_X1 U1068 ( .A1(n1342), .A2(n1205), .ZN(n1341) );
XOR2_X1 U1069 ( .A(n1343), .B(KEYINPUT4), .Z(n1340) );
OR2_X1 U1070 ( .A1(n1205), .A2(n1342), .ZN(n1343) );
XOR2_X1 U1071 ( .A(n1344), .B(n1328), .Z(n1342) );
INV_X1 U1072 ( .A(G143), .ZN(n1328) );
NAND2_X1 U1073 ( .A1(G214), .A2(n1262), .ZN(n1344) );
NOR2_X1 U1074 ( .A1(G953), .A2(G237), .ZN(n1262) );
INV_X1 U1075 ( .A(G131), .ZN(n1205) );
NAND2_X1 U1076 ( .A1(n1345), .A2(KEYINPUT61), .ZN(n1332) );
XNOR2_X1 U1077 ( .A(G104), .B(n1346), .ZN(n1345) );
XNOR2_X1 U1078 ( .A(n1220), .B(G113), .ZN(n1346) );
INV_X1 U1079 ( .A(G122), .ZN(n1220) );
XNOR2_X1 U1080 ( .A(KEYINPUT42), .B(n1074), .ZN(n1331) );
INV_X1 U1081 ( .A(G475), .ZN(n1074) );
endmodule


