//Key = 0111101000001111001010101110111011111111100000110011010111010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370;

XOR2_X1 U758 ( .A(G107), .B(n1045), .Z(G9) );
NOR2_X1 U759 ( .A1(n1046), .A2(n1047), .ZN(G75) );
NOR3_X1 U760 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
NAND3_X1 U761 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1048) );
NAND2_X1 U762 ( .A1(n1054), .A2(n1055), .ZN(n1051) );
NAND2_X1 U763 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND4_X1 U764 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1057) );
NAND2_X1 U765 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND3_X1 U767 ( .A1(n1064), .A2(n1066), .A3(n1067), .ZN(n1056) );
NAND2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NAND2_X1 U769 ( .A1(n1059), .A2(n1070), .ZN(n1069) );
NAND2_X1 U770 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U771 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
INV_X1 U772 ( .A(KEYINPUT61), .ZN(n1074) );
NAND2_X1 U773 ( .A1(n1060), .A2(n1076), .ZN(n1071) );
NAND2_X1 U774 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U775 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U776 ( .A1(n1058), .A2(n1073), .ZN(n1068) );
NAND4_X1 U777 ( .A1(n1058), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1073) );
NAND2_X1 U778 ( .A1(n1059), .A2(n1084), .ZN(n1083) );
NAND2_X1 U779 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U780 ( .A1(KEYINPUT61), .A2(n1075), .ZN(n1086) );
NAND2_X1 U781 ( .A1(KEYINPUT56), .A2(n1087), .ZN(n1085) );
OR3_X1 U782 ( .A1(n1088), .A2(KEYINPUT56), .A3(n1059), .ZN(n1082) );
NAND2_X1 U783 ( .A1(n1060), .A2(n1089), .ZN(n1081) );
NAND2_X1 U784 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U786 ( .A(KEYINPUT36), .B(n1094), .ZN(n1090) );
INV_X1 U787 ( .A(n1095), .ZN(n1054) );
AND3_X1 U788 ( .A1(n1096), .A2(n1052), .A3(n1053), .ZN(n1046) );
NAND4_X1 U789 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1052) );
NOR4_X1 U790 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1100) );
NOR2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NOR2_X1 U792 ( .A1(G469), .A2(n1107), .ZN(n1103) );
NOR2_X1 U793 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U794 ( .A1(KEYINPUT13), .A2(n1110), .ZN(n1109) );
AND2_X1 U795 ( .A1(n1106), .A2(KEYINPUT13), .ZN(n1108) );
OR2_X1 U796 ( .A1(KEYINPUT48), .A2(n1110), .ZN(n1106) );
XNOR2_X1 U797 ( .A(n1111), .B(KEYINPUT0), .ZN(n1110) );
XNOR2_X1 U798 ( .A(n1112), .B(n1113), .ZN(n1102) );
NAND3_X1 U799 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1101) );
XOR2_X1 U800 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U801 ( .A1(KEYINPUT33), .A2(G472), .ZN(n1117) );
XOR2_X1 U802 ( .A(n1119), .B(KEYINPUT52), .Z(n1114) );
NAND2_X1 U803 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR3_X1 U804 ( .A1(n1092), .A2(n1122), .A3(n1079), .ZN(n1099) );
INV_X1 U805 ( .A(n1123), .ZN(n1122) );
OR2_X1 U806 ( .A1(n1121), .A2(n1120), .ZN(n1098) );
XNOR2_X1 U807 ( .A(n1124), .B(KEYINPUT37), .ZN(n1121) );
XNOR2_X1 U808 ( .A(KEYINPUT53), .B(n1125), .ZN(n1097) );
XNOR2_X1 U809 ( .A(n1049), .B(KEYINPUT15), .ZN(n1096) );
INV_X1 U810 ( .A(G952), .ZN(n1049) );
XOR2_X1 U811 ( .A(n1126), .B(n1127), .Z(G72) );
XOR2_X1 U812 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U813 ( .A1(n1130), .A2(G953), .ZN(n1129) );
AND2_X1 U814 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR2_X1 U815 ( .A1(n1133), .A2(n1134), .ZN(n1128) );
XOR2_X1 U816 ( .A(n1135), .B(n1136), .Z(n1134) );
XNOR2_X1 U817 ( .A(G140), .B(G125), .ZN(n1136) );
NOR2_X1 U818 ( .A1(G900), .A2(n1137), .ZN(n1133) );
NOR2_X1 U819 ( .A1(n1138), .A2(n1137), .ZN(n1126) );
NOR2_X1 U820 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U821 ( .A(n1141), .B(n1142), .Z(G69) );
XOR2_X1 U822 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U823 ( .A1(G953), .A2(n1145), .ZN(n1144) );
NAND2_X1 U824 ( .A1(G898), .A2(G224), .ZN(n1145) );
NAND2_X1 U825 ( .A1(n1146), .A2(n1147), .ZN(n1143) );
NAND2_X1 U826 ( .A1(G953), .A2(n1148), .ZN(n1147) );
XOR2_X1 U827 ( .A(n1149), .B(n1150), .Z(n1146) );
XOR2_X1 U828 ( .A(n1151), .B(n1152), .Z(n1150) );
XNOR2_X1 U829 ( .A(n1153), .B(n1154), .ZN(n1149) );
XOR2_X1 U830 ( .A(KEYINPUT9), .B(KEYINPUT19), .Z(n1154) );
NOR2_X1 U831 ( .A1(n1155), .A2(G953), .ZN(n1141) );
NOR2_X1 U832 ( .A1(n1156), .A2(n1157), .ZN(G66) );
XNOR2_X1 U833 ( .A(n1158), .B(n1159), .ZN(n1157) );
XNOR2_X1 U834 ( .A(KEYINPUT40), .B(n1160), .ZN(n1159) );
NOR4_X1 U835 ( .A1(KEYINPUT42), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1160) );
NOR2_X1 U836 ( .A1(n1156), .A2(n1164), .ZN(G63) );
XOR2_X1 U837 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND2_X1 U838 ( .A1(n1167), .A2(G478), .ZN(n1165) );
NOR2_X1 U839 ( .A1(n1168), .A2(n1169), .ZN(G60) );
XNOR2_X1 U840 ( .A(n1156), .B(KEYINPUT26), .ZN(n1169) );
NOR3_X1 U841 ( .A1(n1113), .A2(n1170), .A3(n1171), .ZN(n1168) );
AND3_X1 U842 ( .A1(n1172), .A2(G475), .A3(n1167), .ZN(n1171) );
NOR2_X1 U843 ( .A1(n1173), .A2(n1172), .ZN(n1170) );
AND2_X1 U844 ( .A1(n1050), .A2(G475), .ZN(n1173) );
XOR2_X1 U845 ( .A(n1174), .B(n1175), .Z(G6) );
NAND2_X1 U846 ( .A1(KEYINPUT3), .A2(G104), .ZN(n1175) );
NOR2_X1 U847 ( .A1(n1156), .A2(n1176), .ZN(G57) );
XOR2_X1 U848 ( .A(n1177), .B(n1178), .Z(n1176) );
NOR2_X1 U849 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NAND2_X1 U850 ( .A1(n1181), .A2(n1182), .ZN(n1177) );
NAND2_X1 U851 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XOR2_X1 U852 ( .A(n1185), .B(n1186), .Z(n1181) );
NOR2_X1 U853 ( .A1(n1183), .A2(n1184), .ZN(n1186) );
INV_X1 U854 ( .A(KEYINPUT39), .ZN(n1184) );
AND2_X1 U855 ( .A1(n1187), .A2(n1188), .ZN(n1183) );
NAND2_X1 U856 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U857 ( .A(KEYINPUT43), .B(n1191), .Z(n1189) );
OR2_X1 U858 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
NAND2_X1 U859 ( .A1(n1167), .A2(G472), .ZN(n1185) );
NOR2_X1 U860 ( .A1(n1156), .A2(n1192), .ZN(G54) );
XOR2_X1 U861 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U862 ( .A(n1195), .B(n1135), .Z(n1194) );
XOR2_X1 U863 ( .A(n1196), .B(n1197), .Z(n1135) );
XOR2_X1 U864 ( .A(n1198), .B(n1199), .Z(n1193) );
XOR2_X1 U865 ( .A(n1200), .B(KEYINPUT29), .Z(n1199) );
NAND2_X1 U866 ( .A1(KEYINPUT18), .A2(n1201), .ZN(n1200) );
NAND3_X1 U867 ( .A1(n1167), .A2(G469), .A3(KEYINPUT25), .ZN(n1198) );
NOR2_X1 U868 ( .A1(n1156), .A2(n1202), .ZN(G51) );
XOR2_X1 U869 ( .A(n1203), .B(n1204), .Z(n1202) );
NAND2_X1 U870 ( .A1(n1167), .A2(n1120), .ZN(n1204) );
INV_X1 U871 ( .A(n1163), .ZN(n1167) );
NAND2_X1 U872 ( .A1(G902), .A2(n1050), .ZN(n1163) );
NAND3_X1 U873 ( .A1(n1155), .A2(n1132), .A3(n1205), .ZN(n1050) );
XOR2_X1 U874 ( .A(n1131), .B(KEYINPUT31), .Z(n1205) );
AND4_X1 U875 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1132) );
AND3_X1 U876 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1209) );
NAND2_X1 U877 ( .A1(n1058), .A2(n1213), .ZN(n1208) );
NAND2_X1 U878 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND3_X1 U879 ( .A1(n1216), .A2(n1060), .A3(n1217), .ZN(n1215) );
XNOR2_X1 U880 ( .A(n1218), .B(KEYINPUT62), .ZN(n1214) );
AND4_X1 U881 ( .A1(n1174), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1155) );
NOR4_X1 U882 ( .A1(n1045), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1221) );
INV_X1 U883 ( .A(n1225), .ZN(n1224) );
AND3_X1 U884 ( .A1(n1067), .A2(n1226), .A3(n1075), .ZN(n1045) );
AND2_X1 U885 ( .A1(n1227), .A2(n1228), .ZN(n1220) );
NAND3_X1 U886 ( .A1(n1067), .A2(n1226), .A3(n1087), .ZN(n1174) );
NAND2_X1 U887 ( .A1(KEYINPUT1), .A2(n1229), .ZN(n1203) );
XOR2_X1 U888 ( .A(n1230), .B(n1231), .Z(n1229) );
NOR2_X1 U889 ( .A1(KEYINPUT41), .A2(n1232), .ZN(n1231) );
NOR3_X1 U890 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(n1232) );
NOR2_X1 U891 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
XNOR2_X1 U892 ( .A(n1238), .B(n1190), .ZN(n1237) );
NOR3_X1 U893 ( .A1(G125), .A2(n1190), .A3(n1238), .ZN(n1234) );
NOR2_X1 U894 ( .A1(n1137), .A2(G952), .ZN(n1156) );
XNOR2_X1 U895 ( .A(G146), .B(n1206), .ZN(G48) );
NAND3_X1 U896 ( .A1(n1239), .A2(n1217), .A3(n1240), .ZN(n1206) );
INV_X1 U897 ( .A(n1064), .ZN(n1239) );
XNOR2_X1 U898 ( .A(G143), .B(n1131), .ZN(G45) );
NAND3_X1 U899 ( .A1(n1217), .A2(n1241), .A3(n1242), .ZN(n1131) );
NOR3_X1 U900 ( .A1(n1243), .A2(n1115), .A3(n1077), .ZN(n1242) );
XOR2_X1 U901 ( .A(n1244), .B(n1245), .Z(G42) );
NAND2_X1 U902 ( .A1(KEYINPUT30), .A2(G140), .ZN(n1245) );
NAND2_X1 U903 ( .A1(n1218), .A2(n1058), .ZN(n1244) );
AND4_X1 U904 ( .A1(n1217), .A2(n1087), .A3(n1064), .A4(n1065), .ZN(n1218) );
XNOR2_X1 U905 ( .A(G137), .B(n1246), .ZN(G39) );
NAND3_X1 U906 ( .A1(n1216), .A2(n1060), .A3(n1247), .ZN(n1246) );
NOR3_X1 U907 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1247) );
NOR2_X1 U908 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
INV_X1 U909 ( .A(KEYINPUT49), .ZN(n1252) );
NOR2_X1 U910 ( .A1(n1094), .A2(n1253), .ZN(n1251) );
INV_X1 U911 ( .A(n1254), .ZN(n1094) );
NOR2_X1 U912 ( .A1(KEYINPUT49), .A2(n1217), .ZN(n1249) );
NAND2_X1 U913 ( .A1(n1255), .A2(n1256), .ZN(G36) );
NAND2_X1 U914 ( .A1(G134), .A2(n1207), .ZN(n1256) );
XOR2_X1 U915 ( .A(KEYINPUT34), .B(n1257), .Z(n1255) );
NOR2_X1 U916 ( .A1(G134), .A2(n1207), .ZN(n1257) );
NAND4_X1 U917 ( .A1(n1058), .A2(n1217), .A3(n1241), .A4(n1075), .ZN(n1207) );
XNOR2_X1 U918 ( .A(G131), .B(n1212), .ZN(G33) );
NAND4_X1 U919 ( .A1(n1058), .A2(n1217), .A3(n1241), .A4(n1087), .ZN(n1212) );
INV_X1 U920 ( .A(n1248), .ZN(n1058) );
NAND2_X1 U921 ( .A1(n1080), .A2(n1258), .ZN(n1248) );
XNOR2_X1 U922 ( .A(G128), .B(n1211), .ZN(G30) );
NAND4_X1 U923 ( .A1(n1217), .A2(n1216), .A3(n1075), .A4(n1259), .ZN(n1211) );
AND2_X1 U924 ( .A1(n1254), .A2(n1253), .ZN(n1217) );
XNOR2_X1 U925 ( .A(G101), .B(n1219), .ZN(G3) );
NAND4_X1 U926 ( .A1(n1241), .A2(n1060), .A3(n1260), .A4(n1254), .ZN(n1219) );
XNOR2_X1 U927 ( .A(G125), .B(n1210), .ZN(G27) );
NAND4_X1 U928 ( .A1(n1240), .A2(n1059), .A3(n1064), .A4(n1253), .ZN(n1210) );
NAND2_X1 U929 ( .A1(n1261), .A2(n1095), .ZN(n1253) );
NAND4_X1 U930 ( .A1(G953), .A2(G902), .A3(n1262), .A4(n1140), .ZN(n1261) );
INV_X1 U931 ( .A(G900), .ZN(n1140) );
NOR3_X1 U932 ( .A1(n1077), .A2(n1067), .A3(n1088), .ZN(n1240) );
INV_X1 U933 ( .A(n1259), .ZN(n1077) );
XOR2_X1 U934 ( .A(n1228), .B(n1263), .Z(G24) );
NOR2_X1 U935 ( .A1(G122), .A2(KEYINPUT5), .ZN(n1263) );
NAND4_X1 U936 ( .A1(n1064), .A2(n1264), .A3(n1067), .A4(n1265), .ZN(n1228) );
NOR2_X1 U937 ( .A1(n1266), .A2(n1243), .ZN(n1265) );
XNOR2_X1 U938 ( .A(G119), .B(n1227), .ZN(G21) );
NAND3_X1 U939 ( .A1(n1267), .A2(n1060), .A3(n1216), .ZN(n1227) );
NOR2_X1 U940 ( .A1(n1064), .A2(n1067), .ZN(n1216) );
INV_X1 U941 ( .A(n1065), .ZN(n1067) );
XNOR2_X1 U942 ( .A(G116), .B(n1225), .ZN(G18) );
NAND3_X1 U943 ( .A1(n1267), .A2(n1075), .A3(n1241), .ZN(n1225) );
NOR2_X1 U944 ( .A1(n1268), .A2(n1115), .ZN(n1075) );
INV_X1 U945 ( .A(n1264), .ZN(n1115) );
INV_X1 U946 ( .A(n1266), .ZN(n1267) );
XNOR2_X1 U947 ( .A(G113), .B(n1269), .ZN(G15) );
NOR2_X1 U948 ( .A1(n1223), .A2(KEYINPUT54), .ZN(n1269) );
NOR3_X1 U949 ( .A1(n1088), .A2(n1266), .A3(n1062), .ZN(n1223) );
INV_X1 U950 ( .A(n1241), .ZN(n1062) );
NOR2_X1 U951 ( .A1(n1064), .A2(n1065), .ZN(n1241) );
NAND2_X1 U952 ( .A1(n1059), .A2(n1260), .ZN(n1266) );
NOR2_X1 U953 ( .A1(n1270), .A2(n1092), .ZN(n1059) );
INV_X1 U954 ( .A(n1093), .ZN(n1270) );
INV_X1 U955 ( .A(n1087), .ZN(n1088) );
NOR2_X1 U956 ( .A1(n1243), .A2(n1264), .ZN(n1087) );
XOR2_X1 U957 ( .A(G110), .B(n1222), .Z(G12) );
AND3_X1 U958 ( .A1(n1226), .A2(n1065), .A3(n1060), .ZN(n1222) );
NOR2_X1 U959 ( .A1(n1264), .A2(n1268), .ZN(n1060) );
INV_X1 U960 ( .A(n1243), .ZN(n1268) );
XNOR2_X1 U961 ( .A(n1271), .B(n1113), .ZN(n1243) );
NOR2_X1 U962 ( .A1(n1172), .A2(G902), .ZN(n1113) );
XOR2_X1 U963 ( .A(n1272), .B(n1273), .Z(n1172) );
XOR2_X1 U964 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U965 ( .A(n1276), .B(n1277), .ZN(n1272) );
NAND2_X1 U966 ( .A1(KEYINPUT55), .A2(n1278), .ZN(n1277) );
NAND2_X1 U967 ( .A1(KEYINPUT20), .A2(n1279), .ZN(n1276) );
XOR2_X1 U968 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U969 ( .A(n1282), .B(n1283), .Z(n1281) );
NAND2_X1 U970 ( .A1(G214), .A2(n1284), .ZN(n1282) );
XOR2_X1 U971 ( .A(n1285), .B(n1286), .Z(n1280) );
XNOR2_X1 U972 ( .A(n1287), .B(G125), .ZN(n1286) );
INV_X1 U973 ( .A(G131), .ZN(n1287) );
NAND2_X1 U974 ( .A1(KEYINPUT4), .A2(n1288), .ZN(n1285) );
NAND2_X1 U975 ( .A1(KEYINPUT59), .A2(n1112), .ZN(n1271) );
INV_X1 U976 ( .A(G475), .ZN(n1112) );
XNOR2_X1 U977 ( .A(n1289), .B(G478), .ZN(n1264) );
NAND2_X1 U978 ( .A1(n1166), .A2(n1290), .ZN(n1289) );
XOR2_X1 U979 ( .A(n1291), .B(n1292), .Z(n1166) );
XOR2_X1 U980 ( .A(n1293), .B(n1294), .Z(n1292) );
NOR2_X1 U981 ( .A1(G128), .A2(KEYINPUT58), .ZN(n1294) );
NOR3_X1 U982 ( .A1(n1162), .A2(G953), .A3(n1295), .ZN(n1293) );
XNOR2_X1 U983 ( .A(G234), .B(KEYINPUT21), .ZN(n1295) );
INV_X1 U984 ( .A(G217), .ZN(n1162) );
XOR2_X1 U985 ( .A(n1296), .B(n1297), .Z(n1291) );
NOR2_X1 U986 ( .A1(KEYINPUT45), .A2(n1298), .ZN(n1297) );
XOR2_X1 U987 ( .A(n1299), .B(n1275), .Z(n1298) );
XOR2_X1 U988 ( .A(n1300), .B(G107), .Z(n1299) );
NAND2_X1 U989 ( .A1(KEYINPUT14), .A2(n1301), .ZN(n1300) );
XNOR2_X1 U990 ( .A(KEYINPUT46), .B(n1302), .ZN(n1301) );
INV_X1 U991 ( .A(G116), .ZN(n1302) );
XNOR2_X1 U992 ( .A(G134), .B(G143), .ZN(n1296) );
NAND2_X1 U993 ( .A1(n1125), .A2(n1123), .ZN(n1065) );
NAND3_X1 U994 ( .A1(n1303), .A2(n1290), .A3(n1158), .ZN(n1123) );
NAND2_X1 U995 ( .A1(G217), .A2(n1304), .ZN(n1303) );
NAND3_X1 U996 ( .A1(n1305), .A2(n1304), .A3(G217), .ZN(n1125) );
NAND2_X1 U997 ( .A1(n1158), .A2(n1290), .ZN(n1305) );
XNOR2_X1 U998 ( .A(n1306), .B(n1307), .ZN(n1158) );
XOR2_X1 U999 ( .A(n1308), .B(n1309), .Z(n1307) );
XNOR2_X1 U1000 ( .A(n1310), .B(n1311), .ZN(n1309) );
NOR4_X1 U1001 ( .A1(KEYINPUT8), .A2(G953), .A3(n1312), .A4(n1313), .ZN(n1311) );
INV_X1 U1002 ( .A(G234), .ZN(n1312) );
NAND2_X1 U1003 ( .A1(KEYINPUT47), .A2(n1314), .ZN(n1310) );
XNOR2_X1 U1004 ( .A(G119), .B(n1315), .ZN(n1314) );
NAND2_X1 U1005 ( .A1(KEYINPUT35), .A2(n1316), .ZN(n1315) );
INV_X1 U1006 ( .A(G128), .ZN(n1316) );
XOR2_X1 U1007 ( .A(n1317), .B(n1318), .Z(n1306) );
XOR2_X1 U1008 ( .A(KEYINPUT22), .B(G146), .Z(n1318) );
XNOR2_X1 U1009 ( .A(G137), .B(G125), .ZN(n1317) );
AND3_X1 U1010 ( .A1(n1254), .A2(n1064), .A3(n1260), .ZN(n1226) );
AND2_X1 U1011 ( .A1(n1259), .A2(n1319), .ZN(n1260) );
NAND2_X1 U1012 ( .A1(n1095), .A2(n1320), .ZN(n1319) );
NAND4_X1 U1013 ( .A1(G953), .A2(G902), .A3(n1262), .A4(n1148), .ZN(n1320) );
INV_X1 U1014 ( .A(G898), .ZN(n1148) );
NAND3_X1 U1015 ( .A1(n1053), .A2(n1262), .A3(G952), .ZN(n1095) );
NAND2_X1 U1016 ( .A1(G237), .A2(G234), .ZN(n1262) );
XOR2_X1 U1017 ( .A(G953), .B(KEYINPUT32), .Z(n1053) );
NOR2_X1 U1018 ( .A1(n1080), .A2(n1079), .ZN(n1259) );
INV_X1 U1019 ( .A(n1258), .ZN(n1079) );
NAND2_X1 U1020 ( .A1(G214), .A2(n1321), .ZN(n1258) );
XOR2_X1 U1021 ( .A(n1124), .B(n1120), .Z(n1080) );
AND2_X1 U1022 ( .A1(G210), .A2(n1321), .ZN(n1120) );
NAND2_X1 U1023 ( .A1(n1322), .A2(n1290), .ZN(n1321) );
INV_X1 U1024 ( .A(G237), .ZN(n1322) );
NAND2_X1 U1025 ( .A1(n1323), .A2(n1290), .ZN(n1124) );
XOR2_X1 U1026 ( .A(n1230), .B(n1324), .Z(n1323) );
NOR4_X1 U1027 ( .A1(n1325), .A2(n1326), .A3(KEYINPUT23), .A4(n1233), .ZN(n1324) );
AND3_X1 U1028 ( .A1(n1238), .A2(n1236), .A3(n1190), .ZN(n1233) );
NOR3_X1 U1029 ( .A1(n1238), .A2(n1327), .A3(n1328), .ZN(n1326) );
NOR2_X1 U1030 ( .A1(G125), .A2(n1329), .ZN(n1328) );
AND2_X1 U1031 ( .A1(n1238), .A2(n1327), .ZN(n1325) );
AND2_X1 U1032 ( .A1(n1330), .A2(n1329), .ZN(n1327) );
INV_X1 U1033 ( .A(n1190), .ZN(n1329) );
XNOR2_X1 U1034 ( .A(KEYINPUT60), .B(n1236), .ZN(n1330) );
INV_X1 U1035 ( .A(G125), .ZN(n1236) );
NAND2_X1 U1036 ( .A1(G224), .A2(n1137), .ZN(n1238) );
AND2_X1 U1037 ( .A1(n1331), .A2(n1332), .ZN(n1230) );
NAND2_X1 U1038 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
XNOR2_X1 U1039 ( .A(n1151), .B(n1335), .ZN(n1333) );
XOR2_X1 U1040 ( .A(n1336), .B(KEYINPUT7), .Z(n1331) );
NAND2_X1 U1041 ( .A1(n1153), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1042 ( .A(n1335), .B(n1151), .Z(n1337) );
XOR2_X1 U1043 ( .A(n1338), .B(n1339), .Z(n1151) );
NOR2_X1 U1044 ( .A1(KEYINPUT44), .A2(n1340), .ZN(n1339) );
NAND2_X1 U1045 ( .A1(KEYINPUT12), .A2(n1152), .ZN(n1335) );
XOR2_X1 U1046 ( .A(n1341), .B(n1342), .Z(n1152) );
NOR2_X1 U1047 ( .A1(G107), .A2(KEYINPUT16), .ZN(n1342) );
XNOR2_X1 U1048 ( .A(G101), .B(G104), .ZN(n1341) );
INV_X1 U1049 ( .A(n1334), .ZN(n1153) );
XOR2_X1 U1050 ( .A(G110), .B(n1275), .Z(n1334) );
XOR2_X1 U1051 ( .A(G122), .B(KEYINPUT51), .Z(n1275) );
XOR2_X1 U1052 ( .A(G472), .B(n1343), .Z(n1064) );
NOR2_X1 U1053 ( .A1(KEYINPUT17), .A2(n1344), .ZN(n1343) );
XOR2_X1 U1054 ( .A(KEYINPUT63), .B(n1118), .Z(n1344) );
AND2_X1 U1055 ( .A1(n1345), .A2(n1290), .ZN(n1118) );
XOR2_X1 U1056 ( .A(n1346), .B(n1347), .Z(n1345) );
XOR2_X1 U1057 ( .A(KEYINPUT38), .B(n1348), .Z(n1347) );
NOR2_X1 U1058 ( .A1(n1180), .A2(n1349), .ZN(n1348) );
XOR2_X1 U1059 ( .A(KEYINPUT10), .B(n1179), .Z(n1349) );
NOR2_X1 U1060 ( .A1(n1350), .A2(G101), .ZN(n1179) );
AND2_X1 U1061 ( .A1(G210), .A2(n1284), .ZN(n1350) );
AND3_X1 U1062 ( .A1(G210), .A2(n1284), .A3(G101), .ZN(n1180) );
NOR2_X1 U1063 ( .A1(G953), .A2(G237), .ZN(n1284) );
XNOR2_X1 U1064 ( .A(n1191), .B(n1190), .ZN(n1346) );
XOR2_X1 U1065 ( .A(G128), .B(n1351), .Z(n1190) );
NOR2_X1 U1066 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
NOR3_X1 U1067 ( .A1(KEYINPUT24), .A2(G146), .A3(n1354), .ZN(n1353) );
NOR2_X1 U1068 ( .A1(n1283), .A2(n1355), .ZN(n1352) );
INV_X1 U1069 ( .A(KEYINPUT24), .ZN(n1355) );
XNOR2_X1 U1070 ( .A(n1356), .B(n1357), .ZN(n1191) );
XNOR2_X1 U1071 ( .A(KEYINPUT50), .B(n1340), .ZN(n1357) );
INV_X1 U1072 ( .A(G119), .ZN(n1340) );
XOR2_X1 U1073 ( .A(n1338), .B(n1197), .Z(n1356) );
XNOR2_X1 U1074 ( .A(G116), .B(n1274), .ZN(n1338) );
XOR2_X1 U1075 ( .A(G113), .B(KEYINPUT2), .Z(n1274) );
NOR2_X1 U1076 ( .A1(n1093), .A2(n1092), .ZN(n1254) );
NOR2_X1 U1077 ( .A1(n1313), .A2(n1161), .ZN(n1092) );
INV_X1 U1078 ( .A(n1304), .ZN(n1161) );
NAND2_X1 U1079 ( .A1(n1358), .A2(G234), .ZN(n1304) );
XNOR2_X1 U1080 ( .A(G902), .B(KEYINPUT27), .ZN(n1358) );
INV_X1 U1081 ( .A(G221), .ZN(n1313) );
XOR2_X1 U1082 ( .A(n1359), .B(n1105), .Z(n1093) );
INV_X1 U1083 ( .A(G469), .ZN(n1105) );
NAND2_X1 U1084 ( .A1(KEYINPUT57), .A2(n1111), .ZN(n1359) );
NAND2_X1 U1085 ( .A1(n1360), .A2(n1290), .ZN(n1111) );
INV_X1 U1086 ( .A(G902), .ZN(n1290) );
XOR2_X1 U1087 ( .A(n1361), .B(n1362), .Z(n1360) );
XNOR2_X1 U1088 ( .A(n1195), .B(n1201), .ZN(n1362) );
XOR2_X1 U1089 ( .A(n1308), .B(n1363), .Z(n1201) );
NOR2_X1 U1090 ( .A1(n1139), .A2(n1364), .ZN(n1363) );
XNOR2_X1 U1091 ( .A(KEYINPUT11), .B(n1137), .ZN(n1364) );
INV_X1 U1092 ( .A(G953), .ZN(n1137) );
INV_X1 U1093 ( .A(G227), .ZN(n1139) );
XNOR2_X1 U1094 ( .A(G110), .B(n1288), .ZN(n1308) );
INV_X1 U1095 ( .A(G140), .ZN(n1288) );
XOR2_X1 U1096 ( .A(n1365), .B(n1366), .Z(n1195) );
XNOR2_X1 U1097 ( .A(G107), .B(n1278), .ZN(n1366) );
INV_X1 U1098 ( .A(G104), .ZN(n1278) );
NAND2_X1 U1099 ( .A1(KEYINPUT28), .A2(G101), .ZN(n1365) );
XNOR2_X1 U1100 ( .A(n1367), .B(n1197), .ZN(n1361) );
XOR2_X1 U1101 ( .A(G131), .B(n1368), .Z(n1197) );
XNOR2_X1 U1102 ( .A(n1369), .B(G134), .ZN(n1368) );
INV_X1 U1103 ( .A(G137), .ZN(n1369) );
NAND2_X1 U1104 ( .A1(n1370), .A2(KEYINPUT6), .ZN(n1367) );
XOR2_X1 U1105 ( .A(n1196), .B(KEYINPUT29), .Z(n1370) );
XNOR2_X1 U1106 ( .A(G128), .B(n1283), .ZN(n1196) );
XNOR2_X1 U1107 ( .A(n1354), .B(G146), .ZN(n1283) );
INV_X1 U1108 ( .A(G143), .ZN(n1354) );
endmodule


